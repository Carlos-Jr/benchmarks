module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175,
    n176, n177, n178, n179, n180, n181, n182,
    n183, n184, n185, n186, n187, n188, n189,
    n190, n191, n192, n193, n194, n195, n196,
    n197, n198, n199, n200, n201, n202, n203,
    n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n266, n267,
    n268, n269, n270, n271, n272, n273, n274,
    n275, n276, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n322, n323, n324;
  assign n92 = ~pi9  & ~pi10 ;
  assign n93 = pi11  & ~n92;
  assign n94 = ~pi12  & ~n93;
  assign n95 = ~pi13  & n94;
  assign n96 = pi14  & ~n95;
  assign n97 = pi15  & n96;
  assign n98 = ~pi16  & ~n97;
  assign n99 = pi17  & ~n98;
  assign n100 = ~pi18  & ~n99;
  assign n101 = pi19  & ~n100;
  assign n102 = pi20  & n101;
  assign n103 = ~pi21  & ~n102;
  assign n104 = ~pi22  & n103;
  assign n105 = pi23  & ~n104;
  assign n106 = pi24  & n105;
  assign n107 = pi25  & n106;
  assign n108 = ~pi26  & ~n107;
  assign n109 = pi27  & ~n108;
  assign n110 = pi28  & pi29 ;
  assign n111 = n109 & n110;
  assign n112 = pi24  & ~n105;
  assign n113 = ~pi24  & n105;
  assign n114 = ~n112 & ~n113;
  assign n115 = ~pi23  & n104;
  assign n116 = ~n105 & ~n115;
  assign n117 = pi25  & ~n106;
  assign n118 = ~pi25  & n106;
  assign n119 = ~n117 & ~n118;
  assign n120 = pi22  & ~n103;
  assign n121 = ~n104 & ~n120;
  assign n122 = pi21  & n102;
  assign n123 = ~n103 & ~n122;
  assign n124 = ~pi19  & n100;
  assign n125 = ~n101 & ~n124;
  assign n126 = pi18  & n99;
  assign n127 = ~n100 & ~n126;
  assign n128 = pi20  & ~n101;
  assign n129 = ~pi20  & n101;
  assign n130 = ~n128 & ~n129;
  assign n131 = ~pi17  & n98;
  assign n132 = ~n99 & ~n131;
  assign n133 = pi16  & n97;
  assign n134 = ~n98 & ~n133;
  assign n135 = ~pi11  & n92;
  assign n136 = ~n93 & ~n135;
  assign n137 = pi15  & ~n96;
  assign n138 = ~pi15  & n96;
  assign n139 = ~n137 & ~n138;
  assign n140 = ~pi14  & n95;
  assign n141 = ~n96 & ~n140;
  assign n142 = pi13  & ~n94;
  assign n143 = ~n95 & ~n142;
  assign n144 = pi12  & n93;
  assign n145 = ~n94 & ~n144;
  assign n146 = pi26  & n107;
  assign n147 = ~pi27  & ~n146;
  assign n148 = pi0  & pi1 ;
  assign n149 = pi2  & pi3 ;
  assign n150 = pi4  & pi5 ;
  assign n151 = pi6  & pi7 ;
  assign n152 = pi8  & pi28 ;
  assign n153 = pi29  & n152;
  assign n154 = n150 & n151;
  assign n155 = n148 & n149;
  assign n156 = n92 & n155;
  assign n157 = n153 & n154;
  assign n158 = n156 & n157;
  assign n159 = n136 & n158;
  assign n160 = ~n145 & n159;
  assign n161 = ~n143 & n160;
  assign n162 = n141 & n161;
  assign n163 = ~n139 & n162;
  assign n164 = ~n134 & n163;
  assign n165 = n132 & n164;
  assign n166 = ~n127 & n165;
  assign n167 = n125 & n166;
  assign n168 = ~n130 & n167;
  assign n169 = ~n123 & n168;
  assign n170 = ~n121 & n169;
  assign n171 = n116 & n170;
  assign n172 = ~n114 & n171;
  assign n173 = ~n119 & n172;
  assign n174 = ~n109 & ~n147;
  assign n175 = n173 & n174;
  assign n176 = ~n111 & ~n175;
  assign n177 = ~pi1  & ~pi2 ;
  assign n178 = ~pi3  & ~pi4 ;
  assign n179 = ~pi5  & ~pi6 ;
  assign n180 = ~pi7  & ~pi8 ;
  assign n181 = pi9  & ~pi10 ;
  assign n182 = n180 & n181;
  assign n183 = n178 & n179;
  assign n184 = n177 & n183;
  assign n185 = n182 & n184;
  assign n186 = ~n136 & n185;
  assign n187 = n145 & n186;
  assign n188 = n143 & n187;
  assign n189 = ~n141 & n188;
  assign n190 = n139 & n189;
  assign n191 = n134 & n190;
  assign n192 = ~n132 & n191;
  assign n193 = n127 & n192;
  assign n194 = ~n125 & n193;
  assign n195 = n130 & n194;
  assign n196 = n123 & n195;
  assign n197 = n121 & n196;
  assign n198 = ~n116 & n197;
  assign n199 = n114 & n198;
  assign n200 = ~n108 & n119;
  assign n201 = ~n146 & n200;
  assign n202 = n199 & n201;
  assign n203 = n111 & ~n202;
  assign po0  = n176 | n203;
  assign n205 = ~pi39  & ~pi40 ;
  assign n206 = pi41  & ~n205;
  assign n207 = ~pi42  & ~n206;
  assign n208 = ~pi43  & n207;
  assign n209 = pi44  & ~n208;
  assign n210 = pi45  & n209;
  assign n211 = ~pi46  & ~n210;
  assign n212 = pi47  & ~n211;
  assign n213 = ~pi48  & ~n212;
  assign n214 = pi49  & ~n213;
  assign n215 = pi50  & n214;
  assign n216 = ~pi51  & ~n215;
  assign n217 = ~pi52  & n216;
  assign n218 = pi53  & ~n217;
  assign n219 = pi54  & n218;
  assign n220 = pi55  & n219;
  assign n221 = ~pi56  & ~n220;
  assign n222 = pi57  & ~n221;
  assign n223 = pi58  & pi59 ;
  assign n224 = n222 & n223;
  assign n225 = pi0  & ~n224;
  assign n226 = pi54  & ~n218;
  assign n227 = ~pi54  & n218;
  assign n228 = ~n226 & ~n227;
  assign n229 = ~pi53  & n217;
  assign n230 = ~n218 & ~n229;
  assign n231 = pi55  & ~n219;
  assign n232 = ~pi55  & n219;
  assign n233 = ~n231 & ~n232;
  assign n234 = pi52  & ~n216;
  assign n235 = ~n217 & ~n234;
  assign n236 = pi51  & n215;
  assign n237 = ~n216 & ~n236;
  assign n238 = ~pi49  & n213;
  assign n239 = ~n214 & ~n238;
  assign n240 = pi48  & n212;
  assign n241 = ~n213 & ~n240;
  assign n242 = pi50  & ~n214;
  assign n243 = ~pi50  & n214;
  assign n244 = ~n242 & ~n243;
  assign n245 = ~pi47  & n211;
  assign n246 = ~n212 & ~n245;
  assign n247 = pi46  & n210;
  assign n248 = ~n211 & ~n247;
  assign n249 = ~pi41  & n205;
  assign n250 = ~n206 & ~n249;
  assign n251 = pi45  & ~n209;
  assign n252 = ~pi45  & n209;
  assign n253 = ~n251 & ~n252;
  assign n254 = ~pi44  & n208;
  assign n255 = ~n209 & ~n254;
  assign n256 = pi43  & ~n207;
  assign n257 = ~n208 & ~n256;
  assign n258 = pi42  & n206;
  assign n259 = ~n207 & ~n258;
  assign n260 = pi56  & n220;
  assign n261 = ~pi57  & ~n260;
  assign n262 = pi30  & pi31 ;
  assign n263 = pi32  & pi33 ;
  assign n264 = pi34  & pi35 ;
  assign n265 = pi36  & pi37 ;
  assign n266 = pi38  & n265;
  assign n267 = n263 & n264;
  assign n268 = n205 & n262;
  assign n269 = n223 & n268;
  assign n270 = n266 & n267;
  assign n271 = n269 & n270;
  assign n272 = n250 & n271;
  assign n273 = ~n259 & n272;
  assign n274 = ~n257 & n273;
  assign n275 = n255 & n274;
  assign n276 = ~n253 & n275;
  assign n277 = ~n248 & n276;
  assign n278 = n246 & n277;
  assign n279 = ~n241 & n278;
  assign n280 = n239 & n279;
  assign n281 = ~n244 & n280;
  assign n282 = ~n237 & n281;
  assign n283 = ~n235 & n282;
  assign n284 = n230 & n283;
  assign n285 = ~n228 & n284;
  assign n286 = ~n233 & n285;
  assign n287 = ~n222 & ~n261;
  assign n288 = n286 & n287;
  assign n289 = ~pi31  & ~pi32 ;
  assign n290 = ~pi33  & ~pi34 ;
  assign n291 = ~pi35  & ~pi36 ;
  assign n292 = ~pi37  & ~pi38 ;
  assign n293 = pi39  & ~pi40 ;
  assign n294 = n292 & n293;
  assign n295 = n290 & n291;
  assign n296 = n289 & n295;
  assign n297 = n294 & n296;
  assign n298 = ~n250 & n297;
  assign n299 = n259 & n298;
  assign n300 = n257 & n299;
  assign n301 = ~n255 & n300;
  assign n302 = n253 & n301;
  assign n303 = n248 & n302;
  assign n304 = ~n246 & n303;
  assign n305 = n241 & n304;
  assign n306 = ~n239 & n305;
  assign n307 = n244 & n306;
  assign n308 = n237 & n307;
  assign n309 = n235 & n308;
  assign n310 = ~n230 & n309;
  assign n311 = n228 & n310;
  assign n312 = ~n221 & n233;
  assign n313 = ~n260 & n312;
  assign n314 = n311 & n313;
  assign n315 = ~pi0  & ~pi30 ;
  assign n316 = n314 & n315;
  assign n317 = n224 & ~n316;
  assign n318 = ~n288 & ~n317;
  assign n319 = ~n176 & ~n225;
  assign n320 = ~n318 & n319;
  assign po1  = ~n203 & ~n320;
  assign n322 = pi0  & pi30 ;
  assign n323 = n314 & ~n322;
  assign n324 = n224 & ~n323;
  assign po2  = ~po0  & n324;
  assign po3  = 1'b0;
  assign po4  = 1'b0;
  assign po5  = 1'b0;
  assign po6  = 1'b0;
  assign po7  = 1'b0;
  assign po8  = 1'b0;
  assign po9  = 1'b0;
  assign po10  = 1'b0;
  assign po11  = 1'b0;
  assign po12  = 1'b0;
  assign po13  = 1'b0;
  assign po14  = 1'b0;
  assign po15  = 1'b0;
  assign po16  = 1'b0;
  assign po17  = 1'b0;
  assign po18  = 1'b0;
  assign po19  = 1'b0;
  assign po20  = 1'b0;
  assign po21  = 1'b0;
  assign po22  = 1'b0;
  assign po23  = 1'b0;
  assign po24  = 1'b0;
  assign po25  = 1'b0;
  assign po26  = 1'b0;
  assign po27  = 1'b0;
  assign po28  = 1'b0;
  assign po29  = 1'b0;
endmodule
