module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n404,
    n405, n406, n407, n408, n409, n411, n412,
    n413, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575,
    n576, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n660, n661;
  assign n22 = ~pi3  & ~pi5 ;
  assign n23 = ~pi1  & pi9 ;
  assign n24 = ~pi0  & pi9 ;
  assign n25 = pi1  & ~n24;
  assign n26 = ~n23 & ~n25;
  assign n27 = n22 & n26;
  assign n28 = pi1  & ~pi9 ;
  assign n29 = pi0  & ~pi9 ;
  assign n30 = ~pi1  & ~n29;
  assign n31 = ~pi7  & ~n30;
  assign n32 = ~n28 & n31;
  assign n33 = ~n27 & ~n32;
  assign n34 = ~pi2  & ~n33;
  assign n35 = ~pi2  & ~pi3 ;
  assign n36 = pi9  & ~n35;
  assign n37 = pi0  & pi3 ;
  assign n38 = ~n36 & ~n37;
  assign n39 = ~pi1  & ~n38;
  assign n40 = pi1  & ~pi3 ;
  assign n41 = ~pi2  & ~pi5 ;
  assign n42 = ~pi0  & ~n41;
  assign n43 = pi1  & pi2 ;
  assign n44 = ~n42 & ~n43;
  assign n45 = ~pi9  & ~n44;
  assign n46 = ~n40 & ~n45;
  assign n47 = ~n39 & n46;
  assign n48 = ~pi7  & ~n47;
  assign n49 = ~n34 & ~n48;
  assign n50 = ~pi8  & ~n49;
  assign n51 = ~pi7  & pi9 ;
  assign n52 = ~pi5  & pi8 ;
  assign n53 = pi7  & n52;
  assign n54 = ~n51 & ~n53;
  assign n55 = pi1  & ~n54;
  assign n56 = pi1  & ~pi7 ;
  assign n57 = ~pi5  & ~pi9 ;
  assign n58 = ~n56 & n57;
  assign n59 = ~n55 & ~n58;
  assign n60 = pi0  & ~pi2 ;
  assign n61 = ~n59 & n60;
  assign n62 = ~pi0  & ~pi9 ;
  assign n63 = ~pi1  & pi2 ;
  assign n64 = n62 & n63;
  assign n65 = n53 & n64;
  assign n66 = ~n61 & ~n65;
  assign n67 = ~pi3  & ~n66;
  assign n68 = ~n50 & ~n67;
  assign n69 = ~pi6  & ~n68;
  assign n70 = ~pi1  & ~pi2 ;
  assign n71 = ~pi0  & n70;
  assign n72 = ~pi3  & ~pi8 ;
  assign n73 = ~pi1  & ~pi9 ;
  assign n74 = pi1  & pi9 ;
  assign n75 = ~n73 & ~n74;
  assign n76 = n72 & ~n75;
  assign n77 = n71 & n76;
  assign n78 = ~pi1  & ~n24;
  assign n79 = ~pi8  & ~n78;
  assign n80 = n29 & n63;
  assign n81 = ~n79 & ~n80;
  assign n82 = ~pi5  & ~n81;
  assign n83 = pi5  & pi6 ;
  assign n84 = pi6  & pi9 ;
  assign n85 = n71 & n84;
  assign n86 = pi0  & pi9 ;
  assign n87 = ~n62 & ~n86;
  assign n88 = pi5  & ~n87;
  assign n89 = n43 & n88;
  assign n90 = ~n85 & ~n89;
  assign n91 = ~n83 & n90;
  assign n92 = pi8  & ~n91;
  assign n93 = ~n82 & ~n92;
  assign n94 = pi3  & ~n93;
  assign n95 = ~pi2  & ~n29;
  assign n96 = pi6  & ~n95;
  assign n97 = pi1  & ~n87;
  assign n98 = n35 & n97;
  assign n99 = ~n96 & ~n98;
  assign n100 = pi5  & ~n99;
  assign n101 = pi2  & ~pi9 ;
  assign n102 = ~pi2  & pi9 ;
  assign n103 = ~n101 & ~n102;
  assign n104 = ~pi0  & ~pi3 ;
  assign n105 = pi6  & ~n73;
  assign n106 = n104 & n105;
  assign n107 = n103 & n106;
  assign n108 = ~n100 & ~n107;
  assign n109 = pi8  & ~n108;
  assign n110 = pi1  & ~pi8 ;
  assign n111 = pi2  & ~pi3 ;
  assign n112 = n23 & n111;
  assign n113 = ~n110 & ~n112;
  assign n114 = ~pi0  & ~n113;
  assign n115 = pi2  & pi9 ;
  assign n116 = pi3  & ~pi6 ;
  assign n117 = pi2  & pi3 ;
  assign n118 = ~n116 & ~n117;
  assign n119 = n73 & n118;
  assign n120 = ~n115 & ~n119;
  assign n121 = ~pi8  & ~n120;
  assign n122 = ~n114 & ~n121;
  assign n123 = ~pi5  & ~n122;
  assign n124 = ~n109 & ~n123;
  assign n125 = ~n94 & n124;
  assign n126 = ~n77 & n125;
  assign n127 = ~pi7  & ~n126;
  assign n128 = ~n69 & ~n127;
  assign n129 = ~pi4  & ~n128;
  assign n130 = ~pi0  & ~pi2 ;
  assign n131 = ~pi8  & ~pi9 ;
  assign n132 = ~pi6  & n131;
  assign n133 = pi4  & pi8 ;
  assign n134 = pi6  & n133;
  assign n135 = ~n132 & ~n134;
  assign n136 = pi5  & ~n135;
  assign n137 = ~pi6  & pi9 ;
  assign n138 = ~pi5  & pi6 ;
  assign n139 = ~n137 & ~n138;
  assign n140 = ~pi4  & pi9 ;
  assign n141 = ~pi8  & ~n140;
  assign n142 = ~n139 & n141;
  assign n143 = ~n136 & ~n142;
  assign n144 = ~pi1  & ~pi3 ;
  assign n145 = ~n143 & n144;
  assign n146 = ~pi7  & n145;
  assign n147 = n130 & n146;
  assign po0  = n129 | n147;
  assign n149 = pi8  & n86;
  assign n150 = ~n131 & ~n149;
  assign n151 = pi5  & ~n150;
  assign n152 = ~n60 & ~n101;
  assign n153 = n151 & n152;
  assign n154 = ~pi8  & n57;
  assign n155 = ~n52 & ~n84;
  assign n156 = pi6  & pi8 ;
  assign n157 = pi0  & ~n156;
  assign n158 = ~n29 & ~n157;
  assign n159 = ~n155 & n158;
  assign n160 = ~n154 & ~n159;
  assign n161 = pi2  & ~n160;
  assign n162 = ~n153 & ~n161;
  assign n163 = ~pi4  & ~n162;
  assign n164 = pi4  & pi9 ;
  assign n165 = pi5  & ~pi8 ;
  assign n166 = ~n133 & ~n165;
  assign n167 = ~pi6  & ~n166;
  assign n168 = ~n164 & ~n167;
  assign n169 = ~n137 & ~n168;
  assign n170 = n130 & n169;
  assign n171 = ~n163 & ~n170;
  assign n172 = ~pi1  & ~n171;
  assign n173 = ~n155 & n157;
  assign n174 = ~pi0  & pi5 ;
  assign n175 = ~pi8  & pi9 ;
  assign n176 = n174 & n175;
  assign n177 = ~n173 & ~n176;
  assign n178 = ~pi2  & ~n177;
  assign n179 = ~pi6  & ~pi8 ;
  assign n180 = pi2  & ~pi5 ;
  assign n181 = ~pi6  & ~n180;
  assign n182 = n52 & ~n60;
  assign n183 = ~n181 & n182;
  assign n184 = ~n179 & ~n183;
  assign n185 = ~pi9  & ~n184;
  assign n186 = ~n178 & ~n185;
  assign n187 = pi1  & ~n186;
  assign n188 = ~pi6  & pi8 ;
  assign n189 = n101 & n188;
  assign n190 = ~n187 & ~n189;
  assign n191 = ~pi4  & ~n190;
  assign n192 = ~n172 & ~n191;
  assign n193 = ~pi3  & ~n192;
  assign n194 = ~pi2  & pi8 ;
  assign n195 = pi0  & n194;
  assign n196 = pi0  & ~pi5 ;
  assign n197 = ~n195 & ~n196;
  assign n198 = ~n174 & n197;
  assign n199 = pi1  & ~n198;
  assign n200 = ~pi2  & ~pi8 ;
  assign n201 = ~n35 & ~n200;
  assign n202 = ~pi0  & n201;
  assign n203 = pi5  & n200;
  assign n204 = ~n52 & ~n72;
  assign n205 = pi0  & n204;
  assign n206 = ~n203 & ~n205;
  assign n207 = ~pi1  & ~n206;
  assign n208 = ~n202 & ~n207;
  assign n209 = ~n199 & n208;
  assign n210 = ~pi6  & ~n209;
  assign n211 = pi2  & n116;
  assign n212 = pi3  & ~n211;
  assign n213 = ~pi1  & ~pi8 ;
  assign n214 = ~n43 & ~n213;
  assign n215 = n212 & n214;
  assign n216 = ~pi0  & pi8 ;
  assign n217 = pi0  & pi1 ;
  assign n218 = ~pi1  & ~pi6 ;
  assign n219 = ~pi2  & ~n218;
  assign n220 = ~n217 & n219;
  assign n221 = ~n216 & n220;
  assign n222 = ~n215 & ~n221;
  assign n223 = ~pi5  & ~n222;
  assign n224 = ~pi9  & ~n223;
  assign n225 = ~n210 & n224;
  assign n226 = ~pi4  & ~n225;
  assign n227 = pi1  & pi5 ;
  assign n228 = pi3  & ~pi8 ;
  assign n229 = n70 & n228;
  assign n230 = ~n227 & ~n229;
  assign n231 = pi0  & ~n230;
  assign n232 = pi5  & ~n35;
  assign n233 = ~n231 & ~n232;
  assign n234 = pi6  & ~n233;
  assign n235 = pi3  & n43;
  assign n236 = ~pi6  & ~n165;
  assign n237 = n235 & ~n236;
  assign n238 = pi9  & ~n237;
  assign n239 = ~n234 & n238;
  assign n240 = n226 & ~n239;
  assign n241 = ~n193 & ~n240;
  assign n242 = ~pi7  & ~n241;
  assign n243 = n28 & n194;
  assign n244 = n95 & ~n217;
  assign n245 = ~pi0  & ~n43;
  assign n246 = pi2  & ~n245;
  assign n247 = ~pi8  & ~n246;
  assign n248 = ~n244 & n247;
  assign n249 = ~n243 & ~n248;
  assign n250 = pi7  & ~n249;
  assign n251 = ~n64 & ~n250;
  assign n252 = n22 & ~n251;
  assign n253 = ~pi4  & n252;
  assign n254 = ~pi6  & n253;
  assign po1  = n242 | n254;
  assign n256 = n76 & n84;
  assign n257 = ~pi3  & pi9 ;
  assign n258 = ~n73 & ~n257;
  assign n259 = pi3  & ~n175;
  assign n260 = ~pi6  & ~n259;
  assign n261 = n258 & n260;
  assign n262 = pi3  & ~n194;
  assign n263 = pi5  & ~n262;
  assign n264 = pi3  & ~n180;
  assign n265 = pi8  & ~n264;
  assign n266 = ~n263 & ~n265;
  assign n267 = pi1  & ~n266;
  assign n268 = ~pi3  & n138;
  assign n269 = n213 & n268;
  assign n270 = ~n267 & ~n269;
  assign n271 = ~pi9  & ~n270;
  assign n272 = ~pi1  & n201;
  assign n273 = pi2  & ~n188;
  assign n274 = ~n272 & ~n273;
  assign n275 = pi5  & ~n274;
  assign n276 = pi1  & pi8 ;
  assign n277 = pi6  & ~n276;
  assign n278 = ~pi9  & ~n277;
  assign n279 = ~pi2  & ~n278;
  assign n280 = ~pi8  & n23;
  assign n281 = ~n279 & ~n280;
  assign n282 = pi3  & ~n281;
  assign n283 = ~n275 & ~n282;
  assign n284 = ~n271 & n283;
  assign n285 = ~n261 & n284;
  assign n286 = ~n256 & n285;
  assign n287 = ~pi4  & ~n286;
  assign n288 = pi6  & ~pi8 ;
  assign n289 = pi8  & pi9 ;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~pi5  & ~n290;
  assign n292 = ~pi3  & pi4 ;
  assign n293 = ~n291 & n292;
  assign n294 = n70 & n293;
  assign n295 = ~n287 & ~n294;
  assign n296 = ~pi0  & ~n295;
  assign n297 = ~pi5  & n115;
  assign n298 = ~n151 & ~n297;
  assign n299 = pi1  & ~n298;
  assign n300 = ~n131 & ~n289;
  assign n301 = ~n73 & ~n300;
  assign n302 = pi2  & ~n301;
  assign n303 = ~n299 & ~n302;
  assign n304 = ~pi3  & ~n303;
  assign n305 = ~pi1  & pi8 ;
  assign n306 = n36 & n305;
  assign n307 = ~n41 & ~n229;
  assign n308 = n131 & ~n307;
  assign n309 = ~n306 & ~n308;
  assign n310 = pi0  & ~n309;
  assign n311 = ~n304 & ~n310;
  assign n312 = ~pi6  & ~n311;
  assign n313 = pi6  & ~n23;
  assign n314 = ~n28 & ~n313;
  assign n315 = pi8  & ~n314;
  assign n316 = ~n76 & ~n315;
  assign n317 = ~pi2  & ~n316;
  assign n318 = pi2  & n74;
  assign n319 = ~n305 & ~n318;
  assign n320 = pi6  & ~n319;
  assign n321 = pi2  & ~n300;
  assign n322 = ~n194 & ~n321;
  assign n323 = ~n320 & n322;
  assign n324 = pi3  & ~n323;
  assign n325 = ~n317 & ~n324;
  assign n326 = n196 & ~n325;
  assign n327 = ~n312 & ~n326;
  assign n328 = ~pi4  & ~n327;
  assign n329 = ~n296 & ~n328;
  assign n330 = ~pi7  & ~n329;
  assign n331 = ~pi5  & ~pi6 ;
  assign n332 = n29 & n213;
  assign n333 = ~n51 & ~n175;
  assign n334 = n97 & n333;
  assign n335 = ~n332 & ~n334;
  assign n336 = n331 & ~n335;
  assign n337 = ~pi4  & n336;
  assign n338 = n35 & n337;
  assign po2  = n330 | n338;
  assign n340 = pi6  & ~n35;
  assign n341 = pi3  & ~pi9 ;
  assign n342 = ~n340 & ~n341;
  assign n343 = ~pi4  & ~n342;
  assign n344 = ~pi6  & ~n289;
  assign n345 = ~n83 & ~n331;
  assign n346 = ~pi2  & ~n345;
  assign n347 = ~n344 & n346;
  assign n348 = n292 & n347;
  assign n349 = ~n343 & ~n348;
  assign n350 = ~pi1  & ~n349;
  assign n351 = ~pi6  & ~n228;
  assign n352 = pi3  & ~pi5 ;
  assign n353 = ~n351 & ~n352;
  assign n354 = pi3  & ~n353;
  assign n355 = ~pi5  & n288;
  assign n356 = n155 & ~n165;
  assign n357 = n321 & n356;
  assign n358 = ~n355 & ~n357;
  assign n359 = ~n354 & n358;
  assign n360 = pi1  & ~n359;
  assign n361 = pi2  & n138;
  assign n362 = ~n360 & ~n361;
  assign n363 = ~pi4  & ~n362;
  assign n364 = ~n350 & ~n363;
  assign n365 = ~pi0  & ~n364;
  assign n366 = n203 & n218;
  assign n367 = ~n268 & ~n366;
  assign n368 = ~pi9  & ~n367;
  assign n369 = pi2  & ~n204;
  assign n370 = pi5  & n194;
  assign n371 = ~n369 & ~n370;
  assign n372 = ~pi9  & ~n371;
  assign n373 = ~pi2  & pi3 ;
  assign n374 = n102 & n165;
  assign n375 = ~n373 & ~n374;
  assign n376 = ~n372 & n375;
  assign n377 = ~n353 & n376;
  assign n378 = pi1  & ~n377;
  assign n379 = ~n368 & ~n378;
  assign n380 = pi0  & ~n379;
  assign n381 = ~pi9  & n138;
  assign n382 = n276 & n381;
  assign n383 = ~n116 & ~n381;
  assign n384 = ~pi8  & ~n383;
  assign n385 = ~n138 & ~n211;
  assign n386 = n36 & ~n385;
  assign n387 = ~n384 & ~n386;
  assign n388 = ~pi1  & ~n387;
  assign n389 = ~n57 & ~n179;
  assign n390 = ~pi2  & ~n389;
  assign n391 = pi5  & pi9 ;
  assign n392 = ~pi6  & ~n391;
  assign n393 = pi5  & pi8 ;
  assign n394 = ~n74 & ~n393;
  assign n395 = n392 & ~n394;
  assign n396 = ~n390 & ~n395;
  assign n397 = pi3  & ~n396;
  assign n398 = ~n388 & ~n397;
  assign n399 = ~n382 & n398;
  assign n400 = ~n380 & n399;
  assign n401 = ~pi4  & ~n400;
  assign n402 = ~n365 & ~n401;
  assign po3  = ~pi7  & ~n402;
  assign n404 = ~pi4  & n246;
  assign n405 = pi3  & ~pi4 ;
  assign n406 = ~n292 & ~n405;
  assign n407 = n71 & ~n406;
  assign n408 = ~n404 & ~n407;
  assign n409 = ~pi7  & n83;
  assign po4  = ~n408 & n409;
  assign n411 = ~n71 & n405;
  assign n412 = n71 & n292;
  assign n413 = ~n411 & ~n412;
  assign po5  = n409 & ~n413;
  assign n415 = pi6  & ~n300;
  assign n416 = n103 & n415;
  assign n417 = ~pi0  & n115;
  assign n418 = ~pi9  & n213;
  assign n419 = ~n417 & ~n418;
  assign n420 = pi5  & ~n419;
  assign n421 = pi5  & n74;
  assign n422 = ~pi1  & ~pi5 ;
  assign n423 = pi2  & ~n422;
  assign n424 = ~pi6  & ~n423;
  assign n425 = ~pi9  & n424;
  assign n426 = ~n421 & ~n425;
  assign n427 = pi0  & ~n426;
  assign n428 = ~pi0  & ~n57;
  assign n429 = pi2  & n428;
  assign n430 = ~n427 & ~n429;
  assign n431 = pi8  & ~n430;
  assign n432 = ~n420 & ~n431;
  assign n433 = ~n416 & n432;
  assign n434 = ~pi7  & ~n433;
  assign n435 = pi7  & ~pi9 ;
  assign n436 = pi8  & ~n435;
  assign n437 = pi2  & ~n436;
  assign n438 = ~n28 & ~n437;
  assign n439 = n245 & ~n438;
  assign n440 = pi7  & ~n305;
  assign n441 = ~pi2  & n440;
  assign n442 = ~n150 & n441;
  assign n443 = ~n439 & ~n442;
  assign n444 = n331 & ~n443;
  assign n445 = ~n434 & ~n444;
  assign n446 = ~pi3  & ~n445;
  assign n447 = pi2  & n28;
  assign n448 = ~pi1  & ~n131;
  assign n449 = ~n28 & ~n448;
  assign n450 = pi0  & n449;
  assign n451 = ~n447 & ~n450;
  assign n452 = ~pi0  & ~pi6 ;
  assign n453 = n75 & ~n213;
  assign n454 = n452 & n453;
  assign n455 = n451 & ~n454;
  assign n456 = ~pi5  & ~n455;
  assign n457 = pi0  & n156;
  assign n458 = ~n110 & ~n457;
  assign n459 = ~pi2  & ~n458;
  assign n460 = ~pi8  & n217;
  assign n461 = ~n459 & ~n460;
  assign n462 = pi9  & ~n461;
  assign n463 = ~pi0  & ~pi8 ;
  assign n464 = ~n196 & ~n463;
  assign n465 = n28 & n464;
  assign n466 = ~n462 & ~n465;
  assign n467 = ~n456 & n466;
  assign n468 = pi3  & ~n467;
  assign n469 = n24 & ~n181;
  assign n470 = ~pi2  & pi5 ;
  assign n471 = ~n87 & n470;
  assign n472 = ~n469 & ~n471;
  assign n473 = ~pi8  & ~n472;
  assign n474 = pi2  & ~n131;
  assign n475 = ~n149 & ~n474;
  assign n476 = pi6  & ~n475;
  assign n477 = ~n473 & ~n476;
  assign n478 = pi1  & ~n477;
  assign n479 = ~pi9  & n288;
  assign n480 = n29 & ~n389;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~pi2  & ~n481;
  assign n483 = pi2  & pi8 ;
  assign n484 = n24 & n483;
  assign n485 = ~n482 & ~n484;
  assign n486 = ~pi1  & ~n485;
  assign n487 = ~n478 & ~n486;
  assign n488 = ~n468 & n487;
  assign n489 = ~pi7  & ~n488;
  assign n490 = ~n446 & ~n489;
  assign n491 = ~pi4  & ~n490;
  assign n492 = ~n83 & ~n412;
  assign n493 = ~pi7  & ~n492;
  assign po6  = ~n491 & ~n493;
  assign n495 = ~pi0  & n415;
  assign n496 = n95 & n344;
  assign n497 = ~n495 & ~n496;
  assign n498 = pi3  & ~n497;
  assign n499 = ~pi0  & n200;
  assign n500 = ~n457 & ~n499;
  assign n501 = ~pi9  & ~n500;
  assign n502 = ~pi6  & ~n72;
  assign n503 = n474 & ~n502;
  assign n504 = ~n501 & ~n503;
  assign n505 = ~n498 & n504;
  assign n506 = ~pi1  & ~n505;
  assign n507 = n373 & n479;
  assign n508 = pi0  & pi8 ;
  assign n509 = pi3  & ~n289;
  assign n510 = ~n508 & ~n509;
  assign n511 = ~pi6  & ~n510;
  assign n512 = pi8  & n257;
  assign n513 = ~n511 & ~n512;
  assign n514 = pi2  & ~n513;
  assign n515 = ~pi3  & n132;
  assign n516 = ~pi3  & pi8 ;
  assign n517 = ~n84 & ~n516;
  assign n518 = pi0  & ~n517;
  assign n519 = ~n260 & ~n415;
  assign n520 = ~n511 & n519;
  assign n521 = ~n518 & ~n520;
  assign n522 = ~pi2  & ~n521;
  assign n523 = ~n515 & ~n522;
  assign n524 = ~n514 & n523;
  assign n525 = pi1  & ~n524;
  assign n526 = ~n507 & ~n525;
  assign n527 = ~n506 & n526;
  assign n528 = ~pi5  & ~n527;
  assign n529 = ~pi2  & ~n37;
  assign n530 = ~n117 & n300;
  assign n531 = pi5  & ~n530;
  assign n532 = ~n529 & n531;
  assign n533 = ~pi8  & n101;
  assign n534 = n37 & n533;
  assign n535 = ~n532 & ~n534;
  assign n536 = ~pi1  & ~n535;
  assign n537 = pi8  & n391;
  assign n538 = n117 & n537;
  assign n539 = pi5  & n373;
  assign n540 = ~n101 & ~n264;
  assign n541 = n42 & ~n540;
  assign n542 = ~n539 & ~n541;
  assign n543 = ~pi8  & ~n542;
  assign n544 = pi0  & ~n103;
  assign n545 = ~pi9  & n174;
  assign n546 = ~n544 & ~n545;
  assign n547 = pi8  & ~n546;
  assign n548 = n115 & n165;
  assign n549 = ~n547 & ~n548;
  assign n550 = ~pi3  & ~n549;
  assign n551 = ~pi9  & n539;
  assign n552 = ~n550 & ~n551;
  assign n553 = ~n543 & n552;
  assign n554 = pi1  & ~n553;
  assign n555 = ~n538 & ~n554;
  assign n556 = ~n536 & n555;
  assign n557 = ~pi6  & ~n556;
  assign n558 = ~n528 & ~n557;
  assign n559 = ~pi7  & ~n558;
  assign n560 = ~pi0  & n483;
  assign n561 = ~n195 & ~n560;
  assign n562 = ~n499 & n561;
  assign n563 = ~pi9  & ~n562;
  assign n564 = n115 & n463;
  assign n565 = ~n563 & ~n564;
  assign n566 = ~pi1  & ~n565;
  assign n567 = n74 & n499;
  assign n568 = ~n566 & ~n567;
  assign n569 = ~pi6  & n22;
  assign n570 = ~n568 & n569;
  assign n571 = ~n32 & ~n200;
  assign n572 = n570 & n571;
  assign n573 = ~n559 & ~n572;
  assign n574 = ~pi4  & ~n573;
  assign n575 = ~pi7  & n331;
  assign n576 = n412 & n575;
  assign po7  = ~n574 & ~n576;
  assign n578 = n75 & ~n422;
  assign n579 = n111 & ~n578;
  assign n580 = ~pi2  & ~n227;
  assign n581 = ~n352 & n580;
  assign n582 = n258 & n581;
  assign n583 = ~n579 & ~n582;
  assign n584 = n26 & ~n47;
  assign n585 = n152 & n584;
  assign n586 = n583 & ~n585;
  assign n587 = ~pi8  & ~n586;
  assign n588 = n144 & n196;
  assign n589 = ~n104 & n581;
  assign n590 = ~n588 & ~n589;
  assign n591 = pi8  & ~n590;
  assign n592 = pi2  & ~n196;
  assign n593 = n267 & n592;
  assign n594 = ~n591 & ~n593;
  assign n595 = ~pi9  & ~n594;
  assign n596 = ~n22 & ~n470;
  assign n597 = pi1  & ~n596;
  assign n598 = n201 & n597;
  assign n599 = ~pi2  & ~n174;
  assign n600 = n272 & n599;
  assign n601 = ~n598 & ~n600;
  assign n602 = pi9  & ~n601;
  assign n603 = ~n595 & ~n602;
  assign n604 = ~n587 & n603;
  assign n605 = ~pi6  & ~n604;
  assign n606 = ~n289 & ~n448;
  assign n607 = pi6  & n606;
  assign n608 = ~n218 & n273;
  assign n609 = ~n448 & ~n484;
  assign n610 = n246 & n609;
  assign n611 = ~n313 & ~n610;
  assign n612 = pi0  & ~n611;
  assign n613 = ~n608 & ~n612;
  assign n614 = ~n607 & n613;
  assign n615 = n352 & ~n614;
  assign n616 = ~n605 & ~n615;
  assign n617 = ~pi7  & ~n616;
  assign n618 = ~n570 & ~n617;
  assign n619 = ~pi4  & ~n618;
  assign n620 = ~pi5  & ~pi7 ;
  assign n621 = n412 & n620;
  assign po8  = ~n619 & ~n621;
  assign n623 = n196 & n211;
  assign n624 = ~pi7  & ~n623;
  assign n625 = ~n448 & ~n624;
  assign n626 = ~pi2  & n144;
  assign n627 = ~pi7  & ~n626;
  assign n628 = pi0  & ~n627;
  assign n629 = pi4  & ~n626;
  assign n630 = ~pi3  & ~n57;
  assign n631 = n216 & ~n517;
  assign n632 = ~n630 & ~n631;
  assign n633 = ~pi2  & ~n632;
  assign n634 = ~pi6  & ~n537;
  assign n635 = ~pi3  & ~n634;
  assign n636 = ~n289 & n331;
  assign n637 = n117 & n636;
  assign n638 = ~n635 & ~n637;
  assign n639 = ~n633 & n638;
  assign n640 = pi1  & ~n639;
  assign n641 = ~pi5  & ~n111;
  assign n642 = pi6  & ~n641;
  assign n643 = pi7  & ~n111;
  assign n644 = n216 & ~n392;
  assign n645 = ~n84 & ~n644;
  assign n646 = pi3  & n645;
  assign n647 = n292 & ~n331;
  assign n648 = ~pi2  & ~n647;
  assign n649 = ~n646 & n648;
  assign n650 = ~n266 & n630;
  assign n651 = n474 & n650;
  assign n652 = ~n649 & ~n651;
  assign n653 = ~pi1  & ~n652;
  assign n654 = ~n643 & ~n653;
  assign n655 = ~n642 & n654;
  assign n656 = ~n640 & n655;
  assign n657 = ~n629 & n656;
  assign n658 = ~n628 & n657;
  assign po9  = ~n625 & n658;
  assign n660 = n405 & n610;
  assign n661 = ~n412 & ~n660;
  assign po10  = n575 & ~n661;
endmodule
