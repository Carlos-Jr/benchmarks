module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n709, n710, n711, n712, n713,
    n714, n715, n716, n717, n718, n719, n720,
    n721, n722, n723, n724, n725, n726, n727,
    n728, n729, n730, n731, n732, n733, n734,
    n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755,
    n756, n757, n758, n759, n760, n761, n762,
    n763, n764, n765, n766, n767, n768, n769,
    n770, n771, n772, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n795, n796, n797,
    n798, n799, n800, n801, n802, n803, n804,
    n805, n806, n807, n808, n809, n810, n811,
    n812, n813, n814, n815, n816, n817, n818,
    n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853,
    n854, n855, n856, n857, n858, n859, n860,
    n861, n862, n863, n864, n865, n866, n867,
    n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944,
    n945, n946, n947, n948, n949, n950, n951,
    n952, n953, n954, n955, n956, n957, n958,
    n959, n960, n961, n962, n963, n964, n965,
    n966, n967, n968, n969, n970, n971, n972,
    n973, n974, n975, n976, n977, n978, n979,
    n980, n981, n982, n983, n984, n985, n986,
    n987, n988, n989, n990, n991, n992, n993,
    n994, n995, n996, n997, n998, n999, n1000,
    n1001, n1002, n1003, n1004, n1005, n1006,
    n1007, n1008, n1009, n1010, n1011, n1012,
    n1013, n1014, n1015, n1016, n1017, n1018,
    n1019, n1020, n1021, n1022, n1023, n1024,
    n1025, n1026, n1027, n1028, n1029, n1030,
    n1031, n1032, n1033, n1034, n1035, n1036,
    n1037, n1038, n1039, n1040, n1041, n1042,
    n1043, n1044, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1059, n1060,
    n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1083, n1084,
    n1085, n1086, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1105, n1106, n1107, n1108,
    n1109, n1110, n1111, n1112, n1113, n1114,
    n1115, n1116, n1117, n1118, n1119, n1120,
    n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1145,
    n1146, n1147, n1148, n1149, n1150, n1151,
    n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163,
    n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175,
    n1176, n1177, n1178, n1179, n1180, n1181,
    n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193,
    n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235,
    n1236, n1237, n1238, n1239, n1240, n1241,
    n1242, n1243, n1244, n1245, n1246, n1247,
    n1248, n1249, n1250, n1251, n1252, n1253,
    n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265,
    n1266, n1267, n1268, n1269, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1277,
    n1278, n1279, n1280, n1281, n1282, n1283,
    n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361,
    n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391,
    n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421,
    n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451,
    n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542,
    n1543, n1544, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639,
    n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1910, n1911, n1912,
    n1914, n1915, n1916, n1918, n1919, n1920,
    n1922, n1923, n1924, n1925, n1926, n1927,
    n1928, n1929, n1930, n1931, n1932, n1933,
    n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945,
    n1946, n1947, n1948, n1949, n1950, n1951,
    n1952, n1953, n1954, n1955, n1956, n1957,
    n1958, n1959, n1960, n1961, n1962, n1963,
    n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975,
    n1976, n1977, n1978, n1979, n1980, n1981,
    n1982, n1983, n1984, n1985, n1986, n1987,
    n1988, n1989, n1990, n1991, n1992, n1993,
    n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2082, n2083, n2084,
    n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2097, n2098,
    n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111,
    n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153,
    n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213,
    n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2264, n2265, n2266, n2267,
    n2268, n2269, n2270, n2271, n2272, n2273,
    n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285,
    n2286, n2287, n2288, n2289, n2290, n2291,
    n2292, n2293, n2294, n2295, n2296, n2297,
    n2298, n2299, n2300, n2301, n2302, n2303,
    n2304, n2305, n2306, n2307, n2308, n2309,
    n2310, n2311, n2312, n2313, n2314, n2315,
    n2316, n2317, n2318, n2319, n2320, n2321,
    n2322, n2323, n2324, n2325, n2326, n2327,
    n2328, n2329, n2330, n2331, n2332, n2333,
    n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345,
    n2346, n2347, n2348, n2349, n2350, n2351,
    n2352, n2353, n2354, n2355, n2356, n2357,
    n2358, n2359, n2360, n2361, n2362, n2363,
    n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375,
    n2376, n2377, n2378, n2379, n2380, n2381,
    n2382, n2383, n2384, n2385, n2386, n2387,
    n2388, n2389, n2390, n2391, n2392, n2393,
    n2394, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405,
    n2406, n2407, n2408, n2409, n2410, n2411,
    n2412, n2413, n2414, n2415, n2416, n2417,
    n2418, n2419, n2420, n2421, n2422, n2423,
    n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435,
    n2436, n2437, n2438, n2439, n2440, n2441,
    n2442, n2443, n2444, n2445, n2446, n2447,
    n2448, n2449, n2450, n2451, n2452, n2453,
    n2454, n2455, n2456, n2457, n2458, n2459,
    n2460, n2461, n2462, n2463, n2464, n2465,
    n2466, n2467, n2468, n2469, n2470, n2471,
    n2472, n2473, n2474, n2475, n2476, n2477,
    n2478, n2479, n2480, n2481, n2482, n2483,
    n2484, n2485, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495,
    n2496, n2497, n2498, n2499, n2500, n2501,
    n2502, n2503, n2504, n2505, n2506, n2507,
    n2508, n2509, n2510, n2511, n2512, n2513,
    n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531,
    n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561,
    n2562, n2563, n2564, n2565, n2566, n2567,
    n2568, n2569, n2570, n2571, n2572, n2573,
    n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2591,
    n2592, n2593, n2594, n2595, n2596, n2597,
    n2598, n2599, n2600, n2601, n2602, n2603,
    n2604, n2605, n2606, n2607, n2608, n2609,
    n2610, n2611, n2612, n2613, n2614, n2615,
    n2616, n2617, n2618, n2619, n2620, n2621,
    n2622, n2623, n2624, n2625, n2626, n2627,
    n2628, n2629, n2630, n2631, n2632, n2633,
    n2634, n2635, n2636, n2637, n2638, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645,
    n2646, n2647, n2648, n2649, n2650, n2651,
    n2652, n2653, n2654, n2655, n2656, n2657,
    n2658, n2659, n2660, n2661, n2662, n2663,
    n2664, n2665, n2666, n2667, n2668, n2669,
    n2670, n2671, n2672, n2673, n2674, n2675,
    n2676, n2677, n2678, n2679, n2680, n2681,
    n2682, n2683, n2684, n2685, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2693,
    n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705,
    n2706, n2707, n2708, n2709, n2710, n2711,
    n2712, n2713, n2714, n2715, n2716, n2717,
    n2718, n2719, n2720, n2721, n2722, n2723,
    n2724, n2725, n2726, n2727, n2728, n2729,
    n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2761, n2763,
    n2766, n2767, n2768, n2769, n2770, n2771,
    n2772, n2773, n2774, n2775, n2776, n2777,
    n2778, n2779, n2780, n2781, n2782, n2783,
    n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795,
    n2796, n2797, n2798, n2799, n2800, n2801,
    n2802, n2803, n2804, n2805, n2806, n2807,
    n2808, n2809, n2810, n2812, n2813, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821,
    n2823, n2824, n2825, n2826, n2827, n2828,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2862, n2863, n2864, n2865, n2866,
    n2868, n2869, n2871, n2872, n2874, n2875,
    n2876, n2877, n2879, n2880, n2881, n2883,
    n2884, n2886, n2887, n2888, n2890, n2891,
    n2892, n2894, n2895, n2896, n2897, n2899,
    n2900, n2902, n2903, n2904, n2905, n2906,
    n2907, n2909, n2910, n2912, n2913, n2914,
    n2915, n2917, n2918, n2919, n2920, n2921,
    n2922, n2923, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2935,
    n2936, n2937, n2938, n2940, n2941, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2954, n2955, n2956,
    n2957, n2958, n2959, n2960, n2961, n2962,
    n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2972, n2973, n2974, n2976,
    n2977, n2978, n2979, n2981, n2982, n2983,
    n2984, n2985, n2986, n2988, n2989, n2991,
    n2992, n2994, n2995, n2996, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3006,
    n3007, n3008, n3010, n3011, n3013, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3026, n3027, n3029,
    n3030, n3032, n3033, n3035, n3036, n3038,
    n3039, n3041, n3042, n3044, n3045, n3048,
    n3050, n3051, n3053, n3055, n3056, n3058,
    n3059, n3061, n3062, n3063, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3107,
    n3116, n3117, n3118, n3119, n3121, n3125;
  assign po12 = 1'b1;
  assign n291 = pi122 & pi127;
  assign n292 = ~pi82 & ~n291;
  assign n293 = ~pi38 & ~pi50;
  assign n294 = ~pi42 & ~pi44;
  assign n295 = ~pi40 & n294;
  assign n296 = ~pi40 & ~pi42;
  assign n297 = ~pi38 & ~pi40;
  assign n298 = ~pi42 & ~pi50;
  assign n299 = n297 & n298;
  assign n300 = ~pi42 & n297;
  assign n301 = ~pi38 & n296;
  assign n302 = ~pi50 & n2767;
  assign n303 = n293 & n296;
  assign n304 = ~pi44 & n2766;
  assign n305 = ~pi50 & n294;
  assign n306 = n297 & n305;
  assign n307 = n294 & n297;
  assign n308 = ~pi50 & n307;
  assign n309 = n293 & n295;
  assign n310 = ~pi41 & ~pi46;
  assign n311 = ~pi43 & n310;
  assign n312 = ~pi47 & ~pi48;
  assign n313 = ~pi45 & n312;
  assign n314 = ~pi43 & ~pi47;
  assign n315 = n310 & n314;
  assign n316 = ~pi45 & ~pi48;
  assign n317 = n315 & n316;
  assign n318 = n311 & n313;
  assign n319 = ~pi46 & ~pi50;
  assign n320 = ~pi50 & n310;
  assign n321 = ~pi41 & n319;
  assign n322 = ~pi43 & n312;
  assign n323 = ~pi48 & n314;
  assign n324 = n310 & n2771;
  assign n325 = n311 & n312;
  assign n326 = ~pi50 & n2772;
  assign n327 = n2770 & n2771;
  assign n328 = ~pi38 & ~pi46;
  assign n329 = ~pi46 & n293;
  assign n330 = ~pi50 & n328;
  assign n331 = ~pi40 & n2774;
  assign n332 = n297 & n319;
  assign n333 = n294 & n2775;
  assign n334 = n295 & n319;
  assign n335 = ~pi38 & n334;
  assign n336 = ~pi46 & n2768;
  assign n337 = n295 & n2774;
  assign n338 = ~pi41 & ~pi43;
  assign n339 = ~pi47 & n338;
  assign n340 = n2768 & n310;
  assign n341 = n307 & n2770;
  assign n342 = ~pi43 & n2777;
  assign n343 = n2776 & n338;
  assign n344 = ~pi47 & n2778;
  assign n345 = n2768 & n315;
  assign n346 = n314 & n2777;
  assign n347 = n2776 & n339;
  assign n348 = ~pi48 & n2779;
  assign n349 = ~pi48 & n2766;
  assign n350 = n315 & n349;
  assign n351 = ~pi44 & n350;
  assign n352 = n2768 & n2772;
  assign n353 = n2766 & n315;
  assign n354 = ~pi44 & ~pi48;
  assign n355 = n353 & n354;
  assign n356 = n307 & n2773;
  assign n357 = ~pi45 & n2780;
  assign n358 = n316 & n2779;
  assign n359 = n313 & n2778;
  assign n360 = n316 & n339;
  assign n361 = n2776 & n360;
  assign n362 = n2768 & n2769;
  assign n363 = ~pi2 & ~pi20;
  assign n364 = ~pi15 & ~pi49;
  assign n365 = ~pi15 & ~pi20;
  assign n366 = ~pi2 & n365;
  assign n367 = ~pi49 & n366;
  assign n368 = n363 & n364;
  assign n369 = ~pi24 & ~pi49;
  assign n370 = n366 & n369;
  assign n371 = ~pi24 & n2782;
  assign n372 = ~n291 & n2783;
  assign n373 = n2781 & n372;
  assign n374 = ~pi2 & n316;
  assign n375 = n314 & n374;
  assign n376 = ~pi15 & n369;
  assign n377 = ~pi24 & n364;
  assign n378 = ~pi20 & n2784;
  assign n379 = n365 & n369;
  assign n380 = ~pi41 & n2774;
  assign n381 = ~pi38 & n2770;
  assign n382 = n293 & n310;
  assign n383 = n2785 & n2786;
  assign n384 = n295 & n383;
  assign n385 = n314 & n316;
  assign n386 = n2785 & n385;
  assign n387 = ~pi2 & n295;
  assign n388 = n2786 & n387;
  assign n389 = n386 & n388;
  assign n390 = n2781 & n2783;
  assign n391 = ~pi2 & ~pi45;
  assign n392 = n312 & n391;
  assign n393 = ~pi49 & n365;
  assign n394 = ~pi24 & ~pi45;
  assign n395 = ~pi2 & ~pi48;
  assign n396 = n394 & n395;
  assign n397 = ~pi45 & n2783;
  assign n398 = n2785 & n391;
  assign n399 = n2782 & n394;
  assign n400 = ~pi48 & n2788;
  assign n401 = n316 & n2783;
  assign n402 = n393 & n396;
  assign n403 = ~pi47 & n2789;
  assign n404 = ~pi2 & n312;
  assign n405 = n2785 & n404;
  assign n406 = ~pi45 & n405;
  assign n407 = n2785 & n392;
  assign n408 = n2778 & n2790;
  assign n409 = n375 & n384;
  assign n410 = pi82 & ~n2787;
  assign n411 = ~n291 & ~n410;
  assign n412 = ~n292 & ~n373;
  assign n413 = ~pi65 & ~n291;
  assign n414 = ~n410 & n413;
  assign n415 = ~pi65 & n2791;
  assign n416 = ~pi24 & n316;
  assign n417 = n315 & n416;
  assign n418 = ~pi50 & n297;
  assign n419 = n294 & n364;
  assign n420 = n418 & n419;
  assign n421 = n2781 & n2784;
  assign n422 = ~pi45 & n369;
  assign n423 = ~pi49 & n394;
  assign n424 = n312 & n338;
  assign n425 = n2794 & n424;
  assign n426 = ~pi15 & n2776;
  assign n427 = n425 & n426;
  assign n428 = ~pi48 & n2794;
  assign n429 = n316 & n369;
  assign n430 = n314 & n2795;
  assign n431 = n2771 & n2794;
  assign n432 = n2779 & n2795;
  assign n433 = ~pi44 & n418;
  assign n434 = ~pi24 & ~pi42;
  assign n435 = n433 & n434;
  assign n436 = n2769 & n435;
  assign n437 = ~pi24 & n2781;
  assign n438 = n2769 & n434;
  assign n439 = n433 & n438;
  assign n440 = n2780 & n394;
  assign n441 = ~pi49 & n2798;
  assign n442 = n2781 & n369;
  assign n443 = n2768 & n369;
  assign n444 = n2769 & n443;
  assign n445 = n2780 & n2794;
  assign n446 = n2777 & n2796;
  assign n447 = ~pi15 & n2797;
  assign n448 = ~pi15 & n2795;
  assign n449 = n2779 & n448;
  assign n450 = ~pi15 & n312;
  assign n451 = n338 & n450;
  assign n452 = n2794 & n451;
  assign n453 = n2776 & n452;
  assign n454 = n364 & n2798;
  assign n455 = n417 & n420;
  assign n456 = ~pi20 & pi82;
  assign n457 = n2793 & n456;
  assign n458 = pi2 & ~n292;
  assign n459 = pi82 & ~n2781;
  assign n460 = ~pi82 & n291;
  assign n461 = pi82 & ~n2785;
  assign n462 = ~n460 & ~n461;
  assign n463 = n365 & n2797;
  assign n464 = n2781 & n2785;
  assign n465 = ~pi44 & n393;
  assign n466 = n2766 & n465;
  assign n467 = n417 & n466;
  assign n468 = n312 & n394;
  assign n469 = n393 & n468;
  assign n470 = n2778 & n469;
  assign n471 = ~pi20 & n2793;
  assign n472 = pi82 & ~n2799;
  assign n473 = ~n460 & ~n472;
  assign n474 = ~n459 & n462;
  assign n475 = pi2 & ~n2800;
  assign n476 = ~n457 & n458;
  assign n477 = ~n2792 & ~n2801;
  assign po17 = ~pi129 & ~n477;
  assign n479 = ~pi3 & ~pi129;
  assign n480 = pi5 & ~pi54;
  assign n481 = ~pi5 & ~pi6;
  assign n482 = ~pi7 & ~pi12;
  assign n483 = ~pi6 & ~pi12;
  assign n484 = ~pi5 & ~pi7;
  assign n485 = n483 & n484;
  assign n486 = n481 & n482;
  assign n487 = ~pi16 & pi54;
  assign n488 = n2802 & n487;
  assign n489 = ~pi4 & ~pi19;
  assign n490 = ~pi4 & ~pi18;
  assign n491 = ~pi19 & n490;
  assign n492 = ~pi18 & n489;
  assign n493 = ~pi25 & pi28;
  assign n494 = ~pi25 & ~pi29;
  assign n495 = pi28 & n494;
  assign n496 = ~pi29 & n493;
  assign n497 = n2803 & n2804;
  assign n498 = n488 & n497;
  assign n499 = ~pi10 & ~pi22;
  assign n500 = ~pi9 & ~pi14;
  assign n501 = ~pi9 & ~pi10;
  assign n502 = ~pi22 & n501;
  assign n503 = ~pi9 & n499;
  assign n504 = ~pi14 & n2805;
  assign n505 = n499 & n500;
  assign n506 = ~pi13 & n2806;
  assign n507 = ~pi8 & ~pi21;
  assign n508 = ~pi8 & ~pi17;
  assign n509 = ~pi21 & n508;
  assign n510 = ~pi17 & ~pi21;
  assign n511 = ~pi8 & n510;
  assign n512 = ~pi17 & n507;
  assign n513 = ~pi11 & ~pi59;
  assign n514 = ~pi11 & n507;
  assign n515 = ~pi17 & ~pi59;
  assign n516 = n514 & n515;
  assign n517 = ~pi8 & ~pi11;
  assign n518 = n510 & n517;
  assign n519 = ~pi59 & n518;
  assign n520 = n2807 & n513;
  assign n521 = n506 & n2808;
  assign n522 = n488 & n2808;
  assign n523 = n506 & n522;
  assign n524 = ~pi29 & n523;
  assign n525 = n2803 & n493;
  assign n526 = n524 & n525;
  assign n527 = ~pi6 & ~pi7;
  assign n528 = ~pi7 & n483;
  assign n529 = ~pi12 & n527;
  assign n530 = n2804 & n2810;
  assign n531 = n506 & n530;
  assign n532 = ~pi5 & n2803;
  assign n533 = n487 & n532;
  assign n534 = n2808 & n533;
  assign n535 = n531 & n534;
  assign n536 = n498 & n521;
  assign n537 = ~n480 & ~n2809;
  assign n538 = ~pi129 & ~n537;
  assign n539 = ~pi3 & n538;
  assign n540 = n479 & ~n537;
  assign n541 = pi6 & ~pi54;
  assign n542 = pi25 & ~pi28;
  assign n543 = pi25 & ~pi29;
  assign n544 = ~pi28 & n543;
  assign n545 = ~pi28 & ~pi29;
  assign n546 = pi25 & n545;
  assign n547 = ~pi29 & n542;
  assign n548 = n2803 & n2812;
  assign n549 = n488 & n548;
  assign n550 = n2803 & n542;
  assign n551 = n524 & n550;
  assign n552 = ~pi12 & n2812;
  assign n553 = n484 & n552;
  assign n554 = n506 & n553;
  assign n555 = ~pi6 & n2803;
  assign n556 = n487 & n555;
  assign n557 = n2808 & n556;
  assign n558 = n554 & n557;
  assign n559 = n521 & n549;
  assign n560 = ~n541 & ~n2813;
  assign n561 = ~pi129 & ~n560;
  assign n562 = ~pi3 & n561;
  assign n563 = n479 & ~n560;
  assign n564 = pi13 & ~pi54;
  assign n565 = ~pi25 & ~pi28;
  assign n566 = ~pi25 & pi29;
  assign n567 = ~pi28 & n566;
  assign n568 = pi29 & n565;
  assign n569 = n2803 & n2815;
  assign n570 = n488 & n569;
  assign n571 = n523 & n569;
  assign n572 = ~pi13 & n2803;
  assign n573 = n487 & n572;
  assign n574 = n2808 & n573;
  assign n575 = ~pi5 & n483;
  assign n576 = n2815 & n575;
  assign n577 = ~pi7 & n2806;
  assign n578 = n576 & n577;
  assign n579 = n574 & n578;
  assign n580 = ~pi4 & ~pi16;
  assign n581 = ~pi18 & ~pi19;
  assign n582 = ~pi16 & n2803;
  assign n583 = ~pi16 & n489;
  assign n584 = ~pi18 & n583;
  assign n585 = n580 & n581;
  assign n586 = n487 & n2803;
  assign n587 = pi54 & n583;
  assign n588 = n487 & n489;
  assign n589 = ~pi18 & n2819;
  assign n590 = pi54 & n2817;
  assign n591 = n2815 & n2818;
  assign n592 = ~pi7 & ~pi13;
  assign n593 = n481 & n592;
  assign n594 = n2806 & n593;
  assign n595 = ~pi12 & n594;
  assign n596 = ~pi12 & n593;
  assign n597 = n575 & n592;
  assign n598 = ~pi13 & n2802;
  assign n599 = n2806 & n2821;
  assign n600 = n2802 & n506;
  assign n601 = n2808 & n2820;
  assign n602 = n591 & n601;
  assign n603 = n2803 & n2806;
  assign n604 = n2815 & n603;
  assign n605 = n487 & n592;
  assign n606 = n575 & n605;
  assign n607 = n2808 & n606;
  assign n608 = n604 & n607;
  assign n609 = n521 & n570;
  assign n610 = ~n564 & ~n2816;
  assign n611 = ~pi129 & ~n610;
  assign n612 = ~pi3 & n611;
  assign n613 = n479 & ~n610;
  assign n614 = ~pi15 & ~n363;
  assign n615 = n2778 & n614;
  assign n616 = n369 & n615;
  assign n617 = n313 & n616;
  assign n618 = ~n363 & n2784;
  assign n619 = n2781 & n618;
  assign n620 = n313 & n618;
  assign n621 = n2778 & n620;
  assign n622 = ~n363 & n2793;
  assign n623 = pi15 & ~n2797;
  assign n624 = ~n2823 & ~n623;
  assign n625 = pi82 & ~n624;
  assign n626 = pi15 & n460;
  assign n627 = pi82 & ~n2793;
  assign n628 = ~pi70 & ~n291;
  assign n629 = ~n291 & ~n627;
  assign n630 = ~pi70 & n629;
  assign n631 = ~n627 & n628;
  assign n632 = ~n626 & ~n2824;
  assign n633 = ~n625 & ~n626;
  assign n634 = ~n2824 & n633;
  assign n635 = ~n625 & n632;
  assign po30 = ~pi129 & ~n2825;
  assign n637 = pi17 & ~pi54;
  assign n638 = ~pi7 & n481;
  assign n639 = ~pi12 & n565;
  assign n640 = n638 & n639;
  assign n641 = n506 & n640;
  assign n642 = ~pi17 & ~pi18;
  assign n643 = ~pi17 & pi54;
  assign n644 = ~pi16 & n643;
  assign n645 = n2803 & n644;
  assign n646 = n2819 & n642;
  assign n647 = ~pi29 & pi59;
  assign n648 = n514 & n647;
  assign n649 = n2826 & n648;
  assign n650 = n514 & n643;
  assign n651 = n565 & n647;
  assign n652 = n2802 & n651;
  assign n653 = n2817 & n652;
  assign n654 = n2802 & n545;
  assign n655 = ~pi25 & pi59;
  assign n656 = n643 & n655;
  assign n657 = n514 & n656;
  assign n658 = n654 & n657;
  assign n659 = n2817 & n658;
  assign n660 = n650 & n653;
  assign n661 = n506 & n2827;
  assign n662 = pi59 & n545;
  assign n663 = n2803 & n662;
  assign n664 = n514 & n663;
  assign n665 = ~pi16 & ~pi25;
  assign n666 = n482 & n665;
  assign n667 = n481 & n643;
  assign n668 = n666 & n667;
  assign n669 = n506 & n668;
  assign n670 = n664 & n669;
  assign n671 = n641 & n649;
  assign n672 = ~n637 & ~n2828;
  assign n673 = ~pi129 & ~n672;
  assign n674 = ~pi3 & n673;
  assign n675 = n479 & ~n672;
  assign n676 = pi0 & ~pi113;
  assign n677 = pi0 & ~pi123;
  assign n678 = ~pi113 & n677;
  assign n679 = ~pi123 & n676;
  assign n680 = n2817 & n593;
  assign n681 = ~pi11 & ~pi12;
  assign n682 = ~pi21 & n681;
  assign n683 = n508 & n682;
  assign n684 = n2807 & n681;
  assign n685 = n2806 & n2831;
  assign n686 = n499 & n593;
  assign n687 = n2817 & n686;
  assign n688 = n500 & n2831;
  assign n689 = n687 & n688;
  assign n690 = n508 & n681;
  assign n691 = ~pi21 & n2817;
  assign n692 = n690 & n691;
  assign n693 = n2817 & n2831;
  assign n694 = n594 & n2833;
  assign n695 = n680 & n685;
  assign n696 = ~pi61 & ~pi118;
  assign n697 = ~n2832 & n696;
  assign n698 = ~n2830 & ~n697;
  assign po18 = ~pi129 & ~n698;
  assign n700 = n583 & n642;
  assign n701 = ~pi17 & n2817;
  assign n702 = ~pi5 & ~pi22;
  assign n703 = n483 & n702;
  assign n704 = ~pi17 & n702;
  assign n705 = n483 & n704;
  assign n706 = n2817 & n705;
  assign n707 = n2834 & n703;
  assign n708 = ~pi9 & ~pi11;
  assign n709 = ~pi13 & n507;
  assign n710 = ~pi7 & n709;
  assign n711 = n507 & n592;
  assign n712 = pi7 & ~n507;
  assign n713 = ~pi14 & ~n712;
  assign n714 = n2836 & n713;
  assign n715 = ~pi14 & n2836;
  assign n716 = n708 & n2837;
  assign n717 = ~pi13 & ~pi14;
  assign n718 = n527 & n717;
  assign n719 = ~pi12 & n2807;
  assign n720 = n718 & n719;
  assign n721 = n702 & n708;
  assign n722 = n2817 & n721;
  assign n723 = n720 & n722;
  assign n724 = n703 & n708;
  assign n725 = ~pi18 & ~pi21;
  assign n726 = n508 & n725;
  assign n727 = n507 & n642;
  assign n728 = ~pi14 & n592;
  assign n729 = n583 & n728;
  assign n730 = n2839 & n729;
  assign n731 = n724 & n730;
  assign n732 = n708 & n728;
  assign n733 = n2807 & n703;
  assign n734 = n732 & n733;
  assign n735 = n2817 & n734;
  assign n736 = n702 & n717;
  assign n737 = n708 & n736;
  assign n738 = n2807 & n2810;
  assign n739 = n2817 & n738;
  assign n740 = n737 & n739;
  assign n741 = n2835 & n716;
  assign n742 = pi54 & ~n2838;
  assign n743 = ~pi0 & ~n742;
  assign n744 = ~n2836 & ~n713;
  assign n745 = ~pi7 & n507;
  assign n746 = pi8 & pi21;
  assign n747 = ~pi13 & ~n746;
  assign n748 = ~n745 & ~n747;
  assign n749 = ~pi10 & ~n748;
  assign n750 = pi14 & ~n2836;
  assign n751 = pi13 & ~n507;
  assign n752 = ~pi7 & ~n746;
  assign n753 = ~n751 & n752;
  assign n754 = ~n709 & ~n753;
  assign n755 = ~pi10 & ~n754;
  assign n756 = ~n750 & n755;
  assign n757 = ~n744 & n749;
  assign n758 = ~n2837 & ~n2840;
  assign n759 = ~pi10 & n2837;
  assign n760 = n2835 & ~n759;
  assign n761 = ~pi7 & pi13;
  assign n762 = n507 & n761;
  assign n763 = ~n745 & n747;
  assign n764 = ~n712 & ~n745;
  assign n765 = n747 & n764;
  assign n766 = ~n712 & n763;
  assign n767 = ~n762 & ~n2841;
  assign n768 = ~pi14 & ~n767;
  assign n769 = ~pi13 & pi14;
  assign n770 = n745 & n769;
  assign n771 = ~n768 & ~n770;
  assign n772 = ~pi10 & ~n771;
  assign n773 = ~pi14 & ~n748;
  assign n774 = ~n2836 & ~n773;
  assign n775 = ~n2836 & ~n712;
  assign n776 = ~pi14 & ~n775;
  assign n777 = ~pi10 & ~n776;
  assign n778 = ~n774 & n777;
  assign n779 = ~n2837 & n2840;
  assign n780 = pi10 & n717;
  assign n781 = ~pi14 & n507;
  assign n782 = pi10 & n592;
  assign n783 = n781 & n782;
  assign n784 = n745 & n780;
  assign n785 = ~n2842 & ~n2843;
  assign n786 = n702 & ~n785;
  assign n787 = n2817 & n786;
  assign n788 = ~pi17 & n787;
  assign n789 = n483 & n788;
  assign n790 = n2835 & ~n785;
  assign n791 = ~n758 & n760;
  assign n792 = ~pi56 & ~n702;
  assign n793 = n708 & ~n792;
  assign n794 = ~n2844 & n793;
  assign n795 = ~pi56 & n702;
  assign n796 = ~n708 & ~n795;
  assign n797 = pi54 & ~n796;
  assign n798 = n702 & ~n708;
  assign n799 = ~pi56 & n798;
  assign n800 = ~n708 & n795;
  assign n801 = ~n2844 & ~n792;
  assign n802 = n708 & ~n801;
  assign n803 = ~n2845 & ~n802;
  assign n804 = pi54 & ~n803;
  assign n805 = ~n794 & n797;
  assign n806 = ~n743 & ~n2846;
  assign n807 = ~pi129 & ~n806;
  assign n808 = ~pi3 & n807;
  assign n809 = n479 & ~n806;
  assign n810 = ~pi12 & ~pi14;
  assign n811 = n499 & n810;
  assign n812 = n499 & n681;
  assign n813 = n781 & n812;
  assign n814 = n514 & n811;
  assign n815 = n507 & n681;
  assign n816 = n2817 & n815;
  assign n817 = ~pi14 & n593;
  assign n818 = n499 & n817;
  assign n819 = n816 & n818;
  assign n820 = n681 & n781;
  assign n821 = n687 & n820;
  assign n822 = n593 & n2848;
  assign n823 = n2817 & n822;
  assign n824 = n680 & n2848;
  assign n825 = n643 & ~n2849;
  assign n826 = ~pi1 & ~n825;
  assign n827 = ~n483 & n484;
  assign n828 = n483 & ~n484;
  assign n829 = ~n827 & ~n828;
  assign n830 = ~n481 & ~n482;
  assign n831 = ~pi13 & ~n830;
  assign n832 = pi5 & ~n483;
  assign n833 = pi6 & pi12;
  assign n834 = ~pi7 & ~n833;
  assign n835 = ~n575 & n834;
  assign n836 = ~n575 & ~n832;
  assign n837 = n834 & n836;
  assign n838 = ~n832 & n835;
  assign n839 = pi7 & n575;
  assign n840 = ~n2850 & ~n839;
  assign n841 = ~pi13 & ~n840;
  assign n842 = ~n829 & n831;
  assign n843 = pi13 & n2802;
  assign n844 = n575 & n761;
  assign n845 = ~pi9 & ~n2852;
  assign n846 = pi13 & ~n2802;
  assign n847 = ~n483 & ~n484;
  assign n848 = ~n830 & ~n847;
  assign n849 = ~n846 & n848;
  assign n850 = ~pi13 & ~n847;
  assign n851 = ~n2802 & ~n850;
  assign n852 = ~n2821 & ~n830;
  assign n853 = ~n851 & n852;
  assign n854 = ~n2851 & ~n2852;
  assign n855 = ~n2821 & n849;
  assign n856 = ~pi9 & ~n2853;
  assign n857 = ~n2851 & n845;
  assign n858 = pi9 & ~n2821;
  assign n859 = ~pi14 & pi54;
  assign n860 = pi54 & n499;
  assign n861 = ~pi14 & n860;
  assign n862 = n499 & n859;
  assign n863 = n2817 & n2855;
  assign n864 = n514 & n2834;
  assign n865 = n2855 & n864;
  assign n866 = n518 & n863;
  assign n867 = ~n858 & n2855;
  assign n868 = n864 & n867;
  assign n869 = ~n858 & n2856;
  assign n870 = ~pi9 & n2853;
  assign n871 = pi9 & n2821;
  assign n872 = ~n870 & ~n871;
  assign n873 = n2817 & ~n872;
  assign n874 = n518 & n873;
  assign n875 = n859 & n874;
  assign n876 = n499 & n875;
  assign n877 = n2856 & ~n872;
  assign n878 = ~n2854 & n2857;
  assign n879 = ~n826 & ~n2858;
  assign n880 = ~pi129 & ~n879;
  assign n881 = ~pi3 & n880;
  assign n882 = n479 & ~n879;
  assign n883 = pi4 & ~pi54;
  assign n884 = ~pi11 & n489;
  assign n885 = n487 & n884;
  assign n886 = n2839 & n885;
  assign n887 = pi54 & n864;
  assign n888 = n518 & n2818;
  assign n889 = n2817 & n650;
  assign n890 = pi10 & ~pi22;
  assign n891 = n500 & n890;
  assign n892 = n2821 & n891;
  assign n893 = n2860 & n892;
  assign n894 = ~n883 & ~n893;
  assign n895 = ~pi129 & ~n894;
  assign n896 = ~pi3 & n895;
  assign n897 = n479 & ~n894;
  assign n898 = pi7 & ~pi54;
  assign n899 = n484 & n506;
  assign n900 = ~pi6 & n681;
  assign n901 = ~pi11 & n483;
  assign n902 = n2819 & n2862;
  assign n903 = pi8 & ~pi21;
  assign n904 = pi8 & ~pi17;
  assign n905 = n725 & n904;
  assign n906 = n642 & n903;
  assign n907 = n902 & n2863;
  assign n908 = ~pi7 & n489;
  assign n909 = n487 & n908;
  assign n910 = n2863 & n909;
  assign n911 = ~pi5 & n2862;
  assign n912 = n506 & n911;
  assign n913 = n910 & n912;
  assign n914 = n484 & n903;
  assign n915 = n484 & n2863;
  assign n916 = n642 & n914;
  assign n917 = n506 & n2865;
  assign n918 = n902 & n917;
  assign n919 = n2819 & n725;
  assign n920 = n484 & n904;
  assign n921 = n2862 & n920;
  assign n922 = n902 & n2865;
  assign n923 = n919 & n921;
  assign n924 = n506 & n2866;
  assign n925 = n899 & n907;
  assign n926 = ~n898 & ~n2864;
  assign n927 = ~pi129 & ~n926;
  assign n928 = ~pi3 & n927;
  assign n929 = n479 & ~n926;
  assign n930 = pi8 & ~pi54;
  assign n931 = n517 & n642;
  assign n932 = pi21 & n2819;
  assign n933 = ~pi11 & pi21;
  assign n934 = n642 & n933;
  assign n935 = ~pi8 & n489;
  assign n936 = n487 & n935;
  assign n937 = n934 & n936;
  assign n938 = pi21 & n642;
  assign n939 = pi21 & n931;
  assign n940 = n517 & n938;
  assign n941 = n2819 & n2869;
  assign n942 = pi21 & n517;
  assign n943 = n2826 & n942;
  assign n944 = n931 & n932;
  assign n945 = n2820 & n2868;
  assign n946 = ~n930 & ~n945;
  assign n947 = ~pi129 & ~n946;
  assign n948 = ~pi3 & n947;
  assign n949 = n479 & ~n946;
  assign n950 = pi9 & ~pi54;
  assign n951 = n2803 & n506;
  assign n952 = pi11 & n2807;
  assign n953 = n488 & n952;
  assign n954 = n499 & n717;
  assign n955 = pi11 & n484;
  assign n956 = n483 & n955;
  assign n957 = n954 & n956;
  assign n958 = ~pi9 & n489;
  assign n959 = n487 & n958;
  assign n960 = n2839 & n959;
  assign n961 = n957 & n960;
  assign n962 = pi11 & n2803;
  assign n963 = n2803 & n952;
  assign n964 = n2807 & n962;
  assign n965 = n488 & n2872;
  assign n966 = n506 & n965;
  assign n967 = n499 & n2819;
  assign n968 = ~pi9 & pi11;
  assign n969 = n717 & n968;
  assign n970 = n2802 & n969;
  assign n971 = n2839 & n970;
  assign n972 = n967 & n971;
  assign n973 = n951 & n953;
  assign n974 = ~n950 & ~n2871;
  assign n975 = ~pi129 & ~n974;
  assign n976 = ~pi3 & n975;
  assign n977 = n479 & ~n974;
  assign n978 = pi10 & ~pi54;
  assign n979 = n2805 & n2839;
  assign n980 = ~pi11 & ~pi13;
  assign n981 = pi14 & n980;
  assign n982 = n2802 & n981;
  assign n983 = ~pi11 & n2802;
  assign n984 = n484 & n2862;
  assign n985 = n487 & n769;
  assign n986 = n2819 & n769;
  assign n987 = n489 & n985;
  assign n988 = n2874 & n2875;
  assign n989 = n2819 & n982;
  assign n990 = ~pi10 & n489;
  assign n991 = n487 & n990;
  assign n992 = n2839 & n991;
  assign n993 = ~pi9 & ~pi22;
  assign n994 = n769 & n993;
  assign n995 = n2874 & n994;
  assign n996 = n992 & n995;
  assign n997 = n979 & n2874;
  assign n998 = n2875 & n997;
  assign n999 = n979 & n2875;
  assign n1000 = n2874 & n999;
  assign n1001 = n979 & n2876;
  assign n1002 = ~n978 & ~n2877;
  assign n1003 = ~pi129 & ~n1002;
  assign n1004 = ~pi3 & n1003;
  assign n1005 = n479 & ~n1002;
  assign n1006 = pi11 & ~pi54;
  assign n1007 = ~pi10 & ~pi14;
  assign n1008 = pi22 & n1007;
  assign n1009 = ~pi10 & ~pi11;
  assign n1010 = pi22 & n1009;
  assign n1011 = n500 & n1010;
  assign n1012 = n708 & n1008;
  assign n1013 = n2819 & n2839;
  assign n1014 = n487 & n500;
  assign n1015 = n489 & n1014;
  assign n1016 = n2839 & n1010;
  assign n1017 = n1015 & n1016;
  assign n1018 = n2879 & n1013;
  assign n1019 = ~pi10 & pi22;
  assign n1020 = n500 & n1019;
  assign n1021 = n2821 & n1020;
  assign n1022 = n2860 & n1021;
  assign n1023 = n2839 & n2879;
  assign n1024 = n2819 & n2821;
  assign n1025 = n1023 & n1024;
  assign n1026 = n2821 & n2880;
  assign n1027 = ~n1006 & ~n2881;
  assign n1028 = ~pi129 & ~n1027;
  assign n1029 = ~pi3 & n1028;
  assign n1030 = n479 & ~n1027;
  assign n1031 = pi12 & ~pi54;
  assign n1032 = pi18 & n593;
  assign n1033 = n2819 & n1032;
  assign n1034 = ~pi12 & n489;
  assign n1035 = n487 & n1034;
  assign n1036 = pi18 & n2807;
  assign n1037 = n1035 & n1036;
  assign n1038 = ~pi11 & n594;
  assign n1039 = n1037 & n1038;
  assign n1040 = n2831 & n1032;
  assign n1041 = n2806 & n2819;
  assign n1042 = n1040 & n1041;
  assign n1043 = pi18 & n681;
  assign n1044 = n2819 & n1043;
  assign n1045 = pi18 & n2819;
  assign n1046 = n2831 & n1045;
  assign n1047 = n2807 & n1044;
  assign n1048 = n594 & n2884;
  assign n1049 = n685 & n1033;
  assign n1050 = ~n1031 & ~n2883;
  assign n1051 = ~pi129 & ~n1050;
  assign n1052 = ~pi3 & n1051;
  assign n1053 = n479 & ~n1050;
  assign n1054 = pi14 & ~pi54;
  assign n1055 = pi13 & n500;
  assign n1056 = n2802 & n1055;
  assign n1057 = n860 & n1056;
  assign n1058 = ~pi16 & n859;
  assign n1059 = n489 & n1058;
  assign n1060 = n2839 & n1059;
  assign n1061 = ~pi9 & pi13;
  assign n1062 = n499 & n1061;
  assign n1063 = n2874 & n1062;
  assign n1064 = n1060 & n1063;
  assign n1065 = n489 & n2855;
  assign n1066 = ~pi16 & n1061;
  assign n1067 = n2839 & n1066;
  assign n1068 = n583 & n1061;
  assign n1069 = n489 & n1066;
  assign n1070 = n2839 & n2855;
  assign n1071 = n2887 & n1070;
  assign n1072 = n1065 & n1067;
  assign n1073 = n2874 & n2888;
  assign n1074 = n864 & n1057;
  assign n1075 = ~n1054 & ~n2886;
  assign n1076 = ~pi129 & ~n1075;
  assign n1077 = ~pi3 & n1076;
  assign n1078 = n479 & ~n1075;
  assign n1079 = pi16 & ~pi54;
  assign n1080 = ~pi5 & pi6;
  assign n1081 = pi6 & ~pi12;
  assign n1082 = ~pi5 & n1081;
  assign n1083 = ~pi12 & n1080;
  assign n1084 = n592 & n2890;
  assign n1085 = n482 & n1080;
  assign n1086 = n506 & n1085;
  assign n1087 = n2806 & n1084;
  assign n1088 = n2860 & n1081;
  assign n1089 = n899 & n1088;
  assign n1090 = n2860 & n2891;
  assign n1091 = ~n1079 & ~n2892;
  assign n1092 = ~pi129 & ~n1091;
  assign n1093 = ~pi3 & n1092;
  assign n1094 = n479 & ~n1091;
  assign n1095 = pi18 & ~pi54;
  assign n1096 = pi16 & pi54;
  assign n1097 = pi16 & n650;
  assign n1098 = n518 & n1096;
  assign n1099 = n2803 & n1096;
  assign n1100 = n518 & n1099;
  assign n1101 = pi16 & n643;
  assign n1102 = n2803 & n1101;
  assign n1103 = n514 & n1102;
  assign n1104 = n2803 & n2894;
  assign n1105 = n2803 & n2820;
  assign n1106 = n2802 & n951;
  assign n1107 = n2894 & n2896;
  assign n1108 = n2820 & n2895;
  assign n1109 = ~n1095 & ~n2897;
  assign n1110 = ~pi129 & ~n1109;
  assign n1111 = ~pi3 & n1110;
  assign n1112 = n479 & ~n1109;
  assign n1113 = pi19 & ~pi54;
  assign n1114 = pi17 & ~pi18;
  assign n1115 = n489 & n1114;
  assign n1116 = n487 & n1115;
  assign n1117 = pi17 & n514;
  assign n1118 = n2818 & n1117;
  assign n1119 = pi17 & pi54;
  assign n1120 = n514 & n1119;
  assign n1121 = n2817 & n1120;
  assign n1122 = n514 & n1116;
  assign n1123 = pi17 & n487;
  assign n1124 = n514 & n1123;
  assign n1125 = n2896 & n1124;
  assign n1126 = n2820 & n2899;
  assign n1127 = ~n1113 & ~n2900;
  assign n1128 = ~pi129 & ~n1127;
  assign n1129 = ~pi3 & n1128;
  assign n1130 = n479 & ~n1127;
  assign n1131 = pi2 & n2799;
  assign n1132 = pi20 & ~n2793;
  assign n1133 = ~n1131 & ~n1132;
  assign n1134 = pi82 & ~n1133;
  assign n1135 = pi20 & n460;
  assign n1136 = ~pi71 & ~n291;
  assign n1137 = ~n291 & ~n472;
  assign n1138 = ~pi71 & n1137;
  assign n1139 = ~n472 & n1136;
  assign n1140 = ~n1135 & ~n2902;
  assign n1141 = ~n1134 & ~n1135;
  assign n1142 = ~n2902 & n1141;
  assign n1143 = ~n1134 & n1140;
  assign po35 = ~pi129 & ~n2903;
  assign n1145 = pi21 & ~pi54;
  assign n1146 = ~pi4 & pi19;
  assign n1147 = ~pi21 & n1146;
  assign n1148 = pi19 & ~pi21;
  assign n1149 = ~pi21 & pi54;
  assign n1150 = pi19 & n1149;
  assign n1151 = pi54 & n1148;
  assign n1152 = n580 & n2904;
  assign n1153 = n487 & n1147;
  assign n1154 = n517 & n580;
  assign n1155 = n580 & n642;
  assign n1156 = n517 & n1155;
  assign n1157 = n642 & n1154;
  assign n1158 = n2904 & n2906;
  assign n1159 = n931 & n2905;
  assign n1160 = n2820 & n2907;
  assign n1161 = ~n1145 & ~n1160;
  assign n1162 = ~pi129 & ~n1161;
  assign n1163 = ~pi3 & n1162;
  assign n1164 = n479 & ~n1161;
  assign n1165 = pi22 & ~pi54;
  assign n1166 = pi5 & ~pi14;
  assign n1167 = pi5 & n728;
  assign n1168 = pi5 & ~pi7;
  assign n1169 = n717 & n1168;
  assign n1170 = n592 & n1166;
  assign n1171 = n902 & n2909;
  assign n1172 = ~pi22 & n489;
  assign n1173 = n487 & n1172;
  assign n1174 = n2839 & n1173;
  assign n1175 = n501 & n717;
  assign n1176 = n2862 & n1168;
  assign n1177 = n1175 & n1176;
  assign n1178 = n1174 & n1177;
  assign n1179 = n979 & n2909;
  assign n1180 = n902 & n1179;
  assign n1181 = n2819 & n2909;
  assign n1182 = n2862 & n979;
  assign n1183 = n1181 & n1182;
  assign n1184 = n979 & n1171;
  assign n1185 = ~n1165 & ~n2910;
  assign n1186 = ~pi129 & ~n1185;
  assign n1187 = ~pi3 & n1186;
  assign n1188 = n479 & ~n1185;
  assign n1189 = n392 & n393;
  assign n1190 = n2778 & n1189;
  assign n1191 = n2781 & n2782;
  assign n1192 = pi82 & ~n2912;
  assign n1193 = pi63 & ~n291;
  assign n1194 = ~n291 & ~n1192;
  assign n1195 = pi63 & n1194;
  assign n1196 = ~n1192 & n1193;
  assign n1197 = ~pi24 & ~n2781;
  assign n1198 = pi24 & ~pi45;
  assign n1199 = n2780 & n1198;
  assign n1200 = ~n1197 & ~n1199;
  assign n1201 = pi82 & ~n1200;
  assign n1202 = pi82 & ~n2782;
  assign n1203 = ~pi24 & n291;
  assign n1204 = ~n1202 & n1203;
  assign n1205 = ~pi129 & ~n1204;
  assign n1206 = n291 & ~n1202;
  assign n1207 = ~n459 & ~n1206;
  assign n1208 = ~pi24 & ~n1207;
  assign n1209 = pi24 & pi82;
  assign n1210 = n294 & n1209;
  assign n1211 = n418 & n1210;
  assign n1212 = ~pi44 & pi82;
  assign n1213 = n1198 & n1212;
  assign n1214 = n350 & n1213;
  assign n1215 = pi24 & n1212;
  assign n1216 = n2769 & n1215;
  assign n1217 = n2766 & n1216;
  assign n1218 = n2769 & n1211;
  assign n1219 = ~pi129 & ~n2914;
  assign n1220 = ~n1208 & n1219;
  assign n1221 = ~n1201 & n1205;
  assign n1222 = ~n2913 & n1219;
  assign n1223 = ~n1208 & n1222;
  assign n1224 = ~n2913 & n2915;
  assign n1225 = ~pi53 & pi58;
  assign n1226 = pi53 & ~pi58;
  assign n1227 = ~n1225 & ~n1226;
  assign n1228 = ~pi96 & ~pi110;
  assign n1229 = ~pi85 & ~n1228;
  assign n1230 = pi85 & ~pi116;
  assign n1231 = pi100 & ~n1230;
  assign n1232 = pi85 & pi116;
  assign n1233 = ~pi85 & ~pi96;
  assign n1234 = ~pi85 & ~pi110;
  assign n1235 = ~pi96 & n1234;
  assign n1236 = ~pi110 & n1233;
  assign n1237 = ~n1232 & ~n2917;
  assign n1238 = pi100 & ~n1237;
  assign n1239 = ~n1229 & n1231;
  assign n1240 = pi25 & ~pi116;
  assign n1241 = pi85 & n1240;
  assign n1242 = pi25 & n1230;
  assign n1243 = ~n2918 & ~n2919;
  assign n1244 = ~pi26 & ~n1243;
  assign n1245 = ~pi39 & ~pi52;
  assign n1246 = ~pi51 & ~pi52;
  assign n1247 = ~pi39 & n1246;
  assign n1248 = ~pi51 & n1245;
  assign n1249 = pi116 & n2920;
  assign n1250 = ~pi85 & ~n1249;
  assign n1251 = pi26 & n1250;
  assign n1252 = ~pi25 & ~pi116;
  assign n1253 = n1251 & ~n1252;
  assign n1254 = ~n1244 & ~n1253;
  assign n1255 = ~pi27 & ~n1254;
  assign n1256 = ~pi26 & ~pi85;
  assign n1257 = ~n1240 & ~n1249;
  assign n1258 = pi27 & ~n1257;
  assign n1259 = pi27 & ~n2920;
  assign n1260 = ~pi95 & ~pi100;
  assign n1261 = ~pi97 & n1260;
  assign n1262 = ~pi110 & ~n1261;
  assign n1263 = pi25 & ~n1262;
  assign n1264 = ~n1259 & n1263;
  assign n1265 = ~n1258 & ~n1264;
  assign n1266 = n1256 & ~n1265;
  assign n1267 = pi26 & pi116;
  assign n1268 = ~n1263 & ~n1267;
  assign n1269 = ~n2920 & ~n1268;
  assign n1270 = pi26 & n1240;
  assign n1271 = ~n1269 & ~n1270;
  assign n1272 = ~pi85 & ~n1271;
  assign n1273 = ~n1244 & ~n1272;
  assign n1274 = ~pi27 & ~n1273;
  assign n1275 = n2920 & n1263;
  assign n1276 = ~n1258 & ~n1275;
  assign n1277 = n1256 & ~n1276;
  assign n1278 = ~n1274 & ~n1277;
  assign n1279 = ~n1255 & ~n1266;
  assign n1280 = ~pi53 & ~n2921;
  assign n1281 = n1227 & ~n1280;
  assign n1282 = ~pi53 & ~pi58;
  assign n1283 = ~pi26 & ~pi27;
  assign n1284 = ~pi85 & n1283;
  assign n1285 = pi25 & ~pi26;
  assign n1286 = ~pi116 & n1285;
  assign n1287 = ~pi26 & n1240;
  assign n1288 = ~pi27 & ~pi85;
  assign n1289 = n2922 & n1288;
  assign n1290 = n1240 & n1284;
  assign n1291 = ~n1282 & ~n2923;
  assign n1292 = n479 & ~n1291;
  assign n1293 = pi53 & ~pi85;
  assign n1294 = ~pi27 & n1293;
  assign n1295 = n2922 & n1294;
  assign n1296 = ~n1280 & ~n1295;
  assign n1297 = ~pi58 & ~n1296;
  assign n1298 = n1225 & n1288;
  assign n1299 = n2922 & n1298;
  assign n1300 = ~n1297 & ~n1299;
  assign n1301 = ~pi129 & ~n1300;
  assign n1302 = ~pi3 & n1301;
  assign n1303 = n479 & ~n1300;
  assign n1304 = ~n1281 & n1292;
  assign n1305 = ~pi26 & ~n2920;
  assign n1306 = ~pi27 & n2920;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1262 & ~n1307;
  assign n1309 = pi26 & pi27;
  assign n1310 = pi26 & ~pi27;
  assign n1311 = ~pi26 & pi27;
  assign n1312 = ~n1310 & ~n1311;
  assign n1313 = ~n1283 & ~n1309;
  assign n1314 = ~pi116 & ~n2925;
  assign n1315 = ~n1308 & ~n1314;
  assign n1316 = pi28 & ~n1315;
  assign n1317 = ~pi26 & pi95;
  assign n1318 = ~pi100 & n1317;
  assign n1319 = pi95 & ~pi96;
  assign n1320 = ~pi26 & ~pi100;
  assign n1321 = ~pi110 & n1320;
  assign n1322 = n1319 & n1321;
  assign n1323 = n1228 & n1318;
  assign n1324 = pi26 & n1249;
  assign n1325 = n2920 & n1267;
  assign n1326 = ~n2926 & ~n2927;
  assign n1327 = ~pi27 & ~n1326;
  assign n1328 = pi27 & pi116;
  assign n1329 = n1305 & n1328;
  assign n1330 = ~pi85 & ~n1329;
  assign n1331 = ~n1327 & n1330;
  assign n1332 = ~n1316 & n1331;
  assign n1333 = pi100 & pi116;
  assign n1334 = ~pi28 & ~pi116;
  assign n1335 = n1283 & ~n1334;
  assign n1336 = ~n1333 & n1335;
  assign n1337 = pi85 & ~n1336;
  assign n1338 = ~pi53 & ~n1337;
  assign n1339 = ~n1327 & ~n1329;
  assign n1340 = ~n1316 & n1339;
  assign n1341 = ~pi85 & ~n1340;
  assign n1342 = pi28 & ~pi116;
  assign n1343 = ~pi100 & pi116;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = pi85 & n1283;
  assign n1346 = pi85 & ~n1344;
  assign n1347 = n1283 & n1346;
  assign n1348 = ~n1344 & n1345;
  assign n1349 = ~n1341 & ~n2928;
  assign n1350 = ~pi53 & ~n1349;
  assign n1351 = ~n1332 & n1338;
  assign n1352 = pi53 & ~pi116;
  assign n1353 = ~pi27 & pi28;
  assign n1354 = n1256 & n1353;
  assign n1355 = ~pi116 & n1353;
  assign n1356 = pi53 & n1256;
  assign n1357 = ~pi26 & n1293;
  assign n1358 = n1355 & n2930;
  assign n1359 = n1352 & n1354;
  assign n1360 = ~n2929 & ~n2931;
  assign n1361 = ~pi58 & ~n1360;
  assign n1362 = ~pi26 & ~pi53;
  assign n1363 = ~pi85 & n1362;
  assign n1364 = pi58 & ~pi116;
  assign n1365 = pi58 & n1355;
  assign n1366 = n1353 & n1364;
  assign n1367 = n1225 & n1256;
  assign n1368 = n1355 & n1367;
  assign n1369 = n1363 & n2932;
  assign n1370 = ~n1361 & ~n2933;
  assign n1371 = ~pi129 & ~n1370;
  assign n1372 = ~pi3 & n1371;
  assign n1373 = n479 & ~n1370;
  assign n1374 = pi27 & n1250;
  assign n1375 = ~pi85 & pi95;
  assign n1376 = n1228 & n1375;
  assign n1377 = pi95 & ~n1230;
  assign n1378 = n1228 & n1377;
  assign n1379 = ~n1232 & ~n1378;
  assign n1380 = ~n1232 & ~n1376;
  assign n1381 = ~pi100 & ~n1328;
  assign n1382 = ~pi110 & ~n1230;
  assign n1383 = n1319 & ~n1328;
  assign n1384 = ~n1328 & n1382;
  assign n1385 = n1319 & n1384;
  assign n1386 = n1382 & n1383;
  assign n1387 = ~pi27 & n1232;
  assign n1388 = ~n2936 & ~n1387;
  assign n1389 = ~pi100 & ~n1388;
  assign n1390 = ~n2935 & n1381;
  assign n1391 = ~n1374 & ~n2937;
  assign n1392 = ~pi26 & n479;
  assign n1393 = ~pi26 & n1282;
  assign n1394 = n479 & n1393;
  assign n1395 = n1282 & n1392;
  assign n1396 = ~pi129 & ~n1391;
  assign n1397 = ~pi3 & n1396;
  assign n1398 = n1393 & n1397;
  assign n1399 = ~n1391 & n2938;
  assign n1400 = ~pi96 & ~n1267;
  assign n1401 = ~n1267 & n1382;
  assign n1402 = ~pi96 & n1401;
  assign n1403 = n1382 & n1400;
  assign n1404 = ~pi26 & n1232;
  assign n1405 = ~n2940 & ~n1404;
  assign n1406 = pi100 & ~n1405;
  assign n1407 = n2918 & ~n1267;
  assign n1408 = ~n1251 & ~n2941;
  assign n1409 = ~pi27 & ~pi53;
  assign n1410 = ~pi58 & n1409;
  assign n1411 = n479 & n1410;
  assign n1412 = ~pi129 & ~n1408;
  assign n1413 = ~pi3 & n1412;
  assign n1414 = n1410 & n1413;
  assign n1415 = ~n1408 & n1411;
  assign n1416 = pi97 & ~n1228;
  assign n1417 = ~pi29 & ~pi97;
  assign n1418 = n1260 & ~n1417;
  assign n1419 = ~pi96 & pi97;
  assign n1420 = pi97 & ~pi110;
  assign n1421 = ~pi96 & n1420;
  assign n1422 = pi97 & n1228;
  assign n1423 = ~pi110 & n1419;
  assign n1424 = pi29 & ~pi97;
  assign n1425 = ~n2943 & ~n1424;
  assign n1426 = n1260 & ~n1425;
  assign n1427 = ~n1416 & n1418;
  assign n1428 = pi29 & pi110;
  assign n1429 = ~pi58 & ~n1428;
  assign n1430 = pi29 & ~n1262;
  assign n1431 = n1228 & n1260;
  assign n1432 = n1260 & n2943;
  assign n1433 = pi97 & n1431;
  assign n1434 = ~pi58 & ~n2945;
  assign n1435 = ~n1430 & n1434;
  assign n1436 = ~n2944 & n1429;
  assign n1437 = pi97 & pi116;
  assign n1438 = pi29 & ~pi116;
  assign n1439 = pi58 & ~n1438;
  assign n1440 = pi58 & ~n1437;
  assign n1441 = ~n1438 & n1440;
  assign n1442 = ~n1437 & n1439;
  assign n1443 = ~pi53 & ~n2947;
  assign n1444 = ~n2944 & ~n1428;
  assign n1445 = ~pi58 & ~n1444;
  assign n1446 = ~n1437 & ~n1438;
  assign n1447 = pi58 & ~n1446;
  assign n1448 = ~n1445 & ~n1447;
  assign n1449 = ~pi53 & ~n1448;
  assign n1450 = ~n2946 & n1443;
  assign n1451 = n1226 & n1438;
  assign n1452 = ~n2948 & ~n1451;
  assign n1453 = ~pi27 & ~n1452;
  assign n1454 = pi27 & n1282;
  assign n1455 = pi27 & n1438;
  assign n1456 = n1282 & n1455;
  assign n1457 = n1438 & n1454;
  assign n1458 = ~n1453 & ~n2949;
  assign n1459 = ~pi85 & ~n1458;
  assign n1460 = pi85 & n1438;
  assign n1461 = pi85 & n1410;
  assign n1462 = n1438 & n1461;
  assign n1463 = n1410 & n1460;
  assign n1464 = ~n1459 & ~n2950;
  assign n1465 = ~pi26 & ~n1464;
  assign n1466 = pi26 & n1288;
  assign n1467 = ~pi85 & n1310;
  assign n1468 = n1282 & n1288;
  assign n1469 = pi26 & n1468;
  assign n1470 = pi26 & n1282;
  assign n1471 = n1288 & n1470;
  assign n1472 = ~pi85 & n1282;
  assign n1473 = n1310 & n1472;
  assign n1474 = n1282 & n2951;
  assign n1475 = n1438 & n2952;
  assign n1476 = ~n1465 & ~n1475;
  assign n1477 = ~pi129 & ~n1476;
  assign n1478 = ~pi3 & n1477;
  assign n1479 = n479 & ~n1476;
  assign n1480 = pi82 & ~n295;
  assign n1481 = ~pi43 & n2790;
  assign n1482 = n2771 & n2788;
  assign n1483 = n314 & n2789;
  assign n1484 = n310 & n2954;
  assign n1485 = n393 & n394;
  assign n1486 = n311 & n404;
  assign n1487 = n1485 & n1486;
  assign n1488 = n315 & n2789;
  assign n1489 = n2772 & n2788;
  assign n1490 = ~pi50 & n2955;
  assign n1491 = n2773 & n2788;
  assign n1492 = pi82 & ~n2956;
  assign n1493 = n291 & ~n1492;
  assign n1494 = ~n1480 & ~n1493;
  assign n1495 = ~pi38 & ~n1494;
  assign n1496 = n295 & n2770;
  assign n1497 = n2954 & n1496;
  assign n1498 = ~pi41 & n2954;
  assign n1499 = n339 & n2789;
  assign n1500 = n338 & n2790;
  assign n1501 = n334 & n2958;
  assign n1502 = ~pi50 & n295;
  assign n1503 = n315 & n1502;
  assign n1504 = n2789 & n1503;
  assign n1505 = n295 & n2956;
  assign n1506 = pi82 & ~n2957;
  assign n1507 = pi74 & ~n291;
  assign n1508 = ~n291 & ~n1506;
  assign n1509 = pi74 & n1508;
  assign n1510 = ~n1506 & n1507;
  assign n1511 = pi38 & pi82;
  assign n1512 = ~pi42 & n1212;
  assign n1513 = ~pi40 & n1512;
  assign n1514 = n296 & n1212;
  assign n1515 = pi38 & n2960;
  assign n1516 = pi38 & n296;
  assign n1517 = n1212 & n1516;
  assign n1518 = n295 & n1511;
  assign n1519 = ~pi129 & ~n2961;
  assign n1520 = ~n2959 & n1519;
  assign po53 = ~n1495 & n1520;
  assign n1522 = pi82 & ~n294;
  assign n1523 = n2786 & n2954;
  assign n1524 = n2774 & n2958;
  assign n1525 = pi82 & ~n2962;
  assign n1526 = n291 & ~n1525;
  assign n1527 = ~n1522 & ~n1526;
  assign n1528 = ~pi40 & ~n1527;
  assign n1529 = n293 & n294;
  assign n1530 = n315 & n1529;
  assign n1531 = n294 & n2962;
  assign n1532 = n294 & n2774;
  assign n1533 = n2958 & n1532;
  assign n1534 = n2789 & n1530;
  assign n1535 = pi82 & ~n2963;
  assign n1536 = pi73 & ~n291;
  assign n1537 = ~n291 & ~n1535;
  assign n1538 = pi73 & n1537;
  assign n1539 = ~n1535 & n1536;
  assign n1540 = pi40 & pi82;
  assign n1541 = pi40 & n1512;
  assign n1542 = n294 & n1540;
  assign n1543 = ~pi129 & ~n2965;
  assign n1544 = ~n2964 & n1543;
  assign po55 = ~n1528 & n1544;
  assign n1546 = pi82 & ~n2776;
  assign n1547 = pi82 & ~n2954;
  assign n1548 = n291 & ~n1547;
  assign n1549 = ~n1546 & ~n1548;
  assign n1550 = ~pi41 & ~n1549;
  assign n1551 = n314 & n319;
  assign n1552 = n314 & n2776;
  assign n1553 = n307 & n1551;
  assign n1554 = n2776 & n2954;
  assign n1555 = n2789 & n2966;
  assign n1556 = pi82 & ~n2967;
  assign n1557 = pi76 & ~n291;
  assign n1558 = ~n291 & ~n1556;
  assign n1559 = pi76 & n1558;
  assign n1560 = ~n1556 & n1557;
  assign n1561 = pi41 & pi82;
  assign n1562 = pi41 & n1512;
  assign n1563 = n294 & n1561;
  assign n1564 = ~pi40 & pi41;
  assign n1565 = n2774 & n1564;
  assign n1566 = n1512 & n1565;
  assign n1567 = n2775 & n2969;
  assign n1568 = ~pi129 & ~n2970;
  assign n1569 = ~n2968 & n1568;
  assign n1570 = ~n1550 & n1568;
  assign n1571 = ~n2968 & n1570;
  assign n1572 = ~n1550 & n1569;
  assign n1573 = n2775 & n339;
  assign n1574 = ~pi40 & n2962;
  assign n1575 = n2775 & n2958;
  assign n1576 = n2789 & n1573;
  assign n1577 = pi82 & ~n2972;
  assign n1578 = ~pi72 & ~n291;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = ~n1522 & ~n1579;
  assign n1581 = pi42 & ~n1212;
  assign n1582 = ~n292 & n1581;
  assign n1583 = ~n1580 & ~n1582;
  assign n1584 = pi44 & pi82;
  assign n1585 = n291 & ~n1577;
  assign n1586 = ~n1584 & ~n1585;
  assign n1587 = ~pi42 & ~n1586;
  assign n1588 = n315 & n433;
  assign n1589 = n2789 & n1588;
  assign n1590 = ~pi44 & n2972;
  assign n1591 = n433 & n2955;
  assign n1592 = pi82 & ~n2973;
  assign n1593 = pi72 & ~n291;
  assign n1594 = ~n291 & ~n1592;
  assign n1595 = pi72 & n1594;
  assign n1596 = ~n1592 & n1593;
  assign n1597 = pi42 & n1212;
  assign n1598 = ~pi129 & ~n1597;
  assign n1599 = ~n2974 & n1598;
  assign n1600 = ~n1587 & n1599;
  assign n1601 = ~pi129 & ~n1583;
  assign n1602 = pi82 & ~n2777;
  assign n1603 = pi82 & ~n2790;
  assign n1604 = n291 & ~n1603;
  assign n1605 = ~n1602 & ~n1604;
  assign n1606 = ~pi43 & ~n1605;
  assign n1607 = ~pi47 & n2777;
  assign n1608 = n2789 & n1607;
  assign n1609 = n2777 & n2790;
  assign n1610 = pi82 & ~n2976;
  assign n1611 = pi77 & ~n291;
  assign n1612 = ~n291 & ~n1610;
  assign n1613 = pi77 & n1612;
  assign n1614 = ~n1610 & n1611;
  assign n1615 = n2786 & n2960;
  assign n1616 = pi82 & n2776;
  assign n1617 = ~pi41 & pi43;
  assign n1618 = n1616 & n1617;
  assign n1619 = pi43 & n296;
  assign n1620 = pi43 & n2960;
  assign n1621 = n1212 & n1619;
  assign n1622 = n2786 & n2979;
  assign n1623 = pi43 & n1615;
  assign n1624 = ~pi129 & ~n2978;
  assign n1625 = ~n2977 & n1624;
  assign n1626 = ~n1606 & n1624;
  assign n1627 = ~n2977 & n1626;
  assign n1628 = ~n1606 & n1625;
  assign n1629 = ~pi42 & n2972;
  assign n1630 = n353 & n2789;
  assign n1631 = pi82 & ~n2981;
  assign n1632 = ~pi67 & ~n291;
  assign n1633 = pi44 & n291;
  assign n1634 = pi67 & ~n291;
  assign n1635 = ~pi44 & n291;
  assign n1636 = ~n1634 & ~n1635;
  assign n1637 = ~n1632 & ~n1633;
  assign n1638 = ~n1631 & ~n2982;
  assign n1639 = ~pi129 & ~n1584;
  assign po59 = ~n1638 & n1639;
  assign n1641 = ~pi48 & n2783;
  assign n1642 = n2779 & n1641;
  assign n1643 = n2778 & n405;
  assign n1644 = n2780 & n2783;
  assign n1645 = pi82 & ~n2983;
  assign n1646 = pi68 & ~n291;
  assign n1647 = ~n291 & ~n1645;
  assign n1648 = pi68 & n1647;
  assign n1649 = ~n1645 & n1646;
  assign n1650 = pi82 & ~n2783;
  assign n1651 = n291 & ~n1650;
  assign n1652 = pi82 & ~n2780;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = ~pi45 & ~n1653;
  assign n1655 = pi45 & n1212;
  assign n1656 = pi45 & n2767;
  assign n1657 = n1212 & n1656;
  assign n1658 = n2767 & n1655;
  assign n1659 = pi45 & pi82;
  assign n1660 = n2780 & n1659;
  assign n1661 = n2773 & n2985;
  assign n1662 = ~pi129 & ~n2986;
  assign n1663 = ~n1654 & n1662;
  assign n1664 = ~n2984 & n1662;
  assign n1665 = ~n1654 & n1664;
  assign n1666 = ~n2984 & n1663;
  assign n1667 = ~pi75 & ~n291;
  assign n1668 = pi82 & ~n2958;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = n2776 & ~n1669;
  assign n1671 = pi82 & ~n2768;
  assign n1672 = ~n460 & ~n1671;
  assign n1673 = pi46 & ~n1672;
  assign n1674 = ~pi82 & n1667;
  assign n1675 = ~n1673 & ~n1674;
  assign n1676 = ~n1670 & n1675;
  assign n1677 = n291 & ~n1668;
  assign n1678 = ~n1671 & ~n1677;
  assign n1679 = ~pi46 & ~n1678;
  assign n1680 = n2768 & n2958;
  assign n1681 = pi82 & ~n1680;
  assign n1682 = pi75 & ~n291;
  assign n1683 = ~n291 & ~n1681;
  assign n1684 = pi75 & n1683;
  assign n1685 = ~n1681 & n1682;
  assign n1686 = pi46 & n1212;
  assign n1687 = pi46 & pi82;
  assign n1688 = n2768 & n1687;
  assign n1689 = n2766 & n1686;
  assign n1690 = ~pi129 & ~n2989;
  assign n1691 = ~n2988 & n1690;
  assign n1692 = ~n1679 & n1691;
  assign n1693 = ~pi129 & ~n1676;
  assign n1694 = pi82 & ~n2778;
  assign n1695 = pi82 & ~n2789;
  assign n1696 = n291 & ~n1695;
  assign n1697 = ~n1694 & ~n1696;
  assign n1698 = ~pi47 & ~n1697;
  assign n1699 = n2778 & n2789;
  assign n1700 = pi82 & ~n1699;
  assign n1701 = pi64 & ~n291;
  assign n1702 = ~n291 & ~n1700;
  assign n1703 = pi64 & n1702;
  assign n1704 = ~n1700 & n1701;
  assign n1705 = n2774 & n338;
  assign n1706 = pi47 & n296;
  assign n1707 = n1212 & n1706;
  assign n1708 = pi47 & n338;
  assign n1709 = n1616 & n1708;
  assign n1710 = ~pi43 & pi47;
  assign n1711 = n1615 & n1710;
  assign n1712 = n2774 & n1708;
  assign n1713 = n2960 & n1712;
  assign n1714 = n2960 & n1708;
  assign n1715 = n2774 & n1714;
  assign n1716 = n1705 & n1707;
  assign n1717 = ~pi129 & ~n2992;
  assign n1718 = ~n2991 & n1717;
  assign n1719 = ~n1698 & n1717;
  assign n1720 = ~n2991 & n1719;
  assign n1721 = ~n1698 & n1718;
  assign n1722 = ~pi2 & ~pi47;
  assign n1723 = n1485 & n1722;
  assign n1724 = n2778 & n1723;
  assign n1725 = n2779 & n2788;
  assign n1726 = pi82 & ~n2994;
  assign n1727 = pi62 & ~n291;
  assign n1728 = ~n291 & ~n1726;
  assign n1729 = pi62 & n1728;
  assign n1730 = ~n1726 & n1727;
  assign n1731 = pi82 & ~n2788;
  assign n1732 = n291 & ~n1731;
  assign n1733 = pi82 & ~n2779;
  assign n1734 = ~n1732 & ~n1733;
  assign n1735 = ~pi48 & ~n1734;
  assign n1736 = pi48 & n1212;
  assign n1737 = n314 & n2770;
  assign n1738 = pi48 & n2767;
  assign n1739 = n1212 & n1738;
  assign n1740 = n1737 & n1739;
  assign n1741 = n2766 & n1736;
  assign n1742 = n315 & n1741;
  assign n1743 = pi48 & n314;
  assign n1744 = n1212 & n1743;
  assign n1745 = n2767 & n2770;
  assign n1746 = n1744 & n1745;
  assign n1747 = n353 & n1736;
  assign n1748 = ~pi129 & ~n2996;
  assign n1749 = ~n1735 & n1748;
  assign n1750 = ~n2995 & n1748;
  assign n1751 = ~n1735 & n1750;
  assign n1752 = ~n2995 & n1749;
  assign n1753 = pi49 & ~n2798;
  assign n1754 = ~n2797 & ~n1753;
  assign n1755 = n2769 & ~n366;
  assign n1756 = ~n366 & n443;
  assign n1757 = n315 & n1756;
  assign n1758 = n316 & n1757;
  assign n1759 = ~n366 & n2797;
  assign n1760 = n443 & n1755;
  assign n1761 = ~n1753 & ~n2998;
  assign n1762 = pi82 & ~n1761;
  assign n1763 = n1202 & ~n1754;
  assign n1764 = pi49 & n460;
  assign n1765 = pi82 & ~n2797;
  assign n1766 = ~pi69 & ~n291;
  assign n1767 = ~n291 & ~n1765;
  assign n1768 = ~pi69 & n1767;
  assign n1769 = ~n1765 & n1766;
  assign n1770 = ~n1764 & ~n3000;
  assign n1771 = ~n2999 & ~n1764;
  assign n1772 = ~n3000 & n1771;
  assign n1773 = ~n2999 & n1770;
  assign po64 = ~pi129 & ~n3001;
  assign n1775 = ~n460 & ~n1511;
  assign n1776 = ~n1480 & n1775;
  assign n1777 = pi50 & ~n1776;
  assign n1778 = ~pi66 & ~n291;
  assign n1779 = pi82 & ~n2955;
  assign n1780 = ~n1778 & ~n1779;
  assign n1781 = ~n1671 & ~n1780;
  assign n1782 = ~n1777 & ~n1781;
  assign n1783 = n307 & n315;
  assign n1784 = n295 & n328;
  assign n1785 = n2958 & n1784;
  assign n1786 = n2789 & n1783;
  assign n1787 = pi82 & ~n3002;
  assign n1788 = pi66 & ~n291;
  assign n1789 = ~n291 & ~n1787;
  assign n1790 = pi66 & n1789;
  assign n1791 = ~n1787 & n1788;
  assign n1792 = pi82 & ~n307;
  assign n1793 = n291 & ~n1779;
  assign n1794 = ~n1792 & ~n1793;
  assign n1795 = ~pi50 & ~n1794;
  assign n1796 = pi50 & n1212;
  assign n1797 = pi50 & n2767;
  assign n1798 = n1212 & n1797;
  assign n1799 = pi50 & pi82;
  assign n1800 = n307 & n1799;
  assign n1801 = n2767 & n1796;
  assign n1802 = ~pi129 & ~n3004;
  assign n1803 = ~n1795 & n1802;
  assign n1804 = ~n3003 & n1803;
  assign n1805 = ~n3003 & n1802;
  assign n1806 = ~n1795 & n1805;
  assign n1807 = ~pi129 & ~n1782;
  assign n1808 = ~pi129 & ~n2791;
  assign n1809 = pi59 & ~pi116;
  assign n1810 = ~n1227 & n1809;
  assign n1811 = ~pi96 & n1262;
  assign n1812 = ~pi59 & ~n1262;
  assign n1813 = n1282 & ~n1812;
  assign n1814 = ~n1811 & n1813;
  assign n1815 = ~pi116 & ~n1227;
  assign n1816 = ~n1262 & n1282;
  assign n1817 = ~n1815 & ~n1816;
  assign n1818 = pi59 & ~n1817;
  assign n1819 = pi96 & n1282;
  assign n1820 = n1262 & n1282;
  assign n1821 = pi96 & n1820;
  assign n1822 = n1262 & n1819;
  assign n1823 = ~n1818 & ~n3006;
  assign n1824 = ~n1810 & ~n1814;
  assign n1825 = ~pi85 & ~n3007;
  assign n1826 = pi85 & n1282;
  assign n1827 = n1809 & n1826;
  assign n1828 = ~n1825 & ~n1827;
  assign n1829 = ~pi27 & ~n1828;
  assign n1830 = ~pi85 & n1809;
  assign n1831 = pi27 & n1472;
  assign n1832 = n1809 & n1831;
  assign n1833 = pi27 & n1809;
  assign n1834 = n1472 & n1833;
  assign n1835 = n1454 & n1830;
  assign n1836 = ~n1829 & ~n3008;
  assign n1837 = ~pi26 & ~n1836;
  assign n1838 = n2952 & n1809;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = ~pi129 & ~n1839;
  assign n1841 = ~pi3 & n1840;
  assign n1842 = n479 & ~n1839;
  assign n1843 = ~pi58 & ~n1431;
  assign n1844 = ~pi53 & pi97;
  assign n1845 = ~n1843 & n1844;
  assign n1846 = ~n1352 & ~n1845;
  assign n1847 = n479 & ~n1364;
  assign n1848 = n1284 & n1847;
  assign n1849 = pi58 & pi116;
  assign n1850 = ~pi58 & ~pi96;
  assign n1851 = ~pi58 & ~pi110;
  assign n1852 = ~pi96 & n1851;
  assign n1853 = ~pi58 & n1228;
  assign n1854 = ~pi110 & n1850;
  assign n1855 = n1260 & n3010;
  assign n1856 = ~n1849 & ~n1855;
  assign n1857 = ~pi53 & ~n1856;
  assign n1858 = pi97 & n1857;
  assign n1859 = n1844 & ~n1856;
  assign n1860 = ~pi116 & n1226;
  assign n1861 = ~n3011 & ~n1860;
  assign n1862 = ~pi129 & ~n1861;
  assign n1863 = ~pi3 & n1862;
  assign n1864 = n1288 & n1863;
  assign n1865 = ~pi26 & n1864;
  assign n1866 = n1288 & n1392;
  assign n1867 = ~n1861 & n1866;
  assign n1868 = ~n1846 & n1848;
  assign n1869 = ~pi85 & n1262;
  assign n1870 = ~pi85 & ~n1261;
  assign n1871 = ~pi110 & n1870;
  assign n1872 = n1234 & ~n1261;
  assign n1873 = pi96 & n3013;
  assign n1874 = ~n1230 & ~n1873;
  assign n1875 = n1392 & n1410;
  assign n1876 = ~pi129 & ~n1874;
  assign n1877 = ~pi3 & n1876;
  assign n1878 = n1410 & n1877;
  assign n1879 = ~pi26 & n1878;
  assign n1880 = ~n1874 & n1875;
  assign n1881 = pi131 & pi132;
  assign n1882 = pi132 & pi133;
  assign n1883 = pi131 & n1882;
  assign n1884 = pi133 & n1881;
  assign n1885 = ~pi136 & ~pi137;
  assign n1886 = pi82 & pi138;
  assign n1887 = pi82 & ~pi136;
  assign n1888 = ~pi137 & pi138;
  assign n1889 = n1887 & n1888;
  assign n1890 = pi82 & ~pi137;
  assign n1891 = ~pi136 & n1890;
  assign n1892 = ~pi137 & n1887;
  assign n1893 = pi138 & n3017;
  assign n1894 = n1885 & n1886;
  assign n1895 = pi138 & n3015;
  assign n1896 = n3017 & n1895;
  assign n1897 = n3015 & n3016;
  assign n1898 = ~pi3 & ~pi110;
  assign n1899 = ~n3015 & ~n1898;
  assign n1900 = ~pi3 & ~n3015;
  assign n1901 = ~pi110 & n1900;
  assign n1902 = ~n3015 & n1898;
  assign n1903 = n3015 & ~n3016;
  assign n1904 = ~n3019 & ~n1903;
  assign n1905 = ~n3018 & ~n1899;
  assign n1906 = pi95 & ~n3020;
  assign n1907 = pi143 & n3018;
  assign n1908 = ~n1906 & ~n1907;
  assign po110 = ~pi129 & ~n1908;
  assign n1910 = pi96 & ~n3020;
  assign n1911 = pi146 & n3018;
  assign n1912 = ~n1910 & ~n1911;
  assign po111 = ~pi129 & ~n1912;
  assign n1914 = pi97 & ~n3020;
  assign n1915 = pi145 & n3018;
  assign n1916 = ~n1914 & ~n1915;
  assign po112 = ~pi129 & ~n1916;
  assign n1918 = pi100 & ~n3020;
  assign n1919 = pi144 & n3018;
  assign n1920 = ~n1918 & ~n1919;
  assign po115 = ~pi129 & ~n1920;
  assign n1922 = pi136 & ~pi137;
  assign n1923 = pi99 & n1922;
  assign n1924 = ~pi136 & pi137;
  assign n1925 = ~pi112 & n1924;
  assign n1926 = ~n1923 & ~n1925;
  assign n1927 = pi138 & ~n1926;
  assign n1928 = ~pi32 & pi136;
  assign n1929 = ~pi84 & ~pi136;
  assign n1930 = pi137 & ~n1929;
  assign n1931 = pi84 & ~pi136;
  assign n1932 = pi32 & pi136;
  assign n1933 = ~n1931 & ~n1932;
  assign n1934 = pi137 & ~n1933;
  assign n1935 = ~n1928 & n1930;
  assign n1936 = pi68 & pi136;
  assign n1937 = pi73 & ~pi136;
  assign n1938 = ~pi137 & ~n1937;
  assign n1939 = ~pi68 & pi136;
  assign n1940 = ~pi73 & ~pi136;
  assign n1941 = ~n1939 & ~n1940;
  assign n1942 = ~pi137 & ~n1941;
  assign n1943 = ~n1936 & n1938;
  assign n1944 = ~n3021 & ~n3022;
  assign n1945 = ~pi138 & ~n1944;
  assign n1946 = ~n1927 & ~n1945;
  assign n1947 = ~pi30 & ~pi109;
  assign n1948 = ~pi60 & pi109;
  assign n1949 = pi30 & ~pi109;
  assign n1950 = pi60 & pi109;
  assign n1951 = ~n1949 & ~n1950;
  assign n1952 = ~n1947 & ~n1948;
  assign n1953 = ~pi106 & ~n1949;
  assign n1954 = ~n1950 & n1953;
  assign n1955 = ~pi106 & n3023;
  assign n1956 = ~pi88 & pi106;
  assign n1957 = ~pi129 & ~n1956;
  assign n1958 = ~pi106 & ~n3023;
  assign n1959 = pi88 & pi106;
  assign n1960 = ~n1958 & ~n1959;
  assign n1961 = ~pi129 & ~n1960;
  assign n1962 = ~n3024 & n1957;
  assign n1963 = ~pi31 & ~pi109;
  assign n1964 = ~pi30 & pi109;
  assign n1965 = pi30 & pi109;
  assign n1966 = pi31 & ~pi109;
  assign n1967 = ~n1965 & ~n1966;
  assign n1968 = ~n1963 & ~n1964;
  assign n1969 = ~pi106 & ~n1966;
  assign n1970 = ~n1965 & n1969;
  assign n1971 = ~pi106 & n3026;
  assign n1972 = ~pi89 & pi106;
  assign n1973 = ~pi129 & ~n1972;
  assign n1974 = pi89 & pi106;
  assign n1975 = ~pi106 & ~n3026;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = ~pi129 & ~n1976;
  assign n1978 = ~n3027 & n1973;
  assign n1979 = ~pi32 & ~pi109;
  assign n1980 = ~pi31 & pi109;
  assign n1981 = pi31 & pi109;
  assign n1982 = pi32 & ~pi109;
  assign n1983 = ~n1981 & ~n1982;
  assign n1984 = ~n1979 & ~n1980;
  assign n1985 = ~pi106 & ~n1982;
  assign n1986 = ~n1981 & n1985;
  assign n1987 = ~pi106 & n3029;
  assign n1988 = ~pi99 & pi106;
  assign n1989 = ~pi129 & ~n1988;
  assign n1990 = pi99 & pi106;
  assign n1991 = ~pi106 & ~n3029;
  assign n1992 = ~n1990 & ~n1991;
  assign n1993 = ~pi129 & ~n1992;
  assign n1994 = ~n3030 & n1989;
  assign n1995 = ~pi33 & ~pi109;
  assign n1996 = ~pi32 & pi109;
  assign n1997 = pi32 & pi109;
  assign n1998 = pi33 & ~pi109;
  assign n1999 = ~n1997 & ~n1998;
  assign n2000 = ~n1995 & ~n1996;
  assign n2001 = ~pi106 & ~n1998;
  assign n2002 = ~n1997 & n2001;
  assign n2003 = ~pi106 & n3032;
  assign n2004 = ~pi90 & pi106;
  assign n2005 = ~pi129 & ~n2004;
  assign n2006 = pi90 & pi106;
  assign n2007 = ~pi106 & ~n3032;
  assign n2008 = ~n2006 & ~n2007;
  assign n2009 = ~pi129 & ~n2008;
  assign n2010 = ~n3033 & n2005;
  assign n2011 = ~pi34 & ~pi109;
  assign n2012 = ~pi33 & pi109;
  assign n2013 = pi33 & pi109;
  assign n2014 = pi34 & ~pi109;
  assign n2015 = ~n2013 & ~n2014;
  assign n2016 = ~n2011 & ~n2012;
  assign n2017 = ~pi106 & ~n2014;
  assign n2018 = ~n2013 & n2017;
  assign n2019 = ~pi106 & n3035;
  assign n2020 = ~pi91 & pi106;
  assign n2021 = ~pi129 & ~n2020;
  assign n2022 = pi91 & pi106;
  assign n2023 = ~pi106 & ~n3035;
  assign n2024 = ~n2022 & ~n2023;
  assign n2025 = ~pi129 & ~n2024;
  assign n2026 = ~n3036 & n2021;
  assign n2027 = ~pi35 & ~pi109;
  assign n2028 = ~pi34 & pi109;
  assign n2029 = pi34 & pi109;
  assign n2030 = pi35 & ~pi109;
  assign n2031 = ~n2029 & ~n2030;
  assign n2032 = ~n2027 & ~n2028;
  assign n2033 = ~pi106 & ~n2030;
  assign n2034 = ~n2029 & n2033;
  assign n2035 = ~pi106 & n3038;
  assign n2036 = ~pi92 & pi106;
  assign n2037 = ~pi129 & ~n2036;
  assign n2038 = pi92 & pi106;
  assign n2039 = ~pi106 & ~n3038;
  assign n2040 = ~n2038 & ~n2039;
  assign n2041 = ~pi129 & ~n2040;
  assign n2042 = ~n3039 & n2037;
  assign n2043 = ~pi36 & ~pi109;
  assign n2044 = ~pi35 & pi109;
  assign n2045 = pi35 & pi109;
  assign n2046 = pi36 & ~pi109;
  assign n2047 = ~n2045 & ~n2046;
  assign n2048 = ~n2043 & ~n2044;
  assign n2049 = ~pi106 & ~n2046;
  assign n2050 = ~n2045 & n2049;
  assign n2051 = ~pi106 & n3041;
  assign n2052 = ~pi98 & pi106;
  assign n2053 = ~pi129 & ~n2052;
  assign n2054 = pi98 & pi106;
  assign n2055 = ~pi106 & ~n3041;
  assign n2056 = ~n2054 & ~n2055;
  assign n2057 = ~pi129 & ~n2056;
  assign n2058 = ~n3042 & n2053;
  assign n2059 = ~pi37 & ~pi109;
  assign n2060 = ~pi36 & pi109;
  assign n2061 = pi36 & pi109;
  assign n2062 = pi37 & ~pi109;
  assign n2063 = ~n2061 & ~n2062;
  assign n2064 = ~n2059 & ~n2060;
  assign n2065 = ~pi106 & ~n2062;
  assign n2066 = ~n2061 & n2065;
  assign n2067 = ~pi106 & n3044;
  assign n2068 = ~pi93 & pi106;
  assign n2069 = ~pi129 & ~n2068;
  assign n2070 = pi93 & pi106;
  assign n2071 = ~pi106 & ~n3044;
  assign n2072 = ~n2070 & ~n2071;
  assign n2073 = ~pi129 & ~n2072;
  assign n2074 = ~n3045 & n2069;
  assign n2075 = pi109 & n1246;
  assign n2076 = pi39 & ~n2075;
  assign n2077 = ~pi51 & pi109;
  assign n2078 = n1245 & n2077;
  assign n2079 = ~pi106 & ~n2078;
  assign n2080 = ~n2076 & n2079;
  assign po54 = ~pi129 & ~n2080;
  assign n2082 = pi52 & ~n2077;
  assign n2083 = ~pi106 & ~n2075;
  assign n2084 = ~n2082 & n2083;
  assign po67 = ~pi129 & ~n2084;
  assign n2086 = ~pi23 & pi55;
  assign n2087 = pi61 & ~pi129;
  assign n2088 = ~pi129 & ~n2086;
  assign n2089 = pi61 & n2088;
  assign n2090 = ~n2086 & n2087;
  assign n2091 = pi51 & ~pi109;
  assign n2092 = ~pi106 & ~n2077;
  assign n2093 = ~n2077 & ~n2091;
  assign n2094 = ~pi106 & n2093;
  assign n2095 = ~n2091 & n2092;
  assign po66 = ~pi129 & ~n3048;
  assign n2097 = ~pi123 & ~pi129;
  assign n2098 = pi114 & ~pi122;
  assign po70 = n2097 & n2098;
  assign n2100 = ~pi117 & ~pi122;
  assign n2101 = pi60 & ~n2100;
  assign n2102 = pi123 & n2100;
  assign n2103 = ~n2101 & ~n2102;
  assign n2104 = ~pi114 & ~pi122;
  assign n2105 = pi123 & ~pi129;
  assign n2106 = ~pi114 & pi123;
  assign n2107 = ~pi122 & n2106;
  assign n2108 = ~pi129 & n2107;
  assign n2109 = n2104 & n2105;
  assign n2110 = ~pi27 & n1393;
  assign n2111 = ~pi26 & n1410;
  assign n2112 = n1393 & n3013;
  assign n2113 = ~pi27 & n2112;
  assign n2114 = n3013 & n3050;
  assign n2115 = ~n1232 & ~n3051;
  assign n2116 = ~pi129 & ~n2115;
  assign n2117 = ~pi3 & n2116;
  assign n2118 = n479 & ~n2115;
  assign n2119 = n1283 & n1364;
  assign n2120 = ~pi58 & ~n2925;
  assign n2121 = pi116 & ~n2925;
  assign n2122 = ~pi58 & n2121;
  assign n2123 = n2920 & n2122;
  assign n2124 = ~pi58 & pi116;
  assign n2125 = n2920 & n2124;
  assign n2126 = ~n2925 & n2125;
  assign n2127 = n1249 & n2120;
  assign n2128 = ~n2119 & ~n3053;
  assign n2129 = ~pi53 & ~pi85;
  assign n2130 = n479 & n2129;
  assign n2131 = ~pi129 & ~n2128;
  assign n2132 = ~pi3 & n2131;
  assign n2133 = ~pi53 & n2132;
  assign n2134 = ~pi85 & n2133;
  assign n2135 = ~n2128 & n2130;
  assign n2136 = ~pi26 & pi37;
  assign n2137 = n1282 & n2136;
  assign n2138 = ~pi26 & pi58;
  assign n2139 = pi26 & ~pi58;
  assign n2140 = pi116 & n2139;
  assign n2141 = ~pi58 & n1267;
  assign n2142 = ~n2138 & ~n3055;
  assign n2143 = pi94 & ~n2142;
  assign n2144 = pi37 & ~pi116;
  assign n2145 = ~n2138 & ~n2144;
  assign n2146 = ~n1364 & ~n2145;
  assign n2147 = ~n2143 & ~n2146;
  assign n2148 = ~pi53 & ~n2147;
  assign n2149 = ~pi58 & n2136;
  assign n2150 = ~n2148 & ~n2149;
  assign n2151 = ~pi85 & ~n2150;
  assign n2152 = ~n2137 & ~n2151;
  assign n2153 = n1472 & n2136;
  assign n2154 = ~pi85 & n2137;
  assign n2155 = pi27 & ~n3056;
  assign n2156 = n479 & ~n2155;
  assign n2157 = ~pi27 & ~n2152;
  assign n2158 = ~n3056 & ~n2157;
  assign n2159 = ~pi129 & ~n2158;
  assign n2160 = ~pi3 & n2159;
  assign n2161 = n479 & ~n2158;
  assign n2162 = ~n2152 & n2156;
  assign n2163 = ~pi116 & n1363;
  assign n2164 = pi85 & ~n1362;
  assign n2165 = pi26 & pi53;
  assign n2166 = ~pi58 & ~n2165;
  assign n2167 = ~pi85 & ~n2165;
  assign n2168 = ~n1362 & ~n2167;
  assign n2169 = ~pi58 & ~n2168;
  assign n2170 = ~n2164 & n2166;
  assign n2171 = ~n2163 & ~n3058;
  assign n2172 = pi57 & ~n2171;
  assign n2173 = pi58 & pi60;
  assign n2174 = pi60 & n1849;
  assign n2175 = pi116 & n2173;
  assign n2176 = n1363 & n3059;
  assign n2177 = ~n2172 & ~n2176;
  assign n2178 = ~pi27 & ~n2177;
  assign n2179 = pi57 & ~pi58;
  assign n2180 = n1363 & n2179;
  assign n2181 = ~n2178 & ~n2180;
  assign n2182 = ~pi129 & ~n2181;
  assign n2183 = ~pi3 & n2182;
  assign n2184 = n479 & ~n2181;
  assign n2185 = pi136 & ~pi138;
  assign n2186 = pi31 & n2185;
  assign n2187 = pi115 & pi138;
  assign n2188 = ~pi87 & ~pi138;
  assign n2189 = ~pi136 & ~n2188;
  assign n2190 = ~pi115 & pi138;
  assign n2191 = pi87 & ~pi138;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = ~pi136 & ~n2192;
  assign n2194 = ~n2187 & n2189;
  assign n2195 = ~n2186 & ~n3061;
  assign n2196 = pi137 & ~n2195;
  assign n2197 = pi62 & ~pi138;
  assign n2198 = ~pi89 & pi138;
  assign n2199 = pi136 & ~n2198;
  assign n2200 = pi89 & pi138;
  assign n2201 = ~pi62 & ~pi138;
  assign n2202 = ~n2200 & ~n2201;
  assign n2203 = pi136 & ~n2202;
  assign n2204 = ~n2197 & n2199;
  assign n2205 = pi72 & ~pi138;
  assign n2206 = ~pi119 & pi138;
  assign n2207 = ~pi136 & ~n2206;
  assign n2208 = pi119 & pi138;
  assign n2209 = ~pi72 & ~pi138;
  assign n2210 = ~n2208 & ~n2209;
  assign n2211 = ~pi136 & ~n2210;
  assign n2212 = ~n2205 & n2207;
  assign n2213 = ~n3062 & ~n3063;
  assign n2214 = ~pi137 & ~n2213;
  assign n2215 = ~n2196 & ~n2214;
  assign n2216 = ~pi142 & n3018;
  assign n2217 = ~pi94 & ~n3018;
  assign n2218 = ~pi129 & ~n2217;
  assign n2219 = pi94 & ~n3018;
  assign n2220 = pi142 & n3018;
  assign n2221 = ~n2219 & ~n2220;
  assign n2222 = ~pi129 & ~n2221;
  assign n2223 = ~n2216 & n2218;
  assign n2224 = pi37 & n2185;
  assign n2225 = ~pi96 & pi138;
  assign n2226 = ~pi82 & ~pi138;
  assign n2227 = ~pi136 & ~n2226;
  assign n2228 = pi96 & pi138;
  assign n2229 = pi82 & ~pi138;
  assign n2230 = ~n2228 & ~n2229;
  assign n2231 = ~pi136 & ~n2230;
  assign n2232 = ~n2225 & n2227;
  assign n2233 = ~n2224 & ~n3065;
  assign n2234 = pi137 & ~n2233;
  assign n2235 = pi65 & ~pi138;
  assign n2236 = ~pi93 & pi138;
  assign n2237 = pi136 & ~n2236;
  assign n2238 = ~pi65 & ~pi138;
  assign n2239 = pi93 & pi138;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = pi136 & ~n2240;
  assign n2242 = ~n2235 & n2237;
  assign n2243 = pi77 & ~pi138;
  assign n2244 = ~pi124 & pi138;
  assign n2245 = ~pi136 & ~n2244;
  assign n2246 = pi124 & pi138;
  assign n2247 = ~pi77 & ~pi138;
  assign n2248 = ~n2246 & ~n2247;
  assign n2249 = ~pi136 & ~n2248;
  assign n2250 = ~n2243 & n2245;
  assign n2251 = ~n3066 & ~n3067;
  assign n2252 = ~pi137 & ~n2251;
  assign n2253 = ~n2234 & ~n2252;
  assign n2254 = pi35 & n2185;
  assign n2255 = ~pi100 & pi138;
  assign n2256 = ~pi80 & ~pi138;
  assign n2257 = ~pi136 & ~n2256;
  assign n2258 = pi80 & ~pi138;
  assign n2259 = pi100 & pi138;
  assign n2260 = ~n2258 & ~n2259;
  assign n2261 = ~pi136 & ~n2260;
  assign n2262 = ~n2255 & n2257;
  assign n2263 = ~n2254 & ~n3068;
  assign n2264 = pi137 & ~n2263;
  assign n2265 = pi70 & ~pi138;
  assign n2266 = ~pi92 & pi138;
  assign n2267 = pi136 & ~n2266;
  assign n2268 = pi92 & pi138;
  assign n2269 = ~pi70 & ~pi138;
  assign n2270 = ~n2268 & ~n2269;
  assign n2271 = pi136 & ~n2270;
  assign n2272 = ~n2265 & n2267;
  assign n2273 = pi75 & ~pi138;
  assign n2274 = ~pi125 & pi138;
  assign n2275 = ~pi136 & ~n2274;
  assign n2276 = pi125 & pi138;
  assign n2277 = ~pi75 & ~pi138;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = ~pi136 & ~n2278;
  assign n2280 = ~n2273 & n2275;
  assign n2281 = ~n3069 & ~n3070;
  assign n2282 = ~pi137 & ~n2281;
  assign n2283 = ~n2264 & ~n2282;
  assign n2284 = pi36 & n2185;
  assign n2285 = ~pi97 & pi138;
  assign n2286 = ~pi81 & ~pi138;
  assign n2287 = ~pi136 & ~n2286;
  assign n2288 = pi81 & ~pi138;
  assign n2289 = pi97 & pi138;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = ~pi136 & ~n2290;
  assign n2292 = ~n2285 & n2287;
  assign n2293 = ~n2284 & ~n3071;
  assign n2294 = pi137 & ~n2293;
  assign n2295 = pi71 & ~pi138;
  assign n2296 = ~pi98 & pi138;
  assign n2297 = pi136 & ~n2296;
  assign n2298 = pi98 & pi138;
  assign n2299 = ~pi71 & ~pi138;
  assign n2300 = ~n2298 & ~n2299;
  assign n2301 = pi136 & ~n2300;
  assign n2302 = ~n2295 & n2297;
  assign n2303 = pi76 & ~pi138;
  assign n2304 = ~pi23 & pi138;
  assign n2305 = ~pi136 & ~n2304;
  assign n2306 = ~pi76 & ~pi138;
  assign n2307 = pi23 & pi138;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = ~pi136 & ~n2308;
  assign n2310 = ~n2303 & n2305;
  assign n2311 = ~n3072 & ~n3073;
  assign n2312 = ~pi137 & ~n2311;
  assign n2313 = ~n2294 & ~n2312;
  assign n2314 = pi30 & n2185;
  assign n2315 = ~pi111 & pi138;
  assign n2316 = ~pi86 & ~pi138;
  assign n2317 = ~pi136 & ~n2316;
  assign n2318 = pi86 & ~pi138;
  assign n2319 = pi111 & pi138;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = ~pi136 & ~n2320;
  assign n2322 = ~n2315 & n2317;
  assign n2323 = ~n2314 & ~n3074;
  assign n2324 = pi137 & ~n2323;
  assign n2325 = pi64 & ~pi138;
  assign n2326 = ~pi88 & pi138;
  assign n2327 = pi136 & ~n2326;
  assign n2328 = pi88 & pi138;
  assign n2329 = ~pi64 & ~pi138;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = pi136 & ~n2330;
  assign n2332 = ~n2325 & n2327;
  assign n2333 = pi67 & ~pi138;
  assign n2334 = ~pi120 & pi138;
  assign n2335 = ~pi136 & ~n2334;
  assign n2336 = pi120 & pi138;
  assign n2337 = ~pi67 & ~pi138;
  assign n2338 = ~n2336 & ~n2337;
  assign n2339 = ~pi136 & ~n2338;
  assign n2340 = ~n2333 & n2335;
  assign n2341 = ~n3075 & ~n3076;
  assign n2342 = ~pi137 & ~n2341;
  assign n2343 = ~n2324 & ~n2342;
  assign n2344 = ~pi139 & n3016;
  assign n2345 = ~pi129 & n3015;
  assign n2346 = ~pi111 & ~n3016;
  assign n2347 = n2345 & ~n2346;
  assign n2348 = pi111 & ~n3016;
  assign n2349 = pi82 & n1888;
  assign n2350 = pi138 & n1890;
  assign n2351 = ~pi136 & pi139;
  assign n2352 = n3077 & n2351;
  assign n2353 = ~n2348 & ~n2352;
  assign n2354 = n3015 & ~n2353;
  assign n2355 = ~pi129 & n2354;
  assign n2356 = n2345 & ~n2353;
  assign n2357 = ~n2344 & n2347;
  assign n2358 = pi112 & ~n3016;
  assign n2359 = ~pi141 & n3016;
  assign n2360 = n2345 & ~n2359;
  assign n2361 = ~pi136 & pi141;
  assign n2362 = n3077 & n2361;
  assign n2363 = ~pi112 & ~n3016;
  assign n2364 = ~n2362 & ~n2363;
  assign n2365 = n3015 & ~n2364;
  assign n2366 = ~pi129 & n2365;
  assign n2367 = n2345 & ~n2364;
  assign n2368 = ~n2358 & n2360;
  assign n2369 = pi115 & ~n3016;
  assign n2370 = ~pi140 & n3016;
  assign n2371 = n2345 & ~n2370;
  assign n2372 = ~pi136 & pi140;
  assign n2373 = n3077 & n2372;
  assign n2374 = ~pi115 & ~n3016;
  assign n2375 = ~n2373 & ~n2374;
  assign n2376 = n3015 & ~n2375;
  assign n2377 = ~pi129 & n2376;
  assign n2378 = n2345 & ~n2375;
  assign n2379 = ~n2369 & n2371;
  assign n2380 = ~pi137 & ~pi138;
  assign n2381 = pi136 & n2380;
  assign n2382 = ~pi138 & n1922;
  assign n2383 = ~pi138 & n3015;
  assign n2384 = n1922 & n2383;
  assign n2385 = n3015 & n3081;
  assign n2386 = pi140 & n3082;
  assign n2387 = ~pi62 & ~n3082;
  assign n2388 = ~pi129 & ~n2387;
  assign n2389 = pi62 & ~n3082;
  assign n2390 = ~pi140 & n1922;
  assign n2391 = n2383 & n2390;
  assign n2392 = ~n2389 & ~n2391;
  assign n2393 = ~pi129 & ~n2392;
  assign n2394 = ~n2386 & n2388;
  assign n2395 = pi142 & n3082;
  assign n2396 = ~pi63 & ~n3082;
  assign n2397 = ~pi129 & ~n2396;
  assign n2398 = pi63 & ~n3082;
  assign n2399 = ~pi142 & n1922;
  assign n2400 = n2383 & n2399;
  assign n2401 = ~n2398 & ~n2400;
  assign n2402 = ~pi129 & ~n2401;
  assign n2403 = ~n2395 & n2397;
  assign n2404 = pi139 & n3082;
  assign n2405 = ~pi64 & ~n3082;
  assign n2406 = ~pi129 & ~n2405;
  assign n2407 = pi64 & ~n3082;
  assign n2408 = ~pi139 & n1922;
  assign n2409 = n2383 & n2408;
  assign n2410 = ~n2407 & ~n2409;
  assign n2411 = ~pi129 & ~n2410;
  assign n2412 = ~n2404 & n2406;
  assign n2413 = pi146 & n3082;
  assign n2414 = ~pi65 & ~n3082;
  assign n2415 = ~pi129 & ~n2414;
  assign n2416 = pi65 & ~n3082;
  assign n2417 = ~pi146 & n1922;
  assign n2418 = n2383 & n2417;
  assign n2419 = ~n2416 & ~n2418;
  assign n2420 = ~pi129 & ~n2419;
  assign n2421 = ~n2413 & n2415;
  assign n2422 = n1885 & n2383;
  assign n2423 = pi143 & n2422;
  assign n2424 = ~pi66 & ~n2422;
  assign n2425 = ~pi129 & ~n2424;
  assign n2426 = pi66 & ~n2422;
  assign n2427 = ~pi143 & n2422;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = ~pi129 & ~n2428;
  assign n2430 = ~n2423 & n2425;
  assign n2431 = pi139 & n2422;
  assign n2432 = ~pi67 & ~n2422;
  assign n2433 = ~pi129 & ~n2432;
  assign n2434 = pi67 & ~n2422;
  assign n2435 = ~pi139 & n2422;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = ~pi129 & ~n2436;
  assign n2438 = ~n2431 & n2433;
  assign n2439 = pi141 & n3082;
  assign n2440 = ~pi68 & ~n3082;
  assign n2441 = ~pi129 & ~n2440;
  assign n2442 = pi68 & ~n3082;
  assign n2443 = ~pi141 & n1922;
  assign n2444 = n2383 & n2443;
  assign n2445 = ~n2442 & ~n2444;
  assign n2446 = ~pi129 & ~n2445;
  assign n2447 = ~n2439 & n2441;
  assign n2448 = pi143 & n3082;
  assign n2449 = ~pi69 & ~n3082;
  assign n2450 = ~pi129 & ~n2449;
  assign n2451 = pi69 & ~n3082;
  assign n2452 = ~pi143 & n1922;
  assign n2453 = n2383 & n2452;
  assign n2454 = ~n2451 & ~n2453;
  assign n2455 = ~pi129 & ~n2454;
  assign n2456 = ~n2448 & n2450;
  assign n2457 = pi144 & n3082;
  assign n2458 = ~pi70 & ~n3082;
  assign n2459 = ~pi129 & ~n2458;
  assign n2460 = pi70 & ~n3082;
  assign n2461 = ~pi144 & n1922;
  assign n2462 = n2383 & n2461;
  assign n2463 = ~n2460 & ~n2462;
  assign n2464 = ~pi129 & ~n2463;
  assign n2465 = ~n2457 & n2459;
  assign n2466 = pi145 & n3082;
  assign n2467 = ~pi71 & ~n3082;
  assign n2468 = ~pi129 & ~n2467;
  assign n2469 = pi71 & ~n3082;
  assign n2470 = ~pi145 & n1922;
  assign n2471 = n2383 & n2470;
  assign n2472 = ~n2469 & ~n2471;
  assign n2473 = ~pi129 & ~n2472;
  assign n2474 = ~n2466 & n2468;
  assign n2475 = pi140 & n2422;
  assign n2476 = ~pi72 & ~n2422;
  assign n2477 = ~pi129 & ~n2476;
  assign n2478 = pi72 & ~n2422;
  assign n2479 = ~pi140 & n2422;
  assign n2480 = ~n2478 & ~n2479;
  assign n2481 = ~pi129 & ~n2480;
  assign n2482 = ~n2475 & n2477;
  assign n2483 = pi141 & n2422;
  assign n2484 = ~pi73 & ~n2422;
  assign n2485 = ~pi129 & ~n2484;
  assign n2486 = pi73 & ~n2422;
  assign n2487 = ~pi141 & n2422;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = ~pi129 & ~n2488;
  assign n2490 = ~n2483 & n2485;
  assign n2491 = pi142 & n2422;
  assign n2492 = ~pi74 & ~n2422;
  assign n2493 = ~pi129 & ~n2492;
  assign n2494 = pi74 & ~n2422;
  assign n2495 = ~pi142 & n2422;
  assign n2496 = ~n2494 & ~n2495;
  assign n2497 = ~pi129 & ~n2496;
  assign n2498 = ~n2491 & n2493;
  assign n2499 = pi144 & n2422;
  assign n2500 = ~pi75 & ~n2422;
  assign n2501 = ~pi129 & ~n2500;
  assign n2502 = pi75 & ~n2422;
  assign n2503 = ~pi144 & n2422;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = ~pi129 & ~n2504;
  assign n2506 = ~n2499 & n2501;
  assign n2507 = pi145 & n2422;
  assign n2508 = ~pi76 & ~n2422;
  assign n2509 = ~pi129 & ~n2508;
  assign n2510 = pi76 & ~n2422;
  assign n2511 = ~pi145 & n2422;
  assign n2512 = ~n2510 & ~n2511;
  assign n2513 = ~pi129 & ~n2512;
  assign n2514 = ~n2507 & n2509;
  assign n2515 = pi146 & n2422;
  assign n2516 = ~pi77 & ~n2422;
  assign n2517 = ~pi129 & ~n2516;
  assign n2518 = pi77 & ~n2422;
  assign n2519 = ~pi146 & n2422;
  assign n2520 = ~n2518 & ~n2519;
  assign n2521 = ~pi129 & ~n2520;
  assign n2522 = ~n2515 & n2517;
  assign n2523 = n1924 & n2383;
  assign n2524 = ~pi142 & n2523;
  assign n2525 = ~pi78 & ~n2523;
  assign n2526 = ~pi129 & ~n2525;
  assign n2527 = pi78 & ~n2523;
  assign n2528 = pi142 & n2523;
  assign n2529 = ~n2527 & ~n2528;
  assign n2530 = ~pi129 & ~n2529;
  assign n2531 = ~n2524 & n2526;
  assign n2532 = ~pi143 & n2523;
  assign n2533 = ~pi79 & ~n2523;
  assign n2534 = ~pi129 & ~n2533;
  assign n2535 = pi79 & ~n2523;
  assign n2536 = pi143 & n2523;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = ~pi129 & ~n2537;
  assign n2539 = ~n2532 & n2534;
  assign n2540 = ~pi144 & n2523;
  assign n2541 = ~pi80 & ~n2523;
  assign n2542 = ~pi129 & ~n2541;
  assign n2543 = pi80 & ~n2523;
  assign n2544 = pi144 & n2523;
  assign n2545 = ~n2543 & ~n2544;
  assign n2546 = ~pi129 & ~n2545;
  assign n2547 = ~n2540 & n2542;
  assign n2548 = ~pi145 & n2523;
  assign n2549 = ~pi81 & ~n2523;
  assign n2550 = ~pi129 & ~n2549;
  assign n2551 = pi81 & ~n2523;
  assign n2552 = pi145 & n2523;
  assign n2553 = ~n2551 & ~n2552;
  assign n2554 = ~pi129 & ~n2553;
  assign n2555 = ~n2548 & n2550;
  assign n2556 = ~pi146 & n2523;
  assign n2557 = ~pi82 & ~n2523;
  assign n2558 = ~pi129 & ~n2557;
  assign n2559 = pi82 & ~n2523;
  assign n2560 = pi146 & n2523;
  assign n2561 = ~n2559 & ~n2560;
  assign n2562 = ~pi129 & ~n2561;
  assign n2563 = ~n2556 & n2558;
  assign n2564 = ~pi141 & n2523;
  assign n2565 = ~pi84 & ~n2523;
  assign n2566 = ~pi129 & ~n2565;
  assign n2567 = pi84 & ~n2523;
  assign n2568 = pi141 & n2523;
  assign n2569 = ~n2567 & ~n2568;
  assign n2570 = ~pi129 & ~n2569;
  assign n2571 = ~n2564 & n2566;
  assign n2572 = ~pi139 & n2523;
  assign n2573 = ~pi86 & ~n2523;
  assign n2574 = ~pi129 & ~n2573;
  assign n2575 = pi86 & ~n2523;
  assign n2576 = pi139 & n2523;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = ~pi129 & ~n2577;
  assign n2579 = ~n2572 & n2574;
  assign n2580 = ~pi140 & n2523;
  assign n2581 = ~pi87 & ~n2523;
  assign n2582 = ~pi129 & ~n2581;
  assign n2583 = pi87 & ~n2523;
  assign n2584 = pi140 & n2523;
  assign n2585 = ~n2583 & ~n2584;
  assign n2586 = ~pi129 & ~n2585;
  assign n2587 = ~n2580 & n2582;
  assign n2588 = pi137 & n2185;
  assign n2589 = pi136 & pi137;
  assign n2590 = n2383 & n2589;
  assign n2591 = n3015 & n2588;
  assign n2592 = ~pi139 & n3107;
  assign n2593 = ~pi88 & ~n3107;
  assign n2594 = ~pi129 & ~n2593;
  assign n2595 = pi88 & ~n3107;
  assign n2596 = pi139 & n3107;
  assign n2597 = ~n2595 & ~n2596;
  assign n2598 = ~pi129 & ~n2597;
  assign n2599 = ~n2592 & n2594;
  assign n2600 = ~pi140 & n3107;
  assign n2601 = ~pi89 & ~n3107;
  assign n2602 = ~pi129 & ~n2601;
  assign n2603 = pi89 & ~n3107;
  assign n2604 = pi140 & n3107;
  assign n2605 = ~n2603 & ~n2604;
  assign n2606 = ~pi129 & ~n2605;
  assign n2607 = ~n2600 & n2602;
  assign n2608 = ~pi142 & n3107;
  assign n2609 = ~pi90 & ~n3107;
  assign n2610 = ~pi129 & ~n2609;
  assign n2611 = pi90 & ~n3107;
  assign n2612 = pi142 & n3107;
  assign n2613 = ~n2611 & ~n2612;
  assign n2614 = ~pi129 & ~n2613;
  assign n2615 = ~n2608 & n2610;
  assign n2616 = ~pi143 & n3107;
  assign n2617 = ~pi91 & ~n3107;
  assign n2618 = ~pi129 & ~n2617;
  assign n2619 = pi91 & ~n3107;
  assign n2620 = pi143 & n3107;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = ~pi129 & ~n2621;
  assign n2623 = ~n2616 & n2618;
  assign n2624 = ~pi144 & n3107;
  assign n2625 = ~pi92 & ~n3107;
  assign n2626 = ~pi129 & ~n2625;
  assign n2627 = pi92 & ~n3107;
  assign n2628 = pi144 & n3107;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = ~pi129 & ~n2629;
  assign n2631 = ~n2624 & n2626;
  assign n2632 = ~pi146 & n3107;
  assign n2633 = ~pi93 & ~n3107;
  assign n2634 = ~pi129 & ~n2633;
  assign n2635 = pi93 & ~n3107;
  assign n2636 = pi146 & n3107;
  assign n2637 = ~n2635 & ~n2636;
  assign n2638 = ~pi129 & ~n2637;
  assign n2639 = ~n2632 & n2634;
  assign n2640 = ~pi145 & n3107;
  assign n2641 = ~pi98 & ~n3107;
  assign n2642 = ~pi129 & ~n2641;
  assign n2643 = pi98 & ~n3107;
  assign n2644 = pi145 & n3107;
  assign n2645 = ~n2643 & ~n2644;
  assign n2646 = ~pi129 & ~n2645;
  assign n2647 = ~n2640 & n2642;
  assign n2648 = ~pi141 & n3107;
  assign n2649 = ~pi99 & ~n3107;
  assign n2650 = ~pi129 & ~n2649;
  assign n2651 = pi99 & ~n3107;
  assign n2652 = pi141 & n3107;
  assign n2653 = ~n2651 & ~n2652;
  assign n2654 = ~pi129 & ~n2653;
  assign n2655 = ~n2648 & n2650;
  assign n2656 = pi91 & n1922;
  assign n2657 = pi95 & n1924;
  assign n2658 = ~n2656 & ~n2657;
  assign n2659 = pi138 & ~n2658;
  assign n2660 = ~pi34 & pi136;
  assign n2661 = ~pi79 & ~pi136;
  assign n2662 = pi137 & ~n2661;
  assign n2663 = pi79 & ~pi136;
  assign n2664 = pi34 & pi136;
  assign n2665 = ~n2663 & ~n2664;
  assign n2666 = pi137 & ~n2665;
  assign n2667 = ~n2660 & n2662;
  assign n2668 = pi69 & pi136;
  assign n2669 = pi66 & ~pi136;
  assign n2670 = ~pi137 & ~n2669;
  assign n2671 = ~pi69 & pi136;
  assign n2672 = ~pi66 & ~pi136;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = ~pi137 & ~n2673;
  assign n2675 = ~n2668 & n2670;
  assign n2676 = ~n3116 & ~n3117;
  assign n2677 = ~pi138 & ~n2676;
  assign n2678 = ~n2659 & ~n2677;
  assign n2679 = pi90 & n1922;
  assign n2680 = pi94 & n1924;
  assign n2681 = ~n2679 & ~n2680;
  assign n2682 = pi138 & ~n2681;
  assign n2683 = ~pi33 & pi136;
  assign n2684 = ~pi78 & ~pi136;
  assign n2685 = pi137 & ~n2684;
  assign n2686 = pi78 & ~pi136;
  assign n2687 = pi33 & pi136;
  assign n2688 = ~n2686 & ~n2687;
  assign n2689 = pi137 & ~n2688;
  assign n2690 = ~n2683 & n2685;
  assign n2691 = pi63 & pi136;
  assign n2692 = pi74 & ~pi136;
  assign n2693 = ~pi137 & ~n2692;
  assign n2694 = ~pi63 & pi136;
  assign n2695 = ~pi74 & ~pi136;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = ~pi137 & ~n2696;
  assign n2698 = ~n2691 & n2693;
  assign n2699 = ~n3118 & ~n3119;
  assign n2700 = ~pi138 & ~n2699;
  assign n2701 = ~n2682 & ~n2700;
  assign n2702 = ~pi26 & n2920;
  assign n2703 = pi116 & n479;
  assign n2704 = ~n2925 & n2703;
  assign n2705 = ~n2920 & n1311;
  assign n2706 = ~n1310 & ~n2705;
  assign n2707 = ~pi129 & ~n2706;
  assign n2708 = ~pi3 & n2707;
  assign n2709 = pi116 & n2708;
  assign n2710 = n2703 & ~n2706;
  assign n2711 = ~n2702 & n2704;
  assign n2712 = ~pi4 & ~pi9;
  assign n2713 = ~pi4 & ~pi12;
  assign n2714 = ~pi7 & ~pi9;
  assign n2715 = n2713 & n2714;
  assign n2716 = ~pi4 & ~pi7;
  assign n2717 = ~pi9 & ~pi12;
  assign n2718 = n2716 & n2717;
  assign n2719 = n482 & n2712;
  assign n2720 = pi54 & n479;
  assign n2721 = ~pi129 & ~n3121;
  assign n2722 = ~pi3 & n2721;
  assign n2723 = pi54 & n2722;
  assign n2724 = ~n3121 & n2720;
  assign n2725 = pi122 & ~pi129;
  assign n2726 = ~pi54 & pi118;
  assign n2727 = pi54 & ~pi59;
  assign n2728 = n2815 & n2727;
  assign n2729 = ~n2726 & ~n2728;
  assign po133 = ~pi129 & ~n2729;
  assign n2731 = ~pi97 & n1225;
  assign n2732 = ~n1226 & ~n2731;
  assign n2733 = ~pi129 & ~n2732;
  assign n2734 = ~pi3 & n2733;
  assign n2735 = pi116 & n2734;
  assign n2736 = n2703 & ~n2732;
  assign n2737 = ~pi11 & ~pi22;
  assign n2738 = pi54 & n2737;
  assign n2739 = ~pi54 & pi113;
  assign n2740 = n479 & ~n2739;
  assign n2741 = ~pi54 & ~pi113;
  assign n2742 = pi54 & ~n2737;
  assign n2743 = ~n2741 & ~n2742;
  assign n2744 = ~pi129 & ~n2743;
  assign n2745 = ~pi3 & n2744;
  assign n2746 = n479 & ~n2743;
  assign n2747 = ~n2738 & n2740;
  assign n2748 = ~pi110 & ~pi120;
  assign n2749 = ~pi3 & n2748;
  assign n2750 = ~pi120 & n1898;
  assign n2751 = ~pi111 & ~pi129;
  assign n2752 = ~pi129 & ~n3125;
  assign n2753 = ~pi111 & n2752;
  assign n2754 = ~n3125 & n2751;
  assign n2755 = ~pi129 & ~pi134;
  assign n2756 = ~pi129 & ~pi135;
  assign n2757 = ~pi96 & pi125;
  assign n2758 = ~pi3 & ~n2757;
  assign po140 = ~pi129 & ~n2758;
  assign po134 = ~pi129 & ~n1260;
  assign n2761 = pi81 & pi120;
  assign po136 = ~pi129 & n2761;
  assign n2763 = ~pi126 & pi132;
  assign po141 = pi133 & n2763;
  assign po139 = pi57 & ~pi129;
  assign n2766 = n303 | n299 | n302;
  assign n2767 = n300 | n301;
  assign n2768 = n304 | n306 | n308 | n309;
  assign n2769 = n317 | n318;
  assign n2770 = n320 | n321;
  assign n2771 = n322 | n323;
  assign n2772 = n324 | n325;
  assign n2773 = n326 | n327;
  assign n2774 = n329 | n330;
  assign n2775 = n331 | n332;
  assign n2776 = n333 | n335 | n336 | n337;
  assign n2777 = n340 | n341;
  assign n2778 = n342 | n343;
  assign n2779 = n344 | n345 | n346 | n347;
  assign n2780 = n352 | n348 | n351 | n355 | n356;
  assign n2781 = n359 | n357 | n358 | n361 | n362;
  assign n2782 = n367 | n368;
  assign n2783 = n370 | n371;
  assign n2784 = n376 | n377;
  assign n2785 = n378 | n379;
  assign n2786 = n382 | n380 | n381;
  assign n2787 = n389 | n390 | n408 | n409;
  assign n2788 = n399 | n397 | n398;
  assign n2789 = n402 | n400 | n401;
  assign n2790 = n407 | n403 | n406;
  assign n2791 = n411 | ~n412;
  assign n2792 = n414 | n415;
  assign n2793 = n421 | n427 | n447 | n449 | n455 | n453 | n454;
  assign n2794 = n422 | n423;
  assign n2795 = n428 | n429;
  assign n2796 = n430 | n431;
  assign n2797 = n442 | n432 | n441 | n446 | n444 | n445;
  assign n2798 = n436 | n437 | n439 | n440;
  assign n2799 = n467 | n463 | n464 | n470 | n471;
  assign n2800 = n473 | n474;
  assign n2801 = n475 | n476;
  assign n2802 = n485 | n486;
  assign n2803 = n491 | n492;
  assign n2804 = n495 | n496;
  assign n2805 = n502 | n503;
  assign n2806 = n504 | n505;
  assign n2807 = n512 | n509 | n511;
  assign n2808 = n520 | n516 | n519;
  assign n2809 = n536 | n526 | n535;
  assign n2810 = n528 | n529;
  assign po20 = n539 | n540;
  assign n2812 = n547 | n544 | n546;
  assign n2813 = n559 | n551 | n558;
  assign po21 = n562 | n563;
  assign n2815 = n567 | n568;
  assign n2816 = n602 | n571 | n579 | n608 | n609;
  assign n2817 = n585 | n582 | n584;
  assign n2818 = n590 | n586 | n589;
  assign n2819 = n587 | n588;
  assign n2820 = n600 | n595 | n599;
  assign n2821 = n598 | n596 | n597;
  assign po28 = n612 | n613;
  assign n2823 = n617 | n619 | n621 | n622;
  assign n2824 = n630 | n631;
  assign n2825 = n634 | n635;
  assign n2826 = n645 | n646;
  assign n2827 = n659 | n660;
  assign n2828 = n671 | n661 | n670;
  assign po32 = n674 | n675;
  assign n2830 = n678 | n679;
  assign n2831 = n683 | n684;
  assign n2832 = n695 | n689 | n694;
  assign n2833 = n692 | n693;
  assign n2834 = n700 | n701;
  assign n2835 = n706 | n707;
  assign n2836 = n710 | n711;
  assign n2837 = n714 | n715;
  assign n2838 = n735 | n723 | n731 | n740 | n741;
  assign n2839 = n726 | n727;
  assign n2840 = n756 | n757;
  assign n2841 = n765 | n766;
  assign n2842 = n779 | n772 | n778;
  assign n2843 = n783 | n784;
  assign n2844 = n791 | n789 | n790;
  assign n2845 = n799 | n800;
  assign n2846 = n804 | n805;
  assign n2847 = n808 | n809;
  assign n2848 = n813 | n814;
  assign n2849 = n819 | n821 | n823 | n824;
  assign n2850 = n837 | n838;
  assign n2851 = n841 | n842;
  assign n2852 = n843 | n844;
  assign n2853 = n855 | n853 | ~n854;
  assign n2854 = n856 | n857;
  assign n2855 = n861 | n862;
  assign n2856 = n865 | n866;
  assign n2857 = n868 | n869;
  assign n2858 = n878 | n876 | n877;
  assign n2859 = n881 | n882;
  assign n2860 = n886 | n887 | n888 | n889;
  assign po19 = n896 | n897;
  assign n2862 = n900 | n901;
  assign n2863 = n905 | n906;
  assign n2864 = n913 | n918 | n924 | n925;
  assign n2865 = n915 | n916;
  assign n2866 = n922 | n923;
  assign po22 = n928 | n929;
  assign n2868 = n937 | n941 | n943 | n944;
  assign n2869 = n939 | n940;
  assign po23 = n948 | n949;
  assign n2871 = n961 | n966 | n972 | n973;
  assign n2872 = n963 | n964;
  assign po24 = n976 | n977;
  assign n2874 = n983 | n984;
  assign n2875 = n986 | n987;
  assign n2876 = n988 | n989;
  assign n2877 = n996 | n998 | n1000 | n1001;
  assign po25 = n1004 | n1005;
  assign n2879 = n1011 | n1012;
  assign n2880 = n1017 | n1018;
  assign n2881 = n1026 | n1022 | n1025;
  assign po26 = n1029 | n1030;
  assign n2883 = n1039 | n1042 | n1048 | n1049;
  assign n2884 = n1046 | n1047;
  assign po27 = n1052 | n1053;
  assign n2886 = n1074 | n1064 | n1073;
  assign n2887 = n1068 | n1069;
  assign n2888 = n1071 | n1072;
  assign po29 = n1077 | n1078;
  assign n2890 = n1082 | n1083;
  assign n2891 = n1086 | n1087;
  assign n2892 = n1089 | n1090;
  assign po31 = n1093 | n1094;
  assign n2894 = n1097 | n1098;
  assign n2895 = n1104 | n1100 | n1103;
  assign n2896 = n1105 | n1106;
  assign n2897 = n1107 | n1108;
  assign po33 = n1111 | n1112;
  assign n2899 = n1122 | n1118 | n1121;
  assign n2900 = n1125 | n1126;
  assign po34 = n1129 | n1130;
  assign n2902 = n1138 | n1139;
  assign n2903 = n1142 | n1143;
  assign n2904 = n1150 | n1151;
  assign n2905 = n1152 | n1153;
  assign n2906 = n1156 | n1157;
  assign n2907 = n1158 | n1159;
  assign po36 = n1163 | n1164;
  assign n2909 = n1170 | n1167 | n1169;
  assign n2910 = n1178 | n1180 | n1183 | n1184;
  assign po37 = n1187 | n1188;
  assign n2912 = n1190 | n1191;
  assign n2913 = n1195 | n1196;
  assign n2914 = n1218 | n1214 | n1217;
  assign n2915 = n1220 | n1221;
  assign po39 = n1223 | n1224;
  assign n2917 = n1235 | n1236;
  assign n2918 = n1238 | n1239;
  assign n2919 = n1241 | n1242;
  assign n2920 = n1247 | n1248;
  assign n2921 = n1278 | n1279;
  assign n2922 = n1286 | n1287;
  assign n2923 = n1289 | n1290;
  assign po40 = n1304 | n1302 | n1303;
  assign n2925 = n1312 | ~n1313;
  assign n2926 = n1322 | n1323;
  assign n2927 = n1324 | n1325;
  assign n2928 = n1347 | n1348;
  assign n2929 = n1350 | n1351;
  assign n2930 = n1356 | n1357;
  assign n2931 = n1358 | n1359;
  assign n2932 = n1365 | n1366;
  assign n2933 = n1368 | n1369;
  assign po43 = n1372 | n1373;
  assign n2935 = n1379 | n1380;
  assign n2936 = n1385 | n1386;
  assign n2937 = n1389 | n1390;
  assign n2938 = n1394 | n1395;
  assign po42 = n1398 | n1399;
  assign n2940 = n1402 | n1403;
  assign n2941 = n1406 | n1407;
  assign po41 = n1414 | n1415;
  assign n2943 = n1423 | n1421 | n1422;
  assign n2944 = n1426 | n1427;
  assign n2945 = n1432 | n1433;
  assign n2946 = n1435 | n1436;
  assign n2947 = n1441 | n1442;
  assign n2948 = n1449 | n1450;
  assign n2949 = n1456 | n1457;
  assign n2950 = n1462 | n1463;
  assign n2951 = n1466 | n1467;
  assign n2952 = n1469 | n1471 | n1473 | n1474;
  assign po44 = n1478 | n1479;
  assign n2954 = n1483 | n1481 | n1482;
  assign n2955 = n1484 | n1487 | n1488 | n1489;
  assign n2956 = n1490 | n1491;
  assign n2957 = n1497 | n1501 | n1504 | n1505;
  assign n2958 = n1500 | n1498 | n1499;
  assign n2959 = n1509 | n1510;
  assign n2960 = n1513 | n1514;
  assign n2961 = n1518 | n1515 | n1517;
  assign n2962 = n1523 | n1524;
  assign n2963 = n1534 | n1531 | n1533;
  assign n2964 = n1538 | n1539;
  assign n2965 = n1541 | n1542;
  assign n2966 = n1552 | n1553;
  assign n2967 = n1554 | n1555;
  assign n2968 = n1559 | n1560;
  assign n2969 = n1562 | n1563;
  assign n2970 = n1566 | n1567;
  assign po56 = n1571 | n1572;
  assign n2972 = n1576 | n1574 | n1575;
  assign n2973 = n1591 | n1589 | n1590;
  assign n2974 = n1595 | n1596;
  assign po57 = n1600 | n1601;
  assign n2976 = n1608 | n1609;
  assign n2977 = n1613 | n1614;
  assign n2978 = n1623 | n1618 | n1622;
  assign n2979 = n1620 | n1621;
  assign po58 = n1627 | n1628;
  assign n2981 = n1629 | n1630;
  assign n2982 = n1636 | ~n1637;
  assign n2983 = n1644 | n1642 | n1643;
  assign n2984 = n1648 | n1649;
  assign n2985 = n1657 | n1658;
  assign n2986 = n1660 | n1661;
  assign po60 = n1665 | n1666;
  assign n2988 = n1684 | n1685;
  assign n2989 = n1688 | n1689;
  assign po61 = n1692 | n1693;
  assign n2991 = n1703 | n1704;
  assign n2992 = n1713 | n1709 | n1711 | n1715 | n1716;
  assign po62 = n1720 | n1721;
  assign n2994 = n1724 | n1725;
  assign n2995 = n1729 | n1730;
  assign n2996 = n1740 | n1742 | n1746 | n1747;
  assign po63 = n1751 | n1752;
  assign n2998 = n1760 | n1758 | n1759;
  assign n2999 = n1762 | n1763;
  assign n3000 = n1768 | n1769;
  assign n3001 = n1772 | n1773;
  assign n3002 = n1785 | n1786;
  assign n3003 = n1790 | n1791;
  assign n3004 = n1801 | n1798 | n1800;
  assign po65 = n1807 | n1804 | n1806;
  assign n3006 = n1821 | n1822;
  assign n3007 = n1823 | n1824;
  assign n3008 = n1835 | n1832 | n1834;
  assign po74 = n1841 | n1842;
  assign n3010 = n1854 | n1852 | n1853;
  assign n3011 = n1858 | n1859;
  assign po68 = n1868 | n1865 | n1867;
  assign n3013 = n1872 | n1869 | n1871;
  assign po100 = n1879 | n1880;
  assign n3015 = n1883 | n1884;
  assign n3016 = n1894 | n1889 | n1893;
  assign n3017 = n1891 | n1892;
  assign n3018 = n1896 | n1897;
  assign n3019 = n1901 | n1902;
  assign n3020 = n1904 | ~n1905;
  assign n3021 = n1934 | n1935;
  assign n3022 = n1942 | n1943;
  assign n3023 = n1951 | ~n1952;
  assign n3024 = n1954 | n1955;
  assign po45 = n1961 | n1962;
  assign n3026 = n1967 | ~n1968;
  assign n3027 = n1970 | n1971;
  assign po46 = n1977 | n1978;
  assign n3029 = n1983 | ~n1984;
  assign n3030 = n1986 | n1987;
  assign po47 = n1993 | n1994;
  assign n3032 = n1999 | ~n2000;
  assign n3033 = n2002 | n2003;
  assign po48 = n2009 | n2010;
  assign n3035 = n2015 | ~n2016;
  assign n3036 = n2018 | n2019;
  assign po49 = n2025 | n2026;
  assign n3038 = n2031 | ~n2032;
  assign n3039 = n2034 | n2035;
  assign po50 = n2041 | n2042;
  assign n3041 = n2047 | ~n2048;
  assign n3042 = n2050 | n2051;
  assign po51 = n2057 | n2058;
  assign n3044 = n2063 | ~n2064;
  assign n3045 = n2066 | n2067;
  assign po52 = n2073 | n2074;
  assign po38 = n2089 | n2090;
  assign n3048 = n2094 | n2095;
  assign po76 = n2108 | n2109;
  assign n3050 = n2110 | n2111;
  assign n3051 = n2113 | n2114;
  assign po121 = n2117 | n2118;
  assign n3053 = n2127 | n2123 | n2126;
  assign po73 = n2134 | n2135;
  assign n3055 = n2140 | n2141;
  assign n3056 = n2153 | n2154;
  assign po71 = n2162 | n2160 | n2161;
  assign n3058 = n2169 | n2170;
  assign n3059 = n2174 | n2175;
  assign po72 = n2183 | n2184;
  assign n3061 = n2193 | n2194;
  assign n3062 = n2203 | n2204;
  assign n3063 = n2211 | n2212;
  assign po109 = n2222 | n2223;
  assign n3065 = n2231 | n2232;
  assign n3066 = n2241 | n2242;
  assign n3067 = n2249 | n2250;
  assign n3068 = n2261 | n2262;
  assign n3069 = n2271 | n2272;
  assign n3070 = n2279 | n2280;
  assign n3071 = n2291 | n2292;
  assign n3072 = n2301 | n2302;
  assign n3073 = n2309 | n2310;
  assign n3074 = n2321 | n2322;
  assign n3075 = n2331 | n2332;
  assign n3076 = n2339 | n2340;
  assign n3077 = n2349 | n2350;
  assign po126 = n2357 | n2355 | n2356;
  assign po127 = n2368 | n2366 | n2367;
  assign po130 = n2379 | n2377 | n2378;
  assign n3081 = n2381 | n2382;
  assign n3082 = n2384 | n2385;
  assign n3083 = n2393 | n2394;
  assign n3084 = n2402 | n2403;
  assign n3085 = n2411 | n2412;
  assign n3086 = n2420 | n2421;
  assign n3087 = n2429 | n2430;
  assign n3088 = n2437 | n2438;
  assign n3089 = n2446 | n2447;
  assign n3090 = n2455 | n2456;
  assign n3091 = n2464 | n2465;
  assign n3092 = n2473 | n2474;
  assign n3093 = n2481 | n2482;
  assign n3094 = n2489 | n2490;
  assign n3095 = n2497 | n2498;
  assign n3096 = n2505 | n2506;
  assign n3097 = n2513 | n2514;
  assign n3098 = n2521 | n2522;
  assign po93 = n2530 | n2531;
  assign po94 = n2538 | n2539;
  assign po95 = n2546 | n2547;
  assign po96 = n2554 | n2555;
  assign po97 = n2562 | n2563;
  assign po99 = n2570 | n2571;
  assign po101 = n2578 | n2579;
  assign po102 = n2586 | n2587;
  assign n3107 = n2590 | n2591;
  assign po103 = n2598 | n2599;
  assign po104 = n2606 | n2607;
  assign po105 = n2614 | n2615;
  assign po106 = n2622 | n2623;
  assign po107 = n2630 | n2631;
  assign po108 = n2638 | n2639;
  assign po113 = n2646 | n2647;
  assign po114 = n2654 | n2655;
  assign n3116 = n2666 | n2667;
  assign n3117 = n2674 | n2675;
  assign n3118 = n2689 | n2690;
  assign n3119 = n2697 | n2698;
  assign po124 = n2711 | n2709 | n2710;
  assign n3121 = n2719 | n2715 | n2718;
  assign po131 = n2723 | n2724;
  assign po125 = n2735 | n2736;
  assign po128 = n2747 | n2745 | n2746;
  assign n3125 = n2749 | n2750;
  assign po135 = n2753 | n2754;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
  assign po15 = ~n2847;
  assign po16 = ~n2859;
  assign po69 = ~n1808;
  assign po75 = ~n2103;
  assign po77 = ~n3083;
  assign po78 = ~n3084;
  assign po79 = ~n3085;
  assign po80 = ~n3086;
  assign po81 = ~n3087;
  assign po82 = ~n3088;
  assign po83 = ~n3089;
  assign po84 = ~n3090;
  assign po85 = ~n3091;
  assign po86 = ~n3092;
  assign po87 = ~n3093;
  assign po88 = ~n3094;
  assign po89 = ~n3095;
  assign po90 = ~n3096;
  assign po91 = ~n3097;
  assign po92 = ~n3098;
  assign po98 = ~n2215;
  assign po116 = ~n2253;
  assign po117 = ~n2678;
  assign po118 = ~n2701;
  assign po119 = ~n1946;
  assign po120 = ~n2283;
  assign po122 = ~n2313;
  assign po123 = ~n2343;
  assign po129 = ~n2097;
  assign po132 = ~n2725;
  assign po137 = ~n2755;
  assign po138 = ~n2756;
endmodule
