module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n417, n418,
    n419, n420, n421, n422, n424, n425, n426,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497,
    n498, n499, n500, n501, n502, n503, n504,
    n505, n506, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n566, n567, n568,
    n569, n570, n571, n572, n573, n574, n575,
    n576, n577, n578, n579, n580, n581, n582,
    n583, n584, n585, n586, n587, n589, n590,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639,
    n640, n642, n643, n644, n645, n646, n647,
    n648, n649, n650, n651, n652, n653, n654,
    n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n677, n678, n679, n680, n681, n682;
  assign n22 = ~pi5  & pi7 ;
  assign n23 = pi8  & n22;
  assign n24 = ~pi7  & pi9 ;
  assign n25 = ~n23 & ~n24;
  assign n26 = pi1  & ~n25;
  assign n27 = pi1  & ~pi7 ;
  assign n28 = ~pi5  & ~pi9 ;
  assign n29 = ~n27 & n28;
  assign n30 = ~n26 & ~n29;
  assign n31 = pi0  & ~pi2 ;
  assign n32 = ~n30 & n31;
  assign n33 = ~pi0  & ~pi1 ;
  assign n34 = pi2  & ~pi9 ;
  assign n35 = n33 & n34;
  assign n36 = n23 & n35;
  assign n37 = ~n32 & ~n36;
  assign n38 = ~pi3  & ~n37;
  assign n39 = ~pi3  & ~pi5 ;
  assign n40 = ~pi0  & pi9 ;
  assign n41 = pi1  & ~n40;
  assign n42 = ~pi1  & pi9 ;
  assign n43 = n39 & ~n42;
  assign n44 = ~n41 & n43;
  assign n45 = pi0  & ~pi9 ;
  assign n46 = ~pi1  & ~n45;
  assign n47 = pi1  & ~pi9 ;
  assign n48 = ~pi7  & ~n47;
  assign n49 = ~n46 & n48;
  assign n50 = ~n44 & ~n49;
  assign n51 = ~pi2  & ~n50;
  assign n52 = ~pi2  & ~pi3 ;
  assign n53 = pi9  & ~n52;
  assign n54 = pi0  & pi3 ;
  assign n55 = ~n53 & ~n54;
  assign n56 = ~pi1  & ~n55;
  assign n57 = pi1  & ~pi3 ;
  assign n58 = pi1  & pi2 ;
  assign n59 = ~pi2  & ~pi5 ;
  assign n60 = ~pi0  & ~n59;
  assign n61 = ~n58 & ~n60;
  assign n62 = ~pi9  & ~n61;
  assign n63 = ~n56 & ~n57;
  assign n64 = ~n62 & n63;
  assign n65 = ~pi7  & ~n64;
  assign n66 = ~n51 & ~n65;
  assign n67 = ~pi8  & ~n66;
  assign n68 = ~n38 & ~n67;
  assign n69 = ~pi6  & ~n68;
  assign n70 = ~pi1  & ~pi9 ;
  assign n71 = ~pi8  & n70;
  assign n72 = ~pi0  & n52;
  assign n73 = n71 & n72;
  assign n74 = ~pi0  & ~pi2 ;
  assign n75 = n42 & n74;
  assign n76 = ~pi5  & ~n75;
  assign n77 = pi6  & ~n76;
  assign n78 = ~n40 & ~n45;
  assign n79 = pi1  & pi5 ;
  assign n80 = pi2  & n79;
  assign n81 = n78 & n80;
  assign n82 = ~n77 & ~n81;
  assign n83 = pi8  & ~n82;
  assign n84 = ~pi1  & ~n40;
  assign n85 = ~pi8  & ~n84;
  assign n86 = ~pi1  & pi2 ;
  assign n87 = n45 & n86;
  assign n88 = ~n85 & ~n87;
  assign n89 = ~pi5  & ~n88;
  assign n90 = ~n83 & ~n89;
  assign n91 = pi3  & ~n90;
  assign n92 = pi1  & ~pi8 ;
  assign n93 = pi2  & ~pi3 ;
  assign n94 = n42 & n93;
  assign n95 = ~n92 & ~n94;
  assign n96 = ~pi0  & ~n95;
  assign n97 = pi2  & pi9 ;
  assign n98 = ~pi2  & pi6 ;
  assign n99 = pi3  & ~n98;
  assign n100 = n70 & ~n99;
  assign n101 = ~n97 & ~n100;
  assign n102 = ~pi8  & ~n101;
  assign n103 = ~n96 & ~n102;
  assign n104 = ~pi5  & ~n103;
  assign n105 = ~pi2  & ~n45;
  assign n106 = ~pi6  & ~n105;
  assign n107 = ~pi3  & n41;
  assign n108 = n105 & ~n107;
  assign n109 = pi5  & ~n106;
  assign n110 = ~n108 & n109;
  assign n111 = ~pi2  & n47;
  assign n112 = ~n97 & ~n111;
  assign n113 = ~pi0  & ~pi3 ;
  assign n114 = pi6  & n113;
  assign n115 = ~n112 & n114;
  assign n116 = ~n110 & ~n115;
  assign n117 = pi8  & ~n116;
  assign n118 = ~n73 & ~n104;
  assign n119 = ~n117 & n118;
  assign n120 = ~n91 & n119;
  assign n121 = ~pi7  & ~n120;
  assign n122 = ~n69 & ~n121;
  assign n123 = ~pi4  & ~n122;
  assign n124 = ~pi1  & ~pi3 ;
  assign n125 = ~pi6  & pi8 ;
  assign n126 = pi5  & ~n125;
  assign n127 = pi4  & pi8 ;
  assign n128 = ~pi6  & ~pi9 ;
  assign n129 = ~n127 & ~n128;
  assign n130 = n126 & ~n129;
  assign n131 = pi6  & ~pi9 ;
  assign n132 = pi4  & pi9 ;
  assign n133 = ~n131 & ~n132;
  assign n134 = pi5  & pi6 ;
  assign n135 = ~pi8  & ~n134;
  assign n136 = ~n133 & n135;
  assign n137 = ~n130 & ~n136;
  assign n138 = ~pi7  & n74;
  assign n139 = n124 & n138;
  assign n140 = ~n137 & n139;
  assign po0  = n123 | n140;
  assign n142 = n34 & n125;
  assign n143 = ~pi2  & ~pi8 ;
  assign n144 = ~pi0  & ~pi9 ;
  assign n145 = n143 & n144;
  assign n146 = pi0  & pi8 ;
  assign n147 = pi9  & n146;
  assign n148 = pi2  & n147;
  assign n149 = ~n145 & ~n148;
  assign n150 = pi5  & ~n149;
  assign n151 = ~pi8  & n28;
  assign n152 = ~pi5  & pi8 ;
  assign n153 = pi6  & pi9 ;
  assign n154 = ~n152 & ~n153;
  assign n155 = ~pi0  & ~n154;
  assign n156 = pi6  & pi8 ;
  assign n157 = pi9  & n156;
  assign n158 = ~n151 & ~n157;
  assign n159 = ~n155 & n158;
  assign n160 = pi2  & ~n159;
  assign n161 = ~n150 & ~n160;
  assign n162 = ~pi1  & ~n161;
  assign n163 = ~pi0  & pi5 ;
  assign n164 = ~pi8  & pi9 ;
  assign n165 = n163 & n164;
  assign n166 = pi0  & ~n156;
  assign n167 = ~n154 & n166;
  assign n168 = ~n165 & ~n167;
  assign n169 = ~pi2  & ~n168;
  assign n170 = ~pi6  & ~pi8 ;
  assign n171 = ~pi0  & pi6 ;
  assign n172 = ~pi2  & ~n171;
  assign n173 = n152 & ~n172;
  assign n174 = ~n170 & ~n173;
  assign n175 = ~pi9  & ~n174;
  assign n176 = ~n169 & ~n175;
  assign n177 = pi1  & ~n176;
  assign n178 = ~n142 & ~n162;
  assign n179 = ~n177 & n178;
  assign n180 = ~pi4  & ~n179;
  assign n181 = ~pi2  & n33;
  assign n182 = pi5  & ~pi8 ;
  assign n183 = ~n127 & ~n182;
  assign n184 = n128 & ~n183;
  assign n185 = pi4  & n153;
  assign n186 = ~n184 & ~n185;
  assign n187 = n181 & ~n186;
  assign n188 = ~n180 & ~n187;
  assign n189 = ~pi3  & ~n188;
  assign n190 = pi3  & pi8 ;
  assign n191 = ~pi2  & ~n190;
  assign n192 = ~pi0  & ~n191;
  assign n193 = pi5  & n143;
  assign n194 = ~pi3  & ~pi8 ;
  assign n195 = ~n152 & ~n194;
  assign n196 = pi0  & n195;
  assign n197 = ~n193 & ~n196;
  assign n198 = ~pi1  & ~n197;
  assign n199 = ~pi2  & pi8 ;
  assign n200 = pi0  & n199;
  assign n201 = pi0  & ~pi5 ;
  assign n202 = ~n163 & ~n201;
  assign n203 = ~n200 & n202;
  assign n204 = pi1  & ~n203;
  assign n205 = ~n192 & ~n204;
  assign n206 = ~n198 & n205;
  assign n207 = ~pi6  & ~n206;
  assign n208 = ~pi1  & ~pi8 ;
  assign n209 = ~pi2  & ~n208;
  assign n210 = ~pi1  & pi8 ;
  assign n211 = pi6  & n210;
  assign n212 = ~n209 & ~n211;
  assign n213 = pi3  & ~n212;
  assign n214 = ~pi0  & pi8 ;
  assign n215 = pi0  & pi1 ;
  assign n216 = ~pi1  & ~pi6 ;
  assign n217 = ~pi2  & ~n214;
  assign n218 = ~n215 & ~n216;
  assign n219 = n217 & n218;
  assign n220 = ~n213 & ~n219;
  assign n221 = ~pi5  & ~n220;
  assign n222 = ~pi9  & ~n221;
  assign n223 = ~n207 & n222;
  assign n224 = ~pi1  & pi3 ;
  assign n225 = n143 & n224;
  assign n226 = ~n79 & ~n225;
  assign n227 = pi0  & ~n226;
  assign n228 = pi3  & n58;
  assign n229 = ~pi5  & ~n228;
  assign n230 = ~n52 & ~n229;
  assign n231 = ~n227 & ~n230;
  assign n232 = pi6  & ~n231;
  assign n233 = n182 & n228;
  assign n234 = pi9  & ~n233;
  assign n235 = ~n232 & n234;
  assign n236 = ~pi4  & ~n235;
  assign n237 = ~n223 & n236;
  assign n238 = ~n189 & ~n237;
  assign n239 = ~pi7  & ~n238;
  assign n240 = ~pi6  & n39;
  assign n241 = n47 & n199;
  assign n242 = n105 & ~n215;
  assign n243 = pi2  & ~n33;
  assign n244 = ~pi8  & ~n243;
  assign n245 = ~n242 & n244;
  assign n246 = ~n241 & ~n245;
  assign n247 = pi7  & ~n246;
  assign n248 = ~n35 & ~n247;
  assign n249 = ~pi4  & n240;
  assign n250 = ~n248 & n249;
  assign po1  = n239 | n250;
  assign n252 = ~pi8  & ~pi9 ;
  assign n253 = pi8  & pi9 ;
  assign n254 = ~n252 & ~n253;
  assign n255 = ~n70 & ~n254;
  assign n256 = pi2  & ~n255;
  assign n257 = ~pi5  & ~n97;
  assign n258 = pi5  & ~n252;
  assign n259 = ~n147 & n258;
  assign n260 = pi1  & ~n257;
  assign n261 = ~n259 & n260;
  assign n262 = ~n256 & ~n261;
  assign n263 = ~pi3  & ~n262;
  assign n264 = n53 & n210;
  assign n265 = pi5  & ~n224;
  assign n266 = ~pi2  & n252;
  assign n267 = ~n265 & n266;
  assign n268 = ~n264 & ~n267;
  assign n269 = pi0  & ~n268;
  assign n270 = ~n263 & ~n269;
  assign n271 = ~pi6  & ~n270;
  assign n272 = pi6  & ~n42;
  assign n273 = ~n47 & ~n272;
  assign n274 = pi8  & ~n273;
  assign n275 = pi1  & pi9 ;
  assign n276 = ~n70 & ~n275;
  assign n277 = n194 & ~n276;
  assign n278 = ~n274 & ~n277;
  assign n279 = ~pi2  & ~n278;
  assign n280 = pi8  & ~n34;
  assign n281 = pi2  & n275;
  assign n282 = ~n210 & ~n281;
  assign n283 = pi6  & ~n282;
  assign n284 = pi2  & n252;
  assign n285 = ~n280 & ~n284;
  assign n286 = ~n283 & n285;
  assign n287 = pi3  & ~n286;
  assign n288 = ~n279 & ~n287;
  assign n289 = n201 & ~n288;
  assign n290 = ~n271 & ~n289;
  assign n291 = ~pi4  & ~n290;
  assign n292 = pi6  & ~pi8 ;
  assign n293 = ~n253 & ~n292;
  assign n294 = ~pi5  & ~n293;
  assign n295 = ~pi2  & n124;
  assign n296 = ~n294 & n295;
  assign n297 = pi4  & ~n296;
  assign n298 = pi3  & ~n199;
  assign n299 = pi5  & ~n298;
  assign n300 = pi2  & ~pi5 ;
  assign n301 = pi3  & ~n300;
  assign n302 = pi8  & ~n301;
  assign n303 = ~n299 & ~n302;
  assign n304 = pi1  & ~n303;
  assign n305 = ~pi5  & pi6 ;
  assign n306 = ~pi3  & n305;
  assign n307 = n208 & n306;
  assign n308 = ~n304 & ~n307;
  assign n309 = ~pi9  & ~n308;
  assign n310 = pi1  & pi8 ;
  assign n311 = pi6  & ~n310;
  assign n312 = ~pi9  & ~n311;
  assign n313 = ~pi2  & ~n312;
  assign n314 = ~pi8  & n42;
  assign n315 = ~n313 & ~n314;
  assign n316 = pi3  & ~n315;
  assign n317 = ~pi3  & pi9 ;
  assign n318 = pi1  & n317;
  assign n319 = n292 & n318;
  assign n320 = pi3  & ~pi9 ;
  assign n321 = pi3  & ~pi8 ;
  assign n322 = ~n47 & ~n321;
  assign n323 = ~pi6  & ~n320;
  assign n324 = ~n322 & n323;
  assign n325 = pi2  & ~n125;
  assign n326 = pi1  & ~n325;
  assign n327 = pi5  & ~n191;
  assign n328 = ~n326 & n327;
  assign n329 = ~pi4  & ~n319;
  assign n330 = ~n324 & n329;
  assign n331 = ~n328 & n330;
  assign n332 = ~n316 & n331;
  assign n333 = ~n309 & n332;
  assign n334 = ~pi0  & ~n297;
  assign n335 = ~n333 & n334;
  assign n336 = ~n291 & ~n335;
  assign n337 = ~pi7  & ~n336;
  assign n338 = pi7  & n253;
  assign n339 = pi0  & ~n338;
  assign n340 = n41 & ~n339;
  assign n341 = n45 & n208;
  assign n342 = ~n340 & ~n341;
  assign n343 = ~pi5  & ~pi6 ;
  assign n344 = ~pi4  & n52;
  assign n345 = n343 & n344;
  assign n346 = ~n342 & n345;
  assign po2  = n337 | n346;
  assign n348 = pi2  & n305;
  assign n349 = pi5  & pi9 ;
  assign n350 = pi8  & n349;
  assign n351 = ~pi6  & n350;
  assign n352 = ~n151 & ~n351;
  assign n353 = pi2  & ~n352;
  assign n354 = ~pi3  & ~n292;
  assign n355 = ~n126 & ~n354;
  assign n356 = ~n353 & ~n355;
  assign n357 = pi1  & ~n356;
  assign n358 = pi6  & ~n52;
  assign n359 = ~n320 & ~n358;
  assign n360 = ~pi1  & ~n359;
  assign n361 = ~n348 & ~n360;
  assign n362 = ~n357 & n361;
  assign n363 = ~pi4  & ~n362;
  assign n364 = ~pi3  & pi4 ;
  assign n365 = ~pi5  & ~n253;
  assign n366 = ~n134 & ~n343;
  assign n367 = ~pi1  & ~pi2 ;
  assign n368 = n364 & n367;
  assign n369 = ~n365 & n368;
  assign n370 = ~n366 & n369;
  assign n371 = ~n363 & ~n370;
  assign n372 = ~pi0  & ~n371;
  assign n373 = ~pi9  & n305;
  assign n374 = n310 & n373;
  assign n375 = pi2  & ~n195;
  assign n376 = ~pi2  & pi5 ;
  assign n377 = pi8  & n376;
  assign n378 = ~n375 & ~n377;
  assign n379 = ~pi9  & ~n378;
  assign n380 = pi5  & n164;
  assign n381 = ~pi3  & ~n380;
  assign n382 = ~pi2  & ~n381;
  assign n383 = ~pi6  & ~n321;
  assign n384 = pi3  & ~pi5 ;
  assign n385 = ~n383 & ~n384;
  assign n386 = ~n382 & ~n385;
  assign n387 = ~n379 & n386;
  assign n388 = pi1  & ~n387;
  assign n389 = n193 & n216;
  assign n390 = ~n306 & ~n389;
  assign n391 = ~pi9  & ~n390;
  assign n392 = ~n388 & ~n391;
  assign n393 = pi0  & ~n392;
  assign n394 = ~n28 & ~n170;
  assign n395 = ~pi2  & ~n394;
  assign n396 = ~pi6  & ~n349;
  assign n397 = pi5  & pi8 ;
  assign n398 = ~n275 & ~n397;
  assign n399 = n396 & ~n398;
  assign n400 = ~n395 & ~n399;
  assign n401 = pi3  & ~n400;
  assign n402 = pi3  & ~pi6 ;
  assign n403 = pi2  & n402;
  assign n404 = ~n52 & n305;
  assign n405 = ~n403 & ~n404;
  assign n406 = pi9  & ~n405;
  assign n407 = ~n373 & ~n402;
  assign n408 = ~pi8  & ~n407;
  assign n409 = ~n406 & ~n408;
  assign n410 = ~pi1  & ~n409;
  assign n411 = ~n374 & ~n401;
  assign n412 = ~n410 & n411;
  assign n413 = ~n393 & n412;
  assign n414 = ~pi4  & ~n413;
  assign n415 = ~n372 & ~n414;
  assign po3  = ~pi7  & ~n415;
  assign n417 = ~pi4  & n243;
  assign n418 = pi3  & ~pi4 ;
  assign n419 = ~n364 & ~n418;
  assign n420 = n181 & ~n419;
  assign n421 = ~n417 & ~n420;
  assign n422 = ~pi7  & n134;
  assign po4  = ~n421 & n422;
  assign n424 = ~n181 & n418;
  assign n425 = n181 & n364;
  assign n426 = ~n424 & ~n425;
  assign po5  = n422 & ~n426;
  assign n428 = pi4  & n33;
  assign n429 = n52 & n428;
  assign n430 = ~n134 & ~n429;
  assign n431 = ~pi7  & ~n430;
  assign n432 = pi7  & ~pi9 ;
  assign n433 = pi8  & ~n432;
  assign n434 = n86 & ~n433;
  assign n435 = ~n111 & ~n434;
  assign n436 = ~pi0  & ~n435;
  assign n437 = pi1  & n147;
  assign n438 = ~n252 & ~n437;
  assign n439 = ~pi2  & pi7 ;
  assign n440 = ~n438 & n439;
  assign n441 = ~n436 & ~n440;
  assign n442 = n343 & ~n441;
  assign n443 = pi2  & pi8 ;
  assign n444 = ~n143 & ~n443;
  assign n445 = pi6  & ~n254;
  assign n446 = ~n444 & n445;
  assign n447 = ~pi1  & ~pi5 ;
  assign n448 = pi2  & ~n447;
  assign n449 = n128 & ~n448;
  assign n450 = pi5  & n275;
  assign n451 = ~n449 & ~n450;
  assign n452 = pi0  & ~n451;
  assign n453 = ~pi0  & pi2 ;
  assign n454 = ~n28 & n453;
  assign n455 = ~n452 & ~n454;
  assign n456 = pi8  & ~n455;
  assign n457 = pi9  & n453;
  assign n458 = ~n71 & ~n457;
  assign n459 = pi5  & ~n458;
  assign n460 = ~n446 & ~n459;
  assign n461 = ~n456 & n460;
  assign n462 = ~pi7  & ~n461;
  assign n463 = ~n442 & ~n462;
  assign n464 = ~pi3  & ~n463;
  assign n465 = n40 & n443;
  assign n466 = ~pi2  & ~pi9 ;
  assign n467 = ~pi0  & ~n292;
  assign n468 = ~n397 & n466;
  assign n469 = ~n467 & n468;
  assign n470 = ~n465 & ~n469;
  assign n471 = ~pi1  & ~n470;
  assign n472 = n78 & n376;
  assign n473 = ~pi6  & ~n300;
  assign n474 = n40 & ~n473;
  assign n475 = ~n472 & ~n474;
  assign n476 = ~pi8  & ~n475;
  assign n477 = pi2  & ~n252;
  assign n478 = ~n147 & ~n477;
  assign n479 = pi6  & ~n478;
  assign n480 = ~n476 & ~n479;
  assign n481 = pi1  & ~n480;
  assign n482 = n92 & ~n453;
  assign n483 = pi0  & n156;
  assign n484 = ~pi2  & n483;
  assign n485 = ~n482 & ~n484;
  assign n486 = pi9  & ~n485;
  assign n487 = ~pi0  & ~pi6 ;
  assign n488 = ~n208 & n487;
  assign n489 = ~n58 & ~n488;
  assign n490 = n276 & ~n489;
  assign n491 = ~pi1  & ~n252;
  assign n492 = pi0  & ~n491;
  assign n493 = ~n47 & n492;
  assign n494 = ~n490 & ~n493;
  assign n495 = ~pi5  & ~n494;
  assign n496 = ~pi0  & ~pi8 ;
  assign n497 = n47 & ~n201;
  assign n498 = ~n496 & n497;
  assign n499 = ~n486 & ~n498;
  assign n500 = ~n495 & n499;
  assign n501 = pi3  & ~n500;
  assign n502 = ~n471 & ~n481;
  assign n503 = ~n501 & n502;
  assign n504 = ~pi7  & ~n503;
  assign n505 = ~n464 & ~n504;
  assign n506 = ~pi4  & ~n505;
  assign po6  = ~n431 & ~n506;
  assign n508 = n128 & n194;
  assign n509 = n214 & n402;
  assign n510 = ~n292 & ~n509;
  assign n511 = pi9  & ~n510;
  assign n512 = ~pi8  & ~n153;
  assign n513 = pi0  & ~n402;
  assign n514 = ~n131 & ~n513;
  assign n515 = ~n512 & ~n514;
  assign n516 = ~n511 & ~n515;
  assign n517 = ~pi2  & ~n516;
  assign n518 = pi3  & ~n253;
  assign n519 = ~n146 & ~n518;
  assign n520 = ~pi6  & ~n519;
  assign n521 = ~pi3  & n253;
  assign n522 = ~n520 & ~n521;
  assign n523 = pi2  & ~n522;
  assign n524 = ~n508 & ~n517;
  assign n525 = ~n523 & n524;
  assign n526 = pi1  & ~n525;
  assign n527 = n171 & ~n254;
  assign n528 = ~pi6  & ~n253;
  assign n529 = n105 & n528;
  assign n530 = ~n527 & ~n529;
  assign n531 = pi3  & ~n530;
  assign n532 = ~pi0  & n143;
  assign n533 = ~n483 & ~n532;
  assign n534 = ~pi9  & ~n533;
  assign n535 = ~pi6  & ~n194;
  assign n536 = n477 & ~n535;
  assign n537 = ~n534 & ~n536;
  assign n538 = ~n531 & n537;
  assign n539 = ~pi1  & ~n538;
  assign n540 = pi3  & n143;
  assign n541 = n131 & n540;
  assign n542 = ~n539 & ~n541;
  assign n543 = ~n526 & n542;
  assign n544 = ~pi5  & ~n543;
  assign n545 = pi0  & ~n97;
  assign n546 = ~n466 & n545;
  assign n547 = ~pi9  & n163;
  assign n548 = ~n546 & ~n547;
  assign n549 = pi8  & ~n548;
  assign n550 = n97 & n182;
  assign n551 = ~n549 & ~n550;
  assign n552 = ~pi3  & ~n551;
  assign n553 = pi3  & pi5 ;
  assign n554 = ~n34 & ~n553;
  assign n555 = ~pi0  & ~n554;
  assign n556 = pi3  & n376;
  assign n557 = ~n555 & ~n556;
  assign n558 = ~pi8  & ~n557;
  assign n559 = n466 & n553;
  assign n560 = ~n558 & ~n559;
  assign n561 = ~n552 & n560;
  assign n562 = pi1  & ~n561;
  assign n563 = n54 & n284;
  assign n564 = pi2  & pi3 ;
  assign n565 = n254 & ~n564;
  assign n566 = ~pi2  & ~n54;
  assign n567 = pi5  & ~n566;
  assign n568 = ~n565 & n567;
  assign n569 = ~n563 & ~n568;
  assign n570 = ~pi1  & ~n569;
  assign n571 = n350 & n564;
  assign n572 = ~n570 & ~n571;
  assign n573 = ~n562 & n572;
  assign n574 = ~pi6  & ~n573;
  assign n575 = ~n544 & ~n574;
  assign n576 = ~pi7  & ~n575;
  assign n577 = n254 & n453;
  assign n578 = pi8  & n31;
  assign n579 = n432 & n578;
  assign n580 = ~n577 & ~n579;
  assign n581 = n124 & n343;
  assign n582 = ~n580 & n581;
  assign n583 = ~n576 & ~n582;
  assign n584 = ~pi4  & ~n583;
  assign n585 = ~pi5  & ~pi7 ;
  assign n586 = n425 & n585;
  assign n587 = ~pi6  & n586;
  assign po7  = ~n584 & ~n587;
  assign n589 = n124 & n201;
  assign n590 = ~n79 & ~n384;
  assign n591 = ~pi2  & ~n113;
  assign n592 = n590 & n591;
  assign n593 = ~n589 & ~n592;
  assign n594 = pi8  & ~n593;
  assign n595 = ~pi5  & ~n214;
  assign n596 = n58 & ~n553;
  assign n597 = ~n595 & n596;
  assign n598 = ~n594 & ~n597;
  assign n599 = ~pi9  & ~n598;
  assign n600 = ~n300 & ~n553;
  assign n601 = pi1  & ~n298;
  assign n602 = ~n600 & n601;
  assign n603 = ~n163 & n199;
  assign n604 = n224 & n603;
  assign n605 = ~n602 & ~n604;
  assign n606 = pi9  & ~n605;
  assign n607 = n70 & n376;
  assign n608 = ~n318 & ~n607;
  assign n609 = ~pi0  & ~n608;
  assign n610 = n276 & ~n447;
  assign n611 = n93 & ~n610;
  assign n612 = ~pi2  & ~n70;
  assign n613 = ~n317 & n612;
  assign n614 = n590 & n613;
  assign n615 = ~n609 & ~n611;
  assign n616 = ~n614 & n615;
  assign n617 = ~pi8  & ~n616;
  assign n618 = ~n599 & ~n606;
  assign n619 = ~n617 & n618;
  assign n620 = ~pi6  & ~n619;
  assign n621 = ~n47 & n214;
  assign n622 = n272 & ~n621;
  assign n623 = ~pi2  & ~n622;
  assign n624 = ~pi6  & ~n92;
  assign n625 = ~n492 & n624;
  assign n626 = n384 & ~n623;
  assign n627 = ~n625 & n626;
  assign n628 = ~n620 & ~n627;
  assign n629 = ~pi7  & ~n628;
  assign n630 = ~pi0  & ~n444;
  assign n631 = ~n200 & ~n630;
  assign n632 = ~pi9  & ~n631;
  assign n633 = ~pi8  & n457;
  assign n634 = ~n632 & ~n633;
  assign n635 = ~pi1  & ~n634;
  assign n636 = n275 & n532;
  assign n637 = ~n635 & ~n636;
  assign n638 = n240 & ~n637;
  assign n639 = ~n629 & ~n638;
  assign n640 = ~pi4  & ~n639;
  assign po8  = ~n586 & ~n640;
  assign n642 = pi4  & ~n295;
  assign n643 = n365 & n403;
  assign n644 = ~pi6  & ~n350;
  assign n645 = ~pi3  & ~n644;
  assign n646 = ~pi3  & ~n28;
  assign n647 = pi3  & ~n153;
  assign n648 = n214 & ~n647;
  assign n649 = ~n646 & ~n648;
  assign n650 = ~pi2  & ~n649;
  assign n651 = ~n643 & ~n645;
  assign n652 = ~n650 & n651;
  assign n653 = pi1  & ~n652;
  assign n654 = ~n343 & n364;
  assign n655 = n214 & ~n396;
  assign n656 = n647 & ~n655;
  assign n657 = ~pi2  & ~n654;
  assign n658 = ~n656 & n657;
  assign n659 = n93 & ~n252;
  assign n660 = ~n365 & n659;
  assign n661 = ~n658 & ~n660;
  assign n662 = ~pi1  & ~n661;
  assign n663 = n201 & n403;
  assign n664 = ~pi7  & ~n663;
  assign n665 = ~n491 & ~n664;
  assign n666 = pi7  & ~n93;
  assign n667 = ~pi7  & ~n295;
  assign n668 = pi0  & ~n667;
  assign n669 = ~pi5  & ~n93;
  assign n670 = pi6  & ~n669;
  assign n671 = ~n642 & ~n666;
  assign n672 = ~n670 & n671;
  assign n673 = ~n668 & n672;
  assign n674 = ~n665 & n673;
  assign n675 = ~n653 & n674;
  assign po9  = ~n662 & n675;
  assign n677 = pi8  & ~n41;
  assign n678 = pi2  & n418;
  assign n679 = ~n46 & n678;
  assign n680 = ~n677 & n679;
  assign n681 = ~n425 & ~n680;
  assign n682 = ~pi7  & n343;
  assign po10  = ~n681 & n682;
endmodule
