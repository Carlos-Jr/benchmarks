module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 ,
    pi139 , pi140 , pi141 , pi142 , pi143 , pi144 , pi145 ,
    pi146 , pi147 , pi148 , pi149 , pi150 , pi151 , pi152 ,
    pi153 , pi154 , pi155 , pi156 , pi157 , pi158 , pi159 ,
    pi160 , pi161 , pi162 , pi163 , pi164 , pi165 , pi166 ,
    pi167 , pi168 , pi169 , pi170 , pi171 , pi172 , pi173 ,
    pi174 , pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 , pi194 ,
    pi195 , pi196 , pi197 , pi198 , pi199 , pi200 , pi201 ,
    pi202 , pi203 , pi204 , pi205 , pi206 , pi207 , pi208 ,
    pi209 , pi210 , pi211 , pi212 , pi213 , pi214 , pi215 ,
    pi216 , pi217 , pi218 , pi219 , pi220 , pi221 , pi222 ,
    pi223 , pi224 , pi225 , pi226 , pi227 , pi228 , pi229 ,
    pi230 , pi231 , pi232 , pi233 , pi234 , pi235 , pi236 ,
    pi237 , pi238 , pi239 , pi240 , pi241 , pi242 , pi243 ,
    pi244 , pi245 , pi246 , pi247 , pi248 , pi249 , pi250 ,
    pi251 , pi252 , pi253 , pi254 , pi255 , pi256 , pi257 ,
    pi258 , pi259 , pi260 , pi261 , pi262 , pi263 , pi264 ,
    pi265 , pi266 , pi267 , pi268 , pi269 , pi270 , pi271 ,
    pi272 , pi273 , pi274 , pi275 , pi276 , pi277 , pi278 ,
    pi279 , pi280 , pi281 , pi282 , pi283 , pi284 , pi285 ,
    pi286 , pi287 , pi288 , pi289 , pi290 , pi291 , pi292 ,
    pi293 , pi294 , pi295 , pi296 , pi297 , pi298 , pi299 ,
    pi300 , pi301 , pi302 , pi303 , pi304 , pi305 , pi306 ,
    pi307 , pi308 , pi309 , pi310 , pi311 , pi312 , pi313 ,
    pi314 , pi315 , pi316 , pi317 , pi318 , pi319 , pi320 ,
    pi321 , pi322 , pi323 , pi324 , pi325 , pi326 , pi327 ,
    pi328 , pi329 , pi330 , pi331 , pi332 , pi333 , pi334 ,
    pi335 , pi336 , pi337 , pi338 , pi339 , pi340 , pi341 ,
    pi342 , pi343 , pi344 , pi345 , pi346 , pi347 , pi348 ,
    pi349 , pi350 , pi351 , pi352 , pi353 , pi354 , pi355 ,
    pi356 , pi357 , pi358 , pi359 , pi360 , pi361 , pi362 ,
    pi363 , pi364 , pi365 , pi366 , pi367 , pi368 , pi369 ,
    pi370 , pi371 , pi372 , pi373 , pi374 , pi375 , pi376 ,
    pi377 , pi378 , pi379 , pi380 , pi381 , pi382 , pi383 ,
    pi384 , pi385 , pi386 , pi387 , pi388 , pi389 , pi390 ,
    pi391 , pi392 , pi393 , pi394 , pi395 , pi396 , pi397 ,
    pi398 , pi399 , pi400 , pi401 , pi402 , pi403 , pi404 ,
    pi405 , pi406 , pi407 , pi408 , pi409 , pi410 , pi411 ,
    pi412 , pi413 , pi414 , pi415 , pi416 , pi417 , pi418 ,
    pi419 , pi420 , pi421 , pi422 , pi423 , pi424 , pi425 ,
    pi426 , pi427 , pi428 , pi429 , pi430 , pi431 , pi432 ,
    pi433 , pi434 , pi435 , pi436 , pi437 , pi438 , pi439 ,
    pi440 , pi441 , pi442 , pi443 , pi444 , pi445 , pi446 ,
    pi447 , pi448 , pi449 , pi450 , pi451 , pi452 , pi453 ,
    pi454 , pi455 , pi456 , pi457 , pi458 , pi459 , pi460 ,
    pi461 , pi462 , pi463 , pi464 , pi465 , pi466 , pi467 ,
    pi468 , pi469 , pi470 , pi471 , pi472 , pi473 , pi474 ,
    pi475 , pi476 , pi477 , pi478 , pi479 , pi480 , pi481 ,
    pi482 , pi483 , pi484 , pi485 , pi486 , pi487 , pi488 ,
    pi489 , pi490 , pi491 , pi492 , pi493 , pi494 , pi495 ,
    pi496 , pi497 , pi498 , pi499 , pi500 , pi501 , pi502 ,
    pi503 , pi504 , pi505 , pi506 , pi507 , pi508 , pi509 ,
    pi510 , pi511 , pi512 , pi513 , pi514 , pi515 , pi516 ,
    pi517 , pi518 , pi519 , pi520 , pi521 , pi522 , pi523 ,
    pi524 , pi525 , pi526 , pi527 , pi528 , pi529 , pi530 ,
    pi531 , pi532 , pi533 , pi534 , pi535 , pi536 , pi537 ,
    pi538 , pi539 , pi540 , pi541 , pi542 , pi543 , pi544 ,
    pi545 , pi546 , pi547 , pi548 , pi549 , pi550 , pi551 ,
    pi552 , pi553 , pi554 , pi555 , pi556 , pi557 , pi558 ,
    pi559 , pi560 , pi561 , pi562 , pi563 , pi564 , pi565 ,
    pi566 , pi567 , pi568 , pi569 , pi570 , pi571 , pi572 ,
    pi573 , pi574 , pi575 , pi576 , pi577 , pi578 , pi579 ,
    pi580 , pi581 , pi582 , pi583 , pi584 , pi585 , pi586 ,
    pi587 , pi588 , pi589 , pi590 , pi591 , pi592 , pi593 ,
    pi594 , pi595 , pi596 , pi597 , pi598 , pi599 , pi600 ,
    pi601 , pi602 , pi603 , pi604 , pi605 , pi606 , pi607 ,
    pi608 , pi609 , pi610 , pi611 , pi612 , pi613 , pi614 ,
    pi615 , pi616 , pi617 , pi618 , pi619 , pi620 , pi621 ,
    pi622 , pi623 , pi624 , pi625 , pi626 , pi627 , pi628 ,
    pi629 , pi630 , pi631 , pi632 , pi633 , pi634 , pi635 ,
    pi636 , pi637 , pi638 , pi639 , pi640 , pi641 , pi642 ,
    pi643 , pi644 , pi645 , pi646 , pi647 , pi648 , pi649 ,
    pi650 , pi651 , pi652 , pi653 , pi654 , pi655 , pi656 ,
    pi657 , pi658 , pi659 , pi660 , pi661 , pi662 , pi663 ,
    pi664 , pi665 , pi666 , pi667 , pi668 , pi669 , pi670 ,
    pi671 , pi672 , pi673 , pi674 , pi675 , pi676 , pi677 ,
    pi678 , pi679 , pi680 , pi681 , pi682 , pi683 , pi684 ,
    pi685 , pi686 , pi687 , pi688 , pi689 , pi690 , pi691 ,
    pi692 , pi693 , pi694 , pi695 , pi696 , pi697 , pi698 ,
    pi699 , pi700 , pi701 , pi702 , pi703 , pi704 , pi705 ,
    pi706 , pi707 , pi708 , pi709 , pi710 , pi711 , pi712 ,
    pi713 , pi714 , pi715 , pi716 , pi717 , pi718 , pi719 ,
    pi720 , pi721 , pi722 , pi723 , pi724 , pi725 , pi726 ,
    pi727 , pi728 , pi729 , pi730 , pi731 , pi732 , pi733 ,
    pi734 , pi735 , pi736 , pi737 , pi738 , pi739 , pi740 ,
    pi741 , pi742 , pi743 , pi744 , pi745 , pi746 , pi747 ,
    pi748 , pi749 , pi750 , pi751 , pi752 , pi753 , pi754 ,
    pi755 , pi756 , pi757 , pi758 , pi759 , pi760 , pi761 ,
    pi762 , pi763 , pi764 , pi765 , pi766 , pi767 , pi768 ,
    pi769 , pi770 , pi771 , pi772 , pi773 , pi774 , pi775 ,
    pi776 , pi777 , pi778 , pi779 , pi780 , pi781 , pi782 ,
    pi783 , pi784 , pi785 , pi786 , pi787 , pi788 , pi789 ,
    pi790 , pi791 , pi792 , pi793 , pi794 , pi795 , pi796 ,
    pi797 , pi798 , pi799 , pi800 , pi801 , pi802 , pi803 ,
    pi804 , pi805 , pi806 , pi807 , pi808 , pi809 , pi810 ,
    pi811 , pi812 , pi813 , pi814 , pi815 , pi816 , pi817 ,
    pi818 , pi819 , pi820 , pi821 , pi822 , pi823 , pi824 ,
    pi825 , pi826 , pi827 , pi828 , pi829 , pi830 , pi831 ,
    pi832 , pi833 , pi834 , pi835 , pi836 , pi837 , pi838 ,
    pi839 , pi840 , pi841 , pi842 , pi843 , pi844 , pi845 ,
    pi846 , pi847 , pi848 , pi849 , pi850 , pi851 , pi852 ,
    pi853 , pi854 , pi855 , pi856 , pi857 , pi858 , pi859 ,
    pi860 , pi861 , pi862 , pi863 , pi864 , pi865 , pi866 ,
    pi867 , pi868 , pi869 , pi870 , pi871 , pi872 , pi873 ,
    pi874 , pi875 , pi876 , pi877 , pi878 , pi879 , pi880 ,
    pi881 , pi882 , pi883 , pi884 , pi885 , pi886 , pi887 ,
    pi888 , pi889 , pi890 , pi891 , pi892 , pi893 , pi894 ,
    pi895 , pi896 , pi897 , pi898 , pi899 , pi900 , pi901 ,
    pi902 , pi903 , pi904 , pi905 , pi906 , pi907 , pi908 ,
    pi909 , pi910 , pi911 , pi912 , pi913 , pi914 , pi915 ,
    pi916 , pi917 , pi918 , pi919 , pi920 , pi921 , pi922 ,
    pi923 , pi924 , pi925 , pi926 , pi927 , pi928 , pi929 ,
    pi930 , pi931 , pi932 , pi933 , pi934 , pi935 , pi936 ,
    pi937 , pi938 , pi939 , pi940 , pi941 , pi942 , pi943 ,
    pi944 , pi945 , pi946 , pi947 , pi948 , pi949 , pi950 ,
    pi951 , pi952 , pi953 , pi954 , pi955 , pi956 , pi957 ,
    pi958 , pi959 , pi960 , pi961 , pi962 , pi963 , pi964 ,
    pi965 , pi966 , pi967 , pi968 , pi969 , pi970 , pi971 ,
    pi972 , pi973 , pi974 , pi975 , pi976 , pi977 , pi978 ,
    pi979 , pi980 , pi981 , pi982 , pi983 , pi984 , pi985 ,
    pi986 , pi987 , pi988 , pi989 , pi990 , pi991 , pi992 ,
    pi993 , pi994 , pi995 , pi996 , pi997 , pi998 , pi999 ,
    pi1000 ,
    po0  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 , pi130 ,
    pi131 , pi132 , pi133 , pi134 , pi135 , pi136 , pi137 ,
    pi138 , pi139 , pi140 , pi141 , pi142 , pi143 , pi144 ,
    pi145 , pi146 , pi147 , pi148 , pi149 , pi150 , pi151 ,
    pi152 , pi153 , pi154 , pi155 , pi156 , pi157 , pi158 ,
    pi159 , pi160 , pi161 , pi162 , pi163 , pi164 , pi165 ,
    pi166 , pi167 , pi168 , pi169 , pi170 , pi171 , pi172 ,
    pi173 , pi174 , pi175 , pi176 , pi177 , pi178 , pi179 ,
    pi180 , pi181 , pi182 , pi183 , pi184 , pi185 , pi186 ,
    pi187 , pi188 , pi189 , pi190 , pi191 , pi192 , pi193 ,
    pi194 , pi195 , pi196 , pi197 , pi198 , pi199 , pi200 ,
    pi201 , pi202 , pi203 , pi204 , pi205 , pi206 , pi207 ,
    pi208 , pi209 , pi210 , pi211 , pi212 , pi213 , pi214 ,
    pi215 , pi216 , pi217 , pi218 , pi219 , pi220 , pi221 ,
    pi222 , pi223 , pi224 , pi225 , pi226 , pi227 , pi228 ,
    pi229 , pi230 , pi231 , pi232 , pi233 , pi234 , pi235 ,
    pi236 , pi237 , pi238 , pi239 , pi240 , pi241 , pi242 ,
    pi243 , pi244 , pi245 , pi246 , pi247 , pi248 , pi249 ,
    pi250 , pi251 , pi252 , pi253 , pi254 , pi255 , pi256 ,
    pi257 , pi258 , pi259 , pi260 , pi261 , pi262 , pi263 ,
    pi264 , pi265 , pi266 , pi267 , pi268 , pi269 , pi270 ,
    pi271 , pi272 , pi273 , pi274 , pi275 , pi276 , pi277 ,
    pi278 , pi279 , pi280 , pi281 , pi282 , pi283 , pi284 ,
    pi285 , pi286 , pi287 , pi288 , pi289 , pi290 , pi291 ,
    pi292 , pi293 , pi294 , pi295 , pi296 , pi297 , pi298 ,
    pi299 , pi300 , pi301 , pi302 , pi303 , pi304 , pi305 ,
    pi306 , pi307 , pi308 , pi309 , pi310 , pi311 , pi312 ,
    pi313 , pi314 , pi315 , pi316 , pi317 , pi318 , pi319 ,
    pi320 , pi321 , pi322 , pi323 , pi324 , pi325 , pi326 ,
    pi327 , pi328 , pi329 , pi330 , pi331 , pi332 , pi333 ,
    pi334 , pi335 , pi336 , pi337 , pi338 , pi339 , pi340 ,
    pi341 , pi342 , pi343 , pi344 , pi345 , pi346 , pi347 ,
    pi348 , pi349 , pi350 , pi351 , pi352 , pi353 , pi354 ,
    pi355 , pi356 , pi357 , pi358 , pi359 , pi360 , pi361 ,
    pi362 , pi363 , pi364 , pi365 , pi366 , pi367 , pi368 ,
    pi369 , pi370 , pi371 , pi372 , pi373 , pi374 , pi375 ,
    pi376 , pi377 , pi378 , pi379 , pi380 , pi381 , pi382 ,
    pi383 , pi384 , pi385 , pi386 , pi387 , pi388 , pi389 ,
    pi390 , pi391 , pi392 , pi393 , pi394 , pi395 , pi396 ,
    pi397 , pi398 , pi399 , pi400 , pi401 , pi402 , pi403 ,
    pi404 , pi405 , pi406 , pi407 , pi408 , pi409 , pi410 ,
    pi411 , pi412 , pi413 , pi414 , pi415 , pi416 , pi417 ,
    pi418 , pi419 , pi420 , pi421 , pi422 , pi423 , pi424 ,
    pi425 , pi426 , pi427 , pi428 , pi429 , pi430 , pi431 ,
    pi432 , pi433 , pi434 , pi435 , pi436 , pi437 , pi438 ,
    pi439 , pi440 , pi441 , pi442 , pi443 , pi444 , pi445 ,
    pi446 , pi447 , pi448 , pi449 , pi450 , pi451 , pi452 ,
    pi453 , pi454 , pi455 , pi456 , pi457 , pi458 , pi459 ,
    pi460 , pi461 , pi462 , pi463 , pi464 , pi465 , pi466 ,
    pi467 , pi468 , pi469 , pi470 , pi471 , pi472 , pi473 ,
    pi474 , pi475 , pi476 , pi477 , pi478 , pi479 , pi480 ,
    pi481 , pi482 , pi483 , pi484 , pi485 , pi486 , pi487 ,
    pi488 , pi489 , pi490 , pi491 , pi492 , pi493 , pi494 ,
    pi495 , pi496 , pi497 , pi498 , pi499 , pi500 , pi501 ,
    pi502 , pi503 , pi504 , pi505 , pi506 , pi507 , pi508 ,
    pi509 , pi510 , pi511 , pi512 , pi513 , pi514 , pi515 ,
    pi516 , pi517 , pi518 , pi519 , pi520 , pi521 , pi522 ,
    pi523 , pi524 , pi525 , pi526 , pi527 , pi528 , pi529 ,
    pi530 , pi531 , pi532 , pi533 , pi534 , pi535 , pi536 ,
    pi537 , pi538 , pi539 , pi540 , pi541 , pi542 , pi543 ,
    pi544 , pi545 , pi546 , pi547 , pi548 , pi549 , pi550 ,
    pi551 , pi552 , pi553 , pi554 , pi555 , pi556 , pi557 ,
    pi558 , pi559 , pi560 , pi561 , pi562 , pi563 , pi564 ,
    pi565 , pi566 , pi567 , pi568 , pi569 , pi570 , pi571 ,
    pi572 , pi573 , pi574 , pi575 , pi576 , pi577 , pi578 ,
    pi579 , pi580 , pi581 , pi582 , pi583 , pi584 , pi585 ,
    pi586 , pi587 , pi588 , pi589 , pi590 , pi591 , pi592 ,
    pi593 , pi594 , pi595 , pi596 , pi597 , pi598 , pi599 ,
    pi600 , pi601 , pi602 , pi603 , pi604 , pi605 , pi606 ,
    pi607 , pi608 , pi609 , pi610 , pi611 , pi612 , pi613 ,
    pi614 , pi615 , pi616 , pi617 , pi618 , pi619 , pi620 ,
    pi621 , pi622 , pi623 , pi624 , pi625 , pi626 , pi627 ,
    pi628 , pi629 , pi630 , pi631 , pi632 , pi633 , pi634 ,
    pi635 , pi636 , pi637 , pi638 , pi639 , pi640 , pi641 ,
    pi642 , pi643 , pi644 , pi645 , pi646 , pi647 , pi648 ,
    pi649 , pi650 , pi651 , pi652 , pi653 , pi654 , pi655 ,
    pi656 , pi657 , pi658 , pi659 , pi660 , pi661 , pi662 ,
    pi663 , pi664 , pi665 , pi666 , pi667 , pi668 , pi669 ,
    pi670 , pi671 , pi672 , pi673 , pi674 , pi675 , pi676 ,
    pi677 , pi678 , pi679 , pi680 , pi681 , pi682 , pi683 ,
    pi684 , pi685 , pi686 , pi687 , pi688 , pi689 , pi690 ,
    pi691 , pi692 , pi693 , pi694 , pi695 , pi696 , pi697 ,
    pi698 , pi699 , pi700 , pi701 , pi702 , pi703 , pi704 ,
    pi705 , pi706 , pi707 , pi708 , pi709 , pi710 , pi711 ,
    pi712 , pi713 , pi714 , pi715 , pi716 , pi717 , pi718 ,
    pi719 , pi720 , pi721 , pi722 , pi723 , pi724 , pi725 ,
    pi726 , pi727 , pi728 , pi729 , pi730 , pi731 , pi732 ,
    pi733 , pi734 , pi735 , pi736 , pi737 , pi738 , pi739 ,
    pi740 , pi741 , pi742 , pi743 , pi744 , pi745 , pi746 ,
    pi747 , pi748 , pi749 , pi750 , pi751 , pi752 , pi753 ,
    pi754 , pi755 , pi756 , pi757 , pi758 , pi759 , pi760 ,
    pi761 , pi762 , pi763 , pi764 , pi765 , pi766 , pi767 ,
    pi768 , pi769 , pi770 , pi771 , pi772 , pi773 , pi774 ,
    pi775 , pi776 , pi777 , pi778 , pi779 , pi780 , pi781 ,
    pi782 , pi783 , pi784 , pi785 , pi786 , pi787 , pi788 ,
    pi789 , pi790 , pi791 , pi792 , pi793 , pi794 , pi795 ,
    pi796 , pi797 , pi798 , pi799 , pi800 , pi801 , pi802 ,
    pi803 , pi804 , pi805 , pi806 , pi807 , pi808 , pi809 ,
    pi810 , pi811 , pi812 , pi813 , pi814 , pi815 , pi816 ,
    pi817 , pi818 , pi819 , pi820 , pi821 , pi822 , pi823 ,
    pi824 , pi825 , pi826 , pi827 , pi828 , pi829 , pi830 ,
    pi831 , pi832 , pi833 , pi834 , pi835 , pi836 , pi837 ,
    pi838 , pi839 , pi840 , pi841 , pi842 , pi843 , pi844 ,
    pi845 , pi846 , pi847 , pi848 , pi849 , pi850 , pi851 ,
    pi852 , pi853 , pi854 , pi855 , pi856 , pi857 , pi858 ,
    pi859 , pi860 , pi861 , pi862 , pi863 , pi864 , pi865 ,
    pi866 , pi867 , pi868 , pi869 , pi870 , pi871 , pi872 ,
    pi873 , pi874 , pi875 , pi876 , pi877 , pi878 , pi879 ,
    pi880 , pi881 , pi882 , pi883 , pi884 , pi885 , pi886 ,
    pi887 , pi888 , pi889 , pi890 , pi891 , pi892 , pi893 ,
    pi894 , pi895 , pi896 , pi897 , pi898 , pi899 , pi900 ,
    pi901 , pi902 , pi903 , pi904 , pi905 , pi906 , pi907 ,
    pi908 , pi909 , pi910 , pi911 , pi912 , pi913 , pi914 ,
    pi915 , pi916 , pi917 , pi918 , pi919 , pi920 , pi921 ,
    pi922 , pi923 , pi924 , pi925 , pi926 , pi927 , pi928 ,
    pi929 , pi930 , pi931 , pi932 , pi933 , pi934 , pi935 ,
    pi936 , pi937 , pi938 , pi939 , pi940 , pi941 , pi942 ,
    pi943 , pi944 , pi945 , pi946 , pi947 , pi948 , pi949 ,
    pi950 , pi951 , pi952 , pi953 , pi954 , pi955 , pi956 ,
    pi957 , pi958 , pi959 , pi960 , pi961 , pi962 , pi963 ,
    pi964 , pi965 , pi966 , pi967 , pi968 , pi969 , pi970 ,
    pi971 , pi972 , pi973 , pi974 , pi975 , pi976 , pi977 ,
    pi978 , pi979 , pi980 , pi981 , pi982 , pi983 , pi984 ,
    pi985 , pi986 , pi987 , pi988 , pi989 , pi990 , pi991 ,
    pi992 , pi993 , pi994 , pi995 , pi996 , pi997 , pi998 ,
    pi999 , pi1000 ;
  output po0;
  wire n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062,
    n1063, n1064, n1065, n1066, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110,
    n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122,
    n1123, n1124, n1125, n1126, n1127, n1128,
    n1129, n1130, n1131, n1132, n1133, n1134,
    n1135, n1136, n1137, n1138, n1139, n1140,
    n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152,
    n1153, n1154, n1155, n1156, n1157, n1158,
    n1159, n1160, n1161, n1162, n1163, n1164,
    n1165, n1166, n1167, n1168, n1169, n1170,
    n1171, n1172, n1173, n1174, n1175, n1176,
    n1177, n1178, n1179, n1180, n1181, n1182,
    n1183, n1184, n1185, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1204, n1205, n1206,
    n1207, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254,
    n1255, n1256, n1257, n1258, n1259, n1260,
    n1261, n1262, n1263, n1264, n1265, n1266,
    n1267, n1268, n1269, n1270, n1271, n1272,
    n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1299, n1300, n1301, n1302,
    n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1336, n1337, n1338,
    n1339, n1340, n1341, n1342, n1343, n1344,
    n1345, n1346, n1347, n1348, n1349, n1350,
    n1351, n1352, n1353, n1354, n1355, n1356,
    n1357, n1358, n1359, n1360, n1361, n1362,
    n1363, n1364, n1365, n1366, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1384, n1385, n1386,
    n1387, n1388, n1389, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1419, n1420, n1421, n1422,
    n1423, n1424, n1425, n1426, n1427, n1428,
    n1429, n1430, n1431, n1432, n1433, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542,
    n1543, n1544, n1545, n1546, n1547, n1548,
    n1549, n1550, n1551, n1552, n1553, n1554,
    n1555, n1556, n1557, n1558, n1559, n1560,
    n1561, n1562, n1563, n1564, n1565, n1566,
    n1567, n1568, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1577, n1578,
    n1579, n1580, n1581, n1582, n1583, n1584,
    n1585, n1586, n1587, n1588, n1589, n1590,
    n1591, n1592, n1593, n1594, n1595, n1596,
    n1597, n1598, n1599, n1600, n1601, n1602,
    n1603, n1604, n1605, n1606, n1607, n1608,
    n1609, n1610, n1611, n1612, n1613, n1614,
    n1615, n1616, n1617, n1618, n1619, n1620,
    n1621, n1622, n1623, n1624, n1625, n1626,
    n1627, n1628, n1629, n1630, n1631, n1632,
    n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1640, n1641, n1642, n1643, n1644,
    n1645, n1646, n1647, n1648, n1649, n1650,
    n1651, n1652, n1653, n1654, n1655, n1656,
    n1657, n1658, n1659, n1660, n1661, n1662,
    n1663, n1664, n1665, n1666, n1667, n1668,
    n1669, n1670, n1671, n1672, n1673, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680,
    n1681, n1682, n1683, n1684, n1685, n1686,
    n1687, n1688, n1689, n1690, n1691, n1692,
    n1693, n1694, n1695, n1696, n1697, n1698,
    n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710,
    n1711, n1712, n1713, n1714, n1715, n1716,
    n1717, n1718, n1719, n1720, n1721, n1722,
    n1723, n1724, n1725, n1726, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782,
    n1783, n1784, n1785, n1786, n1787, n1788,
    n1789, n1790, n1791, n1792, n1793, n1794,
    n1795, n1796, n1797, n1798, n1799, n1800,
    n1801, n1802, n1803, n1804, n1805, n1806,
    n1807, n1808, n1809, n1810, n1811, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962,
    n1963, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1992,
    n1993, n1994, n1995, n1996, n1997, n1998,
    n1999, n2000, n2001, n2002, n2003, n2004,
    n2005, n2006, n2007, n2008, n2009, n2010,
    n2011, n2012, n2013, n2014, n2015, n2016,
    n2017, n2018, n2019, n2020, n2021, n2022,
    n2023, n2024, n2025, n2026, n2027, n2028,
    n2029, n2030, n2031, n2032, n2033, n2034,
    n2035, n2036, n2037, n2038, n2039, n2040,
    n2041, n2042, n2043, n2044, n2045, n2046,
    n2047, n2048, n2049, n2050, n2051, n2052,
    n2053, n2054, n2055, n2056, n2057, n2058,
    n2059, n2060, n2061, n2062, n2063, n2064,
    n2065, n2066, n2067, n2068, n2069, n2070,
    n2071, n2072, n2073, n2074, n2075, n2076,
    n2077, n2078, n2079, n2080, n2081, n2082,
    n2083, n2084, n2085, n2086, n2087, n2088,
    n2089, n2090, n2091, n2092, n2093, n2094,
    n2095, n2096, n2097, n2098, n2099, n2100,
    n2101, n2102, n2103, n2104, n2105, n2106,
    n2107, n2108, n2109, n2110, n2111, n2112,
    n2113, n2114, n2115, n2116, n2117, n2118,
    n2119, n2120, n2121, n2122, n2123, n2124,
    n2125, n2126, n2127, n2128, n2129, n2130,
    n2131, n2132, n2133, n2134, n2135, n2136,
    n2137, n2138, n2139, n2140, n2141, n2142,
    n2143, n2144, n2145, n2146, n2147, n2148,
    n2149, n2150, n2151, n2152, n2153, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202,
    n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2226,
    n2227, n2228, n2229, n2230, n2231, n2232,
    n2233, n2234, n2235, n2236, n2237, n2238,
    n2239, n2240, n2241, n2242, n2243, n2244,
    n2245, n2246, n2247, n2248, n2249, n2250,
    n2251, n2252, n2253, n2254, n2255, n2256,
    n2257, n2258, n2259, n2260, n2261, n2262,
    n2263, n2264, n2265, n2266, n2267, n2268,
    n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286,
    n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418,
    n2419, n2420, n2421, n2422, n2423, n2424,
    n2425, n2426, n2427, n2428, n2429, n2430,
    n2431, n2432, n2433, n2434, n2435, n2436,
    n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3290, n3291, n3292, n3293, n3294,
    n3295, n3296, n3297, n3298, n3299, n3300,
    n3301, n3302, n3303, n3304, n3305, n3306,
    n3307, n3308, n3309, n3310, n3311, n3312,
    n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330,
    n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3340, n3341, n3342,
    n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3356, n3357, n3358, n3359, n3360,
    n3361, n3362, n3363, n3364, n3365, n3366,
    n3367, n3368, n3369, n3370, n3371, n3372,
    n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384,
    n3385, n3386, n3387, n3388, n3389, n3390,
    n3391, n3392, n3393, n3394, n3395, n3396,
    n3397, n3398, n3399, n3400, n3401, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419, n3420,
    n3421, n3422, n3423, n3424, n3425, n3426,
    n3427, n3428, n3429, n3430, n3431, n3432,
    n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450,
    n3451, n3452, n3453, n3454, n3455, n3456,
    n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474,
    n3475, n3476, n3477, n3478, n3479, n3480,
    n3481, n3482, n3483, n3484, n3485, n3486,
    n3487, n3488, n3489, n3490, n3491, n3492,
    n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510,
    n3511, n3512, n3513, n3514, n3515, n3516,
    n3517, n3518, n3519, n3520, n3521, n3522,
    n3523, n3524, n3525, n3526, n3527, n3528,
    n3529, n3530, n3531, n3532, n3533, n3534,
    n3535, n3536, n3537, n3538, n3539, n3540,
    n3541, n3542, n3543, n3544, n3545, n3546,
    n3547, n3548, n3549, n3550, n3551, n3552,
    n3553, n3554, n3555, n3556, n3557, n3558,
    n3559, n3560, n3561, n3562, n3563, n3564,
    n3565, n3566, n3567, n3568, n3569, n3570,
    n3571, n3572, n3573, n3574, n3575, n3576,
    n3577, n3578, n3579, n3580, n3581, n3582,
    n3583, n3584, n3585, n3586, n3587, n3588,
    n3589, n3590, n3591, n3592, n3593, n3594,
    n3595, n3596, n3597, n3598, n3599, n3600,
    n3601, n3602, n3603, n3604, n3605, n3606,
    n3607, n3608, n3609, n3610, n3611, n3612,
    n3613, n3614, n3615, n3616, n3617, n3618,
    n3619, n3620, n3621, n3622, n3623, n3624,
    n3625, n3626, n3627, n3628, n3629, n3630,
    n3631, n3632, n3633, n3634, n3635, n3636,
    n3637, n3638, n3639, n3640, n3641, n3642,
    n3643, n3644, n3645, n3646, n3647, n3648,
    n3649, n3650, n3651, n3652, n3653, n3654,
    n3655, n3656, n3657, n3658, n3659, n3660,
    n3661, n3662, n3663, n3664, n3665, n3666,
    n3667, n3668, n3669, n3670, n3671, n3672,
    n3673, n3674, n3675, n3676, n3677, n3678,
    n3679, n3680, n3681, n3682, n3683, n3684,
    n3685, n3686, n3687, n3688, n3689, n3690,
    n3691, n3692, n3693, n3694, n3695, n3696,
    n3697, n3698, n3699, n3700, n3701, n3702,
    n3703, n3704, n3705, n3706, n3707, n3708,
    n3709, n3710, n3711, n3712, n3713, n3714,
    n3715, n3716, n3717, n3718, n3719, n3720,
    n3721, n3722, n3723, n3724, n3725, n3726,
    n3727, n3728, n3729, n3730, n3731, n3732,
    n3733, n3734, n3735, n3736, n3737, n3738,
    n3739, n3740, n3741, n3742, n3743, n3744,
    n3745, n3746, n3747, n3748, n3749, n3750,
    n3751, n3752, n3753, n3754, n3755, n3756,
    n3757, n3758, n3759, n3760, n3761, n3762,
    n3763, n3764, n3765, n3766, n3767, n3768,
    n3769, n3770, n3771, n3772, n3773, n3774,
    n3775, n3776, n3777, n3778, n3779, n3780,
    n3781, n3782, n3783, n3784, n3785, n3786,
    n3787, n3788, n3789, n3790, n3791, n3792,
    n3793, n3794, n3795, n3796, n3797, n3798,
    n3799, n3800, n3801, n3802, n3803, n3804,
    n3805, n3806, n3807, n3808, n3809, n3810,
    n3811, n3812, n3813, n3814, n3815, n3816,
    n3817, n3818, n3819, n3820, n3821, n3822,
    n3823, n3824, n3825, n3826, n3827, n3828,
    n3829, n3830, n3831, n3832, n3833, n3834,
    n3835, n3836, n3837, n3838, n3839, n3840,
    n3841, n3842, n3843, n3844, n3845, n3846,
    n3847, n3848, n3849, n3850, n3851, n3852,
    n3853, n3854, n3855, n3856, n3857, n3858,
    n3859, n3860, n3861, n3862, n3863, n3864,
    n3865, n3866, n3867, n3868, n3869, n3870,
    n3871, n3872, n3873, n3874, n3875, n3876,
    n3877, n3878, n3879, n3880, n3881, n3882,
    n3883, n3884, n3885, n3886, n3887, n3888,
    n3889, n3890, n3891, n3892, n3893, n3894,
    n3895, n3896, n3897, n3898, n3899, n3900,
    n3901, n3902, n3903, n3904, n3905, n3906,
    n3907, n3908, n3909, n3910, n3911, n3912,
    n3913, n3914, n3915, n3916, n3917, n3918,
    n3919, n3920, n3921, n3922, n3923, n3924,
    n3925, n3926, n3927, n3928, n3929, n3930,
    n3931, n3932, n3933, n3934, n3935, n3936,
    n3937, n3938, n3939, n3940, n3941, n3942,
    n3943, n3944, n3945, n3946, n3947, n3948,
    n3949, n3950, n3951, n3952, n3953, n3954,
    n3955, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3992, n3993, n3994, n3995, n3996,
    n3997, n3998, n3999, n4000, n4001, n4002,
    n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014,
    n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4023, n4024, n4025, n4026,
    n4027, n4028, n4029, n4030, n4031, n4032,
    n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044,
    n4045, n4046, n4047, n4048, n4049, n4050,
    n4051, n4052, n4053, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4062,
    n4063, n4064, n4065, n4066, n4067, n4068,
    n4069, n4070, n4071, n4072, n4073, n4074,
    n4075, n4076, n4077, n4078, n4079, n4080,
    n4081, n4082, n4083, n4084, n4085, n4086,
    n4087, n4088, n4089, n4090, n4091, n4092,
    n4093, n4094, n4095, n4096, n4097, n4098,
    n4099, n4100, n4101, n4102, n4103, n4104,
    n4105, n4106, n4107, n4108, n4109, n4110,
    n4111, n4112, n4113, n4114, n4115, n4116,
    n4117, n4118, n4119, n4120, n4121, n4122,
    n4123, n4124, n4125, n4126, n4127, n4128,
    n4129, n4130, n4131, n4132, n4133, n4134,
    n4135, n4136, n4137, n4138, n4139, n4140,
    n4141, n4142, n4143, n4144, n4145, n4146,
    n4147, n4148, n4149, n4150, n4151, n4152,
    n4153, n4154, n4155, n4156, n4157, n4158,
    n4159, n4160, n4161, n4162, n4163, n4164,
    n4165, n4166, n4167, n4168, n4169, n4170,
    n4171, n4172, n4173, n4174, n4175, n4176,
    n4177, n4178, n4179, n4180, n4181, n4182,
    n4183, n4184, n4185, n4186, n4187, n4188,
    n4189, n4190, n4191, n4192, n4193, n4194,
    n4195, n4196, n4197, n4198, n4199, n4200,
    n4201, n4202, n4203, n4204, n4205, n4206,
    n4207, n4208, n4209, n4210, n4211, n4212,
    n4213, n4214, n4215, n4216, n4217, n4218,
    n4219, n4220, n4221, n4222, n4223, n4224,
    n4225, n4226, n4227, n4228, n4229, n4230,
    n4231, n4232, n4233, n4234, n4235, n4236,
    n4237, n4238, n4239, n4240, n4241, n4242,
    n4243, n4244, n4245, n4246, n4247, n4248,
    n4249, n4250, n4251, n4252, n4253, n4254,
    n4255, n4256, n4257, n4258, n4259, n4260,
    n4261, n4262, n4263, n4264, n4265, n4266,
    n4267, n4268, n4269, n4270, n4271, n4272,
    n4273, n4274, n4275, n4276, n4277, n4278,
    n4279, n4280, n4281, n4282, n4283, n4284,
    n4285, n4286, n4287, n4288, n4289, n4290,
    n4291, n4292, n4293, n4294, n4295, n4296,
    n4297, n4298, n4299, n4300, n4301, n4302,
    n4303, n4304, n4305, n4306, n4307, n4308,
    n4309, n4310, n4311, n4312, n4313, n4314,
    n4315, n4316, n4317, n4318, n4319, n4320,
    n4321, n4322, n4323, n4324, n4325, n4326,
    n4327, n4328, n4329, n4330, n4331, n4332,
    n4333, n4334, n4335, n4336, n4337, n4338,
    n4339, n4340, n4341, n4342, n4343, n4344,
    n4345, n4346, n4347, n4348, n4349, n4350,
    n4351, n4352, n4353, n4354, n4355, n4356,
    n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596,
    n4597, n4598, n4599, n4600, n4601, n4602,
    n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662,
    n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686,
    n4687, n4688, n4689, n4690, n4691, n4692,
    n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710,
    n4711, n4712, n4713, n4714, n4715, n4716,
    n4717, n4718, n4719, n4720, n4721, n4722,
    n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734,
    n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752,
    n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764,
    n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776,
    n4777, n4778, n4779, n4780, n4781, n4782,
    n4783, n4784, n4785, n4786, n4787, n4788,
    n4789, n4790, n4791, n4792, n4793, n4794,
    n4795, n4796, n4797, n4798, n4799, n4800,
    n4801, n4802, n4803, n4804, n4805, n4806,
    n4807, n4808, n4809, n4810, n4811, n4812,
    n4813, n4814, n4815, n4816, n4817, n4818,
    n4819, n4820, n4821, n4822, n4823, n4824,
    n4825, n4826, n4827, n4828, n4829, n4830,
    n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848,
    n4849, n4850, n4851, n4852, n4853, n4854,
    n4855, n4856, n4857, n4858, n4859, n4860,
    n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878,
    n4879, n4880, n4881, n4882, n4883, n4884,
    n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4901, n4902,
    n4903, n4904, n4905, n4906, n4907, n4908,
    n4909, n4910, n4911, n4912, n4913, n4914,
    n4915, n4916, n4917, n4918, n4919, n4920,
    n4921, n4922, n4923, n4924, n4925, n4926,
    n4927, n4928, n4929, n4930, n4931, n4932,
    n4933, n4934, n4935, n4936, n4937, n4938,
    n4939, n4940, n4941, n4942, n4943, n4944,
    n4945, n4946, n4947, n4948, n4949, n4950,
    n4951, n4952, n4953, n4954, n4955, n4956,
    n4957, n4958, n4959, n4960, n4961, n4962,
    n4963, n4964, n4965, n4966, n4967, n4968,
    n4969, n4970, n4971, n4972, n4973, n4974,
    n4975, n4976, n4977, n4978, n4979, n4980,
    n4981, n4982, n4983, n4984, n4985, n4986,
    n4987, n4988, n4989, n4990, n4991, n4992,
    n4993, n4994, n4995, n4996, n4997, n4998,
    n4999, n5000, n5001, n5002, n5003, n5004,
    n5005, n5006, n5007, n5008, n5009, n5010,
    n5011, n5012, n5013, n5014, n5015, n5016,
    n5017, n5018, n5019, n5020, n5021, n5022,
    n5023, n5024, n5025, n5026, n5027, n5028,
    n5029, n5030, n5031, n5032, n5033, n5034,
    n5035, n5036, n5037, n5038, n5039, n5040,
    n5041, n5042, n5043, n5044, n5045, n5046,
    n5047, n5048, n5049, n5050, n5051, n5052,
    n5053, n5054, n5055, n5056, n5057, n5058,
    n5059, n5060, n5061, n5062, n5063, n5064,
    n5065, n5066, n5067, n5068, n5069, n5070,
    n5071, n5072, n5073, n5074, n5075, n5076,
    n5077, n5078, n5079, n5080, n5081, n5082,
    n5083, n5084, n5085, n5086, n5087, n5088,
    n5089, n5090, n5091, n5092, n5093, n5094,
    n5095, n5096, n5097, n5098, n5099, n5100,
    n5101, n5102, n5103, n5104, n5105, n5106,
    n5107, n5108, n5109, n5110, n5111, n5112,
    n5113, n5114, n5115, n5116, n5117, n5118,
    n5119, n5120, n5121, n5122, n5123, n5124,
    n5125, n5126, n5127, n5128, n5129, n5130,
    n5131, n5132, n5133, n5134, n5135, n5136,
    n5137, n5138, n5139, n5140, n5141, n5142,
    n5143, n5144, n5145, n5146, n5147, n5148,
    n5149, n5150, n5151, n5152, n5153, n5154,
    n5155, n5156, n5157, n5158, n5159, n5160,
    n5161, n5162, n5163, n5164, n5165, n5166,
    n5167, n5168, n5169, n5170, n5171, n5172,
    n5173, n5174, n5175, n5176, n5177, n5178,
    n5179, n5180, n5181, n5182, n5183, n5184,
    n5185, n5186, n5187, n5188, n5189, n5190,
    n5191, n5192, n5193, n5194, n5195, n5196,
    n5197, n5198, n5199, n5200, n5201, n5202,
    n5203, n5204, n5205, n5206, n5207, n5208,
    n5209, n5210, n5211, n5212, n5213, n5214,
    n5215, n5216, n5217, n5218, n5219, n5220,
    n5221, n5222, n5223, n5224, n5225, n5226,
    n5227, n5228, n5229, n5230, n5231, n5232,
    n5233, n5234, n5235, n5236, n5237, n5238,
    n5239, n5240, n5241, n5242, n5243, n5244,
    n5245, n5246, n5247, n5248, n5249, n5250,
    n5251, n5252, n5253, n5254, n5255, n5256,
    n5257, n5258, n5259, n5260, n5261, n5262,
    n5263, n5264, n5265, n5266, n5267, n5268,
    n5269, n5270, n5271, n5272, n5273, n5274,
    n5275, n5276, n5277, n5278, n5279, n5280,
    n5281, n5282, n5283, n5284, n5285, n5286,
    n5287, n5288, n5289, n5290, n5291, n5292,
    n5293, n5294, n5295, n5296, n5297, n5298,
    n5299, n5300, n5301, n5302, n5303, n5304,
    n5305, n5306, n5307, n5308, n5309, n5310,
    n5311, n5312, n5313, n5314, n5315, n5316,
    n5317, n5318, n5319, n5320, n5321, n5322,
    n5323, n5324, n5325, n5326, n5327, n5328,
    n5329, n5330, n5331, n5332, n5333, n5334,
    n5335, n5336, n5337, n5338, n5339, n5340,
    n5341, n5342, n5343, n5344, n5345, n5346,
    n5347, n5348, n5349, n5350, n5351, n5352,
    n5353, n5354, n5355, n5356, n5357, n5358,
    n5359, n5360, n5361, n5362, n5363, n5364,
    n5365, n5366, n5367, n5368, n5369, n5370,
    n5371, n5372, n5373, n5374, n5375, n5376,
    n5377, n5378, n5379, n5380, n5381, n5382,
    n5383, n5384, n5385, n5386, n5387, n5388,
    n5389, n5390, n5391, n5392, n5393, n5394,
    n5395, n5396, n5397, n5398, n5399, n5400,
    n5401, n5402, n5403, n5404, n5405, n5406,
    n5407, n5408, n5409, n5410, n5411, n5412,
    n5413, n5414, n5415, n5416, n5417, n5418,
    n5419, n5420, n5421, n5422, n5423, n5424,
    n5425, n5426, n5427, n5428, n5429, n5430,
    n5431, n5432, n5433, n5434, n5435, n5436,
    n5437, n5438, n5439, n5440, n5441, n5442,
    n5443, n5444, n5445, n5446, n5447, n5448,
    n5449, n5450, n5451, n5452, n5453, n5454,
    n5455, n5456, n5457, n5458, n5459, n5460,
    n5461, n5462, n5463, n5464, n5465, n5466,
    n5467, n5468, n5469, n5470, n5471, n5472,
    n5473, n5474, n5475, n5476, n5477, n5478,
    n5479, n5480, n5481, n5482, n5483, n5484,
    n5485, n5486, n5487, n5488, n5489, n5490,
    n5491, n5492, n5493, n5494, n5495, n5496,
    n5497, n5498, n5499, n5500, n5501, n5502,
    n5503, n5504, n5505, n5506, n5507, n5508,
    n5509, n5510, n5511, n5512, n5513, n5514,
    n5515, n5516, n5517, n5518, n5519, n5520,
    n5521, n5522, n5523, n5524, n5525, n5526,
    n5527, n5528, n5529, n5530, n5531, n5532,
    n5533, n5534, n5535, n5536, n5537, n5538,
    n5539, n5540, n5541, n5542, n5543, n5544,
    n5545, n5546, n5547, n5548, n5549, n5550,
    n5551, n5552, n5553, n5554, n5555, n5556,
    n5557, n5558, n5559, n5560, n5561, n5562,
    n5563, n5564, n5565, n5566, n5567, n5568,
    n5569, n5570, n5571, n5572, n5573, n5574,
    n5575, n5576, n5577, n5578, n5579, n5580,
    n5581, n5582, n5583, n5584, n5585, n5586,
    n5587, n5588, n5589, n5590, n5591, n5592,
    n5593, n5594, n5595, n5596, n5597, n5598,
    n5599, n5600, n5601, n5602, n5603, n5604,
    n5605, n5606, n5607, n5608, n5609, n5610,
    n5611, n5612, n5613, n5614, n5615, n5616,
    n5617, n5618, n5619, n5620, n5621, n5622,
    n5623, n5624, n5625, n5626, n5627, n5628,
    n5629, n5630, n5631, n5632, n5633, n5634,
    n5635, n5636, n5637, n5638, n5639, n5640,
    n5641, n5642, n5643, n5644, n5645, n5646,
    n5647, n5648, n5649, n5650, n5651, n5652,
    n5653, n5654, n5655, n5656, n5657, n5658,
    n5659, n5660, n5661, n5662, n5663, n5664,
    n5665, n5666, n5667, n5668, n5669, n5670,
    n5671, n5672, n5673, n5674, n5675, n5676,
    n5677, n5678, n5679, n5680, n5681, n5682,
    n5683, n5684, n5685, n5686, n5687, n5688,
    n5689, n5690, n5691, n5692, n5693, n5694,
    n5695, n5696, n5697, n5698, n5699, n5700,
    n5701, n5702, n5703, n5704, n5705, n5706,
    n5707, n5708, n5709, n5710, n5711, n5712,
    n5713, n5714, n5715, n5716, n5717, n5718,
    n5719, n5720, n5721, n5722, n5723, n5724,
    n5725, n5726, n5727, n5728, n5729, n5730,
    n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742,
    n5743, n5744, n5745, n5746, n5747, n5748,
    n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772,
    n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802,
    n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844,
    n5845, n5846, n5847, n5848, n5849, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874,
    n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904,
    n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934,
    n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946,
    n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964,
    n5965, n5966, n5967, n5968, n5969, n5970,
    n5971, n5972, n5973, n5974, n5975, n5976,
    n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994,
    n5995, n5996, n5997, n5998, n5999, n6000,
    n6001, n6002, n6003, n6004, n6005, n6006,
    n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030,
    n6031, n6032, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060,
    n6061, n6062, n6063, n6064, n6065, n6066,
    n6067, n6068, n6069, n6070, n6071, n6072,
    n6073, n6074, n6075, n6076, n6077, n6078,
    n6079, n6080, n6081, n6082, n6083, n6084,
    n6085, n6086, n6087, n6088, n6089, n6090,
    n6091, n6092, n6093, n6094, n6095, n6096,
    n6097, n6098, n6099, n6100, n6101, n6102,
    n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114,
    n6115, n6116, n6117, n6118, n6119, n6120,
    n6121, n6122, n6123, n6124, n6125, n6126,
    n6127, n6128, n6129, n6130, n6131, n6132,
    n6133, n6134, n6135, n6136, n6137, n6138,
    n6139, n6140, n6141, n6142, n6143, n6144,
    n6145, n6146, n6147, n6148, n6149, n6150,
    n6151, n6152, n6153, n6154, n6155, n6156,
    n6157, n6158, n6159, n6160, n6161, n6162,
    n6163, n6164, n6165, n6166, n6167, n6168,
    n6169, n6170, n6171, n6172, n6173, n6174,
    n6175, n6176, n6177, n6178, n6179, n6180,
    n6181, n6182, n6183, n6184, n6185, n6186,
    n6187, n6188, n6189, n6190, n6191, n6192,
    n6193, n6194, n6195, n6196, n6197, n6198,
    n6199, n6200, n6201, n6202, n6203, n6204,
    n6205, n6206, n6207, n6208, n6209, n6210,
    n6211, n6212, n6213, n6214, n6215, n6216,
    n6217, n6218, n6219, n6220, n6221, n6222,
    n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234,
    n6235, n6236, n6237, n6238, n6239, n6240,
    n6241, n6242, n6243, n6244, n6245, n6246,
    n6247, n6248, n6249, n6250, n6251, n6252,
    n6253, n6254, n6255, n6256, n6257, n6258,
    n6259, n6260, n6261, n6262, n6263, n6264,
    n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276,
    n6277, n6278, n6279, n6280, n6281, n6282,
    n6283, n6284, n6285, n6286, n6287, n6288,
    n6289, n6290, n6291, n6292, n6293, n6294,
    n6295, n6296, n6297, n6298, n6299, n6300,
    n6301, n6302, n6303, n6304, n6305, n6306,
    n6307, n6308, n6309, n6310, n6311, n6312,
    n6313, n6314, n6315, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6340, n6341, n6342,
    n6343, n6344, n6345, n6346, n6347, n6348,
    n6349, n6350, n6351, n6352, n6353, n6354,
    n6355, n6356, n6357, n6358, n6359, n6360,
    n6361, n6362, n6363, n6364, n6365, n6366,
    n6367, n6368, n6369, n6370, n6371, n6372,
    n6373, n6374, n6375, n6376, n6377, n6378,
    n6379, n6380, n6381, n6382, n6383, n6384,
    n6385, n6386, n6387, n6388, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546,
    n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570,
    n6571, n6572, n6573, n6574, n6575, n6576,
    n6577, n6578, n6579, n6580, n6581, n6582,
    n6583, n6584, n6585, n6586, n6587, n6588,
    n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600,
    n6601, n6602, n6603, n6604, n6605, n6606,
    n6607, n6608, n6609, n6610, n6611, n6612,
    n6613, n6614, n6615, n6616, n6617, n6618,
    n6619, n6620, n6621, n6622, n6623, n6624,
    n6625, n6626, n6627, n6628, n6629, n6630,
    n6631, n6632, n6633, n6634, n6635, n6636,
    n6637, n6638, n6639, n6640, n6641, n6642,
    n6643, n6644, n6645, n6646, n6647, n6648,
    n6649, n6650, n6651, n6652, n6653, n6654,
    n6655, n6656, n6657, n6658, n6659, n6660,
    n6661, n6662, n6663, n6664, n6665, n6666,
    n6667, n6668, n6669, n6670, n6671, n6672,
    n6673, n6674, n6675, n6676, n6677, n6678,
    n6679, n6680, n6681, n6682, n6683, n6684,
    n6685, n6686, n6687, n6688, n6689, n6690,
    n6691, n6692, n6693, n6694, n6695, n6696,
    n6697, n6698, n6699, n6700, n6701, n6702,
    n6703, n6704, n6705, n6706, n6707, n6708,
    n6709, n6710, n6711, n6712, n6713, n6714,
    n6715, n6716, n6717, n6718, n6719, n6720,
    n6721, n6722, n6723, n6724, n6725, n6726,
    n6727, n6728, n6729, n6730, n6731, n6732,
    n6733, n6734, n6735, n6736, n6737, n6738,
    n6739, n6740, n6741, n6742, n6743, n6744,
    n6745, n6746, n6747, n6748, n6749, n6750,
    n6751, n6752, n6753, n6754, n6755, n6756,
    n6757, n6758, n6759, n6760, n6761, n6762,
    n6763, n6764, n6765, n6766, n6767, n6768,
    n6769, n6770, n6771, n6772, n6773, n6774,
    n6775, n6776, n6777, n6778, n6779, n6780,
    n6781, n6782, n6783, n6784, n6785, n6786,
    n6787, n6788, n6789, n6790, n6791, n6792,
    n6793, n6794, n6795, n6796, n6797, n6798,
    n6799, n6800, n6801, n6802, n6803, n6804,
    n6805, n6806, n6807, n6808, n6809, n6810,
    n6811, n6812, n6813, n6814, n6815, n6816,
    n6817, n6818, n6819, n6820, n6821, n6822,
    n6823, n6824, n6825, n6826, n6827, n6828,
    n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6838, n6839, n6840,
    n6841, n6842, n6843, n6844, n6845, n6846,
    n6847, n6848, n6849, n6850, n6851, n6852,
    n6853, n6854, n6855, n6856, n6857, n6858,
    n6859, n6860, n6861, n6862, n6863, n6864,
    n6865, n6866, n6867, n6868, n6869, n6870,
    n6871, n6872, n6873, n6874, n6875, n6876,
    n6877, n6878, n6879, n6880, n6881, n6882,
    n6883, n6884, n6885, n6886, n6887, n6888,
    n6889, n6890, n6891, n6892, n6893, n6894,
    n6895, n6896, n6897, n6898, n6899, n6900,
    n6901, n6902, n6903, n6904, n6905, n6906,
    n6907, n6908, n6909, n6910, n6911, n6912,
    n6913, n6914, n6915, n6916, n6917, n6918,
    n6919, n6920, n6921, n6922, n6923, n6924,
    n6925, n6926, n6927, n6928, n6929, n6930,
    n6931, n6932, n6933, n6934, n6935, n6936,
    n6937, n6938, n6939, n6940, n6941, n6942,
    n6943, n6944, n6945, n6946, n6947, n6948,
    n6949, n6950, n6951, n6952, n6953, n6954,
    n6955, n6956, n6957, n6958, n6959, n6960,
    n6961, n6962, n6963, n6964, n6965, n6966,
    n6967, n6968, n6969, n6970, n6971, n6972,
    n6973, n6974, n6975, n6976, n6977, n6978,
    n6979, n6980, n6981, n6982, n6983, n6984,
    n6985, n6986, n6987, n6988, n6989, n6990,
    n6991, n6992, n6993, n6994, n6995, n6996,
    n6997, n6998, n6999, n7000, n7001, n7002,
    n7003, n7004, n7005, n7006, n7007, n7008,
    n7009, n7010, n7011, n7012, n7013, n7014,
    n7015, n7016, n7017, n7018, n7019, n7020,
    n7021, n7022, n7023, n7024, n7025, n7026,
    n7027, n7028, n7029, n7030, n7031, n7032,
    n7033, n7034, n7035, n7036, n7037, n7038,
    n7039, n7040, n7041, n7042, n7043, n7044,
    n7045, n7046, n7047, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062,
    n7063, n7064, n7065, n7066, n7067, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074,
    n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092,
    n7093, n7094, n7095, n7096, n7097, n7098,
    n7099, n7100, n7101, n7102, n7103, n7104,
    n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116,
    n7117, n7118, n7119, n7120, n7121, n7122,
    n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134,
    n7135, n7136, n7137, n7138, n7139, n7140,
    n7141, n7142, n7143, n7144, n7145, n7146,
    n7147, n7148, n7149, n7150, n7151, n7152,
    n7153, n7154, n7155, n7156, n7157, n7158,
    n7159, n7160, n7161, n7162, n7163, n7164,
    n7165, n7166, n7167, n7168, n7169, n7170,
    n7171, n7172, n7173, n7174, n7175, n7176,
    n7177, n7178, n7179, n7180, n7181, n7182,
    n7183, n7184, n7185, n7186, n7187, n7188,
    n7189, n7190, n7191, n7192, n7193, n7194,
    n7195, n7196, n7197, n7198, n7199, n7200,
    n7201, n7202, n7203, n7204, n7205, n7206,
    n7207, n7208, n7209, n7210, n7211, n7212,
    n7213, n7214, n7215, n7216, n7217, n7218,
    n7219, n7220, n7221, n7222, n7223, n7224,
    n7225, n7226, n7227, n7228, n7229, n7230,
    n7231, n7232, n7233, n7234, n7235, n7236,
    n7237, n7238, n7239, n7240, n7241, n7242,
    n7243, n7244, n7245, n7246, n7247, n7248,
    n7249, n7250, n7251, n7252, n7253, n7254,
    n7255, n7256, n7257, n7258, n7259, n7260,
    n7261, n7262, n7263, n7264, n7265, n7266,
    n7267, n7268, n7269, n7270, n7271, n7272,
    n7273, n7274, n7275, n7276, n7277, n7278,
    n7279, n7280, n7281, n7282, n7283, n7284,
    n7285, n7286, n7287, n7288, n7289, n7290,
    n7291, n7292, n7293, n7294, n7295, n7296,
    n7297, n7298, n7299, n7300, n7301, n7302,
    n7303, n7304, n7305, n7306, n7307, n7308,
    n7309, n7310, n7311, n7312, n7313, n7314,
    n7315, n7316, n7317, n7318, n7319, n7320,
    n7321, n7322, n7323, n7324, n7325, n7326,
    n7327, n7328, n7329, n7330, n7331, n7332,
    n7333, n7334, n7335, n7336, n7337, n7338,
    n7339, n7340, n7341, n7342, n7343, n7344,
    n7345, n7346, n7347, n7348, n7349, n7350,
    n7351, n7352, n7353, n7354, n7355, n7356,
    n7357, n7358, n7359, n7360, n7361, n7362,
    n7363, n7364, n7365, n7366, n7367, n7368,
    n7369, n7370, n7371, n7372, n7373, n7374,
    n7375, n7376, n7377, n7378, n7379, n7380,
    n7381, n7382, n7383, n7384, n7385, n7386,
    n7387, n7388, n7389, n7390, n7391, n7392,
    n7393, n7394, n7395, n7396, n7397, n7398,
    n7399, n7400, n7401, n7402, n7403, n7404,
    n7405, n7406, n7407, n7408, n7409, n7410,
    n7411, n7412, n7413, n7414, n7415, n7416,
    n7417, n7418, n7419, n7420, n7421, n7422,
    n7423, n7424, n7425, n7426, n7427, n7428,
    n7429, n7430, n7431, n7432, n7433, n7434,
    n7435, n7436, n7437, n7438, n7439, n7440,
    n7441, n7442, n7443, n7444, n7445, n7446,
    n7447, n7448, n7449, n7450, n7451, n7452,
    n7453, n7454, n7455, n7456, n7457, n7458,
    n7459, n7460, n7461, n7462, n7463, n7464,
    n7465, n7466, n7467, n7468, n7469, n7470,
    n7471, n7472, n7473, n7474, n7475, n7476,
    n7477, n7478, n7479, n7480, n7481, n7482,
    n7483, n7484, n7485, n7486, n7487, n7488,
    n7489, n7490, n7491, n7492, n7493, n7494,
    n7495, n7496, n7497, n7498, n7499, n7500,
    n7501, n7502, n7503, n7504, n7505, n7506,
    n7507, n7508, n7509, n7510, n7511, n7512,
    n7513, n7514, n7515, n7516, n7517, n7518,
    n7519, n7520, n7521, n7522, n7523, n7524,
    n7525, n7526, n7527, n7528, n7529, n7530,
    n7531, n7532, n7533, n7534, n7535, n7536,
    n7537, n7538, n7539, n7540, n7541, n7542,
    n7543, n7544, n7545, n7546, n7547, n7548,
    n7549, n7550, n7551, n7552, n7553, n7554,
    n7555, n7556, n7557, n7558, n7559, n7560,
    n7561, n7562, n7563, n7564, n7565, n7566,
    n7567, n7568, n7569, n7570, n7571, n7572,
    n7573, n7574, n7575, n7576, n7577, n7578,
    n7579, n7580, n7581, n7582, n7583, n7584,
    n7585, n7586, n7587, n7588, n7589, n7590,
    n7591, n7592, n7593, n7594, n7595, n7596,
    n7597, n7598, n7599, n7600, n7601, n7602,
    n7603, n7604, n7605, n7606, n7607, n7608,
    n7609, n7610, n7611, n7612, n7613, n7614,
    n7615, n7616, n7617, n7618, n7619, n7620,
    n7621, n7622, n7623, n7624, n7625, n7626,
    n7627, n7628, n7629, n7630, n7631, n7632,
    n7633, n7634, n7635, n7636, n7637, n7638,
    n7639, n7640, n7641, n7642, n7643, n7644,
    n7645, n7646, n7647, n7648, n7649, n7650,
    n7651, n7652, n7653, n7654, n7655, n7656,
    n7657, n7658, n7659, n7660, n7661, n7662,
    n7663, n7664, n7665, n7666, n7667, n7668,
    n7669, n7670, n7671, n7672, n7673, n7674,
    n7675, n7676, n7677, n7678, n7679, n7680,
    n7681, n7682, n7683, n7684, n7685, n7686,
    n7687, n7688, n7689, n7690, n7691, n7692,
    n7693, n7694, n7695, n7696, n7697, n7698,
    n7699, n7700, n7701, n7702, n7703, n7704,
    n7705, n7706, n7707, n7708, n7709, n7710,
    n7711, n7712, n7713, n7714, n7715, n7716,
    n7717, n7718, n7719, n7720, n7721, n7722,
    n7723, n7724, n7725, n7726, n7727, n7728,
    n7729, n7730, n7731, n7732, n7733, n7734,
    n7735, n7736, n7737, n7738, n7739, n7740,
    n7741, n7742, n7743, n7744, n7745, n7746,
    n7747, n7748, n7749, n7750, n7751, n7752,
    n7753, n7754, n7755, n7756, n7757, n7758,
    n7759, n7760, n7761, n7762, n7763, n7764,
    n7765, n7766, n7767, n7768, n7769, n7770,
    n7771, n7772, n7773, n7774, n7775, n7776,
    n7777, n7778, n7779, n7780, n7781, n7782,
    n7783, n7784, n7785, n7786, n7787, n7788,
    n7789, n7790, n7791, n7792, n7793, n7794,
    n7795, n7796, n7797, n7798, n7799, n7800,
    n7801, n7802, n7803, n7804, n7805, n7806,
    n7807, n7808, n7809, n7810, n7811, n7812,
    n7813, n7814, n7815, n7816, n7817, n7818,
    n7819, n7820, n7821, n7822, n7823, n7824,
    n7825, n7826, n7827, n7828, n7829, n7830,
    n7831, n7832, n7833, n7834, n7835, n7836,
    n7837, n7838, n7839, n7840, n7841, n7842,
    n7843, n7844, n7845, n7846, n7847, n7848,
    n7849, n7850, n7851, n7852, n7853, n7854,
    n7855, n7856, n7857, n7858, n7859, n7860,
    n7861, n7862, n7863, n7864, n7865, n7866,
    n7867, n7868, n7869, n7870, n7871, n7872,
    n7873, n7874, n7875, n7876, n7877, n7878,
    n7879, n7880, n7881, n7882, n7883, n7884,
    n7885, n7886, n7887, n7888, n7889, n7890,
    n7891, n7892, n7893, n7894, n7895, n7896,
    n7897, n7898, n7899, n7900, n7901, n7902,
    n7903, n7904, n7905, n7906, n7907, n7908,
    n7909, n7910, n7911, n7912, n7913, n7914,
    n7915, n7916, n7917, n7918, n7919, n7920,
    n7921, n7922, n7923, n7924, n7925, n7926,
    n7927, n7928, n7929, n7930, n7931, n7932,
    n7933, n7934, n7935, n7936, n7937, n7938,
    n7939, n7940, n7941, n7942, n7943, n7944,
    n7945, n7946, n7947, n7948, n7949, n7950,
    n7951, n7952, n7953, n7954, n7955, n7956,
    n7957, n7958, n7959, n7960, n7961, n7962,
    n7963, n7964, n7965, n7966, n7967, n7968,
    n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7977, n7978, n7979, n7980,
    n7981, n7982, n7983, n7984, n7985, n7986,
    n7987, n7988, n7989, n7990, n7991, n7992,
    n7993, n7994, n7995, n7996, n7997, n7998,
    n7999, n8000, n8001, n8002, n8003, n8004,
    n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016,
    n8017, n8018, n8019, n8020, n8021, n8022,
    n8023, n8024, n8025, n8026, n8027, n8028,
    n8029, n8030, n8031, n8032, n8033, n8034,
    n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046,
    n8047, n8048, n8049, n8050, n8051, n8052,
    n8053, n8054, n8055, n8056, n8057, n8058,
    n8059, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076,
    n8077, n8078, n8079, n8080, n8081, n8082,
    n8083, n8084, n8085, n8086, n8087, n8088,
    n8089, n8090, n8091, n8092, n8093, n8094,
    n8095, n8096, n8097, n8098, n8099, n8100,
    n8101, n8102, n8103, n8104, n8105, n8106,
    n8107, n8108, n8109, n8110, n8111, n8112,
    n8113, n8114, n8115, n8116, n8117, n8118,
    n8119, n8120, n8121, n8122, n8123, n8124,
    n8125, n8126, n8127, n8128, n8129, n8130,
    n8131, n8132, n8133, n8134, n8135, n8136,
    n8137, n8138, n8139, n8140, n8141, n8142,
    n8143, n8144, n8145, n8146, n8147, n8148,
    n8149, n8150, n8151, n8152, n8153, n8154,
    n8155, n8156, n8157, n8158, n8159, n8160,
    n8161, n8162, n8163, n8164, n8165, n8166,
    n8167, n8168, n8169, n8170, n8171, n8172,
    n8173, n8174, n8175, n8176, n8177, n8178,
    n8179, n8180, n8181, n8182, n8183, n8184,
    n8185, n8186, n8187, n8188, n8189, n8190,
    n8191, n8192, n8193, n8194, n8195, n8196,
    n8197, n8198, n8199, n8200, n8201, n8202,
    n8203, n8204, n8205, n8206, n8207, n8208,
    n8209, n8210, n8211, n8212, n8213, n8214,
    n8215, n8216, n8217, n8218, n8219, n8220,
    n8221, n8222, n8223, n8224, n8225, n8226,
    n8227, n8228, n8229, n8230, n8231, n8232,
    n8233, n8234, n8235, n8236, n8237, n8238,
    n8239, n8240, n8241, n8242, n8243, n8244,
    n8245, n8246, n8247, n8248, n8249, n8250,
    n8251, n8252, n8253, n8254, n8255, n8256,
    n8257, n8258, n8259, n8260, n8261, n8262,
    n8263, n8264, n8265, n8266, n8267, n8268,
    n8269, n8270, n8271, n8272, n8273, n8274,
    n8275, n8276, n8277, n8278, n8279, n8280,
    n8281, n8282, n8283, n8284, n8285, n8286,
    n8287, n8288, n8289, n8290, n8291, n8292,
    n8293, n8294, n8295, n8296, n8297, n8298,
    n8299, n8300, n8301, n8302, n8303, n8304,
    n8305, n8306, n8307, n8308, n8309, n8310,
    n8311, n8312, n8313, n8314, n8315, n8316,
    n8317, n8318, n8319, n8320, n8321, n8322,
    n8323, n8324, n8325, n8326, n8327, n8328,
    n8329, n8330, n8331, n8332, n8333, n8334,
    n8335, n8336, n8337, n8338, n8339, n8340,
    n8341, n8342, n8343, n8344, n8345, n8346,
    n8347, n8348, n8349, n8350, n8351, n8352,
    n8353, n8354, n8355, n8356, n8357, n8358,
    n8359, n8360, n8361, n8362, n8363, n8364,
    n8365, n8366, n8367, n8368, n8369, n8370,
    n8371, n8372, n8373, n8374, n8375, n8376,
    n8377, n8378, n8379, n8380, n8381, n8382,
    n8383, n8384, n8385, n8386, n8387, n8388,
    n8389, n8390, n8391, n8392, n8393, n8394,
    n8395, n8396, n8397, n8398, n8399, n8400,
    n8401, n8402, n8403, n8404, n8405, n8406,
    n8407, n8408, n8409, n8410, n8411, n8412,
    n8413, n8414, n8415, n8416, n8417, n8418,
    n8419, n8420, n8421, n8422, n8423, n8424,
    n8425, n8426, n8427, n8428, n8429, n8430,
    n8431, n8432, n8433, n8434, n8435, n8436,
    n8437, n8438, n8439, n8440, n8441, n8442,
    n8443, n8444, n8445, n8446, n8447, n8448,
    n8449, n8450, n8451, n8452, n8453, n8454,
    n8455, n8456, n8457, n8458, n8459, n8460,
    n8461, n8462, n8463, n8464, n8465, n8466,
    n8467, n8468, n8469, n8470, n8471, n8472,
    n8473, n8474, n8475, n8476, n8477, n8478,
    n8479, n8480, n8481, n8482, n8483, n8484,
    n8485, n8486, n8487, n8488, n8489, n8490,
    n8491, n8492, n8493, n8494, n8495, n8496,
    n8497, n8498, n8499, n8500, n8501, n8502,
    n8503, n8504, n8505, n8506, n8507, n8508,
    n8509, n8510, n8511, n8512, n8513, n8514,
    n8515, n8516, n8517, n8518, n8519, n8520,
    n8521, n8522, n8523, n8524, n8525, n8526,
    n8527, n8528, n8529, n8530, n8531, n8532,
    n8533, n8534, n8535, n8536, n8537, n8538,
    n8539, n8540, n8541, n8542, n8543, n8544,
    n8545, n8546, n8547, n8548, n8549, n8550,
    n8551, n8552, n8553, n8554, n8555, n8556,
    n8557, n8558, n8559, n8560, n8561, n8562,
    n8563, n8564, n8565, n8566, n8567, n8568,
    n8569, n8570, n8571, n8572, n8573, n8574,
    n8575, n8576, n8577, n8578, n8579, n8580,
    n8581, n8582, n8583, n8584, n8585, n8586,
    n8587, n8588, n8589, n8590, n8591, n8592,
    n8593, n8594, n8595, n8596, n8597, n8598,
    n8599, n8600, n8601, n8602, n8603, n8604,
    n8605, n8606, n8607, n8608, n8609, n8610,
    n8611, n8612, n8613, n8614, n8615, n8616,
    n8617, n8618, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658,
    n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8678, n8679, n8680, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688,
    n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706,
    n8707, n8708, n8709, n8710, n8711, n8712,
    n8713, n8714, n8715, n8716, n8717, n8718,
    n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736,
    n8737, n8738, n8739, n8740, n8741, n8742,
    n8743, n8744, n8745, n8746, n8747, n8748,
    n8749, n8750, n8751, n8752, n8753, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766,
    n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778,
    n8779, n8780, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796,
    n8797, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826,
    n8827, n8828, n8829, n8830, n8831, n8832,
    n8833, n8834, n8835, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844,
    n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856,
    n8857, n8858, n8859, n8860, n8861, n8862,
    n8863, n8864, n8865, n8866, n8867, n8868,
    n8869, n8870, n8871, n8872, n8873, n8874,
    n8875, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886,
    n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898,
    n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8906, n8907, n8908, n8909, n8910,
    n8911, n8912, n8913, n8914, n8915, n8916,
    n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8924, n8925, n8926, n8927, n8928,
    n8929, n8930, n8931, n8932, n8933, n8934,
    n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8942, n8943, n8944, n8945, n8946,
    n8947, n8948, n8949, n8950, n8951, n8952,
    n8953, n8954, n8955, n8956, n8957, n8958,
    n8959, n8960, n8961, n8962, n8963, n8964,
    n8965, n8966, n8967, n8968, n8969, n8970,
    n8971, n8972, n8973, n8974, n8975, n8976,
    n8977, n8978, n8979, n8980, n8981, n8982,
    n8983, n8984, n8985, n8986, n8987, n8988,
    n8989, n8990, n8991, n8992, n8993, n8994,
    n8995, n8996, n8997, n8998, n8999, n9000,
    n9001, n9002, n9003, n9004, n9005, n9006,
    n9007, n9008, n9009, n9010, n9011, n9012,
    n9013, n9014, n9015, n9016, n9017, n9018,
    n9019, n9020, n9021, n9022, n9023, n9024,
    n9025, n9026, n9027, n9028, n9029, n9030,
    n9031, n9032, n9033, n9034, n9035, n9036,
    n9037, n9038, n9039, n9040, n9041, n9042,
    n9043, n9044, n9045, n9046, n9047, n9048,
    n9049, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060,
    n9061, n9062, n9063, n9064, n9065, n9066,
    n9067, n9068, n9069, n9070, n9071, n9072,
    n9073, n9074, n9075, n9076, n9077, n9078,
    n9079, n9080, n9081, n9082, n9083, n9084,
    n9085, n9086, n9087, n9088, n9089, n9090,
    n9091, n9092, n9093, n9094, n9095, n9096,
    n9097, n9098, n9099, n9100, n9101, n9102,
    n9103, n9104, n9105, n9106, n9107, n9108,
    n9109, n9110, n9111, n9112, n9113, n9114,
    n9115, n9116, n9117, n9118, n9119, n9120,
    n9121, n9122, n9123, n9124, n9125, n9126,
    n9127, n9128, n9129, n9130, n9131, n9132,
    n9133, n9134, n9135, n9136, n9137, n9138,
    n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9148, n9149, n9150,
    n9151, n9152, n9153, n9154, n9155, n9156,
    n9157, n9158, n9159, n9160, n9161, n9162,
    n9163, n9164, n9165, n9166, n9167, n9168,
    n9169, n9170, n9171, n9172, n9173, n9174,
    n9175, n9176, n9177, n9178, n9179, n9180,
    n9181, n9182, n9183, n9184, n9185, n9186,
    n9187, n9188, n9189, n9190, n9191, n9192,
    n9193, n9194, n9195, n9196, n9197, n9198,
    n9199, n9200, n9201, n9202, n9203, n9204,
    n9205, n9206, n9207, n9208, n9209, n9210,
    n9211, n9212, n9213, n9214, n9215, n9216,
    n9217, n9218, n9219, n9220, n9221, n9222,
    n9223, n9224, n9225, n9226, n9227, n9228,
    n9229, n9230, n9231, n9232, n9233, n9234,
    n9235, n9236, n9237, n9238, n9239, n9240,
    n9241, n9242, n9243, n9244, n9245, n9246,
    n9247, n9248, n9249, n9250, n9251, n9252,
    n9253, n9254, n9255, n9256, n9257, n9258,
    n9259, n9260, n9261, n9262, n9263, n9264,
    n9265, n9266, n9267, n9268, n9269, n9270,
    n9271, n9272, n9273, n9274, n9275, n9276,
    n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9287, n9288,
    n9289, n9290, n9291, n9292, n9293, n9294,
    n9295, n9296, n9297, n9298, n9299, n9300,
    n9301, n9302, n9303, n9304, n9305, n9306,
    n9307, n9308, n9309, n9310, n9311, n9312,
    n9313, n9314, n9315, n9316, n9317, n9318,
    n9319, n9320, n9321, n9322, n9323, n9324,
    n9325, n9326, n9327, n9328, n9329, n9330,
    n9331, n9332, n9333, n9334, n9335, n9336,
    n9337, n9338, n9339, n9340, n9341, n9342,
    n9343, n9344, n9345, n9346, n9347, n9348,
    n9349, n9350, n9351, n9352, n9353, n9354,
    n9355, n9356, n9357, n9358, n9359, n9360,
    n9361, n9362, n9363, n9364, n9365, n9366,
    n9367, n9368, n9369, n9370, n9371, n9372,
    n9373, n9374, n9375, n9376, n9377, n9378,
    n9379, n9380, n9381, n9382, n9383, n9384,
    n9385, n9386, n9387, n9388, n9389, n9390,
    n9391, n9392, n9393, n9394, n9395, n9396,
    n9397, n9398, n9399, n9400, n9401, n9402,
    n9403, n9404, n9405, n9406, n9407, n9408,
    n9409, n9410, n9411, n9412, n9413, n9414,
    n9415, n9416, n9417, n9418, n9419, n9420,
    n9421, n9422, n9423, n9424, n9425, n9426,
    n9427, n9428, n9429, n9430, n9431, n9432,
    n9433, n9434, n9435, n9436, n9437, n9438,
    n9439, n9440, n9441, n9442, n9443, n9444,
    n9445, n9446, n9447, n9448, n9449, n9450,
    n9451, n9452, n9453, n9454, n9455, n9456,
    n9457, n9458, n9459, n9460, n9461, n9462,
    n9463, n9464, n9465, n9466, n9467, n9468,
    n9469, n9470, n9471, n9472, n9473, n9474,
    n9475, n9476, n9477, n9478, n9479, n9480,
    n9481, n9482, n9483, n9484, n9485, n9486,
    n9487, n9488, n9489, n9490, n9491, n9492,
    n9493, n9494, n9495, n9496, n9497, n9498,
    n9499, n9500, n9501, n9502, n9503, n9504,
    n9505, n9506, n9507, n9508, n9509, n9510,
    n9511, n9512, n9513, n9514, n9515, n9516,
    n9517, n9518, n9519, n9520, n9521, n9522,
    n9523, n9524, n9525, n9526, n9527, n9528,
    n9529, n9530, n9531, n9532, n9533, n9534,
    n9535, n9536, n9537, n9538, n9539, n9540,
    n9541, n9542, n9543, n9544, n9545, n9546,
    n9547, n9548, n9549, n9550, n9551, n9552,
    n9553, n9554, n9555, n9556, n9557, n9558,
    n9559, n9560, n9561, n9562, n9563, n9564,
    n9565, n9566, n9567, n9568, n9569, n9570,
    n9571, n9572, n9573, n9574, n9575, n9576,
    n9577, n9578, n9579, n9580, n9581, n9582,
    n9583, n9584, n9585, n9586, n9587, n9588,
    n9589, n9590, n9591, n9592, n9593, n9594,
    n9595, n9596, n9597, n9598, n9599, n9600,
    n9601, n9602, n9603, n9604, n9605, n9606,
    n9607, n9608, n9609, n9610, n9611, n9612,
    n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624,
    n9625, n9626, n9627, n9628, n9629, n9630,
    n9631, n9632, n9633, n9634, n9635, n9636,
    n9637, n9638, n9639, n9640, n9641, n9642,
    n9643, n9644, n9645, n9646, n9647, n9648,
    n9649, n9650, n9651, n9652, n9653, n9654,
    n9655, n9656, n9657, n9658, n9659, n9660,
    n9661, n9662, n9663, n9664, n9665, n9666,
    n9667, n9668, n9669, n9670, n9671, n9672,
    n9673, n9674, n9675, n9676, n9677, n9678,
    n9679, n9680, n9681, n9682, n9683, n9684,
    n9685, n9686, n9687, n9688, n9689, n9690,
    n9691, n9692, n9693, n9694, n9695, n9696,
    n9697, n9698, n9699, n9700, n9701, n9702,
    n9703, n9704, n9705, n9706, n9707, n9708,
    n9709, n9710, n9711, n9712, n9713, n9714,
    n9715, n9716, n9717, n9718, n9719, n9720,
    n9721, n9722, n9723, n9724, n9725, n9726,
    n9727, n9728, n9729, n9730, n9731, n9732,
    n9733, n9734, n9735, n9736, n9737, n9738,
    n9739, n9740, n9741, n9742, n9743, n9744,
    n9745, n9746, n9747, n9748, n9749, n9750,
    n9751, n9752, n9753, n9754, n9755, n9756,
    n9757, n9758, n9759, n9760, n9761, n9762,
    n9763, n9764, n9765, n9766, n9767, n9768,
    n9769, n9770, n9771, n9772, n9773, n9774,
    n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786,
    n9787, n9788, n9789, n9790, n9791, n9792,
    n9793, n9794, n9795, n9796, n9797, n9798,
    n9799, n9800, n9801, n9802, n9803, n9804,
    n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9813, n9814, n9815, n9816,
    n9817, n9818, n9819, n9820, n9821, n9822,
    n9823, n9824, n9825, n9826, n9827, n9828,
    n9829, n9830, n9831, n9832, n9833, n9834,
    n9835, n9836, n9837, n9838, n9839, n9840,
    n9841, n9842, n9843, n9844, n9845, n9846,
    n9847, n9848, n9849, n9850, n9851, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858,
    n9859, n9860, n9861, n9862, n9863, n9864,
    n9865, n9866, n9867, n9868, n9869, n9870,
    n9871, n9872, n9873, n9874, n9875, n9876,
    n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888,
    n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900,
    n9901, n9902, n9903, n9904, n9905, n9906,
    n9907, n9908, n9909, n9910, n9911, n9912,
    n9913, n9914, n9915, n9916, n9917, n9918,
    n9919, n9920, n9921, n9922, n9923, n9924,
    n9925, n9926, n9927, n9928, n9929, n9930,
    n9931, n9932, n9933, n9934, n9935, n9936,
    n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948,
    n9949, n9950, n9951, n9952, n9953, n9954,
    n9955, n9956, n9957, n9958, n9959, n9960,
    n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990,
    n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044,
    n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074,
    n10075, n10076, n10077, n10078, n10079, n10080,
    n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098,
    n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116,
    n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134,
    n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152,
    n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200,
    n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218,
    n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236,
    n10237, n10238, n10239, n10240, n10241, n10242,
    n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254,
    n10255, n10256, n10257, n10258, n10259, n10260,
    n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272,
    n10273, n10274, n10275, n10276, n10277, n10278,
    n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290,
    n10291, n10292, n10293, n10294, n10295, n10296,
    n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10305, n10306, n10307, n10308,
    n10309, n10310, n10311, n10312, n10313, n10314,
    n10315, n10316, n10317, n10318, n10319, n10320,
    n10321, n10322, n10323, n10324, n10325, n10326,
    n10327, n10328, n10329, n10330, n10331, n10332,
    n10333, n10334, n10335, n10336, n10337, n10338,
    n10339, n10340, n10341, n10342, n10343, n10344,
    n10345, n10346, n10347, n10348, n10349, n10350,
    n10351, n10352, n10353, n10354, n10355, n10356,
    n10357, n10358, n10359, n10360, n10361, n10362,
    n10363, n10364, n10365, n10366, n10367, n10368,
    n10369, n10370, n10371, n10372, n10373, n10374,
    n10375, n10376, n10377, n10378, n10379, n10380,
    n10381, n10382, n10383, n10384, n10385, n10386,
    n10387, n10388, n10389, n10390, n10391, n10392,
    n10393, n10394, n10395, n10396, n10397, n10398,
    n10399, n10400, n10401, n10402, n10403, n10404,
    n10405, n10406, n10407, n10408, n10409, n10410,
    n10411, n10412, n10413, n10414, n10415, n10416,
    n10417, n10418, n10419, n10420, n10421, n10422,
    n10423, n10424, n10425, n10426, n10427, n10428,
    n10429, n10430, n10431, n10432, n10433, n10434,
    n10435, n10436, n10437, n10438, n10439, n10440,
    n10441, n10442, n10443, n10444, n10445, n10446,
    n10447, n10448, n10449, n10450, n10451, n10452,
    n10453, n10454, n10455, n10456, n10457, n10458,
    n10459, n10460, n10461, n10462, n10463, n10464,
    n10465, n10466, n10467, n10468, n10469, n10470,
    n10471, n10472, n10473, n10474, n10475, n10476,
    n10477, n10478, n10479, n10480, n10481, n10482,
    n10483, n10484, n10485, n10486, n10487, n10488,
    n10489, n10490, n10491, n10492, n10493, n10494,
    n10495, n10496, n10497, n10498, n10499, n10500,
    n10501, n10502, n10503, n10504, n10505, n10506,
    n10507, n10508, n10509, n10510, n10511, n10512,
    n10513, n10514, n10515, n10516, n10517, n10518,
    n10519, n10520, n10521, n10522, n10523, n10524,
    n10525, n10526, n10527, n10528, n10529, n10530,
    n10531, n10532, n10533, n10534, n10535, n10536,
    n10537, n10538, n10539, n10540, n10541, n10542,
    n10543, n10544, n10545, n10546, n10547, n10548,
    n10549, n10550, n10551, n10552, n10553, n10554,
    n10555, n10556, n10557, n10558, n10559, n10560,
    n10561, n10562, n10563, n10564, n10565, n10566,
    n10567, n10568, n10569, n10570, n10571, n10572,
    n10573, n10574, n10575, n10576, n10577, n10578,
    n10579, n10580, n10581, n10582, n10583, n10584,
    n10585, n10586, n10587, n10588, n10589, n10590,
    n10591, n10592, n10593, n10594, n10595, n10596,
    n10597, n10598, n10599, n10600, n10601, n10602,
    n10603, n10604, n10605, n10606, n10607, n10608,
    n10609, n10610, n10611, n10612, n10613, n10614,
    n10615, n10616, n10617, n10618, n10619, n10620,
    n10621, n10622, n10623, n10624, n10625, n10626,
    n10627, n10628, n10629, n10630, n10631, n10632,
    n10633, n10634, n10635, n10636, n10637, n10638,
    n10639, n10640, n10641, n10642, n10643, n10644,
    n10645, n10646, n10647, n10648, n10649, n10650,
    n10651, n10652, n10653, n10654, n10655, n10656,
    n10657, n10658, n10659, n10660, n10661, n10662,
    n10663, n10664, n10665, n10666, n10667, n10668,
    n10669, n10670, n10671, n10672, n10673, n10674,
    n10675, n10676, n10677, n10678, n10679, n10680,
    n10681, n10682, n10683, n10684, n10685, n10686,
    n10687, n10688, n10689, n10690, n10691, n10692,
    n10693, n10694, n10695, n10696, n10697, n10698,
    n10699, n10700, n10701, n10702, n10703, n10704,
    n10705, n10706, n10707, n10708, n10709, n10710,
    n10711, n10712, n10713, n10714, n10715, n10716,
    n10717, n10718, n10719, n10720, n10721, n10722,
    n10723, n10724, n10725, n10726, n10727, n10728,
    n10729, n10730, n10731, n10732, n10733, n10734,
    n10735, n10736, n10737, n10738, n10739, n10740,
    n10741, n10742, n10743, n10744, n10745, n10746,
    n10747, n10748, n10749, n10750, n10751, n10752,
    n10753, n10754, n10755, n10756, n10757, n10758,
    n10759, n10760, n10761, n10762, n10763, n10764,
    n10765, n10766, n10767, n10768, n10769, n10770,
    n10771, n10772, n10773, n10774, n10775, n10776,
    n10777, n10778, n10779, n10780, n10781, n10782,
    n10783, n10784, n10785, n10786, n10787, n10788,
    n10789, n10790, n10791, n10792, n10793, n10794,
    n10795, n10796, n10797, n10798, n10799, n10800,
    n10801, n10802, n10803, n10804, n10805, n10806,
    n10807, n10808, n10809, n10810, n10811, n10812,
    n10813, n10814, n10815, n10816, n10817, n10818,
    n10819, n10820, n10821, n10822, n10823, n10824,
    n10825, n10826, n10827, n10828, n10829, n10830,
    n10831, n10832, n10833, n10834, n10835, n10836,
    n10837, n10838, n10839, n10840, n10841, n10842,
    n10843, n10844, n10845, n10846, n10847, n10848,
    n10849, n10850, n10851, n10852, n10853, n10854,
    n10855, n10856, n10857, n10858, n10859, n10860,
    n10861, n10862, n10863, n10864, n10865, n10866,
    n10867, n10868, n10869, n10870, n10871, n10872,
    n10873, n10874, n10875, n10876, n10877, n10878,
    n10879, n10880, n10881, n10882, n10883, n10884,
    n10885, n10886, n10887, n10888, n10889, n10890,
    n10891, n10892, n10893, n10894, n10895, n10896,
    n10897, n10898, n10899, n10900, n10901, n10902,
    n10903, n10904, n10905, n10906, n10907, n10908,
    n10909, n10910, n10911, n10912, n10913, n10914,
    n10915, n10916, n10917, n10918, n10919, n10920,
    n10921, n10922, n10923, n10924, n10925, n10926,
    n10927, n10928, n10929, n10930, n10931, n10932,
    n10933, n10934, n10935, n10936, n10937, n10938,
    n10939, n10940, n10941, n10942, n10943, n10944,
    n10945, n10946, n10947, n10948, n10949, n10950,
    n10951, n10952, n10953, n10954, n10955, n10956,
    n10957, n10958, n10959, n10960, n10961, n10962,
    n10963, n10964, n10965, n10966, n10967, n10968,
    n10969, n10970, n10971, n10972, n10973, n10974,
    n10975, n10976, n10977, n10978, n10979, n10980,
    n10981, n10982, n10983, n10984, n10985, n10986,
    n10987, n10988, n10989, n10990, n10991, n10992,
    n10993, n10994, n10995, n10996, n10997, n10998,
    n10999, n11000, n11001, n11002, n11003, n11004,
    n11005, n11006, n11007, n11008, n11009, n11010,
    n11011, n11012, n11013, n11014, n11015, n11016,
    n11017, n11018, n11019, n11020, n11021, n11022,
    n11023, n11024, n11025, n11026, n11027, n11028,
    n11029, n11030, n11031, n11032, n11033, n11034,
    n11035, n11036, n11037, n11038, n11039, n11040,
    n11041, n11042, n11043, n11044, n11045, n11046,
    n11047, n11048, n11049, n11050, n11051, n11052,
    n11053, n11054, n11055, n11056, n11057, n11058,
    n11059, n11060, n11061, n11062, n11063, n11064,
    n11065, n11066, n11067, n11068, n11069, n11070,
    n11071, n11072, n11073, n11074, n11075, n11076,
    n11077, n11078, n11079, n11080, n11081, n11082,
    n11083, n11084, n11085, n11086, n11087, n11088,
    n11089, n11090, n11091, n11092, n11093, n11094,
    n11095, n11096, n11097, n11098, n11099, n11100,
    n11101, n11102, n11103, n11104, n11105, n11106,
    n11107, n11108, n11109, n11110, n11111, n11112,
    n11113, n11114, n11115, n11116, n11117, n11118,
    n11119, n11120, n11121, n11122, n11123, n11124,
    n11125, n11126, n11127, n11128, n11129, n11130,
    n11131, n11132, n11133, n11134, n11135, n11136,
    n11137, n11138, n11139, n11140, n11141, n11142,
    n11143, n11144, n11145, n11146, n11147, n11148,
    n11149, n11150, n11151, n11152, n11153, n11154,
    n11155, n11156, n11157, n11158, n11159, n11160,
    n11161, n11162, n11163, n11164, n11165, n11166,
    n11167, n11168, n11169, n11170, n11171, n11172,
    n11173, n11174, n11175, n11176, n11177, n11178,
    n11179, n11180;
  assign n1003 = pi967  & ~pi968 ;
  assign n1004 = ~pi967  & pi968 ;
  assign n1005 = pi969  & ~n1003;
  assign n1006 = ~n1004 & n1005;
  assign n1007 = ~n1003 & ~n1004;
  assign n1008 = ~pi969  & ~n1007;
  assign n1009 = ~n1006 & ~n1008;
  assign n1010 = pi970  & ~pi971 ;
  assign n1011 = ~pi970  & pi971 ;
  assign n1012 = pi972  & ~n1010;
  assign n1013 = ~n1011 & n1012;
  assign n1014 = ~n1010 & ~n1011;
  assign n1015 = ~pi972  & ~n1014;
  assign n1016 = ~n1013 & ~n1015;
  assign n1017 = ~n1009 & n1016;
  assign n1018 = n1009 & ~n1016;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = pi973  & ~pi974 ;
  assign n1021 = ~pi973  & pi974 ;
  assign n1022 = pi975  & ~n1020;
  assign n1023 = ~n1021 & n1022;
  assign n1024 = ~n1020 & ~n1021;
  assign n1025 = ~pi975  & ~n1024;
  assign n1026 = ~n1023 & ~n1025;
  assign n1027 = pi976  & ~pi977 ;
  assign n1028 = ~pi976  & pi977 ;
  assign n1029 = pi978  & ~n1027;
  assign n1030 = ~n1028 & n1029;
  assign n1031 = ~n1027 & ~n1028;
  assign n1032 = ~pi978  & ~n1031;
  assign n1033 = ~n1030 & ~n1032;
  assign n1034 = ~n1026 & n1033;
  assign n1035 = n1026 & ~n1033;
  assign n1036 = ~n1034 & ~n1035;
  assign n1037 = ~n1019 & ~n1036;
  assign n1038 = pi976  & pi977 ;
  assign n1039 = pi978  & ~n1031;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = pi973  & pi974 ;
  assign n1042 = pi975  & ~n1024;
  assign n1043 = ~n1041 & ~n1042;
  assign n1044 = ~n1040 & ~n1043;
  assign n1045 = ~n1036 & n1044;
  assign n1046 = ~n1026 & ~n1033;
  assign n1047 = n1040 & n1043;
  assign n1048 = ~n1044 & ~n1047;
  assign n1049 = n1046 & n1048;
  assign n1050 = ~n1046 & ~n1048;
  assign n1051 = ~n1045 & ~n1049;
  assign n1052 = ~n1050 & n1051;
  assign n1053 = n1037 & n1052;
  assign n1054 = ~n1037 & ~n1052;
  assign n1055 = ~n1009 & ~n1016;
  assign n1056 = pi970  & pi971 ;
  assign n1057 = pi972  & ~n1014;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = pi967  & pi968 ;
  assign n1060 = pi969  & ~n1007;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = n1058 & ~n1061;
  assign n1063 = ~n1058 & n1061;
  assign n1064 = ~n1062 & ~n1063;
  assign n1065 = n1055 & n1064;
  assign n1066 = ~n1055 & ~n1064;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = ~n1054 & ~n1067;
  assign n1069 = ~n1053 & ~n1068;
  assign n1070 = n1046 & ~n1047;
  assign n1071 = ~n1044 & ~n1070;
  assign n1072 = ~n1069 & ~n1071;
  assign n1073 = n1069 & n1071;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = n1055 & ~n1058;
  assign n1076 = n1061 & ~n1075;
  assign n1077 = ~n1055 & n1058;
  assign n1078 = ~n1076 & ~n1077;
  assign n1079 = ~n1074 & n1078;
  assign n1080 = n1074 & ~n1078;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = pi985  & ~pi986 ;
  assign n1083 = ~pi985  & pi986 ;
  assign n1084 = pi987  & ~n1082;
  assign n1085 = ~n1083 & n1084;
  assign n1086 = ~n1082 & ~n1083;
  assign n1087 = ~pi987  & ~n1086;
  assign n1088 = ~n1085 & ~n1087;
  assign n1089 = pi988  & ~pi989 ;
  assign n1090 = ~pi988  & pi989 ;
  assign n1091 = pi990  & ~n1089;
  assign n1092 = ~n1090 & n1091;
  assign n1093 = ~n1089 & ~n1090;
  assign n1094 = ~pi990  & ~n1093;
  assign n1095 = ~n1092 & ~n1094;
  assign n1096 = ~n1088 & n1095;
  assign n1097 = n1088 & ~n1095;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = pi988  & pi989 ;
  assign n1100 = pi990  & ~n1093;
  assign n1101 = ~n1099 & ~n1100;
  assign n1102 = pi985  & pi986 ;
  assign n1103 = pi987  & ~n1086;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~n1101 & ~n1104;
  assign n1106 = ~n1098 & n1105;
  assign n1107 = ~n1088 & ~n1095;
  assign n1108 = n1101 & n1104;
  assign n1109 = ~n1105 & ~n1108;
  assign n1110 = n1107 & n1109;
  assign n1111 = ~n1107 & ~n1109;
  assign n1112 = ~n1106 & ~n1110;
  assign n1113 = ~n1111 & n1112;
  assign n1114 = pi979  & ~pi980 ;
  assign n1115 = ~pi979  & pi980 ;
  assign n1116 = pi981  & ~n1114;
  assign n1117 = ~n1115 & n1116;
  assign n1118 = ~n1114 & ~n1115;
  assign n1119 = ~pi981  & ~n1118;
  assign n1120 = ~n1117 & ~n1119;
  assign n1121 = pi982  & ~pi983 ;
  assign n1122 = ~pi982  & pi983 ;
  assign n1123 = pi984  & ~n1121;
  assign n1124 = ~n1122 & n1123;
  assign n1125 = ~n1121 & ~n1122;
  assign n1126 = ~pi984  & ~n1125;
  assign n1127 = ~n1124 & ~n1126;
  assign n1128 = ~n1120 & n1127;
  assign n1129 = n1120 & ~n1127;
  assign n1130 = ~n1128 & ~n1129;
  assign n1131 = ~n1098 & ~n1130;
  assign n1132 = ~n1120 & ~n1127;
  assign n1133 = pi982  & pi983 ;
  assign n1134 = pi984  & ~n1125;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = pi979  & pi980 ;
  assign n1137 = pi981  & ~n1118;
  assign n1138 = ~n1136 & ~n1137;
  assign n1139 = n1135 & ~n1138;
  assign n1140 = ~n1135 & n1138;
  assign n1141 = ~n1139 & ~n1140;
  assign n1142 = n1132 & n1141;
  assign n1143 = ~n1132 & ~n1141;
  assign n1144 = ~n1142 & ~n1143;
  assign n1145 = ~n1131 & n1144;
  assign n1146 = n1113 & ~n1145;
  assign n1147 = n1131 & ~n1144;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = n1107 & ~n1108;
  assign n1150 = ~n1105 & ~n1149;
  assign n1151 = ~n1148 & ~n1150;
  assign n1152 = n1148 & n1150;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = n1132 & ~n1135;
  assign n1155 = n1138 & ~n1154;
  assign n1156 = ~n1132 & n1135;
  assign n1157 = ~n1155 & ~n1156;
  assign n1158 = ~n1153 & n1157;
  assign n1159 = n1153 & ~n1157;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = ~n1081 & ~n1160;
  assign n1162 = n1081 & n1160;
  assign n1163 = n1098 & n1130;
  assign n1164 = ~n1131 & ~n1163;
  assign n1165 = n1019 & n1036;
  assign n1166 = ~n1037 & ~n1165;
  assign n1167 = n1164 & n1166;
  assign n1168 = n1131 & ~n1141;
  assign n1169 = ~n1145 & ~n1168;
  assign n1170 = n1113 & ~n1169;
  assign n1171 = ~n1113 & n1169;
  assign n1172 = ~n1170 & ~n1171;
  assign n1173 = n1167 & ~n1172;
  assign n1174 = ~n1167 & n1172;
  assign n1175 = ~n1053 & ~n1054;
  assign n1176 = ~n1067 & n1175;
  assign n1177 = n1067 & ~n1175;
  assign n1178 = ~n1176 & ~n1177;
  assign n1179 = ~n1174 & n1178;
  assign n1180 = ~n1173 & ~n1179;
  assign n1181 = ~n1162 & ~n1180;
  assign n1182 = ~n1161 & ~n1181;
  assign n1183 = ~n1152 & n1157;
  assign n1184 = ~n1151 & ~n1183;
  assign n1185 = ~n1182 & ~n1184;
  assign n1186 = n1182 & n1184;
  assign n1187 = ~n1073 & n1078;
  assign n1188 = ~n1072 & ~n1187;
  assign n1189 = ~n1186 & ~n1188;
  assign n1190 = ~n1185 & ~n1189;
  assign n1191 = ~n1185 & ~n1186;
  assign n1192 = n1188 & ~n1191;
  assign n1193 = ~n1185 & n1189;
  assign n1194 = ~n1192 & ~n1193;
  assign n1195 = ~pi949  & pi950 ;
  assign n1196 = pi949  & ~pi950 ;
  assign n1197 = pi951  & ~n1195;
  assign n1198 = ~n1196 & n1197;
  assign n1199 = ~n1195 & ~n1196;
  assign n1200 = ~pi951  & ~n1199;
  assign n1201 = ~n1198 & ~n1200;
  assign n1202 = ~pi952  & pi953 ;
  assign n1203 = pi952  & ~pi953 ;
  assign n1204 = pi954  & ~n1202;
  assign n1205 = ~n1203 & n1204;
  assign n1206 = ~n1202 & ~n1203;
  assign n1207 = ~pi954  & ~n1206;
  assign n1208 = ~n1205 & ~n1207;
  assign n1209 = ~n1201 & n1208;
  assign n1210 = n1201 & ~n1208;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = ~pi943  & pi944 ;
  assign n1213 = pi943  & ~pi944 ;
  assign n1214 = pi945  & ~n1212;
  assign n1215 = ~n1213 & n1214;
  assign n1216 = ~n1212 & ~n1213;
  assign n1217 = ~pi945  & ~n1216;
  assign n1218 = ~n1215 & ~n1217;
  assign n1219 = ~pi946  & pi947 ;
  assign n1220 = pi946  & ~pi947 ;
  assign n1221 = pi948  & ~n1219;
  assign n1222 = ~n1220 & n1221;
  assign n1223 = ~n1219 & ~n1220;
  assign n1224 = ~pi948  & ~n1223;
  assign n1225 = ~n1222 & ~n1224;
  assign n1226 = ~n1218 & n1225;
  assign n1227 = n1218 & ~n1225;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = ~n1211 & ~n1228;
  assign n1230 = pi952  & pi953 ;
  assign n1231 = pi954  & ~n1206;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = pi949  & pi950 ;
  assign n1234 = pi951  & ~n1199;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = ~n1232 & ~n1235;
  assign n1237 = ~n1211 & n1236;
  assign n1238 = ~n1201 & ~n1208;
  assign n1239 = n1232 & n1235;
  assign n1240 = ~n1236 & ~n1239;
  assign n1241 = n1238 & n1240;
  assign n1242 = ~n1238 & ~n1240;
  assign n1243 = ~n1237 & ~n1241;
  assign n1244 = ~n1242 & n1243;
  assign n1245 = n1229 & n1244;
  assign n1246 = ~n1229 & ~n1244;
  assign n1247 = pi946  & pi947 ;
  assign n1248 = pi948  & ~n1223;
  assign n1249 = ~n1247 & ~n1248;
  assign n1250 = pi943  & pi944 ;
  assign n1251 = pi945  & ~n1216;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = ~n1249 & n1252;
  assign n1254 = n1249 & ~n1252;
  assign n1255 = ~n1253 & ~n1254;
  assign n1256 = ~n1218 & ~n1225;
  assign n1257 = n1255 & n1256;
  assign n1258 = ~n1255 & ~n1256;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = ~n1246 & ~n1259;
  assign n1261 = ~n1245 & ~n1260;
  assign n1262 = n1238 & ~n1239;
  assign n1263 = ~n1236 & ~n1262;
  assign n1264 = ~n1261 & ~n1263;
  assign n1265 = n1261 & n1263;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = ~n1249 & n1256;
  assign n1268 = n1252 & ~n1267;
  assign n1269 = n1249 & ~n1256;
  assign n1270 = ~n1268 & ~n1269;
  assign n1271 = ~n1266 & n1270;
  assign n1272 = n1266 & ~n1270;
  assign n1273 = ~n1271 & ~n1272;
  assign n1274 = ~pi961  & pi962 ;
  assign n1275 = pi961  & ~pi962 ;
  assign n1276 = pi963  & ~n1274;
  assign n1277 = ~n1275 & n1276;
  assign n1278 = ~n1274 & ~n1275;
  assign n1279 = ~pi963  & ~n1278;
  assign n1280 = ~n1277 & ~n1279;
  assign n1281 = ~pi964  & pi965 ;
  assign n1282 = pi964  & ~pi965 ;
  assign n1283 = pi966  & ~n1281;
  assign n1284 = ~n1282 & n1283;
  assign n1285 = ~n1281 & ~n1282;
  assign n1286 = ~pi966  & ~n1285;
  assign n1287 = ~n1284 & ~n1286;
  assign n1288 = ~n1280 & n1287;
  assign n1289 = n1280 & ~n1287;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = ~pi955  & pi956 ;
  assign n1292 = pi955  & ~pi956 ;
  assign n1293 = pi957  & ~n1291;
  assign n1294 = ~n1292 & n1293;
  assign n1295 = ~n1291 & ~n1292;
  assign n1296 = ~pi957  & ~n1295;
  assign n1297 = ~n1294 & ~n1296;
  assign n1298 = ~pi958  & pi959 ;
  assign n1299 = pi958  & ~pi959 ;
  assign n1300 = pi960  & ~n1298;
  assign n1301 = ~n1299 & n1300;
  assign n1302 = ~n1298 & ~n1299;
  assign n1303 = ~pi960  & ~n1302;
  assign n1304 = ~n1301 & ~n1303;
  assign n1305 = ~n1297 & n1304;
  assign n1306 = n1297 & ~n1304;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1290 & ~n1307;
  assign n1309 = pi964  & pi965 ;
  assign n1310 = pi966  & ~n1285;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = pi961  & pi962 ;
  assign n1313 = pi963  & ~n1278;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = n1311 & ~n1314;
  assign n1316 = ~n1311 & n1314;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = n1308 & ~n1317;
  assign n1319 = ~n1280 & ~n1287;
  assign n1320 = n1317 & n1319;
  assign n1321 = ~n1317 & ~n1319;
  assign n1322 = ~n1308 & ~n1320;
  assign n1323 = ~n1321 & n1322;
  assign n1324 = pi958  & pi959 ;
  assign n1325 = pi960  & ~n1302;
  assign n1326 = ~n1324 & ~n1325;
  assign n1327 = pi955  & pi956 ;
  assign n1328 = pi957  & ~n1295;
  assign n1329 = ~n1327 & ~n1328;
  assign n1330 = ~n1326 & ~n1329;
  assign n1331 = ~n1307 & n1330;
  assign n1332 = ~n1297 & ~n1304;
  assign n1333 = n1326 & n1329;
  assign n1334 = ~n1330 & ~n1333;
  assign n1335 = n1332 & n1334;
  assign n1336 = ~n1332 & ~n1334;
  assign n1337 = ~n1331 & ~n1335;
  assign n1338 = ~n1336 & n1337;
  assign n1339 = ~n1323 & n1338;
  assign n1340 = ~n1318 & ~n1339;
  assign n1341 = ~n1311 & n1319;
  assign n1342 = n1314 & ~n1341;
  assign n1343 = n1311 & ~n1319;
  assign n1344 = ~n1342 & ~n1343;
  assign n1345 = ~n1340 & n1344;
  assign n1346 = n1340 & ~n1344;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = n1332 & ~n1333;
  assign n1349 = ~n1330 & ~n1348;
  assign n1350 = n1347 & ~n1349;
  assign n1351 = ~n1347 & n1349;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = n1273 & ~n1352;
  assign n1354 = ~n1273 & n1352;
  assign n1355 = n1290 & n1307;
  assign n1356 = ~n1308 & ~n1355;
  assign n1357 = n1211 & n1228;
  assign n1358 = ~n1229 & ~n1357;
  assign n1359 = n1356 & n1358;
  assign n1360 = ~n1318 & ~n1323;
  assign n1361 = n1338 & n1360;
  assign n1362 = ~n1338 & ~n1360;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = n1359 & n1363;
  assign n1365 = ~n1359 & ~n1363;
  assign n1366 = ~n1245 & ~n1246;
  assign n1367 = ~n1259 & n1366;
  assign n1368 = n1259 & ~n1366;
  assign n1369 = ~n1367 & ~n1368;
  assign n1370 = ~n1365 & n1369;
  assign n1371 = ~n1364 & ~n1370;
  assign n1372 = ~n1354 & n1371;
  assign n1373 = ~n1353 & ~n1372;
  assign n1374 = ~n1346 & ~n1349;
  assign n1375 = ~n1345 & ~n1374;
  assign n1376 = ~n1373 & n1375;
  assign n1377 = n1373 & ~n1375;
  assign n1378 = ~n1376 & ~n1377;
  assign n1379 = ~n1265 & n1270;
  assign n1380 = ~n1264 & ~n1379;
  assign n1381 = n1378 & n1380;
  assign n1382 = ~n1378 & ~n1380;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = n1194 & ~n1383;
  assign n1385 = ~n1194 & n1383;
  assign n1386 = ~n1353 & ~n1354;
  assign n1387 = ~n1371 & n1386;
  assign n1388 = n1371 & ~n1386;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = ~n1161 & ~n1162;
  assign n1391 = ~n1180 & n1390;
  assign n1392 = n1180 & ~n1390;
  assign n1393 = ~n1391 & ~n1392;
  assign n1394 = ~n1389 & ~n1393;
  assign n1395 = n1389 & n1393;
  assign n1396 = ~n1164 & ~n1166;
  assign n1397 = ~n1167 & ~n1396;
  assign n1398 = ~n1356 & ~n1358;
  assign n1399 = ~n1359 & ~n1398;
  assign n1400 = n1397 & n1399;
  assign n1401 = ~n1173 & ~n1174;
  assign n1402 = ~n1178 & n1401;
  assign n1403 = n1178 & ~n1401;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = n1400 & ~n1404;
  assign n1406 = ~n1400 & n1404;
  assign n1407 = ~n1364 & ~n1365;
  assign n1408 = ~n1369 & n1407;
  assign n1409 = n1369 & ~n1407;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1406 & ~n1410;
  assign n1412 = ~n1405 & ~n1411;
  assign n1413 = ~n1395 & n1412;
  assign n1414 = ~n1394 & ~n1413;
  assign n1415 = ~n1385 & n1414;
  assign n1416 = ~n1384 & ~n1415;
  assign n1417 = n1190 & n1416;
  assign n1418 = ~n1190 & ~n1416;
  assign n1419 = ~n1377 & n1380;
  assign n1420 = ~n1376 & ~n1419;
  assign n1421 = ~n1418 & ~n1420;
  assign n1422 = ~n1417 & ~n1421;
  assign n1423 = pi3  & pi4 ;
  assign n1424 = ~pi3  & pi4 ;
  assign n1425 = pi3  & ~pi4 ;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = pi5  & ~n1426;
  assign n1428 = ~n1423 & ~n1427;
  assign n1429 = pi0  & pi1 ;
  assign n1430 = ~pi0  & pi1 ;
  assign n1431 = pi0  & ~pi1 ;
  assign n1432 = ~n1430 & ~n1431;
  assign n1433 = pi2  & ~n1432;
  assign n1434 = ~n1429 & ~n1433;
  assign n1435 = ~n1428 & n1434;
  assign n1436 = n1428 & ~n1434;
  assign n1437 = ~n1435 & ~n1436;
  assign n1438 = pi5  & ~n1424;
  assign n1439 = ~n1425 & n1438;
  assign n1440 = ~pi5  & ~n1426;
  assign n1441 = ~n1439 & ~n1440;
  assign n1442 = ~pi2  & ~n1432;
  assign n1443 = pi2  & ~n1430;
  assign n1444 = ~n1431 & n1443;
  assign n1445 = ~n1442 & ~n1444;
  assign n1446 = ~pi6  & ~n1445;
  assign n1447 = pi6  & n1445;
  assign n1448 = ~n1446 & ~n1447;
  assign n1449 = ~n1441 & ~n1448;
  assign n1450 = pi6  & ~n1445;
  assign n1451 = ~n1449 & ~n1450;
  assign n1452 = ~n1437 & ~n1451;
  assign n1453 = ~n1428 & ~n1434;
  assign n1454 = ~n1452 & ~n1453;
  assign n1455 = ~pi997  & pi998 ;
  assign n1456 = pi997  & ~pi998 ;
  assign n1457 = pi999  & ~n1455;
  assign n1458 = ~n1456 & n1457;
  assign n1459 = ~n1455 & ~n1456;
  assign n1460 = ~pi999  & ~n1459;
  assign n1461 = ~n1458 & ~n1460;
  assign n1462 = n1441 & ~n1448;
  assign n1463 = ~n1441 & n1448;
  assign n1464 = ~n1462 & ~n1463;
  assign n1465 = ~n1461 & ~n1464;
  assign n1466 = n1437 & n1451;
  assign n1467 = ~n1452 & ~n1466;
  assign n1468 = n1465 & n1467;
  assign n1469 = pi997  & pi998 ;
  assign n1470 = pi999  & ~n1459;
  assign n1471 = ~n1469 & ~n1470;
  assign n1472 = ~n1465 & ~n1467;
  assign n1473 = ~n1471 & ~n1472;
  assign n1474 = ~n1468 & ~n1473;
  assign n1475 = ~n1454 & ~n1474;
  assign n1476 = n1454 & n1474;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = ~pi991  & pi992 ;
  assign n1479 = pi991  & ~pi992 ;
  assign n1480 = pi993  & ~n1478;
  assign n1481 = ~n1479 & n1480;
  assign n1482 = ~n1478 & ~n1479;
  assign n1483 = ~pi993  & ~n1482;
  assign n1484 = ~n1481 & ~n1483;
  assign n1485 = ~pi994  & pi995 ;
  assign n1486 = pi994  & ~pi995 ;
  assign n1487 = pi996  & ~n1485;
  assign n1488 = ~n1486 & n1487;
  assign n1489 = ~n1485 & ~n1486;
  assign n1490 = ~pi996  & ~n1489;
  assign n1491 = ~n1488 & ~n1490;
  assign n1492 = ~n1484 & n1491;
  assign n1493 = n1484 & ~n1491;
  assign n1494 = ~n1492 & ~n1493;
  assign n1495 = n1461 & n1464;
  assign n1496 = ~n1465 & ~n1495;
  assign n1497 = ~n1494 & n1496;
  assign n1498 = ~n1468 & ~n1472;
  assign n1499 = n1471 & ~n1498;
  assign n1500 = ~n1471 & n1498;
  assign n1501 = ~n1499 & ~n1500;
  assign n1502 = ~n1497 & ~n1501;
  assign n1503 = n1497 & n1501;
  assign n1504 = pi994  & pi995 ;
  assign n1505 = pi996  & ~n1489;
  assign n1506 = ~n1504 & ~n1505;
  assign n1507 = pi991  & pi992 ;
  assign n1508 = pi993  & ~n1482;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = ~n1506 & ~n1509;
  assign n1511 = ~n1494 & n1510;
  assign n1512 = ~n1484 & ~n1491;
  assign n1513 = n1506 & n1509;
  assign n1514 = ~n1510 & ~n1513;
  assign n1515 = n1512 & n1514;
  assign n1516 = ~n1512 & ~n1514;
  assign n1517 = ~n1511 & ~n1515;
  assign n1518 = ~n1516 & n1517;
  assign n1519 = ~n1503 & ~n1518;
  assign n1520 = ~n1502 & ~n1519;
  assign n1521 = ~n1477 & ~n1520;
  assign n1522 = n1512 & ~n1513;
  assign n1523 = ~n1510 & ~n1522;
  assign n1524 = ~n1521 & ~n1523;
  assign n1525 = n1475 & n1524;
  assign n1526 = pi7  & ~pi8 ;
  assign n1527 = ~pi7  & pi8 ;
  assign n1528 = pi9  & ~n1526;
  assign n1529 = ~n1527 & n1528;
  assign n1530 = ~n1526 & ~n1527;
  assign n1531 = ~pi9  & ~n1530;
  assign n1532 = ~n1529 & ~n1531;
  assign n1533 = pi10  & ~pi11 ;
  assign n1534 = ~pi10  & pi11 ;
  assign n1535 = pi12  & ~n1533;
  assign n1536 = ~n1534 & n1535;
  assign n1537 = ~n1533 & ~n1534;
  assign n1538 = ~pi12  & ~n1537;
  assign n1539 = ~n1536 & ~n1538;
  assign n1540 = ~n1532 & n1539;
  assign n1541 = n1532 & ~n1539;
  assign n1542 = ~n1540 & ~n1541;
  assign n1543 = pi13  & ~pi14 ;
  assign n1544 = ~pi13  & pi14 ;
  assign n1545 = pi15  & ~n1543;
  assign n1546 = ~n1544 & n1545;
  assign n1547 = ~n1543 & ~n1544;
  assign n1548 = ~pi15  & ~n1547;
  assign n1549 = ~n1546 & ~n1548;
  assign n1550 = pi16  & ~pi17 ;
  assign n1551 = ~pi16  & pi17 ;
  assign n1552 = pi18  & ~n1550;
  assign n1553 = ~n1551 & n1552;
  assign n1554 = ~n1550 & ~n1551;
  assign n1555 = ~pi18  & ~n1554;
  assign n1556 = ~n1553 & ~n1555;
  assign n1557 = ~n1549 & n1556;
  assign n1558 = n1549 & ~n1556;
  assign n1559 = ~n1557 & ~n1558;
  assign n1560 = ~n1542 & ~n1559;
  assign n1561 = pi16  & pi17 ;
  assign n1562 = pi18  & ~n1554;
  assign n1563 = ~n1561 & ~n1562;
  assign n1564 = pi13  & pi14 ;
  assign n1565 = pi15  & ~n1547;
  assign n1566 = ~n1564 & ~n1565;
  assign n1567 = ~n1563 & ~n1566;
  assign n1568 = ~n1559 & n1567;
  assign n1569 = ~n1549 & ~n1556;
  assign n1570 = n1563 & n1566;
  assign n1571 = ~n1567 & ~n1570;
  assign n1572 = n1569 & n1571;
  assign n1573 = ~n1569 & ~n1571;
  assign n1574 = ~n1568 & ~n1572;
  assign n1575 = ~n1573 & n1574;
  assign n1576 = n1560 & n1575;
  assign n1577 = ~n1560 & ~n1575;
  assign n1578 = ~n1532 & ~n1539;
  assign n1579 = pi10  & pi11 ;
  assign n1580 = pi12  & ~n1537;
  assign n1581 = ~n1579 & ~n1580;
  assign n1582 = pi7  & pi8 ;
  assign n1583 = pi9  & ~n1530;
  assign n1584 = ~n1582 & ~n1583;
  assign n1585 = n1581 & ~n1584;
  assign n1586 = ~n1581 & n1584;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = n1578 & n1587;
  assign n1589 = ~n1578 & ~n1587;
  assign n1590 = ~n1588 & ~n1589;
  assign n1591 = ~n1577 & ~n1590;
  assign n1592 = ~n1576 & ~n1591;
  assign n1593 = n1569 & ~n1570;
  assign n1594 = ~n1567 & ~n1593;
  assign n1595 = ~n1592 & ~n1594;
  assign n1596 = n1592 & n1594;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = n1578 & ~n1581;
  assign n1599 = n1584 & ~n1598;
  assign n1600 = ~n1578 & n1581;
  assign n1601 = ~n1599 & ~n1600;
  assign n1602 = ~n1597 & n1601;
  assign n1603 = n1597 & ~n1601;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = pi25  & ~pi26 ;
  assign n1606 = ~pi25  & pi26 ;
  assign n1607 = pi27  & ~n1605;
  assign n1608 = ~n1606 & n1607;
  assign n1609 = ~n1605 & ~n1606;
  assign n1610 = ~pi27  & ~n1609;
  assign n1611 = ~n1608 & ~n1610;
  assign n1612 = pi28  & ~pi29 ;
  assign n1613 = ~pi28  & pi29 ;
  assign n1614 = pi30  & ~n1612;
  assign n1615 = ~n1613 & n1614;
  assign n1616 = ~n1612 & ~n1613;
  assign n1617 = ~pi30  & ~n1616;
  assign n1618 = ~n1615 & ~n1617;
  assign n1619 = ~n1611 & n1618;
  assign n1620 = n1611 & ~n1618;
  assign n1621 = ~n1619 & ~n1620;
  assign n1622 = pi28  & pi29 ;
  assign n1623 = pi30  & ~n1616;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = pi25  & pi26 ;
  assign n1626 = pi27  & ~n1609;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = ~n1624 & ~n1627;
  assign n1629 = ~n1621 & n1628;
  assign n1630 = ~n1611 & ~n1618;
  assign n1631 = n1624 & n1627;
  assign n1632 = ~n1628 & ~n1631;
  assign n1633 = n1630 & n1632;
  assign n1634 = ~n1630 & ~n1632;
  assign n1635 = ~n1629 & ~n1633;
  assign n1636 = ~n1634 & n1635;
  assign n1637 = pi19  & ~pi20 ;
  assign n1638 = ~pi19  & pi20 ;
  assign n1639 = pi21  & ~n1637;
  assign n1640 = ~n1638 & n1639;
  assign n1641 = ~n1637 & ~n1638;
  assign n1642 = ~pi21  & ~n1641;
  assign n1643 = ~n1640 & ~n1642;
  assign n1644 = pi22  & ~pi23 ;
  assign n1645 = ~pi22  & pi23 ;
  assign n1646 = pi24  & ~n1644;
  assign n1647 = ~n1645 & n1646;
  assign n1648 = ~n1644 & ~n1645;
  assign n1649 = ~pi24  & ~n1648;
  assign n1650 = ~n1647 & ~n1649;
  assign n1651 = ~n1643 & n1650;
  assign n1652 = n1643 & ~n1650;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = ~n1621 & ~n1653;
  assign n1655 = ~n1643 & ~n1650;
  assign n1656 = pi22  & pi23 ;
  assign n1657 = pi24  & ~n1648;
  assign n1658 = ~n1656 & ~n1657;
  assign n1659 = pi19  & pi20 ;
  assign n1660 = pi21  & ~n1641;
  assign n1661 = ~n1659 & ~n1660;
  assign n1662 = n1658 & ~n1661;
  assign n1663 = ~n1658 & n1661;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = n1655 & n1664;
  assign n1666 = ~n1655 & ~n1664;
  assign n1667 = ~n1665 & ~n1666;
  assign n1668 = ~n1654 & n1667;
  assign n1669 = n1636 & ~n1668;
  assign n1670 = n1654 & ~n1667;
  assign n1671 = ~n1669 & ~n1670;
  assign n1672 = n1630 & ~n1631;
  assign n1673 = ~n1628 & ~n1672;
  assign n1674 = ~n1671 & ~n1673;
  assign n1675 = n1671 & n1673;
  assign n1676 = ~n1674 & ~n1675;
  assign n1677 = n1655 & ~n1658;
  assign n1678 = n1661 & ~n1677;
  assign n1679 = ~n1655 & n1658;
  assign n1680 = ~n1678 & ~n1679;
  assign n1681 = ~n1676 & n1680;
  assign n1682 = n1676 & ~n1680;
  assign n1683 = ~n1681 & ~n1682;
  assign n1684 = ~n1604 & ~n1683;
  assign n1685 = n1604 & n1683;
  assign n1686 = n1621 & n1653;
  assign n1687 = ~n1654 & ~n1686;
  assign n1688 = n1542 & n1559;
  assign n1689 = ~n1560 & ~n1688;
  assign n1690 = n1687 & n1689;
  assign n1691 = n1654 & ~n1664;
  assign n1692 = ~n1668 & ~n1691;
  assign n1693 = n1636 & ~n1692;
  assign n1694 = ~n1636 & n1692;
  assign n1695 = ~n1693 & ~n1694;
  assign n1696 = n1690 & ~n1695;
  assign n1697 = ~n1690 & n1695;
  assign n1698 = ~n1576 & ~n1577;
  assign n1699 = ~n1590 & n1698;
  assign n1700 = n1590 & ~n1698;
  assign n1701 = ~n1699 & ~n1700;
  assign n1702 = ~n1697 & n1701;
  assign n1703 = ~n1696 & ~n1702;
  assign n1704 = ~n1685 & ~n1703;
  assign n1705 = ~n1684 & ~n1704;
  assign n1706 = ~n1675 & n1680;
  assign n1707 = ~n1674 & ~n1706;
  assign n1708 = ~n1705 & ~n1707;
  assign n1709 = n1705 & n1707;
  assign n1710 = ~n1596 & n1601;
  assign n1711 = ~n1595 & ~n1710;
  assign n1712 = ~n1709 & ~n1711;
  assign n1713 = ~n1708 & ~n1712;
  assign n1714 = n1525 & ~n1713;
  assign n1715 = ~n1525 & n1713;
  assign n1716 = ~n1714 & ~n1715;
  assign n1717 = n1477 & n1520;
  assign n1718 = ~n1475 & ~n1524;
  assign n1719 = ~n1525 & ~n1718;
  assign n1720 = ~n1717 & ~n1719;
  assign n1721 = ~n1708 & ~n1709;
  assign n1722 = n1711 & ~n1721;
  assign n1723 = ~n1708 & n1712;
  assign n1724 = ~n1722 & ~n1723;
  assign n1725 = n1720 & ~n1724;
  assign n1726 = ~n1720 & n1724;
  assign n1727 = n1477 & ~n1520;
  assign n1728 = ~n1477 & n1520;
  assign n1729 = ~n1727 & ~n1728;
  assign n1730 = n1523 & n1729;
  assign n1731 = ~n1523 & ~n1729;
  assign n1732 = ~n1730 & ~n1731;
  assign n1733 = ~n1684 & ~n1685;
  assign n1734 = ~n1703 & n1733;
  assign n1735 = n1703 & ~n1733;
  assign n1736 = ~n1734 & ~n1735;
  assign n1737 = ~n1732 & ~n1736;
  assign n1738 = n1732 & n1736;
  assign n1739 = ~n1494 & ~n1496;
  assign n1740 = n1494 & n1496;
  assign n1741 = ~n1739 & ~n1740;
  assign n1742 = ~n1687 & ~n1689;
  assign n1743 = ~n1690 & ~n1742;
  assign n1744 = ~n1741 & n1743;
  assign n1745 = ~n1696 & ~n1697;
  assign n1746 = ~n1701 & n1745;
  assign n1747 = n1701 & ~n1745;
  assign n1748 = ~n1746 & ~n1747;
  assign n1749 = n1744 & ~n1748;
  assign n1750 = ~n1744 & n1748;
  assign n1751 = ~n1502 & ~n1503;
  assign n1752 = ~n1518 & n1751;
  assign n1753 = n1518 & ~n1751;
  assign n1754 = ~n1752 & ~n1753;
  assign n1755 = ~n1750 & ~n1754;
  assign n1756 = ~n1749 & ~n1755;
  assign n1757 = ~n1738 & n1756;
  assign n1758 = ~n1737 & ~n1757;
  assign n1759 = ~n1726 & ~n1758;
  assign n1760 = ~n1725 & ~n1759;
  assign n1761 = n1716 & n1760;
  assign n1762 = ~n1716 & ~n1760;
  assign n1763 = ~n1761 & ~n1762;
  assign n1764 = ~pi37  & pi38 ;
  assign n1765 = pi37  & ~pi38 ;
  assign n1766 = pi39  & ~n1764;
  assign n1767 = ~n1765 & n1766;
  assign n1768 = ~n1764 & ~n1765;
  assign n1769 = ~pi39  & ~n1768;
  assign n1770 = ~n1767 & ~n1769;
  assign n1771 = ~pi40  & pi41 ;
  assign n1772 = pi40  & ~pi41 ;
  assign n1773 = pi42  & ~n1771;
  assign n1774 = ~n1772 & n1773;
  assign n1775 = ~n1771 & ~n1772;
  assign n1776 = ~pi42  & ~n1775;
  assign n1777 = ~n1774 & ~n1776;
  assign n1778 = ~n1770 & n1777;
  assign n1779 = n1770 & ~n1777;
  assign n1780 = ~n1778 & ~n1779;
  assign n1781 = ~pi31  & pi32 ;
  assign n1782 = pi31  & ~pi32 ;
  assign n1783 = pi33  & ~n1781;
  assign n1784 = ~n1782 & n1783;
  assign n1785 = ~n1781 & ~n1782;
  assign n1786 = ~pi33  & ~n1785;
  assign n1787 = ~n1784 & ~n1786;
  assign n1788 = ~pi34  & pi35 ;
  assign n1789 = pi34  & ~pi35 ;
  assign n1790 = pi36  & ~n1788;
  assign n1791 = ~n1789 & n1790;
  assign n1792 = ~n1788 & ~n1789;
  assign n1793 = ~pi36  & ~n1792;
  assign n1794 = ~n1791 & ~n1793;
  assign n1795 = ~n1787 & n1794;
  assign n1796 = n1787 & ~n1794;
  assign n1797 = ~n1795 & ~n1796;
  assign n1798 = ~n1780 & ~n1797;
  assign n1799 = pi40  & pi41 ;
  assign n1800 = pi42  & ~n1775;
  assign n1801 = ~n1799 & ~n1800;
  assign n1802 = pi37  & pi38 ;
  assign n1803 = pi39  & ~n1768;
  assign n1804 = ~n1802 & ~n1803;
  assign n1805 = ~n1801 & ~n1804;
  assign n1806 = ~n1780 & n1805;
  assign n1807 = ~n1770 & ~n1777;
  assign n1808 = n1801 & n1804;
  assign n1809 = ~n1805 & ~n1808;
  assign n1810 = n1807 & n1809;
  assign n1811 = ~n1807 & ~n1809;
  assign n1812 = ~n1806 & ~n1810;
  assign n1813 = ~n1811 & n1812;
  assign n1814 = n1798 & n1813;
  assign n1815 = ~n1798 & ~n1813;
  assign n1816 = pi34  & pi35 ;
  assign n1817 = pi36  & ~n1792;
  assign n1818 = ~n1816 & ~n1817;
  assign n1819 = pi31  & pi32 ;
  assign n1820 = pi33  & ~n1785;
  assign n1821 = ~n1819 & ~n1820;
  assign n1822 = ~n1818 & n1821;
  assign n1823 = n1818 & ~n1821;
  assign n1824 = ~n1822 & ~n1823;
  assign n1825 = ~n1787 & ~n1794;
  assign n1826 = n1824 & n1825;
  assign n1827 = ~n1824 & ~n1825;
  assign n1828 = ~n1826 & ~n1827;
  assign n1829 = ~n1815 & ~n1828;
  assign n1830 = ~n1814 & ~n1829;
  assign n1831 = n1807 & ~n1808;
  assign n1832 = ~n1805 & ~n1831;
  assign n1833 = ~n1830 & ~n1832;
  assign n1834 = n1830 & n1832;
  assign n1835 = ~n1833 & ~n1834;
  assign n1836 = ~n1818 & n1825;
  assign n1837 = n1821 & ~n1836;
  assign n1838 = n1818 & ~n1825;
  assign n1839 = ~n1837 & ~n1838;
  assign n1840 = ~n1835 & n1839;
  assign n1841 = n1835 & ~n1839;
  assign n1842 = ~n1840 & ~n1841;
  assign n1843 = pi49  & ~pi50 ;
  assign n1844 = ~pi49  & pi50 ;
  assign n1845 = pi51  & ~n1843;
  assign n1846 = ~n1844 & n1845;
  assign n1847 = ~n1843 & ~n1844;
  assign n1848 = ~pi51  & ~n1847;
  assign n1849 = ~n1846 & ~n1848;
  assign n1850 = pi52  & ~pi53 ;
  assign n1851 = ~pi52  & pi53 ;
  assign n1852 = pi54  & ~n1850;
  assign n1853 = ~n1851 & n1852;
  assign n1854 = ~n1850 & ~n1851;
  assign n1855 = ~pi54  & ~n1854;
  assign n1856 = ~n1853 & ~n1855;
  assign n1857 = ~n1849 & n1856;
  assign n1858 = n1849 & ~n1856;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = pi52  & pi53 ;
  assign n1861 = pi54  & ~n1854;
  assign n1862 = ~n1860 & ~n1861;
  assign n1863 = pi49  & pi50 ;
  assign n1864 = pi51  & ~n1847;
  assign n1865 = ~n1863 & ~n1864;
  assign n1866 = ~n1862 & ~n1865;
  assign n1867 = ~n1859 & n1866;
  assign n1868 = ~n1849 & ~n1856;
  assign n1869 = n1862 & n1865;
  assign n1870 = ~n1866 & ~n1869;
  assign n1871 = n1868 & n1870;
  assign n1872 = ~n1868 & ~n1870;
  assign n1873 = ~n1867 & ~n1871;
  assign n1874 = ~n1872 & n1873;
  assign n1875 = pi43  & ~pi44 ;
  assign n1876 = ~pi43  & pi44 ;
  assign n1877 = pi45  & ~n1875;
  assign n1878 = ~n1876 & n1877;
  assign n1879 = ~n1875 & ~n1876;
  assign n1880 = ~pi45  & ~n1879;
  assign n1881 = ~n1878 & ~n1880;
  assign n1882 = pi46  & ~pi47 ;
  assign n1883 = ~pi46  & pi47 ;
  assign n1884 = pi48  & ~n1882;
  assign n1885 = ~n1883 & n1884;
  assign n1886 = ~n1882 & ~n1883;
  assign n1887 = ~pi48  & ~n1886;
  assign n1888 = ~n1885 & ~n1887;
  assign n1889 = ~n1881 & n1888;
  assign n1890 = n1881 & ~n1888;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = ~n1859 & ~n1891;
  assign n1893 = ~n1881 & ~n1888;
  assign n1894 = pi46  & pi47 ;
  assign n1895 = pi48  & ~n1886;
  assign n1896 = ~n1894 & ~n1895;
  assign n1897 = pi43  & pi44 ;
  assign n1898 = pi45  & ~n1879;
  assign n1899 = ~n1897 & ~n1898;
  assign n1900 = n1896 & ~n1899;
  assign n1901 = ~n1896 & n1899;
  assign n1902 = ~n1900 & ~n1901;
  assign n1903 = n1893 & n1902;
  assign n1904 = ~n1893 & ~n1902;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = ~n1892 & n1905;
  assign n1907 = n1874 & ~n1906;
  assign n1908 = n1892 & ~n1905;
  assign n1909 = ~n1907 & ~n1908;
  assign n1910 = n1868 & ~n1869;
  assign n1911 = ~n1866 & ~n1910;
  assign n1912 = ~n1909 & ~n1911;
  assign n1913 = n1909 & n1911;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = n1893 & ~n1896;
  assign n1916 = n1899 & ~n1915;
  assign n1917 = ~n1893 & n1896;
  assign n1918 = ~n1916 & ~n1917;
  assign n1919 = ~n1914 & n1918;
  assign n1920 = n1914 & ~n1918;
  assign n1921 = ~n1919 & ~n1920;
  assign n1922 = ~n1842 & ~n1921;
  assign n1923 = n1842 & n1921;
  assign n1924 = n1859 & n1891;
  assign n1925 = ~n1892 & ~n1924;
  assign n1926 = n1780 & n1797;
  assign n1927 = ~n1798 & ~n1926;
  assign n1928 = n1925 & n1927;
  assign n1929 = n1892 & ~n1902;
  assign n1930 = ~n1906 & ~n1929;
  assign n1931 = n1874 & ~n1930;
  assign n1932 = ~n1874 & n1930;
  assign n1933 = ~n1931 & ~n1932;
  assign n1934 = n1928 & ~n1933;
  assign n1935 = ~n1928 & n1933;
  assign n1936 = ~n1814 & ~n1815;
  assign n1937 = ~n1828 & n1936;
  assign n1938 = n1828 & ~n1936;
  assign n1939 = ~n1937 & ~n1938;
  assign n1940 = ~n1935 & n1939;
  assign n1941 = ~n1934 & ~n1940;
  assign n1942 = ~n1923 & ~n1941;
  assign n1943 = ~n1922 & ~n1942;
  assign n1944 = ~n1913 & n1918;
  assign n1945 = ~n1912 & ~n1944;
  assign n1946 = ~n1943 & ~n1945;
  assign n1947 = n1943 & n1945;
  assign n1948 = ~n1834 & n1839;
  assign n1949 = ~n1833 & ~n1948;
  assign n1950 = ~n1947 & ~n1949;
  assign n1951 = ~n1946 & ~n1950;
  assign n1952 = pi55  & ~pi56 ;
  assign n1953 = ~pi55  & pi56 ;
  assign n1954 = pi57  & ~n1952;
  assign n1955 = ~n1953 & n1954;
  assign n1956 = ~n1952 & ~n1953;
  assign n1957 = ~pi57  & ~n1956;
  assign n1958 = ~n1955 & ~n1957;
  assign n1959 = pi58  & ~pi59 ;
  assign n1960 = ~pi58  & pi59 ;
  assign n1961 = pi60  & ~n1959;
  assign n1962 = ~n1960 & n1961;
  assign n1963 = ~n1959 & ~n1960;
  assign n1964 = ~pi60  & ~n1963;
  assign n1965 = ~n1962 & ~n1964;
  assign n1966 = ~n1958 & n1965;
  assign n1967 = n1958 & ~n1965;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = pi61  & ~pi62 ;
  assign n1970 = ~pi61  & pi62 ;
  assign n1971 = pi63  & ~n1969;
  assign n1972 = ~n1970 & n1971;
  assign n1973 = ~n1969 & ~n1970;
  assign n1974 = ~pi63  & ~n1973;
  assign n1975 = ~n1972 & ~n1974;
  assign n1976 = pi64  & ~pi65 ;
  assign n1977 = ~pi64  & pi65 ;
  assign n1978 = pi66  & ~n1976;
  assign n1979 = ~n1977 & n1978;
  assign n1980 = ~n1976 & ~n1977;
  assign n1981 = ~pi66  & ~n1980;
  assign n1982 = ~n1979 & ~n1981;
  assign n1983 = ~n1975 & n1982;
  assign n1984 = n1975 & ~n1982;
  assign n1985 = ~n1983 & ~n1984;
  assign n1986 = ~n1968 & ~n1985;
  assign n1987 = pi64  & pi65 ;
  assign n1988 = pi66  & ~n1980;
  assign n1989 = ~n1987 & ~n1988;
  assign n1990 = pi61  & pi62 ;
  assign n1991 = pi63  & ~n1973;
  assign n1992 = ~n1990 & ~n1991;
  assign n1993 = ~n1989 & ~n1992;
  assign n1994 = ~n1985 & n1993;
  assign n1995 = ~n1975 & ~n1982;
  assign n1996 = n1989 & n1992;
  assign n1997 = ~n1993 & ~n1996;
  assign n1998 = n1995 & n1997;
  assign n1999 = ~n1995 & ~n1997;
  assign n2000 = ~n1994 & ~n1998;
  assign n2001 = ~n1999 & n2000;
  assign n2002 = n1986 & n2001;
  assign n2003 = ~n1986 & ~n2001;
  assign n2004 = ~n1958 & ~n1965;
  assign n2005 = pi58  & pi59 ;
  assign n2006 = pi60  & ~n1963;
  assign n2007 = ~n2005 & ~n2006;
  assign n2008 = pi55  & pi56 ;
  assign n2009 = pi57  & ~n1956;
  assign n2010 = ~n2008 & ~n2009;
  assign n2011 = n2007 & ~n2010;
  assign n2012 = ~n2007 & n2010;
  assign n2013 = ~n2011 & ~n2012;
  assign n2014 = n2004 & n2013;
  assign n2015 = ~n2004 & ~n2013;
  assign n2016 = ~n2014 & ~n2015;
  assign n2017 = ~n2003 & ~n2016;
  assign n2018 = ~n2002 & ~n2017;
  assign n2019 = n1995 & ~n1996;
  assign n2020 = ~n1993 & ~n2019;
  assign n2021 = ~n2018 & ~n2020;
  assign n2022 = n2018 & n2020;
  assign n2023 = ~n2021 & ~n2022;
  assign n2024 = n2004 & ~n2007;
  assign n2025 = n2010 & ~n2024;
  assign n2026 = ~n2004 & n2007;
  assign n2027 = ~n2025 & ~n2026;
  assign n2028 = ~n2023 & n2027;
  assign n2029 = n2023 & ~n2027;
  assign n2030 = ~n2028 & ~n2029;
  assign n2031 = pi73  & ~pi74 ;
  assign n2032 = ~pi73  & pi74 ;
  assign n2033 = pi75  & ~n2031;
  assign n2034 = ~n2032 & n2033;
  assign n2035 = ~n2031 & ~n2032;
  assign n2036 = ~pi75  & ~n2035;
  assign n2037 = ~n2034 & ~n2036;
  assign n2038 = pi76  & ~pi77 ;
  assign n2039 = ~pi76  & pi77 ;
  assign n2040 = pi78  & ~n2038;
  assign n2041 = ~n2039 & n2040;
  assign n2042 = ~n2038 & ~n2039;
  assign n2043 = ~pi78  & ~n2042;
  assign n2044 = ~n2041 & ~n2043;
  assign n2045 = ~n2037 & n2044;
  assign n2046 = n2037 & ~n2044;
  assign n2047 = ~n2045 & ~n2046;
  assign n2048 = pi76  & pi77 ;
  assign n2049 = pi78  & ~n2042;
  assign n2050 = ~n2048 & ~n2049;
  assign n2051 = pi73  & pi74 ;
  assign n2052 = pi75  & ~n2035;
  assign n2053 = ~n2051 & ~n2052;
  assign n2054 = ~n2050 & ~n2053;
  assign n2055 = ~n2047 & n2054;
  assign n2056 = ~n2037 & ~n2044;
  assign n2057 = n2050 & n2053;
  assign n2058 = ~n2054 & ~n2057;
  assign n2059 = n2056 & n2058;
  assign n2060 = ~n2056 & ~n2058;
  assign n2061 = ~n2055 & ~n2059;
  assign n2062 = ~n2060 & n2061;
  assign n2063 = pi67  & ~pi68 ;
  assign n2064 = ~pi67  & pi68 ;
  assign n2065 = pi69  & ~n2063;
  assign n2066 = ~n2064 & n2065;
  assign n2067 = ~n2063 & ~n2064;
  assign n2068 = ~pi69  & ~n2067;
  assign n2069 = ~n2066 & ~n2068;
  assign n2070 = pi70  & ~pi71 ;
  assign n2071 = ~pi70  & pi71 ;
  assign n2072 = pi72  & ~n2070;
  assign n2073 = ~n2071 & n2072;
  assign n2074 = ~n2070 & ~n2071;
  assign n2075 = ~pi72  & ~n2074;
  assign n2076 = ~n2073 & ~n2075;
  assign n2077 = ~n2069 & n2076;
  assign n2078 = n2069 & ~n2076;
  assign n2079 = ~n2077 & ~n2078;
  assign n2080 = ~n2047 & ~n2079;
  assign n2081 = ~n2069 & ~n2076;
  assign n2082 = pi70  & pi71 ;
  assign n2083 = pi72  & ~n2074;
  assign n2084 = ~n2082 & ~n2083;
  assign n2085 = pi67  & pi68 ;
  assign n2086 = pi69  & ~n2067;
  assign n2087 = ~n2085 & ~n2086;
  assign n2088 = n2084 & ~n2087;
  assign n2089 = ~n2084 & n2087;
  assign n2090 = ~n2088 & ~n2089;
  assign n2091 = n2081 & n2090;
  assign n2092 = ~n2081 & ~n2090;
  assign n2093 = ~n2091 & ~n2092;
  assign n2094 = ~n2080 & n2093;
  assign n2095 = n2062 & ~n2094;
  assign n2096 = n2080 & ~n2093;
  assign n2097 = ~n2095 & ~n2096;
  assign n2098 = n2056 & ~n2057;
  assign n2099 = ~n2054 & ~n2098;
  assign n2100 = ~n2097 & ~n2099;
  assign n2101 = n2097 & n2099;
  assign n2102 = ~n2100 & ~n2101;
  assign n2103 = n2081 & ~n2084;
  assign n2104 = n2087 & ~n2103;
  assign n2105 = ~n2081 & n2084;
  assign n2106 = ~n2104 & ~n2105;
  assign n2107 = ~n2102 & n2106;
  assign n2108 = n2102 & ~n2106;
  assign n2109 = ~n2107 & ~n2108;
  assign n2110 = ~n2030 & ~n2109;
  assign n2111 = n2030 & n2109;
  assign n2112 = n2047 & n2079;
  assign n2113 = ~n2080 & ~n2112;
  assign n2114 = n1968 & n1985;
  assign n2115 = ~n1986 & ~n2114;
  assign n2116 = n2113 & n2115;
  assign n2117 = n2080 & ~n2090;
  assign n2118 = ~n2094 & ~n2117;
  assign n2119 = n2062 & ~n2118;
  assign n2120 = ~n2062 & n2118;
  assign n2121 = ~n2119 & ~n2120;
  assign n2122 = n2116 & ~n2121;
  assign n2123 = ~n2116 & n2121;
  assign n2124 = ~n2002 & ~n2003;
  assign n2125 = ~n2016 & n2124;
  assign n2126 = n2016 & ~n2124;
  assign n2127 = ~n2125 & ~n2126;
  assign n2128 = ~n2123 & n2127;
  assign n2129 = ~n2122 & ~n2128;
  assign n2130 = ~n2111 & ~n2129;
  assign n2131 = ~n2110 & ~n2130;
  assign n2132 = ~n2101 & n2106;
  assign n2133 = ~n2100 & ~n2132;
  assign n2134 = ~n2131 & ~n2133;
  assign n2135 = n2131 & n2133;
  assign n2136 = ~n2022 & n2027;
  assign n2137 = ~n2021 & ~n2136;
  assign n2138 = ~n2135 & ~n2137;
  assign n2139 = ~n2134 & ~n2138;
  assign n2140 = ~n2134 & ~n2135;
  assign n2141 = n2137 & ~n2140;
  assign n2142 = ~n2134 & n2138;
  assign n2143 = ~n2141 & ~n2142;
  assign n2144 = ~n1946 & ~n1947;
  assign n2145 = n1949 & ~n2144;
  assign n2146 = ~n1946 & n1950;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~n2143 & ~n2147;
  assign n2149 = n2143 & n2147;
  assign n2150 = ~n1922 & ~n1923;
  assign n2151 = ~n1941 & n2150;
  assign n2152 = n1941 & ~n2150;
  assign n2153 = ~n2151 & ~n2152;
  assign n2154 = ~n2110 & ~n2111;
  assign n2155 = ~n2129 & n2154;
  assign n2156 = n2129 & ~n2154;
  assign n2157 = ~n2155 & ~n2156;
  assign n2158 = ~n2153 & ~n2157;
  assign n2159 = n2153 & n2157;
  assign n2160 = ~n2113 & ~n2115;
  assign n2161 = ~n2116 & ~n2160;
  assign n2162 = ~n1925 & ~n1927;
  assign n2163 = ~n1928 & ~n2162;
  assign n2164 = n2161 & n2163;
  assign n2165 = ~n2122 & ~n2123;
  assign n2166 = ~n2127 & n2165;
  assign n2167 = n2127 & ~n2165;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = n2164 & ~n2168;
  assign n2170 = ~n2164 & n2168;
  assign n2171 = ~n1934 & ~n1935;
  assign n2172 = ~n1939 & n2171;
  assign n2173 = n1939 & ~n2171;
  assign n2174 = ~n2172 & ~n2173;
  assign n2175 = ~n2170 & ~n2174;
  assign n2176 = ~n2169 & ~n2175;
  assign n2177 = ~n2159 & n2176;
  assign n2178 = ~n2158 & ~n2177;
  assign n2179 = ~n2149 & ~n2178;
  assign n2180 = ~n2148 & ~n2179;
  assign n2181 = n2139 & ~n2180;
  assign n2182 = ~n2139 & n2180;
  assign n2183 = ~n2181 & ~n2182;
  assign n2184 = n1951 & n2183;
  assign n2185 = ~n1951 & ~n2183;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = n1763 & ~n2186;
  assign n2188 = ~n1763 & n2186;
  assign n2189 = ~n2148 & ~n2149;
  assign n2190 = ~n2178 & n2189;
  assign n2191 = n2178 & ~n2189;
  assign n2192 = ~n2190 & ~n2191;
  assign n2193 = ~n1725 & ~n1726;
  assign n2194 = n1758 & n2193;
  assign n2195 = ~n1758 & ~n2193;
  assign n2196 = ~n2194 & ~n2195;
  assign n2197 = ~n2192 & n2196;
  assign n2198 = n2192 & ~n2196;
  assign n2199 = ~n1737 & ~n1738;
  assign n2200 = ~n1756 & n2199;
  assign n2201 = n1756 & ~n2199;
  assign n2202 = ~n2200 & ~n2201;
  assign n2203 = ~n2158 & ~n2159;
  assign n2204 = ~n2176 & n2203;
  assign n2205 = n2176 & ~n2203;
  assign n2206 = ~n2204 & ~n2205;
  assign n2207 = ~n2202 & ~n2206;
  assign n2208 = n2202 & n2206;
  assign n2209 = n2161 & ~n2163;
  assign n2210 = ~n2161 & n2163;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = n1741 & ~n1743;
  assign n2213 = ~n1744 & ~n2212;
  assign n2214 = ~n2211 & n2213;
  assign n2215 = ~n2169 & ~n2170;
  assign n2216 = n2174 & n2215;
  assign n2217 = ~n2174 & ~n2215;
  assign n2218 = ~n2216 & ~n2217;
  assign n2219 = n2214 & ~n2218;
  assign n2220 = ~n2214 & n2218;
  assign n2221 = ~n1749 & ~n1750;
  assign n2222 = n1754 & n2221;
  assign n2223 = ~n1754 & ~n2221;
  assign n2224 = ~n2222 & ~n2223;
  assign n2225 = ~n2220 & ~n2224;
  assign n2226 = ~n2219 & ~n2225;
  assign n2227 = ~n2208 & n2226;
  assign n2228 = ~n2207 & ~n2227;
  assign n2229 = ~n2198 & n2228;
  assign n2230 = ~n2197 & ~n2229;
  assign n2231 = ~n2188 & ~n2230;
  assign n2232 = ~n2187 & ~n2231;
  assign n2233 = n1951 & ~n2182;
  assign n2234 = ~n2181 & ~n2233;
  assign n2235 = ~n1715 & n1760;
  assign n2236 = ~n1714 & ~n2235;
  assign n2237 = ~n2234 & n2236;
  assign n2238 = n2234 & ~n2236;
  assign n2239 = ~n2237 & ~n2238;
  assign n2240 = ~n2232 & ~n2239;
  assign n2241 = n2232 & n2239;
  assign n2242 = ~n2240 & ~n2241;
  assign n2243 = ~n1422 & n2242;
  assign n2244 = n1422 & ~n2242;
  assign n2245 = n1190 & ~n1416;
  assign n2246 = ~n1190 & n1416;
  assign n2247 = ~n2245 & ~n2246;
  assign n2248 = n1420 & n2247;
  assign n2249 = ~n1420 & ~n2247;
  assign n2250 = ~n2248 & ~n2249;
  assign n2251 = ~n2187 & ~n2188;
  assign n2252 = ~n2230 & n2251;
  assign n2253 = n2230 & ~n2251;
  assign n2254 = ~n2252 & ~n2253;
  assign n2255 = n2250 & ~n2254;
  assign n2256 = ~n2250 & n2254;
  assign n2257 = ~n2197 & ~n2198;
  assign n2258 = n2228 & n2257;
  assign n2259 = ~n2228 & ~n2257;
  assign n2260 = ~n2258 & ~n2259;
  assign n2261 = ~n1384 & ~n1385;
  assign n2262 = ~n1414 & n2261;
  assign n2263 = n1414 & ~n2261;
  assign n2264 = ~n2262 & ~n2263;
  assign n2265 = n2260 & ~n2264;
  assign n2266 = ~n2260 & n2264;
  assign n2267 = ~n1394 & ~n1395;
  assign n2268 = ~n1412 & n2267;
  assign n2269 = n1412 & ~n2267;
  assign n2270 = ~n2268 & ~n2269;
  assign n2271 = ~n2207 & ~n2208;
  assign n2272 = ~n2226 & n2271;
  assign n2273 = n2226 & ~n2271;
  assign n2274 = ~n2272 & ~n2273;
  assign n2275 = ~n2270 & ~n2274;
  assign n2276 = n2270 & n2274;
  assign n2277 = n1397 & ~n1399;
  assign n2278 = ~n1397 & n1399;
  assign n2279 = ~n2277 & ~n2278;
  assign n2280 = n2211 & ~n2213;
  assign n2281 = ~n2214 & ~n2280;
  assign n2282 = ~n2279 & n2281;
  assign n2283 = ~n2219 & ~n2220;
  assign n2284 = ~n2224 & n2283;
  assign n2285 = n2224 & ~n2283;
  assign n2286 = ~n2284 & ~n2285;
  assign n2287 = n2282 & n2286;
  assign n2288 = ~n2282 & ~n2286;
  assign n2289 = ~n1405 & ~n1406;
  assign n2290 = n1410 & n2289;
  assign n2291 = ~n1410 & ~n2289;
  assign n2292 = ~n2290 & ~n2291;
  assign n2293 = ~n2288 & ~n2292;
  assign n2294 = ~n2287 & ~n2293;
  assign n2295 = ~n2276 & n2294;
  assign n2296 = ~n2275 & ~n2295;
  assign n2297 = ~n2266 & n2296;
  assign n2298 = ~n2265 & ~n2297;
  assign n2299 = ~n2256 & n2298;
  assign n2300 = ~n2255 & ~n2299;
  assign n2301 = ~n2244 & ~n2300;
  assign n2302 = ~n2243 & ~n2301;
  assign n2303 = ~n2232 & ~n2237;
  assign n2304 = ~n2238 & ~n2303;
  assign n2305 = n2302 & ~n2304;
  assign n2306 = ~n2302 & n2304;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = ~pi853  & pi854 ;
  assign n2309 = pi853  & ~pi854 ;
  assign n2310 = pi855  & ~n2308;
  assign n2311 = ~n2309 & n2310;
  assign n2312 = ~n2308 & ~n2309;
  assign n2313 = ~pi855  & ~n2312;
  assign n2314 = ~n2311 & ~n2313;
  assign n2315 = ~pi856  & pi857 ;
  assign n2316 = pi856  & ~pi857 ;
  assign n2317 = pi858  & ~n2315;
  assign n2318 = ~n2316 & n2317;
  assign n2319 = ~n2315 & ~n2316;
  assign n2320 = ~pi858  & ~n2319;
  assign n2321 = ~n2318 & ~n2320;
  assign n2322 = ~n2314 & n2321;
  assign n2323 = n2314 & ~n2321;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~pi847  & pi848 ;
  assign n2326 = pi847  & ~pi848 ;
  assign n2327 = pi849  & ~n2325;
  assign n2328 = ~n2326 & n2327;
  assign n2329 = ~n2325 & ~n2326;
  assign n2330 = ~pi849  & ~n2329;
  assign n2331 = ~n2328 & ~n2330;
  assign n2332 = ~pi850  & pi851 ;
  assign n2333 = pi850  & ~pi851 ;
  assign n2334 = pi852  & ~n2332;
  assign n2335 = ~n2333 & n2334;
  assign n2336 = ~n2332 & ~n2333;
  assign n2337 = ~pi852  & ~n2336;
  assign n2338 = ~n2335 & ~n2337;
  assign n2339 = ~n2331 & n2338;
  assign n2340 = n2331 & ~n2338;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = ~n2324 & ~n2341;
  assign n2343 = pi856  & pi857 ;
  assign n2344 = pi858  & ~n2319;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = pi853  & pi854 ;
  assign n2347 = pi855  & ~n2312;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = ~n2345 & ~n2348;
  assign n2350 = ~n2324 & n2349;
  assign n2351 = ~n2314 & ~n2321;
  assign n2352 = n2345 & n2348;
  assign n2353 = ~n2349 & ~n2352;
  assign n2354 = n2351 & n2353;
  assign n2355 = ~n2351 & ~n2353;
  assign n2356 = ~n2350 & ~n2354;
  assign n2357 = ~n2355 & n2356;
  assign n2358 = n2342 & n2357;
  assign n2359 = ~n2342 & ~n2357;
  assign n2360 = pi850  & pi851 ;
  assign n2361 = pi852  & ~n2336;
  assign n2362 = ~n2360 & ~n2361;
  assign n2363 = pi847  & pi848 ;
  assign n2364 = pi849  & ~n2329;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = ~n2362 & n2365;
  assign n2367 = n2362 & ~n2365;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = ~n2331 & ~n2338;
  assign n2370 = n2368 & n2369;
  assign n2371 = ~n2368 & ~n2369;
  assign n2372 = ~n2370 & ~n2371;
  assign n2373 = ~n2359 & ~n2372;
  assign n2374 = ~n2358 & ~n2373;
  assign n2375 = n2351 & ~n2352;
  assign n2376 = ~n2349 & ~n2375;
  assign n2377 = ~n2374 & ~n2376;
  assign n2378 = n2374 & n2376;
  assign n2379 = ~n2377 & ~n2378;
  assign n2380 = ~n2362 & n2369;
  assign n2381 = n2365 & ~n2380;
  assign n2382 = n2362 & ~n2369;
  assign n2383 = ~n2381 & ~n2382;
  assign n2384 = ~n2379 & n2383;
  assign n2385 = n2379 & ~n2383;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = ~pi865  & pi866 ;
  assign n2388 = pi865  & ~pi866 ;
  assign n2389 = pi867  & ~n2387;
  assign n2390 = ~n2388 & n2389;
  assign n2391 = ~n2387 & ~n2388;
  assign n2392 = ~pi867  & ~n2391;
  assign n2393 = ~n2390 & ~n2392;
  assign n2394 = ~pi868  & pi869 ;
  assign n2395 = pi868  & ~pi869 ;
  assign n2396 = pi870  & ~n2394;
  assign n2397 = ~n2395 & n2396;
  assign n2398 = ~n2394 & ~n2395;
  assign n2399 = ~pi870  & ~n2398;
  assign n2400 = ~n2397 & ~n2399;
  assign n2401 = ~n2393 & n2400;
  assign n2402 = n2393 & ~n2400;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = ~pi859  & pi860 ;
  assign n2405 = pi859  & ~pi860 ;
  assign n2406 = pi861  & ~n2404;
  assign n2407 = ~n2405 & n2406;
  assign n2408 = ~n2404 & ~n2405;
  assign n2409 = ~pi861  & ~n2408;
  assign n2410 = ~n2407 & ~n2409;
  assign n2411 = ~pi862  & pi863 ;
  assign n2412 = pi862  & ~pi863 ;
  assign n2413 = pi864  & ~n2411;
  assign n2414 = ~n2412 & n2413;
  assign n2415 = ~n2411 & ~n2412;
  assign n2416 = ~pi864  & ~n2415;
  assign n2417 = ~n2414 & ~n2416;
  assign n2418 = ~n2410 & n2417;
  assign n2419 = n2410 & ~n2417;
  assign n2420 = ~n2418 & ~n2419;
  assign n2421 = ~n2403 & ~n2420;
  assign n2422 = pi868  & pi869 ;
  assign n2423 = pi870  & ~n2398;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = pi865  & pi866 ;
  assign n2426 = pi867  & ~n2391;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = n2424 & ~n2427;
  assign n2429 = ~n2424 & n2427;
  assign n2430 = ~n2428 & ~n2429;
  assign n2431 = n2421 & ~n2430;
  assign n2432 = ~n2393 & ~n2400;
  assign n2433 = n2430 & n2432;
  assign n2434 = ~n2430 & ~n2432;
  assign n2435 = ~n2421 & ~n2433;
  assign n2436 = ~n2434 & n2435;
  assign n2437 = pi862  & pi863 ;
  assign n2438 = pi864  & ~n2415;
  assign n2439 = ~n2437 & ~n2438;
  assign n2440 = pi859  & pi860 ;
  assign n2441 = pi861  & ~n2408;
  assign n2442 = ~n2440 & ~n2441;
  assign n2443 = ~n2439 & ~n2442;
  assign n2444 = ~n2420 & n2443;
  assign n2445 = ~n2410 & ~n2417;
  assign n2446 = n2439 & n2442;
  assign n2447 = ~n2443 & ~n2446;
  assign n2448 = n2445 & n2447;
  assign n2449 = ~n2445 & ~n2447;
  assign n2450 = ~n2444 & ~n2448;
  assign n2451 = ~n2449 & n2450;
  assign n2452 = ~n2436 & n2451;
  assign n2453 = ~n2431 & ~n2452;
  assign n2454 = ~n2424 & n2432;
  assign n2455 = n2427 & ~n2454;
  assign n2456 = n2424 & ~n2432;
  assign n2457 = ~n2455 & ~n2456;
  assign n2458 = ~n2453 & n2457;
  assign n2459 = n2453 & ~n2457;
  assign n2460 = ~n2458 & ~n2459;
  assign n2461 = n2445 & ~n2446;
  assign n2462 = ~n2443 & ~n2461;
  assign n2463 = n2460 & ~n2462;
  assign n2464 = ~n2460 & n2462;
  assign n2465 = ~n2463 & ~n2464;
  assign n2466 = n2386 & ~n2465;
  assign n2467 = ~n2386 & n2465;
  assign n2468 = n2403 & n2420;
  assign n2469 = ~n2421 & ~n2468;
  assign n2470 = n2324 & n2341;
  assign n2471 = ~n2342 & ~n2470;
  assign n2472 = n2469 & n2471;
  assign n2473 = ~n2431 & ~n2436;
  assign n2474 = n2451 & n2473;
  assign n2475 = ~n2451 & ~n2473;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = n2472 & n2476;
  assign n2478 = ~n2472 & ~n2476;
  assign n2479 = ~n2358 & ~n2359;
  assign n2480 = ~n2372 & n2479;
  assign n2481 = n2372 & ~n2479;
  assign n2482 = ~n2480 & ~n2481;
  assign n2483 = ~n2478 & n2482;
  assign n2484 = ~n2477 & ~n2483;
  assign n2485 = ~n2467 & n2484;
  assign n2486 = ~n2466 & ~n2485;
  assign n2487 = ~n2459 & ~n2462;
  assign n2488 = ~n2458 & ~n2487;
  assign n2489 = ~n2486 & n2488;
  assign n2490 = n2486 & ~n2488;
  assign n2491 = ~n2378 & n2383;
  assign n2492 = ~n2377 & ~n2491;
  assign n2493 = ~n2490 & n2492;
  assign n2494 = ~n2489 & ~n2493;
  assign n2495 = ~pi877  & pi878 ;
  assign n2496 = pi877  & ~pi878 ;
  assign n2497 = pi879  & ~n2495;
  assign n2498 = ~n2496 & n2497;
  assign n2499 = ~n2495 & ~n2496;
  assign n2500 = ~pi879  & ~n2499;
  assign n2501 = ~n2498 & ~n2500;
  assign n2502 = ~pi880  & pi881 ;
  assign n2503 = pi880  & ~pi881 ;
  assign n2504 = pi882  & ~n2502;
  assign n2505 = ~n2503 & n2504;
  assign n2506 = ~n2502 & ~n2503;
  assign n2507 = ~pi882  & ~n2506;
  assign n2508 = ~n2505 & ~n2507;
  assign n2509 = ~n2501 & n2508;
  assign n2510 = n2501 & ~n2508;
  assign n2511 = ~n2509 & ~n2510;
  assign n2512 = ~pi871  & pi872 ;
  assign n2513 = pi871  & ~pi872 ;
  assign n2514 = pi873  & ~n2512;
  assign n2515 = ~n2513 & n2514;
  assign n2516 = ~n2512 & ~n2513;
  assign n2517 = ~pi873  & ~n2516;
  assign n2518 = ~n2515 & ~n2517;
  assign n2519 = ~pi874  & pi875 ;
  assign n2520 = pi874  & ~pi875 ;
  assign n2521 = pi876  & ~n2519;
  assign n2522 = ~n2520 & n2521;
  assign n2523 = ~n2519 & ~n2520;
  assign n2524 = ~pi876  & ~n2523;
  assign n2525 = ~n2522 & ~n2524;
  assign n2526 = ~n2518 & n2525;
  assign n2527 = n2518 & ~n2525;
  assign n2528 = ~n2526 & ~n2527;
  assign n2529 = ~n2511 & ~n2528;
  assign n2530 = pi880  & pi881 ;
  assign n2531 = pi882  & ~n2506;
  assign n2532 = ~n2530 & ~n2531;
  assign n2533 = pi877  & pi878 ;
  assign n2534 = pi879  & ~n2499;
  assign n2535 = ~n2533 & ~n2534;
  assign n2536 = ~n2532 & ~n2535;
  assign n2537 = ~n2511 & n2536;
  assign n2538 = ~n2501 & ~n2508;
  assign n2539 = n2532 & n2535;
  assign n2540 = ~n2536 & ~n2539;
  assign n2541 = n2538 & n2540;
  assign n2542 = ~n2538 & ~n2540;
  assign n2543 = ~n2537 & ~n2541;
  assign n2544 = ~n2542 & n2543;
  assign n2545 = n2529 & n2544;
  assign n2546 = ~n2529 & ~n2544;
  assign n2547 = pi874  & pi875 ;
  assign n2548 = pi876  & ~n2523;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = pi871  & pi872 ;
  assign n2551 = pi873  & ~n2516;
  assign n2552 = ~n2550 & ~n2551;
  assign n2553 = ~n2549 & n2552;
  assign n2554 = n2549 & ~n2552;
  assign n2555 = ~n2553 & ~n2554;
  assign n2556 = ~n2518 & ~n2525;
  assign n2557 = n2555 & n2556;
  assign n2558 = ~n2555 & ~n2556;
  assign n2559 = ~n2557 & ~n2558;
  assign n2560 = ~n2546 & ~n2559;
  assign n2561 = ~n2545 & ~n2560;
  assign n2562 = n2538 & ~n2539;
  assign n2563 = ~n2536 & ~n2562;
  assign n2564 = ~n2561 & ~n2563;
  assign n2565 = n2561 & n2563;
  assign n2566 = ~n2564 & ~n2565;
  assign n2567 = ~n2549 & n2556;
  assign n2568 = n2552 & ~n2567;
  assign n2569 = n2549 & ~n2556;
  assign n2570 = ~n2568 & ~n2569;
  assign n2571 = ~n2566 & n2570;
  assign n2572 = n2566 & ~n2570;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = ~pi889  & pi890 ;
  assign n2575 = pi889  & ~pi890 ;
  assign n2576 = pi891  & ~n2574;
  assign n2577 = ~n2575 & n2576;
  assign n2578 = ~n2574 & ~n2575;
  assign n2579 = ~pi891  & ~n2578;
  assign n2580 = ~n2577 & ~n2579;
  assign n2581 = ~pi892  & pi893 ;
  assign n2582 = pi892  & ~pi893 ;
  assign n2583 = pi894  & ~n2581;
  assign n2584 = ~n2582 & n2583;
  assign n2585 = ~n2581 & ~n2582;
  assign n2586 = ~pi894  & ~n2585;
  assign n2587 = ~n2584 & ~n2586;
  assign n2588 = ~n2580 & n2587;
  assign n2589 = n2580 & ~n2587;
  assign n2590 = ~n2588 & ~n2589;
  assign n2591 = ~pi883  & pi884 ;
  assign n2592 = pi883  & ~pi884 ;
  assign n2593 = pi885  & ~n2591;
  assign n2594 = ~n2592 & n2593;
  assign n2595 = ~n2591 & ~n2592;
  assign n2596 = ~pi885  & ~n2595;
  assign n2597 = ~n2594 & ~n2596;
  assign n2598 = ~pi886  & pi887 ;
  assign n2599 = pi886  & ~pi887 ;
  assign n2600 = pi888  & ~n2598;
  assign n2601 = ~n2599 & n2600;
  assign n2602 = ~n2598 & ~n2599;
  assign n2603 = ~pi888  & ~n2602;
  assign n2604 = ~n2601 & ~n2603;
  assign n2605 = ~n2597 & n2604;
  assign n2606 = n2597 & ~n2604;
  assign n2607 = ~n2605 & ~n2606;
  assign n2608 = ~n2590 & ~n2607;
  assign n2609 = pi892  & pi893 ;
  assign n2610 = pi894  & ~n2585;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = pi889  & pi890 ;
  assign n2613 = pi891  & ~n2578;
  assign n2614 = ~n2612 & ~n2613;
  assign n2615 = n2611 & ~n2614;
  assign n2616 = ~n2611 & n2614;
  assign n2617 = ~n2615 & ~n2616;
  assign n2618 = n2608 & ~n2617;
  assign n2619 = ~n2580 & ~n2587;
  assign n2620 = n2617 & n2619;
  assign n2621 = ~n2617 & ~n2619;
  assign n2622 = ~n2608 & ~n2620;
  assign n2623 = ~n2621 & n2622;
  assign n2624 = pi886  & pi887 ;
  assign n2625 = pi888  & ~n2602;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = pi883  & pi884 ;
  assign n2628 = pi885  & ~n2595;
  assign n2629 = ~n2627 & ~n2628;
  assign n2630 = ~n2626 & ~n2629;
  assign n2631 = ~n2607 & n2630;
  assign n2632 = ~n2597 & ~n2604;
  assign n2633 = n2626 & n2629;
  assign n2634 = ~n2630 & ~n2633;
  assign n2635 = n2632 & n2634;
  assign n2636 = ~n2632 & ~n2634;
  assign n2637 = ~n2631 & ~n2635;
  assign n2638 = ~n2636 & n2637;
  assign n2639 = ~n2623 & n2638;
  assign n2640 = ~n2618 & ~n2639;
  assign n2641 = ~n2611 & n2619;
  assign n2642 = n2614 & ~n2641;
  assign n2643 = n2611 & ~n2619;
  assign n2644 = ~n2642 & ~n2643;
  assign n2645 = ~n2640 & n2644;
  assign n2646 = n2640 & ~n2644;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = n2632 & ~n2633;
  assign n2649 = ~n2630 & ~n2648;
  assign n2650 = n2647 & ~n2649;
  assign n2651 = ~n2647 & n2649;
  assign n2652 = ~n2650 & ~n2651;
  assign n2653 = n2573 & ~n2652;
  assign n2654 = ~n2573 & n2652;
  assign n2655 = n2590 & n2607;
  assign n2656 = ~n2608 & ~n2655;
  assign n2657 = n2511 & n2528;
  assign n2658 = ~n2529 & ~n2657;
  assign n2659 = n2656 & n2658;
  assign n2660 = ~n2618 & ~n2623;
  assign n2661 = n2638 & n2660;
  assign n2662 = ~n2638 & ~n2660;
  assign n2663 = ~n2661 & ~n2662;
  assign n2664 = n2659 & n2663;
  assign n2665 = ~n2659 & ~n2663;
  assign n2666 = ~n2545 & ~n2546;
  assign n2667 = ~n2559 & n2666;
  assign n2668 = n2559 & ~n2666;
  assign n2669 = ~n2667 & ~n2668;
  assign n2670 = ~n2665 & n2669;
  assign n2671 = ~n2664 & ~n2670;
  assign n2672 = ~n2654 & n2671;
  assign n2673 = ~n2653 & ~n2672;
  assign n2674 = ~n2646 & ~n2649;
  assign n2675 = ~n2645 & ~n2674;
  assign n2676 = ~n2673 & n2675;
  assign n2677 = n2673 & ~n2675;
  assign n2678 = ~n2565 & n2570;
  assign n2679 = ~n2564 & ~n2678;
  assign n2680 = ~n2677 & n2679;
  assign n2681 = ~n2676 & ~n2680;
  assign n2682 = ~n2676 & ~n2677;
  assign n2683 = n2679 & n2682;
  assign n2684 = ~n2679 & ~n2682;
  assign n2685 = ~n2683 & ~n2684;
  assign n2686 = ~n2489 & ~n2490;
  assign n2687 = n2492 & n2686;
  assign n2688 = ~n2492 & ~n2686;
  assign n2689 = ~n2687 & ~n2688;
  assign n2690 = ~n2685 & ~n2689;
  assign n2691 = n2685 & n2689;
  assign n2692 = ~n2466 & ~n2467;
  assign n2693 = ~n2484 & n2692;
  assign n2694 = n2484 & ~n2692;
  assign n2695 = ~n2693 & ~n2694;
  assign n2696 = ~n2653 & ~n2654;
  assign n2697 = ~n2671 & n2696;
  assign n2698 = n2671 & ~n2696;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = ~n2695 & ~n2699;
  assign n2701 = n2695 & n2699;
  assign n2702 = ~n2656 & ~n2658;
  assign n2703 = ~n2659 & ~n2702;
  assign n2704 = ~n2469 & ~n2471;
  assign n2705 = ~n2472 & ~n2704;
  assign n2706 = n2703 & n2705;
  assign n2707 = ~n2664 & ~n2665;
  assign n2708 = ~n2669 & n2707;
  assign n2709 = n2669 & ~n2707;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = n2706 & ~n2710;
  assign n2712 = ~n2706 & n2710;
  assign n2713 = ~n2477 & ~n2478;
  assign n2714 = ~n2482 & n2713;
  assign n2715 = n2482 & ~n2713;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = ~n2712 & ~n2716;
  assign n2718 = ~n2711 & ~n2717;
  assign n2719 = ~n2701 & n2718;
  assign n2720 = ~n2700 & ~n2719;
  assign n2721 = ~n2691 & n2720;
  assign n2722 = ~n2690 & ~n2721;
  assign n2723 = ~n2681 & n2722;
  assign n2724 = n2681 & ~n2722;
  assign n2725 = ~n2723 & ~n2724;
  assign n2726 = n2494 & n2725;
  assign n2727 = ~n2494 & ~n2725;
  assign n2728 = ~n2726 & ~n2727;
  assign n2729 = ~pi901  & pi902 ;
  assign n2730 = pi901  & ~pi902 ;
  assign n2731 = pi903  & ~n2729;
  assign n2732 = ~n2730 & n2731;
  assign n2733 = ~n2729 & ~n2730;
  assign n2734 = ~pi903  & ~n2733;
  assign n2735 = ~n2732 & ~n2734;
  assign n2736 = ~pi904  & pi905 ;
  assign n2737 = pi904  & ~pi905 ;
  assign n2738 = pi906  & ~n2736;
  assign n2739 = ~n2737 & n2738;
  assign n2740 = ~n2736 & ~n2737;
  assign n2741 = ~pi906  & ~n2740;
  assign n2742 = ~n2739 & ~n2741;
  assign n2743 = ~n2735 & n2742;
  assign n2744 = n2735 & ~n2742;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = ~pi895  & pi896 ;
  assign n2747 = pi895  & ~pi896 ;
  assign n2748 = pi897  & ~n2746;
  assign n2749 = ~n2747 & n2748;
  assign n2750 = ~n2746 & ~n2747;
  assign n2751 = ~pi897  & ~n2750;
  assign n2752 = ~n2749 & ~n2751;
  assign n2753 = ~pi898  & pi899 ;
  assign n2754 = pi898  & ~pi899 ;
  assign n2755 = pi900  & ~n2753;
  assign n2756 = ~n2754 & n2755;
  assign n2757 = ~n2753 & ~n2754;
  assign n2758 = ~pi900  & ~n2757;
  assign n2759 = ~n2756 & ~n2758;
  assign n2760 = ~n2752 & n2759;
  assign n2761 = n2752 & ~n2759;
  assign n2762 = ~n2760 & ~n2761;
  assign n2763 = ~n2745 & ~n2762;
  assign n2764 = pi904  & pi905 ;
  assign n2765 = pi906  & ~n2740;
  assign n2766 = ~n2764 & ~n2765;
  assign n2767 = pi901  & pi902 ;
  assign n2768 = pi903  & ~n2733;
  assign n2769 = ~n2767 & ~n2768;
  assign n2770 = ~n2766 & ~n2769;
  assign n2771 = ~n2745 & n2770;
  assign n2772 = ~n2735 & ~n2742;
  assign n2773 = n2766 & n2769;
  assign n2774 = ~n2770 & ~n2773;
  assign n2775 = n2772 & n2774;
  assign n2776 = ~n2772 & ~n2774;
  assign n2777 = ~n2771 & ~n2775;
  assign n2778 = ~n2776 & n2777;
  assign n2779 = n2763 & n2778;
  assign n2780 = ~n2763 & ~n2778;
  assign n2781 = pi898  & pi899 ;
  assign n2782 = pi900  & ~n2757;
  assign n2783 = ~n2781 & ~n2782;
  assign n2784 = pi895  & pi896 ;
  assign n2785 = pi897  & ~n2750;
  assign n2786 = ~n2784 & ~n2785;
  assign n2787 = ~n2783 & n2786;
  assign n2788 = n2783 & ~n2786;
  assign n2789 = ~n2787 & ~n2788;
  assign n2790 = ~n2752 & ~n2759;
  assign n2791 = n2789 & n2790;
  assign n2792 = ~n2789 & ~n2790;
  assign n2793 = ~n2791 & ~n2792;
  assign n2794 = ~n2780 & ~n2793;
  assign n2795 = ~n2779 & ~n2794;
  assign n2796 = n2772 & ~n2773;
  assign n2797 = ~n2770 & ~n2796;
  assign n2798 = ~n2795 & ~n2797;
  assign n2799 = n2795 & n2797;
  assign n2800 = ~n2798 & ~n2799;
  assign n2801 = ~n2783 & n2790;
  assign n2802 = n2786 & ~n2801;
  assign n2803 = n2783 & ~n2790;
  assign n2804 = ~n2802 & ~n2803;
  assign n2805 = ~n2800 & n2804;
  assign n2806 = n2800 & ~n2804;
  assign n2807 = ~n2805 & ~n2806;
  assign n2808 = ~pi913  & pi914 ;
  assign n2809 = pi913  & ~pi914 ;
  assign n2810 = pi915  & ~n2808;
  assign n2811 = ~n2809 & n2810;
  assign n2812 = ~n2808 & ~n2809;
  assign n2813 = ~pi915  & ~n2812;
  assign n2814 = ~n2811 & ~n2813;
  assign n2815 = ~pi916  & pi917 ;
  assign n2816 = pi916  & ~pi917 ;
  assign n2817 = pi918  & ~n2815;
  assign n2818 = ~n2816 & n2817;
  assign n2819 = ~n2815 & ~n2816;
  assign n2820 = ~pi918  & ~n2819;
  assign n2821 = ~n2818 & ~n2820;
  assign n2822 = ~n2814 & n2821;
  assign n2823 = n2814 & ~n2821;
  assign n2824 = ~n2822 & ~n2823;
  assign n2825 = ~pi907  & pi908 ;
  assign n2826 = pi907  & ~pi908 ;
  assign n2827 = pi909  & ~n2825;
  assign n2828 = ~n2826 & n2827;
  assign n2829 = ~n2825 & ~n2826;
  assign n2830 = ~pi909  & ~n2829;
  assign n2831 = ~n2828 & ~n2830;
  assign n2832 = ~pi910  & pi911 ;
  assign n2833 = pi910  & ~pi911 ;
  assign n2834 = pi912  & ~n2832;
  assign n2835 = ~n2833 & n2834;
  assign n2836 = ~n2832 & ~n2833;
  assign n2837 = ~pi912  & ~n2836;
  assign n2838 = ~n2835 & ~n2837;
  assign n2839 = ~n2831 & n2838;
  assign n2840 = n2831 & ~n2838;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = ~n2824 & ~n2841;
  assign n2843 = pi916  & pi917 ;
  assign n2844 = pi918  & ~n2819;
  assign n2845 = ~n2843 & ~n2844;
  assign n2846 = pi913  & pi914 ;
  assign n2847 = pi915  & ~n2812;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = n2845 & ~n2848;
  assign n2850 = ~n2845 & n2848;
  assign n2851 = ~n2849 & ~n2850;
  assign n2852 = n2842 & ~n2851;
  assign n2853 = ~n2814 & ~n2821;
  assign n2854 = n2851 & n2853;
  assign n2855 = ~n2851 & ~n2853;
  assign n2856 = ~n2842 & ~n2854;
  assign n2857 = ~n2855 & n2856;
  assign n2858 = pi910  & pi911 ;
  assign n2859 = pi912  & ~n2836;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = pi907  & pi908 ;
  assign n2862 = pi909  & ~n2829;
  assign n2863 = ~n2861 & ~n2862;
  assign n2864 = ~n2860 & ~n2863;
  assign n2865 = ~n2841 & n2864;
  assign n2866 = ~n2831 & ~n2838;
  assign n2867 = n2860 & n2863;
  assign n2868 = ~n2864 & ~n2867;
  assign n2869 = n2866 & n2868;
  assign n2870 = ~n2866 & ~n2868;
  assign n2871 = ~n2865 & ~n2869;
  assign n2872 = ~n2870 & n2871;
  assign n2873 = ~n2857 & n2872;
  assign n2874 = ~n2852 & ~n2873;
  assign n2875 = ~n2845 & n2853;
  assign n2876 = n2848 & ~n2875;
  assign n2877 = n2845 & ~n2853;
  assign n2878 = ~n2876 & ~n2877;
  assign n2879 = ~n2874 & n2878;
  assign n2880 = n2874 & ~n2878;
  assign n2881 = ~n2879 & ~n2880;
  assign n2882 = n2866 & ~n2867;
  assign n2883 = ~n2864 & ~n2882;
  assign n2884 = n2881 & ~n2883;
  assign n2885 = ~n2881 & n2883;
  assign n2886 = ~n2884 & ~n2885;
  assign n2887 = n2807 & ~n2886;
  assign n2888 = ~n2807 & n2886;
  assign n2889 = n2824 & n2841;
  assign n2890 = ~n2842 & ~n2889;
  assign n2891 = n2745 & n2762;
  assign n2892 = ~n2763 & ~n2891;
  assign n2893 = n2890 & n2892;
  assign n2894 = ~n2852 & ~n2857;
  assign n2895 = n2872 & n2894;
  assign n2896 = ~n2872 & ~n2894;
  assign n2897 = ~n2895 & ~n2896;
  assign n2898 = n2893 & n2897;
  assign n2899 = ~n2893 & ~n2897;
  assign n2900 = ~n2779 & ~n2780;
  assign n2901 = ~n2793 & n2900;
  assign n2902 = n2793 & ~n2900;
  assign n2903 = ~n2901 & ~n2902;
  assign n2904 = ~n2899 & n2903;
  assign n2905 = ~n2898 & ~n2904;
  assign n2906 = ~n2888 & n2905;
  assign n2907 = ~n2887 & ~n2906;
  assign n2908 = ~n2880 & ~n2883;
  assign n2909 = ~n2879 & ~n2908;
  assign n2910 = ~n2907 & n2909;
  assign n2911 = n2907 & ~n2909;
  assign n2912 = ~n2799 & n2804;
  assign n2913 = ~n2798 & ~n2912;
  assign n2914 = ~n2911 & n2913;
  assign n2915 = ~n2910 & ~n2914;
  assign n2916 = ~pi925  & pi926 ;
  assign n2917 = pi925  & ~pi926 ;
  assign n2918 = pi927  & ~n2916;
  assign n2919 = ~n2917 & n2918;
  assign n2920 = ~n2916 & ~n2917;
  assign n2921 = ~pi927  & ~n2920;
  assign n2922 = ~n2919 & ~n2921;
  assign n2923 = ~pi928  & pi929 ;
  assign n2924 = pi928  & ~pi929 ;
  assign n2925 = pi930  & ~n2923;
  assign n2926 = ~n2924 & n2925;
  assign n2927 = ~n2923 & ~n2924;
  assign n2928 = ~pi930  & ~n2927;
  assign n2929 = ~n2926 & ~n2928;
  assign n2930 = ~n2922 & n2929;
  assign n2931 = n2922 & ~n2929;
  assign n2932 = ~n2930 & ~n2931;
  assign n2933 = ~pi919  & pi920 ;
  assign n2934 = pi919  & ~pi920 ;
  assign n2935 = pi921  & ~n2933;
  assign n2936 = ~n2934 & n2935;
  assign n2937 = ~n2933 & ~n2934;
  assign n2938 = ~pi921  & ~n2937;
  assign n2939 = ~n2936 & ~n2938;
  assign n2940 = ~pi922  & pi923 ;
  assign n2941 = pi922  & ~pi923 ;
  assign n2942 = pi924  & ~n2940;
  assign n2943 = ~n2941 & n2942;
  assign n2944 = ~n2940 & ~n2941;
  assign n2945 = ~pi924  & ~n2944;
  assign n2946 = ~n2943 & ~n2945;
  assign n2947 = ~n2939 & n2946;
  assign n2948 = n2939 & ~n2946;
  assign n2949 = ~n2947 & ~n2948;
  assign n2950 = ~n2932 & ~n2949;
  assign n2951 = pi928  & pi929 ;
  assign n2952 = pi930  & ~n2927;
  assign n2953 = ~n2951 & ~n2952;
  assign n2954 = pi925  & pi926 ;
  assign n2955 = pi927  & ~n2920;
  assign n2956 = ~n2954 & ~n2955;
  assign n2957 = ~n2953 & ~n2956;
  assign n2958 = ~n2932 & n2957;
  assign n2959 = ~n2922 & ~n2929;
  assign n2960 = n2953 & n2956;
  assign n2961 = ~n2957 & ~n2960;
  assign n2962 = n2959 & n2961;
  assign n2963 = ~n2959 & ~n2961;
  assign n2964 = ~n2958 & ~n2962;
  assign n2965 = ~n2963 & n2964;
  assign n2966 = n2950 & n2965;
  assign n2967 = ~n2950 & ~n2965;
  assign n2968 = pi922  & pi923 ;
  assign n2969 = pi924  & ~n2944;
  assign n2970 = ~n2968 & ~n2969;
  assign n2971 = pi919  & pi920 ;
  assign n2972 = pi921  & ~n2937;
  assign n2973 = ~n2971 & ~n2972;
  assign n2974 = ~n2970 & n2973;
  assign n2975 = n2970 & ~n2973;
  assign n2976 = ~n2974 & ~n2975;
  assign n2977 = ~n2939 & ~n2946;
  assign n2978 = n2976 & n2977;
  assign n2979 = ~n2976 & ~n2977;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = ~n2967 & ~n2980;
  assign n2982 = ~n2966 & ~n2981;
  assign n2983 = n2959 & ~n2960;
  assign n2984 = ~n2957 & ~n2983;
  assign n2985 = ~n2982 & ~n2984;
  assign n2986 = n2982 & n2984;
  assign n2987 = ~n2985 & ~n2986;
  assign n2988 = ~n2970 & n2977;
  assign n2989 = n2973 & ~n2988;
  assign n2990 = n2970 & ~n2977;
  assign n2991 = ~n2989 & ~n2990;
  assign n2992 = ~n2987 & n2991;
  assign n2993 = n2987 & ~n2991;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = ~pi937  & pi938 ;
  assign n2996 = pi937  & ~pi938 ;
  assign n2997 = pi939  & ~n2995;
  assign n2998 = ~n2996 & n2997;
  assign n2999 = ~n2995 & ~n2996;
  assign n3000 = ~pi939  & ~n2999;
  assign n3001 = ~n2998 & ~n3000;
  assign n3002 = ~pi940  & pi941 ;
  assign n3003 = pi940  & ~pi941 ;
  assign n3004 = pi942  & ~n3002;
  assign n3005 = ~n3003 & n3004;
  assign n3006 = ~n3002 & ~n3003;
  assign n3007 = ~pi942  & ~n3006;
  assign n3008 = ~n3005 & ~n3007;
  assign n3009 = ~n3001 & n3008;
  assign n3010 = n3001 & ~n3008;
  assign n3011 = ~n3009 & ~n3010;
  assign n3012 = ~pi931  & pi932 ;
  assign n3013 = pi931  & ~pi932 ;
  assign n3014 = pi933  & ~n3012;
  assign n3015 = ~n3013 & n3014;
  assign n3016 = ~n3012 & ~n3013;
  assign n3017 = ~pi933  & ~n3016;
  assign n3018 = ~n3015 & ~n3017;
  assign n3019 = ~pi934  & pi935 ;
  assign n3020 = pi934  & ~pi935 ;
  assign n3021 = pi936  & ~n3019;
  assign n3022 = ~n3020 & n3021;
  assign n3023 = ~n3019 & ~n3020;
  assign n3024 = ~pi936  & ~n3023;
  assign n3025 = ~n3022 & ~n3024;
  assign n3026 = ~n3018 & n3025;
  assign n3027 = n3018 & ~n3025;
  assign n3028 = ~n3026 & ~n3027;
  assign n3029 = ~n3011 & ~n3028;
  assign n3030 = pi940  & pi941 ;
  assign n3031 = pi942  & ~n3006;
  assign n3032 = ~n3030 & ~n3031;
  assign n3033 = pi937  & pi938 ;
  assign n3034 = pi939  & ~n2999;
  assign n3035 = ~n3033 & ~n3034;
  assign n3036 = n3032 & ~n3035;
  assign n3037 = ~n3032 & n3035;
  assign n3038 = ~n3036 & ~n3037;
  assign n3039 = n3029 & ~n3038;
  assign n3040 = ~n3001 & ~n3008;
  assign n3041 = n3038 & n3040;
  assign n3042 = ~n3038 & ~n3040;
  assign n3043 = ~n3029 & ~n3041;
  assign n3044 = ~n3042 & n3043;
  assign n3045 = pi934  & pi935 ;
  assign n3046 = pi936  & ~n3023;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = pi931  & pi932 ;
  assign n3049 = pi933  & ~n3016;
  assign n3050 = ~n3048 & ~n3049;
  assign n3051 = ~n3047 & ~n3050;
  assign n3052 = ~n3028 & n3051;
  assign n3053 = ~n3018 & ~n3025;
  assign n3054 = n3047 & n3050;
  assign n3055 = ~n3051 & ~n3054;
  assign n3056 = n3053 & n3055;
  assign n3057 = ~n3053 & ~n3055;
  assign n3058 = ~n3052 & ~n3056;
  assign n3059 = ~n3057 & n3058;
  assign n3060 = ~n3044 & n3059;
  assign n3061 = ~n3039 & ~n3060;
  assign n3062 = ~n3032 & n3040;
  assign n3063 = n3035 & ~n3062;
  assign n3064 = n3032 & ~n3040;
  assign n3065 = ~n3063 & ~n3064;
  assign n3066 = ~n3061 & n3065;
  assign n3067 = n3061 & ~n3065;
  assign n3068 = ~n3066 & ~n3067;
  assign n3069 = n3053 & ~n3054;
  assign n3070 = ~n3051 & ~n3069;
  assign n3071 = n3068 & ~n3070;
  assign n3072 = ~n3068 & n3070;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = n2994 & ~n3073;
  assign n3075 = ~n2994 & n3073;
  assign n3076 = n3011 & n3028;
  assign n3077 = ~n3029 & ~n3076;
  assign n3078 = n2932 & n2949;
  assign n3079 = ~n2950 & ~n3078;
  assign n3080 = n3077 & n3079;
  assign n3081 = ~n3039 & ~n3044;
  assign n3082 = n3059 & n3081;
  assign n3083 = ~n3059 & ~n3081;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = n3080 & n3084;
  assign n3086 = ~n3080 & ~n3084;
  assign n3087 = ~n2966 & ~n2967;
  assign n3088 = ~n2980 & n3087;
  assign n3089 = n2980 & ~n3087;
  assign n3090 = ~n3088 & ~n3089;
  assign n3091 = ~n3086 & n3090;
  assign n3092 = ~n3085 & ~n3091;
  assign n3093 = ~n3075 & n3092;
  assign n3094 = ~n3074 & ~n3093;
  assign n3095 = ~n3067 & ~n3070;
  assign n3096 = ~n3066 & ~n3095;
  assign n3097 = ~n3094 & n3096;
  assign n3098 = n3094 & ~n3096;
  assign n3099 = ~n2986 & n2991;
  assign n3100 = ~n2985 & ~n3099;
  assign n3101 = ~n3098 & n3100;
  assign n3102 = ~n3097 & ~n3101;
  assign n3103 = ~n3097 & ~n3098;
  assign n3104 = n3100 & n3103;
  assign n3105 = ~n3100 & ~n3103;
  assign n3106 = ~n3104 & ~n3105;
  assign n3107 = ~n2910 & ~n2911;
  assign n3108 = n2913 & n3107;
  assign n3109 = ~n2913 & ~n3107;
  assign n3110 = ~n3108 & ~n3109;
  assign n3111 = ~n3106 & ~n3110;
  assign n3112 = n3106 & n3110;
  assign n3113 = ~n2887 & ~n2888;
  assign n3114 = ~n2905 & n3113;
  assign n3115 = n2905 & ~n3113;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = ~n3074 & ~n3075;
  assign n3118 = ~n3092 & n3117;
  assign n3119 = n3092 & ~n3117;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = ~n3116 & ~n3120;
  assign n3122 = n3116 & n3120;
  assign n3123 = ~n3077 & ~n3079;
  assign n3124 = ~n3080 & ~n3123;
  assign n3125 = ~n2890 & ~n2892;
  assign n3126 = ~n2893 & ~n3125;
  assign n3127 = n3124 & n3126;
  assign n3128 = ~n3085 & ~n3086;
  assign n3129 = ~n3090 & n3128;
  assign n3130 = n3090 & ~n3128;
  assign n3131 = ~n3129 & ~n3130;
  assign n3132 = n3127 & ~n3131;
  assign n3133 = ~n3127 & n3131;
  assign n3134 = ~n2898 & ~n2899;
  assign n3135 = ~n2903 & n3134;
  assign n3136 = n2903 & ~n3134;
  assign n3137 = ~n3135 & ~n3136;
  assign n3138 = ~n3133 & ~n3137;
  assign n3139 = ~n3132 & ~n3138;
  assign n3140 = ~n3122 & n3139;
  assign n3141 = ~n3121 & ~n3140;
  assign n3142 = ~n3112 & n3141;
  assign n3143 = ~n3111 & ~n3142;
  assign n3144 = ~n3102 & n3143;
  assign n3145 = n3102 & ~n3143;
  assign n3146 = ~n3144 & ~n3145;
  assign n3147 = n2915 & n3146;
  assign n3148 = ~n2915 & ~n3146;
  assign n3149 = ~n3147 & ~n3148;
  assign n3150 = ~n2728 & ~n3149;
  assign n3151 = n2728 & n3149;
  assign n3152 = ~n3111 & ~n3112;
  assign n3153 = ~n3141 & n3152;
  assign n3154 = n3141 & ~n3152;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = ~n2690 & ~n2691;
  assign n3157 = ~n2720 & n3156;
  assign n3158 = n2720 & ~n3156;
  assign n3159 = ~n3157 & ~n3158;
  assign n3160 = ~n3155 & ~n3159;
  assign n3161 = n3155 & n3159;
  assign n3162 = ~n2700 & ~n2701;
  assign n3163 = ~n2718 & n3162;
  assign n3164 = n2718 & ~n3162;
  assign n3165 = ~n3163 & ~n3164;
  assign n3166 = ~n3121 & ~n3122;
  assign n3167 = ~n3139 & n3166;
  assign n3168 = n3139 & ~n3166;
  assign n3169 = ~n3167 & ~n3168;
  assign n3170 = ~n3165 & ~n3169;
  assign n3171 = n3165 & n3169;
  assign n3172 = n3124 & ~n3126;
  assign n3173 = ~n3124 & n3126;
  assign n3174 = ~n3172 & ~n3173;
  assign n3175 = n2703 & ~n2705;
  assign n3176 = ~n2703 & n2705;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = ~n3174 & ~n3177;
  assign n3179 = ~n3132 & ~n3133;
  assign n3180 = n3137 & n3179;
  assign n3181 = ~n3137 & ~n3179;
  assign n3182 = ~n3180 & ~n3181;
  assign n3183 = n3178 & ~n3182;
  assign n3184 = ~n3178 & n3182;
  assign n3185 = ~n2711 & ~n2712;
  assign n3186 = n2716 & n3185;
  assign n3187 = ~n2716 & ~n3185;
  assign n3188 = ~n3186 & ~n3187;
  assign n3189 = ~n3184 & ~n3188;
  assign n3190 = ~n3183 & ~n3189;
  assign n3191 = ~n3171 & n3190;
  assign n3192 = ~n3170 & ~n3191;
  assign n3193 = ~n3161 & n3192;
  assign n3194 = ~n3160 & ~n3193;
  assign n3195 = ~n3151 & n3194;
  assign n3196 = ~n3150 & ~n3195;
  assign n3197 = ~n2915 & ~n3145;
  assign n3198 = ~n3144 & ~n3197;
  assign n3199 = ~n3196 & ~n3198;
  assign n3200 = n3196 & n3198;
  assign n3201 = ~n2494 & ~n2724;
  assign n3202 = ~n2723 & ~n3201;
  assign n3203 = ~n3200 & ~n3202;
  assign n3204 = ~n3199 & ~n3203;
  assign n3205 = ~n2307 & ~n3204;
  assign n3206 = ~n2243 & ~n2244;
  assign n3207 = ~n2300 & n3206;
  assign n3208 = n2300 & ~n3206;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = ~n3196 & n3198;
  assign n3211 = n3196 & ~n3198;
  assign n3212 = ~n3210 & ~n3211;
  assign n3213 = n3202 & n3212;
  assign n3214 = ~n3202 & ~n3212;
  assign n3215 = ~n3213 & ~n3214;
  assign n3216 = ~n3209 & ~n3215;
  assign n3217 = n3209 & n3215;
  assign n3218 = ~n3150 & ~n3151;
  assign n3219 = ~n3194 & n3218;
  assign n3220 = n3194 & ~n3218;
  assign n3221 = ~n3219 & ~n3220;
  assign n3222 = ~n2255 & ~n2256;
  assign n3223 = ~n2298 & n3222;
  assign n3224 = n2298 & ~n3222;
  assign n3225 = ~n3223 & ~n3224;
  assign n3226 = ~n3221 & ~n3225;
  assign n3227 = n3221 & n3225;
  assign n3228 = ~n2265 & ~n2266;
  assign n3229 = n2296 & n3228;
  assign n3230 = ~n2296 & ~n3228;
  assign n3231 = ~n3229 & ~n3230;
  assign n3232 = ~n3160 & ~n3161;
  assign n3233 = n3192 & n3232;
  assign n3234 = ~n3192 & ~n3232;
  assign n3235 = ~n3233 & ~n3234;
  assign n3236 = ~n3231 & ~n3235;
  assign n3237 = n3231 & n3235;
  assign n3238 = ~n3170 & ~n3171;
  assign n3239 = ~n3190 & n3238;
  assign n3240 = n3190 & ~n3238;
  assign n3241 = ~n3239 & ~n3240;
  assign n3242 = ~n2275 & ~n2276;
  assign n3243 = ~n2294 & n3242;
  assign n3244 = n2294 & ~n3242;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = ~n3241 & ~n3245;
  assign n3247 = n3241 & n3245;
  assign n3248 = n3174 & n3177;
  assign n3249 = ~n3178 & ~n3248;
  assign n3250 = n2279 & ~n2281;
  assign n3251 = ~n2282 & ~n3250;
  assign n3252 = n3249 & n3251;
  assign n3253 = ~n2287 & ~n2288;
  assign n3254 = n2292 & n3253;
  assign n3255 = ~n2292 & ~n3253;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = n3252 & ~n3256;
  assign n3258 = ~n3252 & n3256;
  assign n3259 = ~n3183 & ~n3184;
  assign n3260 = n3188 & n3259;
  assign n3261 = ~n3188 & ~n3259;
  assign n3262 = ~n3260 & ~n3261;
  assign n3263 = ~n3258 & ~n3262;
  assign n3264 = ~n3257 & ~n3263;
  assign n3265 = ~n3247 & n3264;
  assign n3266 = ~n3246 & ~n3265;
  assign n3267 = ~n3237 & ~n3266;
  assign n3268 = ~n3236 & ~n3267;
  assign n3269 = ~n3227 & ~n3268;
  assign n3270 = ~n3226 & ~n3269;
  assign n3271 = ~n3217 & n3270;
  assign n3272 = ~n3216 & ~n3271;
  assign n3273 = ~n3205 & ~n3272;
  assign n3274 = n2305 & n3273;
  assign n3275 = ~pi85  & pi86 ;
  assign n3276 = pi85  & ~pi86 ;
  assign n3277 = pi87  & ~n3275;
  assign n3278 = ~n3276 & n3277;
  assign n3279 = ~n3275 & ~n3276;
  assign n3280 = ~pi87  & ~n3279;
  assign n3281 = ~n3278 & ~n3280;
  assign n3282 = ~pi88  & pi89 ;
  assign n3283 = pi88  & ~pi89 ;
  assign n3284 = pi90  & ~n3282;
  assign n3285 = ~n3283 & n3284;
  assign n3286 = ~n3282 & ~n3283;
  assign n3287 = ~pi90  & ~n3286;
  assign n3288 = ~n3285 & ~n3287;
  assign n3289 = ~n3281 & n3288;
  assign n3290 = n3281 & ~n3288;
  assign n3291 = ~n3289 & ~n3290;
  assign n3292 = ~pi79  & pi80 ;
  assign n3293 = pi79  & ~pi80 ;
  assign n3294 = pi81  & ~n3292;
  assign n3295 = ~n3293 & n3294;
  assign n3296 = ~n3292 & ~n3293;
  assign n3297 = ~pi81  & ~n3296;
  assign n3298 = ~n3295 & ~n3297;
  assign n3299 = ~pi82  & pi83 ;
  assign n3300 = pi82  & ~pi83 ;
  assign n3301 = pi84  & ~n3299;
  assign n3302 = ~n3300 & n3301;
  assign n3303 = ~n3299 & ~n3300;
  assign n3304 = ~pi84  & ~n3303;
  assign n3305 = ~n3302 & ~n3304;
  assign n3306 = ~n3298 & n3305;
  assign n3307 = n3298 & ~n3305;
  assign n3308 = ~n3306 & ~n3307;
  assign n3309 = ~n3291 & ~n3308;
  assign n3310 = pi88  & pi89 ;
  assign n3311 = pi90  & ~n3286;
  assign n3312 = ~n3310 & ~n3311;
  assign n3313 = pi85  & pi86 ;
  assign n3314 = pi87  & ~n3279;
  assign n3315 = ~n3313 & ~n3314;
  assign n3316 = ~n3312 & ~n3315;
  assign n3317 = ~n3291 & n3316;
  assign n3318 = ~n3281 & ~n3288;
  assign n3319 = n3312 & n3315;
  assign n3320 = ~n3316 & ~n3319;
  assign n3321 = n3318 & n3320;
  assign n3322 = ~n3318 & ~n3320;
  assign n3323 = ~n3317 & ~n3321;
  assign n3324 = ~n3322 & n3323;
  assign n3325 = n3309 & n3324;
  assign n3326 = ~n3309 & ~n3324;
  assign n3327 = pi82  & pi83 ;
  assign n3328 = pi84  & ~n3303;
  assign n3329 = ~n3327 & ~n3328;
  assign n3330 = pi79  & pi80 ;
  assign n3331 = pi81  & ~n3296;
  assign n3332 = ~n3330 & ~n3331;
  assign n3333 = ~n3329 & n3332;
  assign n3334 = n3329 & ~n3332;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = ~n3298 & ~n3305;
  assign n3337 = n3335 & n3336;
  assign n3338 = ~n3335 & ~n3336;
  assign n3339 = ~n3337 & ~n3338;
  assign n3340 = ~n3326 & ~n3339;
  assign n3341 = ~n3325 & ~n3340;
  assign n3342 = n3318 & ~n3319;
  assign n3343 = ~n3316 & ~n3342;
  assign n3344 = ~n3341 & ~n3343;
  assign n3345 = n3341 & n3343;
  assign n3346 = ~n3344 & ~n3345;
  assign n3347 = ~n3329 & n3336;
  assign n3348 = n3332 & ~n3347;
  assign n3349 = n3329 & ~n3336;
  assign n3350 = ~n3348 & ~n3349;
  assign n3351 = ~n3346 & n3350;
  assign n3352 = n3346 & ~n3350;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = ~pi97  & pi98 ;
  assign n3355 = pi97  & ~pi98 ;
  assign n3356 = pi99  & ~n3354;
  assign n3357 = ~n3355 & n3356;
  assign n3358 = ~n3354 & ~n3355;
  assign n3359 = ~pi99  & ~n3358;
  assign n3360 = ~n3357 & ~n3359;
  assign n3361 = ~pi100  & pi101 ;
  assign n3362 = pi100  & ~pi101 ;
  assign n3363 = pi102  & ~n3361;
  assign n3364 = ~n3362 & n3363;
  assign n3365 = ~n3361 & ~n3362;
  assign n3366 = ~pi102  & ~n3365;
  assign n3367 = ~n3364 & ~n3366;
  assign n3368 = ~n3360 & n3367;
  assign n3369 = n3360 & ~n3367;
  assign n3370 = ~n3368 & ~n3369;
  assign n3371 = ~pi91  & pi92 ;
  assign n3372 = pi91  & ~pi92 ;
  assign n3373 = pi93  & ~n3371;
  assign n3374 = ~n3372 & n3373;
  assign n3375 = ~n3371 & ~n3372;
  assign n3376 = ~pi93  & ~n3375;
  assign n3377 = ~n3374 & ~n3376;
  assign n3378 = ~pi94  & pi95 ;
  assign n3379 = pi94  & ~pi95 ;
  assign n3380 = pi96  & ~n3378;
  assign n3381 = ~n3379 & n3380;
  assign n3382 = ~n3378 & ~n3379;
  assign n3383 = ~pi96  & ~n3382;
  assign n3384 = ~n3381 & ~n3383;
  assign n3385 = ~n3377 & n3384;
  assign n3386 = n3377 & ~n3384;
  assign n3387 = ~n3385 & ~n3386;
  assign n3388 = ~n3370 & ~n3387;
  assign n3389 = pi100  & pi101 ;
  assign n3390 = pi102  & ~n3365;
  assign n3391 = ~n3389 & ~n3390;
  assign n3392 = pi97  & pi98 ;
  assign n3393 = pi99  & ~n3358;
  assign n3394 = ~n3392 & ~n3393;
  assign n3395 = n3391 & ~n3394;
  assign n3396 = ~n3391 & n3394;
  assign n3397 = ~n3395 & ~n3396;
  assign n3398 = n3388 & ~n3397;
  assign n3399 = ~n3360 & ~n3367;
  assign n3400 = n3397 & n3399;
  assign n3401 = ~n3397 & ~n3399;
  assign n3402 = ~n3388 & ~n3400;
  assign n3403 = ~n3401 & n3402;
  assign n3404 = pi94  & pi95 ;
  assign n3405 = pi96  & ~n3382;
  assign n3406 = ~n3404 & ~n3405;
  assign n3407 = pi91  & pi92 ;
  assign n3408 = pi93  & ~n3375;
  assign n3409 = ~n3407 & ~n3408;
  assign n3410 = ~n3406 & ~n3409;
  assign n3411 = ~n3387 & n3410;
  assign n3412 = ~n3377 & ~n3384;
  assign n3413 = n3406 & n3409;
  assign n3414 = ~n3410 & ~n3413;
  assign n3415 = n3412 & n3414;
  assign n3416 = ~n3412 & ~n3414;
  assign n3417 = ~n3411 & ~n3415;
  assign n3418 = ~n3416 & n3417;
  assign n3419 = ~n3403 & n3418;
  assign n3420 = ~n3398 & ~n3419;
  assign n3421 = ~n3391 & n3399;
  assign n3422 = n3394 & ~n3421;
  assign n3423 = n3391 & ~n3399;
  assign n3424 = ~n3422 & ~n3423;
  assign n3425 = ~n3420 & n3424;
  assign n3426 = n3420 & ~n3424;
  assign n3427 = ~n3425 & ~n3426;
  assign n3428 = n3412 & ~n3413;
  assign n3429 = ~n3410 & ~n3428;
  assign n3430 = n3427 & ~n3429;
  assign n3431 = ~n3427 & n3429;
  assign n3432 = ~n3430 & ~n3431;
  assign n3433 = n3353 & ~n3432;
  assign n3434 = ~n3353 & n3432;
  assign n3435 = n3370 & n3387;
  assign n3436 = ~n3388 & ~n3435;
  assign n3437 = n3291 & n3308;
  assign n3438 = ~n3309 & ~n3437;
  assign n3439 = n3436 & n3438;
  assign n3440 = ~n3398 & ~n3403;
  assign n3441 = n3418 & n3440;
  assign n3442 = ~n3418 & ~n3440;
  assign n3443 = ~n3441 & ~n3442;
  assign n3444 = n3439 & n3443;
  assign n3445 = ~n3439 & ~n3443;
  assign n3446 = ~n3325 & ~n3326;
  assign n3447 = ~n3339 & n3446;
  assign n3448 = n3339 & ~n3446;
  assign n3449 = ~n3447 & ~n3448;
  assign n3450 = ~n3445 & n3449;
  assign n3451 = ~n3444 & ~n3450;
  assign n3452 = ~n3434 & n3451;
  assign n3453 = ~n3433 & ~n3452;
  assign n3454 = ~n3426 & ~n3429;
  assign n3455 = ~n3425 & ~n3454;
  assign n3456 = ~n3453 & n3455;
  assign n3457 = n3453 & ~n3455;
  assign n3458 = ~n3345 & n3350;
  assign n3459 = ~n3344 & ~n3458;
  assign n3460 = ~n3457 & n3459;
  assign n3461 = ~n3456 & ~n3460;
  assign n3462 = ~pi109  & pi110 ;
  assign n3463 = pi109  & ~pi110 ;
  assign n3464 = pi111  & ~n3462;
  assign n3465 = ~n3463 & n3464;
  assign n3466 = ~n3462 & ~n3463;
  assign n3467 = ~pi111  & ~n3466;
  assign n3468 = ~n3465 & ~n3467;
  assign n3469 = ~pi112  & pi113 ;
  assign n3470 = pi112  & ~pi113 ;
  assign n3471 = pi114  & ~n3469;
  assign n3472 = ~n3470 & n3471;
  assign n3473 = ~n3469 & ~n3470;
  assign n3474 = ~pi114  & ~n3473;
  assign n3475 = ~n3472 & ~n3474;
  assign n3476 = ~n3468 & n3475;
  assign n3477 = n3468 & ~n3475;
  assign n3478 = ~n3476 & ~n3477;
  assign n3479 = ~pi103  & pi104 ;
  assign n3480 = pi103  & ~pi104 ;
  assign n3481 = pi105  & ~n3479;
  assign n3482 = ~n3480 & n3481;
  assign n3483 = ~n3479 & ~n3480;
  assign n3484 = ~pi105  & ~n3483;
  assign n3485 = ~n3482 & ~n3484;
  assign n3486 = ~pi106  & pi107 ;
  assign n3487 = pi106  & ~pi107 ;
  assign n3488 = pi108  & ~n3486;
  assign n3489 = ~n3487 & n3488;
  assign n3490 = ~n3486 & ~n3487;
  assign n3491 = ~pi108  & ~n3490;
  assign n3492 = ~n3489 & ~n3491;
  assign n3493 = ~n3485 & n3492;
  assign n3494 = n3485 & ~n3492;
  assign n3495 = ~n3493 & ~n3494;
  assign n3496 = ~n3478 & ~n3495;
  assign n3497 = pi112  & pi113 ;
  assign n3498 = pi114  & ~n3473;
  assign n3499 = ~n3497 & ~n3498;
  assign n3500 = pi109  & pi110 ;
  assign n3501 = pi111  & ~n3466;
  assign n3502 = ~n3500 & ~n3501;
  assign n3503 = ~n3499 & ~n3502;
  assign n3504 = ~n3478 & n3503;
  assign n3505 = ~n3468 & ~n3475;
  assign n3506 = n3499 & n3502;
  assign n3507 = ~n3503 & ~n3506;
  assign n3508 = n3505 & n3507;
  assign n3509 = ~n3505 & ~n3507;
  assign n3510 = ~n3504 & ~n3508;
  assign n3511 = ~n3509 & n3510;
  assign n3512 = n3496 & n3511;
  assign n3513 = ~n3496 & ~n3511;
  assign n3514 = pi106  & pi107 ;
  assign n3515 = pi108  & ~n3490;
  assign n3516 = ~n3514 & ~n3515;
  assign n3517 = pi103  & pi104 ;
  assign n3518 = pi105  & ~n3483;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520 = ~n3516 & n3519;
  assign n3521 = n3516 & ~n3519;
  assign n3522 = ~n3520 & ~n3521;
  assign n3523 = ~n3485 & ~n3492;
  assign n3524 = n3522 & n3523;
  assign n3525 = ~n3522 & ~n3523;
  assign n3526 = ~n3524 & ~n3525;
  assign n3527 = ~n3513 & ~n3526;
  assign n3528 = ~n3512 & ~n3527;
  assign n3529 = n3505 & ~n3506;
  assign n3530 = ~n3503 & ~n3529;
  assign n3531 = ~n3528 & ~n3530;
  assign n3532 = n3528 & n3530;
  assign n3533 = ~n3531 & ~n3532;
  assign n3534 = ~n3516 & n3523;
  assign n3535 = n3519 & ~n3534;
  assign n3536 = n3516 & ~n3523;
  assign n3537 = ~n3535 & ~n3536;
  assign n3538 = ~n3533 & n3537;
  assign n3539 = n3533 & ~n3537;
  assign n3540 = ~n3538 & ~n3539;
  assign n3541 = ~pi121  & pi122 ;
  assign n3542 = pi121  & ~pi122 ;
  assign n3543 = pi123  & ~n3541;
  assign n3544 = ~n3542 & n3543;
  assign n3545 = ~n3541 & ~n3542;
  assign n3546 = ~pi123  & ~n3545;
  assign n3547 = ~n3544 & ~n3546;
  assign n3548 = ~pi124  & pi125 ;
  assign n3549 = pi124  & ~pi125 ;
  assign n3550 = pi126  & ~n3548;
  assign n3551 = ~n3549 & n3550;
  assign n3552 = ~n3548 & ~n3549;
  assign n3553 = ~pi126  & ~n3552;
  assign n3554 = ~n3551 & ~n3553;
  assign n3555 = ~n3547 & n3554;
  assign n3556 = n3547 & ~n3554;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = ~pi115  & pi116 ;
  assign n3559 = pi115  & ~pi116 ;
  assign n3560 = pi117  & ~n3558;
  assign n3561 = ~n3559 & n3560;
  assign n3562 = ~n3558 & ~n3559;
  assign n3563 = ~pi117  & ~n3562;
  assign n3564 = ~n3561 & ~n3563;
  assign n3565 = ~pi118  & pi119 ;
  assign n3566 = pi118  & ~pi119 ;
  assign n3567 = pi120  & ~n3565;
  assign n3568 = ~n3566 & n3567;
  assign n3569 = ~n3565 & ~n3566;
  assign n3570 = ~pi120  & ~n3569;
  assign n3571 = ~n3568 & ~n3570;
  assign n3572 = ~n3564 & n3571;
  assign n3573 = n3564 & ~n3571;
  assign n3574 = ~n3572 & ~n3573;
  assign n3575 = ~n3557 & ~n3574;
  assign n3576 = pi124  & pi125 ;
  assign n3577 = pi126  & ~n3552;
  assign n3578 = ~n3576 & ~n3577;
  assign n3579 = pi121  & pi122 ;
  assign n3580 = pi123  & ~n3545;
  assign n3581 = ~n3579 & ~n3580;
  assign n3582 = n3578 & ~n3581;
  assign n3583 = ~n3578 & n3581;
  assign n3584 = ~n3582 & ~n3583;
  assign n3585 = n3575 & ~n3584;
  assign n3586 = ~n3547 & ~n3554;
  assign n3587 = n3584 & n3586;
  assign n3588 = ~n3584 & ~n3586;
  assign n3589 = ~n3575 & ~n3587;
  assign n3590 = ~n3588 & n3589;
  assign n3591 = pi118  & pi119 ;
  assign n3592 = pi120  & ~n3569;
  assign n3593 = ~n3591 & ~n3592;
  assign n3594 = pi115  & pi116 ;
  assign n3595 = pi117  & ~n3562;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = ~n3593 & ~n3596;
  assign n3598 = ~n3574 & n3597;
  assign n3599 = ~n3564 & ~n3571;
  assign n3600 = n3593 & n3596;
  assign n3601 = ~n3597 & ~n3600;
  assign n3602 = n3599 & n3601;
  assign n3603 = ~n3599 & ~n3601;
  assign n3604 = ~n3598 & ~n3602;
  assign n3605 = ~n3603 & n3604;
  assign n3606 = ~n3590 & n3605;
  assign n3607 = ~n3585 & ~n3606;
  assign n3608 = ~n3578 & n3586;
  assign n3609 = n3581 & ~n3608;
  assign n3610 = n3578 & ~n3586;
  assign n3611 = ~n3609 & ~n3610;
  assign n3612 = ~n3607 & n3611;
  assign n3613 = n3607 & ~n3611;
  assign n3614 = ~n3612 & ~n3613;
  assign n3615 = n3599 & ~n3600;
  assign n3616 = ~n3597 & ~n3615;
  assign n3617 = n3614 & ~n3616;
  assign n3618 = ~n3614 & n3616;
  assign n3619 = ~n3617 & ~n3618;
  assign n3620 = n3540 & ~n3619;
  assign n3621 = ~n3540 & n3619;
  assign n3622 = n3557 & n3574;
  assign n3623 = ~n3575 & ~n3622;
  assign n3624 = n3478 & n3495;
  assign n3625 = ~n3496 & ~n3624;
  assign n3626 = n3623 & n3625;
  assign n3627 = ~n3585 & ~n3590;
  assign n3628 = n3605 & n3627;
  assign n3629 = ~n3605 & ~n3627;
  assign n3630 = ~n3628 & ~n3629;
  assign n3631 = n3626 & n3630;
  assign n3632 = ~n3626 & ~n3630;
  assign n3633 = ~n3512 & ~n3513;
  assign n3634 = ~n3526 & n3633;
  assign n3635 = n3526 & ~n3633;
  assign n3636 = ~n3634 & ~n3635;
  assign n3637 = ~n3632 & n3636;
  assign n3638 = ~n3631 & ~n3637;
  assign n3639 = ~n3621 & n3638;
  assign n3640 = ~n3620 & ~n3639;
  assign n3641 = ~n3613 & ~n3616;
  assign n3642 = ~n3612 & ~n3641;
  assign n3643 = ~n3640 & n3642;
  assign n3644 = n3640 & ~n3642;
  assign n3645 = ~n3532 & n3537;
  assign n3646 = ~n3531 & ~n3645;
  assign n3647 = ~n3644 & n3646;
  assign n3648 = ~n3643 & ~n3647;
  assign n3649 = ~n3643 & ~n3644;
  assign n3650 = n3646 & n3649;
  assign n3651 = ~n3646 & ~n3649;
  assign n3652 = ~n3650 & ~n3651;
  assign n3653 = ~n3456 & ~n3457;
  assign n3654 = n3459 & n3653;
  assign n3655 = ~n3459 & ~n3653;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = ~n3652 & ~n3656;
  assign n3658 = n3652 & n3656;
  assign n3659 = ~n3433 & ~n3434;
  assign n3660 = ~n3451 & n3659;
  assign n3661 = n3451 & ~n3659;
  assign n3662 = ~n3660 & ~n3661;
  assign n3663 = ~n3620 & ~n3621;
  assign n3664 = ~n3638 & n3663;
  assign n3665 = n3638 & ~n3663;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = ~n3662 & ~n3666;
  assign n3668 = n3662 & n3666;
  assign n3669 = ~n3623 & ~n3625;
  assign n3670 = ~n3626 & ~n3669;
  assign n3671 = ~n3436 & ~n3438;
  assign n3672 = ~n3439 & ~n3671;
  assign n3673 = n3670 & n3672;
  assign n3674 = ~n3631 & ~n3632;
  assign n3675 = ~n3636 & n3674;
  assign n3676 = n3636 & ~n3674;
  assign n3677 = ~n3675 & ~n3676;
  assign n3678 = n3673 & ~n3677;
  assign n3679 = ~n3673 & n3677;
  assign n3680 = ~n3444 & ~n3445;
  assign n3681 = ~n3449 & n3680;
  assign n3682 = n3449 & ~n3680;
  assign n3683 = ~n3681 & ~n3682;
  assign n3684 = ~n3679 & ~n3683;
  assign n3685 = ~n3678 & ~n3684;
  assign n3686 = ~n3668 & n3685;
  assign n3687 = ~n3667 & ~n3686;
  assign n3688 = ~n3658 & n3687;
  assign n3689 = ~n3657 & ~n3688;
  assign n3690 = ~n3648 & n3689;
  assign n3691 = n3648 & ~n3689;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = n3461 & n3692;
  assign n3694 = ~n3461 & ~n3692;
  assign n3695 = ~n3693 & ~n3694;
  assign n3696 = ~pi133  & pi134 ;
  assign n3697 = pi133  & ~pi134 ;
  assign n3698 = pi135  & ~n3696;
  assign n3699 = ~n3697 & n3698;
  assign n3700 = ~n3696 & ~n3697;
  assign n3701 = ~pi135  & ~n3700;
  assign n3702 = ~n3699 & ~n3701;
  assign n3703 = ~pi136  & pi137 ;
  assign n3704 = pi136  & ~pi137 ;
  assign n3705 = pi138  & ~n3703;
  assign n3706 = ~n3704 & n3705;
  assign n3707 = ~n3703 & ~n3704;
  assign n3708 = ~pi138  & ~n3707;
  assign n3709 = ~n3706 & ~n3708;
  assign n3710 = ~n3702 & n3709;
  assign n3711 = n3702 & ~n3709;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = ~pi127  & pi128 ;
  assign n3714 = pi127  & ~pi128 ;
  assign n3715 = pi129  & ~n3713;
  assign n3716 = ~n3714 & n3715;
  assign n3717 = ~n3713 & ~n3714;
  assign n3718 = ~pi129  & ~n3717;
  assign n3719 = ~n3716 & ~n3718;
  assign n3720 = ~pi130  & pi131 ;
  assign n3721 = pi130  & ~pi131 ;
  assign n3722 = pi132  & ~n3720;
  assign n3723 = ~n3721 & n3722;
  assign n3724 = ~n3720 & ~n3721;
  assign n3725 = ~pi132  & ~n3724;
  assign n3726 = ~n3723 & ~n3725;
  assign n3727 = ~n3719 & n3726;
  assign n3728 = n3719 & ~n3726;
  assign n3729 = ~n3727 & ~n3728;
  assign n3730 = ~n3712 & ~n3729;
  assign n3731 = pi136  & pi137 ;
  assign n3732 = pi138  & ~n3707;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = pi133  & pi134 ;
  assign n3735 = pi135  & ~n3700;
  assign n3736 = ~n3734 & ~n3735;
  assign n3737 = ~n3733 & ~n3736;
  assign n3738 = ~n3712 & n3737;
  assign n3739 = ~n3702 & ~n3709;
  assign n3740 = n3733 & n3736;
  assign n3741 = ~n3737 & ~n3740;
  assign n3742 = n3739 & n3741;
  assign n3743 = ~n3739 & ~n3741;
  assign n3744 = ~n3738 & ~n3742;
  assign n3745 = ~n3743 & n3744;
  assign n3746 = n3730 & n3745;
  assign n3747 = ~n3730 & ~n3745;
  assign n3748 = pi130  & pi131 ;
  assign n3749 = pi132  & ~n3724;
  assign n3750 = ~n3748 & ~n3749;
  assign n3751 = pi127  & pi128 ;
  assign n3752 = pi129  & ~n3717;
  assign n3753 = ~n3751 & ~n3752;
  assign n3754 = ~n3750 & n3753;
  assign n3755 = n3750 & ~n3753;
  assign n3756 = ~n3754 & ~n3755;
  assign n3757 = ~n3719 & ~n3726;
  assign n3758 = n3756 & n3757;
  assign n3759 = ~n3756 & ~n3757;
  assign n3760 = ~n3758 & ~n3759;
  assign n3761 = ~n3747 & ~n3760;
  assign n3762 = ~n3746 & ~n3761;
  assign n3763 = n3739 & ~n3740;
  assign n3764 = ~n3737 & ~n3763;
  assign n3765 = ~n3762 & ~n3764;
  assign n3766 = n3762 & n3764;
  assign n3767 = ~n3765 & ~n3766;
  assign n3768 = ~n3750 & n3757;
  assign n3769 = n3753 & ~n3768;
  assign n3770 = n3750 & ~n3757;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = ~n3767 & n3771;
  assign n3773 = n3767 & ~n3771;
  assign n3774 = ~n3772 & ~n3773;
  assign n3775 = ~pi145  & pi146 ;
  assign n3776 = pi145  & ~pi146 ;
  assign n3777 = pi147  & ~n3775;
  assign n3778 = ~n3776 & n3777;
  assign n3779 = ~n3775 & ~n3776;
  assign n3780 = ~pi147  & ~n3779;
  assign n3781 = ~n3778 & ~n3780;
  assign n3782 = ~pi148  & pi149 ;
  assign n3783 = pi148  & ~pi149 ;
  assign n3784 = pi150  & ~n3782;
  assign n3785 = ~n3783 & n3784;
  assign n3786 = ~n3782 & ~n3783;
  assign n3787 = ~pi150  & ~n3786;
  assign n3788 = ~n3785 & ~n3787;
  assign n3789 = ~n3781 & n3788;
  assign n3790 = n3781 & ~n3788;
  assign n3791 = ~n3789 & ~n3790;
  assign n3792 = ~pi139  & pi140 ;
  assign n3793 = pi139  & ~pi140 ;
  assign n3794 = pi141  & ~n3792;
  assign n3795 = ~n3793 & n3794;
  assign n3796 = ~n3792 & ~n3793;
  assign n3797 = ~pi141  & ~n3796;
  assign n3798 = ~n3795 & ~n3797;
  assign n3799 = ~pi142  & pi143 ;
  assign n3800 = pi142  & ~pi143 ;
  assign n3801 = pi144  & ~n3799;
  assign n3802 = ~n3800 & n3801;
  assign n3803 = ~n3799 & ~n3800;
  assign n3804 = ~pi144  & ~n3803;
  assign n3805 = ~n3802 & ~n3804;
  assign n3806 = ~n3798 & n3805;
  assign n3807 = n3798 & ~n3805;
  assign n3808 = ~n3806 & ~n3807;
  assign n3809 = ~n3791 & ~n3808;
  assign n3810 = pi148  & pi149 ;
  assign n3811 = pi150  & ~n3786;
  assign n3812 = ~n3810 & ~n3811;
  assign n3813 = pi145  & pi146 ;
  assign n3814 = pi147  & ~n3779;
  assign n3815 = ~n3813 & ~n3814;
  assign n3816 = n3812 & ~n3815;
  assign n3817 = ~n3812 & n3815;
  assign n3818 = ~n3816 & ~n3817;
  assign n3819 = n3809 & ~n3818;
  assign n3820 = ~n3781 & ~n3788;
  assign n3821 = n3818 & n3820;
  assign n3822 = ~n3818 & ~n3820;
  assign n3823 = ~n3809 & ~n3821;
  assign n3824 = ~n3822 & n3823;
  assign n3825 = pi142  & pi143 ;
  assign n3826 = pi144  & ~n3803;
  assign n3827 = ~n3825 & ~n3826;
  assign n3828 = pi139  & pi140 ;
  assign n3829 = pi141  & ~n3796;
  assign n3830 = ~n3828 & ~n3829;
  assign n3831 = ~n3827 & ~n3830;
  assign n3832 = ~n3808 & n3831;
  assign n3833 = ~n3798 & ~n3805;
  assign n3834 = n3827 & n3830;
  assign n3835 = ~n3831 & ~n3834;
  assign n3836 = n3833 & n3835;
  assign n3837 = ~n3833 & ~n3835;
  assign n3838 = ~n3832 & ~n3836;
  assign n3839 = ~n3837 & n3838;
  assign n3840 = ~n3824 & n3839;
  assign n3841 = ~n3819 & ~n3840;
  assign n3842 = ~n3812 & n3820;
  assign n3843 = n3815 & ~n3842;
  assign n3844 = n3812 & ~n3820;
  assign n3845 = ~n3843 & ~n3844;
  assign n3846 = ~n3841 & n3845;
  assign n3847 = n3841 & ~n3845;
  assign n3848 = ~n3846 & ~n3847;
  assign n3849 = n3833 & ~n3834;
  assign n3850 = ~n3831 & ~n3849;
  assign n3851 = n3848 & ~n3850;
  assign n3852 = ~n3848 & n3850;
  assign n3853 = ~n3851 & ~n3852;
  assign n3854 = n3774 & ~n3853;
  assign n3855 = ~n3774 & n3853;
  assign n3856 = n3791 & n3808;
  assign n3857 = ~n3809 & ~n3856;
  assign n3858 = n3712 & n3729;
  assign n3859 = ~n3730 & ~n3858;
  assign n3860 = n3857 & n3859;
  assign n3861 = ~n3819 & ~n3824;
  assign n3862 = n3839 & n3861;
  assign n3863 = ~n3839 & ~n3861;
  assign n3864 = ~n3862 & ~n3863;
  assign n3865 = n3860 & n3864;
  assign n3866 = ~n3860 & ~n3864;
  assign n3867 = ~n3746 & ~n3747;
  assign n3868 = ~n3760 & n3867;
  assign n3869 = n3760 & ~n3867;
  assign n3870 = ~n3868 & ~n3869;
  assign n3871 = ~n3866 & n3870;
  assign n3872 = ~n3865 & ~n3871;
  assign n3873 = ~n3855 & n3872;
  assign n3874 = ~n3854 & ~n3873;
  assign n3875 = ~n3847 & ~n3850;
  assign n3876 = ~n3846 & ~n3875;
  assign n3877 = ~n3874 & n3876;
  assign n3878 = n3874 & ~n3876;
  assign n3879 = ~n3766 & n3771;
  assign n3880 = ~n3765 & ~n3879;
  assign n3881 = ~n3878 & n3880;
  assign n3882 = ~n3877 & ~n3881;
  assign n3883 = ~pi157  & pi158 ;
  assign n3884 = pi157  & ~pi158 ;
  assign n3885 = pi159  & ~n3883;
  assign n3886 = ~n3884 & n3885;
  assign n3887 = ~n3883 & ~n3884;
  assign n3888 = ~pi159  & ~n3887;
  assign n3889 = ~n3886 & ~n3888;
  assign n3890 = ~pi160  & pi161 ;
  assign n3891 = pi160  & ~pi161 ;
  assign n3892 = pi162  & ~n3890;
  assign n3893 = ~n3891 & n3892;
  assign n3894 = ~n3890 & ~n3891;
  assign n3895 = ~pi162  & ~n3894;
  assign n3896 = ~n3893 & ~n3895;
  assign n3897 = ~n3889 & n3896;
  assign n3898 = n3889 & ~n3896;
  assign n3899 = ~n3897 & ~n3898;
  assign n3900 = ~pi151  & pi152 ;
  assign n3901 = pi151  & ~pi152 ;
  assign n3902 = pi153  & ~n3900;
  assign n3903 = ~n3901 & n3902;
  assign n3904 = ~n3900 & ~n3901;
  assign n3905 = ~pi153  & ~n3904;
  assign n3906 = ~n3903 & ~n3905;
  assign n3907 = ~pi154  & pi155 ;
  assign n3908 = pi154  & ~pi155 ;
  assign n3909 = pi156  & ~n3907;
  assign n3910 = ~n3908 & n3909;
  assign n3911 = ~n3907 & ~n3908;
  assign n3912 = ~pi156  & ~n3911;
  assign n3913 = ~n3910 & ~n3912;
  assign n3914 = ~n3906 & n3913;
  assign n3915 = n3906 & ~n3913;
  assign n3916 = ~n3914 & ~n3915;
  assign n3917 = ~n3899 & ~n3916;
  assign n3918 = pi160  & pi161 ;
  assign n3919 = pi162  & ~n3894;
  assign n3920 = ~n3918 & ~n3919;
  assign n3921 = pi157  & pi158 ;
  assign n3922 = pi159  & ~n3887;
  assign n3923 = ~n3921 & ~n3922;
  assign n3924 = ~n3920 & ~n3923;
  assign n3925 = ~n3899 & n3924;
  assign n3926 = ~n3889 & ~n3896;
  assign n3927 = n3920 & n3923;
  assign n3928 = ~n3924 & ~n3927;
  assign n3929 = n3926 & n3928;
  assign n3930 = ~n3926 & ~n3928;
  assign n3931 = ~n3925 & ~n3929;
  assign n3932 = ~n3930 & n3931;
  assign n3933 = n3917 & n3932;
  assign n3934 = ~n3917 & ~n3932;
  assign n3935 = pi154  & pi155 ;
  assign n3936 = pi156  & ~n3911;
  assign n3937 = ~n3935 & ~n3936;
  assign n3938 = pi151  & pi152 ;
  assign n3939 = pi153  & ~n3904;
  assign n3940 = ~n3938 & ~n3939;
  assign n3941 = ~n3937 & n3940;
  assign n3942 = n3937 & ~n3940;
  assign n3943 = ~n3941 & ~n3942;
  assign n3944 = ~n3906 & ~n3913;
  assign n3945 = n3943 & n3944;
  assign n3946 = ~n3943 & ~n3944;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = ~n3934 & ~n3947;
  assign n3949 = ~n3933 & ~n3948;
  assign n3950 = n3926 & ~n3927;
  assign n3951 = ~n3924 & ~n3950;
  assign n3952 = ~n3949 & ~n3951;
  assign n3953 = n3949 & n3951;
  assign n3954 = ~n3952 & ~n3953;
  assign n3955 = ~n3937 & n3944;
  assign n3956 = n3940 & ~n3955;
  assign n3957 = n3937 & ~n3944;
  assign n3958 = ~n3956 & ~n3957;
  assign n3959 = ~n3954 & n3958;
  assign n3960 = n3954 & ~n3958;
  assign n3961 = ~n3959 & ~n3960;
  assign n3962 = ~pi169  & pi170 ;
  assign n3963 = pi169  & ~pi170 ;
  assign n3964 = pi171  & ~n3962;
  assign n3965 = ~n3963 & n3964;
  assign n3966 = ~n3962 & ~n3963;
  assign n3967 = ~pi171  & ~n3966;
  assign n3968 = ~n3965 & ~n3967;
  assign n3969 = ~pi172  & pi173 ;
  assign n3970 = pi172  & ~pi173 ;
  assign n3971 = pi174  & ~n3969;
  assign n3972 = ~n3970 & n3971;
  assign n3973 = ~n3969 & ~n3970;
  assign n3974 = ~pi174  & ~n3973;
  assign n3975 = ~n3972 & ~n3974;
  assign n3976 = ~n3968 & n3975;
  assign n3977 = n3968 & ~n3975;
  assign n3978 = ~n3976 & ~n3977;
  assign n3979 = ~pi163  & pi164 ;
  assign n3980 = pi163  & ~pi164 ;
  assign n3981 = pi165  & ~n3979;
  assign n3982 = ~n3980 & n3981;
  assign n3983 = ~n3979 & ~n3980;
  assign n3984 = ~pi165  & ~n3983;
  assign n3985 = ~n3982 & ~n3984;
  assign n3986 = ~pi166  & pi167 ;
  assign n3987 = pi166  & ~pi167 ;
  assign n3988 = pi168  & ~n3986;
  assign n3989 = ~n3987 & n3988;
  assign n3990 = ~n3986 & ~n3987;
  assign n3991 = ~pi168  & ~n3990;
  assign n3992 = ~n3989 & ~n3991;
  assign n3993 = ~n3985 & n3992;
  assign n3994 = n3985 & ~n3992;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = ~n3978 & ~n3995;
  assign n3997 = pi172  & pi173 ;
  assign n3998 = pi174  & ~n3973;
  assign n3999 = ~n3997 & ~n3998;
  assign n4000 = pi169  & pi170 ;
  assign n4001 = pi171  & ~n3966;
  assign n4002 = ~n4000 & ~n4001;
  assign n4003 = n3999 & ~n4002;
  assign n4004 = ~n3999 & n4002;
  assign n4005 = ~n4003 & ~n4004;
  assign n4006 = n3996 & ~n4005;
  assign n4007 = ~n3968 & ~n3975;
  assign n4008 = n4005 & n4007;
  assign n4009 = ~n4005 & ~n4007;
  assign n4010 = ~n3996 & ~n4008;
  assign n4011 = ~n4009 & n4010;
  assign n4012 = pi166  & pi167 ;
  assign n4013 = pi168  & ~n3990;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = pi163  & pi164 ;
  assign n4016 = pi165  & ~n3983;
  assign n4017 = ~n4015 & ~n4016;
  assign n4018 = ~n4014 & ~n4017;
  assign n4019 = ~n3995 & n4018;
  assign n4020 = ~n3985 & ~n3992;
  assign n4021 = n4014 & n4017;
  assign n4022 = ~n4018 & ~n4021;
  assign n4023 = n4020 & n4022;
  assign n4024 = ~n4020 & ~n4022;
  assign n4025 = ~n4019 & ~n4023;
  assign n4026 = ~n4024 & n4025;
  assign n4027 = ~n4011 & n4026;
  assign n4028 = ~n4006 & ~n4027;
  assign n4029 = ~n3999 & n4007;
  assign n4030 = n4002 & ~n4029;
  assign n4031 = n3999 & ~n4007;
  assign n4032 = ~n4030 & ~n4031;
  assign n4033 = ~n4028 & n4032;
  assign n4034 = n4028 & ~n4032;
  assign n4035 = ~n4033 & ~n4034;
  assign n4036 = n4020 & ~n4021;
  assign n4037 = ~n4018 & ~n4036;
  assign n4038 = n4035 & ~n4037;
  assign n4039 = ~n4035 & n4037;
  assign n4040 = ~n4038 & ~n4039;
  assign n4041 = n3961 & ~n4040;
  assign n4042 = ~n3961 & n4040;
  assign n4043 = n3978 & n3995;
  assign n4044 = ~n3996 & ~n4043;
  assign n4045 = n3899 & n3916;
  assign n4046 = ~n3917 & ~n4045;
  assign n4047 = n4044 & n4046;
  assign n4048 = ~n4006 & ~n4011;
  assign n4049 = n4026 & n4048;
  assign n4050 = ~n4026 & ~n4048;
  assign n4051 = ~n4049 & ~n4050;
  assign n4052 = n4047 & n4051;
  assign n4053 = ~n4047 & ~n4051;
  assign n4054 = ~n3933 & ~n3934;
  assign n4055 = ~n3947 & n4054;
  assign n4056 = n3947 & ~n4054;
  assign n4057 = ~n4055 & ~n4056;
  assign n4058 = ~n4053 & n4057;
  assign n4059 = ~n4052 & ~n4058;
  assign n4060 = ~n4042 & n4059;
  assign n4061 = ~n4041 & ~n4060;
  assign n4062 = ~n4034 & ~n4037;
  assign n4063 = ~n4033 & ~n4062;
  assign n4064 = ~n4061 & n4063;
  assign n4065 = n4061 & ~n4063;
  assign n4066 = ~n3953 & n3958;
  assign n4067 = ~n3952 & ~n4066;
  assign n4068 = ~n4065 & n4067;
  assign n4069 = ~n4064 & ~n4068;
  assign n4070 = ~n4064 & ~n4065;
  assign n4071 = n4067 & n4070;
  assign n4072 = ~n4067 & ~n4070;
  assign n4073 = ~n4071 & ~n4072;
  assign n4074 = ~n3877 & ~n3878;
  assign n4075 = n3880 & n4074;
  assign n4076 = ~n3880 & ~n4074;
  assign n4077 = ~n4075 & ~n4076;
  assign n4078 = ~n4073 & ~n4077;
  assign n4079 = n4073 & n4077;
  assign n4080 = ~n3854 & ~n3855;
  assign n4081 = ~n3872 & n4080;
  assign n4082 = n3872 & ~n4080;
  assign n4083 = ~n4081 & ~n4082;
  assign n4084 = ~n4041 & ~n4042;
  assign n4085 = ~n4059 & n4084;
  assign n4086 = n4059 & ~n4084;
  assign n4087 = ~n4085 & ~n4086;
  assign n4088 = ~n4083 & ~n4087;
  assign n4089 = n4083 & n4087;
  assign n4090 = ~n4044 & ~n4046;
  assign n4091 = ~n4047 & ~n4090;
  assign n4092 = ~n3857 & ~n3859;
  assign n4093 = ~n3860 & ~n4092;
  assign n4094 = n4091 & n4093;
  assign n4095 = ~n4052 & ~n4053;
  assign n4096 = ~n4057 & n4095;
  assign n4097 = n4057 & ~n4095;
  assign n4098 = ~n4096 & ~n4097;
  assign n4099 = n4094 & ~n4098;
  assign n4100 = ~n4094 & n4098;
  assign n4101 = ~n3865 & ~n3866;
  assign n4102 = ~n3870 & n4101;
  assign n4103 = n3870 & ~n4101;
  assign n4104 = ~n4102 & ~n4103;
  assign n4105 = ~n4100 & ~n4104;
  assign n4106 = ~n4099 & ~n4105;
  assign n4107 = ~n4089 & n4106;
  assign n4108 = ~n4088 & ~n4107;
  assign n4109 = ~n4079 & n4108;
  assign n4110 = ~n4078 & ~n4109;
  assign n4111 = ~n4069 & n4110;
  assign n4112 = n4069 & ~n4110;
  assign n4113 = ~n4111 & ~n4112;
  assign n4114 = n3882 & n4113;
  assign n4115 = ~n3882 & ~n4113;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = ~n3695 & ~n4116;
  assign n4118 = n3695 & n4116;
  assign n4119 = ~n4078 & ~n4079;
  assign n4120 = ~n4108 & n4119;
  assign n4121 = n4108 & ~n4119;
  assign n4122 = ~n4120 & ~n4121;
  assign n4123 = ~n3657 & ~n3658;
  assign n4124 = ~n3687 & n4123;
  assign n4125 = n3687 & ~n4123;
  assign n4126 = ~n4124 & ~n4125;
  assign n4127 = ~n4122 & ~n4126;
  assign n4128 = n4122 & n4126;
  assign n4129 = ~n3667 & ~n3668;
  assign n4130 = ~n3685 & n4129;
  assign n4131 = n3685 & ~n4129;
  assign n4132 = ~n4130 & ~n4131;
  assign n4133 = ~n4088 & ~n4089;
  assign n4134 = ~n4106 & n4133;
  assign n4135 = n4106 & ~n4133;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = ~n4132 & ~n4136;
  assign n4138 = n4132 & n4136;
  assign n4139 = n4091 & ~n4093;
  assign n4140 = ~n4091 & n4093;
  assign n4141 = ~n4139 & ~n4140;
  assign n4142 = n3670 & ~n3672;
  assign n4143 = ~n3670 & n3672;
  assign n4144 = ~n4142 & ~n4143;
  assign n4145 = ~n4141 & ~n4144;
  assign n4146 = ~n4099 & ~n4100;
  assign n4147 = n4104 & n4146;
  assign n4148 = ~n4104 & ~n4146;
  assign n4149 = ~n4147 & ~n4148;
  assign n4150 = n4145 & ~n4149;
  assign n4151 = ~n4145 & n4149;
  assign n4152 = ~n3678 & ~n3679;
  assign n4153 = n3683 & n4152;
  assign n4154 = ~n3683 & ~n4152;
  assign n4155 = ~n4153 & ~n4154;
  assign n4156 = ~n4151 & ~n4155;
  assign n4157 = ~n4150 & ~n4156;
  assign n4158 = ~n4138 & n4157;
  assign n4159 = ~n4137 & ~n4158;
  assign n4160 = ~n4128 & n4159;
  assign n4161 = ~n4127 & ~n4160;
  assign n4162 = ~n4118 & n4161;
  assign n4163 = ~n4117 & ~n4162;
  assign n4164 = ~n3882 & ~n4112;
  assign n4165 = ~n4111 & ~n4164;
  assign n4166 = ~n4163 & ~n4165;
  assign n4167 = n4163 & n4165;
  assign n4168 = ~n3461 & ~n3691;
  assign n4169 = ~n3690 & ~n4168;
  assign n4170 = ~n4167 & ~n4169;
  assign n4171 = ~n4166 & ~n4170;
  assign n4172 = ~pi181  & pi182 ;
  assign n4173 = pi181  & ~pi182 ;
  assign n4174 = pi183  & ~n4172;
  assign n4175 = ~n4173 & n4174;
  assign n4176 = ~n4172 & ~n4173;
  assign n4177 = ~pi183  & ~n4176;
  assign n4178 = ~n4175 & ~n4177;
  assign n4179 = ~pi184  & pi185 ;
  assign n4180 = pi184  & ~pi185 ;
  assign n4181 = pi186  & ~n4179;
  assign n4182 = ~n4180 & n4181;
  assign n4183 = ~n4179 & ~n4180;
  assign n4184 = ~pi186  & ~n4183;
  assign n4185 = ~n4182 & ~n4184;
  assign n4186 = ~n4178 & n4185;
  assign n4187 = n4178 & ~n4185;
  assign n4188 = ~n4186 & ~n4187;
  assign n4189 = ~pi175  & pi176 ;
  assign n4190 = pi175  & ~pi176 ;
  assign n4191 = pi177  & ~n4189;
  assign n4192 = ~n4190 & n4191;
  assign n4193 = ~n4189 & ~n4190;
  assign n4194 = ~pi177  & ~n4193;
  assign n4195 = ~n4192 & ~n4194;
  assign n4196 = ~pi178  & pi179 ;
  assign n4197 = pi178  & ~pi179 ;
  assign n4198 = pi180  & ~n4196;
  assign n4199 = ~n4197 & n4198;
  assign n4200 = ~n4196 & ~n4197;
  assign n4201 = ~pi180  & ~n4200;
  assign n4202 = ~n4199 & ~n4201;
  assign n4203 = ~n4195 & n4202;
  assign n4204 = n4195 & ~n4202;
  assign n4205 = ~n4203 & ~n4204;
  assign n4206 = ~n4188 & ~n4205;
  assign n4207 = pi184  & pi185 ;
  assign n4208 = pi186  & ~n4183;
  assign n4209 = ~n4207 & ~n4208;
  assign n4210 = pi181  & pi182 ;
  assign n4211 = pi183  & ~n4176;
  assign n4212 = ~n4210 & ~n4211;
  assign n4213 = ~n4209 & ~n4212;
  assign n4214 = ~n4188 & n4213;
  assign n4215 = ~n4178 & ~n4185;
  assign n4216 = n4209 & n4212;
  assign n4217 = ~n4213 & ~n4216;
  assign n4218 = n4215 & n4217;
  assign n4219 = ~n4215 & ~n4217;
  assign n4220 = ~n4214 & ~n4218;
  assign n4221 = ~n4219 & n4220;
  assign n4222 = n4206 & n4221;
  assign n4223 = ~n4206 & ~n4221;
  assign n4224 = pi178  & pi179 ;
  assign n4225 = pi180  & ~n4200;
  assign n4226 = ~n4224 & ~n4225;
  assign n4227 = pi175  & pi176 ;
  assign n4228 = pi177  & ~n4193;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = ~n4226 & n4229;
  assign n4231 = n4226 & ~n4229;
  assign n4232 = ~n4230 & ~n4231;
  assign n4233 = ~n4195 & ~n4202;
  assign n4234 = n4232 & n4233;
  assign n4235 = ~n4232 & ~n4233;
  assign n4236 = ~n4234 & ~n4235;
  assign n4237 = ~n4223 & ~n4236;
  assign n4238 = ~n4222 & ~n4237;
  assign n4239 = n4215 & ~n4216;
  assign n4240 = ~n4213 & ~n4239;
  assign n4241 = ~n4238 & ~n4240;
  assign n4242 = n4238 & n4240;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = ~n4226 & n4233;
  assign n4245 = n4229 & ~n4244;
  assign n4246 = n4226 & ~n4233;
  assign n4247 = ~n4245 & ~n4246;
  assign n4248 = ~n4243 & n4247;
  assign n4249 = n4243 & ~n4247;
  assign n4250 = ~n4248 & ~n4249;
  assign n4251 = ~pi193  & pi194 ;
  assign n4252 = pi193  & ~pi194 ;
  assign n4253 = pi195  & ~n4251;
  assign n4254 = ~n4252 & n4253;
  assign n4255 = ~n4251 & ~n4252;
  assign n4256 = ~pi195  & ~n4255;
  assign n4257 = ~n4254 & ~n4256;
  assign n4258 = ~pi196  & pi197 ;
  assign n4259 = pi196  & ~pi197 ;
  assign n4260 = pi198  & ~n4258;
  assign n4261 = ~n4259 & n4260;
  assign n4262 = ~n4258 & ~n4259;
  assign n4263 = ~pi198  & ~n4262;
  assign n4264 = ~n4261 & ~n4263;
  assign n4265 = ~n4257 & n4264;
  assign n4266 = n4257 & ~n4264;
  assign n4267 = ~n4265 & ~n4266;
  assign n4268 = ~pi187  & pi188 ;
  assign n4269 = pi187  & ~pi188 ;
  assign n4270 = pi189  & ~n4268;
  assign n4271 = ~n4269 & n4270;
  assign n4272 = ~n4268 & ~n4269;
  assign n4273 = ~pi189  & ~n4272;
  assign n4274 = ~n4271 & ~n4273;
  assign n4275 = ~pi190  & pi191 ;
  assign n4276 = pi190  & ~pi191 ;
  assign n4277 = pi192  & ~n4275;
  assign n4278 = ~n4276 & n4277;
  assign n4279 = ~n4275 & ~n4276;
  assign n4280 = ~pi192  & ~n4279;
  assign n4281 = ~n4278 & ~n4280;
  assign n4282 = ~n4274 & n4281;
  assign n4283 = n4274 & ~n4281;
  assign n4284 = ~n4282 & ~n4283;
  assign n4285 = ~n4267 & ~n4284;
  assign n4286 = pi196  & pi197 ;
  assign n4287 = pi198  & ~n4262;
  assign n4288 = ~n4286 & ~n4287;
  assign n4289 = pi193  & pi194 ;
  assign n4290 = pi195  & ~n4255;
  assign n4291 = ~n4289 & ~n4290;
  assign n4292 = n4288 & ~n4291;
  assign n4293 = ~n4288 & n4291;
  assign n4294 = ~n4292 & ~n4293;
  assign n4295 = n4285 & ~n4294;
  assign n4296 = ~n4257 & ~n4264;
  assign n4297 = n4294 & n4296;
  assign n4298 = ~n4294 & ~n4296;
  assign n4299 = ~n4285 & ~n4297;
  assign n4300 = ~n4298 & n4299;
  assign n4301 = pi190  & pi191 ;
  assign n4302 = pi192  & ~n4279;
  assign n4303 = ~n4301 & ~n4302;
  assign n4304 = pi187  & pi188 ;
  assign n4305 = pi189  & ~n4272;
  assign n4306 = ~n4304 & ~n4305;
  assign n4307 = ~n4303 & ~n4306;
  assign n4308 = ~n4284 & n4307;
  assign n4309 = ~n4274 & ~n4281;
  assign n4310 = n4303 & n4306;
  assign n4311 = ~n4307 & ~n4310;
  assign n4312 = n4309 & n4311;
  assign n4313 = ~n4309 & ~n4311;
  assign n4314 = ~n4308 & ~n4312;
  assign n4315 = ~n4313 & n4314;
  assign n4316 = ~n4300 & n4315;
  assign n4317 = ~n4295 & ~n4316;
  assign n4318 = ~n4288 & n4296;
  assign n4319 = n4291 & ~n4318;
  assign n4320 = n4288 & ~n4296;
  assign n4321 = ~n4319 & ~n4320;
  assign n4322 = ~n4317 & n4321;
  assign n4323 = n4317 & ~n4321;
  assign n4324 = ~n4322 & ~n4323;
  assign n4325 = n4309 & ~n4310;
  assign n4326 = ~n4307 & ~n4325;
  assign n4327 = n4324 & ~n4326;
  assign n4328 = ~n4324 & n4326;
  assign n4329 = ~n4327 & ~n4328;
  assign n4330 = n4250 & ~n4329;
  assign n4331 = ~n4250 & n4329;
  assign n4332 = n4267 & n4284;
  assign n4333 = ~n4285 & ~n4332;
  assign n4334 = n4188 & n4205;
  assign n4335 = ~n4206 & ~n4334;
  assign n4336 = n4333 & n4335;
  assign n4337 = ~n4295 & ~n4300;
  assign n4338 = n4315 & n4337;
  assign n4339 = ~n4315 & ~n4337;
  assign n4340 = ~n4338 & ~n4339;
  assign n4341 = n4336 & n4340;
  assign n4342 = ~n4336 & ~n4340;
  assign n4343 = ~n4222 & ~n4223;
  assign n4344 = ~n4236 & n4343;
  assign n4345 = n4236 & ~n4343;
  assign n4346 = ~n4344 & ~n4345;
  assign n4347 = ~n4342 & n4346;
  assign n4348 = ~n4341 & ~n4347;
  assign n4349 = ~n4331 & n4348;
  assign n4350 = ~n4330 & ~n4349;
  assign n4351 = ~n4323 & ~n4326;
  assign n4352 = ~n4322 & ~n4351;
  assign n4353 = ~n4350 & n4352;
  assign n4354 = n4350 & ~n4352;
  assign n4355 = ~n4242 & n4247;
  assign n4356 = ~n4241 & ~n4355;
  assign n4357 = ~n4354 & n4356;
  assign n4358 = ~n4353 & ~n4357;
  assign n4359 = pi199  & ~pi200 ;
  assign n4360 = ~pi199  & pi200 ;
  assign n4361 = pi201  & ~n4359;
  assign n4362 = ~n4360 & n4361;
  assign n4363 = ~n4359 & ~n4360;
  assign n4364 = ~pi201  & ~n4363;
  assign n4365 = ~n4362 & ~n4364;
  assign n4366 = pi202  & ~pi203 ;
  assign n4367 = ~pi202  & pi203 ;
  assign n4368 = pi204  & ~n4366;
  assign n4369 = ~n4367 & n4368;
  assign n4370 = ~n4366 & ~n4367;
  assign n4371 = ~pi204  & ~n4370;
  assign n4372 = ~n4369 & ~n4371;
  assign n4373 = ~n4365 & n4372;
  assign n4374 = n4365 & ~n4372;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = pi205  & ~pi206 ;
  assign n4377 = ~pi205  & pi206 ;
  assign n4378 = pi207  & ~n4376;
  assign n4379 = ~n4377 & n4378;
  assign n4380 = ~n4376 & ~n4377;
  assign n4381 = ~pi207  & ~n4380;
  assign n4382 = ~n4379 & ~n4381;
  assign n4383 = pi208  & ~pi209 ;
  assign n4384 = ~pi208  & pi209 ;
  assign n4385 = pi210  & ~n4383;
  assign n4386 = ~n4384 & n4385;
  assign n4387 = ~n4383 & ~n4384;
  assign n4388 = ~pi210  & ~n4387;
  assign n4389 = ~n4386 & ~n4388;
  assign n4390 = ~n4382 & n4389;
  assign n4391 = n4382 & ~n4389;
  assign n4392 = ~n4390 & ~n4391;
  assign n4393 = ~n4375 & ~n4392;
  assign n4394 = pi208  & pi209 ;
  assign n4395 = pi210  & ~n4387;
  assign n4396 = ~n4394 & ~n4395;
  assign n4397 = pi205  & pi206 ;
  assign n4398 = pi207  & ~n4380;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n4396 & ~n4399;
  assign n4401 = ~n4392 & n4400;
  assign n4402 = ~n4382 & ~n4389;
  assign n4403 = n4396 & n4399;
  assign n4404 = ~n4400 & ~n4403;
  assign n4405 = n4402 & n4404;
  assign n4406 = ~n4402 & ~n4404;
  assign n4407 = ~n4401 & ~n4405;
  assign n4408 = ~n4406 & n4407;
  assign n4409 = n4393 & n4408;
  assign n4410 = ~n4393 & ~n4408;
  assign n4411 = ~n4365 & ~n4372;
  assign n4412 = pi202  & pi203 ;
  assign n4413 = pi204  & ~n4370;
  assign n4414 = ~n4412 & ~n4413;
  assign n4415 = pi199  & pi200 ;
  assign n4416 = pi201  & ~n4363;
  assign n4417 = ~n4415 & ~n4416;
  assign n4418 = n4414 & ~n4417;
  assign n4419 = ~n4414 & n4417;
  assign n4420 = ~n4418 & ~n4419;
  assign n4421 = n4411 & n4420;
  assign n4422 = ~n4411 & ~n4420;
  assign n4423 = ~n4421 & ~n4422;
  assign n4424 = ~n4410 & ~n4423;
  assign n4425 = ~n4409 & ~n4424;
  assign n4426 = n4402 & ~n4403;
  assign n4427 = ~n4400 & ~n4426;
  assign n4428 = ~n4425 & ~n4427;
  assign n4429 = n4425 & n4427;
  assign n4430 = ~n4428 & ~n4429;
  assign n4431 = n4411 & ~n4414;
  assign n4432 = n4417 & ~n4431;
  assign n4433 = ~n4411 & n4414;
  assign n4434 = ~n4432 & ~n4433;
  assign n4435 = ~n4430 & n4434;
  assign n4436 = n4430 & ~n4434;
  assign n4437 = ~n4435 & ~n4436;
  assign n4438 = pi217  & ~pi218 ;
  assign n4439 = ~pi217  & pi218 ;
  assign n4440 = pi219  & ~n4438;
  assign n4441 = ~n4439 & n4440;
  assign n4442 = ~n4438 & ~n4439;
  assign n4443 = ~pi219  & ~n4442;
  assign n4444 = ~n4441 & ~n4443;
  assign n4445 = pi220  & ~pi221 ;
  assign n4446 = ~pi220  & pi221 ;
  assign n4447 = pi222  & ~n4445;
  assign n4448 = ~n4446 & n4447;
  assign n4449 = ~n4445 & ~n4446;
  assign n4450 = ~pi222  & ~n4449;
  assign n4451 = ~n4448 & ~n4450;
  assign n4452 = ~n4444 & n4451;
  assign n4453 = n4444 & ~n4451;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = pi220  & pi221 ;
  assign n4456 = pi222  & ~n4449;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = pi217  & pi218 ;
  assign n4459 = pi219  & ~n4442;
  assign n4460 = ~n4458 & ~n4459;
  assign n4461 = ~n4457 & ~n4460;
  assign n4462 = ~n4454 & n4461;
  assign n4463 = ~n4444 & ~n4451;
  assign n4464 = n4457 & n4460;
  assign n4465 = ~n4461 & ~n4464;
  assign n4466 = n4463 & n4465;
  assign n4467 = ~n4463 & ~n4465;
  assign n4468 = ~n4462 & ~n4466;
  assign n4469 = ~n4467 & n4468;
  assign n4470 = pi211  & ~pi212 ;
  assign n4471 = ~pi211  & pi212 ;
  assign n4472 = pi213  & ~n4470;
  assign n4473 = ~n4471 & n4472;
  assign n4474 = ~n4470 & ~n4471;
  assign n4475 = ~pi213  & ~n4474;
  assign n4476 = ~n4473 & ~n4475;
  assign n4477 = pi214  & ~pi215 ;
  assign n4478 = ~pi214  & pi215 ;
  assign n4479 = pi216  & ~n4477;
  assign n4480 = ~n4478 & n4479;
  assign n4481 = ~n4477 & ~n4478;
  assign n4482 = ~pi216  & ~n4481;
  assign n4483 = ~n4480 & ~n4482;
  assign n4484 = ~n4476 & n4483;
  assign n4485 = n4476 & ~n4483;
  assign n4486 = ~n4484 & ~n4485;
  assign n4487 = ~n4454 & ~n4486;
  assign n4488 = ~n4476 & ~n4483;
  assign n4489 = pi214  & pi215 ;
  assign n4490 = pi216  & ~n4481;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = pi211  & pi212 ;
  assign n4493 = pi213  & ~n4474;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495 = n4491 & ~n4494;
  assign n4496 = ~n4491 & n4494;
  assign n4497 = ~n4495 & ~n4496;
  assign n4498 = n4488 & n4497;
  assign n4499 = ~n4488 & ~n4497;
  assign n4500 = ~n4498 & ~n4499;
  assign n4501 = ~n4487 & n4500;
  assign n4502 = n4469 & ~n4501;
  assign n4503 = n4487 & ~n4500;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = n4463 & ~n4464;
  assign n4506 = ~n4461 & ~n4505;
  assign n4507 = ~n4504 & ~n4506;
  assign n4508 = n4504 & n4506;
  assign n4509 = ~n4507 & ~n4508;
  assign n4510 = n4488 & ~n4491;
  assign n4511 = n4494 & ~n4510;
  assign n4512 = ~n4488 & n4491;
  assign n4513 = ~n4511 & ~n4512;
  assign n4514 = ~n4509 & n4513;
  assign n4515 = n4509 & ~n4513;
  assign n4516 = ~n4514 & ~n4515;
  assign n4517 = ~n4437 & ~n4516;
  assign n4518 = n4437 & n4516;
  assign n4519 = n4454 & n4486;
  assign n4520 = ~n4487 & ~n4519;
  assign n4521 = n4375 & n4392;
  assign n4522 = ~n4393 & ~n4521;
  assign n4523 = n4520 & n4522;
  assign n4524 = n4487 & ~n4497;
  assign n4525 = ~n4501 & ~n4524;
  assign n4526 = n4469 & ~n4525;
  assign n4527 = ~n4469 & n4525;
  assign n4528 = ~n4526 & ~n4527;
  assign n4529 = n4523 & ~n4528;
  assign n4530 = ~n4523 & n4528;
  assign n4531 = ~n4409 & ~n4410;
  assign n4532 = ~n4423 & n4531;
  assign n4533 = n4423 & ~n4531;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = ~n4530 & n4534;
  assign n4536 = ~n4529 & ~n4535;
  assign n4537 = ~n4518 & ~n4536;
  assign n4538 = ~n4517 & ~n4537;
  assign n4539 = ~n4508 & n4513;
  assign n4540 = ~n4507 & ~n4539;
  assign n4541 = ~n4538 & ~n4540;
  assign n4542 = n4538 & n4540;
  assign n4543 = ~n4429 & n4434;
  assign n4544 = ~n4428 & ~n4543;
  assign n4545 = ~n4542 & ~n4544;
  assign n4546 = ~n4541 & ~n4545;
  assign n4547 = ~n4541 & ~n4542;
  assign n4548 = n4544 & ~n4547;
  assign n4549 = ~n4541 & n4545;
  assign n4550 = ~n4548 & ~n4549;
  assign n4551 = ~n4353 & ~n4354;
  assign n4552 = n4356 & n4551;
  assign n4553 = ~n4356 & ~n4551;
  assign n4554 = ~n4552 & ~n4553;
  assign n4555 = n4550 & ~n4554;
  assign n4556 = ~n4550 & n4554;
  assign n4557 = ~n4330 & ~n4331;
  assign n4558 = ~n4348 & n4557;
  assign n4559 = n4348 & ~n4557;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = ~n4517 & ~n4518;
  assign n4562 = ~n4536 & n4561;
  assign n4563 = n4536 & ~n4561;
  assign n4564 = ~n4562 & ~n4563;
  assign n4565 = ~n4560 & ~n4564;
  assign n4566 = n4560 & n4564;
  assign n4567 = ~n4520 & ~n4522;
  assign n4568 = ~n4523 & ~n4567;
  assign n4569 = ~n4333 & ~n4335;
  assign n4570 = ~n4336 & ~n4569;
  assign n4571 = n4568 & n4570;
  assign n4572 = ~n4529 & ~n4530;
  assign n4573 = ~n4534 & n4572;
  assign n4574 = n4534 & ~n4572;
  assign n4575 = ~n4573 & ~n4574;
  assign n4576 = n4571 & ~n4575;
  assign n4577 = ~n4571 & n4575;
  assign n4578 = ~n4341 & ~n4342;
  assign n4579 = ~n4346 & n4578;
  assign n4580 = n4346 & ~n4578;
  assign n4581 = ~n4579 & ~n4580;
  assign n4582 = ~n4577 & ~n4581;
  assign n4583 = ~n4576 & ~n4582;
  assign n4584 = ~n4566 & n4583;
  assign n4585 = ~n4565 & ~n4584;
  assign n4586 = ~n4556 & n4585;
  assign n4587 = ~n4555 & ~n4586;
  assign n4588 = n4546 & ~n4587;
  assign n4589 = ~n4546 & n4587;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = n4358 & n4590;
  assign n4592 = ~n4358 & ~n4590;
  assign n4593 = ~n4591 & ~n4592;
  assign n4594 = ~pi229  & pi230 ;
  assign n4595 = pi229  & ~pi230 ;
  assign n4596 = pi231  & ~n4594;
  assign n4597 = ~n4595 & n4596;
  assign n4598 = ~n4594 & ~n4595;
  assign n4599 = ~pi231  & ~n4598;
  assign n4600 = ~n4597 & ~n4599;
  assign n4601 = ~pi232  & pi233 ;
  assign n4602 = pi232  & ~pi233 ;
  assign n4603 = pi234  & ~n4601;
  assign n4604 = ~n4602 & n4603;
  assign n4605 = ~n4601 & ~n4602;
  assign n4606 = ~pi234  & ~n4605;
  assign n4607 = ~n4604 & ~n4606;
  assign n4608 = ~n4600 & n4607;
  assign n4609 = n4600 & ~n4607;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = ~pi223  & pi224 ;
  assign n4612 = pi223  & ~pi224 ;
  assign n4613 = pi225  & ~n4611;
  assign n4614 = ~n4612 & n4613;
  assign n4615 = ~n4611 & ~n4612;
  assign n4616 = ~pi225  & ~n4615;
  assign n4617 = ~n4614 & ~n4616;
  assign n4618 = ~pi226  & pi227 ;
  assign n4619 = pi226  & ~pi227 ;
  assign n4620 = pi228  & ~n4618;
  assign n4621 = ~n4619 & n4620;
  assign n4622 = ~n4618 & ~n4619;
  assign n4623 = ~pi228  & ~n4622;
  assign n4624 = ~n4621 & ~n4623;
  assign n4625 = ~n4617 & n4624;
  assign n4626 = n4617 & ~n4624;
  assign n4627 = ~n4625 & ~n4626;
  assign n4628 = ~n4610 & ~n4627;
  assign n4629 = pi232  & pi233 ;
  assign n4630 = pi234  & ~n4605;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = pi229  & pi230 ;
  assign n4633 = pi231  & ~n4598;
  assign n4634 = ~n4632 & ~n4633;
  assign n4635 = ~n4631 & ~n4634;
  assign n4636 = ~n4610 & n4635;
  assign n4637 = ~n4600 & ~n4607;
  assign n4638 = n4631 & n4634;
  assign n4639 = ~n4635 & ~n4638;
  assign n4640 = n4637 & n4639;
  assign n4641 = ~n4637 & ~n4639;
  assign n4642 = ~n4636 & ~n4640;
  assign n4643 = ~n4641 & n4642;
  assign n4644 = n4628 & n4643;
  assign n4645 = ~n4628 & ~n4643;
  assign n4646 = pi226  & pi227 ;
  assign n4647 = pi228  & ~n4622;
  assign n4648 = ~n4646 & ~n4647;
  assign n4649 = pi223  & pi224 ;
  assign n4650 = pi225  & ~n4615;
  assign n4651 = ~n4649 & ~n4650;
  assign n4652 = ~n4648 & n4651;
  assign n4653 = n4648 & ~n4651;
  assign n4654 = ~n4652 & ~n4653;
  assign n4655 = ~n4617 & ~n4624;
  assign n4656 = n4654 & n4655;
  assign n4657 = ~n4654 & ~n4655;
  assign n4658 = ~n4656 & ~n4657;
  assign n4659 = ~n4645 & ~n4658;
  assign n4660 = ~n4644 & ~n4659;
  assign n4661 = n4637 & ~n4638;
  assign n4662 = ~n4635 & ~n4661;
  assign n4663 = ~n4660 & ~n4662;
  assign n4664 = n4660 & n4662;
  assign n4665 = ~n4663 & ~n4664;
  assign n4666 = ~n4648 & n4655;
  assign n4667 = n4651 & ~n4666;
  assign n4668 = n4648 & ~n4655;
  assign n4669 = ~n4667 & ~n4668;
  assign n4670 = ~n4665 & n4669;
  assign n4671 = n4665 & ~n4669;
  assign n4672 = ~n4670 & ~n4671;
  assign n4673 = pi241  & ~pi242 ;
  assign n4674 = ~pi241  & pi242 ;
  assign n4675 = pi243  & ~n4673;
  assign n4676 = ~n4674 & n4675;
  assign n4677 = ~n4673 & ~n4674;
  assign n4678 = ~pi243  & ~n4677;
  assign n4679 = ~n4676 & ~n4678;
  assign n4680 = pi244  & ~pi245 ;
  assign n4681 = ~pi244  & pi245 ;
  assign n4682 = pi246  & ~n4680;
  assign n4683 = ~n4681 & n4682;
  assign n4684 = ~n4680 & ~n4681;
  assign n4685 = ~pi246  & ~n4684;
  assign n4686 = ~n4683 & ~n4685;
  assign n4687 = ~n4679 & n4686;
  assign n4688 = n4679 & ~n4686;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = pi244  & pi245 ;
  assign n4691 = pi246  & ~n4684;
  assign n4692 = ~n4690 & ~n4691;
  assign n4693 = pi241  & pi242 ;
  assign n4694 = pi243  & ~n4677;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = ~n4692 & ~n4695;
  assign n4697 = ~n4689 & n4696;
  assign n4698 = ~n4679 & ~n4686;
  assign n4699 = n4692 & n4695;
  assign n4700 = ~n4696 & ~n4699;
  assign n4701 = n4698 & n4700;
  assign n4702 = ~n4698 & ~n4700;
  assign n4703 = ~n4697 & ~n4701;
  assign n4704 = ~n4702 & n4703;
  assign n4705 = pi235  & ~pi236 ;
  assign n4706 = ~pi235  & pi236 ;
  assign n4707 = pi237  & ~n4705;
  assign n4708 = ~n4706 & n4707;
  assign n4709 = ~n4705 & ~n4706;
  assign n4710 = ~pi237  & ~n4709;
  assign n4711 = ~n4708 & ~n4710;
  assign n4712 = pi238  & ~pi239 ;
  assign n4713 = ~pi238  & pi239 ;
  assign n4714 = pi240  & ~n4712;
  assign n4715 = ~n4713 & n4714;
  assign n4716 = ~n4712 & ~n4713;
  assign n4717 = ~pi240  & ~n4716;
  assign n4718 = ~n4715 & ~n4717;
  assign n4719 = ~n4711 & n4718;
  assign n4720 = n4711 & ~n4718;
  assign n4721 = ~n4719 & ~n4720;
  assign n4722 = ~n4689 & ~n4721;
  assign n4723 = ~n4711 & ~n4718;
  assign n4724 = pi238  & pi239 ;
  assign n4725 = pi240  & ~n4716;
  assign n4726 = ~n4724 & ~n4725;
  assign n4727 = pi235  & pi236 ;
  assign n4728 = pi237  & ~n4709;
  assign n4729 = ~n4727 & ~n4728;
  assign n4730 = n4726 & ~n4729;
  assign n4731 = ~n4726 & n4729;
  assign n4732 = ~n4730 & ~n4731;
  assign n4733 = n4723 & n4732;
  assign n4734 = ~n4723 & ~n4732;
  assign n4735 = ~n4733 & ~n4734;
  assign n4736 = ~n4722 & n4735;
  assign n4737 = n4704 & ~n4736;
  assign n4738 = n4722 & ~n4735;
  assign n4739 = ~n4737 & ~n4738;
  assign n4740 = n4698 & ~n4699;
  assign n4741 = ~n4696 & ~n4740;
  assign n4742 = ~n4739 & ~n4741;
  assign n4743 = n4739 & n4741;
  assign n4744 = ~n4742 & ~n4743;
  assign n4745 = n4723 & ~n4726;
  assign n4746 = n4729 & ~n4745;
  assign n4747 = ~n4723 & n4726;
  assign n4748 = ~n4746 & ~n4747;
  assign n4749 = ~n4744 & n4748;
  assign n4750 = n4744 & ~n4748;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = ~n4672 & ~n4751;
  assign n4753 = n4672 & n4751;
  assign n4754 = n4689 & n4721;
  assign n4755 = ~n4722 & ~n4754;
  assign n4756 = n4610 & n4627;
  assign n4757 = ~n4628 & ~n4756;
  assign n4758 = n4755 & n4757;
  assign n4759 = n4722 & ~n4732;
  assign n4760 = ~n4736 & ~n4759;
  assign n4761 = n4704 & ~n4760;
  assign n4762 = ~n4704 & n4760;
  assign n4763 = ~n4761 & ~n4762;
  assign n4764 = n4758 & ~n4763;
  assign n4765 = ~n4758 & n4763;
  assign n4766 = ~n4644 & ~n4645;
  assign n4767 = ~n4658 & n4766;
  assign n4768 = n4658 & ~n4766;
  assign n4769 = ~n4767 & ~n4768;
  assign n4770 = ~n4765 & n4769;
  assign n4771 = ~n4764 & ~n4770;
  assign n4772 = ~n4753 & ~n4771;
  assign n4773 = ~n4752 & ~n4772;
  assign n4774 = ~n4743 & n4748;
  assign n4775 = ~n4742 & ~n4774;
  assign n4776 = ~n4773 & ~n4775;
  assign n4777 = n4773 & n4775;
  assign n4778 = ~n4664 & n4669;
  assign n4779 = ~n4663 & ~n4778;
  assign n4780 = ~n4777 & ~n4779;
  assign n4781 = ~n4776 & ~n4780;
  assign n4782 = pi247  & ~pi248 ;
  assign n4783 = ~pi247  & pi248 ;
  assign n4784 = pi249  & ~n4782;
  assign n4785 = ~n4783 & n4784;
  assign n4786 = ~n4782 & ~n4783;
  assign n4787 = ~pi249  & ~n4786;
  assign n4788 = ~n4785 & ~n4787;
  assign n4789 = pi250  & ~pi251 ;
  assign n4790 = ~pi250  & pi251 ;
  assign n4791 = pi252  & ~n4789;
  assign n4792 = ~n4790 & n4791;
  assign n4793 = ~n4789 & ~n4790;
  assign n4794 = ~pi252  & ~n4793;
  assign n4795 = ~n4792 & ~n4794;
  assign n4796 = ~n4788 & n4795;
  assign n4797 = n4788 & ~n4795;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = pi253  & ~pi254 ;
  assign n4800 = ~pi253  & pi254 ;
  assign n4801 = pi255  & ~n4799;
  assign n4802 = ~n4800 & n4801;
  assign n4803 = ~n4799 & ~n4800;
  assign n4804 = ~pi255  & ~n4803;
  assign n4805 = ~n4802 & ~n4804;
  assign n4806 = pi256  & ~pi257 ;
  assign n4807 = ~pi256  & pi257 ;
  assign n4808 = pi258  & ~n4806;
  assign n4809 = ~n4807 & n4808;
  assign n4810 = ~n4806 & ~n4807;
  assign n4811 = ~pi258  & ~n4810;
  assign n4812 = ~n4809 & ~n4811;
  assign n4813 = ~n4805 & n4812;
  assign n4814 = n4805 & ~n4812;
  assign n4815 = ~n4813 & ~n4814;
  assign n4816 = ~n4798 & ~n4815;
  assign n4817 = pi256  & pi257 ;
  assign n4818 = pi258  & ~n4810;
  assign n4819 = ~n4817 & ~n4818;
  assign n4820 = pi253  & pi254 ;
  assign n4821 = pi255  & ~n4803;
  assign n4822 = ~n4820 & ~n4821;
  assign n4823 = ~n4819 & ~n4822;
  assign n4824 = ~n4815 & n4823;
  assign n4825 = ~n4805 & ~n4812;
  assign n4826 = n4819 & n4822;
  assign n4827 = ~n4823 & ~n4826;
  assign n4828 = n4825 & n4827;
  assign n4829 = ~n4825 & ~n4827;
  assign n4830 = ~n4824 & ~n4828;
  assign n4831 = ~n4829 & n4830;
  assign n4832 = n4816 & n4831;
  assign n4833 = ~n4816 & ~n4831;
  assign n4834 = ~n4788 & ~n4795;
  assign n4835 = pi250  & pi251 ;
  assign n4836 = pi252  & ~n4793;
  assign n4837 = ~n4835 & ~n4836;
  assign n4838 = pi247  & pi248 ;
  assign n4839 = pi249  & ~n4786;
  assign n4840 = ~n4838 & ~n4839;
  assign n4841 = n4837 & ~n4840;
  assign n4842 = ~n4837 & n4840;
  assign n4843 = ~n4841 & ~n4842;
  assign n4844 = n4834 & n4843;
  assign n4845 = ~n4834 & ~n4843;
  assign n4846 = ~n4844 & ~n4845;
  assign n4847 = ~n4833 & ~n4846;
  assign n4848 = ~n4832 & ~n4847;
  assign n4849 = n4825 & ~n4826;
  assign n4850 = ~n4823 & ~n4849;
  assign n4851 = ~n4848 & ~n4850;
  assign n4852 = n4848 & n4850;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = n4834 & ~n4837;
  assign n4855 = n4840 & ~n4854;
  assign n4856 = ~n4834 & n4837;
  assign n4857 = ~n4855 & ~n4856;
  assign n4858 = ~n4853 & n4857;
  assign n4859 = n4853 & ~n4857;
  assign n4860 = ~n4858 & ~n4859;
  assign n4861 = pi265  & ~pi266 ;
  assign n4862 = ~pi265  & pi266 ;
  assign n4863 = pi267  & ~n4861;
  assign n4864 = ~n4862 & n4863;
  assign n4865 = ~n4861 & ~n4862;
  assign n4866 = ~pi267  & ~n4865;
  assign n4867 = ~n4864 & ~n4866;
  assign n4868 = pi268  & ~pi269 ;
  assign n4869 = ~pi268  & pi269 ;
  assign n4870 = pi270  & ~n4868;
  assign n4871 = ~n4869 & n4870;
  assign n4872 = ~n4868 & ~n4869;
  assign n4873 = ~pi270  & ~n4872;
  assign n4874 = ~n4871 & ~n4873;
  assign n4875 = ~n4867 & n4874;
  assign n4876 = n4867 & ~n4874;
  assign n4877 = ~n4875 & ~n4876;
  assign n4878 = pi268  & pi269 ;
  assign n4879 = pi270  & ~n4872;
  assign n4880 = ~n4878 & ~n4879;
  assign n4881 = pi265  & pi266 ;
  assign n4882 = pi267  & ~n4865;
  assign n4883 = ~n4881 & ~n4882;
  assign n4884 = ~n4880 & ~n4883;
  assign n4885 = ~n4877 & n4884;
  assign n4886 = ~n4867 & ~n4874;
  assign n4887 = n4880 & n4883;
  assign n4888 = ~n4884 & ~n4887;
  assign n4889 = n4886 & n4888;
  assign n4890 = ~n4886 & ~n4888;
  assign n4891 = ~n4885 & ~n4889;
  assign n4892 = ~n4890 & n4891;
  assign n4893 = pi259  & ~pi260 ;
  assign n4894 = ~pi259  & pi260 ;
  assign n4895 = pi261  & ~n4893;
  assign n4896 = ~n4894 & n4895;
  assign n4897 = ~n4893 & ~n4894;
  assign n4898 = ~pi261  & ~n4897;
  assign n4899 = ~n4896 & ~n4898;
  assign n4900 = pi262  & ~pi263 ;
  assign n4901 = ~pi262  & pi263 ;
  assign n4902 = pi264  & ~n4900;
  assign n4903 = ~n4901 & n4902;
  assign n4904 = ~n4900 & ~n4901;
  assign n4905 = ~pi264  & ~n4904;
  assign n4906 = ~n4903 & ~n4905;
  assign n4907 = ~n4899 & n4906;
  assign n4908 = n4899 & ~n4906;
  assign n4909 = ~n4907 & ~n4908;
  assign n4910 = ~n4877 & ~n4909;
  assign n4911 = ~n4899 & ~n4906;
  assign n4912 = pi262  & pi263 ;
  assign n4913 = pi264  & ~n4904;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = pi259  & pi260 ;
  assign n4916 = pi261  & ~n4897;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = n4914 & ~n4917;
  assign n4919 = ~n4914 & n4917;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = n4911 & n4920;
  assign n4922 = ~n4911 & ~n4920;
  assign n4923 = ~n4921 & ~n4922;
  assign n4924 = ~n4910 & n4923;
  assign n4925 = n4892 & ~n4924;
  assign n4926 = n4910 & ~n4923;
  assign n4927 = ~n4925 & ~n4926;
  assign n4928 = n4886 & ~n4887;
  assign n4929 = ~n4884 & ~n4928;
  assign n4930 = ~n4927 & ~n4929;
  assign n4931 = n4927 & n4929;
  assign n4932 = ~n4930 & ~n4931;
  assign n4933 = n4911 & ~n4914;
  assign n4934 = n4917 & ~n4933;
  assign n4935 = ~n4911 & n4914;
  assign n4936 = ~n4934 & ~n4935;
  assign n4937 = ~n4932 & n4936;
  assign n4938 = n4932 & ~n4936;
  assign n4939 = ~n4937 & ~n4938;
  assign n4940 = ~n4860 & ~n4939;
  assign n4941 = n4860 & n4939;
  assign n4942 = n4877 & n4909;
  assign n4943 = ~n4910 & ~n4942;
  assign n4944 = n4798 & n4815;
  assign n4945 = ~n4816 & ~n4944;
  assign n4946 = n4943 & n4945;
  assign n4947 = n4910 & ~n4920;
  assign n4948 = ~n4924 & ~n4947;
  assign n4949 = n4892 & ~n4948;
  assign n4950 = ~n4892 & n4948;
  assign n4951 = ~n4949 & ~n4950;
  assign n4952 = n4946 & ~n4951;
  assign n4953 = ~n4946 & n4951;
  assign n4954 = ~n4832 & ~n4833;
  assign n4955 = ~n4846 & n4954;
  assign n4956 = n4846 & ~n4954;
  assign n4957 = ~n4955 & ~n4956;
  assign n4958 = ~n4953 & n4957;
  assign n4959 = ~n4952 & ~n4958;
  assign n4960 = ~n4941 & ~n4959;
  assign n4961 = ~n4940 & ~n4960;
  assign n4962 = ~n4931 & n4936;
  assign n4963 = ~n4930 & ~n4962;
  assign n4964 = ~n4961 & ~n4963;
  assign n4965 = n4961 & n4963;
  assign n4966 = ~n4852 & n4857;
  assign n4967 = ~n4851 & ~n4966;
  assign n4968 = ~n4965 & ~n4967;
  assign n4969 = ~n4964 & ~n4968;
  assign n4970 = ~n4964 & ~n4965;
  assign n4971 = n4967 & ~n4970;
  assign n4972 = ~n4964 & n4968;
  assign n4973 = ~n4971 & ~n4972;
  assign n4974 = ~n4776 & ~n4777;
  assign n4975 = n4779 & ~n4974;
  assign n4976 = ~n4776 & n4780;
  assign n4977 = ~n4975 & ~n4976;
  assign n4978 = ~n4973 & ~n4977;
  assign n4979 = n4973 & n4977;
  assign n4980 = ~n4752 & ~n4753;
  assign n4981 = ~n4771 & n4980;
  assign n4982 = n4771 & ~n4980;
  assign n4983 = ~n4981 & ~n4982;
  assign n4984 = ~n4940 & ~n4941;
  assign n4985 = ~n4959 & n4984;
  assign n4986 = n4959 & ~n4984;
  assign n4987 = ~n4985 & ~n4986;
  assign n4988 = ~n4983 & ~n4987;
  assign n4989 = n4983 & n4987;
  assign n4990 = ~n4943 & ~n4945;
  assign n4991 = ~n4946 & ~n4990;
  assign n4992 = ~n4755 & ~n4757;
  assign n4993 = ~n4758 & ~n4992;
  assign n4994 = n4991 & n4993;
  assign n4995 = ~n4952 & ~n4953;
  assign n4996 = ~n4957 & n4995;
  assign n4997 = n4957 & ~n4995;
  assign n4998 = ~n4996 & ~n4997;
  assign n4999 = n4994 & ~n4998;
  assign n5000 = ~n4994 & n4998;
  assign n5001 = ~n4764 & ~n4765;
  assign n5002 = ~n4769 & n5001;
  assign n5003 = n4769 & ~n5001;
  assign n5004 = ~n5002 & ~n5003;
  assign n5005 = ~n5000 & ~n5004;
  assign n5006 = ~n4999 & ~n5005;
  assign n5007 = ~n4989 & n5006;
  assign n5008 = ~n4988 & ~n5007;
  assign n5009 = ~n4979 & ~n5008;
  assign n5010 = ~n4978 & ~n5009;
  assign n5011 = n4969 & ~n5010;
  assign n5012 = ~n4969 & n5010;
  assign n5013 = ~n5011 & ~n5012;
  assign n5014 = n4781 & n5013;
  assign n5015 = ~n4781 & ~n5013;
  assign n5016 = ~n5014 & ~n5015;
  assign n5017 = ~n4593 & ~n5016;
  assign n5018 = n4593 & n5016;
  assign n5019 = ~n4978 & ~n4979;
  assign n5020 = ~n5008 & n5019;
  assign n5021 = n5008 & ~n5019;
  assign n5022 = ~n5020 & ~n5021;
  assign n5023 = ~n4555 & ~n4556;
  assign n5024 = ~n4585 & n5023;
  assign n5025 = n4585 & ~n5023;
  assign n5026 = ~n5024 & ~n5025;
  assign n5027 = ~n5022 & ~n5026;
  assign n5028 = n5022 & n5026;
  assign n5029 = ~n4565 & ~n4566;
  assign n5030 = ~n4583 & n5029;
  assign n5031 = n4583 & ~n5029;
  assign n5032 = ~n5030 & ~n5031;
  assign n5033 = ~n4988 & ~n4989;
  assign n5034 = ~n5006 & n5033;
  assign n5035 = n5006 & ~n5033;
  assign n5036 = ~n5034 & ~n5035;
  assign n5037 = ~n5032 & ~n5036;
  assign n5038 = n5032 & n5036;
  assign n5039 = n4991 & ~n4993;
  assign n5040 = ~n4991 & n4993;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = n4568 & ~n4570;
  assign n5043 = ~n4568 & n4570;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = ~n5041 & ~n5044;
  assign n5046 = ~n4999 & ~n5000;
  assign n5047 = n5004 & n5046;
  assign n5048 = ~n5004 & ~n5046;
  assign n5049 = ~n5047 & ~n5048;
  assign n5050 = n5045 & ~n5049;
  assign n5051 = ~n5045 & n5049;
  assign n5052 = ~n4576 & ~n4577;
  assign n5053 = n4581 & n5052;
  assign n5054 = ~n4581 & ~n5052;
  assign n5055 = ~n5053 & ~n5054;
  assign n5056 = ~n5051 & ~n5055;
  assign n5057 = ~n5050 & ~n5056;
  assign n5058 = ~n5038 & n5057;
  assign n5059 = ~n5037 & ~n5058;
  assign n5060 = ~n5028 & n5059;
  assign n5061 = ~n5027 & ~n5060;
  assign n5062 = ~n5018 & ~n5061;
  assign n5063 = ~n5017 & ~n5062;
  assign n5064 = n4781 & ~n5012;
  assign n5065 = ~n5011 & ~n5064;
  assign n5066 = n5063 & ~n5065;
  assign n5067 = ~n5063 & n5065;
  assign n5068 = n4546 & n4587;
  assign n5069 = ~n4546 & ~n4587;
  assign n5070 = ~n4358 & ~n5069;
  assign n5071 = ~n5068 & ~n5070;
  assign n5072 = ~n5067 & ~n5071;
  assign n5073 = ~n5066 & ~n5072;
  assign n5074 = ~n5066 & ~n5067;
  assign n5075 = ~n5071 & ~n5074;
  assign n5076 = n5071 & n5074;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = ~n4163 & n4165;
  assign n5079 = n4163 & ~n4165;
  assign n5080 = ~n5078 & ~n5079;
  assign n5081 = n4169 & n5080;
  assign n5082 = ~n4169 & ~n5080;
  assign n5083 = ~n5081 & ~n5082;
  assign n5084 = n5077 & ~n5083;
  assign n5085 = ~n5077 & n5083;
  assign n5086 = ~n4117 & ~n4118;
  assign n5087 = ~n4161 & n5086;
  assign n5088 = n4161 & ~n5086;
  assign n5089 = ~n5087 & ~n5088;
  assign n5090 = ~n5017 & ~n5018;
  assign n5091 = ~n5061 & n5090;
  assign n5092 = n5061 & ~n5090;
  assign n5093 = ~n5091 & ~n5092;
  assign n5094 = ~n5089 & ~n5093;
  assign n5095 = n5089 & n5093;
  assign n5096 = ~n5027 & ~n5028;
  assign n5097 = n5059 & n5096;
  assign n5098 = ~n5059 & ~n5096;
  assign n5099 = ~n5097 & ~n5098;
  assign n5100 = ~n4127 & ~n4128;
  assign n5101 = n4159 & n5100;
  assign n5102 = ~n4159 & ~n5100;
  assign n5103 = ~n5101 & ~n5102;
  assign n5104 = ~n5099 & ~n5103;
  assign n5105 = n5099 & n5103;
  assign n5106 = ~n4137 & ~n4138;
  assign n5107 = ~n4157 & n5106;
  assign n5108 = n4157 & ~n5106;
  assign n5109 = ~n5107 & ~n5108;
  assign n5110 = ~n5037 & ~n5038;
  assign n5111 = ~n5057 & n5110;
  assign n5112 = n5057 & ~n5110;
  assign n5113 = ~n5111 & ~n5112;
  assign n5114 = ~n5109 & ~n5113;
  assign n5115 = n5109 & n5113;
  assign n5116 = n5041 & n5044;
  assign n5117 = ~n5045 & ~n5116;
  assign n5118 = n4141 & n4144;
  assign n5119 = ~n4145 & ~n5118;
  assign n5120 = n5117 & n5119;
  assign n5121 = ~n5050 & ~n5051;
  assign n5122 = n5055 & n5121;
  assign n5123 = ~n5055 & ~n5121;
  assign n5124 = ~n5122 & ~n5123;
  assign n5125 = n5120 & ~n5124;
  assign n5126 = ~n5120 & n5124;
  assign n5127 = ~n4150 & ~n4151;
  assign n5128 = n4155 & n5127;
  assign n5129 = ~n4155 & ~n5127;
  assign n5130 = ~n5128 & ~n5129;
  assign n5131 = ~n5126 & ~n5130;
  assign n5132 = ~n5125 & ~n5131;
  assign n5133 = ~n5115 & n5132;
  assign n5134 = ~n5114 & ~n5133;
  assign n5135 = ~n5105 & ~n5134;
  assign n5136 = ~n5104 & ~n5135;
  assign n5137 = ~n5095 & ~n5136;
  assign n5138 = ~n5094 & ~n5137;
  assign n5139 = ~n5085 & n5138;
  assign n5140 = ~n5084 & ~n5139;
  assign n5141 = ~n5073 & n5140;
  assign n5142 = n5073 & ~n5140;
  assign n5143 = ~n5141 & ~n5142;
  assign n5144 = n4171 & n5143;
  assign n5145 = ~n4171 & ~n5143;
  assign n5146 = ~n5144 & ~n5145;
  assign n5147 = ~pi277  & pi278 ;
  assign n5148 = pi277  & ~pi278 ;
  assign n5149 = pi279  & ~n5147;
  assign n5150 = ~n5148 & n5149;
  assign n5151 = ~n5147 & ~n5148;
  assign n5152 = ~pi279  & ~n5151;
  assign n5153 = ~n5150 & ~n5152;
  assign n5154 = ~pi280  & pi281 ;
  assign n5155 = pi280  & ~pi281 ;
  assign n5156 = pi282  & ~n5154;
  assign n5157 = ~n5155 & n5156;
  assign n5158 = ~n5154 & ~n5155;
  assign n5159 = ~pi282  & ~n5158;
  assign n5160 = ~n5157 & ~n5159;
  assign n5161 = ~n5153 & n5160;
  assign n5162 = n5153 & ~n5160;
  assign n5163 = ~n5161 & ~n5162;
  assign n5164 = ~pi271  & pi272 ;
  assign n5165 = pi271  & ~pi272 ;
  assign n5166 = pi273  & ~n5164;
  assign n5167 = ~n5165 & n5166;
  assign n5168 = ~n5164 & ~n5165;
  assign n5169 = ~pi273  & ~n5168;
  assign n5170 = ~n5167 & ~n5169;
  assign n5171 = ~pi274  & pi275 ;
  assign n5172 = pi274  & ~pi275 ;
  assign n5173 = pi276  & ~n5171;
  assign n5174 = ~n5172 & n5173;
  assign n5175 = ~n5171 & ~n5172;
  assign n5176 = ~pi276  & ~n5175;
  assign n5177 = ~n5174 & ~n5176;
  assign n5178 = ~n5170 & n5177;
  assign n5179 = n5170 & ~n5177;
  assign n5180 = ~n5178 & ~n5179;
  assign n5181 = ~n5163 & ~n5180;
  assign n5182 = pi280  & pi281 ;
  assign n5183 = pi282  & ~n5158;
  assign n5184 = ~n5182 & ~n5183;
  assign n5185 = pi277  & pi278 ;
  assign n5186 = pi279  & ~n5151;
  assign n5187 = ~n5185 & ~n5186;
  assign n5188 = ~n5184 & ~n5187;
  assign n5189 = ~n5163 & n5188;
  assign n5190 = ~n5153 & ~n5160;
  assign n5191 = n5184 & n5187;
  assign n5192 = ~n5188 & ~n5191;
  assign n5193 = n5190 & n5192;
  assign n5194 = ~n5190 & ~n5192;
  assign n5195 = ~n5189 & ~n5193;
  assign n5196 = ~n5194 & n5195;
  assign n5197 = n5181 & n5196;
  assign n5198 = ~n5181 & ~n5196;
  assign n5199 = pi274  & pi275 ;
  assign n5200 = pi276  & ~n5175;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = pi271  & pi272 ;
  assign n5203 = pi273  & ~n5168;
  assign n5204 = ~n5202 & ~n5203;
  assign n5205 = ~n5201 & n5204;
  assign n5206 = n5201 & ~n5204;
  assign n5207 = ~n5205 & ~n5206;
  assign n5208 = ~n5170 & ~n5177;
  assign n5209 = n5207 & n5208;
  assign n5210 = ~n5207 & ~n5208;
  assign n5211 = ~n5209 & ~n5210;
  assign n5212 = ~n5198 & ~n5211;
  assign n5213 = ~n5197 & ~n5212;
  assign n5214 = n5190 & ~n5191;
  assign n5215 = ~n5188 & ~n5214;
  assign n5216 = ~n5213 & ~n5215;
  assign n5217 = n5213 & n5215;
  assign n5218 = ~n5216 & ~n5217;
  assign n5219 = ~n5201 & n5208;
  assign n5220 = n5204 & ~n5219;
  assign n5221 = n5201 & ~n5208;
  assign n5222 = ~n5220 & ~n5221;
  assign n5223 = ~n5218 & n5222;
  assign n5224 = n5218 & ~n5222;
  assign n5225 = ~n5223 & ~n5224;
  assign n5226 = ~pi289  & pi290 ;
  assign n5227 = pi289  & ~pi290 ;
  assign n5228 = pi291  & ~n5226;
  assign n5229 = ~n5227 & n5228;
  assign n5230 = ~n5226 & ~n5227;
  assign n5231 = ~pi291  & ~n5230;
  assign n5232 = ~n5229 & ~n5231;
  assign n5233 = ~pi292  & pi293 ;
  assign n5234 = pi292  & ~pi293 ;
  assign n5235 = pi294  & ~n5233;
  assign n5236 = ~n5234 & n5235;
  assign n5237 = ~n5233 & ~n5234;
  assign n5238 = ~pi294  & ~n5237;
  assign n5239 = ~n5236 & ~n5238;
  assign n5240 = ~n5232 & n5239;
  assign n5241 = n5232 & ~n5239;
  assign n5242 = ~n5240 & ~n5241;
  assign n5243 = ~pi283  & pi284 ;
  assign n5244 = pi283  & ~pi284 ;
  assign n5245 = pi285  & ~n5243;
  assign n5246 = ~n5244 & n5245;
  assign n5247 = ~n5243 & ~n5244;
  assign n5248 = ~pi285  & ~n5247;
  assign n5249 = ~n5246 & ~n5248;
  assign n5250 = ~pi286  & pi287 ;
  assign n5251 = pi286  & ~pi287 ;
  assign n5252 = pi288  & ~n5250;
  assign n5253 = ~n5251 & n5252;
  assign n5254 = ~n5250 & ~n5251;
  assign n5255 = ~pi288  & ~n5254;
  assign n5256 = ~n5253 & ~n5255;
  assign n5257 = ~n5249 & n5256;
  assign n5258 = n5249 & ~n5256;
  assign n5259 = ~n5257 & ~n5258;
  assign n5260 = ~n5242 & ~n5259;
  assign n5261 = pi292  & pi293 ;
  assign n5262 = pi294  & ~n5237;
  assign n5263 = ~n5261 & ~n5262;
  assign n5264 = pi289  & pi290 ;
  assign n5265 = pi291  & ~n5230;
  assign n5266 = ~n5264 & ~n5265;
  assign n5267 = n5263 & ~n5266;
  assign n5268 = ~n5263 & n5266;
  assign n5269 = ~n5267 & ~n5268;
  assign n5270 = n5260 & ~n5269;
  assign n5271 = ~n5232 & ~n5239;
  assign n5272 = n5269 & n5271;
  assign n5273 = ~n5269 & ~n5271;
  assign n5274 = ~n5260 & ~n5272;
  assign n5275 = ~n5273 & n5274;
  assign n5276 = pi286  & pi287 ;
  assign n5277 = pi288  & ~n5254;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = pi283  & pi284 ;
  assign n5280 = pi285  & ~n5247;
  assign n5281 = ~n5279 & ~n5280;
  assign n5282 = ~n5278 & ~n5281;
  assign n5283 = ~n5259 & n5282;
  assign n5284 = ~n5249 & ~n5256;
  assign n5285 = n5278 & n5281;
  assign n5286 = ~n5282 & ~n5285;
  assign n5287 = n5284 & n5286;
  assign n5288 = ~n5284 & ~n5286;
  assign n5289 = ~n5283 & ~n5287;
  assign n5290 = ~n5288 & n5289;
  assign n5291 = ~n5275 & n5290;
  assign n5292 = ~n5270 & ~n5291;
  assign n5293 = ~n5263 & n5271;
  assign n5294 = n5266 & ~n5293;
  assign n5295 = n5263 & ~n5271;
  assign n5296 = ~n5294 & ~n5295;
  assign n5297 = ~n5292 & n5296;
  assign n5298 = n5292 & ~n5296;
  assign n5299 = ~n5297 & ~n5298;
  assign n5300 = n5284 & ~n5285;
  assign n5301 = ~n5282 & ~n5300;
  assign n5302 = n5299 & ~n5301;
  assign n5303 = ~n5299 & n5301;
  assign n5304 = ~n5302 & ~n5303;
  assign n5305 = n5225 & ~n5304;
  assign n5306 = ~n5225 & n5304;
  assign n5307 = n5242 & n5259;
  assign n5308 = ~n5260 & ~n5307;
  assign n5309 = n5163 & n5180;
  assign n5310 = ~n5181 & ~n5309;
  assign n5311 = n5308 & n5310;
  assign n5312 = ~n5270 & ~n5275;
  assign n5313 = n5290 & n5312;
  assign n5314 = ~n5290 & ~n5312;
  assign n5315 = ~n5313 & ~n5314;
  assign n5316 = n5311 & n5315;
  assign n5317 = ~n5311 & ~n5315;
  assign n5318 = ~n5197 & ~n5198;
  assign n5319 = ~n5211 & n5318;
  assign n5320 = n5211 & ~n5318;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = ~n5317 & n5321;
  assign n5323 = ~n5316 & ~n5322;
  assign n5324 = ~n5306 & n5323;
  assign n5325 = ~n5305 & ~n5324;
  assign n5326 = ~n5298 & ~n5301;
  assign n5327 = ~n5297 & ~n5326;
  assign n5328 = ~n5325 & n5327;
  assign n5329 = n5325 & ~n5327;
  assign n5330 = ~n5217 & n5222;
  assign n5331 = ~n5216 & ~n5330;
  assign n5332 = ~n5329 & n5331;
  assign n5333 = ~n5328 & ~n5332;
  assign n5334 = ~pi301  & pi302 ;
  assign n5335 = pi301  & ~pi302 ;
  assign n5336 = pi303  & ~n5334;
  assign n5337 = ~n5335 & n5336;
  assign n5338 = ~n5334 & ~n5335;
  assign n5339 = ~pi303  & ~n5338;
  assign n5340 = ~n5337 & ~n5339;
  assign n5341 = ~pi304  & pi305 ;
  assign n5342 = pi304  & ~pi305 ;
  assign n5343 = pi306  & ~n5341;
  assign n5344 = ~n5342 & n5343;
  assign n5345 = ~n5341 & ~n5342;
  assign n5346 = ~pi306  & ~n5345;
  assign n5347 = ~n5344 & ~n5346;
  assign n5348 = ~n5340 & n5347;
  assign n5349 = n5340 & ~n5347;
  assign n5350 = ~n5348 & ~n5349;
  assign n5351 = ~pi295  & pi296 ;
  assign n5352 = pi295  & ~pi296 ;
  assign n5353 = pi297  & ~n5351;
  assign n5354 = ~n5352 & n5353;
  assign n5355 = ~n5351 & ~n5352;
  assign n5356 = ~pi297  & ~n5355;
  assign n5357 = ~n5354 & ~n5356;
  assign n5358 = ~pi298  & pi299 ;
  assign n5359 = pi298  & ~pi299 ;
  assign n5360 = pi300  & ~n5358;
  assign n5361 = ~n5359 & n5360;
  assign n5362 = ~n5358 & ~n5359;
  assign n5363 = ~pi300  & ~n5362;
  assign n5364 = ~n5361 & ~n5363;
  assign n5365 = ~n5357 & n5364;
  assign n5366 = n5357 & ~n5364;
  assign n5367 = ~n5365 & ~n5366;
  assign n5368 = ~n5350 & ~n5367;
  assign n5369 = pi304  & pi305 ;
  assign n5370 = pi306  & ~n5345;
  assign n5371 = ~n5369 & ~n5370;
  assign n5372 = pi301  & pi302 ;
  assign n5373 = pi303  & ~n5338;
  assign n5374 = ~n5372 & ~n5373;
  assign n5375 = ~n5371 & ~n5374;
  assign n5376 = ~n5350 & n5375;
  assign n5377 = ~n5340 & ~n5347;
  assign n5378 = n5371 & n5374;
  assign n5379 = ~n5375 & ~n5378;
  assign n5380 = n5377 & n5379;
  assign n5381 = ~n5377 & ~n5379;
  assign n5382 = ~n5376 & ~n5380;
  assign n5383 = ~n5381 & n5382;
  assign n5384 = n5368 & n5383;
  assign n5385 = ~n5368 & ~n5383;
  assign n5386 = pi298  & pi299 ;
  assign n5387 = pi300  & ~n5362;
  assign n5388 = ~n5386 & ~n5387;
  assign n5389 = pi295  & pi296 ;
  assign n5390 = pi297  & ~n5355;
  assign n5391 = ~n5389 & ~n5390;
  assign n5392 = ~n5388 & n5391;
  assign n5393 = n5388 & ~n5391;
  assign n5394 = ~n5392 & ~n5393;
  assign n5395 = ~n5357 & ~n5364;
  assign n5396 = n5394 & n5395;
  assign n5397 = ~n5394 & ~n5395;
  assign n5398 = ~n5396 & ~n5397;
  assign n5399 = ~n5385 & ~n5398;
  assign n5400 = ~n5384 & ~n5399;
  assign n5401 = n5377 & ~n5378;
  assign n5402 = ~n5375 & ~n5401;
  assign n5403 = ~n5400 & ~n5402;
  assign n5404 = n5400 & n5402;
  assign n5405 = ~n5403 & ~n5404;
  assign n5406 = ~n5388 & n5395;
  assign n5407 = n5391 & ~n5406;
  assign n5408 = n5388 & ~n5395;
  assign n5409 = ~n5407 & ~n5408;
  assign n5410 = ~n5405 & n5409;
  assign n5411 = n5405 & ~n5409;
  assign n5412 = ~n5410 & ~n5411;
  assign n5413 = ~pi313  & pi314 ;
  assign n5414 = pi313  & ~pi314 ;
  assign n5415 = pi315  & ~n5413;
  assign n5416 = ~n5414 & n5415;
  assign n5417 = ~n5413 & ~n5414;
  assign n5418 = ~pi315  & ~n5417;
  assign n5419 = ~n5416 & ~n5418;
  assign n5420 = ~pi316  & pi317 ;
  assign n5421 = pi316  & ~pi317 ;
  assign n5422 = pi318  & ~n5420;
  assign n5423 = ~n5421 & n5422;
  assign n5424 = ~n5420 & ~n5421;
  assign n5425 = ~pi318  & ~n5424;
  assign n5426 = ~n5423 & ~n5425;
  assign n5427 = ~n5419 & n5426;
  assign n5428 = n5419 & ~n5426;
  assign n5429 = ~n5427 & ~n5428;
  assign n5430 = ~pi307  & pi308 ;
  assign n5431 = pi307  & ~pi308 ;
  assign n5432 = pi309  & ~n5430;
  assign n5433 = ~n5431 & n5432;
  assign n5434 = ~n5430 & ~n5431;
  assign n5435 = ~pi309  & ~n5434;
  assign n5436 = ~n5433 & ~n5435;
  assign n5437 = ~pi310  & pi311 ;
  assign n5438 = pi310  & ~pi311 ;
  assign n5439 = pi312  & ~n5437;
  assign n5440 = ~n5438 & n5439;
  assign n5441 = ~n5437 & ~n5438;
  assign n5442 = ~pi312  & ~n5441;
  assign n5443 = ~n5440 & ~n5442;
  assign n5444 = ~n5436 & n5443;
  assign n5445 = n5436 & ~n5443;
  assign n5446 = ~n5444 & ~n5445;
  assign n5447 = ~n5429 & ~n5446;
  assign n5448 = pi316  & pi317 ;
  assign n5449 = pi318  & ~n5424;
  assign n5450 = ~n5448 & ~n5449;
  assign n5451 = pi313  & pi314 ;
  assign n5452 = pi315  & ~n5417;
  assign n5453 = ~n5451 & ~n5452;
  assign n5454 = n5450 & ~n5453;
  assign n5455 = ~n5450 & n5453;
  assign n5456 = ~n5454 & ~n5455;
  assign n5457 = n5447 & ~n5456;
  assign n5458 = ~n5419 & ~n5426;
  assign n5459 = n5456 & n5458;
  assign n5460 = ~n5456 & ~n5458;
  assign n5461 = ~n5447 & ~n5459;
  assign n5462 = ~n5460 & n5461;
  assign n5463 = pi310  & pi311 ;
  assign n5464 = pi312  & ~n5441;
  assign n5465 = ~n5463 & ~n5464;
  assign n5466 = pi307  & pi308 ;
  assign n5467 = pi309  & ~n5434;
  assign n5468 = ~n5466 & ~n5467;
  assign n5469 = ~n5465 & ~n5468;
  assign n5470 = ~n5446 & n5469;
  assign n5471 = ~n5436 & ~n5443;
  assign n5472 = n5465 & n5468;
  assign n5473 = ~n5469 & ~n5472;
  assign n5474 = n5471 & n5473;
  assign n5475 = ~n5471 & ~n5473;
  assign n5476 = ~n5470 & ~n5474;
  assign n5477 = ~n5475 & n5476;
  assign n5478 = ~n5462 & n5477;
  assign n5479 = ~n5457 & ~n5478;
  assign n5480 = ~n5450 & n5458;
  assign n5481 = n5453 & ~n5480;
  assign n5482 = n5450 & ~n5458;
  assign n5483 = ~n5481 & ~n5482;
  assign n5484 = ~n5479 & n5483;
  assign n5485 = n5479 & ~n5483;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = n5471 & ~n5472;
  assign n5488 = ~n5469 & ~n5487;
  assign n5489 = n5486 & ~n5488;
  assign n5490 = ~n5486 & n5488;
  assign n5491 = ~n5489 & ~n5490;
  assign n5492 = n5412 & ~n5491;
  assign n5493 = ~n5412 & n5491;
  assign n5494 = n5429 & n5446;
  assign n5495 = ~n5447 & ~n5494;
  assign n5496 = n5350 & n5367;
  assign n5497 = ~n5368 & ~n5496;
  assign n5498 = n5495 & n5497;
  assign n5499 = ~n5457 & ~n5462;
  assign n5500 = n5477 & n5499;
  assign n5501 = ~n5477 & ~n5499;
  assign n5502 = ~n5500 & ~n5501;
  assign n5503 = n5498 & n5502;
  assign n5504 = ~n5498 & ~n5502;
  assign n5505 = ~n5384 & ~n5385;
  assign n5506 = ~n5398 & n5505;
  assign n5507 = n5398 & ~n5505;
  assign n5508 = ~n5506 & ~n5507;
  assign n5509 = ~n5504 & n5508;
  assign n5510 = ~n5503 & ~n5509;
  assign n5511 = ~n5493 & n5510;
  assign n5512 = ~n5492 & ~n5511;
  assign n5513 = ~n5485 & ~n5488;
  assign n5514 = ~n5484 & ~n5513;
  assign n5515 = ~n5512 & n5514;
  assign n5516 = n5512 & ~n5514;
  assign n5517 = ~n5404 & n5409;
  assign n5518 = ~n5403 & ~n5517;
  assign n5519 = ~n5516 & n5518;
  assign n5520 = ~n5515 & ~n5519;
  assign n5521 = ~n5515 & ~n5516;
  assign n5522 = n5518 & n5521;
  assign n5523 = ~n5518 & ~n5521;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = ~n5328 & ~n5329;
  assign n5526 = n5331 & n5525;
  assign n5527 = ~n5331 & ~n5525;
  assign n5528 = ~n5526 & ~n5527;
  assign n5529 = ~n5524 & ~n5528;
  assign n5530 = n5524 & n5528;
  assign n5531 = ~n5305 & ~n5306;
  assign n5532 = ~n5323 & n5531;
  assign n5533 = n5323 & ~n5531;
  assign n5534 = ~n5532 & ~n5533;
  assign n5535 = ~n5492 & ~n5493;
  assign n5536 = ~n5510 & n5535;
  assign n5537 = n5510 & ~n5535;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = ~n5534 & ~n5538;
  assign n5540 = n5534 & n5538;
  assign n5541 = ~n5495 & ~n5497;
  assign n5542 = ~n5498 & ~n5541;
  assign n5543 = ~n5308 & ~n5310;
  assign n5544 = ~n5311 & ~n5543;
  assign n5545 = n5542 & n5544;
  assign n5546 = ~n5503 & ~n5504;
  assign n5547 = ~n5508 & n5546;
  assign n5548 = n5508 & ~n5546;
  assign n5549 = ~n5547 & ~n5548;
  assign n5550 = n5545 & ~n5549;
  assign n5551 = ~n5545 & n5549;
  assign n5552 = ~n5316 & ~n5317;
  assign n5553 = ~n5321 & n5552;
  assign n5554 = n5321 & ~n5552;
  assign n5555 = ~n5553 & ~n5554;
  assign n5556 = ~n5551 & ~n5555;
  assign n5557 = ~n5550 & ~n5556;
  assign n5558 = ~n5540 & n5557;
  assign n5559 = ~n5539 & ~n5558;
  assign n5560 = ~n5530 & n5559;
  assign n5561 = ~n5529 & ~n5560;
  assign n5562 = ~n5520 & n5561;
  assign n5563 = n5520 & ~n5561;
  assign n5564 = ~n5562 & ~n5563;
  assign n5565 = n5333 & n5564;
  assign n5566 = ~n5333 & ~n5564;
  assign n5567 = ~n5565 & ~n5566;
  assign n5568 = ~pi325  & pi326 ;
  assign n5569 = pi325  & ~pi326 ;
  assign n5570 = pi327  & ~n5568;
  assign n5571 = ~n5569 & n5570;
  assign n5572 = ~n5568 & ~n5569;
  assign n5573 = ~pi327  & ~n5572;
  assign n5574 = ~n5571 & ~n5573;
  assign n5575 = ~pi328  & pi329 ;
  assign n5576 = pi328  & ~pi329 ;
  assign n5577 = pi330  & ~n5575;
  assign n5578 = ~n5576 & n5577;
  assign n5579 = ~n5575 & ~n5576;
  assign n5580 = ~pi330  & ~n5579;
  assign n5581 = ~n5578 & ~n5580;
  assign n5582 = ~n5574 & n5581;
  assign n5583 = n5574 & ~n5581;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = ~pi319  & pi320 ;
  assign n5586 = pi319  & ~pi320 ;
  assign n5587 = pi321  & ~n5585;
  assign n5588 = ~n5586 & n5587;
  assign n5589 = ~n5585 & ~n5586;
  assign n5590 = ~pi321  & ~n5589;
  assign n5591 = ~n5588 & ~n5590;
  assign n5592 = ~pi322  & pi323 ;
  assign n5593 = pi322  & ~pi323 ;
  assign n5594 = pi324  & ~n5592;
  assign n5595 = ~n5593 & n5594;
  assign n5596 = ~n5592 & ~n5593;
  assign n5597 = ~pi324  & ~n5596;
  assign n5598 = ~n5595 & ~n5597;
  assign n5599 = ~n5591 & n5598;
  assign n5600 = n5591 & ~n5598;
  assign n5601 = ~n5599 & ~n5600;
  assign n5602 = ~n5584 & ~n5601;
  assign n5603 = pi328  & pi329 ;
  assign n5604 = pi330  & ~n5579;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = pi325  & pi326 ;
  assign n5607 = pi327  & ~n5572;
  assign n5608 = ~n5606 & ~n5607;
  assign n5609 = ~n5605 & ~n5608;
  assign n5610 = ~n5584 & n5609;
  assign n5611 = ~n5574 & ~n5581;
  assign n5612 = n5605 & n5608;
  assign n5613 = ~n5609 & ~n5612;
  assign n5614 = n5611 & n5613;
  assign n5615 = ~n5611 & ~n5613;
  assign n5616 = ~n5610 & ~n5614;
  assign n5617 = ~n5615 & n5616;
  assign n5618 = n5602 & n5617;
  assign n5619 = ~n5602 & ~n5617;
  assign n5620 = pi322  & pi323 ;
  assign n5621 = pi324  & ~n5596;
  assign n5622 = ~n5620 & ~n5621;
  assign n5623 = pi319  & pi320 ;
  assign n5624 = pi321  & ~n5589;
  assign n5625 = ~n5623 & ~n5624;
  assign n5626 = ~n5622 & n5625;
  assign n5627 = n5622 & ~n5625;
  assign n5628 = ~n5626 & ~n5627;
  assign n5629 = ~n5591 & ~n5598;
  assign n5630 = n5628 & n5629;
  assign n5631 = ~n5628 & ~n5629;
  assign n5632 = ~n5630 & ~n5631;
  assign n5633 = ~n5619 & ~n5632;
  assign n5634 = ~n5618 & ~n5633;
  assign n5635 = n5611 & ~n5612;
  assign n5636 = ~n5609 & ~n5635;
  assign n5637 = ~n5634 & ~n5636;
  assign n5638 = n5634 & n5636;
  assign n5639 = ~n5637 & ~n5638;
  assign n5640 = ~n5622 & n5629;
  assign n5641 = n5625 & ~n5640;
  assign n5642 = n5622 & ~n5629;
  assign n5643 = ~n5641 & ~n5642;
  assign n5644 = ~n5639 & n5643;
  assign n5645 = n5639 & ~n5643;
  assign n5646 = ~n5644 & ~n5645;
  assign n5647 = pi337  & ~pi338 ;
  assign n5648 = ~pi337  & pi338 ;
  assign n5649 = pi339  & ~n5647;
  assign n5650 = ~n5648 & n5649;
  assign n5651 = ~n5647 & ~n5648;
  assign n5652 = ~pi339  & ~n5651;
  assign n5653 = ~n5650 & ~n5652;
  assign n5654 = pi340  & ~pi341 ;
  assign n5655 = ~pi340  & pi341 ;
  assign n5656 = pi342  & ~n5654;
  assign n5657 = ~n5655 & n5656;
  assign n5658 = ~n5654 & ~n5655;
  assign n5659 = ~pi342  & ~n5658;
  assign n5660 = ~n5657 & ~n5659;
  assign n5661 = ~n5653 & n5660;
  assign n5662 = n5653 & ~n5660;
  assign n5663 = ~n5661 & ~n5662;
  assign n5664 = pi340  & pi341 ;
  assign n5665 = pi342  & ~n5658;
  assign n5666 = ~n5664 & ~n5665;
  assign n5667 = pi337  & pi338 ;
  assign n5668 = pi339  & ~n5651;
  assign n5669 = ~n5667 & ~n5668;
  assign n5670 = ~n5666 & ~n5669;
  assign n5671 = ~n5663 & n5670;
  assign n5672 = ~n5653 & ~n5660;
  assign n5673 = n5666 & n5669;
  assign n5674 = ~n5670 & ~n5673;
  assign n5675 = n5672 & n5674;
  assign n5676 = ~n5672 & ~n5674;
  assign n5677 = ~n5671 & ~n5675;
  assign n5678 = ~n5676 & n5677;
  assign n5679 = pi331  & ~pi332 ;
  assign n5680 = ~pi331  & pi332 ;
  assign n5681 = pi333  & ~n5679;
  assign n5682 = ~n5680 & n5681;
  assign n5683 = ~n5679 & ~n5680;
  assign n5684 = ~pi333  & ~n5683;
  assign n5685 = ~n5682 & ~n5684;
  assign n5686 = pi334  & ~pi335 ;
  assign n5687 = ~pi334  & pi335 ;
  assign n5688 = pi336  & ~n5686;
  assign n5689 = ~n5687 & n5688;
  assign n5690 = ~n5686 & ~n5687;
  assign n5691 = ~pi336  & ~n5690;
  assign n5692 = ~n5689 & ~n5691;
  assign n5693 = ~n5685 & n5692;
  assign n5694 = n5685 & ~n5692;
  assign n5695 = ~n5693 & ~n5694;
  assign n5696 = ~n5663 & ~n5695;
  assign n5697 = ~n5685 & ~n5692;
  assign n5698 = pi334  & pi335 ;
  assign n5699 = pi336  & ~n5690;
  assign n5700 = ~n5698 & ~n5699;
  assign n5701 = pi331  & pi332 ;
  assign n5702 = pi333  & ~n5683;
  assign n5703 = ~n5701 & ~n5702;
  assign n5704 = n5700 & ~n5703;
  assign n5705 = ~n5700 & n5703;
  assign n5706 = ~n5704 & ~n5705;
  assign n5707 = n5697 & n5706;
  assign n5708 = ~n5697 & ~n5706;
  assign n5709 = ~n5707 & ~n5708;
  assign n5710 = ~n5696 & n5709;
  assign n5711 = n5678 & ~n5710;
  assign n5712 = n5696 & ~n5709;
  assign n5713 = ~n5711 & ~n5712;
  assign n5714 = n5672 & ~n5673;
  assign n5715 = ~n5670 & ~n5714;
  assign n5716 = ~n5713 & ~n5715;
  assign n5717 = n5713 & n5715;
  assign n5718 = ~n5716 & ~n5717;
  assign n5719 = n5697 & ~n5700;
  assign n5720 = n5703 & ~n5719;
  assign n5721 = ~n5697 & n5700;
  assign n5722 = ~n5720 & ~n5721;
  assign n5723 = ~n5718 & n5722;
  assign n5724 = n5718 & ~n5722;
  assign n5725 = ~n5723 & ~n5724;
  assign n5726 = ~n5646 & ~n5725;
  assign n5727 = n5646 & n5725;
  assign n5728 = n5663 & n5695;
  assign n5729 = ~n5696 & ~n5728;
  assign n5730 = n5584 & n5601;
  assign n5731 = ~n5602 & ~n5730;
  assign n5732 = n5729 & n5731;
  assign n5733 = n5696 & ~n5706;
  assign n5734 = ~n5710 & ~n5733;
  assign n5735 = n5678 & ~n5734;
  assign n5736 = ~n5678 & n5734;
  assign n5737 = ~n5735 & ~n5736;
  assign n5738 = n5732 & ~n5737;
  assign n5739 = ~n5732 & n5737;
  assign n5740 = ~n5618 & ~n5619;
  assign n5741 = ~n5632 & n5740;
  assign n5742 = n5632 & ~n5740;
  assign n5743 = ~n5741 & ~n5742;
  assign n5744 = ~n5739 & n5743;
  assign n5745 = ~n5738 & ~n5744;
  assign n5746 = ~n5727 & ~n5745;
  assign n5747 = ~n5726 & ~n5746;
  assign n5748 = ~n5717 & n5722;
  assign n5749 = ~n5716 & ~n5748;
  assign n5750 = ~n5747 & ~n5749;
  assign n5751 = n5747 & n5749;
  assign n5752 = ~n5638 & n5643;
  assign n5753 = ~n5637 & ~n5752;
  assign n5754 = ~n5751 & ~n5753;
  assign n5755 = ~n5750 & ~n5754;
  assign n5756 = pi343  & ~pi344 ;
  assign n5757 = ~pi343  & pi344 ;
  assign n5758 = pi345  & ~n5756;
  assign n5759 = ~n5757 & n5758;
  assign n5760 = ~n5756 & ~n5757;
  assign n5761 = ~pi345  & ~n5760;
  assign n5762 = ~n5759 & ~n5761;
  assign n5763 = pi346  & ~pi347 ;
  assign n5764 = ~pi346  & pi347 ;
  assign n5765 = pi348  & ~n5763;
  assign n5766 = ~n5764 & n5765;
  assign n5767 = ~n5763 & ~n5764;
  assign n5768 = ~pi348  & ~n5767;
  assign n5769 = ~n5766 & ~n5768;
  assign n5770 = ~n5762 & n5769;
  assign n5771 = n5762 & ~n5769;
  assign n5772 = ~n5770 & ~n5771;
  assign n5773 = pi349  & ~pi350 ;
  assign n5774 = ~pi349  & pi350 ;
  assign n5775 = pi351  & ~n5773;
  assign n5776 = ~n5774 & n5775;
  assign n5777 = ~n5773 & ~n5774;
  assign n5778 = ~pi351  & ~n5777;
  assign n5779 = ~n5776 & ~n5778;
  assign n5780 = pi352  & ~pi353 ;
  assign n5781 = ~pi352  & pi353 ;
  assign n5782 = pi354  & ~n5780;
  assign n5783 = ~n5781 & n5782;
  assign n5784 = ~n5780 & ~n5781;
  assign n5785 = ~pi354  & ~n5784;
  assign n5786 = ~n5783 & ~n5785;
  assign n5787 = ~n5779 & n5786;
  assign n5788 = n5779 & ~n5786;
  assign n5789 = ~n5787 & ~n5788;
  assign n5790 = ~n5772 & ~n5789;
  assign n5791 = pi352  & pi353 ;
  assign n5792 = pi354  & ~n5784;
  assign n5793 = ~n5791 & ~n5792;
  assign n5794 = pi349  & pi350 ;
  assign n5795 = pi351  & ~n5777;
  assign n5796 = ~n5794 & ~n5795;
  assign n5797 = ~n5793 & ~n5796;
  assign n5798 = ~n5789 & n5797;
  assign n5799 = ~n5779 & ~n5786;
  assign n5800 = n5793 & n5796;
  assign n5801 = ~n5797 & ~n5800;
  assign n5802 = n5799 & n5801;
  assign n5803 = ~n5799 & ~n5801;
  assign n5804 = ~n5798 & ~n5802;
  assign n5805 = ~n5803 & n5804;
  assign n5806 = n5790 & n5805;
  assign n5807 = ~n5790 & ~n5805;
  assign n5808 = ~n5762 & ~n5769;
  assign n5809 = pi346  & pi347 ;
  assign n5810 = pi348  & ~n5767;
  assign n5811 = ~n5809 & ~n5810;
  assign n5812 = pi343  & pi344 ;
  assign n5813 = pi345  & ~n5760;
  assign n5814 = ~n5812 & ~n5813;
  assign n5815 = n5811 & ~n5814;
  assign n5816 = ~n5811 & n5814;
  assign n5817 = ~n5815 & ~n5816;
  assign n5818 = n5808 & n5817;
  assign n5819 = ~n5808 & ~n5817;
  assign n5820 = ~n5818 & ~n5819;
  assign n5821 = ~n5807 & ~n5820;
  assign n5822 = ~n5806 & ~n5821;
  assign n5823 = n5799 & ~n5800;
  assign n5824 = ~n5797 & ~n5823;
  assign n5825 = ~n5822 & ~n5824;
  assign n5826 = n5822 & n5824;
  assign n5827 = ~n5825 & ~n5826;
  assign n5828 = n5808 & ~n5811;
  assign n5829 = n5814 & ~n5828;
  assign n5830 = ~n5808 & n5811;
  assign n5831 = ~n5829 & ~n5830;
  assign n5832 = ~n5827 & n5831;
  assign n5833 = n5827 & ~n5831;
  assign n5834 = ~n5832 & ~n5833;
  assign n5835 = pi361  & ~pi362 ;
  assign n5836 = ~pi361  & pi362 ;
  assign n5837 = pi363  & ~n5835;
  assign n5838 = ~n5836 & n5837;
  assign n5839 = ~n5835 & ~n5836;
  assign n5840 = ~pi363  & ~n5839;
  assign n5841 = ~n5838 & ~n5840;
  assign n5842 = pi364  & ~pi365 ;
  assign n5843 = ~pi364  & pi365 ;
  assign n5844 = pi366  & ~n5842;
  assign n5845 = ~n5843 & n5844;
  assign n5846 = ~n5842 & ~n5843;
  assign n5847 = ~pi366  & ~n5846;
  assign n5848 = ~n5845 & ~n5847;
  assign n5849 = ~n5841 & n5848;
  assign n5850 = n5841 & ~n5848;
  assign n5851 = ~n5849 & ~n5850;
  assign n5852 = pi364  & pi365 ;
  assign n5853 = pi366  & ~n5846;
  assign n5854 = ~n5852 & ~n5853;
  assign n5855 = pi361  & pi362 ;
  assign n5856 = pi363  & ~n5839;
  assign n5857 = ~n5855 & ~n5856;
  assign n5858 = ~n5854 & ~n5857;
  assign n5859 = ~n5851 & n5858;
  assign n5860 = ~n5841 & ~n5848;
  assign n5861 = n5854 & n5857;
  assign n5862 = ~n5858 & ~n5861;
  assign n5863 = n5860 & n5862;
  assign n5864 = ~n5860 & ~n5862;
  assign n5865 = ~n5859 & ~n5863;
  assign n5866 = ~n5864 & n5865;
  assign n5867 = pi355  & ~pi356 ;
  assign n5868 = ~pi355  & pi356 ;
  assign n5869 = pi357  & ~n5867;
  assign n5870 = ~n5868 & n5869;
  assign n5871 = ~n5867 & ~n5868;
  assign n5872 = ~pi357  & ~n5871;
  assign n5873 = ~n5870 & ~n5872;
  assign n5874 = pi358  & ~pi359 ;
  assign n5875 = ~pi358  & pi359 ;
  assign n5876 = pi360  & ~n5874;
  assign n5877 = ~n5875 & n5876;
  assign n5878 = ~n5874 & ~n5875;
  assign n5879 = ~pi360  & ~n5878;
  assign n5880 = ~n5877 & ~n5879;
  assign n5881 = ~n5873 & n5880;
  assign n5882 = n5873 & ~n5880;
  assign n5883 = ~n5881 & ~n5882;
  assign n5884 = ~n5851 & ~n5883;
  assign n5885 = ~n5873 & ~n5880;
  assign n5886 = pi358  & pi359 ;
  assign n5887 = pi360  & ~n5878;
  assign n5888 = ~n5886 & ~n5887;
  assign n5889 = pi355  & pi356 ;
  assign n5890 = pi357  & ~n5871;
  assign n5891 = ~n5889 & ~n5890;
  assign n5892 = n5888 & ~n5891;
  assign n5893 = ~n5888 & n5891;
  assign n5894 = ~n5892 & ~n5893;
  assign n5895 = n5885 & n5894;
  assign n5896 = ~n5885 & ~n5894;
  assign n5897 = ~n5895 & ~n5896;
  assign n5898 = ~n5884 & n5897;
  assign n5899 = n5866 & ~n5898;
  assign n5900 = n5884 & ~n5897;
  assign n5901 = ~n5899 & ~n5900;
  assign n5902 = n5860 & ~n5861;
  assign n5903 = ~n5858 & ~n5902;
  assign n5904 = ~n5901 & ~n5903;
  assign n5905 = n5901 & n5903;
  assign n5906 = ~n5904 & ~n5905;
  assign n5907 = n5885 & ~n5888;
  assign n5908 = n5891 & ~n5907;
  assign n5909 = ~n5885 & n5888;
  assign n5910 = ~n5908 & ~n5909;
  assign n5911 = ~n5906 & n5910;
  assign n5912 = n5906 & ~n5910;
  assign n5913 = ~n5911 & ~n5912;
  assign n5914 = ~n5834 & ~n5913;
  assign n5915 = n5834 & n5913;
  assign n5916 = n5851 & n5883;
  assign n5917 = ~n5884 & ~n5916;
  assign n5918 = n5772 & n5789;
  assign n5919 = ~n5790 & ~n5918;
  assign n5920 = n5917 & n5919;
  assign n5921 = n5884 & ~n5894;
  assign n5922 = ~n5898 & ~n5921;
  assign n5923 = n5866 & ~n5922;
  assign n5924 = ~n5866 & n5922;
  assign n5925 = ~n5923 & ~n5924;
  assign n5926 = n5920 & ~n5925;
  assign n5927 = ~n5920 & n5925;
  assign n5928 = ~n5806 & ~n5807;
  assign n5929 = ~n5820 & n5928;
  assign n5930 = n5820 & ~n5928;
  assign n5931 = ~n5929 & ~n5930;
  assign n5932 = ~n5927 & n5931;
  assign n5933 = ~n5926 & ~n5932;
  assign n5934 = ~n5915 & ~n5933;
  assign n5935 = ~n5914 & ~n5934;
  assign n5936 = ~n5905 & n5910;
  assign n5937 = ~n5904 & ~n5936;
  assign n5938 = ~n5935 & ~n5937;
  assign n5939 = n5935 & n5937;
  assign n5940 = ~n5826 & n5831;
  assign n5941 = ~n5825 & ~n5940;
  assign n5942 = ~n5939 & ~n5941;
  assign n5943 = ~n5938 & ~n5942;
  assign n5944 = ~n5938 & ~n5939;
  assign n5945 = n5941 & ~n5944;
  assign n5946 = ~n5938 & n5942;
  assign n5947 = ~n5945 & ~n5946;
  assign n5948 = ~n5750 & ~n5751;
  assign n5949 = n5753 & ~n5948;
  assign n5950 = ~n5750 & n5754;
  assign n5951 = ~n5949 & ~n5950;
  assign n5952 = ~n5947 & ~n5951;
  assign n5953 = n5947 & n5951;
  assign n5954 = ~n5726 & ~n5727;
  assign n5955 = ~n5745 & n5954;
  assign n5956 = n5745 & ~n5954;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = ~n5914 & ~n5915;
  assign n5959 = ~n5933 & n5958;
  assign n5960 = n5933 & ~n5958;
  assign n5961 = ~n5959 & ~n5960;
  assign n5962 = ~n5957 & ~n5961;
  assign n5963 = n5957 & n5961;
  assign n5964 = ~n5917 & ~n5919;
  assign n5965 = ~n5920 & ~n5964;
  assign n5966 = ~n5729 & ~n5731;
  assign n5967 = ~n5732 & ~n5966;
  assign n5968 = n5965 & n5967;
  assign n5969 = ~n5926 & ~n5927;
  assign n5970 = ~n5931 & n5969;
  assign n5971 = n5931 & ~n5969;
  assign n5972 = ~n5970 & ~n5971;
  assign n5973 = n5968 & ~n5972;
  assign n5974 = ~n5968 & n5972;
  assign n5975 = ~n5738 & ~n5739;
  assign n5976 = ~n5743 & n5975;
  assign n5977 = n5743 & ~n5975;
  assign n5978 = ~n5976 & ~n5977;
  assign n5979 = ~n5974 & ~n5978;
  assign n5980 = ~n5973 & ~n5979;
  assign n5981 = ~n5963 & n5980;
  assign n5982 = ~n5962 & ~n5981;
  assign n5983 = ~n5953 & ~n5982;
  assign n5984 = ~n5952 & ~n5983;
  assign n5985 = n5943 & ~n5984;
  assign n5986 = ~n5943 & n5984;
  assign n5987 = ~n5985 & ~n5986;
  assign n5988 = n5755 & n5987;
  assign n5989 = ~n5755 & ~n5987;
  assign n5990 = ~n5988 & ~n5989;
  assign n5991 = n5567 & ~n5990;
  assign n5992 = ~n5567 & n5990;
  assign n5993 = ~n5952 & ~n5953;
  assign n5994 = ~n5982 & n5993;
  assign n5995 = n5982 & ~n5993;
  assign n5996 = ~n5994 & ~n5995;
  assign n5997 = ~n5529 & ~n5530;
  assign n5998 = ~n5559 & n5997;
  assign n5999 = n5559 & ~n5997;
  assign n6000 = ~n5998 & ~n5999;
  assign n6001 = ~n5996 & ~n6000;
  assign n6002 = n5996 & n6000;
  assign n6003 = ~n5539 & ~n5540;
  assign n6004 = ~n5557 & n6003;
  assign n6005 = n5557 & ~n6003;
  assign n6006 = ~n6004 & ~n6005;
  assign n6007 = ~n5962 & ~n5963;
  assign n6008 = ~n5980 & n6007;
  assign n6009 = n5980 & ~n6007;
  assign n6010 = ~n6008 & ~n6009;
  assign n6011 = ~n6006 & ~n6010;
  assign n6012 = n6006 & n6010;
  assign n6013 = n5965 & ~n5967;
  assign n6014 = ~n5965 & n5967;
  assign n6015 = ~n6013 & ~n6014;
  assign n6016 = n5542 & ~n5544;
  assign n6017 = ~n5542 & n5544;
  assign n6018 = ~n6016 & ~n6017;
  assign n6019 = ~n6015 & ~n6018;
  assign n6020 = ~n5973 & ~n5974;
  assign n6021 = n5978 & n6020;
  assign n6022 = ~n5978 & ~n6020;
  assign n6023 = ~n6021 & ~n6022;
  assign n6024 = n6019 & ~n6023;
  assign n6025 = ~n6019 & n6023;
  assign n6026 = ~n5550 & ~n5551;
  assign n6027 = n5555 & n6026;
  assign n6028 = ~n5555 & ~n6026;
  assign n6029 = ~n6027 & ~n6028;
  assign n6030 = ~n6025 & ~n6029;
  assign n6031 = ~n6024 & ~n6030;
  assign n6032 = ~n6012 & n6031;
  assign n6033 = ~n6011 & ~n6032;
  assign n6034 = ~n6002 & n6033;
  assign n6035 = ~n6001 & ~n6034;
  assign n6036 = ~n5992 & ~n6035;
  assign n6037 = ~n5991 & ~n6036;
  assign n6038 = n5755 & ~n5986;
  assign n6039 = ~n5985 & ~n6038;
  assign n6040 = n6037 & ~n6039;
  assign n6041 = ~n6037 & n6039;
  assign n6042 = ~n5333 & ~n5563;
  assign n6043 = ~n5562 & ~n6042;
  assign n6044 = ~n6041 & ~n6043;
  assign n6045 = ~n6040 & ~n6044;
  assign n6046 = pi391  & ~pi392 ;
  assign n6047 = ~pi391  & pi392 ;
  assign n6048 = pi393  & ~n6046;
  assign n6049 = ~n6047 & n6048;
  assign n6050 = ~n6046 & ~n6047;
  assign n6051 = ~pi393  & ~n6050;
  assign n6052 = ~n6049 & ~n6051;
  assign n6053 = pi394  & ~pi395 ;
  assign n6054 = ~pi394  & pi395 ;
  assign n6055 = pi396  & ~n6053;
  assign n6056 = ~n6054 & n6055;
  assign n6057 = ~n6053 & ~n6054;
  assign n6058 = ~pi396  & ~n6057;
  assign n6059 = ~n6056 & ~n6058;
  assign n6060 = ~n6052 & n6059;
  assign n6061 = n6052 & ~n6059;
  assign n6062 = ~n6060 & ~n6061;
  assign n6063 = pi397  & ~pi398 ;
  assign n6064 = ~pi397  & pi398 ;
  assign n6065 = pi399  & ~n6063;
  assign n6066 = ~n6064 & n6065;
  assign n6067 = ~n6063 & ~n6064;
  assign n6068 = ~pi399  & ~n6067;
  assign n6069 = ~n6066 & ~n6068;
  assign n6070 = pi400  & ~pi401 ;
  assign n6071 = ~pi400  & pi401 ;
  assign n6072 = pi402  & ~n6070;
  assign n6073 = ~n6071 & n6072;
  assign n6074 = ~n6070 & ~n6071;
  assign n6075 = ~pi402  & ~n6074;
  assign n6076 = ~n6073 & ~n6075;
  assign n6077 = ~n6069 & n6076;
  assign n6078 = n6069 & ~n6076;
  assign n6079 = ~n6077 & ~n6078;
  assign n6080 = ~n6062 & ~n6079;
  assign n6081 = pi400  & pi401 ;
  assign n6082 = pi402  & ~n6074;
  assign n6083 = ~n6081 & ~n6082;
  assign n6084 = pi397  & pi398 ;
  assign n6085 = pi399  & ~n6067;
  assign n6086 = ~n6084 & ~n6085;
  assign n6087 = ~n6083 & ~n6086;
  assign n6088 = ~n6079 & n6087;
  assign n6089 = ~n6069 & ~n6076;
  assign n6090 = n6083 & n6086;
  assign n6091 = ~n6087 & ~n6090;
  assign n6092 = n6089 & n6091;
  assign n6093 = ~n6089 & ~n6091;
  assign n6094 = ~n6088 & ~n6092;
  assign n6095 = ~n6093 & n6094;
  assign n6096 = n6080 & n6095;
  assign n6097 = ~n6080 & ~n6095;
  assign n6098 = ~n6052 & ~n6059;
  assign n6099 = pi394  & pi395 ;
  assign n6100 = pi396  & ~n6057;
  assign n6101 = ~n6099 & ~n6100;
  assign n6102 = pi391  & pi392 ;
  assign n6103 = pi393  & ~n6050;
  assign n6104 = ~n6102 & ~n6103;
  assign n6105 = n6101 & ~n6104;
  assign n6106 = ~n6101 & n6104;
  assign n6107 = ~n6105 & ~n6106;
  assign n6108 = n6098 & n6107;
  assign n6109 = ~n6098 & ~n6107;
  assign n6110 = ~n6108 & ~n6109;
  assign n6111 = ~n6097 & ~n6110;
  assign n6112 = ~n6096 & ~n6111;
  assign n6113 = n6089 & ~n6090;
  assign n6114 = ~n6087 & ~n6113;
  assign n6115 = ~n6112 & ~n6114;
  assign n6116 = n6112 & n6114;
  assign n6117 = ~n6115 & ~n6116;
  assign n6118 = n6098 & ~n6101;
  assign n6119 = n6104 & ~n6118;
  assign n6120 = ~n6098 & n6101;
  assign n6121 = ~n6119 & ~n6120;
  assign n6122 = ~n6117 & n6121;
  assign n6123 = n6117 & ~n6121;
  assign n6124 = ~n6122 & ~n6123;
  assign n6125 = pi409  & ~pi410 ;
  assign n6126 = ~pi409  & pi410 ;
  assign n6127 = pi411  & ~n6125;
  assign n6128 = ~n6126 & n6127;
  assign n6129 = ~n6125 & ~n6126;
  assign n6130 = ~pi411  & ~n6129;
  assign n6131 = ~n6128 & ~n6130;
  assign n6132 = pi412  & ~pi413 ;
  assign n6133 = ~pi412  & pi413 ;
  assign n6134 = pi414  & ~n6132;
  assign n6135 = ~n6133 & n6134;
  assign n6136 = ~n6132 & ~n6133;
  assign n6137 = ~pi414  & ~n6136;
  assign n6138 = ~n6135 & ~n6137;
  assign n6139 = ~n6131 & n6138;
  assign n6140 = n6131 & ~n6138;
  assign n6141 = ~n6139 & ~n6140;
  assign n6142 = pi412  & pi413 ;
  assign n6143 = pi414  & ~n6136;
  assign n6144 = ~n6142 & ~n6143;
  assign n6145 = pi409  & pi410 ;
  assign n6146 = pi411  & ~n6129;
  assign n6147 = ~n6145 & ~n6146;
  assign n6148 = ~n6144 & ~n6147;
  assign n6149 = ~n6141 & n6148;
  assign n6150 = ~n6131 & ~n6138;
  assign n6151 = n6144 & n6147;
  assign n6152 = ~n6148 & ~n6151;
  assign n6153 = n6150 & n6152;
  assign n6154 = ~n6150 & ~n6152;
  assign n6155 = ~n6149 & ~n6153;
  assign n6156 = ~n6154 & n6155;
  assign n6157 = pi403  & ~pi404 ;
  assign n6158 = ~pi403  & pi404 ;
  assign n6159 = pi405  & ~n6157;
  assign n6160 = ~n6158 & n6159;
  assign n6161 = ~n6157 & ~n6158;
  assign n6162 = ~pi405  & ~n6161;
  assign n6163 = ~n6160 & ~n6162;
  assign n6164 = pi406  & ~pi407 ;
  assign n6165 = ~pi406  & pi407 ;
  assign n6166 = pi408  & ~n6164;
  assign n6167 = ~n6165 & n6166;
  assign n6168 = ~n6164 & ~n6165;
  assign n6169 = ~pi408  & ~n6168;
  assign n6170 = ~n6167 & ~n6169;
  assign n6171 = ~n6163 & n6170;
  assign n6172 = n6163 & ~n6170;
  assign n6173 = ~n6171 & ~n6172;
  assign n6174 = ~n6141 & ~n6173;
  assign n6175 = ~n6163 & ~n6170;
  assign n6176 = pi406  & pi407 ;
  assign n6177 = pi408  & ~n6168;
  assign n6178 = ~n6176 & ~n6177;
  assign n6179 = pi403  & pi404 ;
  assign n6180 = pi405  & ~n6161;
  assign n6181 = ~n6179 & ~n6180;
  assign n6182 = n6178 & ~n6181;
  assign n6183 = ~n6178 & n6181;
  assign n6184 = ~n6182 & ~n6183;
  assign n6185 = n6175 & n6184;
  assign n6186 = ~n6175 & ~n6184;
  assign n6187 = ~n6185 & ~n6186;
  assign n6188 = ~n6174 & n6187;
  assign n6189 = n6156 & ~n6188;
  assign n6190 = n6174 & ~n6187;
  assign n6191 = ~n6189 & ~n6190;
  assign n6192 = n6150 & ~n6151;
  assign n6193 = ~n6148 & ~n6192;
  assign n6194 = ~n6191 & ~n6193;
  assign n6195 = n6191 & n6193;
  assign n6196 = ~n6194 & ~n6195;
  assign n6197 = n6175 & ~n6178;
  assign n6198 = n6181 & ~n6197;
  assign n6199 = ~n6175 & n6178;
  assign n6200 = ~n6198 & ~n6199;
  assign n6201 = ~n6196 & n6200;
  assign n6202 = n6196 & ~n6200;
  assign n6203 = ~n6201 & ~n6202;
  assign n6204 = ~n6124 & ~n6203;
  assign n6205 = n6124 & n6203;
  assign n6206 = n6141 & n6173;
  assign n6207 = ~n6174 & ~n6206;
  assign n6208 = n6062 & n6079;
  assign n6209 = ~n6080 & ~n6208;
  assign n6210 = n6207 & n6209;
  assign n6211 = n6174 & ~n6184;
  assign n6212 = ~n6188 & ~n6211;
  assign n6213 = n6156 & ~n6212;
  assign n6214 = ~n6156 & n6212;
  assign n6215 = ~n6213 & ~n6214;
  assign n6216 = n6210 & ~n6215;
  assign n6217 = ~n6210 & n6215;
  assign n6218 = ~n6096 & ~n6097;
  assign n6219 = ~n6110 & n6218;
  assign n6220 = n6110 & ~n6218;
  assign n6221 = ~n6219 & ~n6220;
  assign n6222 = ~n6217 & n6221;
  assign n6223 = ~n6216 & ~n6222;
  assign n6224 = ~n6205 & ~n6223;
  assign n6225 = ~n6204 & ~n6224;
  assign n6226 = ~n6195 & n6200;
  assign n6227 = ~n6194 & ~n6226;
  assign n6228 = ~n6225 & ~n6227;
  assign n6229 = n6225 & n6227;
  assign n6230 = ~n6116 & n6121;
  assign n6231 = ~n6115 & ~n6230;
  assign n6232 = ~n6229 & ~n6231;
  assign n6233 = ~n6228 & ~n6232;
  assign n6234 = ~n6228 & ~n6229;
  assign n6235 = n6231 & ~n6234;
  assign n6236 = ~n6228 & n6232;
  assign n6237 = ~n6235 & ~n6236;
  assign n6238 = ~pi373  & pi374 ;
  assign n6239 = pi373  & ~pi374 ;
  assign n6240 = pi375  & ~n6238;
  assign n6241 = ~n6239 & n6240;
  assign n6242 = ~n6238 & ~n6239;
  assign n6243 = ~pi375  & ~n6242;
  assign n6244 = ~n6241 & ~n6243;
  assign n6245 = ~pi376  & pi377 ;
  assign n6246 = pi376  & ~pi377 ;
  assign n6247 = pi378  & ~n6245;
  assign n6248 = ~n6246 & n6247;
  assign n6249 = ~n6245 & ~n6246;
  assign n6250 = ~pi378  & ~n6249;
  assign n6251 = ~n6248 & ~n6250;
  assign n6252 = ~n6244 & n6251;
  assign n6253 = n6244 & ~n6251;
  assign n6254 = ~n6252 & ~n6253;
  assign n6255 = ~pi367  & pi368 ;
  assign n6256 = pi367  & ~pi368 ;
  assign n6257 = pi369  & ~n6255;
  assign n6258 = ~n6256 & n6257;
  assign n6259 = ~n6255 & ~n6256;
  assign n6260 = ~pi369  & ~n6259;
  assign n6261 = ~n6258 & ~n6260;
  assign n6262 = ~pi370  & pi371 ;
  assign n6263 = pi370  & ~pi371 ;
  assign n6264 = pi372  & ~n6262;
  assign n6265 = ~n6263 & n6264;
  assign n6266 = ~n6262 & ~n6263;
  assign n6267 = ~pi372  & ~n6266;
  assign n6268 = ~n6265 & ~n6267;
  assign n6269 = ~n6261 & n6268;
  assign n6270 = n6261 & ~n6268;
  assign n6271 = ~n6269 & ~n6270;
  assign n6272 = ~n6254 & ~n6271;
  assign n6273 = pi376  & pi377 ;
  assign n6274 = pi378  & ~n6249;
  assign n6275 = ~n6273 & ~n6274;
  assign n6276 = pi373  & pi374 ;
  assign n6277 = pi375  & ~n6242;
  assign n6278 = ~n6276 & ~n6277;
  assign n6279 = ~n6275 & ~n6278;
  assign n6280 = ~n6254 & n6279;
  assign n6281 = ~n6244 & ~n6251;
  assign n6282 = n6275 & n6278;
  assign n6283 = ~n6279 & ~n6282;
  assign n6284 = n6281 & n6283;
  assign n6285 = ~n6281 & ~n6283;
  assign n6286 = ~n6280 & ~n6284;
  assign n6287 = ~n6285 & n6286;
  assign n6288 = n6272 & n6287;
  assign n6289 = ~n6272 & ~n6287;
  assign n6290 = pi370  & pi371 ;
  assign n6291 = pi372  & ~n6266;
  assign n6292 = ~n6290 & ~n6291;
  assign n6293 = pi367  & pi368 ;
  assign n6294 = pi369  & ~n6259;
  assign n6295 = ~n6293 & ~n6294;
  assign n6296 = ~n6292 & n6295;
  assign n6297 = n6292 & ~n6295;
  assign n6298 = ~n6296 & ~n6297;
  assign n6299 = ~n6261 & ~n6268;
  assign n6300 = n6298 & n6299;
  assign n6301 = ~n6298 & ~n6299;
  assign n6302 = ~n6300 & ~n6301;
  assign n6303 = ~n6289 & ~n6302;
  assign n6304 = ~n6288 & ~n6303;
  assign n6305 = n6281 & ~n6282;
  assign n6306 = ~n6279 & ~n6305;
  assign n6307 = ~n6304 & ~n6306;
  assign n6308 = n6304 & n6306;
  assign n6309 = ~n6307 & ~n6308;
  assign n6310 = ~n6292 & n6299;
  assign n6311 = n6295 & ~n6310;
  assign n6312 = n6292 & ~n6299;
  assign n6313 = ~n6311 & ~n6312;
  assign n6314 = ~n6309 & n6313;
  assign n6315 = n6309 & ~n6313;
  assign n6316 = ~n6314 & ~n6315;
  assign n6317 = ~pi385  & pi386 ;
  assign n6318 = pi385  & ~pi386 ;
  assign n6319 = pi387  & ~n6317;
  assign n6320 = ~n6318 & n6319;
  assign n6321 = ~n6317 & ~n6318;
  assign n6322 = ~pi387  & ~n6321;
  assign n6323 = ~n6320 & ~n6322;
  assign n6324 = ~pi388  & pi389 ;
  assign n6325 = pi388  & ~pi389 ;
  assign n6326 = pi390  & ~n6324;
  assign n6327 = ~n6325 & n6326;
  assign n6328 = ~n6324 & ~n6325;
  assign n6329 = ~pi390  & ~n6328;
  assign n6330 = ~n6327 & ~n6329;
  assign n6331 = ~n6323 & n6330;
  assign n6332 = n6323 & ~n6330;
  assign n6333 = ~n6331 & ~n6332;
  assign n6334 = ~pi379  & pi380 ;
  assign n6335 = pi379  & ~pi380 ;
  assign n6336 = pi381  & ~n6334;
  assign n6337 = ~n6335 & n6336;
  assign n6338 = ~n6334 & ~n6335;
  assign n6339 = ~pi381  & ~n6338;
  assign n6340 = ~n6337 & ~n6339;
  assign n6341 = ~pi382  & pi383 ;
  assign n6342 = pi382  & ~pi383 ;
  assign n6343 = pi384  & ~n6341;
  assign n6344 = ~n6342 & n6343;
  assign n6345 = ~n6341 & ~n6342;
  assign n6346 = ~pi384  & ~n6345;
  assign n6347 = ~n6344 & ~n6346;
  assign n6348 = ~n6340 & n6347;
  assign n6349 = n6340 & ~n6347;
  assign n6350 = ~n6348 & ~n6349;
  assign n6351 = ~n6333 & ~n6350;
  assign n6352 = pi388  & pi389 ;
  assign n6353 = pi390  & ~n6328;
  assign n6354 = ~n6352 & ~n6353;
  assign n6355 = pi385  & pi386 ;
  assign n6356 = pi387  & ~n6321;
  assign n6357 = ~n6355 & ~n6356;
  assign n6358 = n6354 & ~n6357;
  assign n6359 = ~n6354 & n6357;
  assign n6360 = ~n6358 & ~n6359;
  assign n6361 = n6351 & ~n6360;
  assign n6362 = ~n6323 & ~n6330;
  assign n6363 = n6360 & n6362;
  assign n6364 = ~n6360 & ~n6362;
  assign n6365 = ~n6351 & ~n6363;
  assign n6366 = ~n6364 & n6365;
  assign n6367 = pi382  & pi383 ;
  assign n6368 = pi384  & ~n6345;
  assign n6369 = ~n6367 & ~n6368;
  assign n6370 = pi379  & pi380 ;
  assign n6371 = pi381  & ~n6338;
  assign n6372 = ~n6370 & ~n6371;
  assign n6373 = ~n6369 & ~n6372;
  assign n6374 = ~n6350 & n6373;
  assign n6375 = ~n6340 & ~n6347;
  assign n6376 = n6369 & n6372;
  assign n6377 = ~n6373 & ~n6376;
  assign n6378 = n6375 & n6377;
  assign n6379 = ~n6375 & ~n6377;
  assign n6380 = ~n6374 & ~n6378;
  assign n6381 = ~n6379 & n6380;
  assign n6382 = ~n6366 & n6381;
  assign n6383 = ~n6361 & ~n6382;
  assign n6384 = ~n6354 & n6362;
  assign n6385 = n6357 & ~n6384;
  assign n6386 = n6354 & ~n6362;
  assign n6387 = ~n6385 & ~n6386;
  assign n6388 = ~n6383 & n6387;
  assign n6389 = n6383 & ~n6387;
  assign n6390 = ~n6388 & ~n6389;
  assign n6391 = n6375 & ~n6376;
  assign n6392 = ~n6373 & ~n6391;
  assign n6393 = n6390 & ~n6392;
  assign n6394 = ~n6390 & n6392;
  assign n6395 = ~n6393 & ~n6394;
  assign n6396 = n6316 & ~n6395;
  assign n6397 = ~n6316 & n6395;
  assign n6398 = n6333 & n6350;
  assign n6399 = ~n6351 & ~n6398;
  assign n6400 = n6254 & n6271;
  assign n6401 = ~n6272 & ~n6400;
  assign n6402 = n6399 & n6401;
  assign n6403 = ~n6361 & ~n6366;
  assign n6404 = n6381 & n6403;
  assign n6405 = ~n6381 & ~n6403;
  assign n6406 = ~n6404 & ~n6405;
  assign n6407 = n6402 & n6406;
  assign n6408 = ~n6402 & ~n6406;
  assign n6409 = ~n6288 & ~n6289;
  assign n6410 = ~n6302 & n6409;
  assign n6411 = n6302 & ~n6409;
  assign n6412 = ~n6410 & ~n6411;
  assign n6413 = ~n6408 & n6412;
  assign n6414 = ~n6407 & ~n6413;
  assign n6415 = ~n6397 & n6414;
  assign n6416 = ~n6396 & ~n6415;
  assign n6417 = ~n6389 & ~n6392;
  assign n6418 = ~n6388 & ~n6417;
  assign n6419 = ~n6416 & n6418;
  assign n6420 = n6416 & ~n6418;
  assign n6421 = ~n6419 & ~n6420;
  assign n6422 = ~n6308 & n6313;
  assign n6423 = ~n6307 & ~n6422;
  assign n6424 = n6421 & n6423;
  assign n6425 = ~n6421 & ~n6423;
  assign n6426 = ~n6424 & ~n6425;
  assign n6427 = n6237 & ~n6426;
  assign n6428 = ~n6237 & n6426;
  assign n6429 = ~n6396 & ~n6397;
  assign n6430 = ~n6414 & n6429;
  assign n6431 = n6414 & ~n6429;
  assign n6432 = ~n6430 & ~n6431;
  assign n6433 = ~n6204 & ~n6205;
  assign n6434 = ~n6223 & n6433;
  assign n6435 = n6223 & ~n6433;
  assign n6436 = ~n6434 & ~n6435;
  assign n6437 = ~n6432 & ~n6436;
  assign n6438 = n6432 & n6436;
  assign n6439 = ~n6207 & ~n6209;
  assign n6440 = ~n6210 & ~n6439;
  assign n6441 = ~n6399 & ~n6401;
  assign n6442 = ~n6402 & ~n6441;
  assign n6443 = n6440 & n6442;
  assign n6444 = ~n6216 & ~n6217;
  assign n6445 = ~n6221 & n6444;
  assign n6446 = n6221 & ~n6444;
  assign n6447 = ~n6445 & ~n6446;
  assign n6448 = n6443 & ~n6447;
  assign n6449 = ~n6443 & n6447;
  assign n6450 = ~n6407 & ~n6408;
  assign n6451 = ~n6412 & n6450;
  assign n6452 = n6412 & ~n6450;
  assign n6453 = ~n6451 & ~n6452;
  assign n6454 = ~n6449 & ~n6453;
  assign n6455 = ~n6448 & ~n6454;
  assign n6456 = ~n6438 & n6455;
  assign n6457 = ~n6437 & ~n6456;
  assign n6458 = ~n6428 & n6457;
  assign n6459 = ~n6427 & ~n6458;
  assign n6460 = n6233 & n6459;
  assign n6461 = ~n6233 & ~n6459;
  assign n6462 = ~n6420 & n6423;
  assign n6463 = ~n6419 & ~n6462;
  assign n6464 = ~n6461 & ~n6463;
  assign n6465 = ~n6460 & ~n6464;
  assign n6466 = n6233 & ~n6459;
  assign n6467 = ~n6233 & n6459;
  assign n6468 = ~n6466 & ~n6467;
  assign n6469 = n6463 & n6468;
  assign n6470 = ~n6463 & ~n6468;
  assign n6471 = ~n6469 & ~n6470;
  assign n6472 = ~pi421  & pi422 ;
  assign n6473 = pi421  & ~pi422 ;
  assign n6474 = pi423  & ~n6472;
  assign n6475 = ~n6473 & n6474;
  assign n6476 = ~n6472 & ~n6473;
  assign n6477 = ~pi423  & ~n6476;
  assign n6478 = ~n6475 & ~n6477;
  assign n6479 = ~pi424  & pi425 ;
  assign n6480 = pi424  & ~pi425 ;
  assign n6481 = pi426  & ~n6479;
  assign n6482 = ~n6480 & n6481;
  assign n6483 = ~n6479 & ~n6480;
  assign n6484 = ~pi426  & ~n6483;
  assign n6485 = ~n6482 & ~n6484;
  assign n6486 = ~n6478 & n6485;
  assign n6487 = n6478 & ~n6485;
  assign n6488 = ~n6486 & ~n6487;
  assign n6489 = ~pi415  & pi416 ;
  assign n6490 = pi415  & ~pi416 ;
  assign n6491 = pi417  & ~n6489;
  assign n6492 = ~n6490 & n6491;
  assign n6493 = ~n6489 & ~n6490;
  assign n6494 = ~pi417  & ~n6493;
  assign n6495 = ~n6492 & ~n6494;
  assign n6496 = ~pi418  & pi419 ;
  assign n6497 = pi418  & ~pi419 ;
  assign n6498 = pi420  & ~n6496;
  assign n6499 = ~n6497 & n6498;
  assign n6500 = ~n6496 & ~n6497;
  assign n6501 = ~pi420  & ~n6500;
  assign n6502 = ~n6499 & ~n6501;
  assign n6503 = ~n6495 & n6502;
  assign n6504 = n6495 & ~n6502;
  assign n6505 = ~n6503 & ~n6504;
  assign n6506 = ~n6488 & ~n6505;
  assign n6507 = pi424  & pi425 ;
  assign n6508 = pi426  & ~n6483;
  assign n6509 = ~n6507 & ~n6508;
  assign n6510 = pi421  & pi422 ;
  assign n6511 = pi423  & ~n6476;
  assign n6512 = ~n6510 & ~n6511;
  assign n6513 = ~n6509 & ~n6512;
  assign n6514 = ~n6488 & n6513;
  assign n6515 = ~n6478 & ~n6485;
  assign n6516 = n6509 & n6512;
  assign n6517 = ~n6513 & ~n6516;
  assign n6518 = n6515 & n6517;
  assign n6519 = ~n6515 & ~n6517;
  assign n6520 = ~n6514 & ~n6518;
  assign n6521 = ~n6519 & n6520;
  assign n6522 = n6506 & n6521;
  assign n6523 = ~n6506 & ~n6521;
  assign n6524 = pi418  & pi419 ;
  assign n6525 = pi420  & ~n6500;
  assign n6526 = ~n6524 & ~n6525;
  assign n6527 = pi415  & pi416 ;
  assign n6528 = pi417  & ~n6493;
  assign n6529 = ~n6527 & ~n6528;
  assign n6530 = ~n6526 & n6529;
  assign n6531 = n6526 & ~n6529;
  assign n6532 = ~n6530 & ~n6531;
  assign n6533 = ~n6495 & ~n6502;
  assign n6534 = n6532 & n6533;
  assign n6535 = ~n6532 & ~n6533;
  assign n6536 = ~n6534 & ~n6535;
  assign n6537 = ~n6523 & ~n6536;
  assign n6538 = ~n6522 & ~n6537;
  assign n6539 = n6515 & ~n6516;
  assign n6540 = ~n6513 & ~n6539;
  assign n6541 = ~n6538 & ~n6540;
  assign n6542 = n6538 & n6540;
  assign n6543 = ~n6541 & ~n6542;
  assign n6544 = ~n6526 & n6533;
  assign n6545 = n6529 & ~n6544;
  assign n6546 = n6526 & ~n6533;
  assign n6547 = ~n6545 & ~n6546;
  assign n6548 = ~n6543 & n6547;
  assign n6549 = n6543 & ~n6547;
  assign n6550 = ~n6548 & ~n6549;
  assign n6551 = pi433  & ~pi434 ;
  assign n6552 = ~pi433  & pi434 ;
  assign n6553 = pi435  & ~n6551;
  assign n6554 = ~n6552 & n6553;
  assign n6555 = ~n6551 & ~n6552;
  assign n6556 = ~pi435  & ~n6555;
  assign n6557 = ~n6554 & ~n6556;
  assign n6558 = pi436  & ~pi437 ;
  assign n6559 = ~pi436  & pi437 ;
  assign n6560 = pi438  & ~n6558;
  assign n6561 = ~n6559 & n6560;
  assign n6562 = ~n6558 & ~n6559;
  assign n6563 = ~pi438  & ~n6562;
  assign n6564 = ~n6561 & ~n6563;
  assign n6565 = ~n6557 & n6564;
  assign n6566 = n6557 & ~n6564;
  assign n6567 = ~n6565 & ~n6566;
  assign n6568 = pi436  & pi437 ;
  assign n6569 = pi438  & ~n6562;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = pi433  & pi434 ;
  assign n6572 = pi435  & ~n6555;
  assign n6573 = ~n6571 & ~n6572;
  assign n6574 = ~n6570 & ~n6573;
  assign n6575 = ~n6567 & n6574;
  assign n6576 = ~n6557 & ~n6564;
  assign n6577 = n6570 & n6573;
  assign n6578 = ~n6574 & ~n6577;
  assign n6579 = n6576 & n6578;
  assign n6580 = ~n6576 & ~n6578;
  assign n6581 = ~n6575 & ~n6579;
  assign n6582 = ~n6580 & n6581;
  assign n6583 = pi427  & ~pi428 ;
  assign n6584 = ~pi427  & pi428 ;
  assign n6585 = pi429  & ~n6583;
  assign n6586 = ~n6584 & n6585;
  assign n6587 = ~n6583 & ~n6584;
  assign n6588 = ~pi429  & ~n6587;
  assign n6589 = ~n6586 & ~n6588;
  assign n6590 = pi430  & ~pi431 ;
  assign n6591 = ~pi430  & pi431 ;
  assign n6592 = pi432  & ~n6590;
  assign n6593 = ~n6591 & n6592;
  assign n6594 = ~n6590 & ~n6591;
  assign n6595 = ~pi432  & ~n6594;
  assign n6596 = ~n6593 & ~n6595;
  assign n6597 = ~n6589 & n6596;
  assign n6598 = n6589 & ~n6596;
  assign n6599 = ~n6597 & ~n6598;
  assign n6600 = ~n6567 & ~n6599;
  assign n6601 = ~n6589 & ~n6596;
  assign n6602 = pi430  & pi431 ;
  assign n6603 = pi432  & ~n6594;
  assign n6604 = ~n6602 & ~n6603;
  assign n6605 = pi427  & pi428 ;
  assign n6606 = pi429  & ~n6587;
  assign n6607 = ~n6605 & ~n6606;
  assign n6608 = n6604 & ~n6607;
  assign n6609 = ~n6604 & n6607;
  assign n6610 = ~n6608 & ~n6609;
  assign n6611 = n6601 & n6610;
  assign n6612 = ~n6601 & ~n6610;
  assign n6613 = ~n6611 & ~n6612;
  assign n6614 = ~n6600 & n6613;
  assign n6615 = n6582 & ~n6614;
  assign n6616 = n6600 & ~n6613;
  assign n6617 = ~n6615 & ~n6616;
  assign n6618 = n6576 & ~n6577;
  assign n6619 = ~n6574 & ~n6618;
  assign n6620 = ~n6617 & ~n6619;
  assign n6621 = n6617 & n6619;
  assign n6622 = ~n6620 & ~n6621;
  assign n6623 = n6601 & ~n6604;
  assign n6624 = n6607 & ~n6623;
  assign n6625 = ~n6601 & n6604;
  assign n6626 = ~n6624 & ~n6625;
  assign n6627 = ~n6622 & n6626;
  assign n6628 = n6622 & ~n6626;
  assign n6629 = ~n6627 & ~n6628;
  assign n6630 = ~n6550 & ~n6629;
  assign n6631 = n6550 & n6629;
  assign n6632 = n6567 & n6599;
  assign n6633 = ~n6600 & ~n6632;
  assign n6634 = n6488 & n6505;
  assign n6635 = ~n6506 & ~n6634;
  assign n6636 = n6633 & n6635;
  assign n6637 = n6600 & ~n6610;
  assign n6638 = ~n6614 & ~n6637;
  assign n6639 = n6582 & ~n6638;
  assign n6640 = ~n6582 & n6638;
  assign n6641 = ~n6639 & ~n6640;
  assign n6642 = n6636 & ~n6641;
  assign n6643 = ~n6636 & n6641;
  assign n6644 = ~n6522 & ~n6523;
  assign n6645 = ~n6536 & n6644;
  assign n6646 = n6536 & ~n6644;
  assign n6647 = ~n6645 & ~n6646;
  assign n6648 = ~n6643 & n6647;
  assign n6649 = ~n6642 & ~n6648;
  assign n6650 = ~n6631 & ~n6649;
  assign n6651 = ~n6630 & ~n6650;
  assign n6652 = ~n6621 & n6626;
  assign n6653 = ~n6620 & ~n6652;
  assign n6654 = ~n6651 & ~n6653;
  assign n6655 = n6651 & n6653;
  assign n6656 = ~n6542 & n6547;
  assign n6657 = ~n6541 & ~n6656;
  assign n6658 = ~n6655 & ~n6657;
  assign n6659 = ~n6654 & ~n6658;
  assign n6660 = pi439  & ~pi440 ;
  assign n6661 = ~pi439  & pi440 ;
  assign n6662 = pi441  & ~n6660;
  assign n6663 = ~n6661 & n6662;
  assign n6664 = ~n6660 & ~n6661;
  assign n6665 = ~pi441  & ~n6664;
  assign n6666 = ~n6663 & ~n6665;
  assign n6667 = pi442  & ~pi443 ;
  assign n6668 = ~pi442  & pi443 ;
  assign n6669 = pi444  & ~n6667;
  assign n6670 = ~n6668 & n6669;
  assign n6671 = ~n6667 & ~n6668;
  assign n6672 = ~pi444  & ~n6671;
  assign n6673 = ~n6670 & ~n6672;
  assign n6674 = ~n6666 & n6673;
  assign n6675 = n6666 & ~n6673;
  assign n6676 = ~n6674 & ~n6675;
  assign n6677 = pi445  & ~pi446 ;
  assign n6678 = ~pi445  & pi446 ;
  assign n6679 = pi447  & ~n6677;
  assign n6680 = ~n6678 & n6679;
  assign n6681 = ~n6677 & ~n6678;
  assign n6682 = ~pi447  & ~n6681;
  assign n6683 = ~n6680 & ~n6682;
  assign n6684 = pi448  & ~pi449 ;
  assign n6685 = ~pi448  & pi449 ;
  assign n6686 = pi450  & ~n6684;
  assign n6687 = ~n6685 & n6686;
  assign n6688 = ~n6684 & ~n6685;
  assign n6689 = ~pi450  & ~n6688;
  assign n6690 = ~n6687 & ~n6689;
  assign n6691 = ~n6683 & n6690;
  assign n6692 = n6683 & ~n6690;
  assign n6693 = ~n6691 & ~n6692;
  assign n6694 = ~n6676 & ~n6693;
  assign n6695 = pi448  & pi449 ;
  assign n6696 = pi450  & ~n6688;
  assign n6697 = ~n6695 & ~n6696;
  assign n6698 = pi445  & pi446 ;
  assign n6699 = pi447  & ~n6681;
  assign n6700 = ~n6698 & ~n6699;
  assign n6701 = ~n6697 & ~n6700;
  assign n6702 = ~n6693 & n6701;
  assign n6703 = ~n6683 & ~n6690;
  assign n6704 = n6697 & n6700;
  assign n6705 = ~n6701 & ~n6704;
  assign n6706 = n6703 & n6705;
  assign n6707 = ~n6703 & ~n6705;
  assign n6708 = ~n6702 & ~n6706;
  assign n6709 = ~n6707 & n6708;
  assign n6710 = n6694 & n6709;
  assign n6711 = ~n6694 & ~n6709;
  assign n6712 = ~n6666 & ~n6673;
  assign n6713 = pi442  & pi443 ;
  assign n6714 = pi444  & ~n6671;
  assign n6715 = ~n6713 & ~n6714;
  assign n6716 = pi439  & pi440 ;
  assign n6717 = pi441  & ~n6664;
  assign n6718 = ~n6716 & ~n6717;
  assign n6719 = n6715 & ~n6718;
  assign n6720 = ~n6715 & n6718;
  assign n6721 = ~n6719 & ~n6720;
  assign n6722 = n6712 & n6721;
  assign n6723 = ~n6712 & ~n6721;
  assign n6724 = ~n6722 & ~n6723;
  assign n6725 = ~n6711 & ~n6724;
  assign n6726 = ~n6710 & ~n6725;
  assign n6727 = n6703 & ~n6704;
  assign n6728 = ~n6701 & ~n6727;
  assign n6729 = ~n6726 & ~n6728;
  assign n6730 = n6726 & n6728;
  assign n6731 = ~n6729 & ~n6730;
  assign n6732 = n6712 & ~n6715;
  assign n6733 = n6718 & ~n6732;
  assign n6734 = ~n6712 & n6715;
  assign n6735 = ~n6733 & ~n6734;
  assign n6736 = ~n6731 & n6735;
  assign n6737 = n6731 & ~n6735;
  assign n6738 = ~n6736 & ~n6737;
  assign n6739 = pi457  & ~pi458 ;
  assign n6740 = ~pi457  & pi458 ;
  assign n6741 = pi459  & ~n6739;
  assign n6742 = ~n6740 & n6741;
  assign n6743 = ~n6739 & ~n6740;
  assign n6744 = ~pi459  & ~n6743;
  assign n6745 = ~n6742 & ~n6744;
  assign n6746 = pi460  & ~pi461 ;
  assign n6747 = ~pi460  & pi461 ;
  assign n6748 = pi462  & ~n6746;
  assign n6749 = ~n6747 & n6748;
  assign n6750 = ~n6746 & ~n6747;
  assign n6751 = ~pi462  & ~n6750;
  assign n6752 = ~n6749 & ~n6751;
  assign n6753 = ~n6745 & n6752;
  assign n6754 = n6745 & ~n6752;
  assign n6755 = ~n6753 & ~n6754;
  assign n6756 = pi460  & pi461 ;
  assign n6757 = pi462  & ~n6750;
  assign n6758 = ~n6756 & ~n6757;
  assign n6759 = pi457  & pi458 ;
  assign n6760 = pi459  & ~n6743;
  assign n6761 = ~n6759 & ~n6760;
  assign n6762 = ~n6758 & ~n6761;
  assign n6763 = ~n6755 & n6762;
  assign n6764 = ~n6745 & ~n6752;
  assign n6765 = n6758 & n6761;
  assign n6766 = ~n6762 & ~n6765;
  assign n6767 = n6764 & n6766;
  assign n6768 = ~n6764 & ~n6766;
  assign n6769 = ~n6763 & ~n6767;
  assign n6770 = ~n6768 & n6769;
  assign n6771 = pi451  & ~pi452 ;
  assign n6772 = ~pi451  & pi452 ;
  assign n6773 = pi453  & ~n6771;
  assign n6774 = ~n6772 & n6773;
  assign n6775 = ~n6771 & ~n6772;
  assign n6776 = ~pi453  & ~n6775;
  assign n6777 = ~n6774 & ~n6776;
  assign n6778 = pi454  & ~pi455 ;
  assign n6779 = ~pi454  & pi455 ;
  assign n6780 = pi456  & ~n6778;
  assign n6781 = ~n6779 & n6780;
  assign n6782 = ~n6778 & ~n6779;
  assign n6783 = ~pi456  & ~n6782;
  assign n6784 = ~n6781 & ~n6783;
  assign n6785 = ~n6777 & n6784;
  assign n6786 = n6777 & ~n6784;
  assign n6787 = ~n6785 & ~n6786;
  assign n6788 = ~n6755 & ~n6787;
  assign n6789 = ~n6777 & ~n6784;
  assign n6790 = pi454  & pi455 ;
  assign n6791 = pi456  & ~n6782;
  assign n6792 = ~n6790 & ~n6791;
  assign n6793 = pi451  & pi452 ;
  assign n6794 = pi453  & ~n6775;
  assign n6795 = ~n6793 & ~n6794;
  assign n6796 = n6792 & ~n6795;
  assign n6797 = ~n6792 & n6795;
  assign n6798 = ~n6796 & ~n6797;
  assign n6799 = n6789 & n6798;
  assign n6800 = ~n6789 & ~n6798;
  assign n6801 = ~n6799 & ~n6800;
  assign n6802 = ~n6788 & n6801;
  assign n6803 = n6770 & ~n6802;
  assign n6804 = n6788 & ~n6801;
  assign n6805 = ~n6803 & ~n6804;
  assign n6806 = n6764 & ~n6765;
  assign n6807 = ~n6762 & ~n6806;
  assign n6808 = ~n6805 & ~n6807;
  assign n6809 = n6805 & n6807;
  assign n6810 = ~n6808 & ~n6809;
  assign n6811 = n6789 & ~n6792;
  assign n6812 = n6795 & ~n6811;
  assign n6813 = ~n6789 & n6792;
  assign n6814 = ~n6812 & ~n6813;
  assign n6815 = ~n6810 & n6814;
  assign n6816 = n6810 & ~n6814;
  assign n6817 = ~n6815 & ~n6816;
  assign n6818 = ~n6738 & ~n6817;
  assign n6819 = n6738 & n6817;
  assign n6820 = n6755 & n6787;
  assign n6821 = ~n6788 & ~n6820;
  assign n6822 = n6676 & n6693;
  assign n6823 = ~n6694 & ~n6822;
  assign n6824 = n6821 & n6823;
  assign n6825 = n6788 & ~n6798;
  assign n6826 = ~n6802 & ~n6825;
  assign n6827 = n6770 & ~n6826;
  assign n6828 = ~n6770 & n6826;
  assign n6829 = ~n6827 & ~n6828;
  assign n6830 = n6824 & ~n6829;
  assign n6831 = ~n6824 & n6829;
  assign n6832 = ~n6710 & ~n6711;
  assign n6833 = ~n6724 & n6832;
  assign n6834 = n6724 & ~n6832;
  assign n6835 = ~n6833 & ~n6834;
  assign n6836 = ~n6831 & n6835;
  assign n6837 = ~n6830 & ~n6836;
  assign n6838 = ~n6819 & ~n6837;
  assign n6839 = ~n6818 & ~n6838;
  assign n6840 = ~n6809 & n6814;
  assign n6841 = ~n6808 & ~n6840;
  assign n6842 = ~n6839 & ~n6841;
  assign n6843 = n6839 & n6841;
  assign n6844 = ~n6730 & n6735;
  assign n6845 = ~n6729 & ~n6844;
  assign n6846 = ~n6843 & ~n6845;
  assign n6847 = ~n6842 & ~n6846;
  assign n6848 = ~n6842 & ~n6843;
  assign n6849 = n6845 & ~n6848;
  assign n6850 = ~n6842 & n6846;
  assign n6851 = ~n6849 & ~n6850;
  assign n6852 = ~n6654 & ~n6655;
  assign n6853 = n6657 & ~n6852;
  assign n6854 = ~n6654 & n6658;
  assign n6855 = ~n6853 & ~n6854;
  assign n6856 = ~n6851 & ~n6855;
  assign n6857 = n6851 & n6855;
  assign n6858 = ~n6630 & ~n6631;
  assign n6859 = ~n6649 & n6858;
  assign n6860 = n6649 & ~n6858;
  assign n6861 = ~n6859 & ~n6860;
  assign n6862 = ~n6818 & ~n6819;
  assign n6863 = ~n6837 & n6862;
  assign n6864 = n6837 & ~n6862;
  assign n6865 = ~n6863 & ~n6864;
  assign n6866 = ~n6861 & ~n6865;
  assign n6867 = n6861 & n6865;
  assign n6868 = ~n6821 & ~n6823;
  assign n6869 = ~n6824 & ~n6868;
  assign n6870 = ~n6633 & ~n6635;
  assign n6871 = ~n6636 & ~n6870;
  assign n6872 = n6869 & n6871;
  assign n6873 = ~n6830 & ~n6831;
  assign n6874 = ~n6835 & n6873;
  assign n6875 = n6835 & ~n6873;
  assign n6876 = ~n6874 & ~n6875;
  assign n6877 = n6872 & ~n6876;
  assign n6878 = ~n6872 & n6876;
  assign n6879 = ~n6642 & ~n6643;
  assign n6880 = ~n6647 & n6879;
  assign n6881 = n6647 & ~n6879;
  assign n6882 = ~n6880 & ~n6881;
  assign n6883 = ~n6878 & ~n6882;
  assign n6884 = ~n6877 & ~n6883;
  assign n6885 = ~n6867 & n6884;
  assign n6886 = ~n6866 & ~n6885;
  assign n6887 = ~n6857 & ~n6886;
  assign n6888 = ~n6856 & ~n6887;
  assign n6889 = n6847 & ~n6888;
  assign n6890 = ~n6847 & n6888;
  assign n6891 = ~n6889 & ~n6890;
  assign n6892 = n6659 & n6891;
  assign n6893 = ~n6659 & ~n6891;
  assign n6894 = ~n6892 & ~n6893;
  assign n6895 = ~n6471 & ~n6894;
  assign n6896 = n6471 & n6894;
  assign n6897 = ~n6856 & ~n6857;
  assign n6898 = ~n6886 & n6897;
  assign n6899 = n6886 & ~n6897;
  assign n6900 = ~n6898 & ~n6899;
  assign n6901 = ~n6427 & ~n6428;
  assign n6902 = ~n6457 & n6901;
  assign n6903 = n6457 & ~n6901;
  assign n6904 = ~n6902 & ~n6903;
  assign n6905 = ~n6900 & ~n6904;
  assign n6906 = n6900 & n6904;
  assign n6907 = ~n6437 & ~n6438;
  assign n6908 = ~n6455 & n6907;
  assign n6909 = n6455 & ~n6907;
  assign n6910 = ~n6908 & ~n6909;
  assign n6911 = ~n6866 & ~n6867;
  assign n6912 = ~n6884 & n6911;
  assign n6913 = n6884 & ~n6911;
  assign n6914 = ~n6912 & ~n6913;
  assign n6915 = ~n6910 & ~n6914;
  assign n6916 = n6910 & n6914;
  assign n6917 = n6869 & ~n6871;
  assign n6918 = ~n6869 & n6871;
  assign n6919 = ~n6917 & ~n6918;
  assign n6920 = n6440 & ~n6442;
  assign n6921 = ~n6440 & n6442;
  assign n6922 = ~n6920 & ~n6921;
  assign n6923 = ~n6919 & ~n6922;
  assign n6924 = ~n6877 & ~n6878;
  assign n6925 = n6882 & n6924;
  assign n6926 = ~n6882 & ~n6924;
  assign n6927 = ~n6925 & ~n6926;
  assign n6928 = n6923 & ~n6927;
  assign n6929 = ~n6923 & n6927;
  assign n6930 = ~n6448 & ~n6449;
  assign n6931 = n6453 & n6930;
  assign n6932 = ~n6453 & ~n6930;
  assign n6933 = ~n6931 & ~n6932;
  assign n6934 = ~n6929 & ~n6933;
  assign n6935 = ~n6928 & ~n6934;
  assign n6936 = ~n6916 & n6935;
  assign n6937 = ~n6915 & ~n6936;
  assign n6938 = ~n6906 & n6937;
  assign n6939 = ~n6905 & ~n6938;
  assign n6940 = ~n6896 & ~n6939;
  assign n6941 = ~n6895 & ~n6940;
  assign n6942 = n6659 & ~n6890;
  assign n6943 = ~n6889 & ~n6942;
  assign n6944 = n6941 & ~n6943;
  assign n6945 = ~n6941 & n6943;
  assign n6946 = ~n6944 & ~n6945;
  assign n6947 = ~n6465 & ~n6946;
  assign n6948 = n6465 & n6946;
  assign n6949 = ~n6947 & ~n6948;
  assign n6950 = ~n6040 & ~n6041;
  assign n6951 = ~n6043 & ~n6950;
  assign n6952 = n6043 & n6950;
  assign n6953 = ~n6951 & ~n6952;
  assign n6954 = ~n6949 & ~n6953;
  assign n6955 = n6949 & n6953;
  assign n6956 = ~n5991 & ~n5992;
  assign n6957 = ~n6035 & n6956;
  assign n6958 = n6035 & ~n6956;
  assign n6959 = ~n6957 & ~n6958;
  assign n6960 = ~n6895 & ~n6896;
  assign n6961 = ~n6939 & n6960;
  assign n6962 = n6939 & ~n6960;
  assign n6963 = ~n6961 & ~n6962;
  assign n6964 = ~n6959 & ~n6963;
  assign n6965 = n6959 & n6963;
  assign n6966 = ~n6905 & ~n6906;
  assign n6967 = n6937 & n6966;
  assign n6968 = ~n6937 & ~n6966;
  assign n6969 = ~n6967 & ~n6968;
  assign n6970 = ~n6001 & ~n6002;
  assign n6971 = n6033 & n6970;
  assign n6972 = ~n6033 & ~n6970;
  assign n6973 = ~n6971 & ~n6972;
  assign n6974 = ~n6969 & ~n6973;
  assign n6975 = n6969 & n6973;
  assign n6976 = ~n6011 & ~n6012;
  assign n6977 = ~n6031 & n6976;
  assign n6978 = n6031 & ~n6976;
  assign n6979 = ~n6977 & ~n6978;
  assign n6980 = ~n6915 & ~n6916;
  assign n6981 = ~n6935 & n6980;
  assign n6982 = n6935 & ~n6980;
  assign n6983 = ~n6981 & ~n6982;
  assign n6984 = ~n6979 & ~n6983;
  assign n6985 = n6979 & n6983;
  assign n6986 = n6919 & n6922;
  assign n6987 = ~n6923 & ~n6986;
  assign n6988 = n6015 & n6018;
  assign n6989 = ~n6019 & ~n6988;
  assign n6990 = n6987 & n6989;
  assign n6991 = ~n6928 & ~n6929;
  assign n6992 = n6933 & n6991;
  assign n6993 = ~n6933 & ~n6991;
  assign n6994 = ~n6992 & ~n6993;
  assign n6995 = n6990 & ~n6994;
  assign n6996 = ~n6990 & n6994;
  assign n6997 = ~n6024 & ~n6025;
  assign n6998 = n6029 & n6997;
  assign n6999 = ~n6029 & ~n6997;
  assign n7000 = ~n6998 & ~n6999;
  assign n7001 = ~n6996 & ~n7000;
  assign n7002 = ~n6995 & ~n7001;
  assign n7003 = ~n6985 & n7002;
  assign n7004 = ~n6984 & ~n7003;
  assign n7005 = ~n6975 & ~n7004;
  assign n7006 = ~n6974 & ~n7005;
  assign n7007 = ~n6965 & ~n7006;
  assign n7008 = ~n6964 & ~n7007;
  assign n7009 = ~n6955 & ~n7008;
  assign n7010 = ~n6954 & ~n7009;
  assign n7011 = ~n6465 & ~n6945;
  assign n7012 = ~n6944 & ~n7011;
  assign n7013 = n7010 & ~n7012;
  assign n7014 = ~n7010 & n7012;
  assign n7015 = ~n7013 & ~n7014;
  assign n7016 = n6045 & n7015;
  assign n7017 = ~n6045 & ~n7015;
  assign n7018 = ~n7016 & ~n7017;
  assign n7019 = n5146 & ~n7018;
  assign n7020 = ~n5146 & n7018;
  assign n7021 = ~n6954 & ~n6955;
  assign n7022 = ~n7008 & n7021;
  assign n7023 = n7008 & ~n7021;
  assign n7024 = ~n7022 & ~n7023;
  assign n7025 = ~n5084 & ~n5085;
  assign n7026 = ~n5138 & n7025;
  assign n7027 = n5138 & ~n7025;
  assign n7028 = ~n7026 & ~n7027;
  assign n7029 = ~n7024 & ~n7028;
  assign n7030 = n7024 & n7028;
  assign n7031 = ~n5094 & ~n5095;
  assign n7032 = n5136 & n7031;
  assign n7033 = ~n5136 & ~n7031;
  assign n7034 = ~n7032 & ~n7033;
  assign n7035 = ~n6964 & ~n6965;
  assign n7036 = n7006 & n7035;
  assign n7037 = ~n7006 & ~n7035;
  assign n7038 = ~n7036 & ~n7037;
  assign n7039 = ~n7034 & ~n7038;
  assign n7040 = n7034 & n7038;
  assign n7041 = ~n6974 & ~n6975;
  assign n7042 = ~n7004 & n7041;
  assign n7043 = n7004 & ~n7041;
  assign n7044 = ~n7042 & ~n7043;
  assign n7045 = ~n5104 & ~n5105;
  assign n7046 = ~n5134 & n7045;
  assign n7047 = n5134 & ~n7045;
  assign n7048 = ~n7046 & ~n7047;
  assign n7049 = ~n7044 & ~n7048;
  assign n7050 = n7044 & n7048;
  assign n7051 = ~n5114 & ~n5115;
  assign n7052 = ~n5132 & n7051;
  assign n7053 = n5132 & ~n7051;
  assign n7054 = ~n7052 & ~n7053;
  assign n7055 = ~n6984 & ~n6985;
  assign n7056 = ~n7002 & n7055;
  assign n7057 = n7002 & ~n7055;
  assign n7058 = ~n7056 & ~n7057;
  assign n7059 = ~n7054 & ~n7058;
  assign n7060 = n7054 & n7058;
  assign n7061 = ~n6987 & ~n6989;
  assign n7062 = ~n6990 & ~n7061;
  assign n7063 = ~n5117 & ~n5119;
  assign n7064 = ~n5120 & ~n7063;
  assign n7065 = n7062 & n7064;
  assign n7066 = ~n6995 & ~n6996;
  assign n7067 = ~n7000 & n7066;
  assign n7068 = n7000 & ~n7066;
  assign n7069 = ~n7067 & ~n7068;
  assign n7070 = n7065 & n7069;
  assign n7071 = ~n7065 & ~n7069;
  assign n7072 = ~n5125 & ~n5126;
  assign n7073 = ~n5130 & n7072;
  assign n7074 = n5130 & ~n7072;
  assign n7075 = ~n7073 & ~n7074;
  assign n7076 = ~n7071 & n7075;
  assign n7077 = ~n7070 & ~n7076;
  assign n7078 = ~n7060 & n7077;
  assign n7079 = ~n7059 & ~n7078;
  assign n7080 = ~n7050 & n7079;
  assign n7081 = ~n7049 & ~n7080;
  assign n7082 = ~n7040 & n7081;
  assign n7083 = ~n7039 & ~n7082;
  assign n7084 = ~n7030 & n7083;
  assign n7085 = ~n7029 & ~n7084;
  assign n7086 = ~n7020 & ~n7085;
  assign n7087 = ~n7019 & ~n7086;
  assign n7088 = ~n7010 & ~n7012;
  assign n7089 = n7010 & n7012;
  assign n7090 = ~n6045 & ~n7089;
  assign n7091 = ~n7088 & ~n7090;
  assign n7092 = n7087 & ~n7091;
  assign n7093 = ~n7087 & n7091;
  assign n7094 = ~n4171 & ~n5142;
  assign n7095 = ~n5141 & ~n7094;
  assign n7096 = ~n7093 & ~n7095;
  assign n7097 = ~n7092 & ~n7096;
  assign n7098 = ~n3274 & ~n7097;
  assign n7099 = n3274 & n7097;
  assign n7100 = n2307 & n3204;
  assign n7101 = ~n2305 & ~n3273;
  assign n7102 = ~n3274 & ~n7101;
  assign n7103 = ~n7100 & ~n7102;
  assign n7104 = ~n7092 & ~n7093;
  assign n7105 = ~n7095 & ~n7104;
  assign n7106 = n7095 & n7104;
  assign n7107 = ~n7105 & ~n7106;
  assign n7108 = n7103 & ~n7107;
  assign n7109 = ~n7103 & n7107;
  assign n7110 = ~n3205 & ~n7100;
  assign n7111 = ~n3272 & n7110;
  assign n7112 = n3272 & ~n7110;
  assign n7113 = ~n7111 & ~n7112;
  assign n7114 = ~n7019 & ~n7020;
  assign n7115 = ~n7085 & n7114;
  assign n7116 = n7085 & ~n7114;
  assign n7117 = ~n7115 & ~n7116;
  assign n7118 = ~n7113 & ~n7117;
  assign n7119 = n7113 & n7117;
  assign n7120 = ~n7029 & ~n7030;
  assign n7121 = n7083 & n7120;
  assign n7122 = ~n7083 & ~n7120;
  assign n7123 = ~n7121 & ~n7122;
  assign n7124 = ~n3216 & ~n3217;
  assign n7125 = n3270 & n7124;
  assign n7126 = ~n3270 & ~n7124;
  assign n7127 = ~n7125 & ~n7126;
  assign n7128 = ~n7123 & ~n7127;
  assign n7129 = n7123 & n7127;
  assign n7130 = ~n3226 & ~n3227;
  assign n7131 = n3268 & n7130;
  assign n7132 = ~n3268 & ~n7130;
  assign n7133 = ~n7131 & ~n7132;
  assign n7134 = ~n7039 & ~n7040;
  assign n7135 = ~n7081 & n7134;
  assign n7136 = n7081 & ~n7134;
  assign n7137 = ~n7135 & ~n7136;
  assign n7138 = ~n7133 & ~n7137;
  assign n7139 = n7133 & n7137;
  assign n7140 = ~n7049 & ~n7050;
  assign n7141 = n7079 & n7140;
  assign n7142 = ~n7079 & ~n7140;
  assign n7143 = ~n7141 & ~n7142;
  assign n7144 = ~n3236 & ~n3237;
  assign n7145 = ~n3266 & n7144;
  assign n7146 = n3266 & ~n7144;
  assign n7147 = ~n7145 & ~n7146;
  assign n7148 = n7143 & ~n7147;
  assign n7149 = ~n7143 & n7147;
  assign n7150 = ~n3246 & ~n3247;
  assign n7151 = ~n3264 & n7150;
  assign n7152 = n3264 & ~n7150;
  assign n7153 = ~n7151 & ~n7152;
  assign n7154 = ~n7059 & ~n7060;
  assign n7155 = ~n7077 & n7154;
  assign n7156 = n7077 & ~n7154;
  assign n7157 = ~n7155 & ~n7156;
  assign n7158 = ~n7153 & ~n7157;
  assign n7159 = n7153 & n7157;
  assign n7160 = n7062 & ~n7064;
  assign n7161 = ~n7062 & n7064;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = ~n3249 & ~n3251;
  assign n7164 = ~n3252 & ~n7163;
  assign n7165 = ~n7162 & n7164;
  assign n7166 = ~n7070 & ~n7071;
  assign n7167 = ~n7075 & n7166;
  assign n7168 = n7075 & ~n7166;
  assign n7169 = ~n7167 & ~n7168;
  assign n7170 = n7165 & ~n7169;
  assign n7171 = ~n7165 & n7169;
  assign n7172 = ~n3257 & ~n3258;
  assign n7173 = ~n3262 & n7172;
  assign n7174 = n3262 & ~n7172;
  assign n7175 = ~n7173 & ~n7174;
  assign n7176 = ~n7171 & n7175;
  assign n7177 = ~n7170 & ~n7176;
  assign n7178 = ~n7159 & n7177;
  assign n7179 = ~n7158 & ~n7178;
  assign n7180 = ~n7149 & n7179;
  assign n7181 = ~n7148 & ~n7180;
  assign n7182 = ~n7139 & n7181;
  assign n7183 = ~n7138 & ~n7182;
  assign n7184 = ~n7129 & ~n7183;
  assign n7185 = ~n7128 & ~n7184;
  assign n7186 = ~n7119 & ~n7185;
  assign n7187 = ~n7118 & ~n7186;
  assign n7188 = ~n7109 & ~n7187;
  assign n7189 = ~n7108 & ~n7188;
  assign n7190 = ~n7099 & ~n7189;
  assign n7191 = ~n7098 & ~n7190;
  assign n7192 = ~pi466  & pi467 ;
  assign n7193 = pi466  & ~pi467 ;
  assign n7194 = pi468  & ~n7192;
  assign n7195 = ~n7193 & n7194;
  assign n7196 = ~n7192 & ~n7193;
  assign n7197 = ~pi468  & ~n7196;
  assign n7198 = ~n7195 & ~n7197;
  assign n7199 = ~pi463  & pi464 ;
  assign n7200 = pi463  & ~pi464 ;
  assign n7201 = pi465  & ~n7199;
  assign n7202 = ~n7200 & n7201;
  assign n7203 = ~n7199 & ~n7200;
  assign n7204 = ~pi465  & ~n7203;
  assign n7205 = ~n7202 & ~n7204;
  assign n7206 = ~n7198 & n7205;
  assign n7207 = n7198 & ~n7205;
  assign n7208 = ~n7206 & ~n7207;
  assign n7209 = ~pi469  & pi470 ;
  assign n7210 = pi469  & ~pi470 ;
  assign n7211 = pi471  & ~n7209;
  assign n7212 = ~n7210 & n7211;
  assign n7213 = ~n7209 & ~n7210;
  assign n7214 = ~pi471  & ~n7213;
  assign n7215 = ~n7212 & ~n7214;
  assign n7216 = ~pi472  & pi473 ;
  assign n7217 = pi472  & ~pi473 ;
  assign n7218 = pi474  & ~n7216;
  assign n7219 = ~n7217 & n7218;
  assign n7220 = ~n7216 & ~n7217;
  assign n7221 = ~pi474  & ~n7220;
  assign n7222 = ~n7219 & ~n7221;
  assign n7223 = ~n7215 & n7222;
  assign n7224 = n7215 & ~n7222;
  assign n7225 = ~n7223 & ~n7224;
  assign n7226 = ~n7208 & ~n7225;
  assign n7227 = n7208 & n7225;
  assign n7228 = ~n7226 & ~n7227;
  assign n7229 = ~pi481  & pi482 ;
  assign n7230 = pi481  & ~pi482 ;
  assign n7231 = pi483  & ~n7229;
  assign n7232 = ~n7230 & n7231;
  assign n7233 = ~n7229 & ~n7230;
  assign n7234 = ~pi483  & ~n7233;
  assign n7235 = ~n7232 & ~n7234;
  assign n7236 = ~pi484  & pi485 ;
  assign n7237 = pi484  & ~pi485 ;
  assign n7238 = pi486  & ~n7236;
  assign n7239 = ~n7237 & n7238;
  assign n7240 = ~n7236 & ~n7237;
  assign n7241 = ~pi486  & ~n7240;
  assign n7242 = ~n7239 & ~n7241;
  assign n7243 = ~n7235 & n7242;
  assign n7244 = n7235 & ~n7242;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = ~pi475  & pi476 ;
  assign n7247 = pi475  & ~pi476 ;
  assign n7248 = pi477  & ~n7246;
  assign n7249 = ~n7247 & n7248;
  assign n7250 = ~n7246 & ~n7247;
  assign n7251 = ~pi477  & ~n7250;
  assign n7252 = ~n7249 & ~n7251;
  assign n7253 = ~pi478  & pi479 ;
  assign n7254 = pi478  & ~pi479 ;
  assign n7255 = pi480  & ~n7253;
  assign n7256 = ~n7254 & n7255;
  assign n7257 = ~n7253 & ~n7254;
  assign n7258 = ~pi480  & ~n7257;
  assign n7259 = ~n7256 & ~n7258;
  assign n7260 = ~n7252 & n7259;
  assign n7261 = n7252 & ~n7259;
  assign n7262 = ~n7260 & ~n7261;
  assign n7263 = ~n7245 & ~n7262;
  assign n7264 = n7245 & n7262;
  assign n7265 = ~n7263 & ~n7264;
  assign n7266 = n7228 & n7265;
  assign n7267 = ~n7228 & ~n7265;
  assign n7268 = ~n7266 & ~n7267;
  assign n7269 = ~pi505  & pi506 ;
  assign n7270 = pi505  & ~pi506 ;
  assign n7271 = pi507  & ~n7269;
  assign n7272 = ~n7270 & n7271;
  assign n7273 = ~n7269 & ~n7270;
  assign n7274 = ~pi507  & ~n7273;
  assign n7275 = ~n7272 & ~n7274;
  assign n7276 = ~pi508  & pi509 ;
  assign n7277 = pi508  & ~pi509 ;
  assign n7278 = pi510  & ~n7276;
  assign n7279 = ~n7277 & n7278;
  assign n7280 = ~n7276 & ~n7277;
  assign n7281 = ~pi510  & ~n7280;
  assign n7282 = ~n7279 & ~n7281;
  assign n7283 = ~n7275 & n7282;
  assign n7284 = n7275 & ~n7282;
  assign n7285 = ~n7283 & ~n7284;
  assign n7286 = ~pi499  & pi500 ;
  assign n7287 = pi499  & ~pi500 ;
  assign n7288 = pi501  & ~n7286;
  assign n7289 = ~n7287 & n7288;
  assign n7290 = ~n7286 & ~n7287;
  assign n7291 = ~pi501  & ~n7290;
  assign n7292 = ~n7289 & ~n7291;
  assign n7293 = ~pi502  & pi503 ;
  assign n7294 = pi502  & ~pi503 ;
  assign n7295 = pi504  & ~n7293;
  assign n7296 = ~n7294 & n7295;
  assign n7297 = ~n7293 & ~n7294;
  assign n7298 = ~pi504  & ~n7297;
  assign n7299 = ~n7296 & ~n7298;
  assign n7300 = ~n7292 & n7299;
  assign n7301 = n7292 & ~n7299;
  assign n7302 = ~n7300 & ~n7301;
  assign n7303 = ~n7285 & ~n7302;
  assign n7304 = n7285 & n7302;
  assign n7305 = ~n7303 & ~n7304;
  assign n7306 = ~pi493  & pi494 ;
  assign n7307 = pi493  & ~pi494 ;
  assign n7308 = pi495  & ~n7306;
  assign n7309 = ~n7307 & n7308;
  assign n7310 = ~n7306 & ~n7307;
  assign n7311 = ~pi495  & ~n7310;
  assign n7312 = ~n7309 & ~n7311;
  assign n7313 = ~pi496  & pi497 ;
  assign n7314 = pi496  & ~pi497 ;
  assign n7315 = pi498  & ~n7313;
  assign n7316 = ~n7314 & n7315;
  assign n7317 = ~n7313 & ~n7314;
  assign n7318 = ~pi498  & ~n7317;
  assign n7319 = ~n7316 & ~n7318;
  assign n7320 = ~n7312 & n7319;
  assign n7321 = n7312 & ~n7319;
  assign n7322 = ~n7320 & ~n7321;
  assign n7323 = ~pi487  & pi488 ;
  assign n7324 = pi487  & ~pi488 ;
  assign n7325 = pi489  & ~n7323;
  assign n7326 = ~n7324 & n7325;
  assign n7327 = ~n7323 & ~n7324;
  assign n7328 = ~pi489  & ~n7327;
  assign n7329 = ~n7326 & ~n7328;
  assign n7330 = ~pi490  & pi491 ;
  assign n7331 = pi490  & ~pi491 ;
  assign n7332 = pi492  & ~n7330;
  assign n7333 = ~n7331 & n7332;
  assign n7334 = ~n7330 & ~n7331;
  assign n7335 = ~pi492  & ~n7334;
  assign n7336 = ~n7333 & ~n7335;
  assign n7337 = ~n7329 & n7336;
  assign n7338 = n7329 & ~n7336;
  assign n7339 = ~n7337 & ~n7338;
  assign n7340 = ~n7322 & ~n7339;
  assign n7341 = n7322 & n7339;
  assign n7342 = ~n7340 & ~n7341;
  assign n7343 = n7305 & n7342;
  assign n7344 = ~n7305 & ~n7342;
  assign n7345 = ~n7343 & ~n7344;
  assign n7346 = n7268 & ~n7345;
  assign n7347 = ~n7268 & n7345;
  assign n7348 = ~n7346 & ~n7347;
  assign n7349 = ~pi553  & pi554 ;
  assign n7350 = pi553  & ~pi554 ;
  assign n7351 = pi555  & ~n7349;
  assign n7352 = ~n7350 & n7351;
  assign n7353 = ~n7349 & ~n7350;
  assign n7354 = ~pi555  & ~n7353;
  assign n7355 = ~n7352 & ~n7354;
  assign n7356 = ~pi556  & pi557 ;
  assign n7357 = pi556  & ~pi557 ;
  assign n7358 = pi558  & ~n7356;
  assign n7359 = ~n7357 & n7358;
  assign n7360 = ~n7356 & ~n7357;
  assign n7361 = ~pi558  & ~n7360;
  assign n7362 = ~n7359 & ~n7361;
  assign n7363 = ~n7355 & n7362;
  assign n7364 = n7355 & ~n7362;
  assign n7365 = ~n7363 & ~n7364;
  assign n7366 = ~pi547  & pi548 ;
  assign n7367 = pi547  & ~pi548 ;
  assign n7368 = pi549  & ~n7366;
  assign n7369 = ~n7367 & n7368;
  assign n7370 = ~n7366 & ~n7367;
  assign n7371 = ~pi549  & ~n7370;
  assign n7372 = ~n7369 & ~n7371;
  assign n7373 = ~pi550  & pi551 ;
  assign n7374 = pi550  & ~pi551 ;
  assign n7375 = pi552  & ~n7373;
  assign n7376 = ~n7374 & n7375;
  assign n7377 = ~n7373 & ~n7374;
  assign n7378 = ~pi552  & ~n7377;
  assign n7379 = ~n7376 & ~n7378;
  assign n7380 = ~n7372 & n7379;
  assign n7381 = n7372 & ~n7379;
  assign n7382 = ~n7380 & ~n7381;
  assign n7383 = ~n7365 & ~n7382;
  assign n7384 = n7365 & n7382;
  assign n7385 = ~n7383 & ~n7384;
  assign n7386 = ~pi541  & pi542 ;
  assign n7387 = pi541  & ~pi542 ;
  assign n7388 = pi543  & ~n7386;
  assign n7389 = ~n7387 & n7388;
  assign n7390 = ~n7386 & ~n7387;
  assign n7391 = ~pi543  & ~n7390;
  assign n7392 = ~n7389 & ~n7391;
  assign n7393 = ~pi544  & pi545 ;
  assign n7394 = pi544  & ~pi545 ;
  assign n7395 = pi546  & ~n7393;
  assign n7396 = ~n7394 & n7395;
  assign n7397 = ~n7393 & ~n7394;
  assign n7398 = ~pi546  & ~n7397;
  assign n7399 = ~n7396 & ~n7398;
  assign n7400 = ~n7392 & n7399;
  assign n7401 = n7392 & ~n7399;
  assign n7402 = ~n7400 & ~n7401;
  assign n7403 = ~pi535  & pi536 ;
  assign n7404 = pi535  & ~pi536 ;
  assign n7405 = pi537  & ~n7403;
  assign n7406 = ~n7404 & n7405;
  assign n7407 = ~n7403 & ~n7404;
  assign n7408 = ~pi537  & ~n7407;
  assign n7409 = ~n7406 & ~n7408;
  assign n7410 = ~pi538  & pi539 ;
  assign n7411 = pi538  & ~pi539 ;
  assign n7412 = pi540  & ~n7410;
  assign n7413 = ~n7411 & n7412;
  assign n7414 = ~n7410 & ~n7411;
  assign n7415 = ~pi540  & ~n7414;
  assign n7416 = ~n7413 & ~n7415;
  assign n7417 = ~n7409 & n7416;
  assign n7418 = n7409 & ~n7416;
  assign n7419 = ~n7417 & ~n7418;
  assign n7420 = ~n7402 & ~n7419;
  assign n7421 = n7402 & n7419;
  assign n7422 = ~n7420 & ~n7421;
  assign n7423 = n7385 & n7422;
  assign n7424 = ~n7385 & ~n7422;
  assign n7425 = ~n7423 & ~n7424;
  assign n7426 = ~pi529  & pi530 ;
  assign n7427 = pi529  & ~pi530 ;
  assign n7428 = pi531  & ~n7426;
  assign n7429 = ~n7427 & n7428;
  assign n7430 = ~n7426 & ~n7427;
  assign n7431 = ~pi531  & ~n7430;
  assign n7432 = ~n7429 & ~n7431;
  assign n7433 = ~pi532  & pi533 ;
  assign n7434 = pi532  & ~pi533 ;
  assign n7435 = pi534  & ~n7433;
  assign n7436 = ~n7434 & n7435;
  assign n7437 = ~n7433 & ~n7434;
  assign n7438 = ~pi534  & ~n7437;
  assign n7439 = ~n7436 & ~n7438;
  assign n7440 = ~n7432 & n7439;
  assign n7441 = n7432 & ~n7439;
  assign n7442 = ~n7440 & ~n7441;
  assign n7443 = ~pi523  & pi524 ;
  assign n7444 = pi523  & ~pi524 ;
  assign n7445 = pi525  & ~n7443;
  assign n7446 = ~n7444 & n7445;
  assign n7447 = ~n7443 & ~n7444;
  assign n7448 = ~pi525  & ~n7447;
  assign n7449 = ~n7446 & ~n7448;
  assign n7450 = ~pi526  & pi527 ;
  assign n7451 = pi526  & ~pi527 ;
  assign n7452 = pi528  & ~n7450;
  assign n7453 = ~n7451 & n7452;
  assign n7454 = ~n7450 & ~n7451;
  assign n7455 = ~pi528  & ~n7454;
  assign n7456 = ~n7453 & ~n7455;
  assign n7457 = ~n7449 & n7456;
  assign n7458 = n7449 & ~n7456;
  assign n7459 = ~n7457 & ~n7458;
  assign n7460 = ~n7442 & ~n7459;
  assign n7461 = n7442 & n7459;
  assign n7462 = ~n7460 & ~n7461;
  assign n7463 = ~pi517  & pi518 ;
  assign n7464 = pi517  & ~pi518 ;
  assign n7465 = pi519  & ~n7463;
  assign n7466 = ~n7464 & n7465;
  assign n7467 = ~n7463 & ~n7464;
  assign n7468 = ~pi519  & ~n7467;
  assign n7469 = ~n7466 & ~n7468;
  assign n7470 = ~pi520  & pi521 ;
  assign n7471 = pi520  & ~pi521 ;
  assign n7472 = pi522  & ~n7470;
  assign n7473 = ~n7471 & n7472;
  assign n7474 = ~n7470 & ~n7471;
  assign n7475 = ~pi522  & ~n7474;
  assign n7476 = ~n7473 & ~n7475;
  assign n7477 = ~n7469 & n7476;
  assign n7478 = n7469 & ~n7476;
  assign n7479 = ~n7477 & ~n7478;
  assign n7480 = ~pi511  & pi512 ;
  assign n7481 = pi511  & ~pi512 ;
  assign n7482 = pi513  & ~n7480;
  assign n7483 = ~n7481 & n7482;
  assign n7484 = ~n7480 & ~n7481;
  assign n7485 = ~pi513  & ~n7484;
  assign n7486 = ~n7483 & ~n7485;
  assign n7487 = ~pi514  & pi515 ;
  assign n7488 = pi514  & ~pi515 ;
  assign n7489 = pi516  & ~n7487;
  assign n7490 = ~n7488 & n7489;
  assign n7491 = ~n7487 & ~n7488;
  assign n7492 = ~pi516  & ~n7491;
  assign n7493 = ~n7490 & ~n7492;
  assign n7494 = ~n7486 & n7493;
  assign n7495 = n7486 & ~n7493;
  assign n7496 = ~n7494 & ~n7495;
  assign n7497 = ~n7479 & ~n7496;
  assign n7498 = n7479 & n7496;
  assign n7499 = ~n7497 & ~n7498;
  assign n7500 = n7462 & n7499;
  assign n7501 = ~n7462 & ~n7499;
  assign n7502 = ~n7500 & ~n7501;
  assign n7503 = n7425 & ~n7502;
  assign n7504 = ~n7425 & n7502;
  assign n7505 = ~n7503 & ~n7504;
  assign n7506 = ~n7348 & ~n7505;
  assign n7507 = n7348 & n7505;
  assign n7508 = ~n7506 & ~n7507;
  assign n7509 = ~pi649  & pi650 ;
  assign n7510 = pi649  & ~pi650 ;
  assign n7511 = pi651  & ~n7509;
  assign n7512 = ~n7510 & n7511;
  assign n7513 = ~n7509 & ~n7510;
  assign n7514 = ~pi651  & ~n7513;
  assign n7515 = ~n7512 & ~n7514;
  assign n7516 = ~pi652  & pi653 ;
  assign n7517 = pi652  & ~pi653 ;
  assign n7518 = pi654  & ~n7516;
  assign n7519 = ~n7517 & n7518;
  assign n7520 = ~n7516 & ~n7517;
  assign n7521 = ~pi654  & ~n7520;
  assign n7522 = ~n7519 & ~n7521;
  assign n7523 = ~n7515 & n7522;
  assign n7524 = n7515 & ~n7522;
  assign n7525 = ~n7523 & ~n7524;
  assign n7526 = ~pi643  & pi644 ;
  assign n7527 = pi643  & ~pi644 ;
  assign n7528 = pi645  & ~n7526;
  assign n7529 = ~n7527 & n7528;
  assign n7530 = ~n7526 & ~n7527;
  assign n7531 = ~pi645  & ~n7530;
  assign n7532 = ~n7529 & ~n7531;
  assign n7533 = ~pi646  & pi647 ;
  assign n7534 = pi646  & ~pi647 ;
  assign n7535 = pi648  & ~n7533;
  assign n7536 = ~n7534 & n7535;
  assign n7537 = ~n7533 & ~n7534;
  assign n7538 = ~pi648  & ~n7537;
  assign n7539 = ~n7536 & ~n7538;
  assign n7540 = ~n7532 & n7539;
  assign n7541 = n7532 & ~n7539;
  assign n7542 = ~n7540 & ~n7541;
  assign n7543 = ~n7525 & ~n7542;
  assign n7544 = n7525 & n7542;
  assign n7545 = ~n7543 & ~n7544;
  assign n7546 = ~pi637  & pi638 ;
  assign n7547 = pi637  & ~pi638 ;
  assign n7548 = pi639  & ~n7546;
  assign n7549 = ~n7547 & n7548;
  assign n7550 = ~n7546 & ~n7547;
  assign n7551 = ~pi639  & ~n7550;
  assign n7552 = ~n7549 & ~n7551;
  assign n7553 = ~pi640  & pi641 ;
  assign n7554 = pi640  & ~pi641 ;
  assign n7555 = pi642  & ~n7553;
  assign n7556 = ~n7554 & n7555;
  assign n7557 = ~n7553 & ~n7554;
  assign n7558 = ~pi642  & ~n7557;
  assign n7559 = ~n7556 & ~n7558;
  assign n7560 = ~n7552 & n7559;
  assign n7561 = n7552 & ~n7559;
  assign n7562 = ~n7560 & ~n7561;
  assign n7563 = ~pi631  & pi632 ;
  assign n7564 = pi631  & ~pi632 ;
  assign n7565 = pi633  & ~n7563;
  assign n7566 = ~n7564 & n7565;
  assign n7567 = ~n7563 & ~n7564;
  assign n7568 = ~pi633  & ~n7567;
  assign n7569 = ~n7566 & ~n7568;
  assign n7570 = ~pi634  & pi635 ;
  assign n7571 = pi634  & ~pi635 ;
  assign n7572 = pi636  & ~n7570;
  assign n7573 = ~n7571 & n7572;
  assign n7574 = ~n7570 & ~n7571;
  assign n7575 = ~pi636  & ~n7574;
  assign n7576 = ~n7573 & ~n7575;
  assign n7577 = ~n7569 & n7576;
  assign n7578 = n7569 & ~n7576;
  assign n7579 = ~n7577 & ~n7578;
  assign n7580 = ~n7562 & ~n7579;
  assign n7581 = n7562 & n7579;
  assign n7582 = ~n7580 & ~n7581;
  assign n7583 = n7545 & n7582;
  assign n7584 = ~n7545 & ~n7582;
  assign n7585 = ~n7583 & ~n7584;
  assign n7586 = ~pi625  & pi626 ;
  assign n7587 = pi625  & ~pi626 ;
  assign n7588 = pi627  & ~n7586;
  assign n7589 = ~n7587 & n7588;
  assign n7590 = ~n7586 & ~n7587;
  assign n7591 = ~pi627  & ~n7590;
  assign n7592 = ~n7589 & ~n7591;
  assign n7593 = ~pi628  & pi629 ;
  assign n7594 = pi628  & ~pi629 ;
  assign n7595 = pi630  & ~n7593;
  assign n7596 = ~n7594 & n7595;
  assign n7597 = ~n7593 & ~n7594;
  assign n7598 = ~pi630  & ~n7597;
  assign n7599 = ~n7596 & ~n7598;
  assign n7600 = ~n7592 & n7599;
  assign n7601 = n7592 & ~n7599;
  assign n7602 = ~n7600 & ~n7601;
  assign n7603 = ~pi619  & pi620 ;
  assign n7604 = pi619  & ~pi620 ;
  assign n7605 = pi621  & ~n7603;
  assign n7606 = ~n7604 & n7605;
  assign n7607 = ~n7603 & ~n7604;
  assign n7608 = ~pi621  & ~n7607;
  assign n7609 = ~n7606 & ~n7608;
  assign n7610 = ~pi622  & pi623 ;
  assign n7611 = pi622  & ~pi623 ;
  assign n7612 = pi624  & ~n7610;
  assign n7613 = ~n7611 & n7612;
  assign n7614 = ~n7610 & ~n7611;
  assign n7615 = ~pi624  & ~n7614;
  assign n7616 = ~n7613 & ~n7615;
  assign n7617 = ~n7609 & n7616;
  assign n7618 = n7609 & ~n7616;
  assign n7619 = ~n7617 & ~n7618;
  assign n7620 = ~n7602 & ~n7619;
  assign n7621 = n7602 & n7619;
  assign n7622 = ~n7620 & ~n7621;
  assign n7623 = ~pi613  & pi614 ;
  assign n7624 = pi613  & ~pi614 ;
  assign n7625 = pi615  & ~n7623;
  assign n7626 = ~n7624 & n7625;
  assign n7627 = ~n7623 & ~n7624;
  assign n7628 = ~pi615  & ~n7627;
  assign n7629 = ~n7626 & ~n7628;
  assign n7630 = ~pi616  & pi617 ;
  assign n7631 = pi616  & ~pi617 ;
  assign n7632 = pi618  & ~n7630;
  assign n7633 = ~n7631 & n7632;
  assign n7634 = ~n7630 & ~n7631;
  assign n7635 = ~pi618  & ~n7634;
  assign n7636 = ~n7633 & ~n7635;
  assign n7637 = ~n7629 & n7636;
  assign n7638 = n7629 & ~n7636;
  assign n7639 = ~n7637 & ~n7638;
  assign n7640 = ~pi607  & pi608 ;
  assign n7641 = pi607  & ~pi608 ;
  assign n7642 = pi609  & ~n7640;
  assign n7643 = ~n7641 & n7642;
  assign n7644 = ~n7640 & ~n7641;
  assign n7645 = ~pi609  & ~n7644;
  assign n7646 = ~n7643 & ~n7645;
  assign n7647 = ~pi610  & pi611 ;
  assign n7648 = pi610  & ~pi611 ;
  assign n7649 = pi612  & ~n7647;
  assign n7650 = ~n7648 & n7649;
  assign n7651 = ~n7647 & ~n7648;
  assign n7652 = ~pi612  & ~n7651;
  assign n7653 = ~n7650 & ~n7652;
  assign n7654 = ~n7646 & n7653;
  assign n7655 = n7646 & ~n7653;
  assign n7656 = ~n7654 & ~n7655;
  assign n7657 = ~n7639 & ~n7656;
  assign n7658 = n7639 & n7656;
  assign n7659 = ~n7657 & ~n7658;
  assign n7660 = n7622 & n7659;
  assign n7661 = ~n7622 & ~n7659;
  assign n7662 = ~n7660 & ~n7661;
  assign n7663 = n7585 & ~n7662;
  assign n7664 = ~n7585 & n7662;
  assign n7665 = ~n7663 & ~n7664;
  assign n7666 = ~pi601  & pi602 ;
  assign n7667 = pi601  & ~pi602 ;
  assign n7668 = pi603  & ~n7666;
  assign n7669 = ~n7667 & n7668;
  assign n7670 = ~n7666 & ~n7667;
  assign n7671 = ~pi603  & ~n7670;
  assign n7672 = ~n7669 & ~n7671;
  assign n7673 = ~pi604  & pi605 ;
  assign n7674 = pi604  & ~pi605 ;
  assign n7675 = pi606  & ~n7673;
  assign n7676 = ~n7674 & n7675;
  assign n7677 = ~n7673 & ~n7674;
  assign n7678 = ~pi606  & ~n7677;
  assign n7679 = ~n7676 & ~n7678;
  assign n7680 = ~n7672 & n7679;
  assign n7681 = n7672 & ~n7679;
  assign n7682 = ~n7680 & ~n7681;
  assign n7683 = ~pi595  & pi596 ;
  assign n7684 = pi595  & ~pi596 ;
  assign n7685 = pi597  & ~n7683;
  assign n7686 = ~n7684 & n7685;
  assign n7687 = ~n7683 & ~n7684;
  assign n7688 = ~pi597  & ~n7687;
  assign n7689 = ~n7686 & ~n7688;
  assign n7690 = ~pi598  & pi599 ;
  assign n7691 = pi598  & ~pi599 ;
  assign n7692 = pi600  & ~n7690;
  assign n7693 = ~n7691 & n7692;
  assign n7694 = ~n7690 & ~n7691;
  assign n7695 = ~pi600  & ~n7694;
  assign n7696 = ~n7693 & ~n7695;
  assign n7697 = ~n7689 & n7696;
  assign n7698 = n7689 & ~n7696;
  assign n7699 = ~n7697 & ~n7698;
  assign n7700 = ~n7682 & ~n7699;
  assign n7701 = n7682 & n7699;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = ~pi589  & pi590 ;
  assign n7704 = pi589  & ~pi590 ;
  assign n7705 = pi591  & ~n7703;
  assign n7706 = ~n7704 & n7705;
  assign n7707 = ~n7703 & ~n7704;
  assign n7708 = ~pi591  & ~n7707;
  assign n7709 = ~n7706 & ~n7708;
  assign n7710 = ~pi592  & pi593 ;
  assign n7711 = pi592  & ~pi593 ;
  assign n7712 = pi594  & ~n7710;
  assign n7713 = ~n7711 & n7712;
  assign n7714 = ~n7710 & ~n7711;
  assign n7715 = ~pi594  & ~n7714;
  assign n7716 = ~n7713 & ~n7715;
  assign n7717 = ~n7709 & n7716;
  assign n7718 = n7709 & ~n7716;
  assign n7719 = ~n7717 & ~n7718;
  assign n7720 = ~pi583  & pi584 ;
  assign n7721 = pi583  & ~pi584 ;
  assign n7722 = pi585  & ~n7720;
  assign n7723 = ~n7721 & n7722;
  assign n7724 = ~n7720 & ~n7721;
  assign n7725 = ~pi585  & ~n7724;
  assign n7726 = ~n7723 & ~n7725;
  assign n7727 = ~pi586  & pi587 ;
  assign n7728 = pi586  & ~pi587 ;
  assign n7729 = pi588  & ~n7727;
  assign n7730 = ~n7728 & n7729;
  assign n7731 = ~n7727 & ~n7728;
  assign n7732 = ~pi588  & ~n7731;
  assign n7733 = ~n7730 & ~n7732;
  assign n7734 = ~n7726 & n7733;
  assign n7735 = n7726 & ~n7733;
  assign n7736 = ~n7734 & ~n7735;
  assign n7737 = ~n7719 & ~n7736;
  assign n7738 = n7719 & n7736;
  assign n7739 = ~n7737 & ~n7738;
  assign n7740 = n7702 & n7739;
  assign n7741 = ~n7702 & ~n7739;
  assign n7742 = ~n7740 & ~n7741;
  assign n7743 = ~pi577  & pi578 ;
  assign n7744 = pi577  & ~pi578 ;
  assign n7745 = pi579  & ~n7743;
  assign n7746 = ~n7744 & n7745;
  assign n7747 = ~n7743 & ~n7744;
  assign n7748 = ~pi579  & ~n7747;
  assign n7749 = ~n7746 & ~n7748;
  assign n7750 = ~pi580  & pi581 ;
  assign n7751 = pi580  & ~pi581 ;
  assign n7752 = pi582  & ~n7750;
  assign n7753 = ~n7751 & n7752;
  assign n7754 = ~n7750 & ~n7751;
  assign n7755 = ~pi582  & ~n7754;
  assign n7756 = ~n7753 & ~n7755;
  assign n7757 = ~n7749 & n7756;
  assign n7758 = n7749 & ~n7756;
  assign n7759 = ~n7757 & ~n7758;
  assign n7760 = ~pi571  & pi572 ;
  assign n7761 = pi571  & ~pi572 ;
  assign n7762 = pi573  & ~n7760;
  assign n7763 = ~n7761 & n7762;
  assign n7764 = ~n7760 & ~n7761;
  assign n7765 = ~pi573  & ~n7764;
  assign n7766 = ~n7763 & ~n7765;
  assign n7767 = ~pi574  & pi575 ;
  assign n7768 = pi574  & ~pi575 ;
  assign n7769 = pi576  & ~n7767;
  assign n7770 = ~n7768 & n7769;
  assign n7771 = ~n7767 & ~n7768;
  assign n7772 = ~pi576  & ~n7771;
  assign n7773 = ~n7770 & ~n7772;
  assign n7774 = ~n7766 & n7773;
  assign n7775 = n7766 & ~n7773;
  assign n7776 = ~n7774 & ~n7775;
  assign n7777 = ~n7759 & ~n7776;
  assign n7778 = n7759 & n7776;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = ~pi565  & pi566 ;
  assign n7781 = pi565  & ~pi566 ;
  assign n7782 = pi567  & ~n7780;
  assign n7783 = ~n7781 & n7782;
  assign n7784 = ~n7780 & ~n7781;
  assign n7785 = ~pi567  & ~n7784;
  assign n7786 = ~n7783 & ~n7785;
  assign n7787 = ~pi568  & pi569 ;
  assign n7788 = pi568  & ~pi569 ;
  assign n7789 = pi570  & ~n7787;
  assign n7790 = ~n7788 & n7789;
  assign n7791 = ~n7787 & ~n7788;
  assign n7792 = ~pi570  & ~n7791;
  assign n7793 = ~n7790 & ~n7792;
  assign n7794 = ~n7786 & n7793;
  assign n7795 = n7786 & ~n7793;
  assign n7796 = ~n7794 & ~n7795;
  assign n7797 = ~pi559  & pi560 ;
  assign n7798 = pi559  & ~pi560 ;
  assign n7799 = pi561  & ~n7797;
  assign n7800 = ~n7798 & n7799;
  assign n7801 = ~n7797 & ~n7798;
  assign n7802 = ~pi561  & ~n7801;
  assign n7803 = ~n7800 & ~n7802;
  assign n7804 = ~pi562  & pi563 ;
  assign n7805 = pi562  & ~pi563 ;
  assign n7806 = pi564  & ~n7804;
  assign n7807 = ~n7805 & n7806;
  assign n7808 = ~n7804 & ~n7805;
  assign n7809 = ~pi564  & ~n7808;
  assign n7810 = ~n7807 & ~n7809;
  assign n7811 = ~n7803 & n7810;
  assign n7812 = n7803 & ~n7810;
  assign n7813 = ~n7811 & ~n7812;
  assign n7814 = ~n7796 & ~n7813;
  assign n7815 = n7796 & n7813;
  assign n7816 = ~n7814 & ~n7815;
  assign n7817 = n7779 & n7816;
  assign n7818 = ~n7779 & ~n7816;
  assign n7819 = ~n7817 & ~n7818;
  assign n7820 = n7742 & ~n7819;
  assign n7821 = ~n7742 & n7819;
  assign n7822 = ~n7820 & ~n7821;
  assign n7823 = ~n7665 & ~n7822;
  assign n7824 = n7665 & n7822;
  assign n7825 = ~n7823 & ~n7824;
  assign n7826 = n7508 & n7825;
  assign n7827 = ~n7508 & ~n7825;
  assign n7828 = ~n7826 & ~n7827;
  assign n7829 = pi835  & ~pi836 ;
  assign n7830 = ~pi835  & pi836 ;
  assign n7831 = pi837  & ~n7829;
  assign n7832 = ~n7830 & n7831;
  assign n7833 = ~n7829 & ~n7830;
  assign n7834 = ~pi837  & ~n7833;
  assign n7835 = ~n7832 & ~n7834;
  assign n7836 = pi838  & ~pi839 ;
  assign n7837 = ~pi838  & pi839 ;
  assign n7838 = pi840  & ~n7836;
  assign n7839 = ~n7837 & n7838;
  assign n7840 = ~n7836 & ~n7837;
  assign n7841 = ~pi840  & ~n7840;
  assign n7842 = ~n7839 & ~n7841;
  assign n7843 = ~n7835 & n7842;
  assign n7844 = n7835 & ~n7842;
  assign n7845 = ~n7843 & ~n7844;
  assign n7846 = pi841  & ~pi842 ;
  assign n7847 = ~pi841  & pi842 ;
  assign n7848 = pi843  & ~n7846;
  assign n7849 = ~n7847 & n7848;
  assign n7850 = ~n7846 & ~n7847;
  assign n7851 = ~pi843  & ~n7850;
  assign n7852 = ~n7849 & ~n7851;
  assign n7853 = pi844  & ~pi845 ;
  assign n7854 = ~pi844  & pi845 ;
  assign n7855 = pi846  & ~n7853;
  assign n7856 = ~n7854 & n7855;
  assign n7857 = ~n7853 & ~n7854;
  assign n7858 = ~pi846  & ~n7857;
  assign n7859 = ~n7856 & ~n7858;
  assign n7860 = ~n7852 & n7859;
  assign n7861 = n7852 & ~n7859;
  assign n7862 = ~n7860 & ~n7861;
  assign n7863 = ~n7845 & ~n7862;
  assign n7864 = n7845 & n7862;
  assign n7865 = ~n7863 & ~n7864;
  assign n7866 = pi823  & ~pi824 ;
  assign n7867 = ~pi823  & pi824 ;
  assign n7868 = pi825  & ~n7866;
  assign n7869 = ~n7867 & n7868;
  assign n7870 = ~n7866 & ~n7867;
  assign n7871 = ~pi825  & ~n7870;
  assign n7872 = ~n7869 & ~n7871;
  assign n7873 = pi826  & ~pi827 ;
  assign n7874 = ~pi826  & pi827 ;
  assign n7875 = pi828  & ~n7873;
  assign n7876 = ~n7874 & n7875;
  assign n7877 = ~n7873 & ~n7874;
  assign n7878 = ~pi828  & ~n7877;
  assign n7879 = ~n7876 & ~n7878;
  assign n7880 = ~n7872 & n7879;
  assign n7881 = n7872 & ~n7879;
  assign n7882 = ~n7880 & ~n7881;
  assign n7883 = pi829  & ~pi830 ;
  assign n7884 = ~pi829  & pi830 ;
  assign n7885 = pi831  & ~n7883;
  assign n7886 = ~n7884 & n7885;
  assign n7887 = ~n7883 & ~n7884;
  assign n7888 = ~pi831  & ~n7887;
  assign n7889 = ~n7886 & ~n7888;
  assign n7890 = pi832  & ~pi833 ;
  assign n7891 = ~pi832  & pi833 ;
  assign n7892 = pi834  & ~n7890;
  assign n7893 = ~n7891 & n7892;
  assign n7894 = ~n7890 & ~n7891;
  assign n7895 = ~pi834  & ~n7894;
  assign n7896 = ~n7893 & ~n7895;
  assign n7897 = ~n7889 & n7896;
  assign n7898 = n7889 & ~n7896;
  assign n7899 = ~n7897 & ~n7898;
  assign n7900 = ~n7882 & ~n7899;
  assign n7901 = n7882 & n7899;
  assign n7902 = ~n7900 & ~n7901;
  assign n7903 = n7865 & n7902;
  assign n7904 = ~n7865 & ~n7902;
  assign n7905 = ~n7903 & ~n7904;
  assign n7906 = pi811  & ~pi812 ;
  assign n7907 = ~pi811  & pi812 ;
  assign n7908 = pi813  & ~n7906;
  assign n7909 = ~n7907 & n7908;
  assign n7910 = ~n7906 & ~n7907;
  assign n7911 = ~pi813  & ~n7910;
  assign n7912 = ~n7909 & ~n7911;
  assign n7913 = pi814  & ~pi815 ;
  assign n7914 = ~pi814  & pi815 ;
  assign n7915 = pi816  & ~n7913;
  assign n7916 = ~n7914 & n7915;
  assign n7917 = ~n7913 & ~n7914;
  assign n7918 = ~pi816  & ~n7917;
  assign n7919 = ~n7916 & ~n7918;
  assign n7920 = ~n7912 & n7919;
  assign n7921 = n7912 & ~n7919;
  assign n7922 = ~n7920 & ~n7921;
  assign n7923 = pi817  & ~pi818 ;
  assign n7924 = ~pi817  & pi818 ;
  assign n7925 = pi819  & ~n7923;
  assign n7926 = ~n7924 & n7925;
  assign n7927 = ~n7923 & ~n7924;
  assign n7928 = ~pi819  & ~n7927;
  assign n7929 = ~n7926 & ~n7928;
  assign n7930 = pi820  & ~pi821 ;
  assign n7931 = ~pi820  & pi821 ;
  assign n7932 = pi822  & ~n7930;
  assign n7933 = ~n7931 & n7932;
  assign n7934 = ~n7930 & ~n7931;
  assign n7935 = ~pi822  & ~n7934;
  assign n7936 = ~n7933 & ~n7935;
  assign n7937 = ~n7929 & n7936;
  assign n7938 = n7929 & ~n7936;
  assign n7939 = ~n7937 & ~n7938;
  assign n7940 = ~n7922 & ~n7939;
  assign n7941 = n7922 & n7939;
  assign n7942 = ~n7940 & ~n7941;
  assign n7943 = ~pi805  & pi806 ;
  assign n7944 = pi805  & ~pi806 ;
  assign n7945 = pi807  & ~n7943;
  assign n7946 = ~n7944 & n7945;
  assign n7947 = ~n7943 & ~n7944;
  assign n7948 = ~pi807  & ~n7947;
  assign n7949 = ~n7946 & ~n7948;
  assign n7950 = ~pi808  & pi809 ;
  assign n7951 = pi808  & ~pi809 ;
  assign n7952 = pi810  & ~n7950;
  assign n7953 = ~n7951 & n7952;
  assign n7954 = ~n7950 & ~n7951;
  assign n7955 = ~pi810  & ~n7954;
  assign n7956 = ~n7953 & ~n7955;
  assign n7957 = ~n7949 & n7956;
  assign n7958 = n7949 & ~n7956;
  assign n7959 = ~n7957 & ~n7958;
  assign n7960 = ~pi799  & pi800 ;
  assign n7961 = pi799  & ~pi800 ;
  assign n7962 = pi801  & ~n7960;
  assign n7963 = ~n7961 & n7962;
  assign n7964 = ~n7960 & ~n7961;
  assign n7965 = ~pi801  & ~n7964;
  assign n7966 = ~n7963 & ~n7965;
  assign n7967 = ~pi802  & pi803 ;
  assign n7968 = pi802  & ~pi803 ;
  assign n7969 = pi804  & ~n7967;
  assign n7970 = ~n7968 & n7969;
  assign n7971 = ~n7967 & ~n7968;
  assign n7972 = ~pi804  & ~n7971;
  assign n7973 = ~n7970 & ~n7972;
  assign n7974 = ~n7966 & n7973;
  assign n7975 = n7966 & ~n7973;
  assign n7976 = ~n7974 & ~n7975;
  assign n7977 = ~n7959 & ~n7976;
  assign n7978 = n7959 & n7976;
  assign n7979 = ~n7977 & ~n7978;
  assign n7980 = n7942 & n7979;
  assign n7981 = ~n7942 & ~n7979;
  assign n7982 = ~n7980 & ~n7981;
  assign n7983 = n7905 & ~n7982;
  assign n7984 = ~n7905 & n7982;
  assign n7985 = ~n7983 & ~n7984;
  assign n7986 = pi787  & ~pi788 ;
  assign n7987 = ~pi787  & pi788 ;
  assign n7988 = pi789  & ~n7986;
  assign n7989 = ~n7987 & n7988;
  assign n7990 = ~n7986 & ~n7987;
  assign n7991 = ~pi789  & ~n7990;
  assign n7992 = ~n7989 & ~n7991;
  assign n7993 = pi790  & ~pi791 ;
  assign n7994 = ~pi790  & pi791 ;
  assign n7995 = pi792  & ~n7993;
  assign n7996 = ~n7994 & n7995;
  assign n7997 = ~n7993 & ~n7994;
  assign n7998 = ~pi792  & ~n7997;
  assign n7999 = ~n7996 & ~n7998;
  assign n8000 = ~n7992 & n7999;
  assign n8001 = n7992 & ~n7999;
  assign n8002 = ~n8000 & ~n8001;
  assign n8003 = pi793  & ~pi794 ;
  assign n8004 = ~pi793  & pi794 ;
  assign n8005 = pi795  & ~n8003;
  assign n8006 = ~n8004 & n8005;
  assign n8007 = ~n8003 & ~n8004;
  assign n8008 = ~pi795  & ~n8007;
  assign n8009 = ~n8006 & ~n8008;
  assign n8010 = pi796  & ~pi797 ;
  assign n8011 = ~pi796  & pi797 ;
  assign n8012 = pi798  & ~n8010;
  assign n8013 = ~n8011 & n8012;
  assign n8014 = ~n8010 & ~n8011;
  assign n8015 = ~pi798  & ~n8014;
  assign n8016 = ~n8013 & ~n8015;
  assign n8017 = ~n8009 & n8016;
  assign n8018 = n8009 & ~n8016;
  assign n8019 = ~n8017 & ~n8018;
  assign n8020 = ~n8002 & ~n8019;
  assign n8021 = n8002 & n8019;
  assign n8022 = ~n8020 & ~n8021;
  assign n8023 = pi775  & ~pi776 ;
  assign n8024 = ~pi775  & pi776 ;
  assign n8025 = pi777  & ~n8023;
  assign n8026 = ~n8024 & n8025;
  assign n8027 = ~n8023 & ~n8024;
  assign n8028 = ~pi777  & ~n8027;
  assign n8029 = ~n8026 & ~n8028;
  assign n8030 = pi778  & ~pi779 ;
  assign n8031 = ~pi778  & pi779 ;
  assign n8032 = pi780  & ~n8030;
  assign n8033 = ~n8031 & n8032;
  assign n8034 = ~n8030 & ~n8031;
  assign n8035 = ~pi780  & ~n8034;
  assign n8036 = ~n8033 & ~n8035;
  assign n8037 = ~n8029 & n8036;
  assign n8038 = n8029 & ~n8036;
  assign n8039 = ~n8037 & ~n8038;
  assign n8040 = pi781  & ~pi782 ;
  assign n8041 = ~pi781  & pi782 ;
  assign n8042 = pi783  & ~n8040;
  assign n8043 = ~n8041 & n8042;
  assign n8044 = ~n8040 & ~n8041;
  assign n8045 = ~pi783  & ~n8044;
  assign n8046 = ~n8043 & ~n8045;
  assign n8047 = pi784  & ~pi785 ;
  assign n8048 = ~pi784  & pi785 ;
  assign n8049 = pi786  & ~n8047;
  assign n8050 = ~n8048 & n8049;
  assign n8051 = ~n8047 & ~n8048;
  assign n8052 = ~pi786  & ~n8051;
  assign n8053 = ~n8050 & ~n8052;
  assign n8054 = ~n8046 & n8053;
  assign n8055 = n8046 & ~n8053;
  assign n8056 = ~n8054 & ~n8055;
  assign n8057 = ~n8039 & ~n8056;
  assign n8058 = n8039 & n8056;
  assign n8059 = ~n8057 & ~n8058;
  assign n8060 = n8022 & n8059;
  assign n8061 = ~n8022 & ~n8059;
  assign n8062 = ~n8060 & ~n8061;
  assign n8063 = ~pi769  & pi770 ;
  assign n8064 = pi769  & ~pi770 ;
  assign n8065 = pi771  & ~n8063;
  assign n8066 = ~n8064 & n8065;
  assign n8067 = ~n8063 & ~n8064;
  assign n8068 = ~pi771  & ~n8067;
  assign n8069 = ~n8066 & ~n8068;
  assign n8070 = ~pi772  & pi773 ;
  assign n8071 = pi772  & ~pi773 ;
  assign n8072 = pi774  & ~n8070;
  assign n8073 = ~n8071 & n8072;
  assign n8074 = ~n8070 & ~n8071;
  assign n8075 = ~pi774  & ~n8074;
  assign n8076 = ~n8073 & ~n8075;
  assign n8077 = ~n8069 & n8076;
  assign n8078 = n8069 & ~n8076;
  assign n8079 = ~n8077 & ~n8078;
  assign n8080 = ~pi763  & pi764 ;
  assign n8081 = pi763  & ~pi764 ;
  assign n8082 = pi765  & ~n8080;
  assign n8083 = ~n8081 & n8082;
  assign n8084 = ~n8080 & ~n8081;
  assign n8085 = ~pi765  & ~n8084;
  assign n8086 = ~n8083 & ~n8085;
  assign n8087 = ~pi766  & pi767 ;
  assign n8088 = pi766  & ~pi767 ;
  assign n8089 = pi768  & ~n8087;
  assign n8090 = ~n8088 & n8089;
  assign n8091 = ~n8087 & ~n8088;
  assign n8092 = ~pi768  & ~n8091;
  assign n8093 = ~n8090 & ~n8092;
  assign n8094 = ~n8086 & n8093;
  assign n8095 = n8086 & ~n8093;
  assign n8096 = ~n8094 & ~n8095;
  assign n8097 = ~n8079 & ~n8096;
  assign n8098 = n8079 & n8096;
  assign n8099 = ~n8097 & ~n8098;
  assign n8100 = ~pi757  & pi758 ;
  assign n8101 = pi757  & ~pi758 ;
  assign n8102 = pi759  & ~n8100;
  assign n8103 = ~n8101 & n8102;
  assign n8104 = ~n8100 & ~n8101;
  assign n8105 = ~pi759  & ~n8104;
  assign n8106 = ~n8103 & ~n8105;
  assign n8107 = ~pi760  & pi761 ;
  assign n8108 = pi760  & ~pi761 ;
  assign n8109 = pi762  & ~n8107;
  assign n8110 = ~n8108 & n8109;
  assign n8111 = ~n8107 & ~n8108;
  assign n8112 = ~pi762  & ~n8111;
  assign n8113 = ~n8110 & ~n8112;
  assign n8114 = ~n8106 & n8113;
  assign n8115 = n8106 & ~n8113;
  assign n8116 = ~n8114 & ~n8115;
  assign n8117 = ~pi751  & pi752 ;
  assign n8118 = pi751  & ~pi752 ;
  assign n8119 = pi753  & ~n8117;
  assign n8120 = ~n8118 & n8119;
  assign n8121 = ~n8117 & ~n8118;
  assign n8122 = ~pi753  & ~n8121;
  assign n8123 = ~n8120 & ~n8122;
  assign n8124 = ~pi754  & pi755 ;
  assign n8125 = pi754  & ~pi755 ;
  assign n8126 = pi756  & ~n8124;
  assign n8127 = ~n8125 & n8126;
  assign n8128 = ~n8124 & ~n8125;
  assign n8129 = ~pi756  & ~n8128;
  assign n8130 = ~n8127 & ~n8129;
  assign n8131 = ~n8123 & n8130;
  assign n8132 = n8123 & ~n8130;
  assign n8133 = ~n8131 & ~n8132;
  assign n8134 = ~n8116 & ~n8133;
  assign n8135 = n8116 & n8133;
  assign n8136 = ~n8134 & ~n8135;
  assign n8137 = n8099 & n8136;
  assign n8138 = ~n8099 & ~n8136;
  assign n8139 = ~n8137 & ~n8138;
  assign n8140 = n8062 & ~n8139;
  assign n8141 = ~n8062 & n8139;
  assign n8142 = ~n8140 & ~n8141;
  assign n8143 = ~n7985 & ~n8142;
  assign n8144 = n7985 & n8142;
  assign n8145 = ~n8143 & ~n8144;
  assign n8146 = pi739  & ~pi740 ;
  assign n8147 = ~pi739  & pi740 ;
  assign n8148 = pi741  & ~n8146;
  assign n8149 = ~n8147 & n8148;
  assign n8150 = ~n8146 & ~n8147;
  assign n8151 = ~pi741  & ~n8150;
  assign n8152 = ~n8149 & ~n8151;
  assign n8153 = pi742  & ~pi743 ;
  assign n8154 = ~pi742  & pi743 ;
  assign n8155 = pi744  & ~n8153;
  assign n8156 = ~n8154 & n8155;
  assign n8157 = ~n8153 & ~n8154;
  assign n8158 = ~pi744  & ~n8157;
  assign n8159 = ~n8156 & ~n8158;
  assign n8160 = ~n8152 & n8159;
  assign n8161 = n8152 & ~n8159;
  assign n8162 = ~n8160 & ~n8161;
  assign n8163 = pi745  & ~pi746 ;
  assign n8164 = ~pi745  & pi746 ;
  assign n8165 = pi747  & ~n8163;
  assign n8166 = ~n8164 & n8165;
  assign n8167 = ~n8163 & ~n8164;
  assign n8168 = ~pi747  & ~n8167;
  assign n8169 = ~n8166 & ~n8168;
  assign n8170 = pi748  & ~pi749 ;
  assign n8171 = ~pi748  & pi749 ;
  assign n8172 = pi750  & ~n8170;
  assign n8173 = ~n8171 & n8172;
  assign n8174 = ~n8170 & ~n8171;
  assign n8175 = ~pi750  & ~n8174;
  assign n8176 = ~n8173 & ~n8175;
  assign n8177 = ~n8169 & n8176;
  assign n8178 = n8169 & ~n8176;
  assign n8179 = ~n8177 & ~n8178;
  assign n8180 = ~n8162 & ~n8179;
  assign n8181 = n8162 & n8179;
  assign n8182 = ~n8180 & ~n8181;
  assign n8183 = pi727  & ~pi728 ;
  assign n8184 = ~pi727  & pi728 ;
  assign n8185 = pi729  & ~n8183;
  assign n8186 = ~n8184 & n8185;
  assign n8187 = ~n8183 & ~n8184;
  assign n8188 = ~pi729  & ~n8187;
  assign n8189 = ~n8186 & ~n8188;
  assign n8190 = pi730  & ~pi731 ;
  assign n8191 = ~pi730  & pi731 ;
  assign n8192 = pi732  & ~n8190;
  assign n8193 = ~n8191 & n8192;
  assign n8194 = ~n8190 & ~n8191;
  assign n8195 = ~pi732  & ~n8194;
  assign n8196 = ~n8193 & ~n8195;
  assign n8197 = ~n8189 & n8196;
  assign n8198 = n8189 & ~n8196;
  assign n8199 = ~n8197 & ~n8198;
  assign n8200 = pi733  & ~pi734 ;
  assign n8201 = ~pi733  & pi734 ;
  assign n8202 = pi735  & ~n8200;
  assign n8203 = ~n8201 & n8202;
  assign n8204 = ~n8200 & ~n8201;
  assign n8205 = ~pi735  & ~n8204;
  assign n8206 = ~n8203 & ~n8205;
  assign n8207 = pi736  & ~pi737 ;
  assign n8208 = ~pi736  & pi737 ;
  assign n8209 = pi738  & ~n8207;
  assign n8210 = ~n8208 & n8209;
  assign n8211 = ~n8207 & ~n8208;
  assign n8212 = ~pi738  & ~n8211;
  assign n8213 = ~n8210 & ~n8212;
  assign n8214 = ~n8206 & n8213;
  assign n8215 = n8206 & ~n8213;
  assign n8216 = ~n8214 & ~n8215;
  assign n8217 = ~n8199 & ~n8216;
  assign n8218 = n8199 & n8216;
  assign n8219 = ~n8217 & ~n8218;
  assign n8220 = n8182 & n8219;
  assign n8221 = ~n8182 & ~n8219;
  assign n8222 = ~n8220 & ~n8221;
  assign n8223 = pi715  & ~pi716 ;
  assign n8224 = ~pi715  & pi716 ;
  assign n8225 = pi717  & ~n8223;
  assign n8226 = ~n8224 & n8225;
  assign n8227 = ~n8223 & ~n8224;
  assign n8228 = ~pi717  & ~n8227;
  assign n8229 = ~n8226 & ~n8228;
  assign n8230 = pi718  & ~pi719 ;
  assign n8231 = ~pi718  & pi719 ;
  assign n8232 = pi720  & ~n8230;
  assign n8233 = ~n8231 & n8232;
  assign n8234 = ~n8230 & ~n8231;
  assign n8235 = ~pi720  & ~n8234;
  assign n8236 = ~n8233 & ~n8235;
  assign n8237 = ~n8229 & n8236;
  assign n8238 = n8229 & ~n8236;
  assign n8239 = ~n8237 & ~n8238;
  assign n8240 = pi721  & ~pi722 ;
  assign n8241 = ~pi721  & pi722 ;
  assign n8242 = pi723  & ~n8240;
  assign n8243 = ~n8241 & n8242;
  assign n8244 = ~n8240 & ~n8241;
  assign n8245 = ~pi723  & ~n8244;
  assign n8246 = ~n8243 & ~n8245;
  assign n8247 = pi724  & ~pi725 ;
  assign n8248 = ~pi724  & pi725 ;
  assign n8249 = pi726  & ~n8247;
  assign n8250 = ~n8248 & n8249;
  assign n8251 = ~n8247 & ~n8248;
  assign n8252 = ~pi726  & ~n8251;
  assign n8253 = ~n8250 & ~n8252;
  assign n8254 = ~n8246 & n8253;
  assign n8255 = n8246 & ~n8253;
  assign n8256 = ~n8254 & ~n8255;
  assign n8257 = ~n8239 & ~n8256;
  assign n8258 = n8239 & n8256;
  assign n8259 = ~n8257 & ~n8258;
  assign n8260 = ~pi709  & pi710 ;
  assign n8261 = pi709  & ~pi710 ;
  assign n8262 = pi711  & ~n8260;
  assign n8263 = ~n8261 & n8262;
  assign n8264 = ~n8260 & ~n8261;
  assign n8265 = ~pi711  & ~n8264;
  assign n8266 = ~n8263 & ~n8265;
  assign n8267 = ~pi712  & pi713 ;
  assign n8268 = pi712  & ~pi713 ;
  assign n8269 = pi714  & ~n8267;
  assign n8270 = ~n8268 & n8269;
  assign n8271 = ~n8267 & ~n8268;
  assign n8272 = ~pi714  & ~n8271;
  assign n8273 = ~n8270 & ~n8272;
  assign n8274 = ~n8266 & n8273;
  assign n8275 = n8266 & ~n8273;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = ~pi703  & pi704 ;
  assign n8278 = pi703  & ~pi704 ;
  assign n8279 = pi705  & ~n8277;
  assign n8280 = ~n8278 & n8279;
  assign n8281 = ~n8277 & ~n8278;
  assign n8282 = ~pi705  & ~n8281;
  assign n8283 = ~n8280 & ~n8282;
  assign n8284 = ~pi706  & pi707 ;
  assign n8285 = pi706  & ~pi707 ;
  assign n8286 = pi708  & ~n8284;
  assign n8287 = ~n8285 & n8286;
  assign n8288 = ~n8284 & ~n8285;
  assign n8289 = ~pi708  & ~n8288;
  assign n8290 = ~n8287 & ~n8289;
  assign n8291 = ~n8283 & n8290;
  assign n8292 = n8283 & ~n8290;
  assign n8293 = ~n8291 & ~n8292;
  assign n8294 = ~n8276 & ~n8293;
  assign n8295 = n8276 & n8293;
  assign n8296 = ~n8294 & ~n8295;
  assign n8297 = n8259 & n8296;
  assign n8298 = ~n8259 & ~n8296;
  assign n8299 = ~n8297 & ~n8298;
  assign n8300 = n8222 & ~n8299;
  assign n8301 = ~n8222 & n8299;
  assign n8302 = ~n8300 & ~n8301;
  assign n8303 = ~pi697  & pi698 ;
  assign n8304 = pi697  & ~pi698 ;
  assign n8305 = pi699  & ~n8303;
  assign n8306 = ~n8304 & n8305;
  assign n8307 = ~n8303 & ~n8304;
  assign n8308 = ~pi699  & ~n8307;
  assign n8309 = ~n8306 & ~n8308;
  assign n8310 = ~pi700  & pi701 ;
  assign n8311 = pi700  & ~pi701 ;
  assign n8312 = pi702  & ~n8310;
  assign n8313 = ~n8311 & n8312;
  assign n8314 = ~n8310 & ~n8311;
  assign n8315 = ~pi702  & ~n8314;
  assign n8316 = ~n8313 & ~n8315;
  assign n8317 = ~n8309 & n8316;
  assign n8318 = n8309 & ~n8316;
  assign n8319 = ~n8317 & ~n8318;
  assign n8320 = ~pi691  & pi692 ;
  assign n8321 = pi691  & ~pi692 ;
  assign n8322 = pi693  & ~n8320;
  assign n8323 = ~n8321 & n8322;
  assign n8324 = ~n8320 & ~n8321;
  assign n8325 = ~pi693  & ~n8324;
  assign n8326 = ~n8323 & ~n8325;
  assign n8327 = ~pi694  & pi695 ;
  assign n8328 = pi694  & ~pi695 ;
  assign n8329 = pi696  & ~n8327;
  assign n8330 = ~n8328 & n8329;
  assign n8331 = ~n8327 & ~n8328;
  assign n8332 = ~pi696  & ~n8331;
  assign n8333 = ~n8330 & ~n8332;
  assign n8334 = ~n8326 & n8333;
  assign n8335 = n8326 & ~n8333;
  assign n8336 = ~n8334 & ~n8335;
  assign n8337 = ~n8319 & ~n8336;
  assign n8338 = n8319 & n8336;
  assign n8339 = ~n8337 & ~n8338;
  assign n8340 = ~pi685  & pi686 ;
  assign n8341 = pi685  & ~pi686 ;
  assign n8342 = pi687  & ~n8340;
  assign n8343 = ~n8341 & n8342;
  assign n8344 = ~n8340 & ~n8341;
  assign n8345 = ~pi687  & ~n8344;
  assign n8346 = ~n8343 & ~n8345;
  assign n8347 = ~pi688  & pi689 ;
  assign n8348 = pi688  & ~pi689 ;
  assign n8349 = pi690  & ~n8347;
  assign n8350 = ~n8348 & n8349;
  assign n8351 = ~n8347 & ~n8348;
  assign n8352 = ~pi690  & ~n8351;
  assign n8353 = ~n8350 & ~n8352;
  assign n8354 = ~n8346 & n8353;
  assign n8355 = n8346 & ~n8353;
  assign n8356 = ~n8354 & ~n8355;
  assign n8357 = ~pi679  & pi680 ;
  assign n8358 = pi679  & ~pi680 ;
  assign n8359 = pi681  & ~n8357;
  assign n8360 = ~n8358 & n8359;
  assign n8361 = ~n8357 & ~n8358;
  assign n8362 = ~pi681  & ~n8361;
  assign n8363 = ~n8360 & ~n8362;
  assign n8364 = ~pi682  & pi683 ;
  assign n8365 = pi682  & ~pi683 ;
  assign n8366 = pi684  & ~n8364;
  assign n8367 = ~n8365 & n8366;
  assign n8368 = ~n8364 & ~n8365;
  assign n8369 = ~pi684  & ~n8368;
  assign n8370 = ~n8367 & ~n8369;
  assign n8371 = ~n8363 & n8370;
  assign n8372 = n8363 & ~n8370;
  assign n8373 = ~n8371 & ~n8372;
  assign n8374 = ~n8356 & ~n8373;
  assign n8375 = n8356 & n8373;
  assign n8376 = ~n8374 & ~n8375;
  assign n8377 = n8339 & n8376;
  assign n8378 = ~n8339 & ~n8376;
  assign n8379 = ~n8377 & ~n8378;
  assign n8380 = ~pi673  & pi674 ;
  assign n8381 = pi673  & ~pi674 ;
  assign n8382 = pi675  & ~n8380;
  assign n8383 = ~n8381 & n8382;
  assign n8384 = ~n8380 & ~n8381;
  assign n8385 = ~pi675  & ~n8384;
  assign n8386 = ~n8383 & ~n8385;
  assign n8387 = ~pi676  & pi677 ;
  assign n8388 = pi676  & ~pi677 ;
  assign n8389 = pi678  & ~n8387;
  assign n8390 = ~n8388 & n8389;
  assign n8391 = ~n8387 & ~n8388;
  assign n8392 = ~pi678  & ~n8391;
  assign n8393 = ~n8390 & ~n8392;
  assign n8394 = ~n8386 & n8393;
  assign n8395 = n8386 & ~n8393;
  assign n8396 = ~n8394 & ~n8395;
  assign n8397 = ~pi667  & pi668 ;
  assign n8398 = pi667  & ~pi668 ;
  assign n8399 = pi669  & ~n8397;
  assign n8400 = ~n8398 & n8399;
  assign n8401 = ~n8397 & ~n8398;
  assign n8402 = ~pi669  & ~n8401;
  assign n8403 = ~n8400 & ~n8402;
  assign n8404 = ~pi670  & pi671 ;
  assign n8405 = pi670  & ~pi671 ;
  assign n8406 = pi672  & ~n8404;
  assign n8407 = ~n8405 & n8406;
  assign n8408 = ~n8404 & ~n8405;
  assign n8409 = ~pi672  & ~n8408;
  assign n8410 = ~n8407 & ~n8409;
  assign n8411 = ~n8403 & n8410;
  assign n8412 = n8403 & ~n8410;
  assign n8413 = ~n8411 & ~n8412;
  assign n8414 = ~n8396 & ~n8413;
  assign n8415 = n8396 & n8413;
  assign n8416 = ~n8414 & ~n8415;
  assign n8417 = ~pi661  & pi662 ;
  assign n8418 = pi661  & ~pi662 ;
  assign n8419 = pi663  & ~n8417;
  assign n8420 = ~n8418 & n8419;
  assign n8421 = ~n8417 & ~n8418;
  assign n8422 = ~pi663  & ~n8421;
  assign n8423 = ~n8420 & ~n8422;
  assign n8424 = ~pi664  & pi665 ;
  assign n8425 = pi664  & ~pi665 ;
  assign n8426 = pi666  & ~n8424;
  assign n8427 = ~n8425 & n8426;
  assign n8428 = ~n8424 & ~n8425;
  assign n8429 = ~pi666  & ~n8428;
  assign n8430 = ~n8427 & ~n8429;
  assign n8431 = ~n8423 & n8430;
  assign n8432 = n8423 & ~n8430;
  assign n8433 = ~n8431 & ~n8432;
  assign n8434 = ~pi655  & pi656 ;
  assign n8435 = pi655  & ~pi656 ;
  assign n8436 = pi657  & ~n8434;
  assign n8437 = ~n8435 & n8436;
  assign n8438 = ~n8434 & ~n8435;
  assign n8439 = ~pi657  & ~n8438;
  assign n8440 = ~n8437 & ~n8439;
  assign n8441 = ~pi658  & pi659 ;
  assign n8442 = pi658  & ~pi659 ;
  assign n8443 = pi660  & ~n8441;
  assign n8444 = ~n8442 & n8443;
  assign n8445 = ~n8441 & ~n8442;
  assign n8446 = ~pi660  & ~n8445;
  assign n8447 = ~n8444 & ~n8446;
  assign n8448 = ~n8440 & n8447;
  assign n8449 = n8440 & ~n8447;
  assign n8450 = ~n8448 & ~n8449;
  assign n8451 = ~n8433 & ~n8450;
  assign n8452 = n8433 & n8450;
  assign n8453 = ~n8451 & ~n8452;
  assign n8454 = n8416 & n8453;
  assign n8455 = ~n8416 & ~n8453;
  assign n8456 = ~n8454 & ~n8455;
  assign n8457 = n8379 & ~n8456;
  assign n8458 = ~n8379 & n8456;
  assign n8459 = ~n8457 & ~n8458;
  assign n8460 = ~n8302 & ~n8459;
  assign n8461 = n8302 & n8459;
  assign n8462 = ~n8460 & ~n8461;
  assign n8463 = n8145 & n8462;
  assign n8464 = ~n8145 & ~n8462;
  assign n8465 = ~n8463 & ~n8464;
  assign n8466 = n7828 & ~n8465;
  assign n8467 = ~n7828 & n8465;
  assign n8468 = ~n8466 & ~n8467;
  assign n8469 = ~n7162 & ~n7164;
  assign n8470 = n7162 & n7164;
  assign n8471 = ~n8469 & ~n8470;
  assign n8472 = ~n8468 & ~n8471;
  assign n8473 = n8468 & n8471;
  assign n8474 = ~n8472 & ~n8473;
  assign n8475 = pi1000  & n8474;
  assign n8476 = ~n7170 & ~n7171;
  assign n8477 = ~n7175 & n8476;
  assign n8478 = n7175 & ~n8476;
  assign n8479 = ~n8477 & ~n8478;
  assign n8480 = ~n8472 & n8479;
  assign n8481 = n8472 & ~n8479;
  assign n8482 = ~n8480 & ~n8481;
  assign n8483 = n7828 & n8465;
  assign n8484 = n7905 & n7982;
  assign n8485 = pi844  & pi845 ;
  assign n8486 = pi846  & ~n7857;
  assign n8487 = ~n8485 & ~n8486;
  assign n8488 = pi841  & pi842 ;
  assign n8489 = pi843  & ~n7850;
  assign n8490 = ~n8488 & ~n8489;
  assign n8491 = ~n8487 & ~n8490;
  assign n8492 = ~n7862 & n8491;
  assign n8493 = ~n7852 & ~n7859;
  assign n8494 = n8487 & n8490;
  assign n8495 = ~n8491 & ~n8494;
  assign n8496 = n8493 & n8495;
  assign n8497 = ~n8493 & ~n8495;
  assign n8498 = ~n8492 & ~n8496;
  assign n8499 = ~n8497 & n8498;
  assign n8500 = pi838  & pi839 ;
  assign n8501 = pi840  & ~n7840;
  assign n8502 = ~n8500 & ~n8501;
  assign n8503 = pi835  & pi836 ;
  assign n8504 = pi837  & ~n7833;
  assign n8505 = ~n8503 & ~n8504;
  assign n8506 = n8502 & ~n8505;
  assign n8507 = ~n8502 & n8505;
  assign n8508 = ~n8506 & ~n8507;
  assign n8509 = n7863 & ~n8508;
  assign n8510 = ~n7835 & ~n7842;
  assign n8511 = n8508 & n8510;
  assign n8512 = ~n8508 & ~n8510;
  assign n8513 = ~n8511 & ~n8512;
  assign n8514 = ~n7863 & n8513;
  assign n8515 = ~n8509 & ~n8514;
  assign n8516 = n8499 & ~n8515;
  assign n8517 = ~n8499 & n8515;
  assign n8518 = ~n8516 & ~n8517;
  assign n8519 = n7903 & ~n8518;
  assign n8520 = ~n7903 & n8518;
  assign n8521 = ~n8519 & ~n8520;
  assign n8522 = pi832  & pi833 ;
  assign n8523 = pi834  & ~n7894;
  assign n8524 = ~n8522 & ~n8523;
  assign n8525 = pi829  & pi830 ;
  assign n8526 = pi831  & ~n7887;
  assign n8527 = ~n8525 & ~n8526;
  assign n8528 = ~n8524 & ~n8527;
  assign n8529 = ~n7899 & n8528;
  assign n8530 = ~n7889 & ~n7896;
  assign n8531 = n8524 & n8527;
  assign n8532 = ~n8528 & ~n8531;
  assign n8533 = n8530 & n8532;
  assign n8534 = ~n8530 & ~n8532;
  assign n8535 = ~n8529 & ~n8533;
  assign n8536 = ~n8534 & n8535;
  assign n8537 = ~n7900 & ~n8536;
  assign n8538 = n7900 & n8536;
  assign n8539 = ~n8537 & ~n8538;
  assign n8540 = ~n7872 & ~n7879;
  assign n8541 = pi826  & pi827 ;
  assign n8542 = pi828  & ~n7877;
  assign n8543 = ~n8541 & ~n8542;
  assign n8544 = pi823  & pi824 ;
  assign n8545 = pi825  & ~n7870;
  assign n8546 = ~n8544 & ~n8545;
  assign n8547 = n8543 & ~n8546;
  assign n8548 = ~n8543 & n8546;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = n8540 & n8549;
  assign n8551 = ~n8540 & ~n8549;
  assign n8552 = ~n8550 & ~n8551;
  assign n8553 = n8539 & ~n8552;
  assign n8554 = ~n8539 & n8552;
  assign n8555 = ~n8553 & ~n8554;
  assign n8556 = n8521 & ~n8555;
  assign n8557 = ~n8521 & n8555;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = n8484 & ~n8558;
  assign n8560 = ~n8484 & n8558;
  assign n8561 = ~n8559 & ~n8560;
  assign n8562 = pi820  & pi821 ;
  assign n8563 = pi822  & ~n7934;
  assign n8564 = ~n8562 & ~n8563;
  assign n8565 = pi817  & pi818 ;
  assign n8566 = pi819  & ~n7927;
  assign n8567 = ~n8565 & ~n8566;
  assign n8568 = ~n8564 & ~n8567;
  assign n8569 = ~n7939 & n8568;
  assign n8570 = ~n7929 & ~n7936;
  assign n8571 = n8564 & n8567;
  assign n8572 = ~n8568 & ~n8571;
  assign n8573 = n8570 & n8572;
  assign n8574 = ~n8570 & ~n8572;
  assign n8575 = ~n8569 & ~n8573;
  assign n8576 = ~n8574 & n8575;
  assign n8577 = pi814  & pi815 ;
  assign n8578 = pi816  & ~n7917;
  assign n8579 = ~n8577 & ~n8578;
  assign n8580 = pi811  & pi812 ;
  assign n8581 = pi813  & ~n7910;
  assign n8582 = ~n8580 & ~n8581;
  assign n8583 = n8579 & ~n8582;
  assign n8584 = ~n8579 & n8582;
  assign n8585 = ~n8583 & ~n8584;
  assign n8586 = n7940 & ~n8585;
  assign n8587 = ~n7912 & ~n7919;
  assign n8588 = n8585 & n8587;
  assign n8589 = ~n8585 & ~n8587;
  assign n8590 = ~n8588 & ~n8589;
  assign n8591 = ~n7940 & n8590;
  assign n8592 = ~n8586 & ~n8591;
  assign n8593 = n8576 & ~n8592;
  assign n8594 = ~n8576 & n8592;
  assign n8595 = ~n8593 & ~n8594;
  assign n8596 = n7980 & ~n8595;
  assign n8597 = ~n7980 & n8595;
  assign n8598 = ~n8596 & ~n8597;
  assign n8599 = pi808  & pi809 ;
  assign n8600 = pi810  & ~n7954;
  assign n8601 = ~n8599 & ~n8600;
  assign n8602 = pi805  & pi806 ;
  assign n8603 = pi807  & ~n7947;
  assign n8604 = ~n8602 & ~n8603;
  assign n8605 = ~n8601 & ~n8604;
  assign n8606 = ~n7959 & n8605;
  assign n8607 = ~n7949 & ~n7956;
  assign n8608 = n8601 & n8604;
  assign n8609 = ~n8605 & ~n8608;
  assign n8610 = n8607 & n8609;
  assign n8611 = ~n8607 & ~n8609;
  assign n8612 = ~n8606 & ~n8610;
  assign n8613 = ~n8611 & n8612;
  assign n8614 = ~n7977 & ~n8613;
  assign n8615 = n7977 & n8613;
  assign n8616 = ~n8614 & ~n8615;
  assign n8617 = pi802  & pi803 ;
  assign n8618 = pi804  & ~n7971;
  assign n8619 = ~n8617 & ~n8618;
  assign n8620 = pi799  & pi800 ;
  assign n8621 = pi801  & ~n7964;
  assign n8622 = ~n8620 & ~n8621;
  assign n8623 = ~n8619 & n8622;
  assign n8624 = n8619 & ~n8622;
  assign n8625 = ~n8623 & ~n8624;
  assign n8626 = ~n7966 & ~n7973;
  assign n8627 = n8625 & n8626;
  assign n8628 = ~n8625 & ~n8626;
  assign n8629 = ~n8627 & ~n8628;
  assign n8630 = n8616 & ~n8629;
  assign n8631 = ~n8616 & n8629;
  assign n8632 = ~n8630 & ~n8631;
  assign n8633 = n8598 & ~n8632;
  assign n8634 = ~n8598 & n8632;
  assign n8635 = ~n8633 & ~n8634;
  assign n8636 = n8561 & n8635;
  assign n8637 = ~n8561 & ~n8635;
  assign n8638 = ~n8636 & ~n8637;
  assign n8639 = n8143 & ~n8638;
  assign n8640 = ~n8143 & n8638;
  assign n8641 = ~n8639 & ~n8640;
  assign n8642 = n8062 & n8139;
  assign n8643 = pi796  & pi797 ;
  assign n8644 = pi798  & ~n8014;
  assign n8645 = ~n8643 & ~n8644;
  assign n8646 = pi793  & pi794 ;
  assign n8647 = pi795  & ~n8007;
  assign n8648 = ~n8646 & ~n8647;
  assign n8649 = ~n8645 & ~n8648;
  assign n8650 = ~n8019 & n8649;
  assign n8651 = ~n8009 & ~n8016;
  assign n8652 = n8645 & n8648;
  assign n8653 = ~n8649 & ~n8652;
  assign n8654 = n8651 & n8653;
  assign n8655 = ~n8651 & ~n8653;
  assign n8656 = ~n8650 & ~n8654;
  assign n8657 = ~n8655 & n8656;
  assign n8658 = pi790  & pi791 ;
  assign n8659 = pi792  & ~n7997;
  assign n8660 = ~n8658 & ~n8659;
  assign n8661 = pi787  & pi788 ;
  assign n8662 = pi789  & ~n7990;
  assign n8663 = ~n8661 & ~n8662;
  assign n8664 = n8660 & ~n8663;
  assign n8665 = ~n8660 & n8663;
  assign n8666 = ~n8664 & ~n8665;
  assign n8667 = n8020 & ~n8666;
  assign n8668 = ~n7992 & ~n7999;
  assign n8669 = n8666 & n8668;
  assign n8670 = ~n8666 & ~n8668;
  assign n8671 = ~n8669 & ~n8670;
  assign n8672 = ~n8020 & n8671;
  assign n8673 = ~n8667 & ~n8672;
  assign n8674 = n8657 & ~n8673;
  assign n8675 = ~n8657 & n8673;
  assign n8676 = ~n8674 & ~n8675;
  assign n8677 = n8060 & ~n8676;
  assign n8678 = ~n8060 & n8676;
  assign n8679 = ~n8677 & ~n8678;
  assign n8680 = pi784  & pi785 ;
  assign n8681 = pi786  & ~n8051;
  assign n8682 = ~n8680 & ~n8681;
  assign n8683 = pi781  & pi782 ;
  assign n8684 = pi783  & ~n8044;
  assign n8685 = ~n8683 & ~n8684;
  assign n8686 = ~n8682 & ~n8685;
  assign n8687 = ~n8056 & n8686;
  assign n8688 = ~n8046 & ~n8053;
  assign n8689 = n8682 & n8685;
  assign n8690 = ~n8686 & ~n8689;
  assign n8691 = n8688 & n8690;
  assign n8692 = ~n8688 & ~n8690;
  assign n8693 = ~n8687 & ~n8691;
  assign n8694 = ~n8692 & n8693;
  assign n8695 = ~n8057 & ~n8694;
  assign n8696 = n8057 & n8694;
  assign n8697 = ~n8695 & ~n8696;
  assign n8698 = ~n8029 & ~n8036;
  assign n8699 = pi778  & pi779 ;
  assign n8700 = pi780  & ~n8034;
  assign n8701 = ~n8699 & ~n8700;
  assign n8702 = pi775  & pi776 ;
  assign n8703 = pi777  & ~n8027;
  assign n8704 = ~n8702 & ~n8703;
  assign n8705 = n8701 & ~n8704;
  assign n8706 = ~n8701 & n8704;
  assign n8707 = ~n8705 & ~n8706;
  assign n8708 = n8698 & n8707;
  assign n8709 = ~n8698 & ~n8707;
  assign n8710 = ~n8708 & ~n8709;
  assign n8711 = n8697 & ~n8710;
  assign n8712 = ~n8697 & n8710;
  assign n8713 = ~n8711 & ~n8712;
  assign n8714 = n8679 & ~n8713;
  assign n8715 = ~n8679 & n8713;
  assign n8716 = ~n8714 & ~n8715;
  assign n8717 = n8642 & ~n8716;
  assign n8718 = ~n8642 & n8716;
  assign n8719 = ~n8717 & ~n8718;
  assign n8720 = pi766  & pi767 ;
  assign n8721 = pi768  & ~n8091;
  assign n8722 = ~n8720 & ~n8721;
  assign n8723 = pi763  & pi764 ;
  assign n8724 = pi765  & ~n8084;
  assign n8725 = ~n8723 & ~n8724;
  assign n8726 = ~n8722 & ~n8725;
  assign n8727 = ~n8096 & n8726;
  assign n8728 = ~n8086 & ~n8093;
  assign n8729 = n8722 & n8725;
  assign n8730 = ~n8726 & ~n8729;
  assign n8731 = n8728 & n8730;
  assign n8732 = ~n8728 & ~n8730;
  assign n8733 = ~n8727 & ~n8731;
  assign n8734 = ~n8732 & n8733;
  assign n8735 = ~n8069 & ~n8076;
  assign n8736 = pi772  & pi773 ;
  assign n8737 = pi774  & ~n8074;
  assign n8738 = ~n8736 & ~n8737;
  assign n8739 = pi769  & pi770 ;
  assign n8740 = pi771  & ~n8067;
  assign n8741 = ~n8739 & ~n8740;
  assign n8742 = n8738 & ~n8741;
  assign n8743 = ~n8738 & n8741;
  assign n8744 = ~n8742 & ~n8743;
  assign n8745 = n8735 & n8744;
  assign n8746 = ~n8735 & ~n8744;
  assign n8747 = ~n8097 & ~n8745;
  assign n8748 = ~n8746 & n8747;
  assign n8749 = n8097 & ~n8744;
  assign n8750 = ~n8748 & ~n8749;
  assign n8751 = n8734 & n8750;
  assign n8752 = ~n8734 & ~n8750;
  assign n8753 = ~n8751 & ~n8752;
  assign n8754 = n8137 & n8753;
  assign n8755 = ~n8137 & ~n8753;
  assign n8756 = ~n8754 & ~n8755;
  assign n8757 = pi760  & pi761 ;
  assign n8758 = pi762  & ~n8111;
  assign n8759 = ~n8757 & ~n8758;
  assign n8760 = pi757  & pi758 ;
  assign n8761 = pi759  & ~n8104;
  assign n8762 = ~n8760 & ~n8761;
  assign n8763 = ~n8759 & ~n8762;
  assign n8764 = ~n8116 & n8763;
  assign n8765 = ~n8106 & ~n8113;
  assign n8766 = n8759 & n8762;
  assign n8767 = ~n8763 & ~n8766;
  assign n8768 = n8765 & n8767;
  assign n8769 = ~n8765 & ~n8767;
  assign n8770 = ~n8764 & ~n8768;
  assign n8771 = ~n8769 & n8770;
  assign n8772 = ~n8134 & ~n8771;
  assign n8773 = n8134 & n8771;
  assign n8774 = ~n8772 & ~n8773;
  assign n8775 = pi754  & pi755 ;
  assign n8776 = pi756  & ~n8128;
  assign n8777 = ~n8775 & ~n8776;
  assign n8778 = pi751  & pi752 ;
  assign n8779 = pi753  & ~n8121;
  assign n8780 = ~n8778 & ~n8779;
  assign n8781 = ~n8777 & n8780;
  assign n8782 = n8777 & ~n8780;
  assign n8783 = ~n8781 & ~n8782;
  assign n8784 = ~n8123 & ~n8130;
  assign n8785 = n8783 & n8784;
  assign n8786 = ~n8783 & ~n8784;
  assign n8787 = ~n8785 & ~n8786;
  assign n8788 = n8774 & ~n8787;
  assign n8789 = ~n8774 & n8787;
  assign n8790 = ~n8788 & ~n8789;
  assign n8791 = n8756 & ~n8790;
  assign n8792 = ~n8756 & n8790;
  assign n8793 = ~n8791 & ~n8792;
  assign n8794 = n8719 & n8793;
  assign n8795 = ~n8719 & ~n8793;
  assign n8796 = ~n8794 & ~n8795;
  assign n8797 = n8641 & n8796;
  assign n8798 = ~n8641 & ~n8796;
  assign n8799 = ~n8797 & ~n8798;
  assign n8800 = n8463 & ~n8799;
  assign n8801 = ~n8463 & n8799;
  assign n8802 = ~n8800 & ~n8801;
  assign n8803 = n8222 & n8299;
  assign n8804 = pi748  & pi749 ;
  assign n8805 = pi750  & ~n8174;
  assign n8806 = ~n8804 & ~n8805;
  assign n8807 = pi745  & pi746 ;
  assign n8808 = pi747  & ~n8167;
  assign n8809 = ~n8807 & ~n8808;
  assign n8810 = ~n8806 & ~n8809;
  assign n8811 = ~n8179 & n8810;
  assign n8812 = ~n8169 & ~n8176;
  assign n8813 = n8806 & n8809;
  assign n8814 = ~n8810 & ~n8813;
  assign n8815 = n8812 & n8814;
  assign n8816 = ~n8812 & ~n8814;
  assign n8817 = ~n8811 & ~n8815;
  assign n8818 = ~n8816 & n8817;
  assign n8819 = pi742  & pi743 ;
  assign n8820 = pi744  & ~n8157;
  assign n8821 = ~n8819 & ~n8820;
  assign n8822 = pi739  & pi740 ;
  assign n8823 = pi741  & ~n8150;
  assign n8824 = ~n8822 & ~n8823;
  assign n8825 = n8821 & ~n8824;
  assign n8826 = ~n8821 & n8824;
  assign n8827 = ~n8825 & ~n8826;
  assign n8828 = n8180 & ~n8827;
  assign n8829 = ~n8152 & ~n8159;
  assign n8830 = n8827 & n8829;
  assign n8831 = ~n8827 & ~n8829;
  assign n8832 = ~n8830 & ~n8831;
  assign n8833 = ~n8180 & n8832;
  assign n8834 = ~n8828 & ~n8833;
  assign n8835 = n8818 & ~n8834;
  assign n8836 = ~n8818 & n8834;
  assign n8837 = ~n8835 & ~n8836;
  assign n8838 = n8220 & ~n8837;
  assign n8839 = ~n8220 & n8837;
  assign n8840 = ~n8838 & ~n8839;
  assign n8841 = pi736  & pi737 ;
  assign n8842 = pi738  & ~n8211;
  assign n8843 = ~n8841 & ~n8842;
  assign n8844 = pi733  & pi734 ;
  assign n8845 = pi735  & ~n8204;
  assign n8846 = ~n8844 & ~n8845;
  assign n8847 = ~n8843 & ~n8846;
  assign n8848 = ~n8216 & n8847;
  assign n8849 = ~n8206 & ~n8213;
  assign n8850 = n8843 & n8846;
  assign n8851 = ~n8847 & ~n8850;
  assign n8852 = n8849 & n8851;
  assign n8853 = ~n8849 & ~n8851;
  assign n8854 = ~n8848 & ~n8852;
  assign n8855 = ~n8853 & n8854;
  assign n8856 = ~n8217 & ~n8855;
  assign n8857 = n8217 & n8855;
  assign n8858 = ~n8856 & ~n8857;
  assign n8859 = ~n8189 & ~n8196;
  assign n8860 = pi730  & pi731 ;
  assign n8861 = pi732  & ~n8194;
  assign n8862 = ~n8860 & ~n8861;
  assign n8863 = pi727  & pi728 ;
  assign n8864 = pi729  & ~n8187;
  assign n8865 = ~n8863 & ~n8864;
  assign n8866 = n8862 & ~n8865;
  assign n8867 = ~n8862 & n8865;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = n8859 & n8868;
  assign n8870 = ~n8859 & ~n8868;
  assign n8871 = ~n8869 & ~n8870;
  assign n8872 = n8858 & ~n8871;
  assign n8873 = ~n8858 & n8871;
  assign n8874 = ~n8872 & ~n8873;
  assign n8875 = n8840 & ~n8874;
  assign n8876 = ~n8840 & n8874;
  assign n8877 = ~n8875 & ~n8876;
  assign n8878 = n8803 & ~n8877;
  assign n8879 = ~n8803 & n8877;
  assign n8880 = ~n8878 & ~n8879;
  assign n8881 = pi724  & pi725 ;
  assign n8882 = pi726  & ~n8251;
  assign n8883 = ~n8881 & ~n8882;
  assign n8884 = pi721  & pi722 ;
  assign n8885 = pi723  & ~n8244;
  assign n8886 = ~n8884 & ~n8885;
  assign n8887 = ~n8883 & ~n8886;
  assign n8888 = ~n8256 & n8887;
  assign n8889 = ~n8246 & ~n8253;
  assign n8890 = n8883 & n8886;
  assign n8891 = ~n8887 & ~n8890;
  assign n8892 = n8889 & n8891;
  assign n8893 = ~n8889 & ~n8891;
  assign n8894 = ~n8888 & ~n8892;
  assign n8895 = ~n8893 & n8894;
  assign n8896 = pi718  & pi719 ;
  assign n8897 = pi720  & ~n8234;
  assign n8898 = ~n8896 & ~n8897;
  assign n8899 = pi715  & pi716 ;
  assign n8900 = pi717  & ~n8227;
  assign n8901 = ~n8899 & ~n8900;
  assign n8902 = n8898 & ~n8901;
  assign n8903 = ~n8898 & n8901;
  assign n8904 = ~n8902 & ~n8903;
  assign n8905 = n8257 & ~n8904;
  assign n8906 = ~n8229 & ~n8236;
  assign n8907 = n8904 & n8906;
  assign n8908 = ~n8904 & ~n8906;
  assign n8909 = ~n8907 & ~n8908;
  assign n8910 = ~n8257 & n8909;
  assign n8911 = ~n8905 & ~n8910;
  assign n8912 = n8895 & ~n8911;
  assign n8913 = ~n8895 & n8911;
  assign n8914 = ~n8912 & ~n8913;
  assign n8915 = n8297 & ~n8914;
  assign n8916 = ~n8297 & n8914;
  assign n8917 = ~n8915 & ~n8916;
  assign n8918 = pi712  & pi713 ;
  assign n8919 = pi714  & ~n8271;
  assign n8920 = ~n8918 & ~n8919;
  assign n8921 = pi709  & pi710 ;
  assign n8922 = pi711  & ~n8264;
  assign n8923 = ~n8921 & ~n8922;
  assign n8924 = ~n8920 & ~n8923;
  assign n8925 = ~n8276 & n8924;
  assign n8926 = ~n8266 & ~n8273;
  assign n8927 = n8920 & n8923;
  assign n8928 = ~n8924 & ~n8927;
  assign n8929 = n8926 & n8928;
  assign n8930 = ~n8926 & ~n8928;
  assign n8931 = ~n8925 & ~n8929;
  assign n8932 = ~n8930 & n8931;
  assign n8933 = ~n8294 & ~n8932;
  assign n8934 = n8294 & n8932;
  assign n8935 = ~n8933 & ~n8934;
  assign n8936 = pi706  & pi707 ;
  assign n8937 = pi708  & ~n8288;
  assign n8938 = ~n8936 & ~n8937;
  assign n8939 = pi703  & pi704 ;
  assign n8940 = pi705  & ~n8281;
  assign n8941 = ~n8939 & ~n8940;
  assign n8942 = ~n8938 & n8941;
  assign n8943 = n8938 & ~n8941;
  assign n8944 = ~n8942 & ~n8943;
  assign n8945 = ~n8283 & ~n8290;
  assign n8946 = n8944 & n8945;
  assign n8947 = ~n8944 & ~n8945;
  assign n8948 = ~n8946 & ~n8947;
  assign n8949 = n8935 & ~n8948;
  assign n8950 = ~n8935 & n8948;
  assign n8951 = ~n8949 & ~n8950;
  assign n8952 = n8917 & ~n8951;
  assign n8953 = ~n8917 & n8951;
  assign n8954 = ~n8952 & ~n8953;
  assign n8955 = n8880 & n8954;
  assign n8956 = ~n8880 & ~n8954;
  assign n8957 = ~n8955 & ~n8956;
  assign n8958 = n8460 & ~n8957;
  assign n8959 = ~n8460 & n8957;
  assign n8960 = ~n8958 & ~n8959;
  assign n8961 = n8379 & n8456;
  assign n8962 = pi694  & pi695 ;
  assign n8963 = pi696  & ~n8331;
  assign n8964 = ~n8962 & ~n8963;
  assign n8965 = pi691  & pi692 ;
  assign n8966 = pi693  & ~n8324;
  assign n8967 = ~n8965 & ~n8966;
  assign n8968 = ~n8964 & ~n8967;
  assign n8969 = ~n8336 & n8968;
  assign n8970 = ~n8326 & ~n8333;
  assign n8971 = n8964 & n8967;
  assign n8972 = ~n8968 & ~n8971;
  assign n8973 = n8970 & n8972;
  assign n8974 = ~n8970 & ~n8972;
  assign n8975 = ~n8969 & ~n8973;
  assign n8976 = ~n8974 & n8975;
  assign n8977 = ~n8309 & ~n8316;
  assign n8978 = pi700  & pi701 ;
  assign n8979 = pi702  & ~n8314;
  assign n8980 = ~n8978 & ~n8979;
  assign n8981 = pi697  & pi698 ;
  assign n8982 = pi699  & ~n8307;
  assign n8983 = ~n8981 & ~n8982;
  assign n8984 = n8980 & ~n8983;
  assign n8985 = ~n8980 & n8983;
  assign n8986 = ~n8984 & ~n8985;
  assign n8987 = n8977 & n8986;
  assign n8988 = ~n8977 & ~n8986;
  assign n8989 = ~n8337 & ~n8987;
  assign n8990 = ~n8988 & n8989;
  assign n8991 = n8337 & ~n8986;
  assign n8992 = ~n8990 & ~n8991;
  assign n8993 = n8976 & n8992;
  assign n8994 = ~n8976 & ~n8992;
  assign n8995 = ~n8993 & ~n8994;
  assign n8996 = n8377 & n8995;
  assign n8997 = ~n8377 & ~n8995;
  assign n8998 = ~n8996 & ~n8997;
  assign n8999 = pi688  & pi689 ;
  assign n9000 = pi690  & ~n8351;
  assign n9001 = ~n8999 & ~n9000;
  assign n9002 = pi685  & pi686 ;
  assign n9003 = pi687  & ~n8344;
  assign n9004 = ~n9002 & ~n9003;
  assign n9005 = ~n9001 & ~n9004;
  assign n9006 = ~n8356 & n9005;
  assign n9007 = ~n8346 & ~n8353;
  assign n9008 = n9001 & n9004;
  assign n9009 = ~n9005 & ~n9008;
  assign n9010 = n9007 & n9009;
  assign n9011 = ~n9007 & ~n9009;
  assign n9012 = ~n9006 & ~n9010;
  assign n9013 = ~n9011 & n9012;
  assign n9014 = ~n8374 & ~n9013;
  assign n9015 = n8374 & n9013;
  assign n9016 = ~n9014 & ~n9015;
  assign n9017 = pi682  & pi683 ;
  assign n9018 = pi684  & ~n8368;
  assign n9019 = ~n9017 & ~n9018;
  assign n9020 = pi679  & pi680 ;
  assign n9021 = pi681  & ~n8361;
  assign n9022 = ~n9020 & ~n9021;
  assign n9023 = ~n9019 & n9022;
  assign n9024 = n9019 & ~n9022;
  assign n9025 = ~n9023 & ~n9024;
  assign n9026 = ~n8363 & ~n8370;
  assign n9027 = n9025 & n9026;
  assign n9028 = ~n9025 & ~n9026;
  assign n9029 = ~n9027 & ~n9028;
  assign n9030 = n9016 & ~n9029;
  assign n9031 = ~n9016 & n9029;
  assign n9032 = ~n9030 & ~n9031;
  assign n9033 = n8998 & ~n9032;
  assign n9034 = ~n8998 & n9032;
  assign n9035 = ~n9033 & ~n9034;
  assign n9036 = n8961 & ~n9035;
  assign n9037 = ~n8961 & n9035;
  assign n9038 = ~n9036 & ~n9037;
  assign n9039 = pi670  & pi671 ;
  assign n9040 = pi672  & ~n8408;
  assign n9041 = ~n9039 & ~n9040;
  assign n9042 = pi667  & pi668 ;
  assign n9043 = pi669  & ~n8401;
  assign n9044 = ~n9042 & ~n9043;
  assign n9045 = ~n9041 & ~n9044;
  assign n9046 = ~n8413 & n9045;
  assign n9047 = ~n8403 & ~n8410;
  assign n9048 = n9041 & n9044;
  assign n9049 = ~n9045 & ~n9048;
  assign n9050 = n9047 & n9049;
  assign n9051 = ~n9047 & ~n9049;
  assign n9052 = ~n9046 & ~n9050;
  assign n9053 = ~n9051 & n9052;
  assign n9054 = ~n8386 & ~n8393;
  assign n9055 = pi676  & pi677 ;
  assign n9056 = pi678  & ~n8391;
  assign n9057 = ~n9055 & ~n9056;
  assign n9058 = pi673  & pi674 ;
  assign n9059 = pi675  & ~n8384;
  assign n9060 = ~n9058 & ~n9059;
  assign n9061 = n9057 & ~n9060;
  assign n9062 = ~n9057 & n9060;
  assign n9063 = ~n9061 & ~n9062;
  assign n9064 = n9054 & n9063;
  assign n9065 = ~n9054 & ~n9063;
  assign n9066 = ~n8414 & ~n9064;
  assign n9067 = ~n9065 & n9066;
  assign n9068 = n8414 & ~n9063;
  assign n9069 = ~n9067 & ~n9068;
  assign n9070 = n9053 & n9069;
  assign n9071 = ~n9053 & ~n9069;
  assign n9072 = ~n9070 & ~n9071;
  assign n9073 = n8454 & n9072;
  assign n9074 = ~n8454 & ~n9072;
  assign n9075 = ~n9073 & ~n9074;
  assign n9076 = pi664  & pi665 ;
  assign n9077 = pi666  & ~n8428;
  assign n9078 = ~n9076 & ~n9077;
  assign n9079 = pi661  & pi662 ;
  assign n9080 = pi663  & ~n8421;
  assign n9081 = ~n9079 & ~n9080;
  assign n9082 = ~n9078 & ~n9081;
  assign n9083 = ~n8433 & n9082;
  assign n9084 = ~n8423 & ~n8430;
  assign n9085 = n9078 & n9081;
  assign n9086 = ~n9082 & ~n9085;
  assign n9087 = n9084 & n9086;
  assign n9088 = ~n9084 & ~n9086;
  assign n9089 = ~n9083 & ~n9087;
  assign n9090 = ~n9088 & n9089;
  assign n9091 = ~n8451 & ~n9090;
  assign n9092 = n8451 & n9090;
  assign n9093 = ~n9091 & ~n9092;
  assign n9094 = pi658  & pi659 ;
  assign n9095 = pi660  & ~n8445;
  assign n9096 = ~n9094 & ~n9095;
  assign n9097 = pi655  & pi656 ;
  assign n9098 = pi657  & ~n8438;
  assign n9099 = ~n9097 & ~n9098;
  assign n9100 = ~n9096 & n9099;
  assign n9101 = n9096 & ~n9099;
  assign n9102 = ~n9100 & ~n9101;
  assign n9103 = ~n8440 & ~n8447;
  assign n9104 = n9102 & n9103;
  assign n9105 = ~n9102 & ~n9103;
  assign n9106 = ~n9104 & ~n9105;
  assign n9107 = n9093 & ~n9106;
  assign n9108 = ~n9093 & n9106;
  assign n9109 = ~n9107 & ~n9108;
  assign n9110 = n9075 & ~n9109;
  assign n9111 = ~n9075 & n9109;
  assign n9112 = ~n9110 & ~n9111;
  assign n9113 = n9038 & n9112;
  assign n9114 = ~n9038 & ~n9112;
  assign n9115 = ~n9113 & ~n9114;
  assign n9116 = n8960 & n9115;
  assign n9117 = ~n8960 & ~n9115;
  assign n9118 = ~n9116 & ~n9117;
  assign n9119 = n8802 & ~n9118;
  assign n9120 = ~n8802 & n9118;
  assign n9121 = ~n9119 & ~n9120;
  assign n9122 = n8483 & n9121;
  assign n9123 = ~n8483 & ~n9121;
  assign n9124 = ~n9122 & ~n9123;
  assign n9125 = n7585 & n7662;
  assign n9126 = pi646  & pi647 ;
  assign n9127 = pi648  & ~n7537;
  assign n9128 = ~n9126 & ~n9127;
  assign n9129 = pi643  & pi644 ;
  assign n9130 = pi645  & ~n7530;
  assign n9131 = ~n9129 & ~n9130;
  assign n9132 = ~n9128 & ~n9131;
  assign n9133 = ~n7542 & n9132;
  assign n9134 = ~n7532 & ~n7539;
  assign n9135 = n9128 & n9131;
  assign n9136 = ~n9132 & ~n9135;
  assign n9137 = n9134 & n9136;
  assign n9138 = ~n9134 & ~n9136;
  assign n9139 = ~n9133 & ~n9137;
  assign n9140 = ~n9138 & n9139;
  assign n9141 = ~n7515 & ~n7522;
  assign n9142 = pi652  & pi653 ;
  assign n9143 = pi654  & ~n7520;
  assign n9144 = ~n9142 & ~n9143;
  assign n9145 = pi649  & pi650 ;
  assign n9146 = pi651  & ~n7513;
  assign n9147 = ~n9145 & ~n9146;
  assign n9148 = n9144 & ~n9147;
  assign n9149 = ~n9144 & n9147;
  assign n9150 = ~n9148 & ~n9149;
  assign n9151 = n9141 & n9150;
  assign n9152 = ~n9141 & ~n9150;
  assign n9153 = ~n7543 & ~n9151;
  assign n9154 = ~n9152 & n9153;
  assign n9155 = n7543 & ~n9150;
  assign n9156 = ~n9154 & ~n9155;
  assign n9157 = n9140 & n9156;
  assign n9158 = ~n9140 & ~n9156;
  assign n9159 = ~n9157 & ~n9158;
  assign n9160 = n7583 & n9159;
  assign n9161 = ~n7583 & ~n9159;
  assign n9162 = ~n9160 & ~n9161;
  assign n9163 = pi640  & pi641 ;
  assign n9164 = pi642  & ~n7557;
  assign n9165 = ~n9163 & ~n9164;
  assign n9166 = pi637  & pi638 ;
  assign n9167 = pi639  & ~n7550;
  assign n9168 = ~n9166 & ~n9167;
  assign n9169 = ~n9165 & ~n9168;
  assign n9170 = ~n7562 & n9169;
  assign n9171 = ~n7552 & ~n7559;
  assign n9172 = n9165 & n9168;
  assign n9173 = ~n9169 & ~n9172;
  assign n9174 = n9171 & n9173;
  assign n9175 = ~n9171 & ~n9173;
  assign n9176 = ~n9170 & ~n9174;
  assign n9177 = ~n9175 & n9176;
  assign n9178 = ~n7580 & ~n9177;
  assign n9179 = n7580 & n9177;
  assign n9180 = ~n9178 & ~n9179;
  assign n9181 = pi634  & pi635 ;
  assign n9182 = pi636  & ~n7574;
  assign n9183 = ~n9181 & ~n9182;
  assign n9184 = pi631  & pi632 ;
  assign n9185 = pi633  & ~n7567;
  assign n9186 = ~n9184 & ~n9185;
  assign n9187 = ~n9183 & n9186;
  assign n9188 = n9183 & ~n9186;
  assign n9189 = ~n9187 & ~n9188;
  assign n9190 = ~n7569 & ~n7576;
  assign n9191 = n9189 & n9190;
  assign n9192 = ~n9189 & ~n9190;
  assign n9193 = ~n9191 & ~n9192;
  assign n9194 = n9180 & ~n9193;
  assign n9195 = ~n9180 & n9193;
  assign n9196 = ~n9194 & ~n9195;
  assign n9197 = n9162 & ~n9196;
  assign n9198 = ~n9162 & n9196;
  assign n9199 = ~n9197 & ~n9198;
  assign n9200 = n9125 & ~n9199;
  assign n9201 = ~n9125 & n9199;
  assign n9202 = ~n9200 & ~n9201;
  assign n9203 = pi622  & pi623 ;
  assign n9204 = pi624  & ~n7614;
  assign n9205 = ~n9203 & ~n9204;
  assign n9206 = pi619  & pi620 ;
  assign n9207 = pi621  & ~n7607;
  assign n9208 = ~n9206 & ~n9207;
  assign n9209 = ~n9205 & ~n9208;
  assign n9210 = ~n7619 & n9209;
  assign n9211 = ~n7609 & ~n7616;
  assign n9212 = n9205 & n9208;
  assign n9213 = ~n9209 & ~n9212;
  assign n9214 = n9211 & n9213;
  assign n9215 = ~n9211 & ~n9213;
  assign n9216 = ~n9210 & ~n9214;
  assign n9217 = ~n9215 & n9216;
  assign n9218 = ~n7592 & ~n7599;
  assign n9219 = pi628  & pi629 ;
  assign n9220 = pi630  & ~n7597;
  assign n9221 = ~n9219 & ~n9220;
  assign n9222 = pi625  & pi626 ;
  assign n9223 = pi627  & ~n7590;
  assign n9224 = ~n9222 & ~n9223;
  assign n9225 = n9221 & ~n9224;
  assign n9226 = ~n9221 & n9224;
  assign n9227 = ~n9225 & ~n9226;
  assign n9228 = n9218 & n9227;
  assign n9229 = ~n9218 & ~n9227;
  assign n9230 = ~n7620 & ~n9228;
  assign n9231 = ~n9229 & n9230;
  assign n9232 = n7620 & ~n9227;
  assign n9233 = ~n9231 & ~n9232;
  assign n9234 = n9217 & n9233;
  assign n9235 = ~n9217 & ~n9233;
  assign n9236 = ~n9234 & ~n9235;
  assign n9237 = n7660 & n9236;
  assign n9238 = ~n7660 & ~n9236;
  assign n9239 = ~n9237 & ~n9238;
  assign n9240 = pi616  & pi617 ;
  assign n9241 = pi618  & ~n7634;
  assign n9242 = ~n9240 & ~n9241;
  assign n9243 = pi613  & pi614 ;
  assign n9244 = pi615  & ~n7627;
  assign n9245 = ~n9243 & ~n9244;
  assign n9246 = ~n9242 & ~n9245;
  assign n9247 = ~n7639 & n9246;
  assign n9248 = ~n7629 & ~n7636;
  assign n9249 = n9242 & n9245;
  assign n9250 = ~n9246 & ~n9249;
  assign n9251 = n9248 & n9250;
  assign n9252 = ~n9248 & ~n9250;
  assign n9253 = ~n9247 & ~n9251;
  assign n9254 = ~n9252 & n9253;
  assign n9255 = ~n7657 & ~n9254;
  assign n9256 = n7657 & n9254;
  assign n9257 = ~n9255 & ~n9256;
  assign n9258 = pi610  & pi611 ;
  assign n9259 = pi612  & ~n7651;
  assign n9260 = ~n9258 & ~n9259;
  assign n9261 = pi607  & pi608 ;
  assign n9262 = pi609  & ~n7644;
  assign n9263 = ~n9261 & ~n9262;
  assign n9264 = ~n9260 & n9263;
  assign n9265 = n9260 & ~n9263;
  assign n9266 = ~n9264 & ~n9265;
  assign n9267 = ~n7646 & ~n7653;
  assign n9268 = n9266 & n9267;
  assign n9269 = ~n9266 & ~n9267;
  assign n9270 = ~n9268 & ~n9269;
  assign n9271 = n9257 & ~n9270;
  assign n9272 = ~n9257 & n9270;
  assign n9273 = ~n9271 & ~n9272;
  assign n9274 = n9239 & ~n9273;
  assign n9275 = ~n9239 & n9273;
  assign n9276 = ~n9274 & ~n9275;
  assign n9277 = n9202 & n9276;
  assign n9278 = ~n9202 & ~n9276;
  assign n9279 = ~n9277 & ~n9278;
  assign n9280 = n7823 & ~n9279;
  assign n9281 = ~n7823 & n9279;
  assign n9282 = ~n9280 & ~n9281;
  assign n9283 = n7742 & n7819;
  assign n9284 = pi598  & pi599 ;
  assign n9285 = pi600  & ~n7694;
  assign n9286 = ~n9284 & ~n9285;
  assign n9287 = pi595  & pi596 ;
  assign n9288 = pi597  & ~n7687;
  assign n9289 = ~n9287 & ~n9288;
  assign n9290 = ~n9286 & ~n9289;
  assign n9291 = ~n7699 & n9290;
  assign n9292 = ~n7689 & ~n7696;
  assign n9293 = n9286 & n9289;
  assign n9294 = ~n9290 & ~n9293;
  assign n9295 = n9292 & n9294;
  assign n9296 = ~n9292 & ~n9294;
  assign n9297 = ~n9291 & ~n9295;
  assign n9298 = ~n9296 & n9297;
  assign n9299 = ~n7672 & ~n7679;
  assign n9300 = pi604  & pi605 ;
  assign n9301 = pi606  & ~n7677;
  assign n9302 = ~n9300 & ~n9301;
  assign n9303 = pi601  & pi602 ;
  assign n9304 = pi603  & ~n7670;
  assign n9305 = ~n9303 & ~n9304;
  assign n9306 = n9302 & ~n9305;
  assign n9307 = ~n9302 & n9305;
  assign n9308 = ~n9306 & ~n9307;
  assign n9309 = n9299 & n9308;
  assign n9310 = ~n9299 & ~n9308;
  assign n9311 = ~n7700 & ~n9309;
  assign n9312 = ~n9310 & n9311;
  assign n9313 = n7700 & ~n9308;
  assign n9314 = ~n9312 & ~n9313;
  assign n9315 = n9298 & n9314;
  assign n9316 = ~n9298 & ~n9314;
  assign n9317 = ~n9315 & ~n9316;
  assign n9318 = n7740 & n9317;
  assign n9319 = ~n7740 & ~n9317;
  assign n9320 = ~n9318 & ~n9319;
  assign n9321 = pi592  & pi593 ;
  assign n9322 = pi594  & ~n7714;
  assign n9323 = ~n9321 & ~n9322;
  assign n9324 = pi589  & pi590 ;
  assign n9325 = pi591  & ~n7707;
  assign n9326 = ~n9324 & ~n9325;
  assign n9327 = ~n9323 & ~n9326;
  assign n9328 = ~n7719 & n9327;
  assign n9329 = ~n7709 & ~n7716;
  assign n9330 = n9323 & n9326;
  assign n9331 = ~n9327 & ~n9330;
  assign n9332 = n9329 & n9331;
  assign n9333 = ~n9329 & ~n9331;
  assign n9334 = ~n9328 & ~n9332;
  assign n9335 = ~n9333 & n9334;
  assign n9336 = ~n7737 & ~n9335;
  assign n9337 = n7737 & n9335;
  assign n9338 = ~n9336 & ~n9337;
  assign n9339 = pi586  & pi587 ;
  assign n9340 = pi588  & ~n7731;
  assign n9341 = ~n9339 & ~n9340;
  assign n9342 = pi583  & pi584 ;
  assign n9343 = pi585  & ~n7724;
  assign n9344 = ~n9342 & ~n9343;
  assign n9345 = ~n9341 & n9344;
  assign n9346 = n9341 & ~n9344;
  assign n9347 = ~n9345 & ~n9346;
  assign n9348 = ~n7726 & ~n7733;
  assign n9349 = n9347 & n9348;
  assign n9350 = ~n9347 & ~n9348;
  assign n9351 = ~n9349 & ~n9350;
  assign n9352 = n9338 & ~n9351;
  assign n9353 = ~n9338 & n9351;
  assign n9354 = ~n9352 & ~n9353;
  assign n9355 = n9320 & ~n9354;
  assign n9356 = ~n9320 & n9354;
  assign n9357 = ~n9355 & ~n9356;
  assign n9358 = n9283 & ~n9357;
  assign n9359 = ~n9283 & n9357;
  assign n9360 = ~n9358 & ~n9359;
  assign n9361 = pi574  & pi575 ;
  assign n9362 = pi576  & ~n7771;
  assign n9363 = ~n9361 & ~n9362;
  assign n9364 = pi571  & pi572 ;
  assign n9365 = pi573  & ~n7764;
  assign n9366 = ~n9364 & ~n9365;
  assign n9367 = ~n9363 & ~n9366;
  assign n9368 = ~n7776 & n9367;
  assign n9369 = ~n7766 & ~n7773;
  assign n9370 = n9363 & n9366;
  assign n9371 = ~n9367 & ~n9370;
  assign n9372 = n9369 & n9371;
  assign n9373 = ~n9369 & ~n9371;
  assign n9374 = ~n9368 & ~n9372;
  assign n9375 = ~n9373 & n9374;
  assign n9376 = ~n7749 & ~n7756;
  assign n9377 = pi580  & pi581 ;
  assign n9378 = pi582  & ~n7754;
  assign n9379 = ~n9377 & ~n9378;
  assign n9380 = pi577  & pi578 ;
  assign n9381 = pi579  & ~n7747;
  assign n9382 = ~n9380 & ~n9381;
  assign n9383 = n9379 & ~n9382;
  assign n9384 = ~n9379 & n9382;
  assign n9385 = ~n9383 & ~n9384;
  assign n9386 = n9376 & n9385;
  assign n9387 = ~n9376 & ~n9385;
  assign n9388 = ~n7777 & ~n9386;
  assign n9389 = ~n9387 & n9388;
  assign n9390 = n7777 & ~n9385;
  assign n9391 = ~n9389 & ~n9390;
  assign n9392 = n9375 & n9391;
  assign n9393 = ~n9375 & ~n9391;
  assign n9394 = ~n9392 & ~n9393;
  assign n9395 = n7817 & n9394;
  assign n9396 = ~n7817 & ~n9394;
  assign n9397 = ~n9395 & ~n9396;
  assign n9398 = pi568  & pi569 ;
  assign n9399 = pi570  & ~n7791;
  assign n9400 = ~n9398 & ~n9399;
  assign n9401 = pi565  & pi566 ;
  assign n9402 = pi567  & ~n7784;
  assign n9403 = ~n9401 & ~n9402;
  assign n9404 = ~n9400 & ~n9403;
  assign n9405 = ~n7796 & n9404;
  assign n9406 = ~n7786 & ~n7793;
  assign n9407 = n9400 & n9403;
  assign n9408 = ~n9404 & ~n9407;
  assign n9409 = n9406 & n9408;
  assign n9410 = ~n9406 & ~n9408;
  assign n9411 = ~n9405 & ~n9409;
  assign n9412 = ~n9410 & n9411;
  assign n9413 = ~n7814 & ~n9412;
  assign n9414 = n7814 & n9412;
  assign n9415 = ~n9413 & ~n9414;
  assign n9416 = pi562  & pi563 ;
  assign n9417 = pi564  & ~n7808;
  assign n9418 = ~n9416 & ~n9417;
  assign n9419 = pi559  & pi560 ;
  assign n9420 = pi561  & ~n7801;
  assign n9421 = ~n9419 & ~n9420;
  assign n9422 = ~n9418 & n9421;
  assign n9423 = n9418 & ~n9421;
  assign n9424 = ~n9422 & ~n9423;
  assign n9425 = ~n7803 & ~n7810;
  assign n9426 = n9424 & n9425;
  assign n9427 = ~n9424 & ~n9425;
  assign n9428 = ~n9426 & ~n9427;
  assign n9429 = n9415 & ~n9428;
  assign n9430 = ~n9415 & n9428;
  assign n9431 = ~n9429 & ~n9430;
  assign n9432 = n9397 & ~n9431;
  assign n9433 = ~n9397 & n9431;
  assign n9434 = ~n9432 & ~n9433;
  assign n9435 = n9360 & n9434;
  assign n9436 = ~n9360 & ~n9434;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = n9282 & n9437;
  assign n9439 = ~n9282 & ~n9437;
  assign n9440 = ~n9438 & ~n9439;
  assign n9441 = n7826 & ~n9440;
  assign n9442 = ~n7826 & n9440;
  assign n9443 = ~n9441 & ~n9442;
  assign n9444 = n7425 & n7502;
  assign n9445 = pi550  & pi551 ;
  assign n9446 = pi552  & ~n7377;
  assign n9447 = ~n9445 & ~n9446;
  assign n9448 = pi547  & pi548 ;
  assign n9449 = pi549  & ~n7370;
  assign n9450 = ~n9448 & ~n9449;
  assign n9451 = ~n9447 & ~n9450;
  assign n9452 = ~n7382 & n9451;
  assign n9453 = ~n7372 & ~n7379;
  assign n9454 = n9447 & n9450;
  assign n9455 = ~n9451 & ~n9454;
  assign n9456 = n9453 & n9455;
  assign n9457 = ~n9453 & ~n9455;
  assign n9458 = ~n9452 & ~n9456;
  assign n9459 = ~n9457 & n9458;
  assign n9460 = ~n7355 & ~n7362;
  assign n9461 = pi556  & pi557 ;
  assign n9462 = pi558  & ~n7360;
  assign n9463 = ~n9461 & ~n9462;
  assign n9464 = pi553  & pi554 ;
  assign n9465 = pi555  & ~n7353;
  assign n9466 = ~n9464 & ~n9465;
  assign n9467 = n9463 & ~n9466;
  assign n9468 = ~n9463 & n9466;
  assign n9469 = ~n9467 & ~n9468;
  assign n9470 = n9460 & n9469;
  assign n9471 = ~n9460 & ~n9469;
  assign n9472 = ~n7383 & ~n9470;
  assign n9473 = ~n9471 & n9472;
  assign n9474 = n7383 & ~n9469;
  assign n9475 = ~n9473 & ~n9474;
  assign n9476 = n9459 & n9475;
  assign n9477 = ~n9459 & ~n9475;
  assign n9478 = ~n9476 & ~n9477;
  assign n9479 = n7423 & n9478;
  assign n9480 = ~n7423 & ~n9478;
  assign n9481 = ~n9479 & ~n9480;
  assign n9482 = pi544  & pi545 ;
  assign n9483 = pi546  & ~n7397;
  assign n9484 = ~n9482 & ~n9483;
  assign n9485 = pi541  & pi542 ;
  assign n9486 = pi543  & ~n7390;
  assign n9487 = ~n9485 & ~n9486;
  assign n9488 = ~n9484 & ~n9487;
  assign n9489 = ~n7402 & n9488;
  assign n9490 = ~n7392 & ~n7399;
  assign n9491 = n9484 & n9487;
  assign n9492 = ~n9488 & ~n9491;
  assign n9493 = n9490 & n9492;
  assign n9494 = ~n9490 & ~n9492;
  assign n9495 = ~n9489 & ~n9493;
  assign n9496 = ~n9494 & n9495;
  assign n9497 = ~n7420 & ~n9496;
  assign n9498 = n7420 & n9496;
  assign n9499 = ~n9497 & ~n9498;
  assign n9500 = pi538  & pi539 ;
  assign n9501 = pi540  & ~n7414;
  assign n9502 = ~n9500 & ~n9501;
  assign n9503 = pi535  & pi536 ;
  assign n9504 = pi537  & ~n7407;
  assign n9505 = ~n9503 & ~n9504;
  assign n9506 = ~n9502 & n9505;
  assign n9507 = n9502 & ~n9505;
  assign n9508 = ~n9506 & ~n9507;
  assign n9509 = ~n7409 & ~n7416;
  assign n9510 = n9508 & n9509;
  assign n9511 = ~n9508 & ~n9509;
  assign n9512 = ~n9510 & ~n9511;
  assign n9513 = n9499 & ~n9512;
  assign n9514 = ~n9499 & n9512;
  assign n9515 = ~n9513 & ~n9514;
  assign n9516 = n9481 & ~n9515;
  assign n9517 = ~n9481 & n9515;
  assign n9518 = ~n9516 & ~n9517;
  assign n9519 = n9444 & ~n9518;
  assign n9520 = ~n9444 & n9518;
  assign n9521 = ~n9519 & ~n9520;
  assign n9522 = pi526  & pi527 ;
  assign n9523 = pi528  & ~n7454;
  assign n9524 = ~n9522 & ~n9523;
  assign n9525 = pi523  & pi524 ;
  assign n9526 = pi525  & ~n7447;
  assign n9527 = ~n9525 & ~n9526;
  assign n9528 = ~n9524 & ~n9527;
  assign n9529 = ~n7459 & n9528;
  assign n9530 = ~n7449 & ~n7456;
  assign n9531 = n9524 & n9527;
  assign n9532 = ~n9528 & ~n9531;
  assign n9533 = n9530 & n9532;
  assign n9534 = ~n9530 & ~n9532;
  assign n9535 = ~n9529 & ~n9533;
  assign n9536 = ~n9534 & n9535;
  assign n9537 = ~n7432 & ~n7439;
  assign n9538 = pi532  & pi533 ;
  assign n9539 = pi534  & ~n7437;
  assign n9540 = ~n9538 & ~n9539;
  assign n9541 = pi529  & pi530 ;
  assign n9542 = pi531  & ~n7430;
  assign n9543 = ~n9541 & ~n9542;
  assign n9544 = n9540 & ~n9543;
  assign n9545 = ~n9540 & n9543;
  assign n9546 = ~n9544 & ~n9545;
  assign n9547 = n9537 & n9546;
  assign n9548 = ~n9537 & ~n9546;
  assign n9549 = ~n7460 & ~n9547;
  assign n9550 = ~n9548 & n9549;
  assign n9551 = n7460 & ~n9546;
  assign n9552 = ~n9550 & ~n9551;
  assign n9553 = n9536 & n9552;
  assign n9554 = ~n9536 & ~n9552;
  assign n9555 = ~n9553 & ~n9554;
  assign n9556 = n7500 & n9555;
  assign n9557 = ~n7500 & ~n9555;
  assign n9558 = ~n9556 & ~n9557;
  assign n9559 = pi520  & pi521 ;
  assign n9560 = pi522  & ~n7474;
  assign n9561 = ~n9559 & ~n9560;
  assign n9562 = pi517  & pi518 ;
  assign n9563 = pi519  & ~n7467;
  assign n9564 = ~n9562 & ~n9563;
  assign n9565 = ~n9561 & ~n9564;
  assign n9566 = ~n7479 & n9565;
  assign n9567 = ~n7469 & ~n7476;
  assign n9568 = n9561 & n9564;
  assign n9569 = ~n9565 & ~n9568;
  assign n9570 = n9567 & n9569;
  assign n9571 = ~n9567 & ~n9569;
  assign n9572 = ~n9566 & ~n9570;
  assign n9573 = ~n9571 & n9572;
  assign n9574 = ~n7497 & ~n9573;
  assign n9575 = n7497 & n9573;
  assign n9576 = ~n9574 & ~n9575;
  assign n9577 = pi514  & pi515 ;
  assign n9578 = pi516  & ~n7491;
  assign n9579 = ~n9577 & ~n9578;
  assign n9580 = pi511  & pi512 ;
  assign n9581 = pi513  & ~n7484;
  assign n9582 = ~n9580 & ~n9581;
  assign n9583 = ~n9579 & n9582;
  assign n9584 = n9579 & ~n9582;
  assign n9585 = ~n9583 & ~n9584;
  assign n9586 = ~n7486 & ~n7493;
  assign n9587 = n9585 & n9586;
  assign n9588 = ~n9585 & ~n9586;
  assign n9589 = ~n9587 & ~n9588;
  assign n9590 = n9576 & ~n9589;
  assign n9591 = ~n9576 & n9589;
  assign n9592 = ~n9590 & ~n9591;
  assign n9593 = n9558 & ~n9592;
  assign n9594 = ~n9558 & n9592;
  assign n9595 = ~n9593 & ~n9594;
  assign n9596 = n9521 & n9595;
  assign n9597 = ~n9521 & ~n9595;
  assign n9598 = ~n9596 & ~n9597;
  assign n9599 = n7506 & ~n9598;
  assign n9600 = ~n7506 & n9598;
  assign n9601 = ~n9599 & ~n9600;
  assign n9602 = n7268 & n7345;
  assign n9603 = pi502  & pi503 ;
  assign n9604 = pi504  & ~n7297;
  assign n9605 = ~n9603 & ~n9604;
  assign n9606 = pi499  & pi500 ;
  assign n9607 = pi501  & ~n7290;
  assign n9608 = ~n9606 & ~n9607;
  assign n9609 = ~n9605 & ~n9608;
  assign n9610 = ~n7302 & n9609;
  assign n9611 = ~n7292 & ~n7299;
  assign n9612 = n9605 & n9608;
  assign n9613 = ~n9609 & ~n9612;
  assign n9614 = n9611 & n9613;
  assign n9615 = ~n9611 & ~n9613;
  assign n9616 = ~n9610 & ~n9614;
  assign n9617 = ~n9615 & n9616;
  assign n9618 = ~n7275 & ~n7282;
  assign n9619 = pi508  & pi509 ;
  assign n9620 = pi510  & ~n7280;
  assign n9621 = ~n9619 & ~n9620;
  assign n9622 = pi505  & pi506 ;
  assign n9623 = pi507  & ~n7273;
  assign n9624 = ~n9622 & ~n9623;
  assign n9625 = n9621 & ~n9624;
  assign n9626 = ~n9621 & n9624;
  assign n9627 = ~n9625 & ~n9626;
  assign n9628 = n9618 & n9627;
  assign n9629 = ~n9618 & ~n9627;
  assign n9630 = ~n7303 & ~n9628;
  assign n9631 = ~n9629 & n9630;
  assign n9632 = n7303 & ~n9627;
  assign n9633 = ~n9631 & ~n9632;
  assign n9634 = n9617 & n9633;
  assign n9635 = ~n9617 & ~n9633;
  assign n9636 = ~n9634 & ~n9635;
  assign n9637 = n7343 & n9636;
  assign n9638 = ~n7343 & ~n9636;
  assign n9639 = ~n9637 & ~n9638;
  assign n9640 = pi496  & pi497 ;
  assign n9641 = pi498  & ~n7317;
  assign n9642 = ~n9640 & ~n9641;
  assign n9643 = pi493  & pi494 ;
  assign n9644 = pi495  & ~n7310;
  assign n9645 = ~n9643 & ~n9644;
  assign n9646 = ~n9642 & ~n9645;
  assign n9647 = ~n7322 & n9646;
  assign n9648 = ~n7312 & ~n7319;
  assign n9649 = n9642 & n9645;
  assign n9650 = ~n9646 & ~n9649;
  assign n9651 = n9648 & n9650;
  assign n9652 = ~n9648 & ~n9650;
  assign n9653 = ~n9647 & ~n9651;
  assign n9654 = ~n9652 & n9653;
  assign n9655 = ~n7340 & ~n9654;
  assign n9656 = n7340 & n9654;
  assign n9657 = ~n9655 & ~n9656;
  assign n9658 = pi490  & pi491 ;
  assign n9659 = pi492  & ~n7334;
  assign n9660 = ~n9658 & ~n9659;
  assign n9661 = pi487  & pi488 ;
  assign n9662 = pi489  & ~n7327;
  assign n9663 = ~n9661 & ~n9662;
  assign n9664 = ~n9660 & n9663;
  assign n9665 = n9660 & ~n9663;
  assign n9666 = ~n9664 & ~n9665;
  assign n9667 = ~n7329 & ~n7336;
  assign n9668 = n9666 & n9667;
  assign n9669 = ~n9666 & ~n9667;
  assign n9670 = ~n9668 & ~n9669;
  assign n9671 = n9657 & ~n9670;
  assign n9672 = ~n9657 & n9670;
  assign n9673 = ~n9671 & ~n9672;
  assign n9674 = n9639 & ~n9673;
  assign n9675 = ~n9639 & n9673;
  assign n9676 = ~n9674 & ~n9675;
  assign n9677 = n9602 & ~n9676;
  assign n9678 = ~n9602 & n9676;
  assign n9679 = ~n9677 & ~n9678;
  assign n9680 = pi478  & pi479 ;
  assign n9681 = pi480  & ~n7257;
  assign n9682 = ~n9680 & ~n9681;
  assign n9683 = pi475  & pi476 ;
  assign n9684 = pi477  & ~n7250;
  assign n9685 = ~n9683 & ~n9684;
  assign n9686 = ~n9682 & ~n9685;
  assign n9687 = ~n7262 & n9686;
  assign n9688 = ~n7252 & ~n7259;
  assign n9689 = n9682 & n9685;
  assign n9690 = ~n9686 & ~n9689;
  assign n9691 = n9688 & n9690;
  assign n9692 = ~n9688 & ~n9690;
  assign n9693 = ~n9687 & ~n9691;
  assign n9694 = ~n9692 & n9693;
  assign n9695 = ~n7235 & ~n7242;
  assign n9696 = pi484  & pi485 ;
  assign n9697 = pi486  & ~n7240;
  assign n9698 = ~n9696 & ~n9697;
  assign n9699 = pi481  & pi482 ;
  assign n9700 = pi483  & ~n7233;
  assign n9701 = ~n9699 & ~n9700;
  assign n9702 = n9698 & ~n9701;
  assign n9703 = ~n9698 & n9701;
  assign n9704 = ~n9702 & ~n9703;
  assign n9705 = n9695 & n9704;
  assign n9706 = ~n9695 & ~n9704;
  assign n9707 = ~n7263 & ~n9705;
  assign n9708 = ~n9706 & n9707;
  assign n9709 = n7263 & ~n9704;
  assign n9710 = ~n9708 & ~n9709;
  assign n9711 = n9694 & n9710;
  assign n9712 = ~n9694 & ~n9710;
  assign n9713 = ~n9711 & ~n9712;
  assign n9714 = n7266 & n9713;
  assign n9715 = ~n7266 & ~n9713;
  assign n9716 = ~n9714 & ~n9715;
  assign n9717 = pi472  & pi473 ;
  assign n9718 = pi474  & ~n7220;
  assign n9719 = ~n9717 & ~n9718;
  assign n9720 = pi469  & pi470 ;
  assign n9721 = pi471  & ~n7213;
  assign n9722 = ~n9720 & ~n9721;
  assign n9723 = ~n9719 & ~n9722;
  assign n9724 = ~n7225 & n9723;
  assign n9725 = ~n7215 & ~n7222;
  assign n9726 = n9719 & n9722;
  assign n9727 = ~n9723 & ~n9726;
  assign n9728 = n9725 & n9727;
  assign n9729 = ~n9725 & ~n9727;
  assign n9730 = ~n9724 & ~n9728;
  assign n9731 = ~n9729 & n9730;
  assign n9732 = pi466  & pi467 ;
  assign n9733 = pi468  & ~n7196;
  assign n9734 = ~n9732 & ~n9733;
  assign n9735 = pi463  & pi464 ;
  assign n9736 = pi465  & ~n7203;
  assign n9737 = ~n9735 & ~n9736;
  assign n9738 = ~n7198 & ~n7205;
  assign n9739 = ~n9734 & n9738;
  assign n9740 = n9734 & ~n9738;
  assign n9741 = ~n9739 & ~n9740;
  assign n9742 = ~n9737 & ~n9741;
  assign n9743 = ~n9734 & n9742;
  assign n9744 = n7226 & ~n9743;
  assign n9745 = ~n9731 & ~n9744;
  assign n9746 = n9731 & n9744;
  assign n9747 = ~n9745 & ~n9746;
  assign n9748 = n9737 & n9741;
  assign n9749 = ~n9742 & ~n9748;
  assign n9750 = n9747 & ~n9749;
  assign n9751 = ~n9747 & n9749;
  assign n9752 = ~n9750 & ~n9751;
  assign n9753 = n9716 & ~n9752;
  assign n9754 = ~n9716 & n9752;
  assign n9755 = ~n9753 & ~n9754;
  assign n9756 = n9679 & n9755;
  assign n9757 = ~n9679 & ~n9755;
  assign n9758 = ~n9756 & ~n9757;
  assign n9759 = n9601 & n9758;
  assign n9760 = ~n9601 & ~n9758;
  assign n9761 = ~n9759 & ~n9760;
  assign n9762 = n9443 & ~n9761;
  assign n9763 = ~n9443 & n9761;
  assign n9764 = ~n9762 & ~n9763;
  assign n9765 = n9124 & ~n9764;
  assign n9766 = ~n9124 & n9764;
  assign n9767 = ~n9765 & ~n9766;
  assign n9768 = n8482 & ~n9767;
  assign n9769 = ~n8482 & n9767;
  assign n9770 = ~n9768 & ~n9769;
  assign n9771 = n8475 & n9770;
  assign n9772 = ~n7158 & ~n7159;
  assign n9773 = ~n7177 & n9772;
  assign n9774 = n7177 & ~n9772;
  assign n9775 = ~n9773 & ~n9774;
  assign n9776 = ~n9746 & n9749;
  assign n9777 = ~n9745 & ~n9776;
  assign n9778 = n9725 & ~n9726;
  assign n9779 = ~n9723 & ~n9778;
  assign n9780 = n9777 & ~n9779;
  assign n9781 = ~n9777 & n9779;
  assign n9782 = ~n9780 & ~n9781;
  assign n9783 = n9737 & ~n9739;
  assign n9784 = ~n9740 & ~n9783;
  assign n9785 = ~n9782 & n9784;
  assign n9786 = n9782 & ~n9784;
  assign n9787 = ~n9785 & ~n9786;
  assign n9788 = n9694 & ~n9708;
  assign n9789 = ~n9709 & ~n9788;
  assign n9790 = n9695 & ~n9698;
  assign n9791 = n9701 & ~n9790;
  assign n9792 = ~n9695 & n9698;
  assign n9793 = ~n9791 & ~n9792;
  assign n9794 = ~n9789 & n9793;
  assign n9795 = n9789 & ~n9793;
  assign n9796 = ~n9794 & ~n9795;
  assign n9797 = n9688 & ~n9689;
  assign n9798 = ~n9686 & ~n9797;
  assign n9799 = n9796 & ~n9798;
  assign n9800 = ~n9796 & n9798;
  assign n9801 = ~n9799 & ~n9800;
  assign n9802 = n9787 & ~n9801;
  assign n9803 = ~n9787 & n9801;
  assign n9804 = ~n9802 & ~n9803;
  assign n9805 = ~n9715 & n9752;
  assign n9806 = ~n9714 & ~n9805;
  assign n9807 = n9804 & ~n9806;
  assign n9808 = ~n9804 & n9806;
  assign n9809 = ~n9807 & ~n9808;
  assign n9810 = ~n9655 & ~n9670;
  assign n9811 = ~n9656 & ~n9810;
  assign n9812 = n9648 & ~n9649;
  assign n9813 = ~n9646 & ~n9812;
  assign n9814 = ~n9811 & ~n9813;
  assign n9815 = n9811 & n9813;
  assign n9816 = ~n9814 & ~n9815;
  assign n9817 = ~n9660 & n9667;
  assign n9818 = n9663 & ~n9817;
  assign n9819 = n9660 & ~n9667;
  assign n9820 = ~n9818 & ~n9819;
  assign n9821 = ~n9816 & n9820;
  assign n9822 = n9816 & ~n9820;
  assign n9823 = ~n9821 & ~n9822;
  assign n9824 = n9617 & ~n9631;
  assign n9825 = ~n9632 & ~n9824;
  assign n9826 = n9618 & ~n9621;
  assign n9827 = n9624 & ~n9826;
  assign n9828 = ~n9618 & n9621;
  assign n9829 = ~n9827 & ~n9828;
  assign n9830 = ~n9825 & n9829;
  assign n9831 = n9825 & ~n9829;
  assign n9832 = ~n9830 & ~n9831;
  assign n9833 = n9611 & ~n9612;
  assign n9834 = ~n9609 & ~n9833;
  assign n9835 = n9832 & ~n9834;
  assign n9836 = ~n9832 & n9834;
  assign n9837 = ~n9835 & ~n9836;
  assign n9838 = n9823 & ~n9837;
  assign n9839 = ~n9823 & n9837;
  assign n9840 = ~n9838 & ~n9839;
  assign n9841 = ~n9638 & n9673;
  assign n9842 = ~n9637 & ~n9841;
  assign n9843 = n9840 & ~n9842;
  assign n9844 = ~n9840 & n9842;
  assign n9845 = ~n9843 & ~n9844;
  assign n9846 = ~n9809 & ~n9845;
  assign n9847 = n9809 & n9845;
  assign n9848 = ~n9846 & ~n9847;
  assign n9849 = ~n9678 & ~n9755;
  assign n9850 = ~n9677 & ~n9849;
  assign n9851 = n9848 & ~n9850;
  assign n9852 = ~n9848 & n9850;
  assign n9853 = ~n9851 & ~n9852;
  assign n9854 = ~n9574 & ~n9589;
  assign n9855 = ~n9575 & ~n9854;
  assign n9856 = n9567 & ~n9568;
  assign n9857 = ~n9565 & ~n9856;
  assign n9858 = ~n9855 & ~n9857;
  assign n9859 = n9855 & n9857;
  assign n9860 = ~n9858 & ~n9859;
  assign n9861 = ~n9579 & n9586;
  assign n9862 = n9582 & ~n9861;
  assign n9863 = n9579 & ~n9586;
  assign n9864 = ~n9862 & ~n9863;
  assign n9865 = ~n9860 & n9864;
  assign n9866 = n9860 & ~n9864;
  assign n9867 = ~n9865 & ~n9866;
  assign n9868 = n9536 & ~n9550;
  assign n9869 = ~n9551 & ~n9868;
  assign n9870 = n9537 & ~n9540;
  assign n9871 = n9543 & ~n9870;
  assign n9872 = ~n9537 & n9540;
  assign n9873 = ~n9871 & ~n9872;
  assign n9874 = ~n9869 & n9873;
  assign n9875 = n9869 & ~n9873;
  assign n9876 = ~n9874 & ~n9875;
  assign n9877 = n9530 & ~n9531;
  assign n9878 = ~n9528 & ~n9877;
  assign n9879 = n9876 & ~n9878;
  assign n9880 = ~n9876 & n9878;
  assign n9881 = ~n9879 & ~n9880;
  assign n9882 = n9867 & ~n9881;
  assign n9883 = ~n9867 & n9881;
  assign n9884 = ~n9882 & ~n9883;
  assign n9885 = ~n9557 & n9592;
  assign n9886 = ~n9556 & ~n9885;
  assign n9887 = n9884 & ~n9886;
  assign n9888 = ~n9884 & n9886;
  assign n9889 = ~n9887 & ~n9888;
  assign n9890 = ~n9497 & ~n9512;
  assign n9891 = ~n9498 & ~n9890;
  assign n9892 = n9490 & ~n9491;
  assign n9893 = ~n9488 & ~n9892;
  assign n9894 = ~n9891 & ~n9893;
  assign n9895 = n9891 & n9893;
  assign n9896 = ~n9894 & ~n9895;
  assign n9897 = ~n9502 & n9509;
  assign n9898 = n9505 & ~n9897;
  assign n9899 = n9502 & ~n9509;
  assign n9900 = ~n9898 & ~n9899;
  assign n9901 = ~n9896 & n9900;
  assign n9902 = n9896 & ~n9900;
  assign n9903 = ~n9901 & ~n9902;
  assign n9904 = n9459 & ~n9473;
  assign n9905 = ~n9474 & ~n9904;
  assign n9906 = n9460 & ~n9463;
  assign n9907 = n9466 & ~n9906;
  assign n9908 = ~n9460 & n9463;
  assign n9909 = ~n9907 & ~n9908;
  assign n9910 = ~n9905 & n9909;
  assign n9911 = n9905 & ~n9909;
  assign n9912 = ~n9910 & ~n9911;
  assign n9913 = n9453 & ~n9454;
  assign n9914 = ~n9451 & ~n9913;
  assign n9915 = n9912 & ~n9914;
  assign n9916 = ~n9912 & n9914;
  assign n9917 = ~n9915 & ~n9916;
  assign n9918 = n9903 & ~n9917;
  assign n9919 = ~n9903 & n9917;
  assign n9920 = ~n9918 & ~n9919;
  assign n9921 = ~n9480 & n9515;
  assign n9922 = ~n9479 & ~n9921;
  assign n9923 = n9920 & ~n9922;
  assign n9924 = ~n9920 & n9922;
  assign n9925 = ~n9923 & ~n9924;
  assign n9926 = ~n9889 & ~n9925;
  assign n9927 = n9889 & n9925;
  assign n9928 = ~n9926 & ~n9927;
  assign n9929 = ~n9520 & ~n9595;
  assign n9930 = ~n9519 & ~n9929;
  assign n9931 = n9928 & ~n9930;
  assign n9932 = ~n9928 & n9930;
  assign n9933 = ~n9931 & ~n9932;
  assign n9934 = ~n9853 & ~n9933;
  assign n9935 = n9853 & n9933;
  assign n9936 = ~n9934 & ~n9935;
  assign n9937 = ~n9600 & ~n9758;
  assign n9938 = ~n9599 & ~n9937;
  assign n9939 = n9936 & ~n9938;
  assign n9940 = ~n9936 & n9938;
  assign n9941 = ~n9939 & ~n9940;
  assign n9942 = ~n9413 & ~n9428;
  assign n9943 = ~n9414 & ~n9942;
  assign n9944 = n9406 & ~n9407;
  assign n9945 = ~n9404 & ~n9944;
  assign n9946 = ~n9943 & ~n9945;
  assign n9947 = n9943 & n9945;
  assign n9948 = ~n9946 & ~n9947;
  assign n9949 = ~n9418 & n9425;
  assign n9950 = n9421 & ~n9949;
  assign n9951 = n9418 & ~n9425;
  assign n9952 = ~n9950 & ~n9951;
  assign n9953 = ~n9948 & n9952;
  assign n9954 = n9948 & ~n9952;
  assign n9955 = ~n9953 & ~n9954;
  assign n9956 = n9375 & ~n9389;
  assign n9957 = ~n9390 & ~n9956;
  assign n9958 = n9376 & ~n9379;
  assign n9959 = n9382 & ~n9958;
  assign n9960 = ~n9376 & n9379;
  assign n9961 = ~n9959 & ~n9960;
  assign n9962 = ~n9957 & n9961;
  assign n9963 = n9957 & ~n9961;
  assign n9964 = ~n9962 & ~n9963;
  assign n9965 = n9369 & ~n9370;
  assign n9966 = ~n9367 & ~n9965;
  assign n9967 = n9964 & ~n9966;
  assign n9968 = ~n9964 & n9966;
  assign n9969 = ~n9967 & ~n9968;
  assign n9970 = n9955 & ~n9969;
  assign n9971 = ~n9955 & n9969;
  assign n9972 = ~n9970 & ~n9971;
  assign n9973 = ~n9396 & n9431;
  assign n9974 = ~n9395 & ~n9973;
  assign n9975 = n9972 & ~n9974;
  assign n9976 = ~n9972 & n9974;
  assign n9977 = ~n9975 & ~n9976;
  assign n9978 = ~n9336 & ~n9351;
  assign n9979 = ~n9337 & ~n9978;
  assign n9980 = n9329 & ~n9330;
  assign n9981 = ~n9327 & ~n9980;
  assign n9982 = ~n9979 & ~n9981;
  assign n9983 = n9979 & n9981;
  assign n9984 = ~n9982 & ~n9983;
  assign n9985 = ~n9341 & n9348;
  assign n9986 = n9344 & ~n9985;
  assign n9987 = n9341 & ~n9348;
  assign n9988 = ~n9986 & ~n9987;
  assign n9989 = ~n9984 & n9988;
  assign n9990 = n9984 & ~n9988;
  assign n9991 = ~n9989 & ~n9990;
  assign n9992 = n9298 & ~n9312;
  assign n9993 = ~n9313 & ~n9992;
  assign n9994 = n9299 & ~n9302;
  assign n9995 = n9305 & ~n9994;
  assign n9996 = ~n9299 & n9302;
  assign n9997 = ~n9995 & ~n9996;
  assign n9998 = ~n9993 & n9997;
  assign n9999 = n9993 & ~n9997;
  assign n10000 = ~n9998 & ~n9999;
  assign n10001 = n9292 & ~n9293;
  assign n10002 = ~n9290 & ~n10001;
  assign n10003 = n10000 & ~n10002;
  assign n10004 = ~n10000 & n10002;
  assign n10005 = ~n10003 & ~n10004;
  assign n10006 = n9991 & ~n10005;
  assign n10007 = ~n9991 & n10005;
  assign n10008 = ~n10006 & ~n10007;
  assign n10009 = ~n9319 & n9354;
  assign n10010 = ~n9318 & ~n10009;
  assign n10011 = n10008 & ~n10010;
  assign n10012 = ~n10008 & n10010;
  assign n10013 = ~n10011 & ~n10012;
  assign n10014 = ~n9977 & ~n10013;
  assign n10015 = n9977 & n10013;
  assign n10016 = ~n10014 & ~n10015;
  assign n10017 = ~n9359 & ~n9434;
  assign n10018 = ~n9358 & ~n10017;
  assign n10019 = n10016 & ~n10018;
  assign n10020 = ~n10016 & n10018;
  assign n10021 = ~n10019 & ~n10020;
  assign n10022 = ~n9255 & ~n9270;
  assign n10023 = ~n9256 & ~n10022;
  assign n10024 = n9248 & ~n9249;
  assign n10025 = ~n9246 & ~n10024;
  assign n10026 = ~n10023 & ~n10025;
  assign n10027 = n10023 & n10025;
  assign n10028 = ~n10026 & ~n10027;
  assign n10029 = ~n9260 & n9267;
  assign n10030 = n9263 & ~n10029;
  assign n10031 = n9260 & ~n9267;
  assign n10032 = ~n10030 & ~n10031;
  assign n10033 = ~n10028 & n10032;
  assign n10034 = n10028 & ~n10032;
  assign n10035 = ~n10033 & ~n10034;
  assign n10036 = n9217 & ~n9231;
  assign n10037 = ~n9232 & ~n10036;
  assign n10038 = n9218 & ~n9221;
  assign n10039 = n9224 & ~n10038;
  assign n10040 = ~n9218 & n9221;
  assign n10041 = ~n10039 & ~n10040;
  assign n10042 = ~n10037 & n10041;
  assign n10043 = n10037 & ~n10041;
  assign n10044 = ~n10042 & ~n10043;
  assign n10045 = n9211 & ~n9212;
  assign n10046 = ~n9209 & ~n10045;
  assign n10047 = n10044 & ~n10046;
  assign n10048 = ~n10044 & n10046;
  assign n10049 = ~n10047 & ~n10048;
  assign n10050 = n10035 & ~n10049;
  assign n10051 = ~n10035 & n10049;
  assign n10052 = ~n10050 & ~n10051;
  assign n10053 = ~n9238 & n9273;
  assign n10054 = ~n9237 & ~n10053;
  assign n10055 = n10052 & ~n10054;
  assign n10056 = ~n10052 & n10054;
  assign n10057 = ~n10055 & ~n10056;
  assign n10058 = ~n9178 & ~n9193;
  assign n10059 = ~n9179 & ~n10058;
  assign n10060 = n9171 & ~n9172;
  assign n10061 = ~n9169 & ~n10060;
  assign n10062 = ~n10059 & ~n10061;
  assign n10063 = n10059 & n10061;
  assign n10064 = ~n10062 & ~n10063;
  assign n10065 = ~n9183 & n9190;
  assign n10066 = n9186 & ~n10065;
  assign n10067 = n9183 & ~n9190;
  assign n10068 = ~n10066 & ~n10067;
  assign n10069 = ~n10064 & n10068;
  assign n10070 = n10064 & ~n10068;
  assign n10071 = ~n10069 & ~n10070;
  assign n10072 = n9140 & ~n9154;
  assign n10073 = ~n9155 & ~n10072;
  assign n10074 = n9141 & ~n9144;
  assign n10075 = n9147 & ~n10074;
  assign n10076 = ~n9141 & n9144;
  assign n10077 = ~n10075 & ~n10076;
  assign n10078 = ~n10073 & n10077;
  assign n10079 = n10073 & ~n10077;
  assign n10080 = ~n10078 & ~n10079;
  assign n10081 = n9134 & ~n9135;
  assign n10082 = ~n9132 & ~n10081;
  assign n10083 = n10080 & ~n10082;
  assign n10084 = ~n10080 & n10082;
  assign n10085 = ~n10083 & ~n10084;
  assign n10086 = n10071 & ~n10085;
  assign n10087 = ~n10071 & n10085;
  assign n10088 = ~n10086 & ~n10087;
  assign n10089 = ~n9161 & n9196;
  assign n10090 = ~n9160 & ~n10089;
  assign n10091 = n10088 & ~n10090;
  assign n10092 = ~n10088 & n10090;
  assign n10093 = ~n10091 & ~n10092;
  assign n10094 = ~n10057 & ~n10093;
  assign n10095 = n10057 & n10093;
  assign n10096 = ~n10094 & ~n10095;
  assign n10097 = ~n9201 & ~n9276;
  assign n10098 = ~n9200 & ~n10097;
  assign n10099 = n10096 & ~n10098;
  assign n10100 = ~n10096 & n10098;
  assign n10101 = ~n10099 & ~n10100;
  assign n10102 = ~n10021 & ~n10101;
  assign n10103 = n10021 & n10101;
  assign n10104 = ~n10102 & ~n10103;
  assign n10105 = ~n9281 & ~n9437;
  assign n10106 = ~n9280 & ~n10105;
  assign n10107 = n10104 & ~n10106;
  assign n10108 = ~n10104 & n10106;
  assign n10109 = ~n10107 & ~n10108;
  assign n10110 = ~n9941 & ~n10109;
  assign n10111 = n9941 & n10109;
  assign n10112 = ~n10110 & ~n10111;
  assign n10113 = ~n9442 & ~n9761;
  assign n10114 = ~n9441 & ~n10113;
  assign n10115 = n10112 & ~n10114;
  assign n10116 = ~n10112 & n10114;
  assign n10117 = ~n10115 & ~n10116;
  assign n10118 = ~n9091 & ~n9106;
  assign n10119 = ~n9092 & ~n10118;
  assign n10120 = n9084 & ~n9085;
  assign n10121 = ~n9082 & ~n10120;
  assign n10122 = ~n10119 & ~n10121;
  assign n10123 = n10119 & n10121;
  assign n10124 = ~n10122 & ~n10123;
  assign n10125 = ~n9096 & n9103;
  assign n10126 = n9099 & ~n10125;
  assign n10127 = n9096 & ~n9103;
  assign n10128 = ~n10126 & ~n10127;
  assign n10129 = ~n10124 & n10128;
  assign n10130 = n10124 & ~n10128;
  assign n10131 = ~n10129 & ~n10130;
  assign n10132 = n9053 & ~n9067;
  assign n10133 = ~n9068 & ~n10132;
  assign n10134 = n9054 & ~n9057;
  assign n10135 = n9060 & ~n10134;
  assign n10136 = ~n9054 & n9057;
  assign n10137 = ~n10135 & ~n10136;
  assign n10138 = ~n10133 & n10137;
  assign n10139 = n10133 & ~n10137;
  assign n10140 = ~n10138 & ~n10139;
  assign n10141 = n9047 & ~n9048;
  assign n10142 = ~n9045 & ~n10141;
  assign n10143 = n10140 & ~n10142;
  assign n10144 = ~n10140 & n10142;
  assign n10145 = ~n10143 & ~n10144;
  assign n10146 = n10131 & ~n10145;
  assign n10147 = ~n10131 & n10145;
  assign n10148 = ~n10146 & ~n10147;
  assign n10149 = ~n9074 & n9109;
  assign n10150 = ~n9073 & ~n10149;
  assign n10151 = n10148 & ~n10150;
  assign n10152 = ~n10148 & n10150;
  assign n10153 = ~n10151 & ~n10152;
  assign n10154 = ~n9014 & ~n9029;
  assign n10155 = ~n9015 & ~n10154;
  assign n10156 = n9007 & ~n9008;
  assign n10157 = ~n9005 & ~n10156;
  assign n10158 = ~n10155 & ~n10157;
  assign n10159 = n10155 & n10157;
  assign n10160 = ~n10158 & ~n10159;
  assign n10161 = ~n9019 & n9026;
  assign n10162 = n9022 & ~n10161;
  assign n10163 = n9019 & ~n9026;
  assign n10164 = ~n10162 & ~n10163;
  assign n10165 = ~n10160 & n10164;
  assign n10166 = n10160 & ~n10164;
  assign n10167 = ~n10165 & ~n10166;
  assign n10168 = n8976 & ~n8990;
  assign n10169 = ~n8991 & ~n10168;
  assign n10170 = n8977 & ~n8980;
  assign n10171 = n8983 & ~n10170;
  assign n10172 = ~n8977 & n8980;
  assign n10173 = ~n10171 & ~n10172;
  assign n10174 = ~n10169 & n10173;
  assign n10175 = n10169 & ~n10173;
  assign n10176 = ~n10174 & ~n10175;
  assign n10177 = n8970 & ~n8971;
  assign n10178 = ~n8968 & ~n10177;
  assign n10179 = n10176 & ~n10178;
  assign n10180 = ~n10176 & n10178;
  assign n10181 = ~n10179 & ~n10180;
  assign n10182 = n10167 & ~n10181;
  assign n10183 = ~n10167 & n10181;
  assign n10184 = ~n10182 & ~n10183;
  assign n10185 = ~n8997 & n9032;
  assign n10186 = ~n8996 & ~n10185;
  assign n10187 = n10184 & ~n10186;
  assign n10188 = ~n10184 & n10186;
  assign n10189 = ~n10187 & ~n10188;
  assign n10190 = ~n10153 & ~n10189;
  assign n10191 = n10153 & n10189;
  assign n10192 = ~n10190 & ~n10191;
  assign n10193 = ~n9037 & ~n9112;
  assign n10194 = ~n9036 & ~n10193;
  assign n10195 = n10192 & ~n10194;
  assign n10196 = ~n10192 & n10194;
  assign n10197 = ~n10195 & ~n10196;
  assign n10198 = ~n8933 & ~n8948;
  assign n10199 = ~n8934 & ~n10198;
  assign n10200 = n8926 & ~n8927;
  assign n10201 = ~n8924 & ~n10200;
  assign n10202 = ~n10199 & ~n10201;
  assign n10203 = n10199 & n10201;
  assign n10204 = ~n10202 & ~n10203;
  assign n10205 = ~n8938 & n8945;
  assign n10206 = n8941 & ~n10205;
  assign n10207 = n8938 & ~n8945;
  assign n10208 = ~n10206 & ~n10207;
  assign n10209 = ~n10204 & n10208;
  assign n10210 = n10204 & ~n10208;
  assign n10211 = ~n10209 & ~n10210;
  assign n10212 = n8895 & ~n8910;
  assign n10213 = n8257 & ~n8909;
  assign n10214 = ~n10212 & ~n10213;
  assign n10215 = n8889 & ~n8890;
  assign n10216 = ~n8887 & ~n10215;
  assign n10217 = ~n10214 & ~n10216;
  assign n10218 = n10214 & n10216;
  assign n10219 = ~n10217 & ~n10218;
  assign n10220 = ~n8898 & n8906;
  assign n10221 = n8901 & ~n10220;
  assign n10222 = n8898 & ~n8906;
  assign n10223 = ~n10221 & ~n10222;
  assign n10224 = ~n10219 & n10223;
  assign n10225 = n10219 & ~n10223;
  assign n10226 = ~n10224 & ~n10225;
  assign n10227 = n10211 & n10226;
  assign n10228 = ~n10211 & ~n10226;
  assign n10229 = ~n10227 & ~n10228;
  assign n10230 = ~n8916 & n8951;
  assign n10231 = ~n8915 & ~n10230;
  assign n10232 = n10229 & ~n10231;
  assign n10233 = ~n10229 & n10231;
  assign n10234 = ~n10232 & ~n10233;
  assign n10235 = ~n8856 & ~n8871;
  assign n10236 = ~n8857 & ~n10235;
  assign n10237 = n8849 & ~n8850;
  assign n10238 = ~n8847 & ~n10237;
  assign n10239 = ~n10236 & ~n10238;
  assign n10240 = n10236 & n10238;
  assign n10241 = ~n10239 & ~n10240;
  assign n10242 = n8859 & ~n8862;
  assign n10243 = n8865 & ~n10242;
  assign n10244 = ~n8859 & n8862;
  assign n10245 = ~n10243 & ~n10244;
  assign n10246 = ~n10241 & n10245;
  assign n10247 = n10241 & ~n10245;
  assign n10248 = ~n10246 & ~n10247;
  assign n10249 = n8818 & ~n8833;
  assign n10250 = n8180 & ~n8832;
  assign n10251 = ~n10249 & ~n10250;
  assign n10252 = n8812 & ~n8813;
  assign n10253 = ~n8810 & ~n10252;
  assign n10254 = ~n10251 & ~n10253;
  assign n10255 = n10251 & n10253;
  assign n10256 = ~n10254 & ~n10255;
  assign n10257 = ~n8821 & n8829;
  assign n10258 = n8824 & ~n10257;
  assign n10259 = n8821 & ~n8829;
  assign n10260 = ~n10258 & ~n10259;
  assign n10261 = ~n10256 & n10260;
  assign n10262 = n10256 & ~n10260;
  assign n10263 = ~n10261 & ~n10262;
  assign n10264 = n10248 & n10263;
  assign n10265 = ~n10248 & ~n10263;
  assign n10266 = ~n10264 & ~n10265;
  assign n10267 = ~n8839 & n8874;
  assign n10268 = ~n8838 & ~n10267;
  assign n10269 = n10266 & ~n10268;
  assign n10270 = ~n10266 & n10268;
  assign n10271 = ~n10269 & ~n10270;
  assign n10272 = ~n10234 & ~n10271;
  assign n10273 = n10234 & n10271;
  assign n10274 = ~n10272 & ~n10273;
  assign n10275 = ~n8879 & ~n8954;
  assign n10276 = ~n8878 & ~n10275;
  assign n10277 = n10274 & ~n10276;
  assign n10278 = ~n10274 & n10276;
  assign n10279 = ~n10277 & ~n10278;
  assign n10280 = ~n10197 & ~n10279;
  assign n10281 = n10197 & n10279;
  assign n10282 = ~n10280 & ~n10281;
  assign n10283 = ~n8959 & ~n9115;
  assign n10284 = ~n8958 & ~n10283;
  assign n10285 = n10282 & ~n10284;
  assign n10286 = ~n10282 & n10284;
  assign n10287 = ~n10285 & ~n10286;
  assign n10288 = ~n8772 & ~n8787;
  assign n10289 = ~n8773 & ~n10288;
  assign n10290 = n8765 & ~n8766;
  assign n10291 = ~n8763 & ~n10290;
  assign n10292 = ~n10289 & ~n10291;
  assign n10293 = n10289 & n10291;
  assign n10294 = ~n10292 & ~n10293;
  assign n10295 = ~n8777 & n8784;
  assign n10296 = n8780 & ~n10295;
  assign n10297 = n8777 & ~n8784;
  assign n10298 = ~n10296 & ~n10297;
  assign n10299 = ~n10294 & n10298;
  assign n10300 = n10294 & ~n10298;
  assign n10301 = ~n10299 & ~n10300;
  assign n10302 = n8734 & ~n8748;
  assign n10303 = ~n8749 & ~n10302;
  assign n10304 = n8735 & ~n8738;
  assign n10305 = n8741 & ~n10304;
  assign n10306 = ~n8735 & n8738;
  assign n10307 = ~n10305 & ~n10306;
  assign n10308 = ~n10303 & n10307;
  assign n10309 = n10303 & ~n10307;
  assign n10310 = ~n10308 & ~n10309;
  assign n10311 = n8728 & ~n8729;
  assign n10312 = ~n8726 & ~n10311;
  assign n10313 = n10310 & ~n10312;
  assign n10314 = ~n10310 & n10312;
  assign n10315 = ~n10313 & ~n10314;
  assign n10316 = n10301 & ~n10315;
  assign n10317 = ~n10301 & n10315;
  assign n10318 = ~n10316 & ~n10317;
  assign n10319 = ~n8755 & n8790;
  assign n10320 = ~n8754 & ~n10319;
  assign n10321 = n10318 & ~n10320;
  assign n10322 = ~n10318 & n10320;
  assign n10323 = ~n10321 & ~n10322;
  assign n10324 = ~n8695 & ~n8710;
  assign n10325 = ~n8696 & ~n10324;
  assign n10326 = n8688 & ~n8689;
  assign n10327 = ~n8686 & ~n10326;
  assign n10328 = ~n10325 & ~n10327;
  assign n10329 = n10325 & n10327;
  assign n10330 = ~n10328 & ~n10329;
  assign n10331 = n8698 & ~n8701;
  assign n10332 = n8704 & ~n10331;
  assign n10333 = ~n8698 & n8701;
  assign n10334 = ~n10332 & ~n10333;
  assign n10335 = ~n10330 & n10334;
  assign n10336 = n10330 & ~n10334;
  assign n10337 = ~n10335 & ~n10336;
  assign n10338 = n8657 & ~n8672;
  assign n10339 = n8020 & ~n8671;
  assign n10340 = ~n10338 & ~n10339;
  assign n10341 = n8651 & ~n8652;
  assign n10342 = ~n8649 & ~n10341;
  assign n10343 = ~n10340 & ~n10342;
  assign n10344 = n10340 & n10342;
  assign n10345 = ~n10343 & ~n10344;
  assign n10346 = ~n8660 & n8668;
  assign n10347 = n8663 & ~n10346;
  assign n10348 = n8660 & ~n8668;
  assign n10349 = ~n10347 & ~n10348;
  assign n10350 = ~n10345 & n10349;
  assign n10351 = n10345 & ~n10349;
  assign n10352 = ~n10350 & ~n10351;
  assign n10353 = n10337 & n10352;
  assign n10354 = ~n10337 & ~n10352;
  assign n10355 = ~n10353 & ~n10354;
  assign n10356 = ~n8678 & n8713;
  assign n10357 = ~n8677 & ~n10356;
  assign n10358 = n10355 & ~n10357;
  assign n10359 = ~n10355 & n10357;
  assign n10360 = ~n10358 & ~n10359;
  assign n10361 = ~n10323 & ~n10360;
  assign n10362 = n10323 & n10360;
  assign n10363 = ~n10361 & ~n10362;
  assign n10364 = ~n8718 & ~n8793;
  assign n10365 = ~n8717 & ~n10364;
  assign n10366 = n10363 & ~n10365;
  assign n10367 = ~n10363 & n10365;
  assign n10368 = ~n10366 & ~n10367;
  assign n10369 = ~n8614 & ~n8629;
  assign n10370 = ~n8615 & ~n10369;
  assign n10371 = n8607 & ~n8608;
  assign n10372 = ~n8605 & ~n10371;
  assign n10373 = ~n10370 & ~n10372;
  assign n10374 = n10370 & n10372;
  assign n10375 = ~n10373 & ~n10374;
  assign n10376 = ~n8619 & n8626;
  assign n10377 = n8622 & ~n10376;
  assign n10378 = n8619 & ~n8626;
  assign n10379 = ~n10377 & ~n10378;
  assign n10380 = ~n10375 & n10379;
  assign n10381 = n10375 & ~n10379;
  assign n10382 = ~n10380 & ~n10381;
  assign n10383 = n8576 & ~n8591;
  assign n10384 = n7940 & ~n8590;
  assign n10385 = ~n10383 & ~n10384;
  assign n10386 = n8570 & ~n8571;
  assign n10387 = ~n8568 & ~n10386;
  assign n10388 = ~n10385 & ~n10387;
  assign n10389 = n10385 & n10387;
  assign n10390 = ~n10388 & ~n10389;
  assign n10391 = ~n8579 & n8587;
  assign n10392 = n8582 & ~n10391;
  assign n10393 = n8579 & ~n8587;
  assign n10394 = ~n10392 & ~n10393;
  assign n10395 = ~n10390 & n10394;
  assign n10396 = n10390 & ~n10394;
  assign n10397 = ~n10395 & ~n10396;
  assign n10398 = n10382 & n10397;
  assign n10399 = ~n10382 & ~n10397;
  assign n10400 = ~n10398 & ~n10399;
  assign n10401 = ~n8597 & n8632;
  assign n10402 = ~n8596 & ~n10401;
  assign n10403 = n10400 & ~n10402;
  assign n10404 = ~n10400 & n10402;
  assign n10405 = ~n10403 & ~n10404;
  assign n10406 = ~n8537 & ~n8552;
  assign n10407 = ~n8538 & ~n10406;
  assign n10408 = n8530 & ~n8531;
  assign n10409 = ~n8528 & ~n10408;
  assign n10410 = ~n10407 & ~n10409;
  assign n10411 = n10407 & n10409;
  assign n10412 = ~n10410 & ~n10411;
  assign n10413 = n8540 & ~n8543;
  assign n10414 = n8546 & ~n10413;
  assign n10415 = ~n8540 & n8543;
  assign n10416 = ~n10414 & ~n10415;
  assign n10417 = ~n10412 & n10416;
  assign n10418 = n10412 & ~n10416;
  assign n10419 = ~n10417 & ~n10418;
  assign n10420 = n8499 & ~n8514;
  assign n10421 = n7863 & ~n8513;
  assign n10422 = ~n10420 & ~n10421;
  assign n10423 = n8493 & ~n8494;
  assign n10424 = ~n8491 & ~n10423;
  assign n10425 = ~n10422 & ~n10424;
  assign n10426 = n10422 & n10424;
  assign n10427 = ~n10425 & ~n10426;
  assign n10428 = ~n8502 & n8510;
  assign n10429 = n8505 & ~n10428;
  assign n10430 = n8502 & ~n8510;
  assign n10431 = ~n10429 & ~n10430;
  assign n10432 = ~n10427 & n10431;
  assign n10433 = n10427 & ~n10431;
  assign n10434 = ~n10432 & ~n10433;
  assign n10435 = n10419 & n10434;
  assign n10436 = ~n10419 & ~n10434;
  assign n10437 = ~n10435 & ~n10436;
  assign n10438 = ~n8520 & n8555;
  assign n10439 = ~n8519 & ~n10438;
  assign n10440 = n10437 & ~n10439;
  assign n10441 = ~n10437 & n10439;
  assign n10442 = ~n10440 & ~n10441;
  assign n10443 = ~n10405 & ~n10442;
  assign n10444 = n10405 & n10442;
  assign n10445 = ~n10443 & ~n10444;
  assign n10446 = ~n8560 & ~n8635;
  assign n10447 = ~n8559 & ~n10446;
  assign n10448 = n10445 & ~n10447;
  assign n10449 = ~n10445 & n10447;
  assign n10450 = ~n10448 & ~n10449;
  assign n10451 = ~n10368 & ~n10450;
  assign n10452 = n10368 & n10450;
  assign n10453 = ~n10451 & ~n10452;
  assign n10454 = ~n8640 & ~n8796;
  assign n10455 = ~n8639 & ~n10454;
  assign n10456 = n10453 & ~n10455;
  assign n10457 = ~n10453 & n10455;
  assign n10458 = ~n10456 & ~n10457;
  assign n10459 = ~n10287 & ~n10458;
  assign n10460 = n10287 & n10458;
  assign n10461 = ~n10459 & ~n10460;
  assign n10462 = ~n8801 & ~n9118;
  assign n10463 = ~n8800 & ~n10462;
  assign n10464 = n10461 & ~n10463;
  assign n10465 = ~n10461 & n10463;
  assign n10466 = ~n10464 & ~n10465;
  assign n10467 = ~n10117 & ~n10466;
  assign n10468 = n10117 & n10466;
  assign n10469 = ~n10467 & ~n10468;
  assign n10470 = ~n9123 & n9764;
  assign n10471 = ~n9122 & ~n10470;
  assign n10472 = n10469 & ~n10471;
  assign n10473 = ~n10469 & n10471;
  assign n10474 = ~n10472 & ~n10473;
  assign n10475 = ~n9775 & ~n10474;
  assign n10476 = n9775 & n10474;
  assign n10477 = ~n10475 & ~n10476;
  assign n10478 = ~n8480 & ~n9767;
  assign n10479 = ~n8481 & ~n10478;
  assign n10480 = n10477 & ~n10479;
  assign n10481 = ~n10477 & n10479;
  assign n10482 = ~n10480 & ~n10481;
  assign n10483 = n9771 & n10482;
  assign n10484 = ~n7148 & ~n7149;
  assign n10485 = n7179 & n10484;
  assign n10486 = ~n7179 & ~n10484;
  assign n10487 = ~n10485 & ~n10486;
  assign n10488 = ~n10435 & ~n10439;
  assign n10489 = ~n10436 & ~n10488;
  assign n10490 = ~n10426 & n10431;
  assign n10491 = ~n10425 & ~n10490;
  assign n10492 = n10489 & n10491;
  assign n10493 = ~n10489 & ~n10491;
  assign n10494 = ~n10492 & ~n10493;
  assign n10495 = ~n10411 & n10416;
  assign n10496 = ~n10410 & ~n10495;
  assign n10497 = ~n10494 & n10496;
  assign n10498 = ~n10492 & ~n10496;
  assign n10499 = ~n10493 & n10498;
  assign n10500 = ~n10497 & ~n10499;
  assign n10501 = ~n10398 & ~n10402;
  assign n10502 = ~n10399 & ~n10501;
  assign n10503 = ~n10389 & n10394;
  assign n10504 = ~n10388 & ~n10503;
  assign n10505 = n10502 & n10504;
  assign n10506 = ~n10502 & ~n10504;
  assign n10507 = ~n10505 & ~n10506;
  assign n10508 = ~n10374 & n10379;
  assign n10509 = ~n10373 & ~n10508;
  assign n10510 = ~n10507 & n10509;
  assign n10511 = ~n10505 & ~n10509;
  assign n10512 = ~n10506 & n10511;
  assign n10513 = ~n10510 & ~n10512;
  assign n10514 = ~n10500 & ~n10513;
  assign n10515 = n10500 & n10513;
  assign n10516 = ~n10514 & ~n10515;
  assign n10517 = ~n10444 & n10447;
  assign n10518 = ~n10443 & ~n10517;
  assign n10519 = n10516 & ~n10518;
  assign n10520 = ~n10516 & n10518;
  assign n10521 = ~n10519 & ~n10520;
  assign n10522 = ~n10353 & ~n10357;
  assign n10523 = ~n10354 & ~n10522;
  assign n10524 = ~n10344 & n10349;
  assign n10525 = ~n10343 & ~n10524;
  assign n10526 = n10523 & n10525;
  assign n10527 = ~n10523 & ~n10525;
  assign n10528 = ~n10526 & ~n10527;
  assign n10529 = ~n10329 & n10334;
  assign n10530 = ~n10328 & ~n10529;
  assign n10531 = ~n10528 & n10530;
  assign n10532 = ~n10526 & ~n10530;
  assign n10533 = ~n10527 & n10532;
  assign n10534 = ~n10531 & ~n10533;
  assign n10535 = ~n10317 & n10320;
  assign n10536 = ~n10316 & ~n10535;
  assign n10537 = ~n10309 & ~n10312;
  assign n10538 = ~n10308 & ~n10537;
  assign n10539 = ~n10536 & n10538;
  assign n10540 = n10536 & ~n10538;
  assign n10541 = ~n10539 & ~n10540;
  assign n10542 = ~n10293 & n10298;
  assign n10543 = ~n10292 & ~n10542;
  assign n10544 = n10541 & n10543;
  assign n10545 = ~n10541 & ~n10543;
  assign n10546 = ~n10544 & ~n10545;
  assign n10547 = ~n10534 & n10546;
  assign n10548 = n10534 & ~n10546;
  assign n10549 = ~n10547 & ~n10548;
  assign n10550 = ~n10362 & n10365;
  assign n10551 = ~n10361 & ~n10550;
  assign n10552 = n10549 & ~n10551;
  assign n10553 = ~n10549 & n10551;
  assign n10554 = ~n10552 & ~n10553;
  assign n10555 = n10521 & n10554;
  assign n10556 = ~n10521 & ~n10554;
  assign n10557 = ~n10555 & ~n10556;
  assign n10558 = ~n10452 & n10455;
  assign n10559 = ~n10451 & ~n10558;
  assign n10560 = n10557 & n10559;
  assign n10561 = ~n10557 & ~n10559;
  assign n10562 = ~n10560 & ~n10561;
  assign n10563 = ~n10264 & ~n10268;
  assign n10564 = ~n10265 & ~n10563;
  assign n10565 = ~n10255 & n10260;
  assign n10566 = ~n10254 & ~n10565;
  assign n10567 = n10564 & n10566;
  assign n10568 = ~n10564 & ~n10566;
  assign n10569 = ~n10567 & ~n10568;
  assign n10570 = ~n10240 & n10245;
  assign n10571 = ~n10239 & ~n10570;
  assign n10572 = ~n10569 & n10571;
  assign n10573 = ~n10567 & ~n10571;
  assign n10574 = ~n10568 & n10573;
  assign n10575 = ~n10572 & ~n10574;
  assign n10576 = ~n10227 & ~n10231;
  assign n10577 = ~n10228 & ~n10576;
  assign n10578 = ~n10218 & n10223;
  assign n10579 = ~n10217 & ~n10578;
  assign n10580 = n10577 & n10579;
  assign n10581 = ~n10577 & ~n10579;
  assign n10582 = ~n10580 & ~n10581;
  assign n10583 = ~n10203 & n10208;
  assign n10584 = ~n10202 & ~n10583;
  assign n10585 = ~n10582 & n10584;
  assign n10586 = ~n10580 & ~n10584;
  assign n10587 = ~n10581 & n10586;
  assign n10588 = ~n10585 & ~n10587;
  assign n10589 = ~n10575 & ~n10588;
  assign n10590 = n10575 & n10588;
  assign n10591 = ~n10589 & ~n10590;
  assign n10592 = ~n10273 & n10276;
  assign n10593 = ~n10272 & ~n10592;
  assign n10594 = n10591 & ~n10593;
  assign n10595 = ~n10591 & n10593;
  assign n10596 = ~n10594 & ~n10595;
  assign n10597 = ~n10183 & n10186;
  assign n10598 = ~n10182 & ~n10597;
  assign n10599 = ~n10175 & ~n10178;
  assign n10600 = ~n10174 & ~n10599;
  assign n10601 = ~n10598 & n10600;
  assign n10602 = n10598 & ~n10600;
  assign n10603 = ~n10601 & ~n10602;
  assign n10604 = ~n10159 & n10164;
  assign n10605 = ~n10158 & ~n10604;
  assign n10606 = n10603 & n10605;
  assign n10607 = ~n10603 & ~n10605;
  assign n10608 = ~n10606 & ~n10607;
  assign n10609 = ~n10147 & n10150;
  assign n10610 = ~n10146 & ~n10609;
  assign n10611 = ~n10139 & ~n10142;
  assign n10612 = ~n10138 & ~n10611;
  assign n10613 = ~n10610 & n10612;
  assign n10614 = n10610 & ~n10612;
  assign n10615 = ~n10613 & ~n10614;
  assign n10616 = ~n10123 & n10128;
  assign n10617 = ~n10122 & ~n10616;
  assign n10618 = n10615 & n10617;
  assign n10619 = ~n10615 & ~n10617;
  assign n10620 = ~n10618 & ~n10619;
  assign n10621 = n10608 & n10620;
  assign n10622 = ~n10608 & ~n10620;
  assign n10623 = ~n10621 & ~n10622;
  assign n10624 = ~n10191 & n10194;
  assign n10625 = ~n10190 & ~n10624;
  assign n10626 = n10623 & ~n10625;
  assign n10627 = ~n10623 & n10625;
  assign n10628 = ~n10626 & ~n10627;
  assign n10629 = n10596 & n10628;
  assign n10630 = ~n10596 & ~n10628;
  assign n10631 = ~n10629 & ~n10630;
  assign n10632 = ~n10281 & n10284;
  assign n10633 = ~n10280 & ~n10632;
  assign n10634 = n10631 & n10633;
  assign n10635 = ~n10631 & ~n10633;
  assign n10636 = ~n10634 & ~n10635;
  assign n10637 = ~n10562 & ~n10636;
  assign n10638 = n10562 & n10636;
  assign n10639 = ~n10637 & ~n10638;
  assign n10640 = ~n10460 & n10463;
  assign n10641 = ~n10459 & ~n10640;
  assign n10642 = n10639 & ~n10641;
  assign n10643 = ~n10639 & n10641;
  assign n10644 = ~n10642 & ~n10643;
  assign n10645 = ~n10087 & n10090;
  assign n10646 = ~n10086 & ~n10645;
  assign n10647 = ~n10079 & ~n10082;
  assign n10648 = ~n10078 & ~n10647;
  assign n10649 = ~n10646 & n10648;
  assign n10650 = n10646 & ~n10648;
  assign n10651 = ~n10649 & ~n10650;
  assign n10652 = ~n10063 & n10068;
  assign n10653 = ~n10062 & ~n10652;
  assign n10654 = n10651 & n10653;
  assign n10655 = ~n10651 & ~n10653;
  assign n10656 = ~n10654 & ~n10655;
  assign n10657 = ~n10051 & n10054;
  assign n10658 = ~n10050 & ~n10657;
  assign n10659 = ~n10043 & ~n10046;
  assign n10660 = ~n10042 & ~n10659;
  assign n10661 = ~n10658 & n10660;
  assign n10662 = n10658 & ~n10660;
  assign n10663 = ~n10661 & ~n10662;
  assign n10664 = ~n10027 & n10032;
  assign n10665 = ~n10026 & ~n10664;
  assign n10666 = n10663 & n10665;
  assign n10667 = ~n10663 & ~n10665;
  assign n10668 = ~n10666 & ~n10667;
  assign n10669 = n10656 & n10668;
  assign n10670 = ~n10656 & ~n10668;
  assign n10671 = ~n10669 & ~n10670;
  assign n10672 = ~n10095 & n10098;
  assign n10673 = ~n10094 & ~n10672;
  assign n10674 = n10671 & ~n10673;
  assign n10675 = ~n10671 & n10673;
  assign n10676 = ~n10674 & ~n10675;
  assign n10677 = ~n10007 & n10010;
  assign n10678 = ~n10006 & ~n10677;
  assign n10679 = ~n9999 & ~n10002;
  assign n10680 = ~n9998 & ~n10679;
  assign n10681 = ~n10678 & n10680;
  assign n10682 = n10678 & ~n10680;
  assign n10683 = ~n10681 & ~n10682;
  assign n10684 = ~n9983 & n9988;
  assign n10685 = ~n9982 & ~n10684;
  assign n10686 = n10683 & n10685;
  assign n10687 = ~n10683 & ~n10685;
  assign n10688 = ~n10686 & ~n10687;
  assign n10689 = ~n9971 & n9974;
  assign n10690 = ~n9970 & ~n10689;
  assign n10691 = ~n9963 & ~n9966;
  assign n10692 = ~n9962 & ~n10691;
  assign n10693 = ~n10690 & n10692;
  assign n10694 = n10690 & ~n10692;
  assign n10695 = ~n10693 & ~n10694;
  assign n10696 = ~n9947 & n9952;
  assign n10697 = ~n9946 & ~n10696;
  assign n10698 = n10695 & n10697;
  assign n10699 = ~n10695 & ~n10697;
  assign n10700 = ~n10698 & ~n10699;
  assign n10701 = n10688 & n10700;
  assign n10702 = ~n10688 & ~n10700;
  assign n10703 = ~n10701 & ~n10702;
  assign n10704 = ~n10015 & n10018;
  assign n10705 = ~n10014 & ~n10704;
  assign n10706 = n10703 & ~n10705;
  assign n10707 = ~n10703 & n10705;
  assign n10708 = ~n10706 & ~n10707;
  assign n10709 = n10676 & n10708;
  assign n10710 = ~n10676 & ~n10708;
  assign n10711 = ~n10709 & ~n10710;
  assign n10712 = ~n10103 & n10106;
  assign n10713 = ~n10102 & ~n10712;
  assign n10714 = n10711 & n10713;
  assign n10715 = ~n10711 & ~n10713;
  assign n10716 = ~n10714 & ~n10715;
  assign n10717 = ~n9919 & n9922;
  assign n10718 = ~n9918 & ~n10717;
  assign n10719 = ~n9911 & ~n9914;
  assign n10720 = ~n9910 & ~n10719;
  assign n10721 = ~n10718 & n10720;
  assign n10722 = n10718 & ~n10720;
  assign n10723 = ~n10721 & ~n10722;
  assign n10724 = ~n9895 & n9900;
  assign n10725 = ~n9894 & ~n10724;
  assign n10726 = n10723 & n10725;
  assign n10727 = ~n10723 & ~n10725;
  assign n10728 = ~n10726 & ~n10727;
  assign n10729 = ~n9883 & n9886;
  assign n10730 = ~n9882 & ~n10729;
  assign n10731 = ~n9875 & ~n9878;
  assign n10732 = ~n9874 & ~n10731;
  assign n10733 = ~n10730 & n10732;
  assign n10734 = n10730 & ~n10732;
  assign n10735 = ~n10733 & ~n10734;
  assign n10736 = ~n9859 & n9864;
  assign n10737 = ~n9858 & ~n10736;
  assign n10738 = n10735 & n10737;
  assign n10739 = ~n10735 & ~n10737;
  assign n10740 = ~n10738 & ~n10739;
  assign n10741 = n10728 & n10740;
  assign n10742 = ~n10728 & ~n10740;
  assign n10743 = ~n10741 & ~n10742;
  assign n10744 = ~n9927 & n9930;
  assign n10745 = ~n9926 & ~n10744;
  assign n10746 = n10743 & ~n10745;
  assign n10747 = ~n10743 & n10745;
  assign n10748 = ~n10746 & ~n10747;
  assign n10749 = ~n9839 & n9842;
  assign n10750 = ~n9838 & ~n10749;
  assign n10751 = ~n9831 & ~n9834;
  assign n10752 = ~n9830 & ~n10751;
  assign n10753 = ~n10750 & n10752;
  assign n10754 = n10750 & ~n10752;
  assign n10755 = ~n10753 & ~n10754;
  assign n10756 = ~n9815 & n9820;
  assign n10757 = ~n9814 & ~n10756;
  assign n10758 = n10755 & n10757;
  assign n10759 = ~n10755 & ~n10757;
  assign n10760 = ~n10758 & ~n10759;
  assign n10761 = ~n9803 & n9806;
  assign n10762 = ~n9802 & ~n10761;
  assign n10763 = ~n9795 & ~n9798;
  assign n10764 = ~n9794 & ~n10763;
  assign n10765 = ~n10762 & n10764;
  assign n10766 = n10762 & ~n10764;
  assign n10767 = ~n10765 & ~n10766;
  assign n10768 = ~n9781 & n9784;
  assign n10769 = ~n9780 & ~n10768;
  assign n10770 = n10767 & n10769;
  assign n10771 = ~n10767 & ~n10769;
  assign n10772 = ~n10770 & ~n10771;
  assign n10773 = n10760 & n10772;
  assign n10774 = ~n10760 & ~n10772;
  assign n10775 = ~n10773 & ~n10774;
  assign n10776 = ~n9847 & n9850;
  assign n10777 = ~n9846 & ~n10776;
  assign n10778 = n10775 & ~n10777;
  assign n10779 = ~n10775 & n10777;
  assign n10780 = ~n10778 & ~n10779;
  assign n10781 = n10748 & n10780;
  assign n10782 = ~n10748 & ~n10780;
  assign n10783 = ~n10781 & ~n10782;
  assign n10784 = ~n9935 & n9938;
  assign n10785 = ~n9934 & ~n10784;
  assign n10786 = n10783 & n10785;
  assign n10787 = ~n10783 & ~n10785;
  assign n10788 = ~n10786 & ~n10787;
  assign n10789 = ~n10716 & ~n10788;
  assign n10790 = n10716 & n10788;
  assign n10791 = ~n10789 & ~n10790;
  assign n10792 = ~n10111 & n10114;
  assign n10793 = ~n10110 & ~n10792;
  assign n10794 = n10791 & ~n10793;
  assign n10795 = ~n10791 & n10793;
  assign n10796 = ~n10794 & ~n10795;
  assign n10797 = n10644 & n10796;
  assign n10798 = ~n10644 & ~n10796;
  assign n10799 = ~n10797 & ~n10798;
  assign n10800 = ~n10468 & n10471;
  assign n10801 = ~n10467 & ~n10800;
  assign n10802 = n10799 & n10801;
  assign n10803 = ~n10799 & ~n10801;
  assign n10804 = ~n10802 & ~n10803;
  assign n10805 = ~n10487 & ~n10804;
  assign n10806 = n10487 & n10804;
  assign n10807 = ~n10805 & ~n10806;
  assign n10808 = ~n10476 & n10479;
  assign n10809 = ~n10475 & ~n10808;
  assign n10810 = n10807 & ~n10809;
  assign n10811 = ~n10807 & n10809;
  assign n10812 = ~n10810 & ~n10811;
  assign n10813 = n10483 & ~n10812;
  assign n10814 = ~n7138 & ~n7139;
  assign n10815 = ~n7181 & n10814;
  assign n10816 = n7181 & ~n10814;
  assign n10817 = ~n10815 & ~n10816;
  assign n10818 = ~n10766 & n10769;
  assign n10819 = ~n10765 & ~n10818;
  assign n10820 = ~n10754 & n10757;
  assign n10821 = ~n10753 & ~n10820;
  assign n10822 = ~n10773 & n10777;
  assign n10823 = ~n10774 & ~n10822;
  assign n10824 = ~n10821 & n10823;
  assign n10825 = n10821 & ~n10823;
  assign n10826 = ~n10824 & ~n10825;
  assign n10827 = n10819 & n10826;
  assign n10828 = ~n10819 & ~n10826;
  assign n10829 = ~n10827 & ~n10828;
  assign n10830 = ~n10734 & n10737;
  assign n10831 = ~n10733 & ~n10830;
  assign n10832 = ~n10722 & n10725;
  assign n10833 = ~n10721 & ~n10832;
  assign n10834 = ~n10741 & n10745;
  assign n10835 = ~n10742 & ~n10834;
  assign n10836 = ~n10833 & n10835;
  assign n10837 = n10833 & ~n10835;
  assign n10838 = ~n10836 & ~n10837;
  assign n10839 = n10831 & n10838;
  assign n10840 = ~n10831 & ~n10838;
  assign n10841 = ~n10839 & ~n10840;
  assign n10842 = ~n10829 & ~n10841;
  assign n10843 = n10829 & n10841;
  assign n10844 = ~n10842 & ~n10843;
  assign n10845 = ~n10781 & n10785;
  assign n10846 = ~n10782 & ~n10845;
  assign n10847 = n10844 & ~n10846;
  assign n10848 = ~n10844 & n10846;
  assign n10849 = ~n10847 & ~n10848;
  assign n10850 = ~n10694 & n10697;
  assign n10851 = ~n10693 & ~n10850;
  assign n10852 = ~n10682 & n10685;
  assign n10853 = ~n10681 & ~n10852;
  assign n10854 = ~n10701 & n10705;
  assign n10855 = ~n10702 & ~n10854;
  assign n10856 = ~n10853 & n10855;
  assign n10857 = n10853 & ~n10855;
  assign n10858 = ~n10856 & ~n10857;
  assign n10859 = n10851 & n10858;
  assign n10860 = ~n10851 & ~n10858;
  assign n10861 = ~n10859 & ~n10860;
  assign n10862 = ~n10662 & n10665;
  assign n10863 = ~n10661 & ~n10862;
  assign n10864 = ~n10650 & n10653;
  assign n10865 = ~n10649 & ~n10864;
  assign n10866 = ~n10669 & n10673;
  assign n10867 = ~n10670 & ~n10866;
  assign n10868 = ~n10865 & n10867;
  assign n10869 = n10865 & ~n10867;
  assign n10870 = ~n10868 & ~n10869;
  assign n10871 = n10863 & n10870;
  assign n10872 = ~n10863 & ~n10870;
  assign n10873 = ~n10871 & ~n10872;
  assign n10874 = ~n10861 & ~n10873;
  assign n10875 = n10861 & n10873;
  assign n10876 = ~n10874 & ~n10875;
  assign n10877 = ~n10709 & n10713;
  assign n10878 = ~n10710 & ~n10877;
  assign n10879 = n10876 & ~n10878;
  assign n10880 = ~n10876 & n10878;
  assign n10881 = ~n10879 & ~n10880;
  assign n10882 = ~n10849 & ~n10881;
  assign n10883 = n10849 & n10881;
  assign n10884 = ~n10882 & ~n10883;
  assign n10885 = ~n10790 & ~n10793;
  assign n10886 = ~n10789 & ~n10885;
  assign n10887 = n10884 & n10886;
  assign n10888 = ~n10884 & ~n10886;
  assign n10889 = ~n10887 & ~n10888;
  assign n10890 = ~n10614 & n10617;
  assign n10891 = ~n10613 & ~n10890;
  assign n10892 = ~n10602 & n10605;
  assign n10893 = ~n10601 & ~n10892;
  assign n10894 = ~n10621 & n10625;
  assign n10895 = ~n10622 & ~n10894;
  assign n10896 = ~n10893 & n10895;
  assign n10897 = n10893 & ~n10895;
  assign n10898 = ~n10896 & ~n10897;
  assign n10899 = n10891 & n10898;
  assign n10900 = ~n10891 & ~n10898;
  assign n10901 = ~n10899 & ~n10900;
  assign n10902 = ~n10581 & ~n10586;
  assign n10903 = ~n10568 & ~n10573;
  assign n10904 = ~n10590 & ~n10593;
  assign n10905 = ~n10589 & ~n10904;
  assign n10906 = n10903 & ~n10905;
  assign n10907 = ~n10903 & n10905;
  assign n10908 = ~n10906 & ~n10907;
  assign n10909 = n10902 & n10908;
  assign n10910 = ~n10902 & ~n10908;
  assign n10911 = ~n10909 & ~n10910;
  assign n10912 = ~n10901 & n10911;
  assign n10913 = n10901 & ~n10911;
  assign n10914 = ~n10912 & ~n10913;
  assign n10915 = ~n10629 & n10633;
  assign n10916 = ~n10630 & ~n10915;
  assign n10917 = n10914 & ~n10916;
  assign n10918 = ~n10914 & n10916;
  assign n10919 = ~n10917 & ~n10918;
  assign n10920 = ~n10540 & n10543;
  assign n10921 = ~n10539 & ~n10920;
  assign n10922 = ~n10527 & ~n10532;
  assign n10923 = ~n10547 & n10551;
  assign n10924 = ~n10548 & ~n10923;
  assign n10925 = n10922 & ~n10924;
  assign n10926 = ~n10922 & n10924;
  assign n10927 = ~n10925 & ~n10926;
  assign n10928 = n10921 & n10927;
  assign n10929 = ~n10921 & ~n10927;
  assign n10930 = ~n10928 & ~n10929;
  assign n10931 = ~n10506 & ~n10511;
  assign n10932 = ~n10493 & ~n10498;
  assign n10933 = ~n10515 & ~n10518;
  assign n10934 = ~n10514 & ~n10933;
  assign n10935 = n10932 & ~n10934;
  assign n10936 = ~n10932 & n10934;
  assign n10937 = ~n10935 & ~n10936;
  assign n10938 = n10931 & n10937;
  assign n10939 = ~n10931 & ~n10937;
  assign n10940 = ~n10938 & ~n10939;
  assign n10941 = n10930 & n10940;
  assign n10942 = ~n10930 & ~n10940;
  assign n10943 = ~n10941 & ~n10942;
  assign n10944 = ~n10555 & n10559;
  assign n10945 = ~n10556 & ~n10944;
  assign n10946 = n10943 & ~n10945;
  assign n10947 = ~n10943 & n10945;
  assign n10948 = ~n10946 & ~n10947;
  assign n10949 = ~n10919 & ~n10948;
  assign n10950 = n10919 & n10948;
  assign n10951 = ~n10949 & ~n10950;
  assign n10952 = ~n10638 & ~n10641;
  assign n10953 = ~n10637 & ~n10952;
  assign n10954 = n10951 & n10953;
  assign n10955 = ~n10951 & ~n10953;
  assign n10956 = ~n10954 & ~n10955;
  assign n10957 = ~n10889 & ~n10956;
  assign n10958 = n10889 & n10956;
  assign n10959 = ~n10957 & ~n10958;
  assign n10960 = ~n10797 & n10801;
  assign n10961 = ~n10798 & ~n10960;
  assign n10962 = n10959 & ~n10961;
  assign n10963 = ~n10959 & n10961;
  assign n10964 = ~n10962 & ~n10963;
  assign n10965 = ~n10817 & ~n10964;
  assign n10966 = n10817 & n10964;
  assign n10967 = ~n10965 & ~n10966;
  assign n10968 = ~n10806 & ~n10809;
  assign n10969 = ~n10805 & ~n10968;
  assign n10970 = n10967 & n10969;
  assign n10971 = ~n10967 & ~n10969;
  assign n10972 = ~n10970 & ~n10971;
  assign n10973 = n10813 & n10972;
  assign n10974 = ~n7128 & ~n7129;
  assign n10975 = ~n7183 & n10974;
  assign n10976 = n7183 & ~n10974;
  assign n10977 = ~n10975 & ~n10976;
  assign n10978 = n10922 & n10924;
  assign n10979 = ~n10922 & ~n10924;
  assign n10980 = ~n10921 & ~n10979;
  assign n10981 = ~n10978 & ~n10980;
  assign n10982 = ~n10941 & ~n10945;
  assign n10983 = ~n10942 & ~n10982;
  assign n10984 = n10931 & ~n10936;
  assign n10985 = ~n10935 & ~n10984;
  assign n10986 = n10983 & ~n10985;
  assign n10987 = ~n10983 & n10985;
  assign n10988 = ~n10986 & ~n10987;
  assign n10989 = ~n10981 & ~n10988;
  assign n10990 = n10981 & n10988;
  assign n10991 = ~n10989 & ~n10990;
  assign n10992 = ~n10891 & ~n10897;
  assign n10993 = ~n10896 & ~n10992;
  assign n10994 = ~n10912 & ~n10916;
  assign n10995 = ~n10913 & ~n10994;
  assign n10996 = n10902 & ~n10907;
  assign n10997 = ~n10906 & ~n10996;
  assign n10998 = n10995 & ~n10997;
  assign n10999 = ~n10995 & n10997;
  assign n11000 = ~n10998 & ~n10999;
  assign n11001 = ~n10993 & ~n11000;
  assign n11002 = n10993 & n11000;
  assign n11003 = ~n11001 & ~n11002;
  assign n11004 = ~n10991 & ~n11003;
  assign n11005 = n10991 & n11003;
  assign n11006 = ~n11004 & ~n11005;
  assign n11007 = ~n10950 & ~n10953;
  assign n11008 = ~n10949 & ~n11007;
  assign n11009 = n11006 & ~n11008;
  assign n11010 = ~n11006 & n11008;
  assign n11011 = ~n11009 & ~n11010;
  assign n11012 = ~n10875 & n10878;
  assign n11013 = ~n10874 & ~n11012;
  assign n11014 = ~n10863 & ~n10869;
  assign n11015 = ~n10868 & ~n11014;
  assign n11016 = ~n11013 & n11015;
  assign n11017 = n11013 & ~n11015;
  assign n11018 = ~n11016 & ~n11017;
  assign n11019 = ~n10851 & ~n10857;
  assign n11020 = ~n10856 & ~n11019;
  assign n11021 = n11018 & n11020;
  assign n11022 = ~n11018 & ~n11020;
  assign n11023 = ~n11021 & ~n11022;
  assign n11024 = ~n10843 & n10846;
  assign n11025 = ~n10842 & ~n11024;
  assign n11026 = ~n10831 & ~n10837;
  assign n11027 = ~n10836 & ~n11026;
  assign n11028 = ~n11025 & n11027;
  assign n11029 = n11025 & ~n11027;
  assign n11030 = ~n11028 & ~n11029;
  assign n11031 = ~n10819 & ~n10825;
  assign n11032 = ~n10824 & ~n11031;
  assign n11033 = n11030 & n11032;
  assign n11034 = ~n11030 & ~n11032;
  assign n11035 = ~n11033 & ~n11034;
  assign n11036 = n11023 & n11035;
  assign n11037 = ~n11023 & ~n11035;
  assign n11038 = ~n11036 & ~n11037;
  assign n11039 = ~n10883 & ~n10886;
  assign n11040 = ~n10882 & ~n11039;
  assign n11041 = n11038 & ~n11040;
  assign n11042 = ~n11038 & n11040;
  assign n11043 = ~n11041 & ~n11042;
  assign n11044 = n11011 & n11043;
  assign n11045 = ~n11011 & ~n11043;
  assign n11046 = ~n11044 & ~n11045;
  assign n11047 = ~n10958 & n10961;
  assign n11048 = ~n10957 & ~n11047;
  assign n11049 = n11046 & n11048;
  assign n11050 = ~n11046 & ~n11048;
  assign n11051 = ~n11049 & ~n11050;
  assign n11052 = n10977 & ~n11051;
  assign n11053 = ~n10977 & n11051;
  assign n11054 = ~n11052 & ~n11053;
  assign n11055 = ~n10966 & ~n10969;
  assign n11056 = ~n10965 & ~n11055;
  assign n11057 = n11054 & n11056;
  assign n11058 = ~n11054 & ~n11056;
  assign n11059 = ~n11057 & ~n11058;
  assign n11060 = n10973 & n11059;
  assign n11061 = ~n7118 & ~n7119;
  assign n11062 = n7185 & n11061;
  assign n11063 = ~n7185 & ~n11061;
  assign n11064 = ~n11062 & ~n11063;
  assign n11065 = ~n11025 & ~n11027;
  assign n11066 = n11025 & n11027;
  assign n11067 = ~n11032 & ~n11066;
  assign n11068 = ~n11065 & ~n11067;
  assign n11069 = ~n11013 & ~n11015;
  assign n11070 = n11013 & n11015;
  assign n11071 = ~n11020 & ~n11070;
  assign n11072 = ~n11069 & ~n11071;
  assign n11073 = ~n11036 & n11040;
  assign n11074 = ~n11037 & ~n11073;
  assign n11075 = ~n11072 & n11074;
  assign n11076 = n11072 & ~n11074;
  assign n11077 = ~n11075 & ~n11076;
  assign n11078 = n11068 & n11077;
  assign n11079 = ~n11068 & ~n11077;
  assign n11080 = ~n11078 & ~n11079;
  assign n11081 = ~n10993 & ~n10999;
  assign n11082 = ~n10998 & ~n11081;
  assign n11083 = ~n11005 & ~n11008;
  assign n11084 = ~n11004 & ~n11083;
  assign n11085 = ~n10981 & ~n10987;
  assign n11086 = ~n10986 & ~n11085;
  assign n11087 = n11084 & ~n11086;
  assign n11088 = ~n11084 & n11086;
  assign n11089 = ~n11087 & ~n11088;
  assign n11090 = n11082 & n11089;
  assign n11091 = ~n11082 & ~n11089;
  assign n11092 = ~n11090 & ~n11091;
  assign n11093 = ~n11080 & n11092;
  assign n11094 = n11080 & ~n11092;
  assign n11095 = ~n11093 & ~n11094;
  assign n11096 = ~n11044 & n11048;
  assign n11097 = ~n11045 & ~n11096;
  assign n11098 = n11095 & ~n11097;
  assign n11099 = ~n11095 & n11097;
  assign n11100 = ~n11098 & ~n11099;
  assign n11101 = ~n11064 & ~n11100;
  assign n11102 = n11064 & n11100;
  assign n11103 = ~n11101 & ~n11102;
  assign n11104 = ~n11052 & n11056;
  assign n11105 = ~n11053 & ~n11104;
  assign n11106 = n11103 & ~n11105;
  assign n11107 = ~n11103 & n11105;
  assign n11108 = ~n11106 & ~n11107;
  assign n11109 = n11060 & n11108;
  assign n11110 = ~n7108 & ~n7109;
  assign n11111 = n7187 & n11110;
  assign n11112 = ~n7187 & ~n11110;
  assign n11113 = ~n11111 & ~n11112;
  assign n11114 = ~n11068 & ~n11076;
  assign n11115 = ~n11075 & ~n11114;
  assign n11116 = ~n11093 & ~n11097;
  assign n11117 = ~n11094 & ~n11116;
  assign n11118 = ~n11084 & ~n11086;
  assign n11119 = n11084 & n11086;
  assign n11120 = ~n11082 & ~n11119;
  assign n11121 = ~n11118 & ~n11120;
  assign n11122 = n11117 & ~n11121;
  assign n11123 = ~n11117 & n11121;
  assign n11124 = ~n11122 & ~n11123;
  assign n11125 = ~n11115 & ~n11124;
  assign n11126 = n11115 & n11124;
  assign n11127 = ~n11125 & ~n11126;
  assign n11128 = ~n11113 & ~n11127;
  assign n11129 = n11113 & n11127;
  assign n11130 = ~n11128 & ~n11129;
  assign n11131 = ~n11102 & n11105;
  assign n11132 = ~n11101 & ~n11131;
  assign n11133 = ~n11130 & n11132;
  assign n11134 = ~n11129 & ~n11132;
  assign n11135 = ~n11128 & n11134;
  assign n11136 = ~n11133 & ~n11135;
  assign n11137 = n11109 & ~n11136;
  assign n11138 = ~n11109 & n11136;
  assign n11139 = ~n10813 & ~n10972;
  assign n11140 = ~n10973 & ~n11139;
  assign n11141 = ~n11128 & ~n11134;
  assign n11142 = ~n7098 & ~n7099;
  assign n11143 = n7189 & ~n11142;
  assign n11144 = ~n7098 & n7190;
  assign n11145 = ~n11143 & ~n11144;
  assign n11146 = ~n11115 & ~n11123;
  assign n11147 = ~n11122 & ~n11146;
  assign n11148 = n11145 & ~n11147;
  assign n11149 = ~n11145 & n11147;
  assign n11150 = ~n11148 & ~n11149;
  assign n11151 = n11141 & n11150;
  assign n11152 = ~n11141 & ~n11150;
  assign n11153 = ~n11151 & ~n11152;
  assign n11154 = ~n10483 & n10812;
  assign n11155 = ~n10813 & ~n11154;
  assign n11156 = ~n8475 & ~n9770;
  assign n11157 = ~n9771 & n11156;
  assign n11158 = ~n10482 & n11157;
  assign n11159 = ~n10483 & ~n11158;
  assign n11160 = n11155 & n11159;
  assign n11161 = ~n11140 & ~n11160;
  assign n11162 = ~n10973 & ~n11059;
  assign n11163 = ~pi1000  & ~n8474;
  assign n11164 = n11156 & n11163;
  assign n11165 = ~n9771 & ~n11164;
  assign n11166 = n10482 & n11165;
  assign n11167 = ~n11155 & ~n11166;
  assign n11168 = n11140 & ~n11167;
  assign n11169 = ~n11161 & n11168;
  assign n11170 = ~n11060 & n11169;
  assign n11171 = ~n11162 & n11170;
  assign n11172 = n11108 & n11171;
  assign n11173 = ~n11137 & n11172;
  assign n11174 = ~n11138 & n11173;
  assign n11175 = n11153 & n11174;
  assign n11176 = n11137 & n11153;
  assign n11177 = n11141 & ~n11148;
  assign n11178 = ~n7191 & ~n11149;
  assign n11179 = ~n11177 & n11178;
  assign n11180 = ~n11176 & n11179;
  assign po0 = n11175 | ~n11180;
endmodule
