module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251,
    n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307,
    n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391,
    n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426,
    n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475,
    n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710;
  assign n91 = 1'b1;
  assign n92 = ~pi9  & ~pi10 ;
  assign n93 = pi11  & ~n92;
  assign n94 = ~pi12  & ~pi13 ;
  assign n95 = ~pi12  & ~n93;
  assign n96 = ~pi13  & n95;
  assign n97 = ~n93 & n94;
  assign n98 = pi14  & ~n675;
  assign n99 = pi15  & n98;
  assign n100 = ~pi16  & ~n99;
  assign n101 = pi17  & ~n100;
  assign n102 = ~pi18  & ~n101;
  assign n103 = pi19  & pi20 ;
  assign n104 = pi19  & ~n102;
  assign n105 = pi20  & n104;
  assign n106 = ~n102 & n103;
  assign n107 = ~pi21  & ~n676;
  assign n108 = ~pi22  & n107;
  assign n109 = pi23  & ~n108;
  assign n110 = pi24  & pi25 ;
  assign n111 = pi24  & n109;
  assign n112 = pi25  & n111;
  assign n113 = n109 & n110;
  assign n114 = ~pi26  & ~n677;
  assign n115 = pi27  & pi28 ;
  assign n116 = pi28  & pi29 ;
  assign n117 = pi27  & n116;
  assign n118 = pi29  & n115;
  assign n119 = pi27  & ~n114;
  assign n120 = pi28  & n119;
  assign n121 = pi29  & n120;
  assign n122 = ~n114 & n678;
  assign n123 = pi22  & ~n107;
  assign n124 = ~pi14  & ~pi15 ;
  assign n125 = ~pi14  & n675;
  assign n126 = ~pi15  & n125;
  assign n127 = n675 & n124;
  assign n128 = pi16  & ~n680;
  assign n129 = ~pi3  & ~pi4 ;
  assign n130 = ~pi5  & ~pi6 ;
  assign n131 = n129 & n130;
  assign n132 = ~pi18  & pi19 ;
  assign n133 = ~pi1  & ~pi2 ;
  assign n134 = n132 & n133;
  assign n135 = n131 & n134;
  assign n136 = pi11  & ~pi12 ;
  assign n137 = ~pi13  & pi17 ;
  assign n138 = n136 & n137;
  assign n139 = ~pi7  & ~pi8 ;
  assign n140 = pi9  & ~pi10 ;
  assign n141 = pi9  & pi10 ;
  assign n142 = ~n92 & ~n141;
  assign n143 = pi9  & n139;
  assign n144 = n142 & n143;
  assign n145 = n139 & n140;
  assign n146 = n138 & n681;
  assign n147 = pi20  & ~pi21 ;
  assign n148 = n110 & n147;
  assign n149 = pi26  & n110;
  assign n150 = n148 & ~n149;
  assign n151 = n146 & n150;
  assign n152 = n135 & n151;
  assign n153 = ~n128 & n152;
  assign n154 = ~n100 & n153;
  assign n155 = ~n123 & n154;
  assign n156 = pi26  & n677;
  assign n157 = pi18  & n101;
  assign n158 = ~pi17  & n100;
  assign n159 = ~n101 & ~n158;
  assign n160 = n94 & n133;
  assign n161 = n131 & n160;
  assign n162 = ~pi20  & pi21 ;
  assign n163 = ~n147 & ~n162;
  assign n164 = pi11  & pi20 ;
  assign n165 = n110 & n164;
  assign n166 = n681 & n165;
  assign n167 = ~n163 & n166;
  assign n168 = n161 & n167;
  assign n169 = ~n100 & n168;
  assign n170 = ~n128 & n169;
  assign n171 = ~n159 & n170;
  assign n172 = ~n157 & n171;
  assign n173 = n104 & n172;
  assign n174 = ~n123 & n173;
  assign n175 = pi25  & ~n111;
  assign n176 = ~pi25  & n111;
  assign n177 = ~n175 & ~n176;
  assign n178 = pi24  & ~n109;
  assign n179 = ~pi24  & n109;
  assign n180 = ~n178 & ~n179;
  assign n181 = ~pi23  & n108;
  assign n182 = ~n109 & ~n181;
  assign n183 = ~n108 & ~n123;
  assign n184 = pi21  & n676;
  assign n185 = ~n107 & ~n184;
  assign n186 = pi20  & ~n104;
  assign n187 = ~pi20  & n104;
  assign n188 = ~n186 & ~n187;
  assign n189 = ~pi19  & n102;
  assign n190 = ~n104 & ~n189;
  assign n191 = ~n102 & ~n157;
  assign n192 = pi16  & n99;
  assign n193 = ~n100 & ~n192;
  assign n194 = pi15  & ~n98;
  assign n195 = ~pi15  & n98;
  assign n196 = ~n194 & ~n195;
  assign n197 = ~n98 & ~n125;
  assign n198 = pi13  & ~n95;
  assign n199 = ~n675 & ~n198;
  assign n200 = pi12  & n93;
  assign n201 = ~n95 & ~n200;
  assign n202 = ~pi11  & n92;
  assign n203 = ~n93 & ~n202;
  assign n204 = ~pi3  & n133;
  assign n205 = ~pi4  & n204;
  assign n206 = ~pi5  & n205;
  assign n207 = ~pi6  & n206;
  assign n208 = n131 & n133;
  assign n209 = n681 & n682;
  assign n210 = ~n203 & n209;
  assign n211 = n201 & n210;
  assign n212 = n199 & n211;
  assign n213 = ~n197 & n212;
  assign n214 = n196 & n213;
  assign n215 = n193 & n214;
  assign n216 = ~n159 & n215;
  assign n217 = n191 & n216;
  assign n218 = ~n190 & n217;
  assign n219 = n188 & n218;
  assign n220 = n185 & n219;
  assign n221 = n183 & n220;
  assign n222 = ~n182 & n221;
  assign n223 = n180 & n222;
  assign n224 = n177 & n223;
  assign n225 = n109 & n174;
  assign n226 = ~n156 & n683;
  assign n227 = ~n114 & ~n156;
  assign n228 = n683 & n227;
  assign n229 = n109 & n155;
  assign n230 = ~pi27  & n114;
  assign n231 = ~n119 & ~n230;
  assign n232 = n684 & ~n231;
  assign n233 = n679 & ~n232;
  assign n234 = pi28  & ~n119;
  assign n235 = ~pi28  & n119;
  assign n236 = ~n234 & ~n235;
  assign n237 = ~pi7  & n682;
  assign n238 = ~pi8  & n237;
  assign n239 = n142 & n238;
  assign n240 = ~n203 & n239;
  assign n241 = n201 & n240;
  assign n242 = n199 & n241;
  assign n243 = ~n197 & n242;
  assign n244 = n196 & n243;
  assign n245 = n193 & n244;
  assign n246 = ~n159 & n245;
  assign n247 = n191 & n246;
  assign n248 = ~n190 & n247;
  assign n249 = n188 & n248;
  assign n250 = n185 & n249;
  assign n251 = n183 & n250;
  assign n252 = ~n182 & n251;
  assign n253 = n180 & n252;
  assign n254 = n177 & n253;
  assign n255 = n227 & n254;
  assign n256 = ~n231 & n255;
  assign n257 = n236 & n256;
  assign n258 = pi9  & n257;
  assign n259 = n232 & n236;
  assign n260 = n679 & ~n686;
  assign n261 = n679 & ~n684;
  assign n262 = ~pi39  & ~pi40 ;
  assign n263 = pi41  & ~n262;
  assign n264 = ~pi42  & ~n263;
  assign n265 = ~pi43  & n264;
  assign n266 = pi44  & ~n265;
  assign n267 = pi45  & n266;
  assign n268 = ~pi46  & ~n267;
  assign n269 = pi47  & ~n268;
  assign n270 = ~pi48  & ~n269;
  assign n271 = pi49  & ~n270;
  assign n272 = pi50  & n271;
  assign n273 = ~pi51  & ~n272;
  assign n274 = ~pi52  & n273;
  assign n275 = pi53  & ~n274;
  assign n276 = pi54  & n275;
  assign n277 = pi55  & n276;
  assign n278 = pi56  & n277;
  assign n279 = ~pi56  & ~n277;
  assign n280 = pi57  & n279;
  assign n281 = ~n278 & ~n280;
  assign n282 = pi57  & ~n279;
  assign n283 = ~pi55  & ~n276;
  assign n284 = pi55  & ~n276;
  assign n285 = ~pi55  & n276;
  assign n286 = ~n284 & ~n285;
  assign n287 = ~n277 & ~n283;
  assign n288 = ~pi54  & ~n275;
  assign n289 = pi54  & ~n275;
  assign n290 = ~pi54  & n275;
  assign n291 = ~n289 & ~n290;
  assign n292 = ~n276 & ~n288;
  assign n293 = ~pi50  & ~n271;
  assign n294 = pi47  & ~n266;
  assign n295 = ~pi47  & n266;
  assign n296 = ~n294 & ~n295;
  assign n297 = pi30  & pi31 ;
  assign n298 = n262 & n297;
  assign n299 = ~pi52  & pi53 ;
  assign n300 = pi58  & pi59 ;
  assign n301 = n299 & n300;
  assign n302 = n298 & n301;
  assign n303 = pi36  & pi37 ;
  assign n304 = pi38  & ~pi43 ;
  assign n305 = n303 & n304;
  assign n306 = pi32  & pi33 ;
  assign n307 = pi34  & pi35 ;
  assign n308 = n306 & n307;
  assign n309 = n305 & n308;
  assign n310 = pi41  & ~pi42 ;
  assign n311 = pi45  & ~pi46 ;
  assign n312 = n310 & n311;
  assign n313 = pi44  & ~pi48 ;
  assign n314 = pi49  & ~pi51 ;
  assign n315 = n313 & n314;
  assign n316 = n312 & n315;
  assign n317 = n309 & n316;
  assign n318 = n298 & n308;
  assign n319 = ~pi42  & ~pi43 ;
  assign n320 = pi44  & pi45 ;
  assign n321 = n319 & n320;
  assign n322 = pi38  & pi41 ;
  assign n323 = n303 & n322;
  assign n324 = n321 & n323;
  assign n325 = ~pi46  & ~pi48 ;
  assign n326 = n314 & n325;
  assign n327 = n301 & n326;
  assign n328 = n324 & n327;
  assign n329 = n318 & n328;
  assign n330 = n302 & n317;
  assign n331 = ~n296 & n689;
  assign n332 = pi50  & ~n271;
  assign n333 = ~pi50  & n271;
  assign n334 = ~n272 & ~n293;
  assign n335 = ~n332 & ~n333;
  assign n336 = n331 & n690;
  assign n337 = ~pi53  & n274;
  assign n338 = ~n275 & ~n337;
  assign n339 = pi52  & ~n273;
  assign n340 = ~n274 & ~n339;
  assign n341 = pi51  & n272;
  assign n342 = ~n273 & ~n341;
  assign n343 = ~pi49  & n270;
  assign n344 = ~n271 & ~n343;
  assign n345 = pi48  & n269;
  assign n346 = ~n270 & ~n345;
  assign n347 = ~pi47  & n268;
  assign n348 = ~n269 & ~n347;
  assign n349 = pi46  & n267;
  assign n350 = ~n268 & ~n349;
  assign n351 = pi45  & ~n266;
  assign n352 = ~pi45  & n266;
  assign n353 = ~n351 & ~n352;
  assign n354 = ~pi44  & n265;
  assign n355 = ~n266 & ~n354;
  assign n356 = pi43  & ~n264;
  assign n357 = ~n265 & ~n356;
  assign n358 = pi42  & n263;
  assign n359 = ~n264 & ~n358;
  assign n360 = ~pi41  & n262;
  assign n361 = ~n263 & ~n360;
  assign n362 = n298 & n300;
  assign n363 = pi38  & n303;
  assign n364 = n308 & n363;
  assign n365 = n362 & n364;
  assign n366 = n361 & n365;
  assign n367 = ~n359 & n366;
  assign n368 = ~n357 & n367;
  assign n369 = n355 & n368;
  assign n370 = ~n353 & n369;
  assign n371 = ~n350 & n370;
  assign n372 = n348 & n371;
  assign n373 = ~n346 & n372;
  assign n374 = n344 & n373;
  assign n375 = n690 & n374;
  assign n376 = ~n342 & n375;
  assign n377 = ~n340 & n376;
  assign n378 = n338 & n377;
  assign n379 = ~n293 & n331;
  assign n380 = ~n688 & n691;
  assign n381 = ~n687 & n380;
  assign n382 = ~n282 & n381;
  assign n383 = pi39  & pi40 ;
  assign n384 = ~n262 & ~n383;
  assign n385 = ~n278 & ~n279;
  assign n386 = ~pi57  & n279;
  assign n387 = ~n282 & ~n386;
  assign n388 = pi58  & ~n282;
  assign n389 = ~pi58  & n282;
  assign n390 = ~n388 & ~n389;
  assign n391 = pi30  & ~pi39 ;
  assign n392 = pi59  & n391;
  assign n393 = ~n390 & n392;
  assign n394 = n387 & n393;
  assign n395 = ~n385 & n394;
  assign n396 = ~n687 & n395;
  assign n397 = ~n688 & n396;
  assign n398 = n338 & n397;
  assign n399 = ~n340 & n398;
  assign n400 = ~n342 & n399;
  assign n401 = n690 & n400;
  assign n402 = n344 & n401;
  assign n403 = ~n346 & n402;
  assign n404 = n348 & n403;
  assign n405 = ~n350 & n404;
  assign n406 = ~n353 & n405;
  assign n407 = n355 & n406;
  assign n408 = ~n357 & n407;
  assign n409 = ~n359 & n408;
  assign n410 = n361 & n409;
  assign n411 = ~n384 & n410;
  assign n412 = pi38  & n411;
  assign n413 = pi37  & n412;
  assign n414 = pi36  & n413;
  assign n415 = pi35  & n414;
  assign n416 = pi34  & n415;
  assign n417 = pi33  & n416;
  assign n418 = pi32  & n417;
  assign n419 = pi31  & n418;
  assign n420 = n381 & ~n385;
  assign n421 = n387 & n420;
  assign n422 = n303 & n307;
  assign n423 = n297 & n306;
  assign n424 = n422 & n423;
  assign n425 = pi38  & ~pi39 ;
  assign n426 = pi59  & n425;
  assign n427 = ~n384 & n426;
  assign n428 = n424 & n427;
  assign n429 = n361 & n428;
  assign n430 = ~n359 & n429;
  assign n431 = ~n357 & n430;
  assign n432 = n355 & n431;
  assign n433 = ~n353 & n432;
  assign n434 = ~n350 & n433;
  assign n435 = n348 & n434;
  assign n436 = ~n346 & n435;
  assign n437 = n344 & n436;
  assign n438 = n690 & n437;
  assign n439 = ~n342 & n438;
  assign n440 = ~n340 & n439;
  assign n441 = n338 & n440;
  assign n442 = ~n688 & n441;
  assign n443 = ~n687 & n442;
  assign n444 = ~n385 & n443;
  assign n445 = n387 & n444;
  assign n446 = ~n390 & n445;
  assign n447 = ~n281 & n382;
  assign n448 = pi58  & n282;
  assign n449 = pi59  & n448;
  assign n450 = n282 & n300;
  assign n451 = pi51  & ~n293;
  assign n452 = ~pi33  & ~pi34 ;
  assign n453 = ~pi35  & ~pi36 ;
  assign n454 = n452 & n453;
  assign n455 = ~pi31  & ~pi32 ;
  assign n456 = n299 & n455;
  assign n457 = n454 & n456;
  assign n458 = pi47  & ~pi48 ;
  assign n459 = pi49  & n458;
  assign n460 = ~pi37  & ~pi38 ;
  assign n461 = pi39  & ~pi40 ;
  assign n462 = pi39  & n460;
  assign n463 = n384 & n462;
  assign n464 = n460 & n461;
  assign n465 = n459 & n694;
  assign n466 = n312 & n694;
  assign n467 = n459 & n466;
  assign n468 = n312 & n465;
  assign n469 = n457 & n695;
  assign n470 = ~n356 & n469;
  assign n471 = n266 & n470;
  assign n472 = ~n273 & n471;
  assign n473 = ~pi33  & n455;
  assign n474 = ~pi34  & n473;
  assign n475 = ~pi35  & n474;
  assign n476 = ~pi36  & n475;
  assign n477 = n454 & n455;
  assign n478 = n695 & n696;
  assign n479 = ~n356 & n478;
  assign n480 = n694 & n696;
  assign n481 = ~n361 & n480;
  assign n482 = n359 & n481;
  assign n483 = n357 & n482;
  assign n484 = ~n355 & n483;
  assign n485 = n353 & n484;
  assign n486 = n350 & n485;
  assign n487 = ~n348 & n486;
  assign n488 = n346 & n487;
  assign n489 = ~n344 & n488;
  assign n490 = n266 & n479;
  assign n491 = ~n690 & n697;
  assign n492 = ~n273 & n697;
  assign n493 = ~n690 & ~n341;
  assign n494 = n492 & n493;
  assign n495 = n342 & n491;
  assign n496 = n340 & n698;
  assign n497 = ~n338 & n496;
  assign n498 = ~n451 & n472;
  assign n499 = n688 & n699;
  assign n500 = ~n278 & n499;
  assign n501 = n687 & n499;
  assign n502 = n385 & n501;
  assign n503 = n687 & n500;
  assign n504 = ~pi0  & ~pi30 ;
  assign n505 = n700 & n504;
  assign n506 = ~n387 & n700;
  assign n507 = n504 & n506;
  assign n508 = n693 & ~n507;
  assign n509 = n693 & ~n505;
  assign n510 = n693 & ~n504;
  assign n511 = ~pi37  & n696;
  assign n512 = ~pi38  & n511;
  assign n513 = n384 & n512;
  assign n514 = ~n361 & n513;
  assign n515 = n359 & n514;
  assign n516 = n357 & n515;
  assign n517 = ~n355 & n516;
  assign n518 = n353 & n517;
  assign n519 = n350 & n518;
  assign n520 = ~n348 & n519;
  assign n521 = n346 & n520;
  assign n522 = ~n344 & n521;
  assign n523 = ~n690 & n522;
  assign n524 = n342 & n523;
  assign n525 = n340 & n524;
  assign n526 = ~n338 & n525;
  assign n527 = n688 & n526;
  assign n528 = n687 & n527;
  assign n529 = n385 & n528;
  assign n530 = ~n387 & n529;
  assign n531 = n390 & n530;
  assign n532 = pi39  & n531;
  assign n533 = n390 & n506;
  assign n534 = n693 & ~n702;
  assign n535 = ~n692 & ~n534;
  assign n536 = ~n510 & n535;
  assign n537 = ~n692 & ~n510;
  assign n538 = ~n534 & n537;
  assign n539 = ~n692 & ~n701;
  assign n540 = ~pi23  & ~n123;
  assign n541 = pi14  & n675;
  assign n542 = ~n198 & ~n541;
  assign n543 = ~pi12  & pi15 ;
  assign n544 = pi17  & ~pi26 ;
  assign n545 = n543 & n544;
  assign n546 = n678 & n545;
  assign n547 = n148 & n546;
  assign n548 = pi0  & pi1 ;
  assign n549 = n92 & n548;
  assign n550 = n132 & n549;
  assign n551 = pi6  & pi7 ;
  assign n552 = pi8  & pi11 ;
  assign n553 = n551 & n552;
  assign n554 = pi2  & pi3 ;
  assign n555 = pi4  & pi5 ;
  assign n556 = n554 & n555;
  assign n557 = n553 & n556;
  assign n558 = n550 & n557;
  assign n559 = pi17  & ~pi18 ;
  assign n560 = n543 & n559;
  assign n561 = n553 & n560;
  assign n562 = n678 & n561;
  assign n563 = n549 & n556;
  assign n564 = pi19  & ~pi26 ;
  assign n565 = n110 & n564;
  assign n566 = n147 & n565;
  assign n567 = n563 & n566;
  assign n568 = n562 & n567;
  assign n569 = n547 & n558;
  assign n570 = ~n98 & n704;
  assign n571 = n197 & n704;
  assign n572 = ~n199 & n571;
  assign n573 = ~n542 & n570;
  assign n574 = n100 & n705;
  assign n575 = ~n109 & n574;
  assign n576 = ~pi29  & n120;
  assign n577 = pi29  & ~n120;
  assign n578 = ~n576 & ~n577;
  assign n579 = ~pi9  & ~n578;
  assign n580 = ~n236 & n579;
  assign n581 = n231 & n580;
  assign n582 = ~n227 & n581;
  assign n583 = ~n177 & n582;
  assign n584 = ~n180 & n583;
  assign n585 = n182 & n584;
  assign n586 = ~n183 & n585;
  assign n587 = ~n185 & n586;
  assign n588 = ~n188 & n587;
  assign n589 = n190 & n588;
  assign n590 = ~n191 & n589;
  assign n591 = n159 & n590;
  assign n592 = ~n193 & n591;
  assign n593 = ~n196 & n592;
  assign n594 = n197 & n593;
  assign n595 = ~n199 & n594;
  assign n596 = ~n201 & n595;
  assign n597 = n203 & n596;
  assign n598 = ~n142 & n597;
  assign n599 = pi8  & n598;
  assign n600 = pi7  & n599;
  assign n601 = pi6  & n600;
  assign n602 = pi5  & n601;
  assign n603 = pi4  & n602;
  assign n604 = pi3  & n603;
  assign n605 = pi2  & n604;
  assign n606 = pi1  & n605;
  assign n607 = pi0  & n606;
  assign n608 = pi8  & pi29 ;
  assign n609 = n551 & n608;
  assign n610 = n563 & n609;
  assign n611 = n203 & n610;
  assign n612 = ~n201 & n611;
  assign n613 = ~n199 & n612;
  assign n614 = n197 & n613;
  assign n615 = ~n196 & n614;
  assign n616 = ~n193 & n615;
  assign n617 = n159 & n616;
  assign n618 = ~n191 & n617;
  assign n619 = n190 & n618;
  assign n620 = ~n188 & n619;
  assign n621 = ~n185 & n620;
  assign n622 = ~n183 & n621;
  assign n623 = n182 & n622;
  assign n624 = ~n180 & n623;
  assign n625 = ~n177 & n624;
  assign n626 = ~n227 & n625;
  assign n627 = ~pi28  & ~n119;
  assign n628 = n231 & ~n627;
  assign n629 = n626 & n628;
  assign n630 = n548 & n556;
  assign n631 = pi8  & ~pi9 ;
  assign n632 = n551 & n631;
  assign n633 = ~n142 & n632;
  assign n634 = n630 & n633;
  assign n635 = n203 & n634;
  assign n636 = ~n201 & n635;
  assign n637 = ~n199 & n636;
  assign n638 = n197 & n637;
  assign n639 = ~n196 & n638;
  assign n640 = ~n193 & n639;
  assign n641 = n159 & n640;
  assign n642 = ~n191 & n641;
  assign n643 = n190 & n642;
  assign n644 = ~n188 & n643;
  assign n645 = ~n185 & n644;
  assign n646 = ~n183 & n645;
  assign n647 = n182 & n646;
  assign n648 = ~n180 & n647;
  assign n649 = ~n177 & n648;
  assign n650 = ~n227 & n649;
  assign n651 = n231 & n650;
  assign n652 = ~n236 & n651;
  assign n653 = ~n578 & n652;
  assign n654 = ~n540 & n575;
  assign n655 = ~n679 & ~n706;
  assign n656 = pi0  & ~n693;
  assign n657 = ~n655 & ~n656;
  assign n658 = ~n703 & ~n655;
  assign n659 = ~n656 & n658;
  assign n660 = ~n703 & n657;
  assign po1  = ~n685 & ~n707;
  assign n662 = pi0  & pi30 ;
  assign n663 = n282 & ~n662;
  assign n664 = n506 & ~n662;
  assign n665 = n700 & n663;
  assign n666 = ~n685 & ~n655;
  assign n667 = n693 & n666;
  assign n668 = pi0  & n693;
  assign n669 = pi30  & n668;
  assign n670 = n693 & n662;
  assign n671 = ~n534 & ~n709;
  assign n672 = n693 & ~n708;
  assign n673 = n666 & ~n710;
  assign n674 = ~n708 & n667;
  assign n675 = n96 | n97;
  assign n676 = n105 | n106;
  assign n677 = n112 | n113;
  assign n678 = n117 | n118;
  assign n679 = n121 | n122;
  assign n680 = n126 | n127;
  assign n681 = n144 | n145;
  assign n682 = n207 | n208;
  assign n683 = n224 | n225;
  assign n684 = n229 | n226 | n228;
  assign n685 = n261 | n233 | n260;
  assign n686 = n258 | n259;
  assign n687 = n286 | ~n287;
  assign n688 = n291 | ~n292;
  assign n689 = n329 | n330;
  assign n690 = n334 | ~n335;
  assign n691 = n379 | n336 | n378;
  assign n692 = n419 | n421 | n446 | n447;
  assign n693 = n449 | n450;
  assign n694 = n463 | n464;
  assign n695 = n467 | n468;
  assign n696 = n476 | n477;
  assign n697 = n489 | n490;
  assign n698 = n494 | n495;
  assign n699 = n497 | n498;
  assign n700 = n502 | n503;
  assign n701 = n508 | n509;
  assign n702 = n532 | n533;
  assign n703 = n539 | n536 | n538;
  assign n704 = n568 | n569;
  assign n705 = n572 | n573;
  assign n706 = n607 | n629 | n653 | n654;
  assign n707 = n659 | n660;
  assign n708 = n664 | n665;
  assign n709 = n669 | n670;
  assign n710 = n671 | ~n672;
  assign po2  = n673 | n674;
  assign po0  = ~n666;
  assign po3  = ~n91;
  assign po4  = ~n91;
  assign po5  = ~n91;
  assign po6  = ~n91;
  assign po7  = ~n91;
  assign po8  = ~n91;
  assign po9  = ~n91;
  assign po10  = ~n91;
  assign po11  = ~n91;
  assign po12  = ~n91;
  assign po13  = ~n91;
  assign po14  = ~n91;
  assign po15  = ~n91;
  assign po16  = ~n91;
  assign po17  = ~n91;
  assign po18  = ~n91;
  assign po19  = ~n91;
  assign po20  = ~n91;
  assign po21  = ~n91;
  assign po22  = ~n91;
  assign po23  = ~n91;
  assign po24  = ~n91;
  assign po25  = ~n91;
  assign po26  = ~n91;
  assign po27  = ~n91;
  assign po28  = ~n91;
  assign po29  = ~n91;
endmodule
