module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24 ;
  wire n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591,
    n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3626, n3627,
    n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651,
    n3652, n3653, n3654, n3655, n3656, n3657,
    n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681,
    n3682, n3683, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927,
    n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951,
    n3952, n3953, n3954, n3955, n3956, n3957,
    n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987,
    n3988, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4017,
    n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047,
    n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077,
    n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101,
    n4102, n4103, n4104, n4105, n4106, n4107,
    n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131,
    n4132, n4133, n4134, n4135, n4136, n4137,
    n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161,
    n4162, n4163, n4164, n4165, n4166, n4167,
    n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191,
    n4192, n4193, n4194, n4195, n4196, n4197,
    n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251,
    n4252, n4253, n4254, n4255, n4256, n4257,
    n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317,
    n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341,
    n4342, n4343, n4344, n4345, n4346, n4347,
    n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4375, n4376, n4377,
    n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395,
    n4396, n4397, n4398, n4399, n4400, n4401,
    n4402, n4403, n4404, n4405, n4406, n4407,
    n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431,
    n4432, n4433, n4434, n4435, n4436, n4437,
    n4438, n4439, n4440, n4441, n4442, n4443,
    n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4455,
    n4456, n4457, n4458, n4459, n4460, n4461,
    n4462, n4463, n4464, n4465, n4466, n4467,
    n4468, n4469, n4470, n4471, n4472, n4473,
    n4474, n4475, n4476, n4477, n4478, n4479,
    n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491,
    n4492, n4493, n4494, n4495, n4496, n4497,
    n4498, n4499, n4500, n4501, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4520, n4521,
    n4522, n4523, n4524, n4525, n4526, n4527,
    n4528, n4529, n4530, n4531, n4532, n4533,
    n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551,
    n4552, n4553, n4554, n4555, n4556, n4557,
    n4558, n4559, n4560, n4561, n4562, n4563,
    n4564, n4565, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581,
    n4582, n4583, n4584, n4585, n4586, n4587,
    n4588, n4589, n4590, n4591, n4592, n4593,
    n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611,
    n4612, n4613, n4614, n4615, n4616, n4617,
    n4618, n4619, n4620, n4621, n4622, n4623,
    n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641,
    n4642, n4643, n4644, n4645, n4646, n4647,
    n4648, n4649, n4650, n4651, n4652, n4653,
    n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671,
    n4672, n4673, n4674, n4675, n4676, n4677,
    n4678, n4679, n4680, n4681, n4682, n4683,
    n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737,
    n4738, n4739, n4740, n4741, n4742, n4743,
    n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4763, n4764, n4765, n4766, n4767,
    n4768, n4769, n4770, n4771, n4772, n4773,
    n4774, n4775, n4776, n4777, n4778, n4779,
    n4780, n4781, n4782, n4783, n4784, n4785,
    n4786, n4787, n4788, n4789, n4790, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797,
    n4798, n4799, n4800, n4801, n4802, n4803,
    n4804, n4805, n4806, n4807, n4808, n4809,
    n4810, n4811, n4812, n4813, n4814, n4815,
    n4816, n4817, n4818, n4819, n4820, n4821,
    n4822, n4823, n4824, n4825, n4826, n4827,
    n4828, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845,
    n4846, n4847, n4848, n4849, n4850, n4851,
    n4852, n4853, n4854, n4855, n4856, n4857,
    n4858, n4859, n4860, n4861, n4862, n4863,
    n4864, n4865, n4866, n4867, n4868, n4869,
    n4870, n4871, n4872, n4873, n4874, n4875,
    n4876, n4877, n4878, n4879, n4880, n4881,
    n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4889, n4890, n4891, n4892, n4893,
    n4894, n4895, n4896, n4897, n4898, n4899,
    n4900, n4901, n4902, n4903, n4904, n4905,
    n4906, n4907, n4908, n4909, n4910, n4911,
    n4912, n4913, n4914, n4915, n4916, n4917,
    n4918, n4919, n4920, n4921, n4922, n4923,
    n4924, n4925, n4926, n4927, n4928, n4929,
    n4930, n4931, n4932, n4933, n4934, n4935,
    n4936, n4937, n4938, n4939, n4940, n4941,
    n4942, n4943, n4944, n4945, n4946, n4947,
    n4948, n4949, n4950, n4951, n4952, n4953,
    n4954, n4955, n4956, n4957, n4958, n4959,
    n4960, n4961, n4962, n4963, n4964, n4965,
    n4966, n4967, n4968, n4969, n4970, n4971,
    n4972, n4973, n4974, n4975, n4976, n4977,
    n4978, n4979, n4980, n4981, n4982, n4983,
    n4984, n4985, n4986, n4987, n4988, n4989,
    n4990, n4991, n4992, n4993, n4994, n4995,
    n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5004, n5005, n5006, n5007,
    n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019,
    n5020, n5021, n5022, n5023, n5024, n5025,
    n5026, n5027, n5028, n5029, n5030, n5031,
    n5032, n5033, n5034, n5035, n5036, n5037,
    n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049,
    n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061,
    n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151,
    n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217,
    n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247,
    n5248, n5249, n5250, n5251, n5252, n5253,
    n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271,
    n5272, n5273, n5274, n5275, n5276, n5277,
    n5278, n5279, n5280, n5281, n5282, n5283,
    n5284, n5285, n5286, n5287, n5288, n5289,
    n5290, n5291, n5292, n5293, n5294, n5295,
    n5296, n5297, n5298, n5299, n5300, n5301,
    n5302, n5303, n5304, n5305, n5306, n5307,
    n5308, n5309, n5310, n5311, n5312, n5313,
    n5314, n5315, n5316, n5317, n5318, n5319,
    n5320, n5321, n5322, n5323, n5324, n5325,
    n5326, n5327, n5328, n5329, n5330, n5331,
    n5332, n5333, n5334, n5335, n5336, n5337,
    n5338, n5339, n5340, n5341, n5342, n5343,
    n5344, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5352, n5353, n5354, n5355,
    n5356, n5357, n5358, n5359, n5360, n5361,
    n5362, n5363, n5364, n5365, n5366, n5367,
    n5368, n5369, n5370, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391,
    n5392, n5393, n5394, n5395, n5396, n5397,
    n5398, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409,
    n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421,
    n5422, n5423, n5424, n5425, n5426, n5427,
    n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451,
    n5452, n5453, n5454, n5455, n5456, n5457,
    n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481,
    n5482, n5483, n5484, n5485, n5486, n5487,
    n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499,
    n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511,
    n5512, n5513, n5514, n5515, n5516, n5517,
    n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541,
    n5542, n5543, n5544, n5545, n5546, n5547,
    n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571,
    n5572, n5573, n5574, n5575, n5576, n5577,
    n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601,
    n5602, n5603, n5604, n5605, n5606, n5607,
    n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619,
    n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631,
    n5632, n5633, n5634, n5635, n5636, n5637,
    n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649,
    n5650, n5651, n5652, n5653, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661,
    n5662, n5663, n5664, n5665, n5666, n5667,
    n5668, n5669, n5670, n5671, n5672, n5673,
    n5674, n5675, n5676, n5677, n5678, n5679,
    n5680, n5681, n5682, n5683, n5684, n5685,
    n5686, n5687, n5688, n5689, n5690, n5691,
    n5692, n5693, n5694, n5695, n5696, n5697,
    n5698, n5699, n5700, n5701, n5702, n5703,
    n5704, n5705, n5706, n5707, n5708, n5709,
    n5710, n5711, n5712, n5713, n5714, n5715,
    n5716, n5717, n5718, n5719, n5720, n5721,
    n5722, n5723, n5724, n5725, n5726, n5727,
    n5728, n5729, n5730, n5731, n5732, n5733,
    n5734, n5735, n5736, n5737, n5738, n5739,
    n5740, n5741, n5742, n5743, n5744, n5745,
    n5746, n5747, n5748, n5749, n5750, n5751,
    n5752, n5753, n5754, n5755, n5756, n5757,
    n5758, n5759, n5760, n5761, n5762, n5763,
    n5764, n5765, n5766, n5767, n5768, n5769,
    n5770, n5771, n5772, n5773, n5774, n5775,
    n5776, n5777, n5778, n5779, n5780, n5781,
    n5782, n5783, n5784, n5785, n5786, n5787,
    n5788, n5789, n5790, n5791, n5792, n5793,
    n5794, n5795, n5796, n5797, n5798, n5799,
    n5800, n5801, n5802, n5803, n5804, n5805,
    n5806, n5807, n5808, n5809, n5810, n5811,
    n5812, n5813, n5814, n5815, n5816, n5817,
    n5818, n5819, n5820, n5821, n5822, n5823,
    n5824, n5825, n5826, n5827, n5828, n5829,
    n5830, n5831, n5832, n5833, n5834, n5835,
    n5836, n5837, n5838, n5839, n5840, n5841,
    n5842, n5843, n5844, n5845, n5846, n5847,
    n5848, n5849, n5850, n5851, n5852, n5853,
    n5854, n5855, n5856, n5857, n5858, n5859,
    n5860, n5861, n5862, n5863, n5864, n5865,
    n5866, n5867, n5868, n5869, n5870, n5871,
    n5872, n5873, n5874, n5875, n5876, n5877,
    n5878, n5879, n5880, n5881, n5882, n5883,
    n5884, n5885, n5886, n5887, n5888, n5889,
    n5890, n5891, n5892, n5893, n5894, n5895,
    n5896, n5897, n5898, n5899, n5900, n5901,
    n5902, n5903, n5904, n5905, n5906, n5907,
    n5908, n5909, n5910, n5911, n5912, n5913,
    n5914, n5915, n5916, n5917, n5918, n5919,
    n5920, n5921, n5922, n5923, n5924, n5925,
    n5926, n5927, n5928, n5929, n5930, n5931,
    n5932, n5933, n5934, n5935, n5936, n5937,
    n5938, n5939, n5940, n5941, n5942, n5943,
    n5944, n5945, n5946, n5947, n5948, n5949,
    n5950, n5951, n5952, n5953, n5954, n5955,
    n5956, n5957, n5958, n5959, n5960, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967,
    n5968, n5969, n5970, n5971, n5972, n5973,
    n5974, n5975, n5976, n5977, n5978, n5979,
    n5980, n5981, n5982, n5983, n5984, n5985,
    n5986, n5987, n5988, n5989, n5990, n5991,
    n5992, n5993, n5994, n5995, n5996, n5997,
    n5998, n5999, n6000, n6001, n6002, n6003,
    n6004, n6005, n6006, n6007, n6008, n6009,
    n6010, n6011, n6012, n6013, n6014, n6015,
    n6016, n6017, n6018, n6019, n6020, n6021,
    n6022, n6023, n6024, n6025, n6026, n6027,
    n6028, n6029, n6030, n6031, n6032, n6033,
    n6034, n6035, n6036, n6037, n6038, n6039,
    n6040, n6041, n6042, n6043, n6044, n6045,
    n6046, n6047, n6048, n6049, n6050, n6051,
    n6052, n6053, n6054, n6055, n6056, n6057,
    n6058, n6059, n6060, n6061, n6062, n6063,
    n6064, n6065, n6066, n6067, n6068, n6069,
    n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6077, n6078, n6079, n6080, n6081,
    n6082, n6083, n6084, n6085, n6086, n6087,
    n6088, n6089, n6090, n6091, n6092, n6093,
    n6094, n6095, n6096, n6097, n6098, n6099,
    n6100, n6101, n6102, n6103, n6104, n6105,
    n6106, n6107, n6108, n6109, n6110, n6111,
    n6112, n6113, n6114, n6115, n6116, n6117,
    n6118, n6119, n6120, n6121, n6122, n6123,
    n6124, n6125, n6126, n6127, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6139, n6140, n6141,
    n6142, n6143, n6144, n6145, n6146, n6147,
    n6148, n6149, n6150, n6151, n6152, n6153,
    n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165,
    n6166, n6167, n6168, n6169, n6170, n6171,
    n6172, n6173, n6174, n6175, n6176, n6177,
    n6178, n6179, n6180, n6181, n6182, n6183,
    n6184, n6185, n6186, n6187, n6188, n6189,
    n6190, n6191, n6192, n6193, n6194, n6195,
    n6196, n6197, n6198, n6199, n6200, n6201,
    n6202, n6203, n6204, n6205, n6206, n6207,
    n6208, n6209, n6210, n6211, n6212, n6213,
    n6214, n6215, n6216, n6217, n6218, n6219,
    n6220, n6221, n6222, n6223, n6224, n6225,
    n6226, n6227, n6228, n6229, n6230, n6231,
    n6232, n6233, n6234, n6235, n6236, n6237,
    n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255,
    n6256, n6257, n6258, n6259, n6260, n6261,
    n6262, n6263, n6264, n6265, n6266, n6267,
    n6268, n6269, n6270, n6271, n6272, n6273,
    n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285,
    n6286, n6287, n6288, n6289, n6290, n6291,
    n6292, n6293, n6294, n6295, n6296, n6297,
    n6298, n6299, n6300, n6301, n6302, n6303,
    n6304, n6305, n6306, n6307, n6308, n6309,
    n6310, n6311, n6312, n6313, n6314, n6315,
    n6316, n6317, n6318, n6319, n6320, n6321,
    n6322, n6323, n6324, n6325, n6326, n6327,
    n6328, n6329, n6330, n6331, n6332, n6333,
    n6334, n6335, n6336, n6337, n6338, n6339,
    n6340, n6341, n6342, n6343, n6344, n6345,
    n6346, n6347, n6348, n6349, n6350, n6351,
    n6352, n6353, n6354, n6355, n6356, n6357,
    n6358, n6359, n6360, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369,
    n6370, n6371, n6372, n6373, n6374, n6375,
    n6376, n6377, n6378, n6379, n6380, n6381,
    n6382, n6383, n6384, n6385, n6386, n6387,
    n6388, n6389, n6390, n6391, n6392, n6393,
    n6394, n6395, n6396, n6397, n6398, n6399,
    n6400, n6401, n6402, n6403, n6404, n6405,
    n6406, n6407, n6408, n6409, n6410, n6411,
    n6412, n6413, n6414, n6415, n6416, n6417,
    n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429,
    n6430, n6431, n6432, n6433, n6434, n6435,
    n6436, n6437, n6438, n6439, n6440, n6441,
    n6442, n6443, n6444, n6445, n6446, n6447,
    n6448, n6449, n6450, n6451, n6452, n6453,
    n6454, n6455, n6456, n6457, n6458, n6459,
    n6460, n6461, n6462, n6463, n6464, n6465,
    n6466, n6467, n6468, n6469, n6470, n6471,
    n6472, n6473, n6474, n6475, n6476, n6477,
    n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6485, n6486, n6487, n6488, n6489,
    n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6500, n6501,
    n6502, n6503, n6504, n6505, n6506, n6507,
    n6508, n6509, n6510, n6511, n6512, n6513,
    n6514, n6515, n6516, n6517, n6518, n6519,
    n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531,
    n6532, n6533, n6534, n6535, n6536, n6537,
    n6538, n6539, n6540, n6541, n6542, n6543,
    n6544, n6545, n6546, n6547, n6548, n6549,
    n6550, n6551, n6552, n6553, n6554, n6555,
    n6556, n6557, n6558, n6559, n6560, n6561,
    n6562, n6563, n6564, n6565, n6566, n6567,
    n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579,
    n6580, n6581, n6582, n6583, n6584, n6585,
    n6586, n6587, n6588, n6589, n6590, n6591,
    n6592, n6593, n6594, n6595, n6596, n6597,
    n6598, n6599, n6600, n6601, n6602, n6603,
    n6604, n6605, n6606, n6607, n6608, n6609,
    n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621,
    n6622, n6623, n6624, n6625, n6626, n6627,
    n6628, n6629, n6630, n6631, n6632, n6633,
    n6634, n6635, n6636, n6637, n6638, n6639,
    n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651,
    n6652, n6653, n6654, n6655, n6656, n6657,
    n6658, n6659, n6660, n6661, n6662, n6663,
    n6664, n6665, n6666, n6667, n6668, n6669,
    n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681,
    n6682, n6683, n6684, n6685, n6686, n6687,
    n6688, n6689, n6690, n6691, n6692, n6693,
    n6694, n6695, n6696, n6697, n6698, n6699,
    n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711,
    n6712, n6713, n6714, n6715, n6716, n6717,
    n6718, n6719, n6720, n6721, n6722, n6723,
    n6724, n6725, n6726, n6727, n6728, n6729,
    n6730, n6731, n6732, n6733, n6734, n6735,
    n6736, n6737, n6738, n6739, n6740, n6741,
    n6742, n6743, n6744, n6745, n6746, n6747,
    n6748, n6749, n6750, n6751, n6752, n6753,
    n6754, n6755, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6767, n6768, n6769, n6770, n6771,
    n6772, n6773, n6774, n6775, n6776, n6777,
    n6778, n6779, n6780, n6781, n6782, n6783,
    n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801,
    n6802, n6803, n6804, n6805, n6806, n6807,
    n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843,
    n6844, n6845, n6846, n6847, n6848, n6849,
    n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861,
    n6862, n6863, n6864, n6865, n6866, n6867,
    n6868, n6869, n6870, n6871, n6872, n6873,
    n6875, n6876, n6877, n6878, n6879, n6880,
    n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892,
    n6893, n6894, n6895, n6896, n6897, n6898,
    n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952,
    n6953, n6954, n6955, n6956, n6957, n6958,
    n6959, n6960, n6961, n6962, n6963, n6964,
    n6965, n6966, n6967, n6968, n6969, n6970,
    n6971, n6972, n6973, n6974, n6975, n6976,
    n6977, n6978, n6979, n6980, n6981, n6982,
    n6983, n6984, n6985, n6986, n6987, n6988,
    n6989, n6990, n6991, n6992, n6993, n6994,
    n6995, n6996, n6997, n6998, n6999, n7000,
    n7001, n7002, n7003, n7004, n7005, n7006,
    n7007, n7008, n7009, n7010, n7011, n7012,
    n7013, n7014, n7015, n7016, n7017, n7018,
    n7019, n7020, n7021, n7022, n7023, n7024,
    n7025, n7026, n7027, n7028, n7029, n7030,
    n7031, n7032, n7033, n7034, n7035, n7036,
    n7037, n7038, n7039, n7040, n7041, n7042,
    n7043, n7044, n7045, n7046, n7047, n7048,
    n7049, n7050, n7051, n7052, n7053, n7054,
    n7055, n7056, n7057, n7058, n7059, n7060,
    n7061, n7062, n7063, n7064, n7065, n7066,
    n7067, n7068, n7069, n7070, n7071, n7072,
    n7073, n7074, n7075, n7076, n7077, n7078,
    n7079, n7080, n7081, n7082, n7083, n7084,
    n7085, n7086, n7087, n7088, n7089, n7090,
    n7091, n7092, n7093, n7094, n7095, n7096,
    n7097, n7098, n7099, n7100, n7101, n7102,
    n7103, n7104, n7105, n7106, n7107, n7108,
    n7109, n7110, n7111, n7112, n7113, n7114,
    n7115, n7116, n7117, n7118, n7119, n7120,
    n7121, n7122, n7123, n7124, n7125, n7126,
    n7127, n7128, n7129, n7130, n7131, n7132,
    n7133, n7134, n7135, n7136, n7137, n7138,
    n7139, n7140, n7141, n7142, n7143, n7144,
    n7145, n7146, n7147, n7148, n7149, n7150,
    n7151, n7152, n7153, n7154, n7155, n7156,
    n7157, n7158, n7159, n7160, n7161, n7162,
    n7163, n7164, n7165, n7166, n7167, n7168,
    n7169, n7170, n7171, n7172, n7173, n7174,
    n7175, n7176, n7177, n7178, n7179, n7180,
    n7181, n7182, n7183, n7184, n7185, n7186,
    n7187, n7188, n7189, n7190, n7191, n7192,
    n7193, n7194, n7195, n7196, n7197, n7198,
    n7199, n7200, n7201, n7202, n7203, n7204,
    n7205, n7206, n7207, n7208, n7209, n7210,
    n7211, n7212, n7213, n7214, n7215, n7216,
    n7217, n7218, n7219, n7220, n7221, n7222,
    n7223, n7224, n7225, n7226, n7227, n7228,
    n7229, n7230, n7231, n7232, n7233, n7234,
    n7235, n7236, n7237, n7238, n7239, n7240,
    n7241, n7242, n7243, n7244, n7245, n7246,
    n7247, n7248, n7249, n7250, n7251, n7252,
    n7253, n7254, n7255, n7256, n7257, n7258,
    n7259, n7260, n7261, n7262, n7263, n7264,
    n7265, n7266, n7267, n7268, n7269, n7270,
    n7271, n7272, n7273, n7274, n7275, n7276,
    n7277, n7278, n7279, n7280, n7281, n7282,
    n7283, n7284, n7285, n7286, n7287, n7288,
    n7289, n7290, n7291, n7292, n7293, n7294,
    n7295, n7296, n7297, n7298, n7299, n7300,
    n7301, n7302, n7303, n7304, n7305, n7306,
    n7307, n7308, n7309, n7310, n7311, n7312,
    n7313, n7314, n7315, n7316, n7317, n7318,
    n7319, n7320, n7321, n7322, n7323, n7324,
    n7325, n7326, n7327, n7328, n7329, n7330,
    n7331, n7332, n7333, n7334, n7335, n7336,
    n7337, n7338, n7339, n7340, n7341, n7342,
    n7343, n7344, n7345, n7346, n7347, n7348,
    n7349, n7350, n7351, n7352, n7353, n7354,
    n7355, n7356, n7357, n7358, n7359, n7360,
    n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7370, n7371, n7372,
    n7373, n7374, n7375, n7376, n7377, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390,
    n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7398, n7399, n7400, n7401, n7402,
    n7403, n7404, n7405, n7406, n7407, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414,
    n7415, n7416, n7417, n7418, n7419, n7420,
    n7421, n7422, n7423, n7424, n7425, n7426,
    n7427, n7428, n7429, n7430, n7431, n7432,
    n7433, n7434, n7435, n7436, n7437, n7438,
    n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7448, n7449, n7450,
    n7451, n7452, n7453, n7454, n7455, n7456,
    n7457, n7458, n7459, n7460, n7461, n7462,
    n7463, n7464, n7465, n7466, n7467, n7468,
    n7469, n7470, n7471, n7472, n7473, n7474,
    n7475, n7476, n7477, n7478, n7479, n7480,
    n7481, n7482, n7483, n7484, n7485, n7486,
    n7487, n7488, n7489, n7490, n7491, n7492,
    n7493, n7494, n7495, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504,
    n7505, n7506, n7507, n7508, n7509, n7510,
    n7511, n7512, n7513, n7514, n7515, n7516,
    n7517, n7518, n7519, n7520, n7521, n7522,
    n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534,
    n7535, n7536, n7537, n7538, n7539, n7540,
    n7541, n7542, n7543, n7544, n7545, n7546,
    n7547, n7548, n7549, n7550, n7551, n7552,
    n7553, n7554, n7555, n7556, n7557, n7558,
    n7559, n7560, n7561, n7562, n7563, n7564,
    n7565, n7566, n7567, n7568, n7569, n7570,
    n7571, n7572, n7573, n7574, n7575, n7576,
    n7577, n7578, n7579, n7580, n7581, n7582,
    n7583, n7584, n7585, n7586, n7587, n7588,
    n7589, n7590, n7591, n7592, n7593, n7594,
    n7595, n7596, n7597, n7598, n7599, n7600,
    n7601, n7602, n7603, n7604, n7605, n7606,
    n7607, n7608, n7609, n7610, n7611, n7612,
    n7613, n7614, n7615, n7616, n7617, n7618,
    n7619, n7620, n7621, n7622, n7623, n7624,
    n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636,
    n7637, n7638, n7639, n7640, n7641, n7642,
    n7643, n7644, n7645, n7646, n7647, n7648,
    n7649, n7650, n7651, n7652, n7653, n7654,
    n7655, n7656, n7657, n7658, n7659, n7660,
    n7661, n7662, n7663, n7664, n7665, n7666,
    n7667, n7668, n7669, n7670, n7671, n7672,
    n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7684,
    n7685, n7686, n7687, n7688, n7689, n7690,
    n7691, n7692, n7693, n7694, n7695, n7696,
    n7697, n7698, n7699, n7700, n7701, n7702,
    n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714,
    n7715, n7716, n7717, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726,
    n7727, n7728, n7729, n7730, n7731, n7732,
    n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744,
    n7745, n7746, n7747, n7748, n7749, n7750,
    n7751, n7752, n7753, n7754, n7755, n7756,
    n7757, n7758, n7759, n7760, n7761, n7762,
    n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7786,
    n7787, n7788, n7789, n7790, n7791, n7792,
    n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7813, n7814, n7815, n7816,
    n7817, n7818, n7819, n7820, n7821, n7822,
    n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062,
    n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8090, n8091, n8092,
    n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104,
    n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116,
    n8117, n8118, n8119, n8120, n8121, n8122,
    n8123, n8124, n8125, n8126, n8127, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134,
    n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146,
    n8147, n8148, n8149, n8150, n8151, n8152,
    n8153, n8154, n8155, n8156, n8157, n8158,
    n8159, n8160, n8161, n8162, n8163, n8164,
    n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176,
    n8177, n8178, n8179, n8180, n8181, n8182,
    n8183, n8184, n8185, n8186, n8187, n8188,
    n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206,
    n8207, n8208, n8209, n8210, n8211, n8212,
    n8213, n8214, n8215, n8216, n8217, n8218,
    n8219, n8220, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236,
    n8237, n8238, n8239, n8240, n8241, n8242,
    n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8272,
    n8273, n8274, n8275, n8276, n8277, n8278,
    n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296,
    n8297, n8298, n8299, n8300, n8301, n8302,
    n8303, n8304, n8305, n8306, n8307, n8308,
    n8309, n8310, n8311, n8312, n8313, n8314,
    n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326,
    n8327, n8328, n8329, n8330, n8331, n8332,
    n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356,
    n8357, n8358, n8359, n8360, n8361, n8362,
    n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8371, n8372, n8373, n8374,
    n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386,
    n8387, n8388, n8389, n8390, n8391, n8392,
    n8393, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404,
    n8405, n8407, n8408, n8409, n8410, n8411,
    n8412, n8413, n8414, n8415, n8416, n8417,
    n8418, n8419, n8420, n8421, n8422, n8423,
    n8424, n8425, n8426, n8427, n8428, n8429,
    n8430, n8431, n8432, n8433, n8434, n8435,
    n8436, n8437, n8438, n8439, n8440, n8441,
    n8442, n8443, n8444, n8445, n8446, n8447,
    n8448, n8449, n8450, n8451, n8452, n8453,
    n8454, n8455, n8456, n8457, n8458, n8459,
    n8460, n8461, n8462, n8463, n8464, n8465,
    n8466, n8467, n8468, n8469, n8470, n8471,
    n8472, n8473, n8474, n8475, n8476, n8477,
    n8478, n8479, n8480, n8481, n8482, n8483,
    n8484, n8485, n8486, n8487, n8488, n8489,
    n8490, n8491, n8492, n8493, n8494, n8495,
    n8496, n8497, n8498, n8499, n8500, n8501,
    n8502, n8503, n8504, n8505, n8506, n8507,
    n8508, n8509, n8510, n8511, n8512, n8513,
    n8514, n8515, n8516, n8517, n8518, n8519,
    n8520, n8521, n8522, n8523, n8524, n8525,
    n8526, n8527, n8528, n8529, n8530, n8531,
    n8532, n8533, n8534, n8535, n8536, n8537,
    n8538, n8539, n8540, n8541, n8542, n8543,
    n8544, n8545, n8546, n8547, n8548, n8549,
    n8550, n8551, n8552, n8553, n8554, n8555,
    n8556, n8557, n8558, n8559, n8560, n8561,
    n8562, n8563, n8564, n8565, n8566, n8567,
    n8568, n8569, n8570, n8571, n8572, n8573,
    n8574, n8575, n8576, n8577, n8578, n8579,
    n8580, n8581, n8582, n8583, n8584, n8585,
    n8586, n8587, n8588, n8589, n8590, n8591,
    n8592, n8593, n8594, n8595, n8596, n8597,
    n8598, n8599, n8600, n8601, n8602, n8603,
    n8604, n8605, n8606, n8607, n8608, n8609,
    n8610, n8611, n8612, n8613, n8614, n8615,
    n8616, n8617, n8619, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658,
    n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8678, n8679, n8680, n8681, n8682,
    n8683, n8684, n8685, n8686, n8687, n8688,
    n8689, n8690, n8691, n8692, n8693, n8694,
    n8695, n8696, n8697, n8698, n8699, n8700,
    n8701, n8702, n8703, n8704, n8705, n8706,
    n8707, n8708, n8709, n8710, n8711, n8712,
    n8713, n8714, n8715, n8716, n8717, n8718,
    n8719, n8720, n8721, n8722, n8723, n8724,
    n8725, n8726, n8727, n8728, n8729, n8730,
    n8731, n8732, n8733, n8734, n8735, n8736,
    n8737, n8738, n8739, n8740, n8741, n8742,
    n8743, n8744, n8745, n8746, n8747, n8748,
    n8749, n8750, n8751, n8752, n8753, n8754,
    n8755, n8756, n8757, n8758, n8759, n8760,
    n8761, n8762, n8763, n8764, n8765, n8766,
    n8767, n8768, n8769, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778,
    n8779, n8780, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796,
    n8797, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826,
    n8827, n8828, n8829, n8830, n8831, n8832,
    n8833, n8834, n8835, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844,
    n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856,
    n8857, n8858, n8859, n8860, n8861, n8862,
    n8863, n8864, n8865, n8866, n8867, n8868,
    n8869, n8870, n8871, n8872, n8873, n8874,
    n8875, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886,
    n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898,
    n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8906, n8907, n8908, n8909, n8910,
    n8911, n8912, n8913, n8914, n8915, n8916,
    n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8924, n8925, n8926, n8927, n8928,
    n8929, n8930, n8931, n8932, n8933, n8934,
    n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8942, n8943, n8944, n8945, n8946,
    n8947, n8948, n8949, n8950, n8951, n8952,
    n8953, n8954, n8955, n8956, n8957, n8958,
    n8959, n8960, n8961, n8962, n8963, n8964,
    n8965, n8966, n8967, n8968, n8969, n8970,
    n8971, n8972, n8973, n8974, n8975, n8976,
    n8977, n8978, n8979, n8980, n8981, n8982,
    n8983, n8984, n8985, n8986, n8987, n8988,
    n8989, n8990, n8991, n8992, n8993, n8994,
    n8995, n8996, n8997, n8998, n8999, n9000,
    n9001, n9002, n9003, n9004, n9005, n9006,
    n9007, n9008, n9009, n9010, n9011, n9012,
    n9013, n9014, n9015, n9016, n9017, n9018,
    n9019, n9020, n9021, n9022, n9023, n9024,
    n9025, n9026, n9027, n9028, n9029, n9030,
    n9031, n9032, n9033, n9034, n9035, n9036,
    n9037, n9038, n9039, n9040, n9041, n9042,
    n9043, n9044, n9045, n9046, n9047, n9048,
    n9049, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060,
    n9061, n9062, n9063, n9064, n9065, n9066,
    n9067, n9068, n9069, n9070, n9071, n9072,
    n9073, n9074, n9075, n9076, n9077, n9078,
    n9079, n9080, n9081, n9082, n9083, n9084,
    n9085, n9086, n9087, n9088, n9089, n9090,
    n9091, n9092, n9093, n9094, n9095, n9096,
    n9097, n9098, n9099, n9100, n9101, n9102,
    n9103, n9104, n9105, n9106, n9107, n9108,
    n9109, n9110, n9111, n9112, n9113, n9114,
    n9115, n9116, n9117, n9118, n9119, n9120,
    n9121, n9122, n9123, n9124, n9125, n9126,
    n9127, n9128, n9129, n9130, n9131, n9132,
    n9133, n9134, n9135, n9136, n9137, n9138,
    n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9148, n9149, n9150,
    n9151, n9152, n9153, n9154, n9155, n9156,
    n9157, n9158, n9159, n9160, n9161, n9162,
    n9163, n9164, n9165, n9166, n9167, n9168,
    n9169, n9170, n9171, n9172, n9173, n9174,
    n9175, n9176, n9177, n9178, n9179, n9180,
    n9181, n9182, n9183, n9184, n9185, n9186,
    n9187, n9188, n9189, n9190, n9191, n9192,
    n9193, n9194, n9195, n9196, n9197, n9198,
    n9199, n9200, n9201, n9202, n9203, n9204,
    n9205, n9206, n9207, n9208, n9209, n9210,
    n9211, n9212, n9213, n9214, n9215, n9216,
    n9217, n9218, n9219, n9220, n9221, n9222,
    n9223, n9224, n9225, n9226, n9227, n9228,
    n9229, n9230, n9231, n9232, n9233, n9234,
    n9235, n9236, n9237, n9238, n9239, n9240,
    n9241, n9242, n9243, n9244, n9245, n9246,
    n9247, n9248, n9249, n9250, n9251, n9252,
    n9253, n9254, n9255, n9256, n9257, n9258,
    n9259, n9260, n9261, n9262, n9263, n9264,
    n9265, n9266, n9267, n9268, n9269, n9270,
    n9271, n9272, n9273, n9274, n9275, n9276,
    n9277, n9278, n9279, n9280, n9281, n9282,
    n9283, n9284, n9285, n9286, n9287, n9288,
    n9289, n9290, n9291, n9292, n9293, n9294,
    n9295, n9296, n9297, n9298, n9299, n9300,
    n9301, n9302, n9303, n9304, n9305, n9306,
    n9307, n9308, n9309, n9310, n9311, n9312,
    n9313, n9314, n9315, n9316, n9317, n9318,
    n9319, n9320, n9321, n9322, n9323, n9324,
    n9325, n9326, n9327, n9328, n9329, n9330,
    n9331, n9332, n9333, n9334, n9335, n9336,
    n9337, n9338, n9339, n9340, n9341, n9342,
    n9343, n9344, n9345, n9346, n9347, n9348,
    n9349, n9350, n9351, n9352, n9353, n9354,
    n9355, n9356, n9357, n9358, n9359, n9360,
    n9361, n9362, n9363, n9364, n9365, n9366,
    n9367, n9368, n9369, n9370, n9371, n9372,
    n9373, n9374, n9375, n9376, n9377, n9378,
    n9379, n9380, n9381, n9382, n9383, n9384,
    n9385, n9386, n9387, n9388, n9389, n9390,
    n9391, n9392, n9393, n9394, n9395, n9396,
    n9397, n9398, n9399, n9400, n9401, n9402,
    n9403, n9404, n9405, n9406, n9407, n9408,
    n9409, n9410, n9411, n9412, n9413, n9414,
    n9415, n9416, n9417, n9418, n9419, n9420,
    n9421, n9422, n9423, n9424, n9425, n9426,
    n9427, n9428, n9429, n9430, n9431, n9432,
    n9433, n9434, n9435, n9436, n9437, n9438,
    n9439, n9440, n9441, n9442, n9443, n9444,
    n9445, n9446, n9447, n9448, n9449, n9450,
    n9451, n9452, n9453, n9454, n9455, n9456,
    n9457, n9458, n9459, n9460, n9461, n9462,
    n9463, n9464, n9465, n9466, n9467, n9468,
    n9469, n9470, n9471, n9472, n9473, n9474,
    n9475, n9476, n9477, n9478, n9479, n9480,
    n9481, n9482, n9483, n9484, n9485, n9486,
    n9487, n9488, n9489, n9490, n9491, n9492,
    n9493, n9494, n9495, n9496, n9497, n9498,
    n9499, n9500, n9501, n9502, n9503, n9504,
    n9505, n9506, n9507, n9508, n9509, n9510,
    n9511, n9512, n9513, n9514, n9515, n9516,
    n9517, n9518, n9519, n9520, n9521, n9522,
    n9523, n9524, n9525, n9526, n9527, n9528,
    n9529, n9530, n9531, n9532, n9533, n9534,
    n9535, n9536, n9537, n9538, n9539, n9540,
    n9541, n9542, n9543, n9544, n9545, n9546,
    n9547, n9548, n9549, n9550, n9551, n9552,
    n9553, n9554, n9555, n9556, n9557, n9558,
    n9559, n9560, n9561, n9562, n9563, n9564,
    n9565, n9566, n9567, n9568, n9569, n9570,
    n9571, n9572, n9573, n9574, n9575, n9576,
    n9577, n9578, n9579, n9580, n9581, n9582,
    n9583, n9584, n9585, n9586, n9587, n9588,
    n9589, n9590, n9591, n9592, n9593, n9594,
    n9595, n9596, n9597, n9598, n9599;
  assign n50 = ~pi0  & ~pi1 ;
  assign n51 = ~pi1  & ~pi2 ;
  assign n52 = ~pi0  & n51;
  assign n53 = ~pi2  & n50;
  assign n54 = ~pi3  & n8619;
  assign n55 = ~pi4  & n54;
  assign n56 = ~pi22  & ~n55;
  assign n57 = ~pi5  & ~n56;
  assign n58 = pi5  & n56;
  assign n59 = pi5  & ~n56;
  assign n60 = ~pi5  & n56;
  assign n61 = ~n59 & ~n60;
  assign n62 = ~n57 & ~n58;
  assign n63 = pi4  & pi22 ;
  assign n64 = pi4  & ~n54;
  assign n65 = n56 & ~n64;
  assign n66 = ~n63 & ~n65;
  assign n67 = n8620 & ~n66;
  assign n68 = ~n8620 & n66;
  assign n69 = n8620 & n66;
  assign n70 = ~n8620 & ~n66;
  assign n71 = ~n69 & ~n70;
  assign n72 = ~n67 & ~n68;
  assign n73 = ~pi22  & ~n8619;
  assign n74 = ~pi3  & ~n73;
  assign n75 = pi3  & n73;
  assign n76 = pi3  & ~n73;
  assign n77 = ~pi3  & n73;
  assign n78 = ~n76 & ~n77;
  assign n79 = ~n74 & ~n75;
  assign n80 = pi2  & pi22 ;
  assign n81 = pi2  & ~n50;
  assign n82 = n73 & ~n81;
  assign n83 = ~n80 & ~n82;
  assign n84 = n8622 & ~n83;
  assign n85 = ~n8622 & n83;
  assign n86 = n8622 & n83;
  assign n87 = ~n8622 & ~n83;
  assign n88 = ~n86 & ~n87;
  assign n89 = ~n84 & ~n85;
  assign n90 = n8621 & n8623;
  assign n91 = ~pi5  & n55;
  assign n92 = ~pi6  & n91;
  assign n93 = ~pi7  & n92;
  assign n94 = ~pi8  & n93;
  assign n95 = ~pi9  & n94;
  assign n96 = ~pi10  & n95;
  assign n97 = ~pi11  & n96;
  assign n98 = ~pi12  & n97;
  assign n99 = ~pi13  & n98;
  assign n100 = ~pi14  & n99;
  assign n101 = ~pi22  & ~n100;
  assign n102 = pi15  & ~n101;
  assign n103 = ~pi15  & n101;
  assign n104 = pi15  & pi22 ;
  assign n105 = ~pi15  & n100;
  assign n106 = ~pi22  & ~n105;
  assign n107 = pi15  & ~n100;
  assign n108 = n106 & ~n107;
  assign n109 = ~n104 & ~n108;
  assign n110 = ~n102 & ~n103;
  assign n111 = pi20  & pi22 ;
  assign n112 = ~pi16  & n105;
  assign n113 = ~pi17  & n112;
  assign n114 = ~pi18  & n113;
  assign n115 = ~pi19  & n114;
  assign n116 = pi20  & ~n115;
  assign n117 = ~pi20  & n115;
  assign n118 = ~pi22  & ~n117;
  assign n119 = ~n116 & ~n117;
  assign n120 = ~pi22  & n119;
  assign n121 = ~n116 & n118;
  assign n122 = ~n111 & ~n8625;
  assign n123 = pi21  & ~n118;
  assign n124 = ~pi21  & ~pi22 ;
  assign n125 = ~n117 & n124;
  assign n126 = pi21  & pi22 ;
  assign n127 = ~pi21  & n117;
  assign n128 = pi21  & ~n117;
  assign n129 = ~pi22  & ~n128;
  assign n130 = ~n127 & ~n128;
  assign n131 = ~pi22  & n130;
  assign n132 = ~n127 & n129;
  assign n133 = ~n126 & ~n8626;
  assign n134 = ~n123 & ~n125;
  assign n135 = n122 & ~n8627;
  assign n136 = ~n8624 & n135;
  assign n137 = ~pi22  & ~n112;
  assign n138 = pi17  & ~n137;
  assign n139 = ~pi17  & n137;
  assign n140 = ~n138 & ~n139;
  assign n141 = pi16  & ~n106;
  assign n142 = ~pi16  & n106;
  assign n143 = ~n141 & ~n142;
  assign n144 = n140 & ~n143;
  assign n145 = pi18  & pi22 ;
  assign n146 = ~pi22  & ~n114;
  assign n147 = pi18  & ~n113;
  assign n148 = n146 & ~n147;
  assign n149 = ~n145 & ~n148;
  assign n150 = ~pi19  & ~n146;
  assign n151 = pi19  & n146;
  assign n152 = pi19  & ~n146;
  assign n153 = ~pi19  & n146;
  assign n154 = ~n152 & ~n153;
  assign n155 = ~n150 & ~n151;
  assign n156 = ~n149 & ~n8628;
  assign n157 = n144 & n156;
  assign n158 = n136 & n157;
  assign n159 = n149 & ~n8628;
  assign n160 = ~n140 & n143;
  assign n161 = n159 & n160;
  assign n162 = ~n122 & ~n8627;
  assign n163 = n8624 & n162;
  assign n164 = n161 & n163;
  assign n165 = ~n8624 & n162;
  assign n166 = n161 & n165;
  assign n167 = ~n164 & ~n166;
  assign n168 = ~n158 & n167;
  assign n169 = n149 & n8628;
  assign n170 = ~n140 & ~n143;
  assign n171 = n169 & n170;
  assign n172 = n162 & n171;
  assign n173 = n163 & n171;
  assign n174 = n8624 & n172;
  assign n175 = n140 & n143;
  assign n176 = n156 & n175;
  assign n177 = n136 & n176;
  assign n178 = ~n8629 & ~n177;
  assign n179 = n159 & n170;
  assign n180 = n162 & n179;
  assign n181 = n163 & n179;
  assign n182 = n8624 & n180;
  assign n183 = n165 & n171;
  assign n184 = ~n8624 & n172;
  assign n185 = ~n8630 & ~n8631;
  assign n186 = n178 & n185;
  assign n187 = ~n164 & ~n8630;
  assign n188 = n178 & n187;
  assign n189 = ~n166 & n188;
  assign n190 = ~n8631 & n189;
  assign n191 = ~n158 & n190;
  assign n192 = ~n158 & ~n8631;
  assign n193 = ~n166 & n192;
  assign n194 = n188 & n193;
  assign n195 = n168 & n186;
  assign n196 = n8624 & n135;
  assign n197 = n157 & n196;
  assign n198 = n176 & n196;
  assign n199 = ~n197 & ~n198;
  assign n200 = n8632 & ~n197;
  assign n201 = ~n198 & n200;
  assign n202 = n8632 & n199;
  assign n203 = n144 & n159;
  assign n204 = n196 & n203;
  assign n205 = ~n149 & n8628;
  assign n206 = n175 & n205;
  assign n207 = n163 & n206;
  assign n208 = ~n204 & ~n207;
  assign n209 = n160 & n205;
  assign n210 = n165 & n209;
  assign n211 = n170 & n205;
  assign n212 = n163 & n211;
  assign n213 = ~n210 & ~n212;
  assign n214 = ~n207 & ~n212;
  assign n215 = ~n210 & n214;
  assign n216 = ~n204 & n215;
  assign n217 = ~n204 & ~n210;
  assign n218 = n214 & n217;
  assign n219 = n208 & n213;
  assign n220 = n165 & n211;
  assign n221 = n159 & n175;
  assign n222 = n196 & n221;
  assign n223 = n136 & n221;
  assign n224 = ~n222 & ~n223;
  assign n225 = ~n220 & ~n222;
  assign n226 = ~n223 & n225;
  assign n227 = ~n220 & n224;
  assign n228 = n136 & n203;
  assign n229 = n165 & n206;
  assign n230 = ~n228 & ~n229;
  assign n231 = n8635 & n230;
  assign n232 = n8634 & n8635;
  assign n233 = ~n229 & n232;
  assign n234 = ~n228 & n233;
  assign n235 = n8634 & n231;
  assign n236 = n162 & n203;
  assign n237 = n165 & n203;
  assign n238 = ~n8624 & n236;
  assign n239 = n156 & n160;
  assign n240 = n163 & n239;
  assign n241 = ~n8637 & ~n240;
  assign n242 = n144 & n169;
  assign n243 = n163 & n242;
  assign n244 = n157 & n163;
  assign n245 = ~n243 & ~n244;
  assign n246 = ~n8637 & ~n243;
  assign n247 = ~n240 & ~n244;
  assign n248 = n246 & n247;
  assign n249 = n241 & n245;
  assign n250 = n156 & n170;
  assign n251 = n136 & n250;
  assign n252 = n169 & n175;
  assign n253 = n163 & n252;
  assign n254 = ~n251 & ~n253;
  assign n255 = n165 & n252;
  assign n256 = n157 & n165;
  assign n257 = ~n255 & ~n256;
  assign n258 = n254 & n257;
  assign n259 = n8638 & n258;
  assign n260 = n8636 & n259;
  assign n261 = n8633 & n254;
  assign n262 = n8636 & n261;
  assign n263 = ~n243 & n262;
  assign n264 = ~n244 & n263;
  assign n265 = ~n240 & n264;
  assign n266 = ~n256 & n265;
  assign n267 = ~n255 & n266;
  assign n268 = ~n8637 & n267;
  assign n269 = n8633 & n260;
  assign n270 = n196 & n211;
  assign n271 = n136 & n209;
  assign n272 = ~n270 & ~n271;
  assign n273 = n144 & n205;
  assign n274 = n162 & n273;
  assign n275 = n163 & n273;
  assign n276 = n8624 & n274;
  assign n277 = n135 & n161;
  assign n278 = ~n8640 & ~n277;
  assign n279 = n165 & n221;
  assign n280 = n136 & n179;
  assign n281 = ~n279 & ~n280;
  assign n282 = ~n277 & ~n280;
  assign n283 = ~n8640 & ~n279;
  assign n284 = n282 & n283;
  assign n285 = n278 & n281;
  assign n286 = n272 & n8641;
  assign n287 = n163 & n209;
  assign n288 = n136 & n211;
  assign n289 = n165 & n273;
  assign n290 = ~n8624 & n274;
  assign n291 = ~n288 & ~n8642;
  assign n292 = ~n287 & n291;
  assign n293 = n163 & n203;
  assign n294 = n8624 & n236;
  assign n295 = n163 & n221;
  assign n296 = n179 & n196;
  assign n297 = ~n295 & ~n296;
  assign n298 = ~n8643 & n297;
  assign n299 = n292 & n298;
  assign n300 = ~n287 & ~n8643;
  assign n301 = n272 & n297;
  assign n302 = n291 & n301;
  assign n303 = n300 & n302;
  assign n304 = ~n8640 & n303;
  assign n305 = ~n279 & n304;
  assign n306 = ~n277 & n305;
  assign n307 = ~n280 & n306;
  assign n308 = n286 & n299;
  assign n309 = n196 & n250;
  assign n310 = n165 & n179;
  assign n311 = ~n8624 & n180;
  assign n312 = ~n309 & ~n8645;
  assign n313 = n163 & n176;
  assign n314 = n165 & n176;
  assign n315 = n135 & n239;
  assign n316 = ~n314 & ~n315;
  assign n317 = ~n313 & ~n315;
  assign n318 = ~n314 & n317;
  assign n319 = ~n313 & n316;
  assign n320 = n136 & n239;
  assign n321 = ~n8624 & n315;
  assign n322 = n196 & n239;
  assign n323 = n8624 & n315;
  assign n324 = ~n8645 & ~n313;
  assign n325 = ~n314 & n324;
  assign n326 = ~n309 & n325;
  assign n327 = ~n8648 & n326;
  assign n328 = ~n8647 & n327;
  assign n329 = n312 & n8646;
  assign n330 = n165 & n239;
  assign n331 = n165 & n242;
  assign n332 = ~n330 & ~n331;
  assign n333 = n160 & n169;
  assign n334 = ~n250 & ~n333;
  assign n335 = n162 & ~n334;
  assign n336 = n332 & ~n335;
  assign n337 = n8649 & n336;
  assign n338 = n8644 & n337;
  assign n339 = n165 & n250;
  assign n340 = n165 & n333;
  assign n341 = n163 & n250;
  assign n342 = n163 & n333;
  assign n343 = n8649 & n332;
  assign n344 = n8639 & n343;
  assign n345 = n8644 & n344;
  assign n346 = ~n342 & n345;
  assign n347 = ~n341 & n346;
  assign n348 = ~n340 & n347;
  assign n349 = ~n339 & n348;
  assign n350 = n8639 & n338;
  assign n351 = ~pi22  & ~n92;
  assign n352 = ~pi7  & ~n351;
  assign n353 = pi7  & n351;
  assign n354 = pi7  & ~n351;
  assign n355 = ~pi7  & n351;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n352 & ~n353;
  assign n358 = ~n8650 & ~n8651;
  assign n359 = n196 & n209;
  assign n360 = ~n122 & n8627;
  assign n361 = n8624 & n360;
  assign n362 = n273 & n361;
  assign n363 = ~n359 & ~n362;
  assign n364 = ~n212 & ~n279;
  assign n365 = n161 & n196;
  assign n366 = n8624 & n277;
  assign n367 = ~n198 & ~n8652;
  assign n368 = n364 & n367;
  assign n369 = ~n359 & n364;
  assign n370 = ~n8652 & n369;
  assign n371 = ~n198 & n370;
  assign n372 = ~n362 & n371;
  assign n373 = n363 & n367;
  assign n374 = n364 & n373;
  assign n375 = n363 & n368;
  assign n376 = ~n8624 & n360;
  assign n377 = n250 & n376;
  assign n378 = n122 & n8627;
  assign n379 = n8624 & n378;
  assign n380 = n157 & n379;
  assign n381 = ~n377 & ~n380;
  assign n382 = n221 & n376;
  assign n383 = ~n8624 & n378;
  assign n384 = n209 & n383;
  assign n385 = ~n382 & ~n384;
  assign n386 = n239 & n361;
  assign n387 = n211 & n379;
  assign n388 = ~n386 & ~n387;
  assign n389 = n385 & n388;
  assign n390 = n381 & n389;
  assign n391 = n273 & n383;
  assign n392 = n196 & n206;
  assign n393 = n206 & n383;
  assign n394 = ~n392 & ~n393;
  assign n395 = ~n391 & ~n392;
  assign n396 = ~n393 & n395;
  assign n397 = ~n391 & n394;
  assign n398 = n203 & n379;
  assign n399 = ~n8629 & ~n222;
  assign n400 = ~n398 & n399;
  assign n401 = n8654 & n400;
  assign n402 = n390 & n401;
  assign n403 = n381 & n8654;
  assign n404 = n8653 & n403;
  assign n405 = n385 & n404;
  assign n406 = ~n8629 & n405;
  assign n407 = ~n222 & n406;
  assign n408 = ~n386 & n407;
  assign n409 = ~n387 & n408;
  assign n410 = ~n398 & n409;
  assign n411 = n8653 & n402;
  assign n412 = n221 & n379;
  assign n413 = ~n295 & ~n412;
  assign n414 = n239 & n383;
  assign n415 = n203 & n361;
  assign n416 = ~n414 & ~n415;
  assign n417 = n209 & n361;
  assign n418 = n242 & n376;
  assign n419 = ~n417 & ~n418;
  assign n420 = n416 & n419;
  assign n421 = ~n295 & ~n418;
  assign n422 = ~n415 & n421;
  assign n423 = ~n417 & n422;
  assign n424 = ~n412 & n423;
  assign n425 = ~n414 & n424;
  assign n426 = ~n412 & ~n417;
  assign n427 = n421 & n426;
  assign n428 = n416 & n427;
  assign n429 = n413 & n420;
  assign n430 = n176 & n376;
  assign n431 = n333 & n376;
  assign n432 = ~n430 & ~n431;
  assign n433 = n239 & n379;
  assign n434 = n333 & n383;
  assign n435 = ~n433 & ~n434;
  assign n436 = n211 & n376;
  assign n437 = ~n8643 & ~n436;
  assign n438 = ~n433 & ~n436;
  assign n439 = ~n8643 & ~n434;
  assign n440 = n438 & n439;
  assign n441 = n435 & n437;
  assign n442 = n432 & n8657;
  assign n443 = n252 & n376;
  assign n444 = n136 & n206;
  assign n445 = n136 & n273;
  assign n446 = ~n444 & ~n445;
  assign n447 = ~n443 & n446;
  assign n448 = n242 & n383;
  assign n449 = ~n280 & ~n448;
  assign n450 = n161 & n361;
  assign n451 = ~n228 & ~n450;
  assign n452 = ~n228 & ~n280;
  assign n453 = ~n450 & n452;
  assign n454 = ~n448 & n453;
  assign n455 = ~n448 & ~n450;
  assign n456 = n452 & n455;
  assign n457 = n449 & n451;
  assign n458 = n447 & n8658;
  assign n459 = n442 & n458;
  assign n460 = n8656 & n447;
  assign n461 = n8658 & n460;
  assign n462 = ~n8643 & n461;
  assign n463 = ~n436 & n462;
  assign n464 = ~n430 & n463;
  assign n465 = ~n431 & n464;
  assign n466 = ~n433 & n465;
  assign n467 = ~n434 & n466;
  assign n468 = n8656 & n459;
  assign n469 = n209 & n376;
  assign n470 = ~n229 & ~n469;
  assign n471 = ~n229 & ~n255;
  assign n472 = ~n469 & n471;
  assign n473 = ~n255 & n470;
  assign n474 = n196 & n242;
  assign n475 = n136 & n333;
  assign n476 = ~n158 & ~n475;
  assign n477 = ~n474 & ~n475;
  assign n478 = ~n158 & n477;
  assign n479 = ~n474 & n476;
  assign n480 = n171 & n383;
  assign n481 = ~n207 & ~n315;
  assign n482 = ~n480 & n481;
  assign n483 = n8661 & n482;
  assign n484 = n8660 & n483;
  assign n485 = ~n8631 & ~n253;
  assign n486 = n176 & n379;
  assign n487 = n157 & n361;
  assign n488 = ~n486 & ~n487;
  assign n489 = n485 & n488;
  assign n490 = n252 & n383;
  assign n491 = ~n243 & ~n490;
  assign n492 = n206 & n361;
  assign n493 = n161 & n379;
  assign n494 = ~n492 & ~n493;
  assign n495 = n491 & n494;
  assign n496 = ~n243 & ~n253;
  assign n497 = ~n8631 & n496;
  assign n498 = ~n492 & n497;
  assign n499 = ~n487 & n498;
  assign n500 = ~n486 & n499;
  assign n501 = ~n493 & n500;
  assign n502 = ~n490 & n501;
  assign n503 = n488 & n494;
  assign n504 = n485 & n491;
  assign n505 = n503 & n504;
  assign n506 = n489 & n495;
  assign n507 = n179 & n378;
  assign n508 = n179 & n379;
  assign n509 = n8624 & n507;
  assign n510 = ~n288 & ~n8663;
  assign n511 = n171 & n361;
  assign n512 = ~n220 & ~n511;
  assign n513 = n250 & n383;
  assign n514 = n179 & n360;
  assign n515 = n179 & n376;
  assign n516 = ~n8624 & n514;
  assign n517 = ~n513 & ~n8664;
  assign n518 = n512 & n517;
  assign n519 = ~n220 & ~n288;
  assign n520 = ~n8664 & n519;
  assign n521 = ~n511 & n520;
  assign n522 = ~n8663 & n521;
  assign n523 = ~n513 & n522;
  assign n524 = ~n220 & ~n513;
  assign n525 = ~n511 & ~n8664;
  assign n526 = n510 & n525;
  assign n527 = n524 & n526;
  assign n528 = n510 & n518;
  assign n529 = n8662 & n8665;
  assign n530 = n484 & n529;
  assign n531 = n8659 & n530;
  assign n532 = n8660 & n8661;
  assign n533 = n8665 & n532;
  assign n534 = n8655 & n533;
  assign n535 = n8659 & n534;
  assign n536 = n8662 & n535;
  assign n537 = ~n207 & n536;
  assign n538 = ~n8648 & n537;
  assign n539 = ~n8647 & n538;
  assign n540 = ~n480 & n539;
  assign n541 = n8655 & n531;
  assign n542 = n221 & n383;
  assign n543 = ~n398 & ~n542;
  assign n544 = n250 & n361;
  assign n545 = n196 & n333;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~n542 & ~n545;
  assign n548 = ~n544 & n547;
  assign n549 = ~n398 & n548;
  assign n550 = n543 & n546;
  assign n551 = ~n240 & ~n313;
  assign n552 = n157 & n376;
  assign n553 = ~n341 & ~n552;
  assign n554 = ~n341 & n551;
  assign n555 = ~n552 & n554;
  assign n556 = ~n313 & ~n341;
  assign n557 = ~n240 & ~n552;
  assign n558 = n556 & n557;
  assign n559 = n551 & n553;
  assign n560 = n203 & n383;
  assign n561 = ~n342 & ~n560;
  assign n562 = ~n210 & n561;
  assign n563 = n8668 & n562;
  assign n564 = n8667 & n562;
  assign n565 = n8668 & n564;
  assign n566 = n8667 & n563;
  assign n567 = ~n207 & ~n243;
  assign n568 = ~n197 & ~n279;
  assign n569 = ~n339 & n568;
  assign n570 = ~n339 & n567;
  assign n571 = ~n279 & n570;
  assign n572 = ~n197 & n571;
  assign n573 = n567 & n569;
  assign n574 = ~n8648 & ~n487;
  assign n575 = ~n256 & ~n443;
  assign n576 = ~n251 & ~n474;
  assign n577 = n575 & n576;
  assign n578 = n574 & n575;
  assign n579 = n576 & n578;
  assign n580 = n574 & n577;
  assign n581 = n8670 & n8671;
  assign n582 = n8668 & n576;
  assign n583 = n8670 & n582;
  assign n584 = n8667 & n583;
  assign n585 = ~n342 & n584;
  assign n586 = ~n256 & n585;
  assign n587 = ~n210 & n586;
  assign n588 = ~n443 & n587;
  assign n589 = n574 & n588;
  assign n590 = ~n560 & n589;
  assign n591 = n8669 & n581;
  assign n592 = ~n295 & ~n314;
  assign n593 = ~n387 & ~n412;
  assign n594 = n592 & n593;
  assign n595 = ~n295 & n8672;
  assign n596 = ~n314 & n595;
  assign n597 = ~n387 & n596;
  assign n598 = ~n412 & n597;
  assign n599 = n8672 & n594;
  assign n600 = n179 & n361;
  assign n601 = n8624 & n514;
  assign n602 = ~n469 & ~n8674;
  assign n603 = ~n296 & n602;
  assign n604 = ~n444 & ~n8663;
  assign n605 = ~n444 & n603;
  assign n606 = ~n8663 & n605;
  assign n607 = n603 & n604;
  assign n608 = n252 & n361;
  assign n609 = ~n414 & ~n608;
  assign n610 = n211 & n383;
  assign n611 = ~n8645 & ~n610;
  assign n612 = n609 & n611;
  assign n613 = n196 & n273;
  assign n614 = ~n359 & ~n613;
  assign n615 = ~n229 & ~n340;
  assign n616 = n614 & n615;
  assign n617 = n609 & n615;
  assign n618 = ~n8645 & n617;
  assign n619 = ~n359 & n618;
  assign n620 = ~n613 & n619;
  assign n621 = ~n610 & n620;
  assign n622 = n611 & n614;
  assign n623 = n617 & n622;
  assign n624 = n612 & n616;
  assign n625 = n250 & n379;
  assign n626 = ~n204 & ~n625;
  assign n627 = ~n204 & ~n415;
  assign n628 = ~n625 & n627;
  assign n629 = ~n415 & n626;
  assign n630 = n300 & n8677;
  assign n631 = n8676 & n630;
  assign n632 = n8675 & n631;
  assign n633 = n135 & n171;
  assign n634 = n136 & n171;
  assign n635 = ~n8624 & n633;
  assign n636 = n203 & n376;
  assign n637 = ~n8678 & ~n636;
  assign n638 = ~n8664 & ~n636;
  assign n639 = ~n8678 & n638;
  assign n640 = ~n8664 & n637;
  assign n641 = n211 & n361;
  assign n642 = n171 & n376;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~n330 & ~n492;
  assign n645 = n367 & n644;
  assign n646 = n643 & n645;
  assign n647 = ~n330 & n8679;
  assign n648 = ~n8652 & n647;
  assign n649 = ~n198 & n648;
  assign n650 = ~n642 & n649;
  assign n651 = ~n492 & n650;
  assign n652 = ~n641 & n651;
  assign n653 = n8679 & n646;
  assign n654 = ~n222 & ~n8647;
  assign n655 = ~n493 & n654;
  assign n656 = n161 & n383;
  assign n657 = ~n513 & ~n656;
  assign n658 = n136 & n252;
  assign n659 = ~n270 & ~n658;
  assign n660 = ~n244 & ~n511;
  assign n661 = n659 & n660;
  assign n662 = n657 & n661;
  assign n663 = n655 & n657;
  assign n664 = ~n244 & n663;
  assign n665 = ~n270 & n664;
  assign n666 = ~n658 & n665;
  assign n667 = ~n511 & n666;
  assign n668 = n655 & n662;
  assign n669 = n8680 & n8681;
  assign n670 = n632 & n669;
  assign n671 = n8673 & n8675;
  assign n672 = n300 & n671;
  assign n673 = n8681 & n672;
  assign n674 = n8680 & n673;
  assign n675 = n8676 & n674;
  assign n676 = ~n204 & n675;
  assign n677 = ~n415 & n676;
  assign n678 = ~n625 & n677;
  assign n679 = n8673 & n670;
  assign n680 = ~n240 & ~n271;
  assign n681 = ~n240 & ~n340;
  assign n682 = ~n271 & n681;
  assign n683 = ~n340 & n680;
  assign n684 = ~n8642 & ~n377;
  assign n685 = ~n288 & ~n309;
  assign n686 = n221 & n361;
  assign n687 = ~n511 & ~n686;
  assign n688 = n685 & n687;
  assign n689 = n684 & n687;
  assign n690 = n685 & n689;
  assign n691 = n684 & n688;
  assign n692 = n8683 & n687;
  assign n693 = n291 & n692;
  assign n694 = ~n309 & n693;
  assign n695 = ~n377 & n694;
  assign n696 = n8683 & n8684;
  assign n697 = n179 & n383;
  assign n698 = ~n8624 & n507;
  assign n699 = ~n244 & ~n8686;
  assign n700 = ~n434 & n699;
  assign n701 = ~n487 & ~n658;
  assign n702 = n388 & n701;
  assign n703 = ~n244 & ~n386;
  assign n704 = n701 & n703;
  assign n705 = ~n387 & n704;
  assign n706 = ~n434 & n705;
  assign n707 = ~n8686 & n706;
  assign n708 = ~n387 & ~n434;
  assign n709 = ~n8686 & n708;
  assign n710 = n704 & n709;
  assign n711 = n700 & n702;
  assign n712 = ~n296 & ~n486;
  assign n713 = ~n8652 & n491;
  assign n714 = ~n243 & n712;
  assign n715 = ~n8652 & n714;
  assign n716 = ~n490 & n715;
  assign n717 = n712 & n713;
  assign n718 = ~n8630 & ~n436;
  assign n719 = ~n341 & ~n418;
  assign n720 = n718 & n719;
  assign n721 = n176 & n361;
  assign n722 = ~n469 & ~n721;
  assign n723 = ~n177 & ~n610;
  assign n724 = n722 & n723;
  assign n725 = ~n177 & ~n341;
  assign n726 = ~n8630 & ~n610;
  assign n727 = n725 & n726;
  assign n728 = ~n418 & ~n436;
  assign n729 = n722 & n728;
  assign n730 = n727 & n729;
  assign n731 = n720 & n724;
  assign n732 = n8688 & n8689;
  assign n733 = n8687 & n8689;
  assign n734 = n8688 & n733;
  assign n735 = n8687 & n732;
  assign n736 = n8688 & n722;
  assign n737 = n8685 & n736;
  assign n738 = n8687 & n737;
  assign n739 = ~n8630 & n738;
  assign n740 = ~n341 & n739;
  assign n741 = ~n177 & n740;
  assign n742 = ~n436 & n741;
  assign n743 = ~n418 & n742;
  assign n744 = ~n610 & n743;
  assign n745 = n8685 & n8690;
  assign n746 = ~n450 & ~n625;
  assign n747 = n171 & n379;
  assign n748 = ~n166 & ~n747;
  assign n749 = ~n166 & ~n450;
  assign n750 = ~n625 & ~n747;
  assign n751 = n749 & n750;
  assign n752 = n746 & n748;
  assign n753 = ~n166 & n8635;
  assign n754 = ~n450 & n753;
  assign n755 = ~n747 & n754;
  assign n756 = ~n625 & n755;
  assign n757 = n8635 & n8692;
  assign n758 = ~n8631 & ~n204;
  assign n759 = ~n8631 & ~n362;
  assign n760 = ~n204 & n759;
  assign n761 = ~n362 & n758;
  assign n762 = ~n256 & ~n415;
  assign n763 = ~n270 & ~n8643;
  assign n764 = n762 & n763;
  assign n765 = n8694 & n764;
  assign n766 = ~n513 & ~n642;
  assign n767 = ~n480 & ~n513;
  assign n768 = ~n642 & n767;
  assign n769 = ~n480 & n766;
  assign n770 = n8667 & n8695;
  assign n771 = n765 & n770;
  assign n772 = n762 & n8695;
  assign n773 = n763 & n772;
  assign n774 = n8693 & n773;
  assign n775 = n8667 & n774;
  assign n776 = ~n8631 & n775;
  assign n777 = ~n204 & n776;
  assign n778 = ~n362 & n777;
  assign n779 = n8693 & n771;
  assign n780 = ~n330 & ~n412;
  assign n781 = ~n229 & ~n330;
  assign n782 = ~n412 & n781;
  assign n783 = ~n229 & ~n412;
  assign n784 = ~n330 & n783;
  assign n785 = ~n229 & n780;
  assign n786 = ~n280 & ~n444;
  assign n787 = ~n210 & ~n280;
  assign n788 = ~n444 & n787;
  assign n789 = ~n210 & n786;
  assign n790 = ~n339 & ~n8674;
  assign n791 = ~n414 & n790;
  assign n792 = n8698 & n791;
  assign n793 = n8697 & n8698;
  assign n794 = n791 & n793;
  assign n795 = n8697 & n792;
  assign n796 = n136 & n161;
  assign n797 = ~n8624 & n277;
  assign n798 = n176 & n383;
  assign n799 = ~n8647 & ~n798;
  assign n800 = ~n8647 & ~n8700;
  assign n801 = ~n798 & n800;
  assign n802 = ~n8700 & n799;
  assign n803 = ~n198 & ~n392;
  assign n804 = ~n255 & ~n448;
  assign n805 = ~n198 & ~n448;
  assign n806 = ~n255 & ~n392;
  assign n807 = n805 & n806;
  assign n808 = n803 & n804;
  assign n809 = ~n198 & n806;
  assign n810 = ~n8700 & n809;
  assign n811 = ~n8647 & n810;
  assign n812 = ~n448 & n811;
  assign n813 = ~n798 & n812;
  assign n814 = n8701 & n8702;
  assign n815 = n252 & n379;
  assign n816 = ~n228 & ~n815;
  assign n817 = n242 & n379;
  assign n818 = ~n251 & ~n817;
  assign n819 = n816 & n818;
  assign n820 = n242 & n361;
  assign n821 = n206 & n376;
  assign n822 = ~n820 & ~n821;
  assign n823 = n333 & n379;
  assign n824 = ~n475 & ~n823;
  assign n825 = n822 & n824;
  assign n826 = n818 & n822;
  assign n827 = n816 & n824;
  assign n828 = n826 & n827;
  assign n829 = n819 & n825;
  assign n830 = n8703 & n8704;
  assign n831 = n8699 & n830;
  assign n832 = n8696 & n831;
  assign n833 = n8698 & n822;
  assign n834 = n8697 & n833;
  assign n835 = n791 & n834;
  assign n836 = n816 & n835;
  assign n837 = n8703 & n836;
  assign n838 = n8696 & n837;
  assign n839 = n8691 & n838;
  assign n840 = ~n475 & n839;
  assign n841 = ~n251 & n840;
  assign n842 = ~n817 & n841;
  assign n843 = ~n823 & n842;
  assign n844 = n8691 & n832;
  assign n845 = ~n8682 & ~n8705;
  assign n846 = ~n8666 & ~n845;
  assign n847 = n358 & ~n846;
  assign n848 = ~n358 & n846;
  assign n849 = ~n847 & ~n848;
  assign n850 = pi8  & pi22 ;
  assign n851 = ~pi22  & ~n94;
  assign n852 = pi8  & ~n93;
  assign n853 = n851 & ~n852;
  assign n854 = ~n850 & ~n853;
  assign n855 = ~n8650 & ~n854;
  assign n856 = n849 & ~n854;
  assign n857 = ~n8650 & n856;
  assign n858 = n849 & n855;
  assign n859 = ~n847 & ~n8706;
  assign n860 = ~n359 & ~n544;
  assign n861 = n196 & n252;
  assign n862 = n860 & ~n861;
  assign n863 = ~n658 & ~n721;
  assign n864 = ~n545 & ~n8678;
  assign n865 = n136 & n242;
  assign n866 = ~n475 & ~n865;
  assign n867 = n864 & n866;
  assign n868 = n863 & n867;
  assign n869 = ~n861 & n864;
  assign n870 = n860 & n863;
  assign n871 = n866 & n870;
  assign n872 = n869 & n871;
  assign n873 = n862 & n868;
  assign n874 = ~n430 & ~n552;
  assign n875 = ~n487 & n874;
  assign n876 = n239 & n376;
  assign n877 = ~n514 & ~n876;
  assign n878 = ~n514 & n875;
  assign n879 = ~n876 & n878;
  assign n880 = n875 & n877;
  assign n881 = n171 & n196;
  assign n882 = n8624 & n633;
  assign n883 = ~n377 & ~n8709;
  assign n884 = n161 & n376;
  assign n885 = ~n386 & ~n474;
  assign n886 = ~n884 & n885;
  assign n887 = ~n474 & ~n8709;
  assign n888 = ~n884 & n887;
  assign n889 = ~n377 & n888;
  assign n890 = ~n386 & n889;
  assign n891 = ~n377 & ~n386;
  assign n892 = n888 & n891;
  assign n893 = n883 & n886;
  assign n894 = n8708 & n8710;
  assign n895 = n860 & n864;
  assign n896 = n866 & n895;
  assign n897 = n8710 & n896;
  assign n898 = n8708 & n897;
  assign n899 = ~n861 & n898;
  assign n900 = ~n658 & n899;
  assign n901 = ~n721 & n900;
  assign n902 = n8707 & n894;
  assign n903 = ~n392 & ~n613;
  assign n904 = n157 & n383;
  assign n905 = ~n798 & ~n904;
  assign n906 = n609 & n905;
  assign n907 = n609 & n903;
  assign n908 = n905 & n907;
  assign n909 = n903 & n906;
  assign n910 = n250 & n378;
  assign n911 = ~n433 & ~n910;
  assign n912 = ~n380 & n911;
  assign n913 = n447 & n912;
  assign n914 = n447 & n905;
  assign n915 = n609 & n914;
  assign n916 = n903 & n915;
  assign n917 = ~n433 & n916;
  assign n918 = ~n625 & n917;
  assign n919 = ~n380 & n918;
  assign n920 = ~n513 & n919;
  assign n921 = n8712 & n913;
  assign n922 = ~n486 & ~n507;
  assign n923 = ~n656 & n922;
  assign n924 = ~n486 & n8713;
  assign n925 = ~n8663 & n924;
  assign n926 = ~n8686 & n925;
  assign n927 = ~n656 & n926;
  assign n928 = n8713 & n923;
  assign n929 = ~n493 & ~n560;
  assign n930 = n543 & n929;
  assign n931 = n8714 & n930;
  assign n932 = ~n542 & n8714;
  assign n933 = n8711 & n932;
  assign n934 = ~n493 & n933;
  assign n935 = ~n398 & n934;
  assign n936 = ~n560 & n935;
  assign n937 = n8711 & n931;
  assign n938 = n273 & n376;
  assign n939 = ~n641 & ~n938;
  assign n940 = ~n417 & ~n641;
  assign n941 = ~n938 & n940;
  assign n942 = ~n417 & n939;
  assign n943 = ~n382 & ~n469;
  assign n944 = ~n636 & n943;
  assign n945 = ~n436 & ~n450;
  assign n946 = ~n415 & ~n686;
  assign n947 = n945 & n946;
  assign n948 = ~n382 & ~n415;
  assign n949 = ~n469 & n948;
  assign n950 = ~n636 & ~n686;
  assign n951 = n945 & n950;
  assign n952 = n949 & n951;
  assign n953 = n944 & n947;
  assign n954 = n8716 & n945;
  assign n955 = ~n469 & n954;
  assign n956 = ~n382 & n955;
  assign n957 = ~n636 & n956;
  assign n958 = ~n686 & n957;
  assign n959 = ~n415 & n958;
  assign n960 = n8716 & n8717;
  assign n961 = n446 & n903;
  assign n962 = n8718 & n961;
  assign n963 = n8711 & n8718;
  assign n964 = n446 & n963;
  assign n965 = n903 & n964;
  assign n966 = n8711 & n962;
  assign n967 = n333 & n361;
  assign n968 = ~n511 & ~n967;
  assign n969 = ~n418 & ~n511;
  assign n970 = ~n967 & n969;
  assign n971 = ~n418 & n968;
  assign n972 = ~n418 & n822;
  assign n973 = ~n967 & n972;
  assign n974 = ~n511 & n973;
  assign n975 = n822 & n8720;
  assign n976 = ~n431 & ~n492;
  assign n977 = ~n642 & n976;
  assign n978 = ~n642 & n8721;
  assign n979 = ~n431 & n978;
  assign n980 = ~n492 & n979;
  assign n981 = n8721 & n977;
  assign n982 = ~n362 & n8722;
  assign n983 = n8719 & n8722;
  assign n984 = ~n362 & n983;
  assign n985 = n8719 & n982;
  assign n986 = ~n8715 & ~n8723;
  assign n987 = n8715 & n8723;
  assign n988 = n8715 & ~n8723;
  assign n989 = ~n8715 & n8723;
  assign n990 = ~n988 & ~n989;
  assign n991 = ~n986 & ~n987;
  assign n992 = n8650 & n8724;
  assign n993 = pi10  & pi22 ;
  assign n994 = ~pi22  & ~n96;
  assign n995 = pi10  & ~n95;
  assign n996 = n994 & ~n995;
  assign n997 = ~n993 & ~n996;
  assign n998 = n992 & n997;
  assign n999 = n987 & ~n997;
  assign n1000 = ~pi11  & ~n994;
  assign n1001 = pi11  & n994;
  assign n1002 = pi11  & ~n994;
  assign n1003 = ~pi11  & n994;
  assign n1004 = ~n1002 & ~n1003;
  assign n1005 = ~n1000 & ~n1001;
  assign n1006 = ~n8650 & ~n8725;
  assign n1007 = n8650 & n8725;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = ~n8724 & n8725;
  assign n1010 = ~n8724 & ~n1008;
  assign n1011 = ~n999 & ~n8726;
  assign n1012 = ~n998 & ~n999;
  assign n1013 = ~n8726 & n1012;
  assign n1014 = ~n998 & n1011;
  assign n1015 = ~n859 & n8727;
  assign n1016 = pi14  & pi22 ;
  assign n1017 = pi14  & ~n99;
  assign n1018 = ~n100 & ~n1017;
  assign n1019 = ~pi22  & n1018;
  assign n1020 = n101 & ~n1017;
  assign n1021 = ~n1016 & ~n8728;
  assign n1022 = ~n382 & ~n544;
  assign n1023 = ~n608 & n1022;
  assign n1024 = ~n613 & ~n8709;
  assign n1025 = ~n198 & ~n552;
  assign n1026 = ~n198 & ~n8709;
  assign n1027 = ~n613 & n1026;
  assign n1028 = ~n552 & n1027;
  assign n1029 = ~n198 & ~n613;
  assign n1030 = ~n552 & ~n8709;
  assign n1031 = n1029 & n1030;
  assign n1032 = n1024 & n1025;
  assign n1033 = ~n177 & ~n747;
  assign n1034 = ~n387 & n1033;
  assign n1035 = n8729 & n1034;
  assign n1036 = n1023 & n1035;
  assign n1037 = ~n295 & ~n377;
  assign n1038 = ~n486 & ~n8678;
  assign n1039 = ~n295 & ~n486;
  assign n1040 = ~n377 & ~n8678;
  assign n1041 = n1039 & n1040;
  assign n1042 = n1037 & n1038;
  assign n1043 = ~n295 & n8698;
  assign n1044 = ~n8678 & n1043;
  assign n1045 = ~n377 & n1044;
  assign n1046 = ~n486 & n1045;
  assign n1047 = n8698 & n8730;
  assign n1048 = ~n445 & ~n450;
  assign n1049 = ~n412 & ~n8700;
  assign n1050 = ~n8648 & ~n8700;
  assign n1051 = ~n412 & n1050;
  assign n1052 = ~n8648 & ~n412;
  assign n1053 = ~n8700 & n1052;
  assign n1054 = ~n8648 & n1049;
  assign n1055 = ~n445 & n8732;
  assign n1056 = ~n450 & n1055;
  assign n1057 = n1048 & n8732;
  assign n1058 = ~n341 & ~n656;
  assign n1059 = ~n821 & n946;
  assign n1060 = ~n341 & ~n821;
  assign n1061 = ~n686 & n1060;
  assign n1062 = ~n415 & n1061;
  assign n1063 = ~n656 & n1062;
  assign n1064 = ~n415 & ~n656;
  assign n1065 = ~n686 & n1064;
  assign n1066 = n1060 & n1065;
  assign n1067 = n1058 & n1059;
  assign n1068 = n8733 & n8734;
  assign n1069 = n8731 & n8734;
  assign n1070 = n8733 & n1069;
  assign n1071 = n8731 & n1068;
  assign n1072 = n1036 & n8735;
  assign n1073 = n209 & n379;
  assign n1074 = ~n434 & ~n1073;
  assign n1075 = ~n274 & ~n625;
  assign n1076 = ~n8640 & n1074;
  assign n1077 = ~n8642 & n1076;
  assign n1078 = ~n625 & n1077;
  assign n1079 = n1074 & n1075;
  assign n1080 = ~n166 & ~n8645;
  assign n1081 = ~n8645 & ~n339;
  assign n1082 = ~n166 & n1081;
  assign n1083 = ~n166 & ~n339;
  assign n1084 = ~n8645 & n1083;
  assign n1085 = ~n339 & n1080;
  assign n1086 = n8695 & n8737;
  assign n1087 = n8695 & n8736;
  assign n1088 = n8737 & n1087;
  assign n1089 = n8736 & n1086;
  assign n1090 = ~n313 & ~n392;
  assign n1091 = ~n296 & ~n314;
  assign n1092 = n1090 & n1091;
  assign n1093 = ~n8663 & ~n636;
  assign n1094 = n575 & n1093;
  assign n1095 = ~n256 & n1090;
  assign n1096 = ~n314 & n1095;
  assign n1097 = ~n296 & n1096;
  assign n1098 = ~n443 & n1097;
  assign n1099 = ~n636 & n1098;
  assign n1100 = ~n8663 & n1099;
  assign n1101 = n575 & n1091;
  assign n1102 = n1090 & n1093;
  assign n1103 = n1101 & n1102;
  assign n1104 = n1092 & n1094;
  assign n1105 = ~n158 & ~n197;
  assign n1106 = n135 & n157;
  assign n1107 = ~n8686 & n8740;
  assign n1108 = ~n240 & ~n359;
  assign n1109 = ~n823 & n1108;
  assign n1110 = n1107 & n1109;
  assign n1111 = n8739 & n1110;
  assign n1112 = n1086 & n1107;
  assign n1113 = n8736 & n1112;
  assign n1114 = n8739 & n1113;
  assign n1115 = ~n240 & n1114;
  assign n1116 = ~n359 & n1115;
  assign n1117 = ~n823 & n1116;
  assign n1118 = n8738 & n1111;
  assign n1119 = ~n330 & ~n610;
  assign n1120 = ~n362 & ~n876;
  assign n1121 = n1119 & n1120;
  assign n1122 = n187 & n1119;
  assign n1123 = n1120 & n1122;
  assign n1124 = n187 & n1120;
  assign n1125 = n1119 & n1124;
  assign n1126 = n187 & n1121;
  assign n1127 = n162 & n211;
  assign n1128 = ~n8637 & ~n1127;
  assign n1129 = ~n8647 & ~n384;
  assign n1130 = n1128 & n1129;
  assign n1131 = n300 & n703;
  assign n1132 = ~n212 & ~n8647;
  assign n1133 = ~n8637 & n1132;
  assign n1134 = ~n220 & ~n384;
  assign n1135 = n300 & n1134;
  assign n1136 = n703 & n1135;
  assign n1137 = n1133 & n1136;
  assign n1138 = n1130 & n1131;
  assign n1139 = n703 & n8742;
  assign n1140 = n300 & n1139;
  assign n1141 = ~n212 & n1140;
  assign n1142 = ~n220 & n1141;
  assign n1143 = ~n8637 & n1142;
  assign n1144 = ~n8647 & n1143;
  assign n1145 = ~n384 & n1144;
  assign n1146 = n8742 & n8743;
  assign n1147 = ~n279 & ~n492;
  assign n1148 = ~n279 & n8744;
  assign n1149 = ~n492 & n1148;
  assign n1150 = n8744 & n1147;
  assign n1151 = n8741 & n8745;
  assign n1152 = n1033 & n8745;
  assign n1153 = n1023 & n1152;
  assign n1154 = n8729 & n1153;
  assign n1155 = n8734 & n1154;
  assign n1156 = n8731 & n1155;
  assign n1157 = n8741 & n1156;
  assign n1158 = n8733 & n1157;
  assign n1159 = ~n387 & n1158;
  assign n1160 = n1072 & n8741;
  assign n1161 = n8745 & n1160;
  assign n1162 = n1072 & n1151;
  assign n1163 = n273 & n379;
  assign n1164 = ~n445 & ~n1163;
  assign n1165 = ~n207 & ~n641;
  assign n1166 = ~n207 & ~n445;
  assign n1167 = ~n641 & ~n1163;
  assign n1168 = n1166 & n1167;
  assign n1169 = n1164 & n1165;
  assign n1170 = n332 & n945;
  assign n1171 = ~n8629 & ~n240;
  assign n1172 = n187 & n1171;
  assign n1173 = n945 & n1171;
  assign n1174 = n187 & n332;
  assign n1175 = n1173 & n1174;
  assign n1176 = n1170 & n1172;
  assign n1177 = n8747 & n8748;
  assign n1178 = n945 & n1174;
  assign n1179 = n8676 & n1178;
  assign n1180 = ~n207 & n1179;
  assign n1181 = ~n8629 & n1180;
  assign n1182 = ~n240 & n1181;
  assign n1183 = ~n445 & n1182;
  assign n1184 = ~n641 & n1183;
  assign n1185 = ~n1163 & n1184;
  assign n1186 = n8676 & n1177;
  assign n1187 = ~n339 & ~n412;
  assign n1188 = ~n339 & n8749;
  assign n1189 = ~n412 & n1188;
  assign n1190 = n8749 & n1187;
  assign n1191 = ~n8652 & ~n511;
  assign n1192 = ~n8647 & ~n433;
  assign n1193 = ~n8631 & ~n197;
  assign n1194 = n1192 & n1193;
  assign n1195 = ~n8631 & ~n511;
  assign n1196 = ~n197 & ~n8652;
  assign n1197 = n1195 & n1196;
  assign n1198 = n1192 & n1197;
  assign n1199 = n1191 & n1194;
  assign n1200 = ~n166 & ~n545;
  assign n1201 = ~n166 & ~n342;
  assign n1202 = ~n545 & n1201;
  assign n1203 = ~n342 & n1200;
  assign n1204 = ~n544 & ~n560;
  assign n1205 = ~n177 & ~n636;
  assign n1206 = ~n544 & n1205;
  assign n1207 = ~n560 & n1206;
  assign n1208 = ~n560 & ~n636;
  assign n1209 = ~n177 & ~n544;
  assign n1210 = n1208 & n1209;
  assign n1211 = n1204 & n1205;
  assign n1212 = n8752 & n8753;
  assign n1213 = ~n8637 & ~n377;
  assign n1214 = ~n8637 & ~n313;
  assign n1215 = ~n377 & n1214;
  assign n1216 = ~n313 & n1213;
  assign n1217 = ~n256 & ~n721;
  assign n1218 = ~n256 & ~n486;
  assign n1219 = ~n721 & n1218;
  assign n1220 = ~n486 & n1217;
  assign n1221 = n8754 & n8755;
  assign n1222 = n8752 & n1221;
  assign n1223 = n8753 & n1222;
  assign n1224 = n1212 & n1221;
  assign n1225 = ~n8631 & n8756;
  assign n1226 = ~n8652 & n1225;
  assign n1227 = ~n197 & n1226;
  assign n1228 = ~n8647 & n1227;
  assign n1229 = ~n511 & n1228;
  assign n1230 = ~n433 & n1229;
  assign n1231 = n8751 & n8756;
  assign n1232 = ~n747 & ~n865;
  assign n1233 = ~n391 & ~n475;
  assign n1234 = n1232 & n1233;
  assign n1235 = ~n493 & ~n817;
  assign n1236 = n1120 & n1235;
  assign n1237 = ~n817 & n1232;
  assign n1238 = ~n493 & n1120;
  assign n1239 = n1233 & n1238;
  assign n1240 = n1237 & n1239;
  assign n1241 = n1120 & n1234;
  assign n1242 = ~n817 & n1241;
  assign n1243 = ~n493 & n1242;
  assign n1244 = n1234 & n1236;
  assign n1245 = ~n430 & n8758;
  assign n1246 = ~n431 & n1245;
  assign n1247 = n432 & n8758;
  assign n1248 = ~n228 & ~n314;
  assign n1249 = ~n8686 & ~n967;
  assign n1250 = n1248 & n1249;
  assign n1251 = ~n158 & ~n204;
  assign n1252 = ~n223 & ~n244;
  assign n1253 = n1251 & n1252;
  assign n1254 = n1250 & n1253;
  assign n1255 = ~n480 & ~n904;
  assign n1256 = ~n480 & n574;
  assign n1257 = ~n904 & n1256;
  assign n1258 = n574 & n1255;
  assign n1259 = ~n443 & ~n821;
  assign n1260 = ~n341 & ~n448;
  assign n1261 = n1259 & n1260;
  assign n1262 = n8760 & n1261;
  assign n1263 = n1248 & n1251;
  assign n1264 = n1060 & n1252;
  assign n1265 = n1263 & n1264;
  assign n1266 = ~n443 & ~n448;
  assign n1267 = n1249 & n1266;
  assign n1268 = n8760 & n1267;
  assign n1269 = n1265 & n1268;
  assign n1270 = n1254 & n1262;
  assign n1271 = n8759 & n8761;
  assign n1272 = n8757 & n8761;
  assign n1273 = n8759 & n1272;
  assign n1274 = n8757 & n1271;
  assign n1275 = n8750 & n8759;
  assign n1276 = n1252 & n1275;
  assign n1277 = n1248 & n1276;
  assign n1278 = n1251 & n1277;
  assign n1279 = n8757 & n1278;
  assign n1280 = n8760 & n1279;
  assign n1281 = ~n443 & n1280;
  assign n1282 = n1060 & n1281;
  assign n1283 = ~n967 & n1282;
  assign n1284 = ~n448 & n1283;
  assign n1285 = ~n8686 & n1284;
  assign n1286 = n8750 & n8762;
  assign n1287 = ~n8666 & ~n8763;
  assign n1288 = n8666 & n8763;
  assign n1289 = n8666 & ~n8763;
  assign n1290 = ~n8666 & n8763;
  assign n1291 = ~n1289 & ~n1290;
  assign n1292 = ~n1287 & ~n1288;
  assign n1293 = ~n8746 & ~n1287;
  assign n1294 = ~n8764 & ~n1293;
  assign n1295 = n8746 & ~n8764;
  assign n1296 = n1021 & n8765;
  assign n1297 = n8746 & ~n1288;
  assign n1298 = ~n8764 & ~n1297;
  assign n1299 = ~n8746 & ~n8764;
  assign n1300 = ~n1021 & n8766;
  assign n1301 = ~n1296 & ~n1300;
  assign n1302 = ~pi22  & ~n98;
  assign n1303 = ~pi13  & ~n1302;
  assign n1304 = pi13  & n1302;
  assign n1305 = pi13  & ~n1302;
  assign n1306 = ~pi13  & n1302;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1303 & ~n1304;
  assign n1309 = n8764 & ~n1293;
  assign n1310 = n8767 & n1309;
  assign n1311 = n8746 & ~n8763;
  assign n1312 = n8764 & ~n1297;
  assign n1313 = n8764 & ~n1311;
  assign n1314 = ~n8767 & n8768;
  assign n1315 = ~n1310 & ~n1314;
  assign n1316 = ~n1296 & n1315;
  assign n1317 = ~n1300 & n1316;
  assign n1318 = ~n1296 & ~n1314;
  assign n1319 = ~n1300 & ~n1310;
  assign n1320 = n1318 & n1319;
  assign n1321 = n1301 & n1315;
  assign n1322 = pi12  & pi22 ;
  assign n1323 = pi12  & ~n97;
  assign n1324 = n1302 & ~n1323;
  assign n1325 = ~n1322 & ~n1324;
  assign n1326 = ~n210 & ~n8637;
  assign n1327 = ~n443 & ~n1073;
  assign n1328 = ~n8637 & ~n443;
  assign n1329 = ~n210 & ~n1073;
  assign n1330 = n1328 & n1329;
  assign n1331 = n1326 & n1327;
  assign n1332 = ~n382 & ~n417;
  assign n1333 = ~n393 & ~n433;
  assign n1334 = n300 & n1333;
  assign n1335 = n1332 & n1334;
  assign n1336 = ~n210 & n1334;
  assign n1337 = ~n8637 & n1336;
  assign n1338 = ~n443 & n1337;
  assign n1339 = ~n382 & n1338;
  assign n1340 = ~n417 & n1339;
  assign n1341 = ~n1073 & n1340;
  assign n1342 = n8770 & n1335;
  assign n1343 = ~n391 & ~n444;
  assign n1344 = ~n798 & ~n8709;
  assign n1345 = n206 & n379;
  assign n1346 = ~n658 & ~n1345;
  assign n1347 = n1344 & n1346;
  assign n1348 = n1343 & n1346;
  assign n1349 = n1344 & n1348;
  assign n1350 = n1343 & n1347;
  assign n1351 = ~n295 & ~n686;
  assign n1352 = ~n243 & ~n295;
  assign n1353 = ~n686 & n1352;
  assign n1354 = ~n243 & n1351;
  assign n1355 = ~n255 & ~n8640;
  assign n1356 = ~n220 & ~n636;
  assign n1357 = ~n220 & n1355;
  assign n1358 = ~n636 & n1357;
  assign n1359 = n1355 & n1356;
  assign n1360 = n8773 & n8774;
  assign n1361 = n8772 & n1360;
  assign n1362 = n8771 & n1361;
  assign n1363 = n8750 & n8774;
  assign n1364 = n1344 & n1363;
  assign n1365 = n8773 & n1364;
  assign n1366 = n8771 & n1365;
  assign n1367 = ~n444 & n1366;
  assign n1368 = ~n658 & n1367;
  assign n1369 = ~n1345 & n1368;
  assign n1370 = ~n391 & n1369;
  assign n1371 = n8750 & n1362;
  assign n1372 = ~n244 & ~n8642;
  assign n1373 = ~n384 & ~n513;
  assign n1374 = n1372 & n1373;
  assign n1375 = n576 & n1374;
  assign n1376 = n576 & n8752;
  assign n1377 = ~n244 & n1376;
  assign n1378 = ~n8642 & n1377;
  assign n1379 = ~n513 & n1378;
  assign n1380 = ~n384 & n1379;
  assign n1381 = n8752 & n1375;
  assign n1382 = ~n8631 & ~n865;
  assign n1383 = ~n8631 & n8776;
  assign n1384 = ~n865 & n1383;
  assign n1385 = n8776 & n1382;
  assign n1386 = ~n314 & ~n469;
  assign n1387 = ~n341 & ~n475;
  assign n1388 = ~n469 & ~n475;
  assign n1389 = ~n314 & ~n341;
  assign n1390 = n1388 & n1389;
  assign n1391 = n1386 & n1387;
  assign n1392 = ~n253 & ~n309;
  assign n1393 = n762 & n1392;
  assign n1394 = ~n341 & n1393;
  assign n1395 = ~n314 & n1394;
  assign n1396 = ~n475 & n1395;
  assign n1397 = ~n469 & n1396;
  assign n1398 = n8778 & n1393;
  assign n1399 = n364 & ~n904;
  assign n1400 = ~n387 & ~n625;
  assign n1401 = n1090 & n1400;
  assign n1402 = ~n8678 & ~n938;
  assign n1403 = ~n380 & ~n861;
  assign n1404 = n1402 & n1403;
  assign n1405 = n1401 & n1404;
  assign n1406 = n1399 & n1405;
  assign n1407 = n8779 & n1406;
  assign n1408 = n8777 & n1407;
  assign n1409 = n1090 & n8777;
  assign n1410 = n1399 & n1409;
  assign n1411 = n1403 & n1410;
  assign n1412 = n8779 & n1411;
  assign n1413 = n8775 & n1412;
  assign n1414 = n1402 & n1413;
  assign n1415 = ~n387 & n1414;
  assign n1416 = ~n625 & n1415;
  assign n1417 = n8775 & n1408;
  assign n1418 = ~n8746 & ~n8780;
  assign n1419 = n8746 & n8780;
  assign n1420 = n8746 & ~n8780;
  assign n1421 = ~n8746 & n8780;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = ~n1418 & ~n1419;
  assign n1424 = n8715 & ~n1419;
  assign n1425 = ~n8781 & ~n1424;
  assign n1426 = ~n8715 & ~n8781;
  assign n1427 = ~n1325 & n8782;
  assign n1428 = ~n8715 & ~n1418;
  assign n1429 = ~n8781 & ~n1428;
  assign n1430 = n8715 & ~n8781;
  assign n1431 = n1325 & n8783;
  assign n1432 = ~n1427 & ~n1431;
  assign n1433 = n8781 & ~n1428;
  assign n1434 = n8725 & n1433;
  assign n1435 = n8715 & ~n8780;
  assign n1436 = n8781 & ~n1424;
  assign n1437 = n8781 & ~n1435;
  assign n1438 = ~n8725 & n8784;
  assign n1439 = ~n1434 & ~n1438;
  assign n1440 = ~n1431 & n1439;
  assign n1441 = ~n1427 & n1440;
  assign n1442 = n1432 & n1439;
  assign n1443 = n8769 & n8785;
  assign n1444 = ~n8769 & ~n8785;
  assign n1445 = n8769 & ~n8785;
  assign n1446 = ~n8769 & n8785;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~n1443 & ~n1444;
  assign n1449 = ~pi9  & ~n851;
  assign n1450 = pi9  & n851;
  assign n1451 = pi9  & ~n851;
  assign n1452 = ~pi9  & n851;
  assign n1453 = ~n1451 & ~n1452;
  assign n1454 = ~n1449 & ~n1450;
  assign n1455 = n992 & n8787;
  assign n1456 = n987 & ~n8787;
  assign n1457 = ~n8650 & ~n997;
  assign n1458 = n8650 & n997;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = ~n8724 & n997;
  assign n1461 = ~n8724 & ~n1459;
  assign n1462 = ~n1456 & ~n8788;
  assign n1463 = ~n1455 & ~n1456;
  assign n1464 = ~n8788 & n1463;
  assign n1465 = ~n1455 & n1462;
  assign n1466 = ~n8786 & n8789;
  assign n1467 = ~n1443 & ~n1466;
  assign n1468 = n859 & ~n8727;
  assign n1469 = n8727 & ~n1015;
  assign n1470 = ~n859 & ~n1015;
  assign n1471 = ~n1469 & ~n1470;
  assign n1472 = ~n1015 & ~n1468;
  assign n1473 = ~n1467 & ~n8790;
  assign n1474 = ~n1015 & ~n1473;
  assign n1475 = ~n8650 & ~n8787;
  assign n1476 = ~n1293 & n1475;
  assign n1477 = n1293 & ~n1475;
  assign n1478 = ~n1476 & ~n1477;
  assign n1479 = n1457 & n1478;
  assign n1480 = ~n1457 & ~n1478;
  assign n1481 = ~n1479 & ~n1480;
  assign n1482 = ~n1474 & n1481;
  assign n1483 = n1474 & ~n1481;
  assign n1484 = ~n1482 & ~n1483;
  assign n1485 = ~n1021 & n8764;
  assign n1486 = n1021 & ~n1293;
  assign n1487 = ~n8765 & ~n1486;
  assign n1488 = ~n1293 & ~n1485;
  assign n1489 = ~n1021 & n8768;
  assign n1490 = n8791 & ~n1489;
  assign n1491 = ~n1475 & n1490;
  assign n1492 = n1475 & ~n1490;
  assign n1493 = ~n1491 & ~n1492;
  assign n1494 = ~n8767 & n8782;
  assign n1495 = n8767 & n8783;
  assign n1496 = ~n1494 & ~n1495;
  assign n1497 = ~n1325 & n8784;
  assign n1498 = n1325 & n1433;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = ~n1495 & n1499;
  assign n1501 = ~n1494 & n1500;
  assign n1502 = n1496 & n1499;
  assign n1503 = n1493 & n8792;
  assign n1504 = ~n1491 & ~n1503;
  assign n1505 = n992 & n8725;
  assign n1506 = n987 & ~n8725;
  assign n1507 = ~n8650 & ~n1325;
  assign n1508 = n8650 & n1325;
  assign n1509 = ~n1507 & ~n1508;
  assign n1510 = ~n8724 & n1325;
  assign n1511 = ~n8724 & ~n1509;
  assign n1512 = ~n1506 & ~n8793;
  assign n1513 = ~n1505 & ~n1506;
  assign n1514 = ~n8793 & n1513;
  assign n1515 = ~n1505 & n1512;
  assign n1516 = ~n1021 & n8782;
  assign n1517 = n1021 & n8783;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = n8767 & n1433;
  assign n1520 = ~n8767 & n8784;
  assign n1521 = ~n1519 & ~n1520;
  assign n1522 = ~n1517 & n1521;
  assign n1523 = ~n1516 & n1522;
  assign n1524 = n1518 & n1521;
  assign n1525 = n8794 & n8795;
  assign n1526 = ~n8794 & ~n8795;
  assign n1527 = ~n1525 & ~n1526;
  assign n1528 = ~n1504 & n1527;
  assign n1529 = n1504 & ~n1527;
  assign n1530 = ~n1528 & ~n1529;
  assign n1531 = n1484 & n1530;
  assign n1532 = ~n1482 & ~n1531;
  assign n1533 = ~n1021 & n8781;
  assign n1534 = n1021 & ~n1428;
  assign n1535 = ~n8783 & ~n1534;
  assign n1536 = ~n1428 & ~n1533;
  assign n1537 = ~n1021 & n8784;
  assign n1538 = n8796 & ~n1537;
  assign n1539 = ~n1006 & n1538;
  assign n1540 = n1006 & ~n1538;
  assign n1541 = ~n1539 & ~n1540;
  assign n1542 = n992 & n1325;
  assign n1543 = n987 & ~n1325;
  assign n1544 = ~n8650 & ~n8767;
  assign n1545 = n8650 & n8767;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = ~n8724 & n8767;
  assign n1548 = ~n8724 & ~n1546;
  assign n1549 = ~n1543 & ~n8797;
  assign n1550 = ~n1542 & ~n1543;
  assign n1551 = ~n8797 & n1550;
  assign n1552 = ~n1542 & n1549;
  assign n1553 = n1541 & n8798;
  assign n1554 = ~n1541 & ~n8798;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = ~n1476 & ~n1479;
  assign n1557 = ~n1525 & ~n1528;
  assign n1558 = ~n1556 & ~n1557;
  assign n1559 = n1556 & n1557;
  assign n1560 = ~n1556 & ~n1558;
  assign n1561 = ~n1556 & n1557;
  assign n1562 = ~n1557 & ~n1558;
  assign n1563 = n1556 & ~n1557;
  assign n1564 = ~n8799 & ~n8800;
  assign n1565 = ~n1558 & ~n1559;
  assign n1566 = n1555 & ~n8801;
  assign n1567 = ~n1555 & n8801;
  assign n1568 = ~n8801 & ~n1566;
  assign n1569 = ~n1555 & ~n8801;
  assign n1570 = n1555 & ~n1566;
  assign n1571 = n1555 & n8801;
  assign n1572 = ~n8802 & ~n8803;
  assign n1573 = ~n1566 & ~n1567;
  assign n1574 = ~n1532 & ~n8804;
  assign n1575 = n854 & n992;
  assign n1576 = ~n854 & n987;
  assign n1577 = n8650 & n8787;
  assign n1578 = ~n1475 & ~n1577;
  assign n1579 = ~n8724 & n8787;
  assign n1580 = ~n8724 & ~n1578;
  assign n1581 = ~n1576 & ~n8805;
  assign n1582 = ~n1575 & ~n1576;
  assign n1583 = ~n8805 & n1582;
  assign n1584 = ~n1575 & n1581;
  assign n1585 = ~n8725 & n8782;
  assign n1586 = n8725 & n8783;
  assign n1587 = ~n1585 & ~n1586;
  assign n1588 = ~n997 & n8784;
  assign n1589 = n997 & n1433;
  assign n1590 = ~n1588 & ~n1589;
  assign n1591 = ~n1586 & n1590;
  assign n1592 = ~n1585 & n1591;
  assign n1593 = n1587 & n1590;
  assign n1594 = n8806 & n8807;
  assign n1595 = ~n8806 & ~n8807;
  assign n1596 = ~n1594 & ~n1595;
  assign n1597 = ~n314 & ~n8709;
  assign n1598 = ~n380 & ~n415;
  assign n1599 = ~n415 & n1597;
  assign n1600 = ~n380 & n1599;
  assign n1601 = n1597 & n1598;
  assign n1602 = ~n359 & ~n418;
  assign n1603 = ~n820 & n1602;
  assign n1604 = ~n8648 & ~n658;
  assign n1605 = ~n8648 & ~n823;
  assign n1606 = ~n658 & n1605;
  assign n1607 = ~n823 & n1604;
  assign n1608 = n1603 & n8809;
  assign n1609 = n8808 & n8809;
  assign n1610 = n1603 & n1609;
  assign n1611 = n8808 & n1603;
  assign n1612 = n8809 & n1611;
  assign n1613 = n8808 & n1608;
  assign n1614 = ~n270 & ~n377;
  assign n1615 = ~n341 & ~n377;
  assign n1616 = ~n270 & ~n656;
  assign n1617 = n1615 & n1616;
  assign n1618 = n1058 & n1614;
  assign n1619 = n1120 & n8811;
  assign n1620 = n8670 & n1619;
  assign n1621 = n8670 & n8810;
  assign n1622 = n1120 & n1621;
  assign n1623 = ~n341 & n1622;
  assign n1624 = ~n270 & n1623;
  assign n1625 = ~n377 & n1624;
  assign n1626 = ~n656 & n1625;
  assign n1627 = n8810 & n1620;
  assign n1628 = ~n431 & ~n487;
  assign n1629 = ~n387 & n1628;
  assign n1630 = ~n8629 & ~n8647;
  assign n1631 = n816 & n1630;
  assign n1632 = n1629 & n1631;
  assign n1633 = n8736 & n1632;
  assign n1634 = ~n277 & ~n414;
  assign n1635 = ~n821 & ~n884;
  assign n1636 = ~n514 & n1635;
  assign n1637 = ~n277 & ~n821;
  assign n1638 = ~n414 & n1637;
  assign n1639 = ~n514 & n1638;
  assign n1640 = ~n884 & n1639;
  assign n1641 = n1634 & n1636;
  assign n1642 = ~n560 & ~n1345;
  assign n1643 = ~n223 & ~n287;
  assign n1644 = n615 & n1643;
  assign n1645 = n1642 & n1643;
  assign n1646 = n615 & n1645;
  assign n1647 = n1642 & n1644;
  assign n1648 = n8813 & n8814;
  assign n1649 = ~n8629 & ~n387;
  assign n1650 = ~n8647 & n1649;
  assign n1651 = n615 & n1628;
  assign n1652 = n1650 & n1651;
  assign n1653 = n8736 & n1652;
  assign n1654 = n816 & n1643;
  assign n1655 = n1642 & n1654;
  assign n1656 = n8813 & n1655;
  assign n1657 = n1653 & n1656;
  assign n1658 = n1633 & n1648;
  assign n1659 = ~n475 & ~n8686;
  assign n1660 = ~n204 & ~n382;
  assign n1661 = n1659 & n1660;
  assign n1662 = n722 & n1090;
  assign n1663 = ~n220 & ~n430;
  assign n1664 = n1343 & n1663;
  assign n1665 = n1662 & n1664;
  assign n1666 = n1233 & n1662;
  assign n1667 = ~n220 & n1666;
  assign n1668 = ~n204 & n1667;
  assign n1669 = ~n444 & n1668;
  assign n1670 = ~n382 & n1669;
  assign n1671 = ~n430 & n1670;
  assign n1672 = ~n8686 & n1671;
  assign n1673 = ~n220 & ~n382;
  assign n1674 = ~n204 & ~n8686;
  assign n1675 = n1673 & n1674;
  assign n1676 = ~n430 & ~n444;
  assign n1677 = n1233 & n1676;
  assign n1678 = n1662 & n1677;
  assign n1679 = n1675 & n1678;
  assign n1680 = n1661 & n1665;
  assign n1681 = ~n198 & ~n542;
  assign n1682 = ~n436 & n1681;
  assign n1683 = ~n490 & ~n967;
  assign n1684 = n257 & n1683;
  assign n1685 = n864 & n1684;
  assign n1686 = ~n542 & n864;
  assign n1687 = ~n256 & n1686;
  assign n1688 = ~n255 & n1687;
  assign n1689 = ~n198 & n1688;
  assign n1690 = ~n436 & n1689;
  assign n1691 = ~n967 & n1690;
  assign n1692 = ~n490 & n1691;
  assign n1693 = ~n198 & ~n967;
  assign n1694 = ~n542 & n1693;
  assign n1695 = ~n436 & ~n490;
  assign n1696 = n257 & n1695;
  assign n1697 = n864 & n1696;
  assign n1698 = n1694 & n1697;
  assign n1699 = n1682 & n1685;
  assign n1700 = n8816 & n8817;
  assign n1701 = n8815 & n1700;
  assign n1702 = n8736 & n8814;
  assign n1703 = n816 & n1702;
  assign n1704 = n8817 & n1703;
  assign n1705 = n8813 & n1704;
  assign n1706 = n8816 & n1705;
  assign n1707 = n8812 & n1706;
  assign n1708 = ~n8629 & n1707;
  assign n1709 = ~n8647 & n1708;
  assign n1710 = ~n431 & n1709;
  assign n1711 = ~n487 & n1710;
  assign n1712 = ~n387 & n1711;
  assign n1713 = n8812 & n1701;
  assign n1714 = ~n240 & ~n511;
  assign n1715 = ~n861 & n1714;
  assign n1716 = n1399 & n1715;
  assign n1717 = n8697 & n1716;
  assign n1718 = ~n210 & ~n339;
  assign n1719 = n866 & n1718;
  assign n1720 = n1248 & n1642;
  assign n1721 = n866 & n1642;
  assign n1722 = n1248 & n1721;
  assign n1723 = ~n210 & n1722;
  assign n1724 = ~n339 & n1723;
  assign n1725 = n1248 & n1718;
  assign n1726 = n1721 & n1725;
  assign n1727 = n1719 & n1720;
  assign n1728 = ~n341 & ~n636;
  assign n1729 = ~n164 & ~n1163;
  assign n1730 = n291 & n1729;
  assign n1731 = n1728 & n1730;
  assign n1732 = n8813 & n1731;
  assign n1733 = n8819 & n1732;
  assign n1734 = n8697 & n1399;
  assign n1735 = n291 & n1734;
  assign n1736 = n8813 & n1735;
  assign n1737 = n8819 & n1736;
  assign n1738 = ~n240 & n1737;
  assign n1739 = ~n341 & n1738;
  assign n1740 = ~n164 & n1739;
  assign n1741 = ~n861 & n1740;
  assign n1742 = ~n636 & n1741;
  assign n1743 = ~n511 & n1742;
  assign n1744 = ~n1163 & n1743;
  assign n1745 = ~n861 & n1729;
  assign n1746 = n1399 & n1745;
  assign n1747 = n8697 & n1746;
  assign n1748 = n291 & n1714;
  assign n1749 = n1728 & n1748;
  assign n1750 = n8813 & n1749;
  assign n1751 = n8819 & n1750;
  assign n1752 = n1747 & n1751;
  assign n1753 = n1717 & n1733;
  assign n1754 = ~n204 & ~n359;
  assign n1755 = ~n331 & ~n387;
  assign n1756 = n1754 & n1755;
  assign n1757 = n712 & n1392;
  assign n1758 = n804 & n1757;
  assign n1759 = ~n331 & n1757;
  assign n1760 = ~n255 & n1759;
  assign n1761 = ~n359 & n1760;
  assign n1762 = ~n204 & n1761;
  assign n1763 = ~n387 & n1762;
  assign n1764 = ~n448 & n1763;
  assign n1765 = ~n255 & ~n359;
  assign n1766 = ~n204 & ~n331;
  assign n1767 = n1765 & n1766;
  assign n1768 = ~n387 & ~n448;
  assign n1769 = n1392 & n1768;
  assign n1770 = n712 & n1769;
  assign n1771 = n1767 & n1770;
  assign n1772 = n1756 & n1758;
  assign n1773 = ~n490 & ~n817;
  assign n1774 = ~n223 & ~n815;
  assign n1775 = n1773 & n1774;
  assign n1776 = n446 & n1107;
  assign n1777 = n1775 & n1776;
  assign n1778 = ~n393 & ~n610;
  assign n1779 = ~n280 & n1778;
  assign n1780 = n655 & n1779;
  assign n1781 = ~n280 & ~n490;
  assign n1782 = ~n393 & ~n817;
  assign n1783 = n1781 & n1782;
  assign n1784 = n1776 & n1783;
  assign n1785 = ~n223 & ~n610;
  assign n1786 = ~n815 & n1785;
  assign n1787 = n655 & n1786;
  assign n1788 = n1784 & n1787;
  assign n1789 = n1777 & n1780;
  assign n1790 = n655 & n1107;
  assign n1791 = ~n815 & n1790;
  assign n1792 = n8821 & n1791;
  assign n1793 = n446 & n1792;
  assign n1794 = ~n280 & n1793;
  assign n1795 = ~n223 & n1794;
  assign n1796 = ~n817 & n1795;
  assign n1797 = ~n490 & n1796;
  assign n1798 = ~n610 & n1797;
  assign n1799 = ~n393 & n1798;
  assign n1800 = n8821 & n8822;
  assign n1801 = ~n207 & ~n386;
  assign n1802 = ~n8640 & ~n721;
  assign n1803 = ~n207 & ~n8640;
  assign n1804 = ~n386 & n1803;
  assign n1805 = ~n721 & n1804;
  assign n1806 = n1801 & n1802;
  assign n1807 = n185 & ~n820;
  assign n1808 = n875 & n1807;
  assign n1809 = n8824 & n1808;
  assign n1810 = ~n492 & ~n608;
  assign n1811 = ~n641 & ~n967;
  assign n1812 = ~n492 & ~n641;
  assign n1813 = ~n608 & ~n967;
  assign n1814 = n1812 & n1813;
  assign n1815 = n1810 & n1811;
  assign n1816 = ~n492 & n1402;
  assign n1817 = ~n967 & n1816;
  assign n1818 = ~n641 & n1817;
  assign n1819 = ~n608 & n1818;
  assign n1820 = n1402 & n8825;
  assign n1821 = n300 & n945;
  assign n1822 = n381 & n945;
  assign n1823 = n300 & n1822;
  assign n1824 = n381 & n1821;
  assign n1825 = n8826 & n8827;
  assign n1826 = n1809 & n1825;
  assign n1827 = n8823 & n1826;
  assign n1828 = n381 & n8824;
  assign n1829 = n875 & n1828;
  assign n1830 = n945 & n1829;
  assign n1831 = n8826 & n1830;
  assign n1832 = n300 & n1831;
  assign n1833 = n8823 & n1832;
  assign n1834 = n8820 & n1833;
  assign n1835 = ~n8630 & n1834;
  assign n1836 = ~n8631 & n1835;
  assign n1837 = ~n820 & n1836;
  assign n1838 = n8820 & n1827;
  assign n1839 = ~n8818 & ~n8828;
  assign n1840 = ~n8705 & ~n1839;
  assign n1841 = n8818 & ~n1840;
  assign n1842 = n8705 & n8818;
  assign n1843 = pi6  & pi22 ;
  assign n1844 = pi6  & ~n91;
  assign n1845 = n351 & ~n1844;
  assign n1846 = ~n1843 & ~n1845;
  assign n1847 = ~n8650 & ~n1846;
  assign n1848 = ~n8705 & ~n8818;
  assign n1849 = ~n8818 & n1840;
  assign n1850 = ~n8818 & n8828;
  assign n1851 = ~n8705 & n1850;
  assign n1852 = n8828 & n1848;
  assign n1853 = n1847 & ~n8830;
  assign n1854 = ~n8829 & n1847;
  assign n1855 = ~n8830 & n1854;
  assign n1856 = ~n8829 & ~n1855;
  assign n1857 = ~n8829 & ~n1853;
  assign n1858 = n1596 & ~n8831;
  assign n1859 = ~n1594 & ~n1858;
  assign n1860 = n8682 & n8705;
  assign n1861 = ~n8682 & n8705;
  assign n1862 = n8682 & ~n8705;
  assign n1863 = ~n1861 & ~n1862;
  assign n1864 = ~n845 & ~n1860;
  assign n1865 = ~n1021 & n8832;
  assign n1866 = ~n846 & ~n8832;
  assign n1867 = n8666 & ~n8832;
  assign n1868 = ~n846 & n1021;
  assign n1869 = ~n8833 & ~n1868;
  assign n1870 = ~n846 & ~n1865;
  assign n1871 = n8666 & ~n1860;
  assign n1872 = n8832 & ~n1871;
  assign n1873 = ~n1021 & n1872;
  assign n1874 = n1865 & ~n1871;
  assign n1875 = n8834 & ~n8835;
  assign n1876 = ~n358 & n1875;
  assign n1877 = n358 & ~n1875;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = n8765 & n8767;
  assign n1880 = n8766 & ~n8767;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = n8768 & ~n1325;
  assign n1883 = n1309 & n1325;
  assign n1884 = ~n1882 & ~n1883;
  assign n1885 = ~n1879 & n1884;
  assign n1886 = ~n1880 & n1885;
  assign n1887 = ~n1879 & ~n1882;
  assign n1888 = ~n1880 & ~n1883;
  assign n1889 = n1887 & n1888;
  assign n1890 = n1881 & n1884;
  assign n1891 = n1878 & n8836;
  assign n1892 = ~n1876 & ~n1891;
  assign n1893 = ~n1859 & ~n1892;
  assign n1894 = ~n849 & ~n855;
  assign n1895 = ~n8650 & ~n8706;
  assign n1896 = ~n854 & n1895;
  assign n1897 = n849 & ~n8706;
  assign n1898 = ~n1896 & ~n1897;
  assign n1899 = ~n8706 & ~n1894;
  assign n1900 = n1859 & n1892;
  assign n1901 = ~n1859 & ~n1893;
  assign n1902 = ~n1859 & n1892;
  assign n1903 = ~n1892 & ~n1893;
  assign n1904 = n1859 & ~n1892;
  assign n1905 = ~n8838 & ~n8839;
  assign n1906 = ~n1893 & ~n1900;
  assign n1907 = ~n8837 & ~n8840;
  assign n1908 = ~n1893 & ~n1907;
  assign n1909 = ~n1493 & ~n8792;
  assign n1910 = ~n1503 & ~n1909;
  assign n1911 = ~n1908 & n1910;
  assign n1912 = n1908 & ~n1910;
  assign n1913 = ~n1911 & ~n1912;
  assign n1914 = n1467 & n8790;
  assign n1915 = ~n1467 & ~n1473;
  assign n1916 = ~n8790 & ~n1473;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = ~n1473 & ~n1914;
  assign n1919 = n1913 & ~n8841;
  assign n1920 = ~n1911 & ~n1919;
  assign n1921 = ~n1484 & ~n1530;
  assign n1922 = ~n1531 & ~n1921;
  assign n1923 = ~n1920 & n1922;
  assign n1924 = ~n1913 & n8841;
  assign n1925 = n1913 & ~n1919;
  assign n1926 = ~n8841 & ~n1919;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = ~n1919 & ~n1924;
  assign n1929 = n8651 & n992;
  assign n1930 = ~n8651 & n987;
  assign n1931 = n8650 & n854;
  assign n1932 = ~n855 & ~n1931;
  assign n1933 = n854 & ~n8724;
  assign n1934 = ~n8724 & ~n1932;
  assign n1935 = ~n1930 & ~n8843;
  assign n1936 = ~n1929 & ~n1930;
  assign n1937 = ~n8843 & n1936;
  assign n1938 = ~n1929 & n1935;
  assign n1939 = ~n997 & n8782;
  assign n1940 = n997 & n8783;
  assign n1941 = ~n1939 & ~n1940;
  assign n1942 = n1433 & n8787;
  assign n1943 = n8784 & ~n8787;
  assign n1944 = ~n1942 & ~n1943;
  assign n1945 = ~n1940 & n1944;
  assign n1946 = ~n1939 & n1945;
  assign n1947 = n1941 & n1944;
  assign n1948 = n8844 & n8845;
  assign n1949 = ~n8844 & ~n8845;
  assign n1950 = ~n8844 & n8845;
  assign n1951 = n8844 & ~n8845;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = ~n1948 & ~n1949;
  assign n1954 = ~n8832 & ~n1871;
  assign n1955 = ~n8666 & ~n8832;
  assign n1956 = ~n1021 & n8847;
  assign n1957 = n1021 & n8833;
  assign n1958 = ~n1956 & ~n1957;
  assign n1959 = ~n846 & n8832;
  assign n1960 = n8767 & n1959;
  assign n1961 = ~n8767 & n1872;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = ~n1957 & n1962;
  assign n1964 = ~n1956 & n1963;
  assign n1965 = n1958 & n1962;
  assign n1966 = ~n8846 & n8848;
  assign n1967 = ~n1948 & ~n1966;
  assign n1968 = ~n1878 & ~n8836;
  assign n1969 = ~n1891 & ~n1968;
  assign n1970 = ~n1967 & n1969;
  assign n1971 = ~n1596 & n8831;
  assign n1972 = ~n1858 & ~n1971;
  assign n1973 = n1967 & ~n1969;
  assign n1974 = ~n1967 & ~n1970;
  assign n1975 = n1969 & ~n1970;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = ~n1970 & ~n1973;
  assign n1978 = n1972 & ~n8849;
  assign n1979 = ~n1970 & ~n1978;
  assign n1980 = n8786 & ~n8789;
  assign n1981 = n8789 & ~n1466;
  assign n1982 = n8786 & n8789;
  assign n1983 = ~n8786 & ~n1466;
  assign n1984 = ~n8786 & ~n8789;
  assign n1985 = ~n8850 & ~n8851;
  assign n1986 = ~n1466 & ~n1980;
  assign n1987 = n1979 & n8852;
  assign n1988 = ~n1979 & ~n8852;
  assign n1989 = n8837 & n8840;
  assign n1990 = ~n8840 & ~n1907;
  assign n1991 = n8837 & ~n8840;
  assign n1992 = ~n8837 & ~n1907;
  assign n1993 = ~n8837 & n8840;
  assign n1994 = ~n8853 & ~n8854;
  assign n1995 = ~n1907 & ~n1989;
  assign n1996 = ~n1988 & n8855;
  assign n1997 = ~n1979 & ~n1988;
  assign n1998 = ~n8852 & ~n1988;
  assign n1999 = ~n1997 & ~n1998;
  assign n2000 = ~n1987 & ~n1988;
  assign n2001 = ~n8855 & ~n8856;
  assign n2002 = ~n1988 & ~n2001;
  assign n2003 = ~n1987 & ~n1996;
  assign n2004 = ~n8842 & ~n8857;
  assign n2005 = ~n8829 & ~n8830;
  assign n2006 = n1847 & ~n1855;
  assign n2007 = n1847 & ~n2005;
  assign n2008 = ~n8830 & n8831;
  assign n2009 = ~n1853 & n2005;
  assign n2010 = ~n8858 & ~n8859;
  assign n2011 = n8765 & n1325;
  assign n2012 = n8766 & ~n1325;
  assign n2013 = ~n2011 & ~n2012;
  assign n2014 = n8725 & n1309;
  assign n2015 = ~n8725 & n8768;
  assign n2016 = ~n2014 & ~n2015;
  assign n2017 = ~n2011 & n2016;
  assign n2018 = ~n2012 & n2017;
  assign n2019 = ~n2011 & ~n2015;
  assign n2020 = ~n2012 & ~n2014;
  assign n2021 = n2019 & n2020;
  assign n2022 = n2013 & n2016;
  assign n2023 = ~n2010 & n8860;
  assign n2024 = ~n8620 & ~n8650;
  assign n2025 = ~n8818 & n2024;
  assign n2026 = n8818 & ~n2024;
  assign n2027 = ~n2025 & ~n2026;
  assign n2028 = n8818 & n8828;
  assign n2029 = n8818 & ~n8828;
  assign n2030 = ~n1850 & ~n2029;
  assign n2031 = ~n1839 & ~n2028;
  assign n2032 = ~n1021 & n8861;
  assign n2033 = ~n1840 & ~n8861;
  assign n2034 = n8705 & ~n8861;
  assign n2035 = n1021 & ~n1840;
  assign n2036 = ~n8862 & ~n2035;
  assign n2037 = ~n1840 & ~n2032;
  assign n2038 = n8705 & ~n2028;
  assign n2039 = n8861 & ~n2038;
  assign n2040 = ~n1021 & n2039;
  assign n2041 = n2032 & ~n2038;
  assign n2042 = n8863 & ~n8864;
  assign n2043 = ~n2025 & n2042;
  assign n2044 = ~n2026 & n2043;
  assign n2045 = n2027 & n2042;
  assign n2046 = ~n2025 & ~n8865;
  assign n2047 = n2010 & ~n8860;
  assign n2048 = ~n2023 & ~n2047;
  assign n2049 = ~n2046 & n2048;
  assign n2050 = ~n2023 & ~n2049;
  assign n2051 = ~n8767 & n8847;
  assign n2052 = n8767 & n8833;
  assign n2053 = ~n2051 & ~n2052;
  assign n2054 = ~n1325 & n1872;
  assign n2055 = n1325 & n1959;
  assign n2056 = ~n2054 & ~n2055;
  assign n2057 = ~n2052 & n2056;
  assign n2058 = ~n2051 & n2057;
  assign n2059 = n2053 & n2056;
  assign n2060 = n8725 & n8765;
  assign n2061 = ~n8725 & n8766;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = ~n997 & n8768;
  assign n2064 = n997 & n1309;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = ~n2060 & n2065;
  assign n2067 = ~n2061 & n2066;
  assign n2068 = ~n2060 & ~n2063;
  assign n2069 = ~n2061 & ~n2064;
  assign n2070 = n2068 & n2069;
  assign n2071 = n2062 & n2065;
  assign n2072 = n8866 & n8867;
  assign n2073 = ~n8866 & ~n8867;
  assign n2074 = n8866 & ~n8867;
  assign n2075 = ~n8866 & n8867;
  assign n2076 = ~n2074 & ~n2075;
  assign n2077 = ~n2072 & ~n2073;
  assign n2078 = n8782 & ~n8787;
  assign n2079 = n8783 & n8787;
  assign n2080 = ~n2078 & ~n2079;
  assign n2081 = ~n854 & n8784;
  assign n2082 = n854 & n1433;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = ~n2079 & n2083;
  assign n2085 = ~n2078 & n2084;
  assign n2086 = n2080 & n2083;
  assign n2087 = ~n8868 & n8869;
  assign n2088 = ~n2072 & ~n2087;
  assign n2089 = n8846 & ~n8848;
  assign n2090 = ~n1966 & ~n2089;
  assign n2091 = ~n2088 & n2090;
  assign n2092 = ~n66 & ~n8650;
  assign n2093 = ~n8818 & n2092;
  assign n2094 = n8818 & ~n2092;
  assign n2095 = ~n2093 & ~n2094;
  assign n2096 = ~n8861 & ~n2038;
  assign n2097 = ~n8705 & ~n8861;
  assign n2098 = ~n1021 & n8870;
  assign n2099 = n1021 & n8862;
  assign n2100 = ~n2098 & ~n2099;
  assign n2101 = ~n1840 & n8861;
  assign n2102 = n8767 & n2101;
  assign n2103 = ~n8767 & n2039;
  assign n2104 = ~n2102 & ~n2103;
  assign n2105 = ~n2099 & n2104;
  assign n2106 = ~n2098 & n2105;
  assign n2107 = n2100 & n2104;
  assign n2108 = ~n2093 & n8871;
  assign n2109 = ~n2094 & n2108;
  assign n2110 = n2095 & n8871;
  assign n2111 = ~n2093 & ~n8872;
  assign n2112 = n992 & n1846;
  assign n2113 = n987 & ~n1846;
  assign n2114 = n8650 & n8651;
  assign n2115 = ~n358 & ~n2114;
  assign n2116 = n8651 & ~n8724;
  assign n2117 = ~n8724 & ~n2115;
  assign n2118 = ~n2113 & ~n8873;
  assign n2119 = ~n2112 & ~n2113;
  assign n2120 = ~n8873 & n2119;
  assign n2121 = ~n2112 & n2118;
  assign n2122 = ~n2111 & n8874;
  assign n2123 = n2111 & ~n8874;
  assign n2124 = ~n2122 & ~n2123;
  assign n2125 = n997 & n8765;
  assign n2126 = ~n997 & n8766;
  assign n2127 = ~n2125 & ~n2126;
  assign n2128 = n1309 & n8787;
  assign n2129 = n8768 & ~n8787;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = ~n2125 & n2130;
  assign n2132 = ~n2126 & n2131;
  assign n2133 = ~n2125 & ~n2129;
  assign n2134 = ~n2126 & ~n2128;
  assign n2135 = n2133 & n2134;
  assign n2136 = n2127 & n2130;
  assign n2137 = ~n1325 & n8847;
  assign n2138 = n1325 & n8833;
  assign n2139 = ~n2137 & ~n2138;
  assign n2140 = n8725 & n1959;
  assign n2141 = ~n8725 & n1872;
  assign n2142 = ~n2140 & ~n2141;
  assign n2143 = ~n2138 & n2142;
  assign n2144 = ~n2137 & n2143;
  assign n2145 = n2139 & n2142;
  assign n2146 = n8875 & n8876;
  assign n2147 = ~n8875 & ~n8876;
  assign n2148 = ~n8875 & n8876;
  assign n2149 = n8875 & ~n8876;
  assign n2150 = ~n2148 & ~n2149;
  assign n2151 = ~n2146 & ~n2147;
  assign n2152 = ~n854 & n8782;
  assign n2153 = n854 & n8783;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = n8651 & n1433;
  assign n2156 = ~n8651 & n8784;
  assign n2157 = ~n2155 & ~n2156;
  assign n2158 = ~n2153 & n2157;
  assign n2159 = ~n2152 & n2158;
  assign n2160 = n2154 & n2157;
  assign n2161 = ~n8877 & n8878;
  assign n2162 = ~n2146 & ~n2161;
  assign n2163 = n2124 & ~n2162;
  assign n2164 = ~n2122 & ~n2163;
  assign n2165 = n2088 & ~n2090;
  assign n2166 = ~n2091 & ~n2165;
  assign n2167 = ~n2164 & n2166;
  assign n2168 = ~n2091 & ~n2167;
  assign n2169 = ~n2050 & ~n2168;
  assign n2170 = ~n1972 & n8849;
  assign n2171 = n1972 & ~n1978;
  assign n2172 = ~n8849 & ~n1978;
  assign n2173 = ~n2171 & ~n2172;
  assign n2174 = ~n1978 & ~n2170;
  assign n2175 = n2050 & n2168;
  assign n2176 = ~n2050 & ~n2169;
  assign n2177 = ~n2050 & n2168;
  assign n2178 = ~n2168 & ~n2169;
  assign n2179 = n2050 & ~n2168;
  assign n2180 = ~n8880 & ~n8881;
  assign n2181 = ~n2169 & ~n2175;
  assign n2182 = ~n8879 & ~n8882;
  assign n2183 = ~n2169 & ~n2182;
  assign n2184 = n8855 & ~n8856;
  assign n2185 = ~n8855 & n8856;
  assign n2186 = ~n2184 & ~n2185;
  assign n2187 = ~n2183 & ~n2186;
  assign n2188 = ~n2027 & ~n2042;
  assign n2189 = ~n2026 & n2046;
  assign n2190 = n2042 & ~n8865;
  assign n2191 = ~n2189 & ~n2190;
  assign n2192 = ~n8865 & ~n2188;
  assign n2193 = n8868 & ~n8869;
  assign n2194 = n8869 & ~n2087;
  assign n2195 = n8868 & n8869;
  assign n2196 = ~n8868 & ~n2087;
  assign n2197 = ~n8868 & ~n8869;
  assign n2198 = ~n8884 & ~n8885;
  assign n2199 = ~n2087 & ~n2193;
  assign n2200 = ~n8883 & ~n8886;
  assign n2201 = ~n8622 & ~n8650;
  assign n2202 = ~n295 & ~n625;
  assign n2203 = n332 & n2202;
  assign n2204 = n654 & n1403;
  assign n2205 = n2203 & n2204;
  assign n2206 = ~n210 & ~n8652;
  assign n2207 = ~n511 & n2206;
  assign n2208 = ~n210 & n1191;
  assign n2209 = ~n197 & ~n255;
  assign n2210 = ~n642 & n2209;
  assign n2211 = n8729 & n2210;
  assign n2212 = n8887 & n2211;
  assign n2213 = n332 & n8729;
  assign n2214 = n8887 & n2213;
  assign n2215 = n654 & n2214;
  assign n2216 = n1403 & n2215;
  assign n2217 = ~n295 & n2216;
  assign n2218 = ~n255 & n2217;
  assign n2219 = ~n197 & n2218;
  assign n2220 = ~n642 & n2219;
  assign n2221 = ~n625 & n2220;
  assign n2222 = ~n255 & ~n295;
  assign n2223 = n332 & n2222;
  assign n2224 = n2204 & n2223;
  assign n2225 = ~n197 & ~n642;
  assign n2226 = ~n625 & n2225;
  assign n2227 = n8729 & n2226;
  assign n2228 = n8887 & n2227;
  assign n2229 = n2224 & n2228;
  assign n2230 = n2205 & n2212;
  assign n2231 = ~n391 & ~n821;
  assign n2232 = ~n1345 & n2231;
  assign n2233 = ~n817 & ~n938;
  assign n2234 = ~n8640 & ~n313;
  assign n2235 = n1333 & n2234;
  assign n2236 = n2233 & n2235;
  assign n2237 = ~n8640 & ~n821;
  assign n2238 = ~n1345 & n2237;
  assign n2239 = ~n313 & ~n391;
  assign n2240 = n1333 & n2239;
  assign n2241 = n2233 & n2240;
  assign n2242 = n2238 & n2241;
  assign n2243 = n2232 & n2236;
  assign n2244 = n8632 & n8889;
  assign n2245 = ~n610 & ~n8678;
  assign n2246 = ~n658 & n2245;
  assign n2247 = ~n443 & ~n450;
  assign n2248 = ~n415 & ~n608;
  assign n2249 = ~n798 & ~n815;
  assign n2250 = n2248 & n2249;
  assign n2251 = n2247 & n2250;
  assign n2252 = ~n8678 & ~n815;
  assign n2253 = ~n658 & n2252;
  assign n2254 = ~n443 & n2253;
  assign n2255 = ~n415 & n2254;
  assign n2256 = ~n608 & n2255;
  assign n2257 = ~n450 & n2256;
  assign n2258 = ~n798 & n2257;
  assign n2259 = ~n610 & n2258;
  assign n2260 = ~n658 & ~n798;
  assign n2261 = ~n815 & n2260;
  assign n2262 = ~n415 & ~n610;
  assign n2263 = ~n608 & ~n8678;
  assign n2264 = n2262 & n2263;
  assign n2265 = n2247 & n2264;
  assign n2266 = n2261 & n2265;
  assign n2267 = n2246 & n2251;
  assign n2268 = ~n228 & ~n544;
  assign n2269 = ~n296 & ~n387;
  assign n2270 = ~n228 & ~n387;
  assign n2271 = ~n296 & ~n544;
  assign n2272 = n2270 & n2271;
  assign n2273 = n2268 & n2269;
  assign n2274 = n684 & n1232;
  assign n2275 = n824 & n2274;
  assign n2276 = ~n8642 & n1232;
  assign n2277 = ~n296 & n2276;
  assign n2278 = ~n475 & n2277;
  assign n2279 = ~n228 & n2278;
  assign n2280 = ~n377 & n2279;
  assign n2281 = ~n544 & n2280;
  assign n2282 = ~n387 & n2281;
  assign n2283 = ~n823 & n2282;
  assign n2284 = n8891 & n2275;
  assign n2285 = n8890 & n8892;
  assign n2286 = n2244 & n2285;
  assign n2287 = n1333 & n8890;
  assign n2288 = n8888 & n2287;
  assign n2289 = n8632 & n2288;
  assign n2290 = n8892 & n2289;
  assign n2291 = ~n313 & n2290;
  assign n2292 = ~n8640 & n2291;
  assign n2293 = ~n821 & n2292;
  assign n2294 = ~n938 & n2293;
  assign n2295 = ~n817 & n2294;
  assign n2296 = ~n1345 & n2295;
  assign n2297 = ~n391 & n2296;
  assign n2298 = n8888 & n2286;
  assign n2299 = n8818 & ~n8893;
  assign n2300 = ~n8893 & ~n2299;
  assign n2301 = ~n8818 & ~n8893;
  assign n2302 = n1021 & ~n8818;
  assign n2303 = ~n1021 & n8893;
  assign n2304 = ~n8818 & ~n2303;
  assign n2305 = ~n8894 & ~n2302;
  assign n2306 = n2201 & n8895;
  assign n2307 = ~n2201 & ~n8895;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = ~n8767 & n8870;
  assign n2310 = n8767 & n8862;
  assign n2311 = ~n2309 & ~n2310;
  assign n2312 = ~n1325 & n2039;
  assign n2313 = n1325 & n2101;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = ~n2310 & n2314;
  assign n2316 = ~n2309 & n2315;
  assign n2317 = n2311 & n2314;
  assign n2318 = n2308 & n8896;
  assign n2319 = ~n2306 & ~n2318;
  assign n2320 = n8620 & n992;
  assign n2321 = ~n8620 & n987;
  assign n2322 = n8650 & n1846;
  assign n2323 = ~n1847 & ~n2322;
  assign n2324 = ~n8724 & n1846;
  assign n2325 = ~n8724 & ~n2323;
  assign n2326 = ~n2321 & ~n8897;
  assign n2327 = ~n2320 & ~n2321;
  assign n2328 = ~n8897 & n2327;
  assign n2329 = ~n2320 & n2326;
  assign n2330 = ~n2319 & n8898;
  assign n2331 = n2319 & ~n8898;
  assign n2332 = ~n2330 & ~n2331;
  assign n2333 = n8765 & n8787;
  assign n2334 = n8766 & ~n8787;
  assign n2335 = ~n2333 & ~n2334;
  assign n2336 = ~n854 & n8768;
  assign n2337 = n854 & n1309;
  assign n2338 = ~n2336 & ~n2337;
  assign n2339 = ~n2333 & n2338;
  assign n2340 = ~n2334 & n2339;
  assign n2341 = ~n2333 & ~n2336;
  assign n2342 = ~n2334 & ~n2337;
  assign n2343 = n2341 & n2342;
  assign n2344 = n2335 & n2338;
  assign n2345 = ~n8725 & n8847;
  assign n2346 = n8725 & n8833;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = ~n997 & n1872;
  assign n2349 = n997 & n1959;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = ~n2346 & n2350;
  assign n2352 = ~n2345 & n2351;
  assign n2353 = n2347 & n2350;
  assign n2354 = n8899 & n8900;
  assign n2355 = ~n8899 & ~n8900;
  assign n2356 = ~n8899 & n8900;
  assign n2357 = n8899 & ~n8900;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = ~n2354 & ~n2355;
  assign n2360 = ~n8651 & n8782;
  assign n2361 = n8651 & n8783;
  assign n2362 = ~n2360 & ~n2361;
  assign n2363 = n8784 & ~n1846;
  assign n2364 = n1433 & n1846;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = ~n2361 & n2365;
  assign n2367 = ~n2360 & n2366;
  assign n2368 = n2362 & n2365;
  assign n2369 = ~n8901 & n8902;
  assign n2370 = ~n2354 & ~n2369;
  assign n2371 = n2332 & ~n2370;
  assign n2372 = ~n2330 & ~n2371;
  assign n2373 = n8883 & n8886;
  assign n2374 = ~n8883 & ~n2200;
  assign n2375 = ~n8883 & n8886;
  assign n2376 = ~n8886 & ~n2200;
  assign n2377 = n8883 & ~n8886;
  assign n2378 = ~n8903 & ~n8904;
  assign n2379 = ~n2200 & ~n2373;
  assign n2380 = ~n2372 & ~n8905;
  assign n2381 = ~n2200 & ~n2380;
  assign n2382 = n2046 & ~n2048;
  assign n2383 = ~n2049 & ~n2382;
  assign n2384 = ~n2381 & n2383;
  assign n2385 = n2381 & ~n2383;
  assign n2386 = ~n2384 & ~n2385;
  assign n2387 = n2164 & ~n2166;
  assign n2388 = ~n2167 & ~n2387;
  assign n2389 = n2386 & n2388;
  assign n2390 = ~n2384 & ~n2389;
  assign n2391 = n8879 & n8882;
  assign n2392 = ~n8882 & ~n2182;
  assign n2393 = n8879 & ~n8882;
  assign n2394 = ~n8879 & ~n2182;
  assign n2395 = ~n8879 & n8882;
  assign n2396 = ~n8906 & ~n8907;
  assign n2397 = ~n2182 & ~n2391;
  assign n2398 = ~n2390 & ~n8908;
  assign n2399 = ~n1021 & ~n8893;
  assign n2400 = n8818 & ~n2399;
  assign n2401 = ~n1021 & n8894;
  assign n2402 = ~n8767 & n8893;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = n1021 & n2299;
  assign n2405 = n8767 & ~n8818;
  assign n2406 = n8893 & ~n2405;
  assign n2407 = ~n2404 & ~n2406;
  assign n2408 = ~n2401 & n2407;
  assign n2409 = ~n2400 & n2403;
  assign n2410 = ~n8650 & n8909;
  assign n2411 = n66 & n992;
  assign n2412 = ~n66 & n987;
  assign n2413 = n8620 & n8650;
  assign n2414 = ~n2024 & ~n2413;
  assign n2415 = n8620 & ~n8724;
  assign n2416 = ~n8724 & ~n2414;
  assign n2417 = ~n2412 & ~n8910;
  assign n2418 = ~n2411 & ~n2412;
  assign n2419 = ~n8910 & n2418;
  assign n2420 = ~n2411 & n2417;
  assign n2421 = n2410 & n8911;
  assign n2422 = n854 & n8765;
  assign n2423 = ~n854 & n8766;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = n8651 & n1309;
  assign n2426 = ~n8651 & n8768;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = ~n2422 & n2427;
  assign n2429 = ~n2423 & n2428;
  assign n2430 = ~n2422 & ~n2426;
  assign n2431 = ~n2423 & ~n2425;
  assign n2432 = n2430 & n2431;
  assign n2433 = n2424 & n2427;
  assign n2434 = n8782 & ~n1846;
  assign n2435 = n8783 & n1846;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = n8620 & n1433;
  assign n2438 = ~n8620 & n8784;
  assign n2439 = ~n2437 & ~n2438;
  assign n2440 = ~n2435 & n2439;
  assign n2441 = ~n2434 & n2440;
  assign n2442 = n2436 & n2439;
  assign n2443 = n8912 & n8913;
  assign n2444 = ~n8912 & ~n8913;
  assign n2445 = n8912 & ~n8913;
  assign n2446 = ~n8912 & n8913;
  assign n2447 = ~n2445 & ~n2446;
  assign n2448 = ~n2443 & ~n2444;
  assign n2449 = ~n997 & n8847;
  assign n2450 = n997 & n8833;
  assign n2451 = ~n2449 & ~n2450;
  assign n2452 = n8787 & n1959;
  assign n2453 = ~n8787 & n1872;
  assign n2454 = ~n2452 & ~n2453;
  assign n2455 = ~n2450 & n2454;
  assign n2456 = ~n2449 & n2455;
  assign n2457 = n2451 & n2454;
  assign n2458 = ~n8914 & n8915;
  assign n2459 = ~n2443 & ~n2458;
  assign n2460 = ~n2410 & ~n8911;
  assign n2461 = ~n2421 & ~n2460;
  assign n2462 = ~n2459 & n2461;
  assign n2463 = ~n2421 & ~n2462;
  assign n2464 = ~n2095 & ~n8871;
  assign n2465 = ~n2094 & n2111;
  assign n2466 = n8871 & ~n8872;
  assign n2467 = ~n2465 & ~n2466;
  assign n2468 = ~n8872 & ~n2464;
  assign n2469 = ~n2463 & ~n8916;
  assign n2470 = n2463 & n8916;
  assign n2471 = n2463 & ~n8916;
  assign n2472 = ~n2463 & n8916;
  assign n2473 = ~n2471 & ~n2472;
  assign n2474 = ~n2469 & ~n2470;
  assign n2475 = n8877 & ~n8878;
  assign n2476 = n8878 & ~n2161;
  assign n2477 = n8877 & n8878;
  assign n2478 = ~n8877 & ~n2161;
  assign n2479 = ~n8877 & ~n8878;
  assign n2480 = ~n8918 & ~n8919;
  assign n2481 = ~n2161 & ~n2475;
  assign n2482 = ~n8917 & ~n8920;
  assign n2483 = ~n2469 & ~n2482;
  assign n2484 = ~n2124 & n2162;
  assign n2485 = ~n2163 & ~n2484;
  assign n2486 = ~n2483 & n2485;
  assign n2487 = n2483 & ~n2485;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = n2372 & n8905;
  assign n2490 = ~n2372 & n8905;
  assign n2491 = n2372 & ~n8905;
  assign n2492 = ~n2490 & ~n2491;
  assign n2493 = ~n2380 & ~n2489;
  assign n2494 = n2488 & ~n8921;
  assign n2495 = ~n2486 & ~n2494;
  assign n2496 = ~n2386 & ~n2388;
  assign n2497 = ~n2389 & ~n2496;
  assign n2498 = ~n2495 & n2497;
  assign n2499 = ~n2332 & n2370;
  assign n2500 = ~n2371 & ~n2499;
  assign n2501 = ~n2308 & ~n8896;
  assign n2502 = ~n2318 & ~n2501;
  assign n2503 = n8622 & n992;
  assign n2504 = ~n8622 & n987;
  assign n2505 = n66 & n8650;
  assign n2506 = ~n2092 & ~n2505;
  assign n2507 = n66 & ~n8724;
  assign n2508 = ~n8724 & ~n2506;
  assign n2509 = ~n2504 & ~n8922;
  assign n2510 = ~n2503 & ~n2504;
  assign n2511 = ~n8922 & n2510;
  assign n2512 = ~n2503 & n2509;
  assign n2513 = ~n1325 & n8870;
  assign n2514 = n1325 & n8862;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = n8725 & n2101;
  assign n2517 = ~n8725 & n2039;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = ~n2514 & n2518;
  assign n2520 = ~n2513 & n2519;
  assign n2521 = n2515 & n2518;
  assign n2522 = n8923 & n8924;
  assign n2523 = ~n8923 & ~n8924;
  assign n2524 = n8650 & ~n8909;
  assign n2525 = ~n2410 & ~n2524;
  assign n2526 = ~n2523 & n2525;
  assign n2527 = ~n2522 & ~n2523;
  assign n2528 = n2525 & n2527;
  assign n2529 = ~n2522 & ~n2528;
  assign n2530 = ~n2522 & ~n2526;
  assign n2531 = n2502 & ~n8925;
  assign n2532 = ~n2502 & n8925;
  assign n2533 = n8901 & ~n8902;
  assign n2534 = n8902 & ~n2369;
  assign n2535 = n8901 & n8902;
  assign n2536 = ~n8901 & ~n2369;
  assign n2537 = ~n8901 & ~n8902;
  assign n2538 = ~n8926 & ~n8927;
  assign n2539 = ~n2369 & ~n2533;
  assign n2540 = ~n2532 & ~n8928;
  assign n2541 = ~n2531 & ~n2532;
  assign n2542 = ~n8928 & n2541;
  assign n2543 = ~n2531 & ~n2542;
  assign n2544 = ~n2531 & ~n2540;
  assign n2545 = n2500 & ~n8929;
  assign n2546 = ~n2500 & n8929;
  assign n2547 = ~n2545 & ~n2546;
  assign n2548 = n8917 & n8920;
  assign n2549 = ~n2482 & ~n2548;
  assign n2550 = n2547 & n2549;
  assign n2551 = ~n2545 & ~n2550;
  assign n2552 = ~n2488 & n8921;
  assign n2553 = ~n2494 & ~n2552;
  assign n2554 = ~n2551 & n2553;
  assign n2555 = ~n8787 & n8847;
  assign n2556 = n8787 & n8833;
  assign n2557 = ~n2555 & ~n2556;
  assign n2558 = ~n854 & n1872;
  assign n2559 = n854 & n1959;
  assign n2560 = ~n2558 & ~n2559;
  assign n2561 = ~n2556 & n2560;
  assign n2562 = ~n2555 & n2561;
  assign n2563 = n2557 & n2560;
  assign n2564 = n8651 & n8765;
  assign n2565 = ~n8651 & n8766;
  assign n2566 = ~n2564 & ~n2565;
  assign n2567 = n8768 & ~n1846;
  assign n2568 = n1309 & n1846;
  assign n2569 = ~n2567 & ~n2568;
  assign n2570 = ~n2564 & n2569;
  assign n2571 = ~n2565 & n2570;
  assign n2572 = ~n2564 & ~n2567;
  assign n2573 = ~n2565 & ~n2568;
  assign n2574 = n2572 & n2573;
  assign n2575 = n2566 & n2569;
  assign n2576 = n8930 & n8931;
  assign n2577 = ~n8622 & ~n8781;
  assign n2578 = ~n8622 & n8782;
  assign n2579 = n8622 & ~n1428;
  assign n2580 = ~n1433 & ~n2579;
  assign n2581 = ~n2578 & n2580;
  assign n2582 = n1428 & n2581;
  assign n2583 = n1428 & ~n2577;
  assign n2584 = ~n1325 & ~n8893;
  assign n2585 = n8818 & ~n2584;
  assign n2586 = ~n1325 & n8894;
  assign n2587 = ~n8725 & n8893;
  assign n2588 = ~n2586 & ~n2587;
  assign n2589 = n1325 & n2299;
  assign n2590 = n8725 & ~n8818;
  assign n2591 = n8893 & ~n2590;
  assign n2592 = ~n2589 & ~n2591;
  assign n2593 = ~n2586 & n2592;
  assign n2594 = ~n2585 & n2588;
  assign n2595 = n8932 & n8933;
  assign n2596 = ~n8930 & ~n8931;
  assign n2597 = n8930 & ~n8931;
  assign n2598 = ~n8930 & n8931;
  assign n2599 = ~n2597 & ~n2598;
  assign n2600 = ~n2576 & ~n2596;
  assign n2601 = n2595 & ~n8934;
  assign n2602 = ~n2576 & ~n2601;
  assign n2603 = ~n8767 & ~n8893;
  assign n2604 = n8818 & ~n2603;
  assign n2605 = ~n8767 & n8894;
  assign n2606 = ~n1325 & n8893;
  assign n2607 = ~n2605 & ~n2606;
  assign n2608 = n8767 & n2299;
  assign n2609 = n1325 & ~n8818;
  assign n2610 = n8893 & ~n2609;
  assign n2611 = ~n2608 & ~n2610;
  assign n2612 = ~n2605 & n2611;
  assign n2613 = ~n2604 & n2607;
  assign n2614 = ~n8725 & n8870;
  assign n2615 = n8725 & n8862;
  assign n2616 = ~n2614 & ~n2615;
  assign n2617 = ~n997 & n2039;
  assign n2618 = n997 & n2101;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = ~n2615 & n2619;
  assign n2621 = ~n2614 & n2620;
  assign n2622 = n2616 & n2619;
  assign n2623 = n8935 & n8936;
  assign n2624 = ~n8935 & ~n8936;
  assign n2625 = n8935 & ~n8936;
  assign n2626 = ~n8935 & n8936;
  assign n2627 = ~n2625 & ~n2626;
  assign n2628 = ~n2623 & ~n2624;
  assign n2629 = ~n8620 & n8782;
  assign n2630 = n8620 & n8783;
  assign n2631 = ~n2629 & ~n2630;
  assign n2632 = ~n66 & n8784;
  assign n2633 = n66 & n1433;
  assign n2634 = ~n2632 & ~n2633;
  assign n2635 = ~n2630 & n2634;
  assign n2636 = ~n2629 & n2635;
  assign n2637 = n2631 & n2634;
  assign n2638 = ~n8937 & n8938;
  assign n2639 = ~n2623 & ~n2638;
  assign n2640 = ~n2602 & ~n2639;
  assign n2641 = n2602 & n2639;
  assign n2642 = ~n2602 & ~n2640;
  assign n2643 = ~n2602 & n2639;
  assign n2644 = ~n2639 & ~n2640;
  assign n2645 = n2602 & ~n2639;
  assign n2646 = ~n8939 & ~n8940;
  assign n2647 = ~n2640 & ~n2641;
  assign n2648 = n8914 & ~n8915;
  assign n2649 = n8915 & ~n2458;
  assign n2650 = n8914 & n8915;
  assign n2651 = ~n8914 & ~n2458;
  assign n2652 = ~n8914 & ~n8915;
  assign n2653 = ~n8942 & ~n8943;
  assign n2654 = ~n2458 & ~n2648;
  assign n2655 = ~n8941 & ~n8944;
  assign n2656 = ~n2640 & ~n2655;
  assign n2657 = n2459 & ~n2461;
  assign n2658 = ~n2462 & ~n2657;
  assign n2659 = ~n2656 & n2658;
  assign n2660 = n2656 & ~n2658;
  assign n2661 = ~n2659 & ~n2660;
  assign n2662 = n8928 & ~n2541;
  assign n2663 = n2541 & ~n2542;
  assign n2664 = ~n8928 & ~n2542;
  assign n2665 = ~n2663 & ~n2664;
  assign n2666 = ~n2542 & ~n2662;
  assign n2667 = n2661 & ~n8945;
  assign n2668 = ~n2659 & ~n2667;
  assign n2669 = ~n2547 & ~n2549;
  assign n2670 = ~n2550 & ~n2669;
  assign n2671 = ~n2668 & n2670;
  assign n2672 = n2668 & ~n2670;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = ~n8622 & ~n8724;
  assign n2675 = ~n997 & n8870;
  assign n2676 = n997 & n8862;
  assign n2677 = ~n2675 & ~n2676;
  assign n2678 = n8787 & n2101;
  assign n2679 = ~n8787 & n2039;
  assign n2680 = ~n2678 & ~n2679;
  assign n2681 = ~n2676 & n2680;
  assign n2682 = ~n2675 & n2681;
  assign n2683 = n2677 & n2680;
  assign n2684 = n8765 & n1846;
  assign n2685 = n8766 & ~n1846;
  assign n2686 = ~n2684 & ~n2685;
  assign n2687 = n8620 & n1309;
  assign n2688 = ~n8620 & n8768;
  assign n2689 = ~n2687 & ~n2688;
  assign n2690 = ~n2684 & n2689;
  assign n2691 = ~n2685 & n2690;
  assign n2692 = ~n2684 & ~n2688;
  assign n2693 = ~n2685 & ~n2687;
  assign n2694 = n2692 & n2693;
  assign n2695 = n2686 & n2689;
  assign n2696 = n8946 & n8947;
  assign n2697 = ~n8946 & ~n8947;
  assign n2698 = n8946 & ~n8947;
  assign n2699 = ~n8946 & n8947;
  assign n2700 = ~n2698 & ~n2699;
  assign n2701 = ~n2696 & ~n2697;
  assign n2702 = ~n854 & n8847;
  assign n2703 = n854 & n8833;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = n8651 & n1959;
  assign n2706 = ~n8651 & n1872;
  assign n2707 = ~n2705 & ~n2706;
  assign n2708 = ~n2703 & n2707;
  assign n2709 = ~n2702 & n2708;
  assign n2710 = n2704 & n2707;
  assign n2711 = ~n8948 & n8949;
  assign n2712 = ~n2696 & ~n2711;
  assign n2713 = n8622 & n8650;
  assign n2714 = ~n992 & ~n2713;
  assign n2715 = n8650 & ~n2712;
  assign n2716 = n2714 & n2715;
  assign n2717 = n2674 & ~n2712;
  assign n2718 = ~n2595 & n8934;
  assign n2719 = ~n2601 & ~n2718;
  assign n2720 = ~n2674 & n2712;
  assign n2721 = n8650 & ~n8950;
  assign n2722 = n2714 & n2721;
  assign n2723 = ~n2712 & ~n8950;
  assign n2724 = ~n2722 & ~n2723;
  assign n2725 = ~n8950 & ~n2720;
  assign n2726 = n2719 & ~n8951;
  assign n2727 = ~n8950 & ~n2726;
  assign n2728 = n2525 & ~n2528;
  assign n2729 = n2525 & ~n2527;
  assign n2730 = ~n2523 & n8925;
  assign n2731 = ~n2525 & n2527;
  assign n2732 = ~n8952 & ~n8953;
  assign n2733 = ~n2727 & ~n2732;
  assign n2734 = n2727 & n2732;
  assign n2735 = ~n2727 & n2732;
  assign n2736 = n2727 & ~n2732;
  assign n2737 = ~n2735 & ~n2736;
  assign n2738 = ~n2733 & ~n2734;
  assign n2739 = n8941 & n8944;
  assign n2740 = ~n8941 & ~n2655;
  assign n2741 = ~n8944 & ~n2655;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = ~n2655 & ~n2739;
  assign n2744 = ~n8954 & ~n8955;
  assign n2745 = ~n2733 & ~n2744;
  assign n2746 = ~n2661 & n8945;
  assign n2747 = ~n2667 & ~n2746;
  assign n2748 = ~n2745 & n2747;
  assign n2749 = n2745 & ~n2747;
  assign n2750 = n8954 & n8955;
  assign n2751 = ~n2744 & ~n2750;
  assign n2752 = ~n2719 & n8951;
  assign n2753 = ~n8951 & ~n2726;
  assign n2754 = n2719 & ~n2726;
  assign n2755 = ~n2753 & ~n2754;
  assign n2756 = ~n2726 & ~n2752;
  assign n2757 = ~n8932 & ~n8933;
  assign n2758 = ~n2595 & ~n2757;
  assign n2759 = ~n66 & n8782;
  assign n2760 = n66 & n8783;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = n8622 & n1433;
  assign n2763 = ~n8622 & n8784;
  assign n2764 = ~n2762 & ~n2763;
  assign n2765 = ~n2760 & n2764;
  assign n2766 = ~n2759 & n2765;
  assign n2767 = n2761 & n2764;
  assign n2768 = n2758 & n8957;
  assign n2769 = ~n8725 & ~n8893;
  assign n2770 = n8818 & ~n2769;
  assign n2771 = ~n8725 & n8894;
  assign n2772 = ~n997 & n8893;
  assign n2773 = ~n2771 & ~n2772;
  assign n2774 = n8725 & n2299;
  assign n2775 = n997 & ~n8818;
  assign n2776 = n8893 & ~n2775;
  assign n2777 = ~n2774 & ~n2776;
  assign n2778 = ~n2771 & n2777;
  assign n2779 = ~n2770 & n2773;
  assign n2780 = ~n8787 & n8870;
  assign n2781 = n8787 & n8862;
  assign n2782 = ~n2780 & ~n2781;
  assign n2783 = ~n854 & n2039;
  assign n2784 = n854 & n2101;
  assign n2785 = ~n2783 & ~n2784;
  assign n2786 = ~n2781 & n2785;
  assign n2787 = ~n2780 & n2786;
  assign n2788 = n2782 & n2785;
  assign n2789 = n8958 & n8959;
  assign n2790 = ~n8958 & ~n8959;
  assign n2791 = n8958 & ~n8959;
  assign n2792 = ~n8958 & n8959;
  assign n2793 = ~n2791 & ~n2792;
  assign n2794 = ~n2789 & ~n2790;
  assign n2795 = ~n8651 & n8847;
  assign n2796 = n8651 & n8833;
  assign n2797 = ~n2795 & ~n2796;
  assign n2798 = ~n1846 & n1872;
  assign n2799 = n1846 & n1959;
  assign n2800 = ~n2798 & ~n2799;
  assign n2801 = ~n2796 & n2800;
  assign n2802 = ~n2795 & n2801;
  assign n2803 = n2797 & n2800;
  assign n2804 = ~n8960 & n8961;
  assign n2805 = ~n2789 & ~n2804;
  assign n2806 = ~n2758 & ~n8957;
  assign n2807 = ~n2758 & n8957;
  assign n2808 = n2758 & ~n8957;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = ~n2768 & ~n2806;
  assign n2811 = ~n2805 & ~n8962;
  assign n2812 = ~n2768 & ~n2811;
  assign n2813 = n8937 & ~n8938;
  assign n2814 = n8938 & ~n2638;
  assign n2815 = n8937 & n8938;
  assign n2816 = ~n8937 & ~n2638;
  assign n2817 = ~n8937 & ~n8938;
  assign n2818 = ~n8963 & ~n8964;
  assign n2819 = ~n2638 & ~n2813;
  assign n2820 = ~n2812 & ~n8965;
  assign n2821 = n2812 & n8965;
  assign n2822 = ~n2812 & ~n2820;
  assign n2823 = ~n8965 & ~n2820;
  assign n2824 = ~n2822 & ~n2823;
  assign n2825 = ~n2820 & ~n2821;
  assign n2826 = ~n8956 & ~n8966;
  assign n2827 = n8956 & n8966;
  assign n2828 = ~n2826 & ~n2827;
  assign n2829 = ~n8622 & ~n8764;
  assign n2830 = ~n8622 & n8766;
  assign n2831 = n8622 & ~n1293;
  assign n2832 = ~n1309 & ~n2831;
  assign n2833 = ~n2830 & n2832;
  assign n2834 = n1293 & n2833;
  assign n2835 = n1293 & ~n2829;
  assign n2836 = ~n997 & ~n8893;
  assign n2837 = n8818 & ~n2836;
  assign n2838 = ~n997 & n8894;
  assign n2839 = ~n8787 & n8893;
  assign n2840 = ~n2838 & ~n2839;
  assign n2841 = n997 & n2299;
  assign n2842 = n8787 & ~n8818;
  assign n2843 = n8893 & ~n2842;
  assign n2844 = ~n2841 & ~n2843;
  assign n2845 = ~n2838 & n2844;
  assign n2846 = ~n2837 & n2840;
  assign n2847 = n8967 & n8968;
  assign n2848 = n8620 & n8765;
  assign n2849 = ~n8620 & n8766;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = ~n66 & n8768;
  assign n2852 = n66 & n1309;
  assign n2853 = ~n2851 & ~n2852;
  assign n2854 = ~n2848 & n2853;
  assign n2855 = ~n2849 & n2854;
  assign n2856 = ~n2848 & ~n2851;
  assign n2857 = ~n2849 & ~n2852;
  assign n2858 = n2856 & n2857;
  assign n2859 = n2850 & n2853;
  assign n2860 = n2847 & n8969;
  assign n2861 = ~n2847 & ~n8969;
  assign n2862 = n2847 & ~n8969;
  assign n2863 = ~n2847 & n8969;
  assign n2864 = ~n2862 & ~n2863;
  assign n2865 = ~n2860 & ~n2861;
  assign n2866 = n2577 & ~n8970;
  assign n2867 = ~n2860 & ~n2866;
  assign n2868 = n8948 & ~n8949;
  assign n2869 = ~n2711 & ~n2868;
  assign n2870 = ~n2867 & n2869;
  assign n2871 = n2867 & ~n2869;
  assign n2872 = ~n2870 & ~n2871;
  assign n2873 = n2805 & n8962;
  assign n2874 = ~n2811 & ~n2873;
  assign n2875 = n2872 & n2874;
  assign n2876 = ~n2872 & ~n2874;
  assign n2877 = ~n2875 & ~n2876;
  assign n2878 = ~n2577 & n8970;
  assign n2879 = ~n2866 & ~n2878;
  assign n2880 = ~n854 & n8870;
  assign n2881 = n854 & n8862;
  assign n2882 = ~n2880 & ~n2881;
  assign n2883 = n8651 & n2101;
  assign n2884 = ~n8651 & n2039;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = ~n2881 & n2885;
  assign n2887 = ~n2880 & n2886;
  assign n2888 = n2882 & n2885;
  assign n2889 = ~n1846 & n8847;
  assign n2890 = n1846 & n8833;
  assign n2891 = ~n2889 & ~n2890;
  assign n2892 = n8620 & n1959;
  assign n2893 = ~n8620 & n1872;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = ~n2890 & n2894;
  assign n2896 = ~n2889 & n2895;
  assign n2897 = n2891 & n2894;
  assign n2898 = n8971 & n8972;
  assign n2899 = ~n8971 & ~n8972;
  assign n2900 = n8971 & ~n8972;
  assign n2901 = ~n8971 & n8972;
  assign n2902 = ~n2900 & ~n2901;
  assign n2903 = ~n2898 & ~n2899;
  assign n2904 = n66 & n8765;
  assign n2905 = ~n66 & n8766;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = n8622 & n1309;
  assign n2908 = ~n8622 & n8768;
  assign n2909 = ~n2907 & ~n2908;
  assign n2910 = ~n2904 & n2909;
  assign n2911 = ~n2905 & n2910;
  assign n2912 = ~n2905 & ~n2908;
  assign n2913 = ~n2904 & ~n2907;
  assign n2914 = n2912 & n2913;
  assign n2915 = n2906 & n2909;
  assign n2916 = ~n8973 & n8974;
  assign n2917 = ~n2898 & ~n2916;
  assign n2918 = n8960 & ~n8961;
  assign n2919 = ~n2804 & ~n2918;
  assign n2920 = ~n2917 & n2919;
  assign n2921 = n2917 & ~n2919;
  assign n2922 = ~n2917 & ~n2920;
  assign n2923 = n2919 & ~n2920;
  assign n2924 = ~n2922 & ~n2923;
  assign n2925 = ~n2920 & ~n2921;
  assign n2926 = n2879 & ~n8975;
  assign n2927 = ~n2879 & n8975;
  assign n2928 = ~n2926 & ~n2927;
  assign n2929 = ~n8967 & ~n8968;
  assign n2930 = ~n2847 & ~n2929;
  assign n2931 = ~n8787 & ~n8893;
  assign n2932 = n8818 & ~n2931;
  assign n2933 = ~n8787 & n8894;
  assign n2934 = ~n854 & n8893;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = n8787 & n2299;
  assign n2937 = n854 & ~n8818;
  assign n2938 = n8893 & ~n2937;
  assign n2939 = ~n2936 & ~n2938;
  assign n2940 = ~n2933 & n2939;
  assign n2941 = ~n2932 & n2935;
  assign n2942 = ~n8651 & n8870;
  assign n2943 = n8651 & n8862;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = ~n1846 & n2039;
  assign n2946 = n1846 & n2101;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = ~n2943 & n2947;
  assign n2949 = ~n2942 & n2948;
  assign n2950 = n2944 & n2947;
  assign n2951 = n8976 & n8977;
  assign n2952 = ~n8976 & ~n8977;
  assign n2953 = n8976 & ~n8977;
  assign n2954 = ~n8976 & n8977;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = ~n2951 & ~n2952;
  assign n2957 = ~n8620 & n8847;
  assign n2958 = n8620 & n8833;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = ~n66 & n1872;
  assign n2961 = n66 & n1959;
  assign n2962 = ~n2960 & ~n2961;
  assign n2963 = ~n2958 & n2962;
  assign n2964 = ~n2957 & n2963;
  assign n2965 = n2959 & n2962;
  assign n2966 = ~n8978 & n8979;
  assign n2967 = ~n2951 & ~n2966;
  assign n2968 = n2930 & ~n2967;
  assign n2969 = ~n2930 & n2967;
  assign n2970 = ~n2968 & ~n2969;
  assign n2971 = n8973 & ~n8974;
  assign n2972 = n8974 & ~n2916;
  assign n2973 = n8973 & n8974;
  assign n2974 = ~n8973 & ~n2916;
  assign n2975 = ~n8973 & ~n8974;
  assign n2976 = ~n8980 & ~n8981;
  assign n2977 = ~n2916 & ~n2971;
  assign n2978 = n2970 & ~n8982;
  assign n2979 = ~n2970 & n8982;
  assign n2980 = ~n2978 & ~n2979;
  assign n2981 = ~n8622 & ~n8832;
  assign n2982 = ~n8622 & n8847;
  assign n2983 = n8622 & ~n846;
  assign n2984 = ~n1959 & ~n2983;
  assign n2985 = ~n2982 & n2984;
  assign n2986 = n846 & n2985;
  assign n2987 = n846 & ~n2981;
  assign n2988 = ~n854 & ~n8893;
  assign n2989 = n8818 & ~n2988;
  assign n2990 = ~n854 & n8894;
  assign n2991 = ~n8651 & n8893;
  assign n2992 = ~n2990 & ~n2991;
  assign n2993 = n854 & n2299;
  assign n2994 = n8651 & ~n8818;
  assign n2995 = n8893 & ~n2994;
  assign n2996 = ~n2993 & ~n2995;
  assign n2997 = ~n2990 & n2996;
  assign n2998 = ~n2989 & n2992;
  assign n2999 = n8983 & n8984;
  assign n3000 = ~n8967 & n2999;
  assign n3001 = n2832 & n3000;
  assign n3002 = n2829 & n2999;
  assign n3003 = ~n2829 & ~n2999;
  assign n3004 = n2999 & ~n8985;
  assign n3005 = ~n2829 & n2999;
  assign n3006 = ~n8967 & ~n8985;
  assign n3007 = n2832 & n3006;
  assign n3008 = n2829 & ~n2999;
  assign n3009 = ~n8986 & ~n8987;
  assign n3010 = ~n8985 & ~n3003;
  assign n3011 = ~n1846 & n8870;
  assign n3012 = n1846 & n8862;
  assign n3013 = ~n3011 & ~n3012;
  assign n3014 = n8620 & n2101;
  assign n3015 = ~n8620 & n2039;
  assign n3016 = ~n3014 & ~n3015;
  assign n3017 = ~n3012 & n3016;
  assign n3018 = ~n3011 & n3017;
  assign n3019 = n3013 & n3016;
  assign n3020 = ~n66 & n8847;
  assign n3021 = n66 & n8833;
  assign n3022 = ~n3020 & ~n3021;
  assign n3023 = ~n8622 & n1872;
  assign n3024 = n8622 & n1959;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = ~n3021 & n3025;
  assign n3027 = ~n3020 & n3026;
  assign n3028 = n3022 & n3025;
  assign n3029 = n8989 & n8990;
  assign n3030 = ~n8983 & ~n8984;
  assign n3031 = ~n2999 & ~n3030;
  assign n3032 = ~n8989 & ~n8990;
  assign n3033 = n3031 & ~n3032;
  assign n3034 = ~n3029 & ~n3032;
  assign n3035 = n3031 & n3034;
  assign n3036 = ~n3029 & ~n3035;
  assign n3037 = ~n3029 & ~n3033;
  assign n3038 = ~n8988 & ~n8991;
  assign n3039 = n8988 & n8991;
  assign n3040 = ~n8991 & ~n3038;
  assign n3041 = ~n8988 & ~n3038;
  assign n3042 = ~n3040 & ~n3041;
  assign n3043 = ~n3038 & ~n3039;
  assign n3044 = n8978 & ~n8979;
  assign n3045 = ~n2966 & ~n3044;
  assign n3046 = ~n8992 & n3045;
  assign n3047 = n8992 & ~n3045;
  assign n3048 = ~n8651 & n8894;
  assign n3049 = ~n8818 & n1846;
  assign n3050 = n8893 & ~n3049;
  assign n3051 = n8651 & n8818;
  assign n3052 = n8651 & n2299;
  assign n3053 = ~n3050 & ~n3052;
  assign n3054 = ~n3050 & ~n3051;
  assign n3055 = ~n3048 & n8993;
  assign n3056 = ~n8620 & n8870;
  assign n3057 = n8620 & n8862;
  assign n3058 = ~n3056 & ~n3057;
  assign n3059 = n66 & n2101;
  assign n3060 = ~n66 & n2039;
  assign n3061 = ~n3059 & ~n3060;
  assign n3062 = ~n3057 & n3061;
  assign n3063 = ~n3056 & n3062;
  assign n3064 = n3058 & n3061;
  assign n3065 = n3055 & n8994;
  assign n3066 = ~n8622 & ~n8861;
  assign n3067 = ~n8622 & n8870;
  assign n3068 = n8622 & ~n1840;
  assign n3069 = ~n2101 & ~n3068;
  assign n3070 = ~n3067 & n3069;
  assign n3071 = n1840 & n3070;
  assign n3072 = n1840 & ~n3066;
  assign n3073 = n8620 & ~n8818;
  assign n3074 = n8893 & ~n3073;
  assign n3075 = ~n1846 & ~n8894;
  assign n3076 = ~n3049 & ~n3075;
  assign n3077 = ~n1846 & n8894;
  assign n3078 = n1846 & n2299;
  assign n3079 = ~n3074 & ~n3078;
  assign n3080 = ~n3077 & n3079;
  assign n3081 = ~n3074 & ~n3076;
  assign n3082 = n8995 & n8996;
  assign n3083 = ~n3055 & ~n8994;
  assign n3084 = n3055 & ~n8994;
  assign n3085 = ~n3055 & n8994;
  assign n3086 = ~n3084 & ~n3085;
  assign n3087 = ~n3065 & ~n3083;
  assign n3088 = n3082 & ~n8997;
  assign n3089 = ~n3065 & ~n3088;
  assign n3090 = n3031 & ~n3035;
  assign n3091 = n3031 & ~n3034;
  assign n3092 = ~n3032 & n8991;
  assign n3093 = ~n3031 & n3034;
  assign n3094 = ~n8998 & ~n8999;
  assign n3095 = ~n3089 & ~n3094;
  assign n3096 = n3089 & n3094;
  assign n3097 = ~n8995 & ~n8996;
  assign n3098 = ~n3082 & ~n3097;
  assign n3099 = ~n66 & ~n8893;
  assign n3100 = n8622 & ~n8818;
  assign n3101 = ~n3099 & n3100;
  assign n3102 = ~n3066 & ~n3101;
  assign n3103 = ~n8620 & n8818;
  assign n3104 = ~n3073 & ~n3103;
  assign n3105 = ~n8893 & ~n3104;
  assign n3106 = n66 & ~n8818;
  assign n3107 = n8893 & n3106;
  assign n3108 = ~n8620 & n8894;
  assign n3109 = n8818 & n8893;
  assign n3110 = n66 & ~n3109;
  assign n3111 = ~n3099 & ~n3110;
  assign n3112 = n8893 & ~n3106;
  assign n3113 = n8620 & n2299;
  assign n3114 = ~n9000 & ~n3113;
  assign n3115 = ~n3108 & n3114;
  assign n3116 = ~n8893 & ~n3073;
  assign n3117 = ~n3103 & n3116;
  assign n3118 = ~n9000 & ~n3117;
  assign n3119 = ~n3105 & ~n3107;
  assign n3120 = ~n3101 & ~n9001;
  assign n3121 = ~n8995 & ~n3120;
  assign n3122 = n3069 & n3121;
  assign n3123 = n3066 & n9001;
  assign n3124 = n3101 & n9001;
  assign n3125 = ~n9002 & ~n3124;
  assign n3126 = ~n3101 & ~n9002;
  assign n3127 = ~n3066 & ~n9001;
  assign n3128 = ~n3126 & ~n3127;
  assign n3129 = ~n3102 & n9001;
  assign n3130 = ~n3098 & n9003;
  assign n3131 = n3098 & ~n9003;
  assign n3132 = ~n66 & n8870;
  assign n3133 = n66 & n8862;
  assign n3134 = ~n3132 & ~n3133;
  assign n3135 = n8622 & n2101;
  assign n3136 = ~n8622 & n2039;
  assign n3137 = ~n3135 & ~n3136;
  assign n3138 = n3134 & n3137;
  assign n3139 = ~n3131 & ~n3138;
  assign n3140 = ~n3130 & ~n3135;
  assign n3141 = ~n3136 & n3140;
  assign n3142 = ~n3133 & n3141;
  assign n3143 = ~n3132 & n3142;
  assign n3144 = ~n3131 & ~n3143;
  assign n3145 = ~n3130 & ~n3139;
  assign n3146 = n2981 & ~n9004;
  assign n3147 = ~n2981 & n9004;
  assign n3148 = ~n3082 & n8997;
  assign n3149 = ~n3088 & ~n3148;
  assign n3150 = ~n3088 & ~n3147;
  assign n3151 = ~n3148 & n3150;
  assign n3152 = ~n3147 & n3149;
  assign n3153 = ~n3146 & ~n9005;
  assign n3154 = ~n3096 & ~n3153;
  assign n3155 = n3094 & n3153;
  assign n3156 = ~n3089 & ~n3155;
  assign n3157 = ~n3094 & ~n3153;
  assign n3158 = ~n3156 & ~n3157;
  assign n3159 = ~n3095 & ~n3154;
  assign n3160 = ~n3047 & ~n9006;
  assign n3161 = ~n8992 & ~n9006;
  assign n3162 = n8992 & n9006;
  assign n3163 = ~n2966 & ~n3162;
  assign n3164 = ~n3044 & n3163;
  assign n3165 = ~n3161 & ~n3164;
  assign n3166 = ~n3045 & ~n3161;
  assign n3167 = ~n3162 & ~n3166;
  assign n3168 = ~n3046 & ~n3160;
  assign n3169 = n2980 & ~n9007;
  assign n3170 = ~n8985 & ~n3038;
  assign n3171 = ~n2980 & n9007;
  assign n3172 = ~n3170 & ~n3171;
  assign n3173 = ~n9007 & ~n3170;
  assign n3174 = n9007 & n3170;
  assign n3175 = n2980 & ~n3174;
  assign n3176 = ~n3173 & ~n3175;
  assign n3177 = ~n2980 & ~n3173;
  assign n3178 = ~n3174 & ~n3177;
  assign n3179 = ~n3169 & ~n3172;
  assign n3180 = n2928 & ~n9008;
  assign n3181 = ~n2968 & ~n2978;
  assign n3182 = ~n2928 & n9008;
  assign n3183 = ~n3181 & ~n3182;
  assign n3184 = ~n9008 & ~n3181;
  assign n3185 = n9008 & n3181;
  assign n3186 = n2928 & ~n3185;
  assign n3187 = ~n3184 & ~n3186;
  assign n3188 = ~n2928 & ~n3184;
  assign n3189 = ~n3185 & ~n3188;
  assign n3190 = ~n3180 & ~n3183;
  assign n3191 = n2877 & ~n9009;
  assign n3192 = ~n2920 & ~n2926;
  assign n3193 = ~n2877 & n9009;
  assign n3194 = ~n3192 & ~n3193;
  assign n3195 = ~n9009 & ~n3192;
  assign n3196 = n9009 & n3192;
  assign n3197 = ~n2875 & ~n3196;
  assign n3198 = ~n2876 & n3197;
  assign n3199 = ~n3195 & ~n3198;
  assign n3200 = ~n2877 & ~n3195;
  assign n3201 = ~n3196 & ~n3200;
  assign n3202 = ~n3191 & ~n3194;
  assign n3203 = n2828 & ~n9010;
  assign n3204 = ~n2870 & ~n2875;
  assign n3205 = ~n2828 & n9010;
  assign n3206 = ~n3204 & ~n3205;
  assign n3207 = ~n9010 & ~n3204;
  assign n3208 = n9010 & n3204;
  assign n3209 = n2828 & ~n3208;
  assign n3210 = ~n3207 & ~n3209;
  assign n3211 = ~n2828 & ~n3207;
  assign n3212 = ~n3208 & ~n3211;
  assign n3213 = ~n3203 & ~n3206;
  assign n3214 = n2751 & ~n9011;
  assign n3215 = ~n2820 & ~n2826;
  assign n3216 = ~n2751 & n9011;
  assign n3217 = ~n3215 & ~n3216;
  assign n3218 = ~n9011 & ~n3215;
  assign n3219 = n9011 & n3215;
  assign n3220 = ~n2750 & ~n3219;
  assign n3221 = ~n2744 & n3220;
  assign n3222 = ~n3218 & ~n3221;
  assign n3223 = ~n2751 & ~n3218;
  assign n3224 = ~n3219 & ~n3223;
  assign n3225 = ~n3214 & ~n3217;
  assign n3226 = ~n2749 & ~n9012;
  assign n3227 = ~n2748 & ~n2749;
  assign n3228 = ~n9012 & n3227;
  assign n3229 = ~n2748 & ~n3228;
  assign n3230 = ~n2748 & n9012;
  assign n3231 = ~n2749 & ~n3230;
  assign n3232 = ~n2748 & ~n3226;
  assign n3233 = n2673 & ~n9013;
  assign n3234 = ~n2671 & ~n3233;
  assign n3235 = n2551 & ~n2553;
  assign n3236 = ~n2554 & ~n3235;
  assign n3237 = ~n3234 & n3236;
  assign n3238 = ~n2554 & ~n3237;
  assign n3239 = n2495 & ~n2497;
  assign n3240 = ~n2498 & ~n3239;
  assign n3241 = ~n3238 & n3240;
  assign n3242 = ~n2498 & ~n3241;
  assign n3243 = n2390 & n8908;
  assign n3244 = ~n2390 & n8908;
  assign n3245 = n2390 & ~n8908;
  assign n3246 = ~n3244 & ~n3245;
  assign n3247 = ~n2398 & ~n3243;
  assign n3248 = ~n3242 & ~n9014;
  assign n3249 = ~n2398 & ~n3248;
  assign n3250 = n2183 & n2186;
  assign n3251 = ~n2187 & ~n3250;
  assign n3252 = ~n3249 & n3251;
  assign n3253 = ~n2187 & ~n3252;
  assign n3254 = n8842 & n8857;
  assign n3255 = ~n8842 & ~n2004;
  assign n3256 = ~n8857 & ~n2004;
  assign n3257 = ~n3255 & ~n3256;
  assign n3258 = ~n2004 & ~n3254;
  assign n3259 = ~n3253 & ~n9015;
  assign n3260 = ~n2004 & ~n3259;
  assign n3261 = n1920 & ~n1922;
  assign n3262 = ~n1923 & ~n3261;
  assign n3263 = ~n3260 & n3262;
  assign n3264 = ~n1923 & ~n3263;
  assign n3265 = n1532 & n8804;
  assign n3266 = ~n1532 & n8804;
  assign n3267 = n1532 & ~n8804;
  assign n3268 = ~n3266 & ~n3267;
  assign n3269 = ~n1574 & ~n3265;
  assign n3270 = ~n3264 & ~n9016;
  assign n3271 = ~n1574 & ~n3270;
  assign n3272 = ~n1558 & ~n1566;
  assign n3273 = ~n1539 & ~n1553;
  assign n3274 = n992 & n8767;
  assign n3275 = n987 & ~n8767;
  assign n3276 = ~n8650 & n1021;
  assign n3277 = n8650 & ~n1021;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = ~n8724 & n1021;
  assign n3280 = ~n8724 & n3278;
  assign n3281 = ~n3275 & ~n9017;
  assign n3282 = ~n3274 & ~n3275;
  assign n3283 = ~n9017 & n3282;
  assign n3284 = ~n3274 & n3281;
  assign n3285 = ~n3273 & n9018;
  assign n3286 = n3273 & ~n9018;
  assign n3287 = ~n3285 & ~n3286;
  assign n3288 = ~n1006 & ~n1428;
  assign n3289 = n1507 & n3288;
  assign n3290 = ~n1507 & ~n3288;
  assign n3291 = ~n3289 & ~n3290;
  assign n3292 = n3287 & n3291;
  assign n3293 = ~n3287 & ~n3291;
  assign n3294 = ~n3292 & ~n3293;
  assign n3295 = ~n3272 & n3294;
  assign n3296 = n3272 & ~n3294;
  assign n3297 = ~n3295 & ~n3296;
  assign n3298 = ~n3271 & n3297;
  assign n3299 = n3271 & ~n3297;
  assign n3300 = ~n3298 & ~n3299;
  assign n3301 = n609 & n703;
  assign n3302 = ~n430 & ~n480;
  assign n3303 = n1392 & n3302;
  assign n3304 = n3301 & n3303;
  assign n3305 = ~n8663 & ~n967;
  assign n3306 = ~n865 & n3305;
  assign n3307 = n8683 & n3306;
  assign n3308 = n8658 & n8755;
  assign n3309 = n3307 & n3308;
  assign n3310 = ~n430 & ~n8663;
  assign n3311 = n609 & n3310;
  assign n3312 = n703 & n1392;
  assign n3313 = n3311 & n3312;
  assign n3314 = ~n480 & ~n865;
  assign n3315 = ~n967 & n3314;
  assign n3316 = n8658 & n3315;
  assign n3317 = n8683 & n8755;
  assign n3318 = n3316 & n3317;
  assign n3319 = n3313 & n3318;
  assign n3320 = n3304 & n3309;
  assign n3321 = n8680 & n8771;
  assign n3322 = n9019 & n3321;
  assign n3323 = n703 & n8755;
  assign n3324 = n8683 & n3323;
  assign n3325 = n609 & n3324;
  assign n3326 = n1392 & n3325;
  assign n3327 = n8658 & n3326;
  assign n3328 = n8680 & n3327;
  assign n3329 = n8771 & n3328;
  assign n3330 = n8812 & n3329;
  assign n3331 = ~n865 & n3330;
  assign n3332 = ~n430 & n3331;
  assign n3333 = ~n967 & n3332;
  assign n3334 = ~n8663 & n3333;
  assign n3335 = ~n480 & n3334;
  assign n3336 = n8812 & n3322;
  assign n3337 = ~n3300 & ~n9020;
  assign n3338 = n3264 & n9016;
  assign n3339 = ~n3270 & ~n3338;
  assign n3340 = ~n362 & ~n434;
  assign n3341 = ~n8664 & n3340;
  assign n3342 = ~n474 & ~n721;
  assign n3343 = n701 & n3342;
  assign n3344 = ~n474 & n701;
  assign n3345 = ~n8664 & n3344;
  assign n3346 = ~n362 & n3345;
  assign n3347 = ~n721 & n3346;
  assign n3348 = ~n434 & n3347;
  assign n3349 = ~n362 & ~n474;
  assign n3350 = ~n721 & n3349;
  assign n3351 = ~n434 & ~n8664;
  assign n3352 = n701 & n3351;
  assign n3353 = n3350 & n3352;
  assign n3354 = n3341 & n3343;
  assign n3355 = ~n228 & ~n8645;
  assign n3356 = ~n197 & ~n448;
  assign n3357 = n3355 & n3356;
  assign n3358 = n8774 & n3357;
  assign n3359 = n8734 & n3358;
  assign n3360 = n8734 & n8774;
  assign n3361 = n9021 & n3360;
  assign n3362 = ~n8645 & n3361;
  assign n3363 = ~n197 & n3362;
  assign n3364 = ~n228 & n3363;
  assign n3365 = ~n448 & n3364;
  assign n3366 = n9021 & n3359;
  assign n3367 = ~n251 & ~n342;
  assign n3368 = ~n342 & ~n613;
  assign n3369 = ~n251 & n3368;
  assign n3370 = ~n613 & n3367;
  assign n3371 = ~n339 & ~n431;
  assign n3372 = n1392 & n3371;
  assign n3373 = n9023 & n3372;
  assign n3374 = ~n386 & ~n938;
  assign n3375 = n654 & ~n938;
  assign n3376 = ~n386 & n3375;
  assign n3377 = n654 & n3374;
  assign n3378 = ~n8631 & ~n8637;
  assign n3379 = ~n8637 & ~n542;
  assign n3380 = ~n8631 & n3379;
  assign n3381 = ~n542 & n3378;
  assign n3382 = n9024 & n9025;
  assign n3383 = n3373 & n3382;
  assign n3384 = ~n158 & ~n8642;
  assign n3385 = ~n414 & ~n642;
  assign n3386 = n1233 & n3385;
  assign n3387 = n3384 & n3386;
  assign n3388 = n8733 & n3387;
  assign n3389 = n9023 & n9024;
  assign n3390 = n3385 & n3389;
  assign n3391 = n1233 & n3390;
  assign n3392 = n1392 & n3391;
  assign n3393 = n9025 & n3392;
  assign n3394 = n8733 & n3393;
  assign n3395 = ~n8642 & n3394;
  assign n3396 = ~n339 & n3395;
  assign n3397 = ~n158 & n3396;
  assign n3398 = ~n431 & n3397;
  assign n3399 = n1233 & n3371;
  assign n3400 = n9024 & n3399;
  assign n3401 = n9023 & n9025;
  assign n3402 = n3400 & n3401;
  assign n3403 = n1392 & n3384;
  assign n3404 = n3385 & n3403;
  assign n3405 = n8733 & n3404;
  assign n3406 = n3402 & n3405;
  assign n3407 = n3383 & n3388;
  assign n3408 = ~n288 & ~n398;
  assign n3409 = ~n288 & ~n469;
  assign n3410 = ~n398 & n3409;
  assign n3411 = ~n469 & n3408;
  assign n3412 = ~n313 & ~n417;
  assign n3413 = ~n417 & ~n513;
  assign n3414 = ~n313 & n3413;
  assign n3415 = ~n513 & n3412;
  assign n3416 = ~n223 & n1119;
  assign n3417 = n9028 & n3416;
  assign n3418 = n9027 & n3416;
  assign n3419 = n9028 & n3418;
  assign n3420 = n9027 & n3417;
  assign n3421 = ~n340 & ~n1073;
  assign n3422 = n905 & n1403;
  assign n3423 = n3421 & n3422;
  assign n3424 = n8731 & n3423;
  assign n3425 = n9029 & n3424;
  assign n3426 = n9026 & n3425;
  assign n3427 = n905 & n9027;
  assign n3428 = n9028 & n3427;
  assign n3429 = n1119 & n3428;
  assign n3430 = n8731 & n3429;
  assign n3431 = n1403 & n3430;
  assign n3432 = n9022 & n3431;
  assign n3433 = n9026 & n3432;
  assign n3434 = ~n340 & n3433;
  assign n3435 = ~n223 & n3434;
  assign n3436 = ~n1073 & n3435;
  assign n3437 = n9022 & n3426;
  assign n3438 = ~n3339 & ~n9030;
  assign n3439 = n3260 & ~n3262;
  assign n3440 = ~n3263 & ~n3439;
  assign n3441 = ~n393 & ~n8686;
  assign n3442 = ~n8630 & ~n393;
  assign n3443 = ~n8686 & n3442;
  assign n3444 = ~n8630 & n3441;
  assign n3445 = ~n8630 & n9026;
  assign n3446 = ~n8686 & n3445;
  assign n3447 = ~n393 & n3446;
  assign n3448 = n9026 & n9031;
  assign n3449 = ~n492 & ~n820;
  assign n3450 = ~n625 & ~n1345;
  assign n3451 = ~n492 & ~n625;
  assign n3452 = ~n820 & ~n1345;
  assign n3453 = n3451 & n3452;
  assign n3454 = n3449 & n3450;
  assign n3455 = n1171 & n9033;
  assign n3456 = n298 & n875;
  assign n3457 = n297 & n9028;
  assign n3458 = n875 & n3457;
  assign n3459 = ~n8643 & n3458;
  assign n3460 = n9028 & n3456;
  assign n3461 = ~n8629 & n9034;
  assign n3462 = ~n240 & n3461;
  assign n3463 = ~n492 & n3462;
  assign n3464 = ~n820 & n3463;
  assign n3465 = ~n625 & n3464;
  assign n3466 = ~n1345 & n3465;
  assign n3467 = n3455 & n9034;
  assign n3468 = ~n204 & ~n641;
  assign n3469 = ~n287 & ~n865;
  assign n3470 = ~n362 & ~n823;
  assign n3471 = n3469 & n3470;
  assign n3472 = ~n362 & ~n865;
  assign n3473 = ~n287 & ~n823;
  assign n3474 = n3468 & n3473;
  assign n3475 = n3472 & n3474;
  assign n3476 = n3468 & n3471;
  assign n3477 = ~n287 & n8753;
  assign n3478 = ~n204 & n3477;
  assign n3479 = ~n865 & n3478;
  assign n3480 = ~n641 & n3479;
  assign n3481 = ~n362 & n3480;
  assign n3482 = ~n823 & n3481;
  assign n3483 = n8753 & n9036;
  assign n3484 = ~n288 & ~n633;
  assign n3485 = ~n256 & ~n280;
  assign n3486 = ~n280 & ~n633;
  assign n3487 = ~n256 & ~n288;
  assign n3488 = n3486 & n3487;
  assign n3489 = n3484 & n3485;
  assign n3490 = n567 & n816;
  assign n3491 = n9038 & n3490;
  assign n3492 = ~n387 & ~n480;
  assign n3493 = ~n387 & ~n8664;
  assign n3494 = ~n480 & n3493;
  assign n3495 = ~n480 & ~n8664;
  assign n3496 = ~n387 & n3495;
  assign n3497 = ~n8664 & n3492;
  assign n3498 = n8887 & n9039;
  assign n3499 = n3491 & n3498;
  assign n3500 = n9037 & n3499;
  assign n3501 = n9035 & n3500;
  assign n3502 = n8887 & n9032;
  assign n3503 = n9039 & n3502;
  assign n3504 = n816 & n3503;
  assign n3505 = n9037 & n3504;
  assign n3506 = n9035 & n3505;
  assign n3507 = n567 & n3506;
  assign n3508 = ~n256 & n3507;
  assign n3509 = ~n8709 & n3508;
  assign n3510 = ~n280 & n3509;
  assign n3511 = ~n8678 & n3510;
  assign n3512 = ~n288 & n3511;
  assign n3513 = n9032 & n3501;
  assign n3514 = ~n3440 & ~n9040;
  assign n3515 = n3253 & n9015;
  assign n3516 = ~n3259 & ~n3515;
  assign n3517 = ~n433 & ~n1163;
  assign n3518 = ~n433 & n8691;
  assign n3519 = ~n1163 & n3518;
  assign n3520 = n8691 & n3517;
  assign n3521 = ~n166 & ~n493;
  assign n3522 = ~n544 & ~n865;
  assign n3523 = n3521 & n3522;
  assign n3524 = n300 & n1403;
  assign n3525 = ~n295 & ~n8664;
  assign n3526 = n1642 & n3525;
  assign n3527 = n3524 & n3526;
  assign n3528 = n300 & n3522;
  assign n3529 = n1403 & n1642;
  assign n3530 = n3521 & n3525;
  assign n3531 = n3529 & n3530;
  assign n3532 = n3528 & n3531;
  assign n3533 = n3523 & n3527;
  assign n3534 = n300 & n1642;
  assign n3535 = n8703 & n3534;
  assign n3536 = n1403 & n3535;
  assign n3537 = n3521 & n3536;
  assign n3538 = ~n295 & n3537;
  assign n3539 = ~n865 & n3538;
  assign n3540 = ~n8664 & n3539;
  assign n3541 = ~n544 & n3540;
  assign n3542 = n8703 & n9042;
  assign n3543 = ~n391 & ~n876;
  assign n3544 = ~n279 & ~n445;
  assign n3545 = ~n656 & n3544;
  assign n3546 = ~n876 & n3544;
  assign n3547 = ~n391 & n3546;
  assign n3548 = ~n656 & n3547;
  assign n3549 = ~n656 & n3543;
  assign n3550 = n3544 & n3549;
  assign n3551 = n3543 & n3545;
  assign n3552 = ~n212 & ~n8663;
  assign n3553 = n643 & n3552;
  assign n3554 = n2247 & n3355;
  assign n3555 = ~n212 & ~n8645;
  assign n3556 = ~n228 & n3555;
  assign n3557 = ~n443 & n3556;
  assign n3558 = ~n642 & n3557;
  assign n3559 = ~n641 & n3558;
  assign n3560 = ~n450 & n3559;
  assign n3561 = ~n8663 & n3560;
  assign n3562 = n2247 & n3552;
  assign n3563 = n643 & n3355;
  assign n3564 = n3562 & n3563;
  assign n3565 = n3553 & n3554;
  assign n3566 = ~n8631 & ~n207;
  assign n3567 = ~n331 & ~n398;
  assign n3568 = n3566 & n3567;
  assign n3569 = ~n342 & ~n382;
  assign n3570 = n874 & n3569;
  assign n3571 = ~n382 & ~n398;
  assign n3572 = ~n331 & ~n342;
  assign n3573 = n3571 & n3572;
  assign n3574 = n874 & n3566;
  assign n3575 = n3573 & n3574;
  assign n3576 = n3568 & n3570;
  assign n3577 = n9045 & n9046;
  assign n3578 = n9044 & n9046;
  assign n3579 = n9045 & n3578;
  assign n3580 = n9044 & n3577;
  assign n3581 = n9043 & n9047;
  assign n3582 = n9041 & n9044;
  assign n3583 = n9043 & n3582;
  assign n3584 = n9045 & n3583;
  assign n3585 = ~n342 & n3584;
  assign n3586 = ~n207 & n3585;
  assign n3587 = ~n331 & n3586;
  assign n3588 = ~n8631 & n3587;
  assign n3589 = ~n382 & n3588;
  assign n3590 = n874 & n3589;
  assign n3591 = ~n398 & n3590;
  assign n3592 = n9041 & n3581;
  assign n3593 = ~n3516 & ~n9048;
  assign n3594 = n3249 & ~n3251;
  assign n3595 = ~n3252 & ~n3594;
  assign n3596 = ~n490 & ~n861;
  assign n3597 = ~n448 & ~n490;
  assign n3598 = ~n861 & n3597;
  assign n3599 = ~n448 & n3596;
  assign n3600 = ~n861 & n8716;
  assign n3601 = ~n448 & n3600;
  assign n3602 = ~n490 & n3601;
  assign n3603 = n8716 & n9049;
  assign n3604 = ~n212 & ~n876;
  assign n3605 = ~n418 & ~n445;
  assign n3606 = n1634 & n3605;
  assign n3607 = n3604 & n3606;
  assign n3608 = n8693 & n3607;
  assign n3609 = n9050 & n3608;
  assign n3610 = n722 & n950;
  assign n3611 = ~n656 & ~n1163;
  assign n3612 = n763 & n3611;
  assign n3613 = n950 & n3611;
  assign n3614 = n722 & n763;
  assign n3615 = n3613 & n3614;
  assign n3616 = n3610 & n3612;
  assign n3617 = n8654 & n722;
  assign n3618 = n763 & n3617;
  assign n3619 = ~n636 & n3618;
  assign n3620 = ~n686 & n3619;
  assign n3621 = ~n1163 & n3620;
  assign n3622 = ~n656 & n3621;
  assign n3623 = n8654 & n9051;
  assign n3624 = ~n359 & ~n433;
  assign n3625 = ~n434 & n3624;
  assign n3626 = ~n359 & n435;
  assign n3627 = ~n8630 & ~n821;
  assign n3628 = n1344 & n3627;
  assign n3629 = n291 & n332;
  assign n3630 = n3628 & n3629;
  assign n3631 = n9053 & n3630;
  assign n3632 = n9052 & n3631;
  assign n3633 = n1344 & n1634;
  assign n3634 = n3604 & n3633;
  assign n3635 = n8693 & n3634;
  assign n3636 = n9050 & n3635;
  assign n3637 = n3605 & n3627;
  assign n3638 = n3629 & n3637;
  assign n3639 = n9053 & n3638;
  assign n3640 = n9052 & n3639;
  assign n3641 = n3636 & n3640;
  assign n3642 = n3609 & n3632;
  assign n3643 = n332 & n9053;
  assign n3644 = n3604 & n3643;
  assign n3645 = n1638 & n3644;
  assign n3646 = n1344 & n3645;
  assign n3647 = n291 & n3646;
  assign n3648 = n9052 & n3647;
  assign n3649 = n8672 & n3648;
  assign n3650 = n8693 & n3649;
  assign n3651 = n9050 & n3650;
  assign n3652 = ~n8630 & n3651;
  assign n3653 = ~n445 & n3652;
  assign n3654 = ~n418 & n3653;
  assign n3655 = n8672 & n9054;
  assign n3656 = ~n3595 & ~n9055;
  assign n3657 = n3242 & n9014;
  assign n3658 = ~n3248 & ~n3657;
  assign n3659 = ~n545 & ~n625;
  assign n3660 = ~n545 & n3521;
  assign n3661 = ~n625 & n3660;
  assign n3662 = n3521 & n3659;
  assign n3663 = ~n560 & ~n876;
  assign n3664 = ~n296 & ~n8647;
  assign n3665 = ~n8647 & ~n560;
  assign n3666 = ~n296 & ~n876;
  assign n3667 = n3665 & n3666;
  assign n3668 = n3663 & n3664;
  assign n3669 = n1333 & n9057;
  assign n3670 = n9056 & n3669;
  assign n3671 = n8733 & n8826;
  assign n3672 = n1333 & n9056;
  assign n3673 = n8826 & n3672;
  assign n3674 = n8733 & n3673;
  assign n3675 = ~n296 & n3674;
  assign n3676 = ~n8647 & n3675;
  assign n3677 = ~n876 & n3676;
  assign n3678 = ~n560 & n3677;
  assign n3679 = n3670 & n3671;
  assign n3680 = ~n8652 & n1119;
  assign n3681 = n1119 & n9058;
  assign n3682 = ~n8652 & n3681;
  assign n3683 = n9058 & n3680;
  assign n3684 = ~n251 & ~n552;
  assign n3685 = ~n552 & ~n1073;
  assign n3686 = ~n251 & n3685;
  assign n3687 = ~n1073 & n3684;
  assign n3688 = ~n8629 & ~n270;
  assign n3689 = ~n415 & ~n444;
  assign n3690 = n3688 & n3689;
  assign n3691 = ~n331 & ~n480;
  assign n3692 = n614 & n3691;
  assign n3693 = n3690 & n3692;
  assign n3694 = n9060 & n3693;
  assign n3695 = n9060 & n3691;
  assign n3696 = n8687 & n3695;
  assign n3697 = ~n8629 & n3696;
  assign n3698 = ~n270 & n3697;
  assign n3699 = ~n359 & n3698;
  assign n3700 = ~n613 & n3699;
  assign n3701 = ~n444 & n3700;
  assign n3702 = ~n415 & n3701;
  assign n3703 = n8687 & n3694;
  assign n3704 = ~n197 & ~n414;
  assign n3705 = ~n823 & ~n884;
  assign n3706 = n3704 & n3705;
  assign n3707 = n300 & n685;
  assign n3708 = n300 & ~n309;
  assign n3709 = ~n197 & n3708;
  assign n3710 = ~n288 & n3709;
  assign n3711 = ~n884 & n3710;
  assign n3712 = ~n823 & n3711;
  assign n3713 = ~n414 & n3712;
  assign n3714 = n3706 & n3707;
  assign n3715 = ~n339 & ~n380;
  assign n3716 = ~n341 & n3715;
  assign n3717 = ~n514 & ~n544;
  assign n3718 = ~n280 & ~n8642;
  assign n3719 = n3717 & n3718;
  assign n3720 = n385 & n3719;
  assign n3721 = ~n339 & ~n341;
  assign n3722 = ~n8642 & n3721;
  assign n3723 = ~n280 & ~n514;
  assign n3724 = ~n380 & ~n544;
  assign n3725 = n3723 & n3724;
  assign n3726 = n385 & n3725;
  assign n3727 = n3722 & n3726;
  assign n3728 = n3716 & n3720;
  assign n3729 = n9062 & n9063;
  assign n3730 = n9061 & n3729;
  assign n3731 = ~n514 & n9059;
  assign n3732 = n9061 & n3731;
  assign n3733 = n385 & n3732;
  assign n3734 = n9062 & n3733;
  assign n3735 = ~n341 & n3734;
  assign n3736 = ~n8642 & n3735;
  assign n3737 = ~n339 & n3736;
  assign n3738 = ~n280 & n3737;
  assign n3739 = ~n544 & n3738;
  assign n3740 = ~n380 & n3739;
  assign n3741 = n9059 & n3730;
  assign n3742 = ~n3658 & ~n9064;
  assign n3743 = n3238 & ~n3240;
  assign n3744 = ~n3241 & ~n3743;
  assign n3745 = ~n686 & ~n1163;
  assign n3746 = ~n560 & ~n8678;
  assign n3747 = ~n560 & ~n1163;
  assign n3748 = ~n8678 & ~n686;
  assign n3749 = n3747 & n3748;
  assign n3750 = n3745 & n3746;
  assign n3751 = n701 & n9065;
  assign n3752 = n8634 & n8737;
  assign n3753 = n9027 & n3752;
  assign n3754 = n8737 & n9027;
  assign n3755 = n701 & n3754;
  assign n3756 = n8634 & n3755;
  assign n3757 = ~n8678 & n3756;
  assign n3758 = ~n686 & n3757;
  assign n3759 = ~n1163 & n3758;
  assign n3760 = ~n560 & n3759;
  assign n3761 = n3751 & n3753;
  assign n3762 = ~n8631 & ~n642;
  assign n3763 = ~n1073 & n3762;
  assign n3764 = ~n223 & ~n817;
  assign n3765 = ~n8686 & ~n798;
  assign n3766 = n3764 & n3765;
  assign n3767 = ~n642 & ~n1073;
  assign n3768 = ~n798 & n3767;
  assign n3769 = ~n8631 & ~n817;
  assign n3770 = ~n223 & ~n8686;
  assign n3771 = n3769 & n3770;
  assign n3772 = n3768 & n3771;
  assign n3773 = n3763 & n3766;
  assign n3774 = n8668 & n9067;
  assign n3775 = ~n382 & ~n625;
  assign n3776 = n254 & n3775;
  assign n3777 = n903 & n1635;
  assign n3778 = n254 & n903;
  assign n3779 = ~n382 & n3778;
  assign n3780 = ~n821 & n3779;
  assign n3781 = ~n884 & n3780;
  assign n3782 = ~n625 & n3781;
  assign n3783 = n3776 & n3777;
  assign n3784 = ~n279 & ~n8648;
  assign n3785 = n1033 & n1120;
  assign n3786 = n3784 & n3785;
  assign n3787 = n9068 & n3786;
  assign n3788 = n3774 & n3787;
  assign n3789 = n8659 & n3788;
  assign n3790 = n1033 & n9068;
  assign n3791 = n9066 & n3790;
  assign n3792 = n8659 & n3791;
  assign n3793 = n8668 & n3792;
  assign n3794 = n1120 & n3793;
  assign n3795 = ~n279 & n3794;
  assign n3796 = ~n8631 & n3795;
  assign n3797 = ~n8648 & n3796;
  assign n3798 = ~n223 & n3797;
  assign n3799 = ~n642 & n3798;
  assign n3800 = ~n817 & n3799;
  assign n3801 = ~n1073 & n3800;
  assign n3802 = ~n798 & n3801;
  assign n3803 = ~n8686 & n3802;
  assign n3804 = n9066 & n3789;
  assign n3805 = ~n3744 & ~n9069;
  assign n3806 = n3234 & ~n3236;
  assign n3807 = ~n3237 & ~n3806;
  assign n3808 = ~n967 & n1333;
  assign n3809 = n8667 & n9039;
  assign n3810 = n3808 & n3809;
  assign n3811 = ~n823 & ~n1345;
  assign n3812 = ~n820 & n3811;
  assign n3813 = ~n721 & ~n904;
  assign n3814 = ~n721 & n3812;
  assign n3815 = ~n904 & n3814;
  assign n3816 = ~n820 & n3813;
  assign n3817 = n3811 & n3816;
  assign n3818 = n3812 & n3813;
  assign n3819 = ~n560 & n657;
  assign n3820 = ~n380 & ~n492;
  assign n3821 = ~n552 & ~n8686;
  assign n3822 = n3820 & n3821;
  assign n3823 = n3819 & n3822;
  assign n3824 = n9050 & n3823;
  assign n3825 = n9070 & n3824;
  assign n3826 = n657 & n3821;
  assign n3827 = n9070 & n3826;
  assign n3828 = n9039 & n3827;
  assign n3829 = n1333 & n3828;
  assign n3830 = n9050 & n3829;
  assign n3831 = n8667 & n3830;
  assign n3832 = ~n492 & n3831;
  assign n3833 = ~n967 & n3832;
  assign n3834 = ~n380 & n3833;
  assign n3835 = ~n560 & n3834;
  assign n3836 = ~n560 & ~n967;
  assign n3837 = n1333 & n3836;
  assign n3838 = n8667 & n3837;
  assign n3839 = n9039 & n3838;
  assign n3840 = n657 & n3820;
  assign n3841 = n3821 & n3840;
  assign n3842 = n9050 & n3841;
  assign n3843 = n9070 & n3842;
  assign n3844 = n3839 & n3843;
  assign n3845 = n3810 & n3825;
  assign n3846 = ~n295 & ~n342;
  assign n3847 = ~n412 & ~n436;
  assign n3848 = n1251 & n3847;
  assign n3849 = n3846 & n3848;
  assign n3850 = ~n255 & ~n8678;
  assign n3851 = ~n434 & n3850;
  assign n3852 = ~n222 & ~n296;
  assign n3853 = n816 & n3852;
  assign n3854 = n3851 & n3853;
  assign n3855 = n297 & n816;
  assign n3856 = n3847 & n3855;
  assign n3857 = ~n255 & ~n342;
  assign n3858 = ~n8678 & n3857;
  assign n3859 = ~n222 & ~n434;
  assign n3860 = n1251 & n3859;
  assign n3861 = n3858 & n3860;
  assign n3862 = n3856 & n3861;
  assign n3863 = n3849 & n3854;
  assign n3864 = n8670 & n9068;
  assign n3865 = n9072 & n3864;
  assign n3866 = n8685 & n8744;
  assign n3867 = n8685 & n3865;
  assign n3868 = n8744 & n3867;
  assign n3869 = n3865 & n3866;
  assign n3870 = n297 & n1251;
  assign n3871 = n3847 & n3870;
  assign n3872 = n9068 & n3871;
  assign n3873 = n816 & n3872;
  assign n3874 = n8685 & n3873;
  assign n3875 = n8670 & n3874;
  assign n3876 = n9071 & n3875;
  assign n3877 = n8744 & n3876;
  assign n3878 = ~n342 & n3877;
  assign n3879 = ~n255 & n3878;
  assign n3880 = ~n222 & n3879;
  assign n3881 = ~n8678 & n3880;
  assign n3882 = ~n434 & n3881;
  assign n3883 = n9071 & n9073;
  assign n3884 = ~n3807 & ~n9074;
  assign n3885 = ~n2673 & n9013;
  assign n3886 = ~n3233 & ~n3885;
  assign n3887 = ~n180 & ~n544;
  assign n3888 = ~n1073 & n3887;
  assign n3889 = ~n8630 & n1643;
  assign n3890 = ~n8645 & n3889;
  assign n3891 = ~n544 & n3890;
  assign n3892 = ~n1073 & n3891;
  assign n3893 = n1643 & n3888;
  assign n3894 = ~n309 & ~n938;
  assign n3895 = ~n256 & ~n545;
  assign n3896 = ~n384 & n3895;
  assign n3897 = ~n256 & ~n309;
  assign n3898 = ~n545 & n3897;
  assign n3899 = ~n938 & n3898;
  assign n3900 = ~n384 & n3899;
  assign n3901 = ~n384 & ~n545;
  assign n3902 = ~n938 & n3897;
  assign n3903 = n3901 & n3902;
  assign n3904 = n3894 & n3896;
  assign n3905 = n211 & n378;
  assign n3906 = ~n8709 & ~n3905;
  assign n3907 = ~n492 & ~n865;
  assign n3908 = ~n492 & ~n3905;
  assign n3909 = ~n865 & ~n8709;
  assign n3910 = n3908 & n3909;
  assign n3911 = n3906 & n3907;
  assign n3912 = n9076 & n9077;
  assign n3913 = n9075 & n9076;
  assign n3914 = ~n8709 & n3913;
  assign n3915 = ~n865 & n3914;
  assign n3916 = ~n492 & n3915;
  assign n3917 = ~n387 & n3916;
  assign n3918 = ~n610 & n3917;
  assign n3919 = n9075 & n9077;
  assign n3920 = n9076 & n3919;
  assign n3921 = n9075 & n3912;
  assign n3922 = ~n8637 & ~n8640;
  assign n3923 = ~n295 & ~n8700;
  assign n3924 = n3922 & n3923;
  assign n3925 = n609 & n3821;
  assign n3926 = n3924 & n3925;
  assign n3927 = ~n228 & n576;
  assign n3928 = ~n398 & ~n641;
  assign n3929 = ~n884 & n3928;
  assign n3930 = n8760 & n3929;
  assign n3931 = n3927 & n3930;
  assign n3932 = ~n295 & ~n398;
  assign n3933 = n609 & n3932;
  assign n3934 = n3821 & n3922;
  assign n3935 = n3933 & n3934;
  assign n3936 = ~n641 & ~n8700;
  assign n3937 = ~n884 & n3936;
  assign n3938 = n8760 & n3937;
  assign n3939 = n3927 & n3938;
  assign n3940 = n3935 & n3939;
  assign n3941 = n3926 & n3931;
  assign n3942 = n9052 & n9079;
  assign n3943 = n576 & n3821;
  assign n3944 = n609 & n3943;
  assign n3945 = n9052 & n3944;
  assign n3946 = n9078 & n3945;
  assign n3947 = n8760 & n3946;
  assign n3948 = ~n295 & n3947;
  assign n3949 = ~n8640 & n3948;
  assign n3950 = ~n8637 & n3949;
  assign n3951 = ~n8700 & n3950;
  assign n3952 = ~n228 & n3951;
  assign n3953 = ~n884 & n3952;
  assign n3954 = ~n641 & n3953;
  assign n3955 = ~n398 & n3954;
  assign n3956 = n9078 & n3942;
  assign n3957 = ~n3886 & ~n9080;
  assign n3958 = n9012 & ~n3227;
  assign n3959 = ~n9012 & ~n3228;
  assign n3960 = ~n9012 & ~n3227;
  assign n3961 = n3227 & ~n3228;
  assign n3962 = n9012 & n3227;
  assign n3963 = ~n9081 & ~n9082;
  assign n3964 = ~n3228 & ~n3958;
  assign n3965 = n447 & n8668;
  assign n3966 = n1603 & n9024;
  assign n3967 = n3965 & n3966;
  assign n3968 = ~n430 & ~n608;
  assign n3969 = ~n253 & ~n430;
  assign n3970 = ~n608 & n3969;
  assign n3971 = ~n253 & n3968;
  assign n3972 = ~n253 & n1355;
  assign n3973 = ~n430 & n3972;
  assign n3974 = ~n608 & n3973;
  assign n3975 = n1355 & n9084;
  assign n3976 = ~n610 & n1074;
  assign n3977 = n385 & ~n610;
  assign n3978 = n1074 & n3977;
  assign n3979 = n385 & n3976;
  assign n3980 = n9085 & n9086;
  assign n3981 = n1074 & n9024;
  assign n3982 = n447 & n3981;
  assign n3983 = n1603 & n3982;
  assign n3984 = n9085 & n3983;
  assign n3985 = n8668 & n3984;
  assign n3986 = n385 & n3985;
  assign n3987 = ~n610 & n3986;
  assign n3988 = n3967 & n3980;
  assign n3989 = n8658 & n8808;
  assign n3990 = n3808 & n3989;
  assign n3991 = ~n197 & ~n8700;
  assign n3992 = ~n8674 & ~n1345;
  assign n3993 = n3991 & n3992;
  assign n3994 = n8661 & n3993;
  assign n3995 = n8688 & n3994;
  assign n3996 = n8658 & n8661;
  assign n3997 = n8808 & n3996;
  assign n3998 = ~n8700 & ~n1345;
  assign n3999 = ~n8674 & n3998;
  assign n4000 = ~n197 & ~n967;
  assign n4001 = n1333 & n4000;
  assign n4002 = n3999 & n4001;
  assign n4003 = n8688 & n4002;
  assign n4004 = n3997 & n4003;
  assign n4005 = n3990 & n3995;
  assign n4006 = n9087 & n9088;
  assign n4007 = n8661 & n8808;
  assign n4008 = n8688 & n4007;
  assign n4009 = n1333 & n4008;
  assign n4010 = n9066 & n4009;
  assign n4011 = n8658 & n4010;
  assign n4012 = n9087 & n4011;
  assign n4013 = ~n197 & n4012;
  assign n4014 = ~n8700 & n4013;
  assign n4015 = ~n967 & n4014;
  assign n4016 = ~n8674 & n4015;
  assign n4017 = ~n1345 & n4016;
  assign n4018 = n9066 & n4006;
  assign n4019 = ~n9083 & n9089;
  assign n4020 = n3886 & n9080;
  assign n4021 = ~n3957 & ~n4020;
  assign n4022 = ~n3957 & ~n4019;
  assign n4023 = ~n4020 & n4022;
  assign n4024 = ~n4019 & n4021;
  assign n4025 = ~n3957 & ~n9090;
  assign n4026 = n3807 & n9074;
  assign n4027 = ~n3884 & ~n4026;
  assign n4028 = ~n3884 & ~n4025;
  assign n4029 = ~n4026 & n4028;
  assign n4030 = ~n4025 & n4027;
  assign n4031 = ~n3884 & ~n9091;
  assign n4032 = n3744 & n9069;
  assign n4033 = ~n3805 & ~n4032;
  assign n4034 = ~n4031 & n4033;
  assign n4035 = ~n3805 & ~n4034;
  assign n4036 = n3658 & n9064;
  assign n4037 = ~n3742 & ~n4036;
  assign n4038 = ~n4035 & n4037;
  assign n4039 = ~n3742 & ~n4038;
  assign n4040 = n3595 & n9055;
  assign n4041 = ~n3656 & ~n4040;
  assign n4042 = ~n3656 & ~n4039;
  assign n4043 = ~n4040 & n4042;
  assign n4044 = ~n4039 & n4041;
  assign n4045 = ~n3656 & ~n9092;
  assign n4046 = n3516 & n9048;
  assign n4047 = ~n9048 & ~n3593;
  assign n4048 = ~n3516 & ~n3593;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = ~n3593 & ~n4046;
  assign n4051 = ~n4045 & ~n9093;
  assign n4052 = ~n3593 & ~n4051;
  assign n4053 = n3440 & n9040;
  assign n4054 = ~n3514 & ~n4053;
  assign n4055 = ~n3514 & ~n4052;
  assign n4056 = ~n4053 & n4055;
  assign n4057 = ~n4052 & n4054;
  assign n4058 = ~n3514 & ~n9094;
  assign n4059 = n3339 & n9030;
  assign n4060 = ~n3438 & ~n4059;
  assign n4061 = ~n4058 & n4060;
  assign n4062 = ~n3438 & ~n4061;
  assign n4063 = n3300 & n9020;
  assign n4064 = ~n3337 & ~n4063;
  assign n4065 = ~n3337 & ~n4062;
  assign n4066 = ~n4063 & n4065;
  assign n4067 = ~n4062 & n4064;
  assign n4068 = ~n3337 & ~n9095;
  assign n4069 = ~n3295 & ~n3298;
  assign n4070 = ~n3285 & ~n3292;
  assign n4071 = ~n1006 & ~n3289;
  assign n4072 = n8650 & n1021;
  assign n4073 = n8724 & ~n1021;
  assign n4074 = n8650 & ~n4073;
  assign n4075 = n8724 & ~n4072;
  assign n4076 = n987 & ~n1021;
  assign n4077 = ~n9096 & ~n4076;
  assign n4078 = ~n1544 & n4077;
  assign n4079 = n1544 & ~n4077;
  assign n4080 = ~n4078 & ~n4079;
  assign n4081 = ~n4071 & ~n4078;
  assign n4082 = ~n4079 & n4081;
  assign n4083 = ~n4071 & n4080;
  assign n4084 = n4071 & ~n4080;
  assign n4085 = ~n4071 & ~n9097;
  assign n4086 = ~n4078 & ~n9097;
  assign n4087 = ~n4079 & n4086;
  assign n4088 = ~n4085 & ~n4087;
  assign n4089 = ~n9097 & ~n4084;
  assign n4090 = ~n4070 & ~n9098;
  assign n4091 = n4070 & n9098;
  assign n4092 = ~n4070 & n9098;
  assign n4093 = n4070 & ~n9098;
  assign n4094 = ~n4092 & ~n4093;
  assign n4095 = ~n4090 & ~n4091;
  assign n4096 = ~n4069 & ~n9099;
  assign n4097 = n4069 & n9099;
  assign n4098 = ~n4096 & ~n4097;
  assign n4099 = n187 & n272;
  assign n4100 = n394 & n1252;
  assign n4101 = n4099 & n4100;
  assign n4102 = ~n342 & ~n625;
  assign n4103 = ~n279 & ~n436;
  assign n4104 = n4102 & n4103;
  assign n4105 = n9025 & n4104;
  assign n4106 = n4101 & n4105;
  assign n4107 = n8665 & n4106;
  assign n4108 = n9037 & n4107;
  assign n4109 = ~n613 & ~n1163;
  assign n4110 = ~n798 & ~n967;
  assign n4111 = ~n474 & n4110;
  assign n4112 = ~n474 & ~n613;
  assign n4113 = ~n967 & n4112;
  assign n4114 = ~n1163 & n4113;
  assign n4115 = ~n798 & n4114;
  assign n4116 = ~n474 & ~n1163;
  assign n4117 = ~n613 & ~n967;
  assign n4118 = ~n798 & n4117;
  assign n4119 = n4116 & n4118;
  assign n4120 = n4109 & n4111;
  assign n4121 = ~n431 & ~n747;
  assign n4122 = ~n8674 & n4121;
  assign n4123 = ~n198 & ~n8648;
  assign n4124 = n449 & n4123;
  assign n4125 = n381 & n4124;
  assign n4126 = ~n8648 & ~n747;
  assign n4127 = ~n8674 & n4126;
  assign n4128 = ~n431 & ~n448;
  assign n4129 = ~n198 & ~n280;
  assign n4130 = n4128 & n4129;
  assign n4131 = n381 & n4130;
  assign n4132 = n4127 & n4131;
  assign n4133 = n4122 & n4125;
  assign n4134 = n381 & n9100;
  assign n4135 = ~n8648 & n4134;
  assign n4136 = ~n198 & n4135;
  assign n4137 = ~n280 & n4136;
  assign n4138 = ~n431 & n4137;
  assign n4139 = ~n8674 & n4138;
  assign n4140 = ~n747 & n4139;
  assign n4141 = ~n448 & n4140;
  assign n4142 = n9100 & n9101;
  assign n4143 = n9087 & n9102;
  assign n4144 = n187 & n1252;
  assign n4145 = n272 & n4144;
  assign n4146 = n8665 & n4145;
  assign n4147 = n9037 & n4146;
  assign n4148 = n9087 & n4147;
  assign n4149 = n9102 & n4148;
  assign n4150 = n9025 & n4149;
  assign n4151 = ~n342 & n4150;
  assign n4152 = ~n279 & n4151;
  assign n4153 = ~n392 & n4152;
  assign n4154 = ~n436 & n4153;
  assign n4155 = ~n625 & n4154;
  assign n4156 = ~n393 & n4155;
  assign n4157 = n4108 & n4143;
  assign n4158 = ~n4098 & ~n9103;
  assign n4159 = n4098 & n9103;
  assign n4160 = ~n4158 & ~n4159;
  assign n4161 = ~n4068 & n4160;
  assign n4162 = n4068 & ~n4160;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = ~n4158 & ~n4161;
  assign n4165 = ~n164 & ~n490;
  assign n4166 = ~n222 & ~n817;
  assign n4167 = n4165 & n4166;
  assign n4168 = n1344 & n3922;
  assign n4169 = n816 & n860;
  assign n4170 = n4168 & n4169;
  assign n4171 = n860 & n1344;
  assign n4172 = n816 & n3922;
  assign n4173 = n4167 & n4172;
  assign n4174 = n4171 & n4173;
  assign n4175 = n4167 & n4170;
  assign n4176 = ~n223 & ~n820;
  assign n4177 = ~n8629 & ~n223;
  assign n4178 = ~n820 & n4177;
  assign n4179 = ~n8629 & n4176;
  assign n4180 = ~n8629 & ~n295;
  assign n4181 = ~n314 & n4180;
  assign n4182 = ~n223 & n4181;
  assign n4183 = ~n820 & n4182;
  assign n4184 = n592 & n9105;
  assign n4185 = ~n270 & ~n1163;
  assign n4186 = ~n8663 & ~n1163;
  assign n4187 = ~n270 & n4186;
  assign n4188 = ~n8663 & n4185;
  assign n4189 = ~n270 & n9023;
  assign n4190 = ~n8663 & n4189;
  assign n4191 = ~n1163 & n4190;
  assign n4192 = n9023 & n9107;
  assign n4193 = n9106 & n9108;
  assign n4194 = n9104 & n4193;
  assign n4195 = n8685 & n8816;
  assign n4196 = n4194 & n4195;
  assign n4197 = n860 & n9059;
  assign n4198 = n4165 & n4197;
  assign n4199 = n4166 & n4198;
  assign n4200 = n1344 & n4199;
  assign n4201 = n9106 & n4200;
  assign n4202 = n9108 & n4201;
  assign n4203 = n816 & n4202;
  assign n4204 = n8685 & n4203;
  assign n4205 = n8816 & n4204;
  assign n4206 = ~n8640 & n4205;
  assign n4207 = ~n8637 & n4206;
  assign n4208 = n9059 & n4196;
  assign n4209 = ~n1021 & n8767;
  assign n4210 = n1021 & ~n8767;
  assign n4211 = n1021 & n8767;
  assign n4212 = ~n1021 & ~n8767;
  assign n4213 = ~n4211 & ~n4212;
  assign n4214 = ~n4209 & ~n4210;
  assign n4215 = ~n986 & n9110;
  assign n4216 = ~n986 & ~n9110;
  assign n4217 = n986 & n9110;
  assign n4218 = n986 & ~n9110;
  assign n4219 = ~n4215 & ~n4218;
  assign n4220 = ~n4216 & ~n4217;
  assign n4221 = ~n8650 & n9111;
  assign n4222 = ~n8650 & ~n4215;
  assign n4223 = ~n4090 & ~n4096;
  assign n4224 = n4086 & ~n4223;
  assign n4225 = ~n4086 & n4223;
  assign n4226 = ~n4224 & ~n4225;
  assign n4227 = n9112 & n4226;
  assign n4228 = ~n9112 & ~n4226;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = ~n9109 & ~n4229;
  assign n4231 = n9109 & n4229;
  assign n4232 = ~n4230 & ~n4231;
  assign n4233 = ~n4164 & ~n4230;
  assign n4234 = ~n4231 & n4233;
  assign n4235 = ~n4164 & n4232;
  assign n4236 = n4164 & ~n4232;
  assign n4237 = ~n4164 & ~n9113;
  assign n4238 = ~n4230 & ~n9113;
  assign n4239 = ~n4231 & n4238;
  assign n4240 = ~n4237 & ~n4239;
  assign n4241 = ~n9113 & ~n4236;
  assign n4242 = n4163 & ~n9114;
  assign n4243 = n4062 & ~n4064;
  assign n4244 = ~n4062 & ~n9095;
  assign n4245 = ~n4063 & n4068;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = ~n9095 & ~n4243;
  assign n4248 = n4163 & ~n9115;
  assign n4249 = n4058 & ~n4060;
  assign n4250 = ~n4061 & ~n4249;
  assign n4251 = ~n9115 & n4250;
  assign n4252 = n4052 & ~n4054;
  assign n4253 = ~n4052 & ~n9094;
  assign n4254 = ~n4053 & n4058;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = ~n9094 & ~n4252;
  assign n4257 = n4250 & ~n9116;
  assign n4258 = n4045 & n9093;
  assign n4259 = ~n4045 & ~n4051;
  assign n4260 = ~n9093 & ~n4051;
  assign n4261 = ~n4259 & ~n4260;
  assign n4262 = ~n4051 & ~n4258;
  assign n4263 = ~n9116 & ~n9117;
  assign n4264 = n4039 & ~n4041;
  assign n4265 = ~n4039 & ~n9092;
  assign n4266 = ~n4040 & n4045;
  assign n4267 = ~n4265 & ~n4266;
  assign n4268 = ~n9092 & ~n4264;
  assign n4269 = ~n9117 & ~n9118;
  assign n4270 = n4035 & ~n4037;
  assign n4271 = ~n4038 & ~n4270;
  assign n4272 = ~n9118 & n4271;
  assign n4273 = n4031 & ~n4033;
  assign n4274 = ~n4034 & ~n4273;
  assign n4275 = n4271 & n4274;
  assign n4276 = n4025 & ~n4027;
  assign n4277 = ~n4025 & ~n9091;
  assign n4278 = ~n4026 & n4031;
  assign n4279 = ~n4277 & ~n4278;
  assign n4280 = ~n9091 & ~n4276;
  assign n4281 = n4274 & ~n9119;
  assign n4282 = ~n4274 & n9119;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = n9083 & ~n9089;
  assign n4285 = ~n4019 & ~n4284;
  assign n4286 = n9119 & n4285;
  assign n4287 = n4019 & ~n4021;
  assign n4288 = ~n4019 & ~n9090;
  assign n4289 = ~n4020 & n4025;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = ~n9090 & ~n4287;
  assign n4292 = ~n9119 & ~n9120;
  assign n4293 = ~n4285 & ~n9120;
  assign n4294 = n9119 & n4293;
  assign n4295 = ~n4292 & ~n4294;
  assign n4296 = ~n4286 & ~n9120;
  assign n4297 = ~n4282 & ~n9121;
  assign n4298 = ~n4281 & n4297;
  assign n4299 = n4283 & ~n9121;
  assign n4300 = ~n4281 & ~n9122;
  assign n4301 = ~n4271 & ~n4274;
  assign n4302 = ~n4275 & ~n4301;
  assign n4303 = ~n4300 & ~n4301;
  assign n4304 = ~n4275 & n4303;
  assign n4305 = ~n4300 & n4302;
  assign n4306 = ~n4275 & ~n9123;
  assign n4307 = n9118 & ~n4271;
  assign n4308 = ~n4272 & ~n4307;
  assign n4309 = ~n4306 & n4308;
  assign n4310 = ~n4272 & ~n4309;
  assign n4311 = n9117 & n9118;
  assign n4312 = ~n4269 & ~n4311;
  assign n4313 = ~n4310 & n4312;
  assign n4314 = ~n4269 & ~n4313;
  assign n4315 = n9116 & n9117;
  assign n4316 = ~n4263 & ~n4315;
  assign n4317 = ~n4314 & n4316;
  assign n4318 = ~n4263 & ~n4317;
  assign n4319 = ~n4250 & n9116;
  assign n4320 = ~n4257 & ~n4319;
  assign n4321 = ~n4318 & n4320;
  assign n4322 = ~n4257 & ~n4321;
  assign n4323 = n9115 & ~n4250;
  assign n4324 = ~n4251 & ~n4323;
  assign n4325 = ~n4322 & n4324;
  assign n4326 = ~n4251 & ~n4325;
  assign n4327 = ~n4163 & n9115;
  assign n4328 = ~n4248 & ~n4327;
  assign n4329 = ~n4326 & n4328;
  assign n4330 = ~n4248 & ~n4329;
  assign n4331 = ~n4163 & n9114;
  assign n4332 = ~n4242 & ~n4331;
  assign n4333 = ~n4330 & n4332;
  assign n4334 = ~n4242 & ~n4333;
  assign n4335 = n905 & n1120;
  assign n4336 = n790 & n4335;
  assign n4337 = ~n204 & ~n560;
  assign n4338 = ~n387 & ~n1073;
  assign n4339 = ~n387 & ~n560;
  assign n4340 = ~n204 & ~n1073;
  assign n4341 = n4339 & n4340;
  assign n4342 = n4337 & n4338;
  assign n4343 = n1603 & n9124;
  assign n4344 = n4336 & n4343;
  assign n4345 = n8776 & n4344;
  assign n4346 = ~n8629 & ~n296;
  assign n4347 = ~n8645 & ~n493;
  assign n4348 = ~n207 & n4347;
  assign n4349 = ~n207 & ~n493;
  assign n4350 = ~n8629 & ~n8645;
  assign n4351 = ~n296 & n4350;
  assign n4352 = n4349 & n4351;
  assign n4353 = n4346 & n4348;
  assign n4354 = ~n207 & n8754;
  assign n4355 = ~n8629 & n4354;
  assign n4356 = ~n8645 & n4355;
  assign n4357 = ~n296 & n4356;
  assign n4358 = ~n493 & n4357;
  assign n4359 = n8754 & n9125;
  assign n4360 = n9052 & n9126;
  assign n4361 = n4345 & n4360;
  assign n4362 = n905 & n1603;
  assign n4363 = n9052 & n4362;
  assign n4364 = n8888 & n4363;
  assign n4365 = n9126 & n4364;
  assign n4366 = n8776 & n4365;
  assign n4367 = n1120 & n4366;
  assign n4368 = ~n204 & n4367;
  assign n4369 = n790 & n4368;
  assign n4370 = ~n387 & n4369;
  assign n4371 = ~n1073 & n4370;
  assign n4372 = ~n560 & n4371;
  assign n4373 = n8888 & n4361;
  assign n4374 = n4238 & n9127;
  assign n4375 = ~n4238 & ~n9127;
  assign n4376 = ~n4374 & ~n4375;
  assign n4377 = ~n9114 & ~n4376;
  assign n4378 = n9114 & n4376;
  assign n4379 = ~n4377 & ~n4378;
  assign n4380 = ~n4334 & n4379;
  assign n4381 = n4334 & ~n4379;
  assign n4382 = ~n4380 & ~n4381;
  assign n4383 = n90 & n4382;
  assign n4384 = ~n8621 & n8623;
  assign n4385 = ~n4376 & n4384;
  assign n4386 = ~n66 & n8622;
  assign n4387 = n66 & ~n8622;
  assign n4388 = n66 & n8622;
  assign n4389 = ~n66 & ~n8622;
  assign n4390 = ~n4388 & ~n4389;
  assign n4391 = ~n4386 & ~n4387;
  assign n4392 = n8621 & ~n8623;
  assign n4393 = ~n8623 & ~n9128;
  assign n4394 = n8621 & n4393;
  assign n4395 = ~n9128 & n4392;
  assign n4396 = n4163 & n9129;
  assign n4397 = ~n8623 & n9128;
  assign n4398 = ~n9114 & n4397;
  assign n4399 = ~n4396 & ~n4398;
  assign n4400 = ~n4385 & n4399;
  assign n4401 = ~n4383 & n4400;
  assign n4402 = ~n8620 & ~n4401;
  assign n4403 = n8620 & n4401;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = ~n854 & n8787;
  assign n4406 = n854 & ~n8787;
  assign n4407 = n854 & n8787;
  assign n4408 = ~n854 & ~n8787;
  assign n4409 = ~n4407 & ~n4408;
  assign n4410 = ~n4405 & ~n4406;
  assign n4411 = ~n997 & n8725;
  assign n4412 = n997 & ~n8725;
  assign n4413 = n997 & n8725;
  assign n4414 = ~n997 & ~n8725;
  assign n4415 = ~n4413 & ~n4414;
  assign n4416 = ~n4411 & ~n4412;
  assign n4417 = n9130 & n9131;
  assign n4418 = n4300 & ~n4302;
  assign n4419 = ~n4300 & ~n9123;
  assign n4420 = ~n4301 & n4306;
  assign n4421 = ~n4419 & ~n4420;
  assign n4422 = ~n9123 & ~n4418;
  assign n4423 = n4417 & ~n9132;
  assign n4424 = n9130 & ~n9131;
  assign n4425 = n4271 & n4424;
  assign n4426 = ~n997 & n8787;
  assign n4427 = n997 & ~n8787;
  assign n4428 = n997 & n8787;
  assign n4429 = ~n997 & ~n8787;
  assign n4430 = ~n4428 & ~n4429;
  assign n4431 = ~n4426 & ~n4427;
  assign n4432 = ~n9130 & n9133;
  assign n4433 = n4274 & n4432;
  assign n4434 = ~n9130 & n9131;
  assign n4435 = ~n9130 & ~n9133;
  assign n4436 = n9131 & n4435;
  assign n4437 = ~n9133 & n4434;
  assign n4438 = ~n9119 & n9134;
  assign n4439 = ~n4433 & ~n4438;
  assign n4440 = ~n4425 & ~n4433;
  assign n4441 = ~n4438 & n4440;
  assign n4442 = ~n4425 & n4439;
  assign n4443 = ~n4417 & n9135;
  assign n4444 = n9132 & n9135;
  assign n4445 = ~n4443 & ~n4444;
  assign n4446 = ~n4423 & n9135;
  assign n4447 = n8725 & ~n9136;
  assign n4448 = ~n8725 & n9136;
  assign n4449 = ~n4447 & ~n4448;
  assign n4450 = n8725 & ~n1325;
  assign n4451 = ~n8725 & n1325;
  assign n4452 = n8725 & n1325;
  assign n4453 = ~n8725 & ~n1325;
  assign n4454 = ~n4452 & ~n4453;
  assign n4455 = ~n4450 & ~n4451;
  assign n4456 = ~n1021 & ~n4285;
  assign n4457 = n9137 & n4456;
  assign n4458 = ~n4285 & n9120;
  assign n4459 = n4285 & ~n9120;
  assign n4460 = ~n4021 & n4285;
  assign n4461 = ~n4458 & ~n9138;
  assign n4462 = n9110 & n9137;
  assign n4463 = ~n4461 & n4462;
  assign n4464 = n8767 & ~n1325;
  assign n4465 = ~n8767 & n1325;
  assign n4466 = n8767 & n1325;
  assign n4467 = ~n8767 & ~n1325;
  assign n4468 = ~n4466 & ~n4467;
  assign n4469 = ~n4464 & ~n4465;
  assign n4470 = ~n9137 & n9139;
  assign n4471 = ~n4285 & n4470;
  assign n4472 = ~n9110 & n9137;
  assign n4473 = ~n9120 & n4472;
  assign n4474 = ~n4471 & ~n4473;
  assign n4475 = ~n4463 & n4474;
  assign n4476 = n4457 & ~n4475;
  assign n4477 = ~n4457 & n4475;
  assign n4478 = ~n4285 & n9137;
  assign n4479 = n4475 & ~n4478;
  assign n4480 = ~n1021 & ~n4478;
  assign n4481 = ~n1021 & ~n4475;
  assign n4482 = ~n1021 & ~n4481;
  assign n4483 = ~n4475 & ~n4481;
  assign n4484 = ~n4482 & ~n4483;
  assign n4485 = n4480 & ~n4484;
  assign n4486 = ~n1021 & n4479;
  assign n4487 = ~n4480 & n4484;
  assign n4488 = ~n9140 & ~n4487;
  assign n4489 = ~n4476 & ~n4477;
  assign n4490 = n4449 & n9141;
  assign n4491 = n4417 & ~n4461;
  assign n4492 = ~n4285 & n4432;
  assign n4493 = ~n9120 & n4424;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495 = ~n4491 & n4494;
  assign n4496 = ~n4285 & n9130;
  assign n4497 = ~n8725 & ~n4496;
  assign n4498 = ~n8725 & ~n4495;
  assign n4499 = n8725 & n4495;
  assign n4500 = ~n4498 & ~n4499;
  assign n4501 = n4497 & n4500;
  assign n4502 = n4495 & n4497;
  assign n4503 = ~n9119 & ~n9138;
  assign n4504 = n9119 & n9138;
  assign n4505 = n9119 & ~n9138;
  assign n4506 = ~n9119 & n9138;
  assign n4507 = ~n4505 & ~n4506;
  assign n4508 = ~n4503 & ~n4504;
  assign n4509 = n4417 & n9143;
  assign n4510 = ~n9119 & n4424;
  assign n4511 = ~n9120 & n4432;
  assign n4512 = ~n4285 & n9134;
  assign n4513 = ~n4511 & ~n4512;
  assign n4514 = ~n4510 & n4513;
  assign n4515 = ~n4417 & n4514;
  assign n4516 = ~n9143 & n4514;
  assign n4517 = ~n4515 & ~n4516;
  assign n4518 = ~n4509 & n4514;
  assign n4519 = n8725 & ~n9144;
  assign n4520 = ~n8725 & n9144;
  assign n4521 = ~n4519 & ~n4520;
  assign n4522 = n9142 & n4521;
  assign n4523 = n9142 & ~n9144;
  assign n4524 = n4478 & n9145;
  assign n4525 = ~n4283 & n9121;
  assign n4526 = ~n9121 & ~n9122;
  assign n4527 = ~n4282 & n4300;
  assign n4528 = ~n4526 & ~n4527;
  assign n4529 = ~n9122 & ~n4525;
  assign n4530 = n4417 & ~n9146;
  assign n4531 = n4274 & n4424;
  assign n4532 = ~n9120 & n9134;
  assign n4533 = ~n9119 & n4432;
  assign n4534 = ~n4532 & ~n4533;
  assign n4535 = ~n4531 & ~n4532;
  assign n4536 = ~n4533 & n4535;
  assign n4537 = ~n4531 & n4534;
  assign n4538 = ~n4530 & n9147;
  assign n4539 = ~n8725 & ~n4538;
  assign n4540 = n8725 & n4538;
  assign n4541 = ~n4539 & ~n4540;
  assign n4542 = ~n4478 & ~n9145;
  assign n4543 = n9145 & ~n4524;
  assign n4544 = ~n4478 & n9145;
  assign n4545 = n4478 & ~n4524;
  assign n4546 = n4478 & ~n9145;
  assign n4547 = ~n9148 & ~n9149;
  assign n4548 = ~n4524 & ~n4542;
  assign n4549 = n4541 & ~n9150;
  assign n4550 = ~n4524 & ~n4549;
  assign n4551 = ~n4449 & ~n9141;
  assign n4552 = ~n4490 & ~n4551;
  assign n4553 = ~n4550 & n4552;
  assign n4554 = ~n4490 & ~n4553;
  assign n4555 = n4306 & ~n4308;
  assign n4556 = ~n4309 & ~n4555;
  assign n4557 = n4417 & n4556;
  assign n4558 = ~n9118 & n4424;
  assign n4559 = n4271 & n4432;
  assign n4560 = n4274 & n9134;
  assign n4561 = ~n4559 & ~n4560;
  assign n4562 = ~n4558 & n4561;
  assign n4563 = ~n4557 & n4562;
  assign n4564 = ~n8725 & ~n4563;
  assign n4565 = n8725 & n4563;
  assign n4566 = ~n4564 & ~n4565;
  assign n4567 = ~n1021 & ~n4479;
  assign n4568 = n4462 & n9143;
  assign n4569 = ~n9119 & n4472;
  assign n4570 = ~n9120 & n4470;
  assign n4571 = ~n9137 & ~n9139;
  assign n4572 = n9110 & ~n9137;
  assign n4573 = ~n9139 & n4572;
  assign n4574 = n9110 & n4571;
  assign n4575 = ~n4285 & n9151;
  assign n4576 = ~n4570 & ~n4575;
  assign n4577 = ~n4569 & n4576;
  assign n4578 = ~n4462 & n4577;
  assign n4579 = ~n9143 & n4577;
  assign n4580 = ~n4578 & ~n4579;
  assign n4581 = ~n4568 & n4577;
  assign n4582 = n4567 & n9152;
  assign n4583 = ~n4567 & ~n9152;
  assign n4584 = n4479 & ~n9152;
  assign n4585 = ~n1021 & n4584;
  assign n4586 = n1021 & ~n9152;
  assign n4587 = ~n1021 & n9152;
  assign n4588 = ~n4586 & ~n4587;
  assign n4589 = n9140 & n4588;
  assign n4590 = n9140 & ~n9152;
  assign n4591 = ~n9140 & ~n4588;
  assign n4592 = ~n9153 & ~n4591;
  assign n4593 = ~n4582 & ~n4583;
  assign n4594 = n4566 & n9154;
  assign n4595 = ~n4566 & ~n9154;
  assign n4596 = ~n4594 & ~n4595;
  assign n4597 = n4554 & ~n4596;
  assign n4598 = ~n4554 & n4596;
  assign n4599 = ~n4597 & ~n4598;
  assign n4600 = n8620 & ~n1846;
  assign n4601 = ~n8620 & n1846;
  assign n4602 = n8620 & n1846;
  assign n4603 = ~n8620 & ~n1846;
  assign n4604 = ~n4602 & ~n4603;
  assign n4605 = ~n4600 & ~n4601;
  assign n4606 = n8651 & ~n854;
  assign n4607 = ~n8651 & n854;
  assign n4608 = n8651 & n854;
  assign n4609 = ~n8651 & ~n854;
  assign n4610 = ~n4608 & ~n4609;
  assign n4611 = ~n4606 & ~n4607;
  assign n4612 = n9155 & n9156;
  assign n4613 = n4318 & ~n4320;
  assign n4614 = ~n4321 & ~n4613;
  assign n4615 = n4612 & n4614;
  assign n4616 = n9155 & ~n9156;
  assign n4617 = n4250 & n4616;
  assign n4618 = n8651 & ~n1846;
  assign n4619 = ~n8651 & n1846;
  assign n4620 = n8651 & n1846;
  assign n4621 = ~n8651 & ~n1846;
  assign n4622 = ~n4620 & ~n4621;
  assign n4623 = ~n4618 & ~n4619;
  assign n4624 = ~n9155 & ~n9157;
  assign n4625 = ~n9155 & n9156;
  assign n4626 = ~n9157 & n4625;
  assign n4627 = n9156 & n4624;
  assign n4628 = ~n9117 & n9158;
  assign n4629 = ~n9155 & n9157;
  assign n4630 = ~n9116 & n4629;
  assign n4631 = ~n4628 & ~n4630;
  assign n4632 = ~n4617 & n4631;
  assign n4633 = ~n4614 & n4632;
  assign n4634 = ~n4612 & n4632;
  assign n4635 = ~n4633 & ~n4634;
  assign n4636 = ~n4615 & n4632;
  assign n4637 = n854 & ~n9159;
  assign n4638 = ~n854 & n9159;
  assign n4639 = ~n4637 & ~n4638;
  assign n4640 = n4599 & n4639;
  assign n4641 = ~n4599 & ~n4639;
  assign n4642 = n4599 & ~n4640;
  assign n4643 = n4639 & ~n4640;
  assign n4644 = ~n4642 & ~n4643;
  assign n4645 = ~n4640 & ~n4641;
  assign n4646 = n4314 & ~n4316;
  assign n4647 = ~n4317 & ~n4646;
  assign n4648 = n4612 & n4647;
  assign n4649 = ~n9116 & n4616;
  assign n4650 = ~n9117 & n4629;
  assign n4651 = ~n9118 & n9158;
  assign n4652 = ~n4650 & ~n4651;
  assign n4653 = ~n4649 & n4652;
  assign n4654 = ~n4648 & n4653;
  assign n4655 = ~n854 & ~n4654;
  assign n4656 = ~n4654 & ~n4655;
  assign n4657 = n854 & ~n4654;
  assign n4658 = ~n854 & ~n4655;
  assign n4659 = ~n854 & n4654;
  assign n4660 = ~n9161 & ~n9162;
  assign n4661 = n4550 & ~n4552;
  assign n4662 = ~n4553 & ~n4661;
  assign n4663 = n4660 & ~n4662;
  assign n4664 = ~n4660 & n4662;
  assign n4665 = n4310 & ~n4312;
  assign n4666 = ~n4313 & ~n4665;
  assign n4667 = n4612 & n4666;
  assign n4668 = ~n9117 & n4616;
  assign n4669 = ~n9118 & n4629;
  assign n4670 = n4271 & n9158;
  assign n4671 = ~n4669 & ~n4670;
  assign n4672 = ~n4668 & n4671;
  assign n4673 = ~n4666 & n4672;
  assign n4674 = ~n4612 & n4672;
  assign n4675 = ~n4673 & ~n4674;
  assign n4676 = ~n4667 & n4672;
  assign n4677 = n854 & ~n9163;
  assign n4678 = ~n854 & n9163;
  assign n4679 = ~n4677 & ~n4678;
  assign n4680 = ~n4541 & n9150;
  assign n4681 = ~n9150 & ~n4549;
  assign n4682 = ~n4541 & ~n9150;
  assign n4683 = n4541 & ~n4549;
  assign n4684 = n4541 & n9150;
  assign n4685 = ~n9164 & ~n9165;
  assign n4686 = ~n4549 & ~n4680;
  assign n4687 = n4679 & ~n9166;
  assign n4688 = ~n4679 & n9166;
  assign n4689 = ~n9166 & ~n4687;
  assign n4690 = ~n4679 & ~n9166;
  assign n4691 = n4679 & ~n4687;
  assign n4692 = n4679 & n9166;
  assign n4693 = ~n9167 & ~n9168;
  assign n4694 = ~n4687 & ~n4688;
  assign n4695 = n4556 & n4612;
  assign n4696 = ~n9118 & n4616;
  assign n4697 = n4271 & n4629;
  assign n4698 = n4274 & n9158;
  assign n4699 = ~n4697 & ~n4698;
  assign n4700 = ~n4696 & n4699;
  assign n4701 = ~n4695 & n4700;
  assign n4702 = ~n854 & ~n4701;
  assign n4703 = ~n4701 & ~n4702;
  assign n4704 = n854 & ~n4701;
  assign n4705 = ~n854 & ~n4702;
  assign n4706 = ~n854 & n4701;
  assign n4707 = ~n9170 & ~n9171;
  assign n4708 = ~n8725 & ~n9142;
  assign n4709 = n9144 & n4708;
  assign n4710 = ~n9144 & ~n4708;
  assign n4711 = ~n9142 & ~n4521;
  assign n4712 = ~n9145 & ~n4711;
  assign n4713 = ~n4709 & ~n4710;
  assign n4714 = n4707 & ~n9172;
  assign n4715 = ~n4707 & n9172;
  assign n4716 = ~n9132 & n4612;
  assign n4717 = n4271 & n4616;
  assign n4718 = n4274 & n4629;
  assign n4719 = ~n9119 & n9158;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = ~n4717 & ~n4718;
  assign n4722 = ~n4719 & n4721;
  assign n4723 = ~n4717 & n4720;
  assign n4724 = ~n4612 & n9173;
  assign n4725 = n9132 & n9173;
  assign n4726 = ~n4724 & ~n4725;
  assign n4727 = ~n4716 & n9173;
  assign n4728 = n854 & ~n9174;
  assign n4729 = ~n854 & n9174;
  assign n4730 = ~n4728 & ~n4729;
  assign n4731 = ~n8725 & n4496;
  assign n4732 = ~n4495 & n4731;
  assign n4733 = n4495 & ~n4731;
  assign n4734 = ~n4497 & ~n4500;
  assign n4735 = ~n9142 & ~n4734;
  assign n4736 = ~n4732 & ~n4733;
  assign n4737 = n4730 & n9175;
  assign n4738 = ~n4461 & n4612;
  assign n4739 = ~n4285 & n4629;
  assign n4740 = ~n9120 & n4616;
  assign n4741 = ~n4739 & ~n4740;
  assign n4742 = ~n4738 & n4741;
  assign n4743 = ~n4285 & n9155;
  assign n4744 = ~n854 & ~n4743;
  assign n4745 = ~n854 & ~n4742;
  assign n4746 = ~n854 & ~n4745;
  assign n4747 = ~n4742 & ~n4745;
  assign n4748 = ~n4746 & ~n4747;
  assign n4749 = n4744 & ~n4748;
  assign n4750 = n4742 & n4744;
  assign n4751 = n9143 & n4612;
  assign n4752 = ~n9119 & n4616;
  assign n4753 = ~n9120 & n4629;
  assign n4754 = ~n4285 & n9158;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = ~n4752 & n4755;
  assign n4757 = ~n9143 & n4756;
  assign n4758 = ~n4612 & n4756;
  assign n4759 = ~n4757 & ~n4758;
  assign n4760 = ~n4751 & n4756;
  assign n4761 = n854 & ~n9177;
  assign n4762 = ~n854 & n9177;
  assign n4763 = ~n4761 & ~n4762;
  assign n4764 = n9176 & n4763;
  assign n4765 = n9176 & ~n9177;
  assign n4766 = n4496 & n9178;
  assign n4767 = ~n9146 & n4612;
  assign n4768 = n4274 & n4616;
  assign n4769 = ~n9120 & n9158;
  assign n4770 = ~n9119 & n4629;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = ~n4768 & ~n4769;
  assign n4773 = ~n4770 & n4772;
  assign n4774 = ~n4768 & n4771;
  assign n4775 = ~n4767 & n9179;
  assign n4776 = ~n854 & ~n4775;
  assign n4777 = ~n854 & ~n4776;
  assign n4778 = ~n854 & n4775;
  assign n4779 = ~n4775 & ~n4776;
  assign n4780 = n854 & ~n4775;
  assign n4781 = ~n9180 & ~n9181;
  assign n4782 = ~n4496 & ~n9178;
  assign n4783 = n9178 & ~n4766;
  assign n4784 = ~n4496 & n9178;
  assign n4785 = n4496 & ~n4766;
  assign n4786 = n4496 & ~n9178;
  assign n4787 = ~n9182 & ~n9183;
  assign n4788 = ~n4766 & ~n4782;
  assign n4789 = ~n4781 & ~n9184;
  assign n4790 = ~n4766 & ~n4789;
  assign n4791 = ~n4730 & ~n9175;
  assign n4792 = ~n4737 & ~n4791;
  assign n4793 = ~n4790 & n4792;
  assign n4794 = ~n4737 & ~n4793;
  assign n4795 = ~n4715 & n4794;
  assign n4796 = ~n4707 & ~n4715;
  assign n4797 = n9172 & ~n4715;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = ~n4714 & ~n4715;
  assign n4800 = ~n4794 & ~n9185;
  assign n4801 = ~n4715 & ~n4800;
  assign n4802 = ~n4714 & ~n4795;
  assign n4803 = ~n9169 & ~n9186;
  assign n4804 = ~n4687 & ~n4803;
  assign n4805 = ~n4664 & n4804;
  assign n4806 = ~n4660 & ~n4664;
  assign n4807 = n4662 & ~n4664;
  assign n4808 = ~n4806 & ~n4807;
  assign n4809 = ~n4663 & ~n4664;
  assign n4810 = ~n4804 & ~n9187;
  assign n4811 = ~n4664 & ~n4810;
  assign n4812 = ~n4663 & ~n4805;
  assign n4813 = ~n9160 & ~n9188;
  assign n4814 = ~n4640 & ~n4813;
  assign n4815 = ~n4594 & ~n4598;
  assign n4816 = n4417 & n4666;
  assign n4817 = ~n9117 & n4424;
  assign n4818 = ~n9118 & n4432;
  assign n4819 = n4271 & n9134;
  assign n4820 = ~n4818 & ~n4819;
  assign n4821 = ~n4817 & n4820;
  assign n4822 = ~n4816 & n4821;
  assign n4823 = ~n8725 & ~n4822;
  assign n4824 = n8725 & n4822;
  assign n4825 = ~n4823 & ~n4824;
  assign n4826 = n4456 & n9153;
  assign n4827 = ~n4285 & n9153;
  assign n4828 = n4456 & n4584;
  assign n4829 = ~n4456 & ~n9153;
  assign n4830 = ~n9189 & ~n4829;
  assign n4831 = ~n1021 & ~n4830;
  assign n4832 = n4462 & ~n9146;
  assign n4833 = n4274 & n4472;
  assign n4834 = ~n9120 & n9151;
  assign n4835 = ~n9119 & n4470;
  assign n4836 = ~n4834 & ~n4835;
  assign n4837 = ~n4833 & ~n4834;
  assign n4838 = ~n4835 & n4837;
  assign n4839 = ~n4833 & n4836;
  assign n4840 = ~n4832 & n9190;
  assign n4841 = n4831 & ~n4840;
  assign n4842 = ~n4831 & n4840;
  assign n4843 = ~n1021 & ~n4840;
  assign n4844 = ~n4840 & ~n4843;
  assign n4845 = n1021 & ~n4840;
  assign n4846 = ~n1021 & ~n4843;
  assign n4847 = ~n1021 & n4840;
  assign n4848 = ~n9191 & ~n9192;
  assign n4849 = ~n9189 & ~n4848;
  assign n4850 = ~n4829 & n4849;
  assign n4851 = n4830 & ~n4848;
  assign n4852 = ~n4848 & ~n9193;
  assign n4853 = ~n9189 & ~n9193;
  assign n4854 = ~n4829 & n4840;
  assign n4855 = ~n4829 & n9194;
  assign n4856 = ~n4852 & ~n4855;
  assign n4857 = ~n4830 & n4848;
  assign n4858 = ~n9193 & ~n4857;
  assign n4859 = ~n4841 & ~n4842;
  assign n4860 = n4825 & ~n9195;
  assign n4861 = ~n4825 & n9195;
  assign n4862 = n4825 & ~n4860;
  assign n4863 = ~n9195 & ~n4860;
  assign n4864 = ~n4862 & ~n4863;
  assign n4865 = ~n4860 & ~n4861;
  assign n4866 = n4815 & n9196;
  assign n4867 = ~n4815 & ~n9196;
  assign n4868 = ~n4866 & ~n4867;
  assign n4869 = n4322 & ~n4324;
  assign n4870 = ~n4325 & ~n4869;
  assign n4871 = n4612 & n4870;
  assign n4872 = ~n9115 & n4616;
  assign n4873 = n4250 & n4629;
  assign n4874 = ~n9116 & n9158;
  assign n4875 = ~n4873 & ~n4874;
  assign n4876 = ~n4872 & n4875;
  assign n4877 = ~n4870 & n4876;
  assign n4878 = ~n4612 & n4876;
  assign n4879 = ~n4877 & ~n4878;
  assign n4880 = ~n4871 & n4876;
  assign n4881 = n854 & ~n9197;
  assign n4882 = ~n854 & n9197;
  assign n4883 = ~n4881 & ~n4882;
  assign n4884 = n4868 & n4883;
  assign n4885 = ~n4868 & ~n4883;
  assign n4886 = n4868 & ~n4884;
  assign n4887 = n4883 & ~n4884;
  assign n4888 = ~n4886 & ~n4887;
  assign n4889 = ~n4884 & ~n4885;
  assign n4890 = ~n4814 & ~n9198;
  assign n4891 = n4814 & n9198;
  assign n4892 = ~n4814 & ~n4890;
  assign n4893 = ~n9198 & ~n4890;
  assign n4894 = ~n4892 & ~n4893;
  assign n4895 = ~n4890 & ~n4891;
  assign n4896 = n4404 & ~n9199;
  assign n4897 = n4330 & ~n4332;
  assign n4898 = ~n4333 & ~n4897;
  assign n4899 = n90 & n4898;
  assign n4900 = ~n9114 & n4384;
  assign n4901 = n4163 & n4397;
  assign n4902 = ~n9115 & n9129;
  assign n4903 = ~n4901 & ~n4902;
  assign n4904 = ~n4900 & n4903;
  assign n4905 = ~n4899 & n4904;
  assign n4906 = ~n8620 & ~n4905;
  assign n4907 = n8620 & n4905;
  assign n4908 = ~n4906 & ~n4907;
  assign n4909 = n9160 & n9188;
  assign n4910 = ~n9188 & ~n4813;
  assign n4911 = ~n9160 & ~n4813;
  assign n4912 = ~n4910 & ~n4911;
  assign n4913 = ~n4813 & ~n4909;
  assign n4914 = n4908 & ~n9200;
  assign n4915 = n4326 & ~n4328;
  assign n4916 = ~n4329 & ~n4915;
  assign n4917 = n90 & n4916;
  assign n4918 = n4163 & n4384;
  assign n4919 = n4250 & n9129;
  assign n4920 = ~n9115 & n4397;
  assign n4921 = ~n4919 & ~n4920;
  assign n4922 = ~n4918 & n4921;
  assign n4923 = ~n90 & n4922;
  assign n4924 = ~n4916 & n4922;
  assign n4925 = ~n4923 & ~n4924;
  assign n4926 = ~n4917 & n4922;
  assign n4927 = n8620 & ~n9201;
  assign n4928 = ~n8620 & n9201;
  assign n4929 = ~n4927 & ~n4928;
  assign n4930 = n4804 & ~n9187;
  assign n4931 = ~n4804 & n9187;
  assign n4932 = ~n4930 & ~n4931;
  assign n4933 = n4929 & ~n4932;
  assign n4934 = n90 & n4870;
  assign n4935 = ~n9115 & n4384;
  assign n4936 = n4250 & n4397;
  assign n4937 = ~n9116 & n9129;
  assign n4938 = ~n4936 & ~n4937;
  assign n4939 = ~n4935 & n4938;
  assign n4940 = ~n90 & n4939;
  assign n4941 = ~n4870 & n4939;
  assign n4942 = ~n4940 & ~n4941;
  assign n4943 = ~n4934 & n4939;
  assign n4944 = n8620 & ~n9202;
  assign n4945 = ~n8620 & n9202;
  assign n4946 = ~n4944 & ~n4945;
  assign n4947 = n9169 & n9186;
  assign n4948 = ~n9186 & ~n4803;
  assign n4949 = n9169 & ~n9186;
  assign n4950 = ~n9169 & ~n4803;
  assign n4951 = ~n9169 & n9186;
  assign n4952 = ~n9203 & ~n9204;
  assign n4953 = ~n4803 & ~n4947;
  assign n4954 = n4946 & ~n9205;
  assign n4955 = n90 & n4614;
  assign n4956 = n4250 & n4384;
  assign n4957 = ~n9117 & n9129;
  assign n4958 = ~n9116 & n4397;
  assign n4959 = ~n4957 & ~n4958;
  assign n4960 = ~n4956 & n4959;
  assign n4961 = ~n90 & n4960;
  assign n4962 = ~n4614 & n4960;
  assign n4963 = ~n4961 & ~n4962;
  assign n4964 = ~n4955 & n4960;
  assign n4965 = n8620 & ~n9206;
  assign n4966 = ~n8620 & n9206;
  assign n4967 = ~n4965 & ~n4966;
  assign n4968 = n4794 & ~n9185;
  assign n4969 = ~n4794 & n9185;
  assign n4970 = ~n4968 & ~n4969;
  assign n4971 = n4967 & ~n4970;
  assign n4972 = n90 & n4647;
  assign n4973 = ~n9116 & n4384;
  assign n4974 = ~n9117 & n4397;
  assign n4975 = ~n9118 & n9129;
  assign n4976 = ~n4974 & ~n4975;
  assign n4977 = ~n4973 & n4976;
  assign n4978 = ~n4972 & n4977;
  assign n4979 = ~n8620 & ~n4978;
  assign n4980 = n8620 & n4978;
  assign n4981 = ~n4979 & ~n4980;
  assign n4982 = n4790 & ~n4792;
  assign n4983 = ~n4793 & ~n4982;
  assign n4984 = n4981 & n4983;
  assign n4985 = n90 & n4666;
  assign n4986 = ~n9117 & n4384;
  assign n4987 = ~n9118 & n4397;
  assign n4988 = n4271 & n9129;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 = ~n4986 & n4989;
  assign n4991 = ~n90 & n4990;
  assign n4992 = ~n4666 & n4990;
  assign n4993 = ~n4991 & ~n4992;
  assign n4994 = ~n4985 & n4990;
  assign n4995 = n8620 & ~n9207;
  assign n4996 = ~n8620 & n9207;
  assign n4997 = ~n4995 & ~n4996;
  assign n4998 = n4781 & n9184;
  assign n4999 = ~n9184 & ~n4789;
  assign n5000 = ~n4781 & ~n4789;
  assign n5001 = ~n4999 & ~n5000;
  assign n5002 = ~n4789 & ~n4998;
  assign n5003 = n4997 & ~n9208;
  assign n5004 = n90 & n4556;
  assign n5005 = ~n9118 & n4384;
  assign n5006 = n4271 & n4397;
  assign n5007 = n4274 & n9129;
  assign n5008 = ~n5006 & ~n5007;
  assign n5009 = ~n5005 & n5008;
  assign n5010 = ~n5004 & n5009;
  assign n5011 = ~n8620 & ~n5010;
  assign n5012 = n8620 & n5010;
  assign n5013 = ~n5011 & ~n5012;
  assign n5014 = ~n854 & ~n9176;
  assign n5015 = n9177 & n5014;
  assign n5016 = ~n9177 & ~n5014;
  assign n5017 = ~n9176 & ~n4763;
  assign n5018 = ~n9178 & ~n5017;
  assign n5019 = ~n5015 & ~n5016;
  assign n5020 = n5013 & n9209;
  assign n5021 = n90 & ~n9132;
  assign n5022 = n4271 & n4384;
  assign n5023 = n4274 & n4397;
  assign n5024 = ~n9119 & n9129;
  assign n5025 = ~n5023 & ~n5024;
  assign n5026 = ~n5022 & ~n5023;
  assign n5027 = ~n5024 & n5026;
  assign n5028 = ~n5022 & n5025;
  assign n5029 = ~n90 & n9210;
  assign n5030 = n9132 & n9210;
  assign n5031 = ~n5029 & ~n5030;
  assign n5032 = ~n5021 & n9210;
  assign n5033 = n8620 & ~n9211;
  assign n5034 = ~n8620 & n9211;
  assign n5035 = ~n5033 & ~n5034;
  assign n5036 = ~n854 & n4743;
  assign n5037 = ~n4742 & n5036;
  assign n5038 = n4742 & ~n5036;
  assign n5039 = ~n4744 & n4748;
  assign n5040 = ~n9176 & ~n5039;
  assign n5041 = ~n5037 & ~n5038;
  assign n5042 = n5035 & n9212;
  assign n5043 = n90 & ~n4461;
  assign n5044 = ~n4285 & n4397;
  assign n5045 = ~n9120 & n4384;
  assign n5046 = ~n5044 & ~n5045;
  assign n5047 = ~n5043 & n5046;
  assign n5048 = n8623 & ~n4285;
  assign n5049 = ~n8620 & ~n5048;
  assign n5050 = ~n8620 & ~n5047;
  assign n5051 = n8620 & n5047;
  assign n5052 = ~n5050 & ~n5051;
  assign n5053 = n5049 & n5052;
  assign n5054 = n5047 & n5049;
  assign n5055 = n90 & n9143;
  assign n5056 = ~n9119 & n4384;
  assign n5057 = ~n9120 & n4397;
  assign n5058 = ~n4285 & n9129;
  assign n5059 = ~n5057 & ~n5058;
  assign n5060 = ~n5056 & n5059;
  assign n5061 = ~n90 & n5060;
  assign n5062 = ~n9143 & n5060;
  assign n5063 = ~n5061 & ~n5062;
  assign n5064 = ~n5055 & n5060;
  assign n5065 = n8620 & ~n9214;
  assign n5066 = ~n8620 & n9214;
  assign n5067 = ~n5065 & ~n5066;
  assign n5068 = n9213 & n5067;
  assign n5069 = n9213 & ~n9214;
  assign n5070 = n4743 & n9215;
  assign n5071 = n90 & ~n9146;
  assign n5072 = n4274 & n4384;
  assign n5073 = ~n9120 & n9129;
  assign n5074 = ~n9119 & n4397;
  assign n5075 = ~n5073 & ~n5074;
  assign n5076 = ~n5072 & ~n5073;
  assign n5077 = ~n5074 & n5076;
  assign n5078 = ~n5072 & n5075;
  assign n5079 = ~n5071 & n9216;
  assign n5080 = ~n8620 & ~n5079;
  assign n5081 = n8620 & n5079;
  assign n5082 = ~n5080 & ~n5081;
  assign n5083 = ~n4743 & ~n9215;
  assign n5084 = n9215 & ~n5070;
  assign n5085 = ~n4743 & n9215;
  assign n5086 = n4743 & ~n5070;
  assign n5087 = n4743 & ~n9215;
  assign n5088 = ~n9217 & ~n9218;
  assign n5089 = ~n5070 & ~n5083;
  assign n5090 = n5082 & ~n9219;
  assign n5091 = ~n5070 & ~n5090;
  assign n5092 = ~n5035 & ~n9212;
  assign n5093 = ~n5042 & ~n5092;
  assign n5094 = ~n5091 & n5093;
  assign n5095 = ~n5042 & ~n5094;
  assign n5096 = ~n5013 & ~n9209;
  assign n5097 = ~n5020 & ~n5096;
  assign n5098 = ~n5095 & n5097;
  assign n5099 = ~n5020 & ~n5098;
  assign n5100 = ~n4997 & n9208;
  assign n5101 = ~n9208 & ~n5003;
  assign n5102 = n4997 & ~n5003;
  assign n5103 = ~n5101 & ~n5102;
  assign n5104 = ~n5003 & ~n5100;
  assign n5105 = ~n5099 & ~n9220;
  assign n5106 = ~n5003 & ~n5105;
  assign n5107 = ~n4981 & ~n4983;
  assign n5108 = ~n4984 & ~n5107;
  assign n5109 = ~n5106 & n5108;
  assign n5110 = ~n4984 & ~n5109;
  assign n5111 = ~n4967 & n4970;
  assign n5112 = ~n4970 & ~n4971;
  assign n5113 = n4967 & ~n4971;
  assign n5114 = ~n5112 & ~n5113;
  assign n5115 = ~n4971 & ~n5111;
  assign n5116 = ~n5110 & ~n9221;
  assign n5117 = ~n4971 & ~n5116;
  assign n5118 = ~n4946 & n9205;
  assign n5119 = ~n9205 & ~n4954;
  assign n5120 = ~n4946 & ~n9205;
  assign n5121 = n4946 & ~n4954;
  assign n5122 = n4946 & n9205;
  assign n5123 = ~n9222 & ~n9223;
  assign n5124 = ~n4954 & ~n5118;
  assign n5125 = ~n5117 & ~n9224;
  assign n5126 = ~n4954 & ~n5125;
  assign n5127 = ~n4929 & n4932;
  assign n5128 = ~n4933 & ~n5127;
  assign n5129 = ~n5126 & n5128;
  assign n5130 = ~n4933 & ~n5129;
  assign n5131 = ~n4908 & n9200;
  assign n5132 = n4908 & ~n4914;
  assign n5133 = ~n9200 & ~n4914;
  assign n5134 = ~n5132 & ~n5133;
  assign n5135 = ~n4914 & ~n5131;
  assign n5136 = ~n5130 & ~n9225;
  assign n5137 = ~n4914 & ~n5136;
  assign n5138 = ~n4404 & n9199;
  assign n5139 = n4404 & ~n4896;
  assign n5140 = ~n9199 & ~n4896;
  assign n5141 = ~n5139 & ~n5140;
  assign n5142 = ~n4896 & ~n5138;
  assign n5143 = ~n5137 & ~n9226;
  assign n5144 = ~n4896 & ~n5143;
  assign n5145 = ~n4377 & ~n4380;
  assign n5146 = ~n475 & n1252;
  assign n5147 = ~n253 & ~n861;
  assign n5148 = ~n8664 & n5147;
  assign n5149 = n9025 & n5148;
  assign n5150 = n5146 & n5149;
  assign n5151 = ~n444 & ~n8700;
  assign n5152 = ~n331 & ~n341;
  assign n5153 = ~n8674 & n5152;
  assign n5154 = ~n8700 & n5152;
  assign n5155 = ~n444 & n5154;
  assign n5156 = ~n8674 & n5155;
  assign n5157 = ~n341 & ~n444;
  assign n5158 = ~n331 & ~n8700;
  assign n5159 = ~n8674 & n5158;
  assign n5160 = n5157 & n5159;
  assign n5161 = n5151 & n5153;
  assign n5162 = ~n8648 & ~n1163;
  assign n5163 = ~n545 & ~n967;
  assign n5164 = n5162 & n5163;
  assign n5165 = ~n798 & ~n820;
  assign n5166 = ~n433 & ~n686;
  assign n5167 = n5165 & n5166;
  assign n5168 = n5164 & n5167;
  assign n5169 = n9227 & n5168;
  assign n5170 = ~n475 & ~n1163;
  assign n5171 = ~n1163 & n5146;
  assign n5172 = n1252 & n5170;
  assign n5173 = n9227 & n9228;
  assign n5174 = n9025 & n5173;
  assign n5175 = ~n253 & n5174;
  assign n5176 = ~n8648 & n5175;
  assign n5177 = ~n861 & n5176;
  assign n5178 = ~n545 & n5177;
  assign n5179 = ~n8664 & n5178;
  assign n5180 = ~n820 & n5179;
  assign n5181 = ~n686 & n5180;
  assign n5182 = ~n967 & n5181;
  assign n5183 = ~n433 & n5182;
  assign n5184 = ~n798 & n5183;
  assign n5185 = ~n8648 & ~n545;
  assign n5186 = ~n861 & ~n967;
  assign n5187 = n5185 & n5186;
  assign n5188 = n9025 & n5187;
  assign n5189 = n9228 & n5188;
  assign n5190 = ~n253 & ~n8664;
  assign n5191 = n5165 & n5190;
  assign n5192 = n5166 & n5191;
  assign n5193 = n9227 & n5192;
  assign n5194 = n5189 & n5193;
  assign n5195 = n5150 & n5169;
  assign n5196 = ~n8640 & ~n431;
  assign n5197 = ~n271 & ~n8640;
  assign n5198 = ~n431 & n5197;
  assign n5199 = ~n271 & n5196;
  assign n5200 = ~n210 & ~n256;
  assign n5201 = ~n658 & ~n904;
  assign n5202 = n5200 & n5201;
  assign n5203 = n9060 & n5202;
  assign n5204 = n9230 & n5203;
  assign n5205 = ~n164 & ~n177;
  assign n5206 = ~n8645 & ~n938;
  assign n5207 = n1119 & n5206;
  assign n5208 = n5205 & n5207;
  assign n5209 = n8656 & n5208;
  assign n5210 = ~n210 & ~n8645;
  assign n5211 = ~n658 & ~n938;
  assign n5212 = n5210 & n5211;
  assign n5213 = n9060 & n5212;
  assign n5214 = n9230 & n5213;
  assign n5215 = ~n256 & ~n904;
  assign n5216 = n1119 & n5215;
  assign n5217 = n5205 & n5216;
  assign n5218 = n8656 & n5217;
  assign n5219 = n5214 & n5218;
  assign n5220 = n5204 & n5209;
  assign n5221 = n8655 & n9231;
  assign n5222 = n8656 & n9060;
  assign n5223 = n1119 & n5222;
  assign n5224 = n8655 & n5223;
  assign n5225 = n9229 & n5224;
  assign n5226 = n9230 & n5225;
  assign n5227 = ~n164 & n5226;
  assign n5228 = ~n256 & n5227;
  assign n5229 = ~n210 & n5228;
  assign n5230 = ~n8645 & n5229;
  assign n5231 = ~n177 & n5230;
  assign n5232 = ~n658 & n5231;
  assign n5233 = ~n938 & n5232;
  assign n5234 = ~n904 & n5233;
  assign n5235 = n9229 & n5221;
  assign n5236 = n4374 & n9232;
  assign n5237 = ~n4374 & ~n9232;
  assign n5238 = ~n4374 & n9232;
  assign n5239 = n4374 & ~n9232;
  assign n5240 = ~n5238 & ~n5239;
  assign n5241 = ~n5236 & ~n5237;
  assign n5242 = ~n4376 & n9233;
  assign n5243 = n4376 & ~n9233;
  assign n5244 = n4376 & n9232;
  assign n5245 = ~n5242 & ~n9234;
  assign n5246 = ~n5145 & n5245;
  assign n5247 = n5145 & ~n5245;
  assign n5248 = ~n5246 & ~n5247;
  assign n5249 = n90 & n5248;
  assign n5250 = n4384 & n9233;
  assign n5251 = ~n4376 & n4397;
  assign n5252 = ~n9114 & n9129;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = ~n5250 & n5253;
  assign n5255 = ~n5249 & n5254;
  assign n5256 = ~n8620 & ~n5255;
  assign n5257 = n8620 & n5255;
  assign n5258 = ~n5256 & ~n5257;
  assign n5259 = ~n4884 & ~n4890;
  assign n5260 = n4612 & n4916;
  assign n5261 = n4163 & n4616;
  assign n5262 = n4250 & n9158;
  assign n5263 = ~n9115 & n4629;
  assign n5264 = ~n5262 & ~n5263;
  assign n5265 = ~n5261 & n5264;
  assign n5266 = ~n4916 & n5265;
  assign n5267 = ~n4612 & n5265;
  assign n5268 = ~n5266 & ~n5267;
  assign n5269 = ~n5260 & n5265;
  assign n5270 = n854 & ~n9235;
  assign n5271 = ~n854 & n9235;
  assign n5272 = ~n5270 & ~n5271;
  assign n5273 = ~n4860 & ~n4867;
  assign n5274 = n4417 & n4647;
  assign n5275 = ~n9116 & n4424;
  assign n5276 = ~n9117 & n4432;
  assign n5277 = ~n9118 & n9134;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = ~n5275 & n5278;
  assign n5280 = ~n5274 & n5279;
  assign n5281 = ~n8725 & ~n5280;
  assign n5282 = n8725 & n5280;
  assign n5283 = ~n5281 & ~n5282;
  assign n5284 = ~n1021 & n9120;
  assign n5285 = ~n9132 & n4462;
  assign n5286 = n4271 & n4472;
  assign n5287 = n4274 & n4470;
  assign n5288 = ~n9119 & n9151;
  assign n5289 = ~n5287 & ~n5288;
  assign n5290 = ~n5286 & ~n5287;
  assign n5291 = ~n5288 & n5290;
  assign n5292 = ~n5286 & n5289;
  assign n5293 = ~n5285 & n9236;
  assign n5294 = n5284 & ~n5293;
  assign n5295 = ~n5284 & n5293;
  assign n5296 = ~n1021 & ~n9120;
  assign n5297 = ~n1021 & ~n5293;
  assign n5298 = n5296 & ~n5297;
  assign n5299 = n5293 & n5296;
  assign n5300 = n5296 & ~n9237;
  assign n5301 = n1021 & n5293;
  assign n5302 = ~n5297 & ~n5301;
  assign n5303 = ~n9237 & n5302;
  assign n5304 = ~n5300 & ~n5303;
  assign n5305 = ~n5294 & ~n5295;
  assign n5306 = ~n9194 & ~n9238;
  assign n5307 = n9194 & n9238;
  assign n5308 = ~n9194 & ~n5306;
  assign n5309 = ~n9238 & ~n5306;
  assign n5310 = ~n5308 & ~n5309;
  assign n5311 = ~n5306 & ~n5307;
  assign n5312 = n5283 & ~n9239;
  assign n5313 = ~n5283 & n9239;
  assign n5314 = n5283 & ~n5312;
  assign n5315 = ~n9239 & ~n5312;
  assign n5316 = ~n5314 & ~n5315;
  assign n5317 = ~n5312 & ~n5313;
  assign n5318 = ~n5273 & ~n9240;
  assign n5319 = n5273 & n9240;
  assign n5320 = ~n5273 & n9240;
  assign n5321 = n5273 & ~n9240;
  assign n5322 = ~n5320 & ~n5321;
  assign n5323 = ~n5318 & ~n5319;
  assign n5324 = n5272 & ~n9241;
  assign n5325 = ~n5272 & n9241;
  assign n5326 = ~n5324 & ~n5325;
  assign n5327 = ~n5259 & n5326;
  assign n5328 = n5259 & ~n5326;
  assign n5329 = ~n5327 & ~n5328;
  assign n5330 = n5258 & n5329;
  assign n5331 = ~n5258 & ~n5329;
  assign n5332 = ~n5330 & ~n5331;
  assign n5333 = ~n5144 & n5332;
  assign n5334 = n5144 & ~n5332;
  assign n5335 = ~n5333 & ~n5334;
  assign n5336 = pi0  & ~pi22 ;
  assign n5337 = pi1  & ~n5336;
  assign n5338 = ~pi1  & n5336;
  assign n5339 = ~n5337 & ~n5338;
  assign n5340 = n83 & n5339;
  assign n5341 = ~n83 & ~n5339;
  assign n5342 = ~n83 & n5339;
  assign n5343 = n83 & ~n5339;
  assign n5344 = ~n5342 & ~n5343;
  assign n5345 = ~n5340 & ~n5341;
  assign n5346 = pi0  & ~n9242;
  assign n5347 = n602 & n3302;
  assign n5348 = n3811 & n5347;
  assign n5349 = ~n377 & ~n815;
  assign n5350 = ~n436 & n5349;
  assign n5351 = n1237 & n5350;
  assign n5352 = ~n377 & ~n480;
  assign n5353 = ~n815 & ~n817;
  assign n5354 = n5352 & n5353;
  assign n5355 = ~n430 & ~n436;
  assign n5356 = n1232 & n5355;
  assign n5357 = n602 & n3811;
  assign n5358 = n5356 & n5357;
  assign n5359 = n5354 & n5358;
  assign n5360 = n5348 & n5351;
  assign n5361 = n9021 & n9050;
  assign n5362 = n9243 & n5361;
  assign n5363 = n8713 & n5362;
  assign n5364 = ~n815 & n1232;
  assign n5365 = n8713 & n5364;
  assign n5366 = n8639 & n5365;
  assign n5367 = n9021 & n5366;
  assign n5368 = n9050 & n5367;
  assign n5369 = n3811 & n5368;
  assign n5370 = n602 & n5369;
  assign n5371 = ~n436 & n5370;
  assign n5372 = ~n430 & n5371;
  assign n5373 = ~n377 & n5372;
  assign n5374 = ~n817 & n5373;
  assign n5375 = ~n480 & n5374;
  assign n5376 = n8639 & n5363;
  assign n5377 = n5236 & n9244;
  assign n5378 = ~n229 & ~n8637;
  assign n5379 = n272 & n860;
  assign n5380 = n5378 & n5379;
  assign n5381 = n292 & n8824;
  assign n5382 = n5380 & n5381;
  assign n5383 = n8649 & n8708;
  assign n5384 = n5382 & n5383;
  assign n5385 = n8633 & n8713;
  assign n5386 = n8722 & n5385;
  assign n5387 = n8633 & n860;
  assign n5388 = n8824 & n5387;
  assign n5389 = n272 & n5388;
  assign n5390 = n8649 & n5389;
  assign n5391 = n291 & n5390;
  assign n5392 = n8713 & n5391;
  assign n5393 = n8722 & n5392;
  assign n5394 = n8708 & n5393;
  assign n5395 = n5378 & n5394;
  assign n5396 = ~n287 & n5395;
  assign n5397 = n5384 & n5386;
  assign n5398 = n5377 & n9245;
  assign n5399 = ~n5377 & ~n9245;
  assign n5400 = ~n5377 & n9245;
  assign n5401 = n5377 & ~n9245;
  assign n5402 = ~n5400 & ~n5401;
  assign n5403 = ~n5398 & ~n5399;
  assign n5404 = ~n5236 & ~n9244;
  assign n5405 = ~n5377 & ~n5404;
  assign n5406 = n9246 & ~n5405;
  assign n5407 = n9233 & ~n5405;
  assign n5408 = ~n5242 & ~n5246;
  assign n5409 = ~n9233 & n5405;
  assign n5410 = ~n9233 & n9244;
  assign n5411 = ~n5407 & ~n9247;
  assign n5412 = ~n5408 & n5411;
  assign n5413 = ~n5407 & ~n5412;
  assign n5414 = ~n9246 & n5405;
  assign n5415 = n9245 & n5405;
  assign n5416 = ~n5406 & ~n9248;
  assign n5417 = ~n5413 & n5416;
  assign n5418 = ~n5406 & ~n5417;
  assign n5419 = n8636 & n8713;
  assign n5420 = n8718 & n5419;
  assign n5421 = ~n359 & n8722;
  assign n5422 = ~n362 & n5421;
  assign n5423 = n363 & n8722;
  assign n5424 = ~n172 & ~n884;
  assign n5425 = n8644 & n5424;
  assign n5426 = n9249 & n5425;
  assign n5427 = n8718 & n9249;
  assign n5428 = n8713 & n5427;
  assign n5429 = n8636 & n5428;
  assign n5430 = n8644 & n5429;
  assign n5431 = ~n8629 & n5430;
  assign n5432 = ~n8631 & n5431;
  assign n5433 = ~n884 & n5432;
  assign n5434 = n5420 & n5426;
  assign n5435 = ~n5398 & ~n9250;
  assign n5436 = n5398 & n9250;
  assign n5437 = ~n5435 & ~n5436;
  assign n5438 = n9246 & ~n5437;
  assign n5439 = ~n9246 & n5437;
  assign n5440 = ~n9246 & n9250;
  assign n5441 = ~n5438 & ~n9251;
  assign n5442 = ~n5418 & n5441;
  assign n5443 = n5418 & ~n5441;
  assign n5444 = ~n5442 & ~n5443;
  assign n5445 = n5346 & n5444;
  assign n5446 = pi0  & n9242;
  assign n5447 = ~n5437 & n5446;
  assign n5448 = ~pi0  & ~n5339;
  assign n5449 = n9246 & n5448;
  assign n5450 = n50 & ~n9242;
  assign n5451 = pi2  & n50;
  assign n5452 = ~n5405 & n9252;
  assign n5453 = ~n5449 & ~n5452;
  assign n5454 = ~n5447 & n5453;
  assign n5455 = ~n5346 & n5454;
  assign n5456 = ~n5444 & n5454;
  assign n5457 = ~n5455 & ~n5456;
  assign n5458 = ~n5445 & n5454;
  assign n5459 = n83 & ~n9253;
  assign n5460 = ~n83 & n9253;
  assign n5461 = ~n5459 & ~n5460;
  assign n5462 = n5335 & n5461;
  assign n5463 = n5137 & n9226;
  assign n5464 = ~n5143 & ~n5463;
  assign n5465 = n5413 & ~n5416;
  assign n5466 = ~n5417 & ~n5465;
  assign n5467 = n5346 & n5466;
  assign n5468 = n9246 & n5446;
  assign n5469 = ~n5405 & n5448;
  assign n5470 = n9233 & n9252;
  assign n5471 = ~n5469 & ~n5470;
  assign n5472 = ~n5468 & n5471;
  assign n5473 = ~n5346 & n5472;
  assign n5474 = ~n5466 & n5472;
  assign n5475 = ~n5473 & ~n5474;
  assign n5476 = ~n5467 & n5472;
  assign n5477 = n83 & ~n9254;
  assign n5478 = ~n83 & n9254;
  assign n5479 = ~n5477 & ~n5478;
  assign n5480 = n5464 & n5479;
  assign n5481 = n5130 & n9225;
  assign n5482 = ~n5136 & ~n5481;
  assign n5483 = n5408 & ~n5411;
  assign n5484 = ~n5412 & ~n5483;
  assign n5485 = n5346 & n5484;
  assign n5486 = ~n5405 & n5446;
  assign n5487 = n9233 & n5448;
  assign n5488 = ~n4376 & n9252;
  assign n5489 = ~n5487 & ~n5488;
  assign n5490 = ~n5486 & n5489;
  assign n5491 = ~n5346 & n5490;
  assign n5492 = ~n5484 & n5490;
  assign n5493 = ~n5491 & ~n5492;
  assign n5494 = ~n5485 & n5490;
  assign n5495 = n83 & ~n9255;
  assign n5496 = ~n83 & n9255;
  assign n5497 = ~n5495 & ~n5496;
  assign n5498 = n5482 & n5497;
  assign n5499 = ~n5482 & ~n5497;
  assign n5500 = n5482 & ~n5498;
  assign n5501 = n5497 & ~n5498;
  assign n5502 = ~n5500 & ~n5501;
  assign n5503 = ~n5498 & ~n5499;
  assign n5504 = n5126 & ~n5128;
  assign n5505 = ~n5129 & ~n5504;
  assign n5506 = n5117 & n9224;
  assign n5507 = ~n5125 & ~n5506;
  assign n5508 = n5110 & n9221;
  assign n5509 = ~n5116 & ~n5508;
  assign n5510 = n5106 & ~n5108;
  assign n5511 = ~n5109 & ~n5510;
  assign n5512 = n5099 & n9220;
  assign n5513 = ~n5099 & ~n5105;
  assign n5514 = ~n9220 & ~n5105;
  assign n5515 = ~n5513 & ~n5514;
  assign n5516 = ~n5105 & ~n5512;
  assign n5517 = n5095 & ~n5097;
  assign n5518 = ~n5098 & ~n5517;
  assign n5519 = ~n9117 & n9252;
  assign n5520 = ~n83 & ~n5519;
  assign n5521 = n4614 & n5346;
  assign n5522 = n4250 & n5446;
  assign n5523 = ~n9116 & n5448;
  assign n5524 = ~n5522 & ~n5523;
  assign n5525 = ~n5521 & n5524;
  assign n5526 = ~n5520 & n5525;
  assign n5527 = ~n83 & ~n5525;
  assign n5528 = n83 & ~n5525;
  assign n5529 = n5520 & n5525;
  assign n5530 = ~n5528 & ~n5529;
  assign n5531 = ~n5526 & ~n5527;
  assign n5532 = n5518 & ~n9258;
  assign n5533 = n5091 & ~n5093;
  assign n5534 = ~n5094 & ~n5533;
  assign n5535 = ~n5082 & n9219;
  assign n5536 = ~n9219 & ~n5090;
  assign n5537 = n5082 & ~n5090;
  assign n5538 = ~n5536 & ~n5537;
  assign n5539 = ~n5090 & ~n5535;
  assign n5540 = ~n8620 & ~n9213;
  assign n5541 = n9214 & n5540;
  assign n5542 = ~n9214 & ~n5540;
  assign n5543 = ~n5541 & ~n5542;
  assign n5544 = ~n8620 & n5048;
  assign n5545 = ~n5047 & n5544;
  assign n5546 = n5047 & ~n5544;
  assign n5547 = ~n5049 & ~n5052;
  assign n5548 = ~n9213 & ~n5547;
  assign n5549 = ~n5545 & ~n5546;
  assign n5550 = n9119 & n9120;
  assign n5551 = n5446 & ~n5550;
  assign n5552 = n9119 & n4461;
  assign n5553 = n5346 & ~n5552;
  assign n5554 = ~n9120 & n5448;
  assign n5555 = ~n8619 & ~n4285;
  assign n5556 = ~n83 & ~n5555;
  assign n5557 = ~n5554 & n5556;
  assign n5558 = ~n5553 & n5557;
  assign n5559 = pi0  & ~n4285;
  assign n5560 = ~n83 & n5346;
  assign n5561 = n9143 & n5560;
  assign n5562 = ~n9119 & n5446;
  assign n5563 = ~n4285 & n9252;
  assign n5564 = ~n5554 & ~n5563;
  assign n5565 = ~n5562 & n5564;
  assign n5566 = ~n83 & ~n5565;
  assign n5567 = ~n4461 & n5560;
  assign n5568 = ~n9120 & n5446;
  assign n5569 = ~n4285 & n5448;
  assign n5570 = ~n83 & ~n5569;
  assign n5571 = ~n5568 & n5570;
  assign n5572 = ~n5567 & n5571;
  assign n5573 = ~n5566 & n5572;
  assign n5574 = ~n5561 & n5573;
  assign n5575 = ~n5559 & n5574;
  assign n5576 = ~n5552 & n5560;
  assign n5577 = ~n50 & ~n4285;
  assign n5578 = ~n83 & ~n5577;
  assign n5579 = ~n5568 & n5578;
  assign n5580 = ~n5576 & n5579;
  assign n5581 = ~n5566 & n5580;
  assign n5582 = ~n5551 & n5558;
  assign n5583 = ~n5048 & ~n9261;
  assign n5584 = ~n9146 & n5346;
  assign n5585 = ~n9119 & n5448;
  assign n5586 = n4274 & n5446;
  assign n5587 = ~n5585 & ~n5586;
  assign n5588 = ~n5584 & n5587;
  assign n5589 = n83 & ~n5588;
  assign n5590 = n50 & ~n9120;
  assign n5591 = ~n83 & ~n5590;
  assign n5592 = n5588 & n5591;
  assign n5593 = ~n9120 & n9252;
  assign n5594 = ~n5586 & ~n5593;
  assign n5595 = ~n5585 & n5594;
  assign n5596 = ~n5584 & n5595;
  assign n5597 = ~n83 & ~n5596;
  assign n5598 = n83 & n5596;
  assign n5599 = ~n5597 & ~n5598;
  assign n5600 = ~n5589 & ~n5592;
  assign n5601 = ~n5583 & n9262;
  assign n5602 = n9260 & n5601;
  assign n5603 = ~n9260 & ~n5601;
  assign n5604 = ~n9132 & n5346;
  assign n5605 = n4271 & n5446;
  assign n5606 = n4274 & n5448;
  assign n5607 = ~n9119 & n9252;
  assign n5608 = ~n5606 & ~n5607;
  assign n5609 = ~n5605 & ~n5606;
  assign n5610 = ~n5607 & n5609;
  assign n5611 = ~n5605 & n5608;
  assign n5612 = ~n5604 & n9263;
  assign n5613 = ~n83 & ~n5612;
  assign n5614 = n83 & n5612;
  assign n5615 = ~n5613 & ~n5614;
  assign n5616 = ~n83 & ~n9263;
  assign n5617 = ~n9132 & n5560;
  assign n5618 = ~n5603 & ~n5617;
  assign n5619 = ~n5614 & n5618;
  assign n5620 = ~n5616 & n5619;
  assign n5621 = ~n5603 & n5615;
  assign n5622 = ~n5602 & ~n9264;
  assign n5623 = ~n5543 & n5622;
  assign n5624 = n5543 & ~n5622;
  assign n5625 = n4556 & n5346;
  assign n5626 = ~n9118 & n5446;
  assign n5627 = n4271 & n5448;
  assign n5628 = n4274 & n9252;
  assign n5629 = ~n5627 & ~n5628;
  assign n5630 = ~n5626 & n5629;
  assign n5631 = ~n5625 & n5630;
  assign n5632 = ~n83 & ~n5631;
  assign n5633 = ~n5631 & ~n5632;
  assign n5634 = n83 & ~n5631;
  assign n5635 = ~n83 & ~n5632;
  assign n5636 = ~n83 & n5631;
  assign n5637 = ~n9265 & ~n9266;
  assign n5638 = ~n5624 & n5637;
  assign n5639 = ~n9213 & ~n5067;
  assign n5640 = n5622 & n5637;
  assign n5641 = ~n9215 & ~n5640;
  assign n5642 = ~n5639 & n5641;
  assign n5643 = ~n5622 & ~n5637;
  assign n5644 = ~n5642 & ~n5643;
  assign n5645 = ~n5623 & ~n5638;
  assign n5646 = ~n9259 & ~n9267;
  assign n5647 = n4666 & n5346;
  assign n5648 = ~n9117 & n5446;
  assign n5649 = ~n9118 & n5448;
  assign n5650 = n4271 & n9252;
  assign n5651 = ~n5649 & ~n5650;
  assign n5652 = ~n5648 & n5651;
  assign n5653 = ~n5647 & n5652;
  assign n5654 = n83 & ~n5653;
  assign n5655 = ~n83 & n5653;
  assign n5656 = ~n5654 & ~n5655;
  assign n5657 = ~n5646 & n5656;
  assign n5658 = n9259 & n9267;
  assign n5659 = ~n83 & ~n5652;
  assign n5660 = n83 & n5653;
  assign n5661 = n4666 & n5560;
  assign n5662 = ~n5658 & ~n5661;
  assign n5663 = ~n5660 & n5662;
  assign n5664 = ~n5659 & n5663;
  assign n5665 = ~n5646 & ~n5664;
  assign n5666 = ~n9267 & ~n5656;
  assign n5667 = n9267 & n5656;
  assign n5668 = ~n9259 & ~n5667;
  assign n5669 = ~n5666 & ~n5668;
  assign n5670 = ~n5657 & ~n5658;
  assign n5671 = n5534 & ~n9268;
  assign n5672 = n4647 & n5346;
  assign n5673 = ~n9116 & n5446;
  assign n5674 = ~n9117 & n5448;
  assign n5675 = ~n9118 & n9252;
  assign n5676 = ~n5674 & ~n5675;
  assign n5677 = ~n5673 & n5676;
  assign n5678 = ~n5672 & n5677;
  assign n5679 = ~n83 & ~n5678;
  assign n5680 = ~n5678 & ~n5679;
  assign n5681 = n83 & ~n5678;
  assign n5682 = ~n83 & ~n5679;
  assign n5683 = ~n83 & n5678;
  assign n5684 = ~n9269 & ~n9270;
  assign n5685 = ~n5671 & n5684;
  assign n5686 = ~n5534 & n9268;
  assign n5687 = ~n5518 & n9258;
  assign n5688 = ~n5686 & ~n5687;
  assign n5689 = ~n5685 & n5688;
  assign n5690 = n9268 & n5684;
  assign n5691 = ~n5094 & ~n5690;
  assign n5692 = ~n5533 & n5691;
  assign n5693 = ~n9268 & ~n5684;
  assign n5694 = ~n5692 & ~n5693;
  assign n5695 = ~n5685 & ~n5686;
  assign n5696 = n5518 & ~n9271;
  assign n5697 = ~n5518 & n9271;
  assign n5698 = ~n5519 & ~n5523;
  assign n5699 = ~n5522 & n5698;
  assign n5700 = ~n83 & ~n5699;
  assign n5701 = ~n5521 & n5699;
  assign n5702 = n83 & n5701;
  assign n5703 = n4614 & n5560;
  assign n5704 = ~n5697 & ~n5703;
  assign n5705 = ~n5702 & n5704;
  assign n5706 = ~n5700 & n5705;
  assign n5707 = ~n9258 & ~n5697;
  assign n5708 = ~n5696 & ~n9272;
  assign n5709 = ~n5532 & ~n5689;
  assign n5710 = ~n9257 & ~n9273;
  assign n5711 = n9257 & n9273;
  assign n5712 = n4870 & n5346;
  assign n5713 = ~n9115 & n5446;
  assign n5714 = n4250 & n5448;
  assign n5715 = ~n9116 & n9252;
  assign n5716 = ~n5714 & ~n5715;
  assign n5717 = ~n5713 & n5716;
  assign n5718 = ~n5712 & n5717;
  assign n5719 = ~n83 & ~n5718;
  assign n5720 = n83 & n5718;
  assign n5721 = ~n5719 & ~n5720;
  assign n5722 = ~n83 & ~n5717;
  assign n5723 = n4870 & n5560;
  assign n5724 = ~n5711 & ~n5723;
  assign n5725 = ~n5720 & n5724;
  assign n5726 = ~n5722 & n5725;
  assign n5727 = ~n5711 & n5721;
  assign n5728 = ~n5710 & ~n9274;
  assign n5729 = n5511 & ~n5728;
  assign n5730 = ~n5511 & n5728;
  assign n5731 = n4916 & n5346;
  assign n5732 = n4163 & n5446;
  assign n5733 = ~n9115 & n5448;
  assign n5734 = ~n5732 & ~n5733;
  assign n5735 = ~n5731 & n5734;
  assign n5736 = n4250 & n9252;
  assign n5737 = ~n83 & ~n5736;
  assign n5738 = n5735 & n5737;
  assign n5739 = n83 & ~n5735;
  assign n5740 = ~n5738 & ~n5739;
  assign n5741 = ~n5733 & ~n5736;
  assign n5742 = ~n5732 & n5741;
  assign n5743 = ~n83 & ~n5742;
  assign n5744 = ~n5731 & n5742;
  assign n5745 = n83 & n5744;
  assign n5746 = n4916 & n5560;
  assign n5747 = ~n5730 & ~n5746;
  assign n5748 = ~n5745 & n5747;
  assign n5749 = ~n5743 & n5748;
  assign n5750 = ~n5730 & ~n5740;
  assign n5751 = ~n5729 & ~n9275;
  assign n5752 = ~n5509 & n5751;
  assign n5753 = n5509 & ~n5751;
  assign n5754 = n4898 & n5346;
  assign n5755 = ~n9114 & n5446;
  assign n5756 = n4163 & n5448;
  assign n5757 = ~n9115 & n9252;
  assign n5758 = ~n5756 & ~n5757;
  assign n5759 = ~n5755 & n5758;
  assign n5760 = ~n5754 & n5759;
  assign n5761 = n83 & ~n5760;
  assign n5762 = ~n83 & n5760;
  assign n5763 = ~n5761 & ~n5762;
  assign n5764 = ~n5753 & n5763;
  assign n5765 = ~n5752 & ~n5764;
  assign n5766 = n5507 & n5765;
  assign n5767 = ~n5507 & ~n5765;
  assign n5768 = n4382 & n5346;
  assign n5769 = ~n4376 & n5446;
  assign n5770 = ~n9114 & n5448;
  assign n5771 = ~n5769 & ~n5770;
  assign n5772 = ~n5768 & n5771;
  assign n5773 = n4163 & n9252;
  assign n5774 = ~n83 & ~n5773;
  assign n5775 = n5772 & n5774;
  assign n5776 = n83 & ~n5772;
  assign n5777 = ~n5770 & ~n5773;
  assign n5778 = ~n5769 & n5777;
  assign n5779 = ~n5768 & n5778;
  assign n5780 = ~n83 & ~n5779;
  assign n5781 = n83 & n5779;
  assign n5782 = ~n5780 & ~n5781;
  assign n5783 = ~n5775 & ~n5776;
  assign n5784 = ~n5767 & n9276;
  assign n5785 = ~n5766 & ~n5784;
  assign n5786 = ~n5505 & n5785;
  assign n5787 = n5505 & ~n5785;
  assign n5788 = n5248 & n5346;
  assign n5789 = n9233 & n5446;
  assign n5790 = ~n4376 & n5448;
  assign n5791 = ~n9114 & n9252;
  assign n5792 = ~n5790 & ~n5791;
  assign n5793 = ~n5789 & n5792;
  assign n5794 = ~n5788 & n5793;
  assign n5795 = ~n83 & ~n5794;
  assign n5796 = ~n5794 & ~n5795;
  assign n5797 = n83 & ~n5794;
  assign n5798 = ~n83 & ~n5795;
  assign n5799 = ~n83 & n5794;
  assign n5800 = ~n9277 & ~n9278;
  assign n5801 = ~n5787 & n5800;
  assign n5802 = n5785 & n5800;
  assign n5803 = ~n5129 & ~n5802;
  assign n5804 = ~n5504 & n5803;
  assign n5805 = ~n5785 & ~n5800;
  assign n5806 = ~n5804 & ~n5805;
  assign n5807 = ~n5786 & ~n5801;
  assign n5808 = ~n9256 & ~n9279;
  assign n5809 = ~n5498 & ~n5808;
  assign n5810 = ~n5464 & ~n5479;
  assign n5811 = n5464 & ~n5480;
  assign n5812 = n5479 & ~n5480;
  assign n5813 = ~n5811 & ~n5812;
  assign n5814 = ~n5480 & ~n5810;
  assign n5815 = ~n5809 & ~n9280;
  assign n5816 = ~n5480 & ~n5815;
  assign n5817 = ~n5335 & ~n5461;
  assign n5818 = ~n5462 & ~n5817;
  assign n5819 = ~n5816 & n5818;
  assign n5820 = ~n5462 & ~n5819;
  assign n5821 = ~n5438 & ~n5442;
  assign n5822 = ~n228 & ~n271;
  assign n5823 = ~n8652 & ~n656;
  assign n5824 = n5822 & n5823;
  assign n5825 = ~n434 & ~n480;
  assign n5826 = n1033 & n3408;
  assign n5827 = n5825 & n5826;
  assign n5828 = n1033 & n5825;
  assign n5829 = ~n8652 & n5828;
  assign n5830 = ~n228 & n5829;
  assign n5831 = ~n288 & n5830;
  assign n5832 = ~n271 & n5831;
  assign n5833 = ~n398 & n5832;
  assign n5834 = ~n656 & n5833;
  assign n5835 = ~n8652 & ~n398;
  assign n5836 = ~n271 & ~n656;
  assign n5837 = n5835 & n5836;
  assign n5838 = ~n228 & ~n288;
  assign n5839 = n1033 & n5838;
  assign n5840 = n5825 & n5839;
  assign n5841 = n5837 & n5840;
  assign n5842 = n5824 & n5827;
  assign n5843 = ~n391 & ~n560;
  assign n5844 = n803 & n5843;
  assign n5845 = n3421 & n3811;
  assign n5846 = n5844 & n5845;
  assign n5847 = ~n243 & ~n542;
  assign n5848 = ~n384 & n5847;
  assign n5849 = n8732 & n5848;
  assign n5850 = ~n243 & ~n384;
  assign n5851 = ~n198 & ~n391;
  assign n5852 = n5850 & n5851;
  assign n5853 = n5845 & n5852;
  assign n5854 = ~n392 & ~n560;
  assign n5855 = ~n542 & n5854;
  assign n5856 = n8732 & n5855;
  assign n5857 = n5853 & n5856;
  assign n5858 = n5846 & n5849;
  assign n5859 = n9108 & n9282;
  assign n5860 = n9281 & n5859;
  assign n5861 = ~n542 & n8732;
  assign n5862 = n9108 & n5861;
  assign n5863 = n8823 & n5862;
  assign n5864 = n9281 & n5863;
  assign n5865 = n3811 & n5864;
  assign n5866 = ~n243 & n5865;
  assign n5867 = ~n340 & n5866;
  assign n5868 = ~n392 & n5867;
  assign n5869 = ~n198 & n5868;
  assign n5870 = ~n1073 & n5869;
  assign n5871 = ~n391 & n5870;
  assign n5872 = ~n384 & n5871;
  assign n5873 = ~n560 & n5872;
  assign n5874 = n8823 & n5860;
  assign n5875 = ~n5436 & ~n9283;
  assign n5876 = ~n5437 & ~n9283;
  assign n5877 = ~n5437 & n5875;
  assign n5878 = n5437 & n9283;
  assign n5879 = ~n9284 & ~n5878;
  assign n5880 = ~n5821 & n5879;
  assign n5881 = n5821 & ~n5879;
  assign n5882 = ~n5880 & ~n5881;
  assign n5883 = n5346 & n5882;
  assign n5884 = n5446 & n5875;
  assign n5885 = n5446 & ~n9283;
  assign n5886 = ~n5437 & n5448;
  assign n5887 = n9246 & n9252;
  assign n5888 = ~n5886 & ~n5887;
  assign n5889 = ~n9285 & n5888;
  assign n5890 = ~n5883 & n5889;
  assign n5891 = ~n83 & ~n5890;
  assign n5892 = ~n5890 & ~n5891;
  assign n5893 = n83 & ~n5890;
  assign n5894 = ~n83 & ~n5891;
  assign n5895 = ~n83 & n5890;
  assign n5896 = ~n9286 & ~n9287;
  assign n5897 = ~n5330 & ~n5333;
  assign n5898 = ~n5324 & ~n5327;
  assign n5899 = n4612 & n4898;
  assign n5900 = ~n9114 & n4616;
  assign n5901 = n4163 & n4629;
  assign n5902 = ~n9115 & n9158;
  assign n5903 = ~n5901 & ~n5902;
  assign n5904 = ~n5900 & n5903;
  assign n5905 = ~n5899 & n5904;
  assign n5906 = ~n854 & ~n5905;
  assign n5907 = ~n5905 & ~n5906;
  assign n5908 = n854 & ~n5905;
  assign n5909 = ~n854 & ~n5906;
  assign n5910 = ~n854 & n5905;
  assign n5911 = ~n9288 & ~n9289;
  assign n5912 = ~n5312 & ~n5318;
  assign n5913 = ~n1021 & n9119;
  assign n5914 = n4462 & n4556;
  assign n5915 = ~n9118 & n4472;
  assign n5916 = n4271 & n4470;
  assign n5917 = n4274 & n9151;
  assign n5918 = ~n5916 & ~n5917;
  assign n5919 = ~n5915 & n5918;
  assign n5920 = ~n5914 & n5919;
  assign n5921 = n5913 & ~n5920;
  assign n5922 = ~n5913 & n5920;
  assign n5923 = ~n5921 & ~n5922;
  assign n5924 = ~n9237 & ~n5306;
  assign n5925 = n5923 & ~n5924;
  assign n5926 = ~n5923 & n5924;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = n4417 & n4614;
  assign n5929 = n4250 & n4424;
  assign n5930 = ~n9117 & n9134;
  assign n5931 = ~n9116 & n4432;
  assign n5932 = ~n5930 & ~n5931;
  assign n5933 = ~n5929 & n5932;
  assign n5934 = ~n4417 & n5933;
  assign n5935 = ~n4614 & n5933;
  assign n5936 = ~n5934 & ~n5935;
  assign n5937 = ~n5928 & n5933;
  assign n5938 = n8725 & ~n9290;
  assign n5939 = ~n8725 & n9290;
  assign n5940 = ~n5938 & ~n5939;
  assign n5941 = n5927 & n5940;
  assign n5942 = ~n5927 & ~n5940;
  assign n5943 = n5927 & ~n5941;
  assign n5944 = n5940 & ~n5941;
  assign n5945 = ~n5943 & ~n5944;
  assign n5946 = ~n5941 & ~n5942;
  assign n5947 = ~n5912 & ~n9291;
  assign n5948 = n5912 & n9291;
  assign n5949 = ~n5912 & ~n5947;
  assign n5950 = ~n9291 & ~n5947;
  assign n5951 = ~n5949 & ~n5950;
  assign n5952 = ~n5947 & ~n5948;
  assign n5953 = ~n5911 & ~n9292;
  assign n5954 = n5911 & n9292;
  assign n5955 = ~n5911 & ~n5953;
  assign n5956 = ~n9292 & ~n5953;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = ~n5953 & ~n5954;
  assign n5959 = n5898 & n9293;
  assign n5960 = ~n5898 & ~n9293;
  assign n5961 = ~n5959 & ~n5960;
  assign n5962 = n90 & n5484;
  assign n5963 = n4384 & ~n5405;
  assign n5964 = n4397 & n9233;
  assign n5965 = ~n4376 & n9129;
  assign n5966 = ~n5964 & ~n5965;
  assign n5967 = ~n5963 & n5966;
  assign n5968 = ~n90 & n5967;
  assign n5969 = ~n5484 & n5967;
  assign n5970 = ~n5968 & ~n5969;
  assign n5971 = ~n5962 & n5967;
  assign n5972 = n8620 & ~n9294;
  assign n5973 = ~n8620 & n9294;
  assign n5974 = ~n5972 & ~n5973;
  assign n5975 = n5961 & n5974;
  assign n5976 = ~n5961 & ~n5974;
  assign n5977 = n5961 & ~n5975;
  assign n5978 = n5974 & ~n5975;
  assign n5979 = ~n5977 & ~n5978;
  assign n5980 = ~n5975 & ~n5976;
  assign n5981 = ~n5897 & ~n9295;
  assign n5982 = n5897 & n9295;
  assign n5983 = ~n5897 & ~n5981;
  assign n5984 = ~n9295 & ~n5981;
  assign n5985 = ~n5983 & ~n5984;
  assign n5986 = ~n5981 & ~n5982;
  assign n5987 = ~n5896 & ~n9296;
  assign n5988 = n5896 & n9296;
  assign n5989 = ~n5896 & ~n5987;
  assign n5990 = ~n9296 & ~n5987;
  assign n5991 = ~n5989 & ~n5990;
  assign n5992 = ~n5987 & ~n5988;
  assign n5993 = n5820 & n9297;
  assign n5994 = ~n5820 & ~n9297;
  assign n5995 = ~n5993 & ~n5994;
  assign n5996 = n8809 & n8887;
  assign n5997 = n9230 & n5996;
  assign n5998 = ~n251 & ~n490;
  assign n5999 = ~n362 & ~n490;
  assign n6000 = ~n251 & n5999;
  assign n6001 = ~n362 & n5998;
  assign n6002 = n1251 & n5825;
  assign n6003 = n9298 & n6002;
  assign n6004 = n8779 & n6003;
  assign n6005 = n5997 & n6004;
  assign n6006 = n8749 & n6005;
  assign n6007 = n8809 & n5825;
  assign n6008 = n1251 & n6007;
  assign n6009 = n8887 & n6008;
  assign n6010 = n9043 & n6009;
  assign n6011 = n8779 & n6010;
  assign n6012 = n8749 & n6011;
  assign n6013 = n9230 & n6012;
  assign n6014 = ~n251 & n6013;
  assign n6015 = ~n362 & n6014;
  assign n6016 = ~n490 & n6015;
  assign n6017 = n9043 & n6006;
  assign n6018 = ~n5995 & n9299;
  assign n6019 = n5995 & ~n9299;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = n5816 & ~n5818;
  assign n6022 = ~n5819 & ~n6021;
  assign n6023 = ~n8645 & ~n560;
  assign n6024 = ~n158 & ~n884;
  assign n6025 = ~n158 & ~n560;
  assign n6026 = ~n8645 & ~n884;
  assign n6027 = n6025 & n6026;
  assign n6028 = n6023 & n6024;
  assign n6029 = ~n279 & ~n8645;
  assign n6030 = ~n8648 & n6029;
  assign n6031 = ~n158 & n6030;
  assign n6032 = ~n884 & n6031;
  assign n6033 = ~n560 & n6032;
  assign n6034 = n3784 & n9300;
  assign n6035 = ~n8642 & ~n393;
  assign n6036 = ~n210 & ~n243;
  assign n6037 = ~n243 & ~n393;
  assign n6038 = ~n210 & ~n8642;
  assign n6039 = n6037 & n6038;
  assign n6040 = n6035 & n6036;
  assign n6041 = n1048 & n3385;
  assign n6042 = ~n8631 & ~n198;
  assign n6043 = n5825 & n6042;
  assign n6044 = n6041 & n6043;
  assign n6045 = n9302 & n6044;
  assign n6046 = n3385 & n5825;
  assign n6047 = n9301 & n6046;
  assign n6048 = ~n243 & n6047;
  assign n6049 = ~n8642 & n6048;
  assign n6050 = ~n210 & n6049;
  assign n6051 = ~n8631 & n6050;
  assign n6052 = ~n198 & n6051;
  assign n6053 = ~n445 & n6052;
  assign n6054 = ~n450 & n6053;
  assign n6055 = ~n393 & n6054;
  assign n6056 = n9301 & n6045;
  assign n6057 = ~n377 & ~n861;
  assign n6058 = ~n255 & ~n391;
  assign n6059 = n6057 & n6058;
  assign n6060 = ~n255 & n9303;
  assign n6061 = ~n861 & n6060;
  assign n6062 = ~n377 & n6061;
  assign n6063 = ~n391 & n6062;
  assign n6064 = n9303 & n6059;
  assign n6065 = ~n280 & ~n487;
  assign n6066 = n178 & n6065;
  assign n6067 = n8739 & n6066;
  assign n6068 = n178 & n9227;
  assign n6069 = n8739 & n6068;
  assign n6070 = ~n280 & n6069;
  assign n6071 = ~n487 & n6070;
  assign n6072 = n9227 & n6067;
  assign n6073 = ~n821 & n9230;
  assign n6074 = ~n240 & ~n721;
  assign n6075 = ~n166 & ~n721;
  assign n6076 = ~n240 & n6075;
  assign n6077 = ~n166 & n6074;
  assign n6078 = n4166 & n5166;
  assign n6079 = n9306 & n6078;
  assign n6080 = n3927 & n6079;
  assign n6081 = n6073 & n6080;
  assign n6082 = n8744 & n6081;
  assign n6083 = n9305 & n6082;
  assign n6084 = n576 & n4166;
  assign n6085 = n9304 & n6084;
  assign n6086 = n9230 & n6085;
  assign n6087 = n9305 & n6086;
  assign n6088 = n8744 & n6087;
  assign n6089 = ~n240 & n6088;
  assign n6090 = ~n166 & n6089;
  assign n6091 = ~n228 & n6090;
  assign n6092 = ~n821 & n6091;
  assign n6093 = ~n686 & n6092;
  assign n6094 = ~n721 & n6093;
  assign n6095 = ~n433 & n6094;
  assign n6096 = n9304 & n6083;
  assign n6097 = ~n6022 & n9307;
  assign n6098 = n6022 & ~n9307;
  assign n6099 = n5809 & ~n5812;
  assign n6100 = ~n5811 & n6099;
  assign n6101 = n5809 & n9280;
  assign n6102 = ~n5815 & ~n9308;
  assign n6103 = n9256 & n9279;
  assign n6104 = ~n244 & ~n904;
  assign n6105 = n272 & n6104;
  assign n6106 = ~n415 & ~n904;
  assign n6107 = ~n244 & ~n608;
  assign n6108 = n6106 & n6107;
  assign n6109 = n272 & n6108;
  assign n6110 = n2248 & n6105;
  assign n6111 = n9039 & n9309;
  assign n6112 = n272 & n9039;
  assign n6113 = n9045 & n6112;
  assign n6114 = ~n244 & n6113;
  assign n6115 = ~n415 & n6114;
  assign n6116 = ~n608 & n6115;
  assign n6117 = ~n904 & n6116;
  assign n6118 = n9045 & n6111;
  assign n6119 = ~n220 & ~n330;
  assign n6120 = n9106 & n6119;
  assign n6121 = n8758 & n9106;
  assign n6122 = ~n220 & n6121;
  assign n6123 = ~n330 & n6122;
  assign n6124 = n8758 & n6119;
  assign n6125 = n9106 & n6124;
  assign n6126 = n8758 & n6120;
  assign n6127 = n864 & n3847;
  assign n6128 = n3821 & n6042;
  assign n6129 = n6127 & n6128;
  assign n6130 = ~n296 & ~n469;
  assign n6131 = ~n253 & n6130;
  assign n6132 = ~n164 & ~n340;
  assign n6133 = n1344 & n6132;
  assign n6134 = ~n296 & n6132;
  assign n6135 = ~n253 & ~n469;
  assign n6136 = n1344 & n6135;
  assign n6137 = n6134 & n6136;
  assign n6138 = n6131 & n6133;
  assign n6139 = n6129 & n9312;
  assign n6140 = n9062 & n6139;
  assign n6141 = n9311 & n6140;
  assign n6142 = n864 & n3821;
  assign n6143 = n3847 & n6142;
  assign n6144 = n1344 & n6143;
  assign n6145 = n9311 & n6144;
  assign n6146 = n9310 & n6145;
  assign n6147 = n9062 & n6146;
  assign n6148 = ~n253 & n6147;
  assign n6149 = ~n164 & n6148;
  assign n6150 = ~n340 & n6149;
  assign n6151 = ~n8631 & n6150;
  assign n6152 = ~n296 & n6151;
  assign n6153 = ~n198 & n6152;
  assign n6154 = ~n469 & n6153;
  assign n6155 = n9310 & n6141;
  assign n6156 = ~n5808 & ~n9313;
  assign n6157 = ~n5808 & ~n6103;
  assign n6158 = ~n9313 & n6157;
  assign n6159 = ~n6103 & n6156;
  assign n6160 = ~n6102 & ~n9314;
  assign n6161 = n6102 & n9314;
  assign n6162 = ~n251 & ~n393;
  assign n6163 = n945 & n6162;
  assign n6164 = n3605 & n6163;
  assign n6165 = ~n398 & ~n823;
  assign n6166 = ~n513 & n6165;
  assign n6167 = n9056 & n6166;
  assign n6168 = ~n398 & ~n513;
  assign n6169 = n3605 & n6168;
  assign n6170 = n945 & n6169;
  assign n6171 = ~n393 & ~n823;
  assign n6172 = ~n251 & n6171;
  assign n6173 = n9056 & n6172;
  assign n6174 = n6170 & n6173;
  assign n6175 = n6164 & n6167;
  assign n6176 = n945 & n9056;
  assign n6177 = n8819 & n6176;
  assign n6178 = ~n445 & n6177;
  assign n6179 = ~n251 & n6178;
  assign n6180 = ~n418 & n6179;
  assign n6181 = ~n823 & n6180;
  assign n6182 = ~n398 & n6181;
  assign n6183 = ~n513 & n6182;
  assign n6184 = ~n393 & n6183;
  assign n6185 = n8819 & n9315;
  assign n6186 = ~n197 & ~n382;
  assign n6187 = n8760 & n6186;
  assign n6188 = n8760 & n9316;
  assign n6189 = ~n197 & n6188;
  assign n6190 = ~n382 & n6189;
  assign n6191 = n9316 & n6187;
  assign n6192 = ~n417 & ~n448;
  assign n6193 = ~n686 & ~n8686;
  assign n6194 = ~n610 & ~n8686;
  assign n6195 = ~n686 & n6194;
  assign n6196 = ~n610 & n6193;
  assign n6197 = ~n417 & ~n686;
  assign n6198 = ~n448 & n6197;
  assign n6199 = ~n8686 & n6198;
  assign n6200 = ~n610 & n6199;
  assign n6201 = n6192 & n9318;
  assign n6202 = ~n288 & ~n492;
  assign n6203 = ~n8643 & ~n386;
  assign n6204 = ~n8643 & ~n492;
  assign n6205 = ~n288 & ~n386;
  assign n6206 = n6204 & n6205;
  assign n6207 = n6202 & n6203;
  assign n6208 = n1192 & n1251;
  assign n6209 = n5205 & n6208;
  assign n6210 = n9320 & n6209;
  assign n6211 = n1251 & n9319;
  assign n6212 = ~n8643 & n6211;
  assign n6213 = ~n164 & n6212;
  assign n6214 = ~n177 & n6213;
  assign n6215 = ~n288 & n6214;
  assign n6216 = ~n8647 & n6215;
  assign n6217 = ~n492 & n6216;
  assign n6218 = ~n386 & n6217;
  assign n6219 = ~n433 & n6218;
  assign n6220 = n9319 & n6210;
  assign n6221 = ~n486 & ~n876;
  assign n6222 = ~n474 & n6221;
  assign n6223 = n567 & n1663;
  assign n6224 = n659 & n5165;
  assign n6225 = n6223 & n6224;
  assign n6226 = ~n220 & ~n474;
  assign n6227 = ~n876 & n6226;
  assign n6228 = ~n430 & ~n486;
  assign n6229 = n567 & n6228;
  assign n6230 = n6224 & n6229;
  assign n6231 = n6227 & n6230;
  assign n6232 = n6222 & n6225;
  assign n6233 = n9075 & n9322;
  assign n6234 = n9321 & n6233;
  assign n6235 = n9075 & n9317;
  assign n6236 = n9321 & n6235;
  assign n6237 = n567 & n6236;
  assign n6238 = ~n220 & n6237;
  assign n6239 = ~n474 & n6238;
  assign n6240 = ~n270 & n6239;
  assign n6241 = ~n658 & n6240;
  assign n6242 = ~n876 & n6241;
  assign n6243 = ~n430 & n6242;
  assign n6244 = ~n820 & n6243;
  assign n6245 = ~n486 & n6244;
  assign n6246 = ~n798 & n6245;
  assign n6247 = n9317 & n6234;
  assign n6248 = ~n6161 & n9323;
  assign n6249 = ~n6160 & ~n9323;
  assign n6250 = ~n6161 & ~n6249;
  assign n6251 = ~n6102 & n9323;
  assign n6252 = n6102 & ~n9323;
  assign n6253 = ~n9314 & ~n6252;
  assign n6254 = ~n6251 & ~n6253;
  assign n6255 = ~n6160 & ~n6248;
  assign n6256 = ~n6098 & n9324;
  assign n6257 = ~n9307 & ~n6098;
  assign n6258 = n6022 & ~n6098;
  assign n6259 = ~n6257 & ~n6258;
  assign n6260 = ~n6097 & ~n6098;
  assign n6261 = ~n9324 & ~n9325;
  assign n6262 = ~n6098 & ~n6261;
  assign n6263 = ~n6097 & ~n6256;
  assign n6264 = n6020 & ~n9326;
  assign n6265 = ~n6020 & n9326;
  assign n6266 = ~n6264 & ~n6265;
  assign n6267 = ~n9325 & ~n6261;
  assign n6268 = n9324 & ~n9325;
  assign n6269 = ~n9324 & ~n6261;
  assign n6270 = ~n9324 & n9325;
  assign n6271 = ~n9327 & ~n9328;
  assign n6272 = n6266 & ~n6271;
  assign n6273 = ~n6266 & n6271;
  assign n6274 = n6266 & ~n6272;
  assign n6275 = n6266 & n6271;
  assign n6276 = ~n6271 & ~n6272;
  assign n6277 = ~n6266 & ~n6271;
  assign n6278 = ~n9329 & ~n9330;
  assign n6279 = ~n6272 & ~n6273;
  assign n6280 = ~pi22  & ~pi23 ;
  assign n6281 = pi22  & pi23 ;
  assign n6282 = pi22  & ~pi23 ;
  assign n6283 = ~pi22  & pi23 ;
  assign n6284 = ~n6282 & ~n6283;
  assign n6285 = ~n6280 & ~n6281;
  assign n6286 = ~n9331 & ~n9332;
  assign n6287 = ~n6019 & ~n6264;
  assign n6288 = ~n5987 & ~n5994;
  assign n6289 = ~n9284 & ~n5880;
  assign n6290 = ~n487 & ~n821;
  assign n6291 = n1093 & n6290;
  assign n6292 = n385 & n3385;
  assign n6293 = n3847 & n6292;
  assign n6294 = n385 & n6290;
  assign n6295 = n1093 & n3385;
  assign n6296 = n3847 & n6295;
  assign n6297 = n6294 & n6296;
  assign n6298 = n6291 & n6293;
  assign n6299 = n3385 & n3847;
  assign n6300 = n8710 & n6299;
  assign n6301 = n385 & n6300;
  assign n6302 = ~n636 & n6301;
  assign n6303 = ~n821 & n6302;
  assign n6304 = ~n487 & n6303;
  assign n6305 = ~n8663 & n6304;
  assign n6306 = n8710 & n9333;
  assign n6307 = n602 & n687;
  assign n6308 = ~n625 & ~n1163;
  assign n6309 = ~n418 & ~n486;
  assign n6310 = n6308 & n6309;
  assign n6311 = n1074 & n6310;
  assign n6312 = n687 & n1074;
  assign n6313 = n602 & n6312;
  assign n6314 = n6310 & n6313;
  assign n6315 = n6307 & n6311;
  assign n6316 = n8890 & n9335;
  assign n6317 = n8759 & n9335;
  assign n6318 = n8890 & n6317;
  assign n6319 = n8759 & n6316;
  assign n6320 = n9334 & n9336;
  assign n6321 = n8759 & n6312;
  assign n6322 = n8890 & n6321;
  assign n6323 = n9334 & n6322;
  assign n6324 = n9071 & n6323;
  assign n6325 = n602 & n6324;
  assign n6326 = ~n418 & n6325;
  assign n6327 = ~n486 & n6326;
  assign n6328 = ~n625 & n6327;
  assign n6329 = ~n1163 & n6328;
  assign n6330 = n9071 & n6320;
  assign n6331 = ~n5875 & n9337;
  assign n6332 = n9283 & n9337;
  assign n6333 = n5875 & ~n9337;
  assign n6334 = ~n9283 & ~n9337;
  assign n6335 = n9283 & ~n9337;
  assign n6336 = ~n9283 & n9337;
  assign n6337 = ~n6335 & ~n6336;
  assign n6338 = ~n9338 & ~n9339;
  assign n6339 = ~n6289 & ~n9340;
  assign n6340 = n6289 & n9340;
  assign n6341 = ~n6339 & ~n6340;
  assign n6342 = n5346 & n6341;
  assign n6343 = n5446 & ~n9337;
  assign n6344 = n5448 & n5875;
  assign n6345 = n5448 & ~n9283;
  assign n6346 = ~n5437 & n9252;
  assign n6347 = ~n9341 & ~n6346;
  assign n6348 = ~n6343 & n6347;
  assign n6349 = ~n6342 & n6348;
  assign n6350 = ~n83 & ~n6349;
  assign n6351 = ~n6349 & ~n6350;
  assign n6352 = n83 & ~n6349;
  assign n6353 = ~n83 & ~n6350;
  assign n6354 = ~n83 & n6349;
  assign n6355 = ~n9342 & ~n9343;
  assign n6356 = ~n5975 & ~n5981;
  assign n6357 = ~n5953 & ~n5960;
  assign n6358 = n4382 & n4612;
  assign n6359 = ~n4376 & n4616;
  assign n6360 = n4163 & n9158;
  assign n6361 = ~n9114 & n4629;
  assign n6362 = ~n6360 & ~n6361;
  assign n6363 = ~n6359 & n6362;
  assign n6364 = ~n6358 & n6363;
  assign n6365 = ~n854 & ~n6364;
  assign n6366 = ~n6364 & ~n6365;
  assign n6367 = n854 & ~n6364;
  assign n6368 = ~n854 & ~n6365;
  assign n6369 = ~n854 & n6364;
  assign n6370 = ~n9344 & ~n9345;
  assign n6371 = ~n5941 & ~n5947;
  assign n6372 = n4417 & n4870;
  assign n6373 = ~n9115 & n4424;
  assign n6374 = n4250 & n4432;
  assign n6375 = ~n9116 & n9134;
  assign n6376 = ~n6374 & ~n6375;
  assign n6377 = ~n6373 & n6376;
  assign n6378 = ~n4417 & n6377;
  assign n6379 = ~n4870 & n6377;
  assign n6380 = ~n6378 & ~n6379;
  assign n6381 = ~n6372 & n6377;
  assign n6382 = n8725 & ~n9346;
  assign n6383 = ~n8725 & n9346;
  assign n6384 = ~n6382 & ~n6383;
  assign n6385 = ~n1021 & ~n4274;
  assign n6386 = n4462 & n4666;
  assign n6387 = ~n9117 & n4472;
  assign n6388 = ~n9118 & n4470;
  assign n6389 = n4271 & n9151;
  assign n6390 = ~n6388 & ~n6389;
  assign n6391 = ~n6387 & n6390;
  assign n6392 = ~n6386 & n6391;
  assign n6393 = n6385 & ~n6392;
  assign n6394 = ~n6385 & n6392;
  assign n6395 = ~n6393 & ~n6394;
  assign n6396 = ~n1021 & ~n9119;
  assign n6397 = n5920 & n6396;
  assign n6398 = ~n5925 & ~n6397;
  assign n6399 = n6395 & ~n6398;
  assign n6400 = ~n6395 & n6398;
  assign n6401 = ~n6398 & ~n6399;
  assign n6402 = ~n6395 & ~n6398;
  assign n6403 = n6395 & ~n6399;
  assign n6404 = n6395 & n6398;
  assign n6405 = ~n9347 & ~n9348;
  assign n6406 = ~n6399 & ~n6400;
  assign n6407 = n6384 & ~n9349;
  assign n6408 = ~n6384 & n9349;
  assign n6409 = ~n9349 & ~n6407;
  assign n6410 = ~n6384 & ~n9349;
  assign n6411 = n6384 & ~n6407;
  assign n6412 = n6384 & n9349;
  assign n6413 = ~n9350 & ~n9351;
  assign n6414 = ~n6407 & ~n6408;
  assign n6415 = ~n6371 & ~n9352;
  assign n6416 = n6371 & n9352;
  assign n6417 = ~n6371 & ~n6415;
  assign n6418 = ~n6371 & n9352;
  assign n6419 = ~n9352 & ~n6415;
  assign n6420 = n6371 & ~n9352;
  assign n6421 = ~n9353 & ~n9354;
  assign n6422 = ~n6415 & ~n6416;
  assign n6423 = ~n6370 & ~n9355;
  assign n6424 = n6370 & n9355;
  assign n6425 = ~n6370 & ~n6423;
  assign n6426 = ~n9355 & ~n6423;
  assign n6427 = ~n6425 & ~n6426;
  assign n6428 = ~n6423 & ~n6424;
  assign n6429 = n6357 & n9356;
  assign n6430 = ~n6357 & ~n9356;
  assign n6431 = ~n6429 & ~n6430;
  assign n6432 = n90 & n5466;
  assign n6433 = n4384 & n9246;
  assign n6434 = n4397 & ~n5405;
  assign n6435 = n9129 & n9233;
  assign n6436 = ~n6434 & ~n6435;
  assign n6437 = ~n6433 & n6436;
  assign n6438 = ~n90 & n6437;
  assign n6439 = ~n5466 & n6437;
  assign n6440 = ~n6438 & ~n6439;
  assign n6441 = ~n6432 & n6437;
  assign n6442 = n8620 & ~n9357;
  assign n6443 = ~n8620 & n9357;
  assign n6444 = ~n6442 & ~n6443;
  assign n6445 = n6431 & n6444;
  assign n6446 = ~n6431 & ~n6444;
  assign n6447 = n6431 & ~n6445;
  assign n6448 = n6444 & ~n6445;
  assign n6449 = ~n6447 & ~n6448;
  assign n6450 = ~n6445 & ~n6446;
  assign n6451 = ~n6356 & ~n9358;
  assign n6452 = n6356 & n9358;
  assign n6453 = ~n6356 & ~n6451;
  assign n6454 = ~n9358 & ~n6451;
  assign n6455 = ~n6453 & ~n6454;
  assign n6456 = ~n6451 & ~n6452;
  assign n6457 = ~n6355 & ~n9359;
  assign n6458 = n6355 & n9359;
  assign n6459 = ~n6355 & ~n6457;
  assign n6460 = ~n9359 & ~n6457;
  assign n6461 = ~n6459 & ~n6460;
  assign n6462 = ~n6457 & ~n6458;
  assign n6463 = n6288 & n9360;
  assign n6464 = ~n6288 & ~n9360;
  assign n6465 = ~n6463 & ~n6464;
  assign n6466 = ~n330 & ~n444;
  assign n6467 = ~n398 & n6466;
  assign n6468 = n385 & n1392;
  assign n6469 = n6467 & n6468;
  assign n6470 = ~n229 & ~n287;
  assign n6471 = ~n938 & n6470;
  assign n6472 = ~n817 & n6471;
  assign n6473 = n2233 & n6470;
  assign n6474 = ~n314 & n3604;
  assign n6475 = n9361 & n6474;
  assign n6476 = n6469 & n6475;
  assign n6477 = n4185 & n5146;
  assign n6478 = n6073 & n6477;
  assign n6479 = ~n314 & ~n330;
  assign n6480 = ~n270 & n6479;
  assign n6481 = n9228 & n6480;
  assign n6482 = n9361 & n6481;
  assign n6483 = ~n398 & ~n444;
  assign n6484 = n385 & n6483;
  assign n6485 = n1392 & n3604;
  assign n6486 = n6484 & n6485;
  assign n6487 = n6073 & n6486;
  assign n6488 = n6482 & n6487;
  assign n6489 = n6476 & n6478;
  assign n6490 = n9035 & n9362;
  assign n6491 = n9035 & n6485;
  assign n6492 = n9303 & n6491;
  assign n6493 = n385 & n6492;
  assign n6494 = n9361 & n6493;
  assign n6495 = n9230 & n6494;
  assign n6496 = n9228 & n6495;
  assign n6497 = ~n314 & n6496;
  assign n6498 = ~n330 & n6497;
  assign n6499 = ~n270 & n6498;
  assign n6500 = ~n444 & n6499;
  assign n6501 = ~n821 & n6500;
  assign n6502 = ~n398 & n6501;
  assign n6503 = n9303 & n6490;
  assign n6504 = ~n6465 & n9363;
  assign n6505 = n6465 & ~n9363;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = ~n6287 & n6506;
  assign n6508 = n6287 & ~n6506;
  assign n6509 = ~n6507 & ~n6508;
  assign n6510 = n6272 & n6509;
  assign n6511 = ~n6272 & ~n6509;
  assign n6512 = ~n6510 & ~n6511;
  assign n6513 = n6286 & ~n6512;
  assign n6514 = n6286 & ~n6509;
  assign n6515 = ~n6286 & n6512;
  assign n6516 = ~n9364 & ~n6515;
  assign n6517 = ~n6505 & ~n6507;
  assign n6518 = ~n6457 & ~n6464;
  assign n6519 = n9337 & n6339;
  assign n6520 = n9283 & ~n5880;
  assign n6521 = ~n5875 & ~n5880;
  assign n6522 = ~n9337 & n9365;
  assign n6523 = n9283 & ~n6339;
  assign n6524 = ~n9337 & ~n6523;
  assign n6525 = n9337 & ~n6339;
  assign n6526 = ~n6524 & ~n6525;
  assign n6527 = ~n6519 & ~n6522;
  assign n6528 = n5346 & n9366;
  assign n6529 = n9252 & n5875;
  assign n6530 = n9252 & ~n9283;
  assign n6531 = n5448 & ~n9337;
  assign n6532 = ~n9367 & ~n6531;
  assign n6533 = ~n6528 & n6532;
  assign n6534 = ~n83 & ~n6533;
  assign n6535 = ~n6533 & ~n6534;
  assign n6536 = n83 & ~n6533;
  assign n6537 = ~n83 & ~n6534;
  assign n6538 = ~n83 & n6533;
  assign n6539 = ~n9368 & ~n9369;
  assign n6540 = ~n6445 & ~n6451;
  assign n6541 = ~n6423 & ~n6430;
  assign n6542 = n4612 & n5248;
  assign n6543 = n4616 & n9233;
  assign n6544 = ~n4376 & n4629;
  assign n6545 = ~n9114 & n9158;
  assign n6546 = ~n6544 & ~n6545;
  assign n6547 = ~n6543 & n6546;
  assign n6548 = ~n6542 & n6547;
  assign n6549 = ~n854 & ~n6548;
  assign n6550 = ~n6548 & ~n6549;
  assign n6551 = n854 & ~n6548;
  assign n6552 = ~n854 & ~n6549;
  assign n6553 = ~n854 & n6548;
  assign n6554 = ~n9370 & ~n9371;
  assign n6555 = ~n6407 & ~n6415;
  assign n6556 = n4417 & n4916;
  assign n6557 = n4163 & n4424;
  assign n6558 = n4250 & n9134;
  assign n6559 = ~n9115 & n4432;
  assign n6560 = ~n6558 & ~n6559;
  assign n6561 = ~n6557 & n6560;
  assign n6562 = ~n4417 & n6561;
  assign n6563 = ~n4916 & n6561;
  assign n6564 = ~n6562 & ~n6563;
  assign n6565 = ~n6556 & n6561;
  assign n6566 = n8725 & ~n9372;
  assign n6567 = ~n8725 & n9372;
  assign n6568 = ~n6566 & ~n6567;
  assign n6569 = ~n1021 & ~n4271;
  assign n6570 = n4462 & n4647;
  assign n6571 = ~n9116 & n4472;
  assign n6572 = ~n9117 & n4470;
  assign n6573 = ~n9118 & n9151;
  assign n6574 = ~n6572 & ~n6573;
  assign n6575 = ~n6571 & n6574;
  assign n6576 = ~n6570 & n6575;
  assign n6577 = n6569 & ~n6576;
  assign n6578 = ~n6569 & n6576;
  assign n6579 = ~n6577 & ~n6578;
  assign n6580 = ~n1021 & n4274;
  assign n6581 = ~n1021 & n6392;
  assign n6582 = n4274 & n6581;
  assign n6583 = n6392 & n6580;
  assign n6584 = ~n6399 & ~n9373;
  assign n6585 = n6579 & ~n6584;
  assign n6586 = ~n6579 & n6584;
  assign n6587 = ~n6584 & ~n6585;
  assign n6588 = ~n6579 & ~n6584;
  assign n6589 = n6579 & ~n6585;
  assign n6590 = n6579 & n6584;
  assign n6591 = ~n9374 & ~n9375;
  assign n6592 = ~n6585 & ~n6586;
  assign n6593 = n6568 & ~n9376;
  assign n6594 = ~n6568 & n9376;
  assign n6595 = ~n9376 & ~n6593;
  assign n6596 = ~n6568 & ~n9376;
  assign n6597 = n6568 & ~n6593;
  assign n6598 = n6568 & n9376;
  assign n6599 = ~n9377 & ~n9378;
  assign n6600 = ~n6593 & ~n6594;
  assign n6601 = ~n6555 & ~n9379;
  assign n6602 = n6555 & n9379;
  assign n6603 = ~n6555 & ~n6601;
  assign n6604 = ~n6555 & n9379;
  assign n6605 = ~n9379 & ~n6601;
  assign n6606 = n6555 & ~n9379;
  assign n6607 = ~n9380 & ~n9381;
  assign n6608 = ~n6601 & ~n6602;
  assign n6609 = ~n6554 & ~n9382;
  assign n6610 = n6554 & n9382;
  assign n6611 = ~n6554 & ~n6609;
  assign n6612 = ~n9382 & ~n6609;
  assign n6613 = ~n6611 & ~n6612;
  assign n6614 = ~n6609 & ~n6610;
  assign n6615 = n6541 & n9383;
  assign n6616 = ~n6541 & ~n9383;
  assign n6617 = ~n6615 & ~n6616;
  assign n6618 = n90 & n5444;
  assign n6619 = n4384 & ~n5437;
  assign n6620 = n4397 & n9246;
  assign n6621 = n9129 & ~n5405;
  assign n6622 = ~n6620 & ~n6621;
  assign n6623 = ~n6619 & n6622;
  assign n6624 = ~n90 & n6623;
  assign n6625 = ~n5444 & n6623;
  assign n6626 = ~n6624 & ~n6625;
  assign n6627 = ~n6618 & n6623;
  assign n6628 = n8620 & ~n9384;
  assign n6629 = ~n8620 & n9384;
  assign n6630 = ~n6628 & ~n6629;
  assign n6631 = n6617 & n6630;
  assign n6632 = ~n6617 & ~n6630;
  assign n6633 = n6617 & ~n6631;
  assign n6634 = n6630 & ~n6631;
  assign n6635 = ~n6633 & ~n6634;
  assign n6636 = ~n6631 & ~n6632;
  assign n6637 = ~n6540 & ~n9385;
  assign n6638 = n6540 & n9385;
  assign n6639 = ~n6540 & ~n6637;
  assign n6640 = ~n9385 & ~n6637;
  assign n6641 = ~n6639 & ~n6640;
  assign n6642 = ~n6637 & ~n6638;
  assign n6643 = ~n6539 & ~n9386;
  assign n6644 = n6539 & n9386;
  assign n6645 = ~n6539 & ~n6643;
  assign n6646 = ~n9386 & ~n6643;
  assign n6647 = ~n6645 & ~n6646;
  assign n6648 = ~n6643 & ~n6644;
  assign n6649 = ~n6518 & ~n9387;
  assign n6650 = n6518 & n9387;
  assign n6651 = ~n6518 & n9387;
  assign n6652 = n6518 & ~n9387;
  assign n6653 = ~n6651 & ~n6652;
  assign n6654 = ~n6649 & ~n6650;
  assign n6655 = ~n240 & ~n279;
  assign n6656 = ~n279 & ~n384;
  assign n6657 = ~n240 & n6656;
  assign n6658 = ~n384 & n6655;
  assign n6659 = n1801 & n4165;
  assign n6660 = ~n207 & n4165;
  assign n6661 = ~n240 & n6660;
  assign n6662 = ~n279 & n6661;
  assign n6663 = ~n386 & n6662;
  assign n6664 = ~n384 & n6663;
  assign n6665 = n9389 & n6659;
  assign n6666 = ~n288 & ~n1163;
  assign n6667 = n254 & n6666;
  assign n6668 = n1332 & n6667;
  assign n6669 = ~n865 & ~n876;
  assign n6670 = ~n436 & n6669;
  assign n6671 = n8773 & n6670;
  assign n6672 = ~n288 & ~n436;
  assign n6673 = n254 & n6672;
  assign n6674 = n1332 & n6673;
  assign n6675 = ~n1163 & n6669;
  assign n6676 = n8773 & n6675;
  assign n6677 = n6674 & n6676;
  assign n6678 = n6668 & n6671;
  assign n6679 = n9390 & n9391;
  assign n6680 = n8757 & n6679;
  assign n6681 = n254 & n8773;
  assign n6682 = n8757 & n6681;
  assign n6683 = n9390 & n6682;
  assign n6684 = n9310 & n6683;
  assign n6685 = ~n288 & n6684;
  assign n6686 = ~n865 & n6685;
  assign n6687 = ~n436 & n6686;
  assign n6688 = ~n382 & n6687;
  assign n6689 = ~n876 & n6688;
  assign n6690 = ~n417 & n6689;
  assign n6691 = ~n1163 & n6690;
  assign n6692 = n9310 & n6680;
  assign n6693 = ~n9388 & ~n9392;
  assign n6694 = n9388 & n9392;
  assign n6695 = ~n6693 & ~n6694;
  assign n6696 = ~n6517 & ~n6694;
  assign n6697 = ~n6693 & n6696;
  assign n6698 = ~n6517 & n6695;
  assign n6699 = n6517 & ~n6695;
  assign n6700 = ~n6517 & ~n9393;
  assign n6701 = ~n6693 & ~n9393;
  assign n6702 = ~n6694 & n6701;
  assign n6703 = ~n6700 & ~n6702;
  assign n6704 = ~n9393 & ~n6699;
  assign n6705 = ~n6510 & n9394;
  assign n6706 = n6510 & ~n9394;
  assign n6707 = ~n6705 & ~n6706;
  assign n6708 = n9331 & ~n6512;
  assign n6709 = ~n9332 & ~n6708;
  assign n6710 = n6707 & ~n6709;
  assign n6711 = ~n6707 & n6709;
  assign n6712 = ~n6710 & ~n6711;
  assign n6713 = ~n6707 & n6708;
  assign n6714 = ~n9332 & ~n6713;
  assign n6715 = ~n6643 & ~n6649;
  assign n6716 = ~n6631 & ~n6637;
  assign n6717 = n5346 & ~n9365;
  assign n6718 = ~n9252 & ~n6717;
  assign n6719 = n9252 & ~n9337;
  assign n6720 = n5346 & n6524;
  assign n6721 = ~n6719 & ~n6720;
  assign n6722 = ~n9337 & ~n6718;
  assign n6723 = ~n83 & ~n9395;
  assign n6724 = ~n9395 & ~n6723;
  assign n6725 = n83 & ~n9395;
  assign n6726 = ~n83 & ~n6723;
  assign n6727 = ~n83 & n9395;
  assign n6728 = ~n9396 & ~n9397;
  assign n6729 = ~n6609 & ~n6616;
  assign n6730 = n4612 & n5484;
  assign n6731 = n4616 & ~n5405;
  assign n6732 = n4629 & n9233;
  assign n6733 = ~n4376 & n9158;
  assign n6734 = ~n6732 & ~n6733;
  assign n6735 = ~n6731 & n6734;
  assign n6736 = ~n6730 & n6735;
  assign n6737 = ~n854 & ~n6736;
  assign n6738 = ~n6736 & ~n6737;
  assign n6739 = n854 & ~n6736;
  assign n6740 = ~n854 & ~n6737;
  assign n6741 = ~n854 & n6736;
  assign n6742 = ~n9398 & ~n9399;
  assign n6743 = ~n6593 & ~n6601;
  assign n6744 = n4417 & n4898;
  assign n6745 = ~n9114 & n4424;
  assign n6746 = n4163 & n4432;
  assign n6747 = ~n9115 & n9134;
  assign n6748 = ~n6746 & ~n6747;
  assign n6749 = ~n6745 & n6748;
  assign n6750 = ~n4417 & n6749;
  assign n6751 = ~n4898 & n6749;
  assign n6752 = ~n6750 & ~n6751;
  assign n6753 = ~n6744 & n6749;
  assign n6754 = n8725 & ~n9400;
  assign n6755 = ~n8725 & n9400;
  assign n6756 = ~n6754 & ~n6755;
  assign n6757 = ~n1021 & n9118;
  assign n6758 = n4462 & n4614;
  assign n6759 = n4250 & n4472;
  assign n6760 = ~n9117 & n9151;
  assign n6761 = ~n9116 & n4470;
  assign n6762 = ~n6760 & ~n6761;
  assign n6763 = ~n6759 & n6762;
  assign n6764 = ~n6758 & n6763;
  assign n6765 = n6757 & ~n6764;
  assign n6766 = ~n6757 & n6764;
  assign n6767 = ~n6765 & ~n6766;
  assign n6768 = ~n1021 & n4271;
  assign n6769 = ~n1021 & n6576;
  assign n6770 = n4271 & n6769;
  assign n6771 = n6576 & n6768;
  assign n6772 = ~n6585 & ~n9401;
  assign n6773 = n6767 & ~n6772;
  assign n6774 = ~n6767 & n6772;
  assign n6775 = ~n6772 & ~n6773;
  assign n6776 = ~n6767 & ~n6772;
  assign n6777 = n6767 & ~n6773;
  assign n6778 = n6767 & n6772;
  assign n6779 = ~n9402 & ~n9403;
  assign n6780 = ~n6773 & ~n6774;
  assign n6781 = n6756 & ~n9404;
  assign n6782 = ~n6756 & n9404;
  assign n6783 = ~n6781 & ~n6782;
  assign n6784 = ~n6743 & n6783;
  assign n6785 = n6743 & ~n6783;
  assign n6786 = ~n6784 & ~n6785;
  assign n6787 = ~n6742 & n6786;
  assign n6788 = n6742 & ~n6786;
  assign n6789 = ~n6742 & ~n6787;
  assign n6790 = n6786 & ~n6787;
  assign n6791 = ~n6789 & ~n6790;
  assign n6792 = ~n6787 & ~n6788;
  assign n6793 = n6729 & n9405;
  assign n6794 = ~n6729 & ~n9405;
  assign n6795 = ~n6793 & ~n6794;
  assign n6796 = n90 & n5882;
  assign n6797 = n4384 & n5875;
  assign n6798 = n4384 & ~n9283;
  assign n6799 = n4397 & ~n5437;
  assign n6800 = n9129 & n9246;
  assign n6801 = ~n6799 & ~n6800;
  assign n6802 = ~n9406 & n6801;
  assign n6803 = ~n90 & n6802;
  assign n6804 = ~n5882 & n6802;
  assign n6805 = ~n6803 & ~n6804;
  assign n6806 = ~n6796 & n6802;
  assign n6807 = n8620 & ~n9407;
  assign n6808 = ~n8620 & n9407;
  assign n6809 = ~n6807 & ~n6808;
  assign n6810 = n6795 & n6809;
  assign n6811 = ~n6795 & ~n6809;
  assign n6812 = ~n6810 & ~n6811;
  assign n6813 = ~n6728 & n6812;
  assign n6814 = n6728 & ~n6812;
  assign n6815 = ~n6813 & ~n6814;
  assign n6816 = ~n6716 & n6815;
  assign n6817 = n6716 & ~n6815;
  assign n6818 = ~n6816 & ~n6817;
  assign n6819 = ~n6715 & n6818;
  assign n6820 = n6715 & ~n6818;
  assign n6821 = ~n6819 & ~n6820;
  assign n6822 = n8662 & n8733;
  assign n6823 = n9319 & n6822;
  assign n6824 = ~n545 & ~n721;
  assign n6825 = ~n434 & n6824;
  assign n6826 = ~n340 & ~n817;
  assign n6827 = n272 & n6826;
  assign n6828 = n6825 & n6827;
  assign n6829 = n791 & n6474;
  assign n6830 = ~n434 & ~n545;
  assign n6831 = n272 & n6830;
  assign n6832 = n3604 & n6831;
  assign n6833 = ~n721 & ~n817;
  assign n6834 = ~n314 & ~n340;
  assign n6835 = n6833 & n6834;
  assign n6836 = n791 & n6835;
  assign n6837 = n6832 & n6836;
  assign n6838 = n6828 & n6829;
  assign n6839 = n9037 & n9408;
  assign n6840 = n6823 & n6839;
  assign n6841 = n3604 & n9319;
  assign n6842 = n272 & n6841;
  assign n6843 = n791 & n6842;
  assign n6844 = n9037 & n6843;
  assign n6845 = n8888 & n6844;
  assign n6846 = n8662 & n6845;
  assign n6847 = n8733 & n6846;
  assign n6848 = ~n340 & n6847;
  assign n6849 = ~n314 & n6848;
  assign n6850 = ~n545 & n6849;
  assign n6851 = ~n721 & n6850;
  assign n6852 = ~n817 & n6851;
  assign n6853 = ~n434 & n6852;
  assign n6854 = n8888 & n6840;
  assign n6855 = n6821 & ~n9409;
  assign n6856 = ~n6821 & n9409;
  assign n6857 = ~n9409 & ~n6855;
  assign n6858 = n6821 & ~n6855;
  assign n6859 = ~n6857 & ~n6858;
  assign n6860 = ~n6855 & ~n6856;
  assign n6861 = ~n6701 & ~n9410;
  assign n6862 = n6701 & ~n6858;
  assign n6863 = ~n6857 & n6862;
  assign n6864 = n6701 & n9410;
  assign n6865 = ~n6861 & ~n9411;
  assign n6866 = n6706 & n6865;
  assign n6867 = ~n6706 & ~n6865;
  assign n6868 = n6865 & ~n6866;
  assign n6869 = n6706 & ~n6866;
  assign n6870 = ~n6868 & ~n6869;
  assign n6871 = ~n6866 & ~n6867;
  assign n6872 = n6714 & ~n9412;
  assign n6873 = ~n6714 & n9412;
  assign po3  = ~n6872 & ~n6873;
  assign n6875 = ~n6855 & ~n6861;
  assign n6876 = ~n6816 & ~n6819;
  assign n6877 = ~n6810 & ~n6813;
  assign n6878 = ~n6787 & ~n6794;
  assign n6879 = n4612 & n5466;
  assign n6880 = n4616 & n9246;
  assign n6881 = n4629 & ~n5405;
  assign n6882 = n9158 & n9233;
  assign n6883 = ~n6881 & ~n6882;
  assign n6884 = ~n6880 & n6883;
  assign n6885 = ~n6879 & n6884;
  assign n6886 = ~n854 & ~n6885;
  assign n6887 = ~n854 & ~n6886;
  assign n6888 = ~n854 & n6885;
  assign n6889 = ~n6885 & ~n6886;
  assign n6890 = n854 & ~n6885;
  assign n6891 = ~n9413 & ~n9414;
  assign n6892 = ~n6781 & ~n6784;
  assign n6893 = n4382 & n4417;
  assign n6894 = ~n4376 & n4424;
  assign n6895 = n4163 & n9134;
  assign n6896 = ~n9114 & n4432;
  assign n6897 = ~n6895 & ~n6896;
  assign n6898 = ~n6894 & n6897;
  assign n6899 = ~n6893 & n6898;
  assign n6900 = ~n8725 & ~n6899;
  assign n6901 = n8725 & n6899;
  assign n6902 = ~n6900 & ~n6901;
  assign n6903 = n4462 & n4870;
  assign n6904 = ~n9115 & n4472;
  assign n6905 = n4250 & n4470;
  assign n6906 = ~n9116 & n9151;
  assign n6907 = ~n6905 & ~n6906;
  assign n6908 = ~n6904 & n6907;
  assign n6909 = ~n6903 & n6908;
  assign n6910 = ~n1021 & ~n6909;
  assign n6911 = ~n6909 & ~n6910;
  assign n6912 = n1021 & ~n6909;
  assign n6913 = ~n1021 & ~n6910;
  assign n6914 = ~n1021 & n6909;
  assign n6915 = ~n9415 & ~n9416;
  assign n6916 = ~n83 & ~n1021;
  assign n6917 = ~n1021 & ~n9117;
  assign n6918 = ~n83 & n6917;
  assign n6919 = ~n9117 & n6916;
  assign n6920 = n83 & ~n6917;
  assign n6921 = ~n83 & ~n9417;
  assign n6922 = ~n9117 & ~n9417;
  assign n6923 = ~n1021 & n6922;
  assign n6924 = ~n6921 & ~n6923;
  assign n6925 = ~n9417 & ~n6920;
  assign n6926 = ~n6915 & ~n9418;
  assign n6927 = n6915 & n9418;
  assign n6928 = ~n6915 & ~n6926;
  assign n6929 = ~n9418 & ~n6926;
  assign n6930 = ~n6928 & ~n6929;
  assign n6931 = ~n6926 & ~n6927;
  assign n6932 = ~n1021 & ~n9118;
  assign n6933 = n6764 & n6932;
  assign n6934 = ~n6773 & ~n6933;
  assign n6935 = ~n9419 & ~n6934;
  assign n6936 = n9419 & n6934;
  assign n6937 = n9419 & ~n6934;
  assign n6938 = ~n9419 & n6934;
  assign n6939 = ~n6937 & ~n6938;
  assign n6940 = ~n6935 & ~n6936;
  assign n6941 = n6902 & ~n9420;
  assign n6942 = ~n6902 & n9420;
  assign n6943 = ~n9420 & ~n6941;
  assign n6944 = ~n6902 & ~n9420;
  assign n6945 = n6902 & ~n6941;
  assign n6946 = n6902 & n9420;
  assign n6947 = ~n9421 & ~n9422;
  assign n6948 = ~n6941 & ~n6942;
  assign n6949 = ~n6892 & ~n9423;
  assign n6950 = n6892 & n9423;
  assign n6951 = ~n6892 & n9423;
  assign n6952 = n6892 & ~n9423;
  assign n6953 = ~n6951 & ~n6952;
  assign n6954 = ~n6949 & ~n6950;
  assign n6955 = ~n6891 & ~n9424;
  assign n6956 = n6891 & n9424;
  assign n6957 = ~n6955 & ~n6956;
  assign n6958 = ~n6878 & n6957;
  assign n6959 = n6878 & ~n6957;
  assign n6960 = ~n6958 & ~n6959;
  assign n6961 = n90 & n6341;
  assign n6962 = n4384 & ~n9337;
  assign n6963 = n4397 & n5875;
  assign n6964 = n4397 & ~n9283;
  assign n6965 = n9129 & ~n5437;
  assign n6966 = ~n9425 & ~n6965;
  assign n6967 = ~n6962 & n6966;
  assign n6968 = ~n6961 & n6967;
  assign n6969 = ~n8620 & ~n6968;
  assign n6970 = n8620 & n6968;
  assign n6971 = ~n6969 & ~n6970;
  assign n6972 = n6960 & n6971;
  assign n6973 = ~n6960 & ~n6971;
  assign n6974 = ~n6972 & ~n6973;
  assign n6975 = ~n6877 & n6974;
  assign n6976 = n6877 & ~n6974;
  assign n6977 = ~n6975 & ~n6976;
  assign n6978 = n6876 & ~n6977;
  assign n6979 = ~n6876 & n6977;
  assign n6980 = ~n6978 & ~n6979;
  assign n6981 = n1403 & n4165;
  assign n6982 = n1233 & n6981;
  assign n6983 = ~n313 & ~n331;
  assign n6984 = ~n747 & ~n821;
  assign n6985 = n6983 & n6984;
  assign n6986 = n3812 & n6985;
  assign n6987 = n822 & n3811;
  assign n6988 = n4165 & n6987;
  assign n6989 = ~n313 & ~n747;
  assign n6990 = ~n331 & n6989;
  assign n6991 = n1233 & n1403;
  assign n6992 = n6990 & n6991;
  assign n6993 = n6988 & n6992;
  assign n6994 = n6982 & n6986;
  assign n6995 = n8681 & n9426;
  assign n6996 = n8659 & n6995;
  assign n6997 = n822 & n4165;
  assign n6998 = n1233 & n6997;
  assign n6999 = n9078 & n6998;
  assign n7000 = n8681 & n6999;
  assign n7001 = n8659 & n7000;
  assign n7002 = n1403 & n7001;
  assign n7003 = n3811 & n7002;
  assign n7004 = ~n313 & n7003;
  assign n7005 = ~n331 & n7004;
  assign n7006 = ~n747 & n7005;
  assign n7007 = n9078 & n6996;
  assign n7008 = ~n6980 & n9427;
  assign n7009 = n6980 & ~n9427;
  assign n7010 = ~n7008 & ~n7009;
  assign n7011 = ~n6875 & n7010;
  assign n7012 = n6875 & ~n7010;
  assign n7013 = ~n7011 & ~n7012;
  assign n7014 = ~n6866 & ~n7013;
  assign n7015 = n6866 & n7013;
  assign n7016 = ~n7014 & ~n7015;
  assign n7017 = n6713 & n9412;
  assign n7018 = ~n9332 & ~n7017;
  assign n7019 = n7016 & ~n7018;
  assign n7020 = ~n7016 & n7018;
  assign n7021 = ~n7019 & ~n7020;
  assign n7022 = ~n7009 & ~n7011;
  assign n7023 = ~n6975 & ~n6979;
  assign n7024 = ~n6958 & ~n6972;
  assign n7025 = n90 & n9366;
  assign n7026 = n9129 & n5875;
  assign n7027 = n9129 & ~n9283;
  assign n7028 = n4397 & ~n9337;
  assign n7029 = ~n9428 & ~n7028;
  assign n7030 = ~n7025 & n7029;
  assign n7031 = ~n8620 & ~n7030;
  assign n7032 = n8620 & n7030;
  assign n7033 = ~n7031 & ~n7032;
  assign n7034 = ~n6949 & ~n6955;
  assign n7035 = n4612 & n5444;
  assign n7036 = n4616 & ~n5437;
  assign n7037 = n4629 & n9246;
  assign n7038 = n9158 & ~n5405;
  assign n7039 = ~n7037 & ~n7038;
  assign n7040 = ~n7036 & n7039;
  assign n7041 = ~n7035 & n7040;
  assign n7042 = ~n854 & ~n7041;
  assign n7043 = ~n7041 & ~n7042;
  assign n7044 = n854 & ~n7041;
  assign n7045 = ~n854 & ~n7042;
  assign n7046 = ~n854 & n7041;
  assign n7047 = ~n9429 & ~n9430;
  assign n7048 = ~n6935 & ~n6941;
  assign n7049 = n4417 & n5248;
  assign n7050 = n4424 & n9233;
  assign n7051 = ~n4376 & n4432;
  assign n7052 = ~n9114 & n9134;
  assign n7053 = ~n7051 & ~n7052;
  assign n7054 = ~n7050 & n7053;
  assign n7055 = ~n7049 & n7054;
  assign n7056 = ~n8725 & ~n7055;
  assign n7057 = n8725 & n7055;
  assign n7058 = ~n7056 & ~n7057;
  assign n7059 = n4462 & n4916;
  assign n7060 = n4163 & n4472;
  assign n7061 = n4250 & n9151;
  assign n7062 = ~n9115 & n4470;
  assign n7063 = ~n7061 & ~n7062;
  assign n7064 = ~n7060 & n7063;
  assign n7065 = ~n4462 & n7064;
  assign n7066 = ~n4916 & n7064;
  assign n7067 = ~n7065 & ~n7066;
  assign n7068 = ~n7059 & n7064;
  assign n7069 = n1021 & ~n9431;
  assign n7070 = ~n1021 & n9431;
  assign n7071 = ~n7069 & ~n7070;
  assign n7072 = ~n9417 & ~n6926;
  assign n7073 = ~n1021 & ~n9116;
  assign n7074 = ~n83 & n7073;
  assign n7075 = ~n9116 & n6916;
  assign n7076 = n83 & ~n7073;
  assign n7077 = ~n83 & ~n9432;
  assign n7078 = ~n9116 & ~n9432;
  assign n7079 = ~n1021 & n7078;
  assign n7080 = ~n7077 & ~n7079;
  assign n7081 = ~n9432 & ~n7076;
  assign n7082 = ~n7072 & ~n9433;
  assign n7083 = n7072 & n9433;
  assign n7084 = ~n7072 & ~n7082;
  assign n7085 = ~n9433 & ~n7082;
  assign n7086 = ~n7084 & ~n7085;
  assign n7087 = ~n7082 & ~n7083;
  assign n7088 = n7071 & ~n9434;
  assign n7089 = ~n7071 & n9434;
  assign n7090 = ~n9434 & ~n7088;
  assign n7091 = n7071 & ~n7088;
  assign n7092 = ~n7090 & ~n7091;
  assign n7093 = ~n7088 & ~n7089;
  assign n7094 = n7058 & ~n9435;
  assign n7095 = ~n7058 & ~n7091;
  assign n7096 = ~n7090 & n7095;
  assign n7097 = ~n7058 & n9435;
  assign n7098 = ~n7094 & ~n9436;
  assign n7099 = ~n7048 & n7098;
  assign n7100 = n7048 & ~n7098;
  assign n7101 = ~n7048 & ~n7099;
  assign n7102 = n7098 & ~n7099;
  assign n7103 = ~n7101 & ~n7102;
  assign n7104 = ~n7099 & ~n7100;
  assign n7105 = ~n7047 & ~n9437;
  assign n7106 = n7047 & ~n7102;
  assign n7107 = ~n7101 & n7106;
  assign n7108 = n7047 & n9437;
  assign n7109 = ~n7105 & ~n9438;
  assign n7110 = ~n7034 & n7109;
  assign n7111 = n7034 & ~n7109;
  assign n7112 = ~n7034 & ~n7110;
  assign n7113 = n7109 & ~n7110;
  assign n7114 = ~n7112 & ~n7113;
  assign n7115 = ~n7110 & ~n7111;
  assign n7116 = n7033 & ~n9439;
  assign n7117 = ~n7033 & ~n7113;
  assign n7118 = ~n7112 & n7117;
  assign n7119 = ~n7033 & n9439;
  assign n7120 = ~n7116 & ~n9440;
  assign n7121 = ~n7024 & n7120;
  assign n7122 = n7024 & ~n7120;
  assign n7123 = ~n7121 & ~n7122;
  assign n7124 = ~n7023 & n7123;
  assign n7125 = n7023 & ~n7123;
  assign n7126 = ~n7124 & ~n7125;
  assign n7127 = n178 & n3521;
  assign n7128 = ~n340 & ~n492;
  assign n7129 = ~n380 & n7128;
  assign n7130 = ~n340 & n3820;
  assign n7131 = n9361 & n9441;
  assign n7132 = n7127 & n7131;
  assign n7133 = ~n204 & ~n313;
  assign n7134 = ~n197 & ~n480;
  assign n7135 = n7133 & n7134;
  assign n7136 = n291 & n1248;
  assign n7137 = n7135 & n7136;
  assign n7138 = n9044 & n7137;
  assign n7139 = n7132 & n7138;
  assign n7140 = n9229 & n7139;
  assign n7141 = n178 & n1248;
  assign n7142 = n9441 & n7141;
  assign n7143 = n9044 & n7142;
  assign n7144 = n291 & n7143;
  assign n7145 = n9334 & n7144;
  assign n7146 = n9229 & n7145;
  assign n7147 = n9361 & n7146;
  assign n7148 = n3521 & n7147;
  assign n7149 = ~n313 & n7148;
  assign n7150 = ~n197 & n7149;
  assign n7151 = ~n204 & n7150;
  assign n7152 = ~n480 & n7151;
  assign n7153 = n9334 & n7140;
  assign n7154 = ~n7126 & n9442;
  assign n7155 = n7126 & ~n9442;
  assign n7156 = ~n7154 & ~n7155;
  assign n7157 = ~n7022 & n7156;
  assign n7158 = n7022 & ~n7156;
  assign n7159 = ~n7157 & ~n7158;
  assign n7160 = ~n7015 & ~n7159;
  assign n7161 = n7015 & n7159;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = ~n7016 & n7017;
  assign n7164 = ~n9332 & ~n7163;
  assign n7165 = n7162 & ~n7164;
  assign n7166 = ~n7162 & n7164;
  assign n7167 = ~n7165 & ~n7166;
  assign n7168 = ~n7155 & ~n7157;
  assign n7169 = ~n7121 & ~n7124;
  assign n7170 = ~n7110 & ~n7116;
  assign n7171 = ~n7099 & ~n7105;
  assign n7172 = n90 & ~n9365;
  assign n7173 = ~n9129 & ~n7172;
  assign n7174 = n9129 & ~n9337;
  assign n7175 = n90 & n6524;
  assign n7176 = ~n7174 & ~n7175;
  assign n7177 = ~n9337 & ~n7173;
  assign n7178 = n8620 & ~n9443;
  assign n7179 = ~n8620 & n9443;
  assign n7180 = ~n7178 & ~n7179;
  assign n7181 = ~n7171 & ~n7180;
  assign n7182 = n7171 & n7180;
  assign n7183 = ~n7181 & ~n7182;
  assign n7184 = n4612 & n5882;
  assign n7185 = n4616 & n5875;
  assign n7186 = n4616 & ~n9283;
  assign n7187 = n4629 & ~n5437;
  assign n7188 = n9158 & n9246;
  assign n7189 = ~n7187 & ~n7188;
  assign n7190 = ~n9444 & n7189;
  assign n7191 = ~n7184 & n7190;
  assign n7192 = ~n854 & ~n7191;
  assign n7193 = ~n7191 & ~n7192;
  assign n7194 = n854 & ~n7191;
  assign n7195 = ~n854 & ~n7192;
  assign n7196 = ~n854 & n7191;
  assign n7197 = ~n9445 & ~n9446;
  assign n7198 = ~n7088 & ~n7094;
  assign n7199 = n4417 & n5484;
  assign n7200 = n4424 & ~n5405;
  assign n7201 = n4432 & n9233;
  assign n7202 = ~n4376 & n9134;
  assign n7203 = ~n7201 & ~n7202;
  assign n7204 = ~n7200 & n7203;
  assign n7205 = ~n7199 & n7204;
  assign n7206 = ~n8725 & ~n7205;
  assign n7207 = n8725 & n7205;
  assign n7208 = ~n7206 & ~n7207;
  assign n7209 = n4462 & n4898;
  assign n7210 = ~n9114 & n4472;
  assign n7211 = n4163 & n4470;
  assign n7212 = ~n9115 & n9151;
  assign n7213 = ~n7211 & ~n7212;
  assign n7214 = ~n7210 & n7213;
  assign n7215 = ~n4462 & n7214;
  assign n7216 = ~n4898 & n7214;
  assign n7217 = ~n7215 & ~n7216;
  assign n7218 = ~n7209 & n7214;
  assign n7219 = n1021 & ~n9447;
  assign n7220 = ~n1021 & n9447;
  assign n7221 = ~n7219 & ~n7220;
  assign n7222 = ~n9432 & ~n7082;
  assign n7223 = ~n1021 & n4250;
  assign n7224 = ~n83 & n7223;
  assign n7225 = n4250 & n6916;
  assign n7226 = n83 & ~n7223;
  assign n7227 = ~n83 & ~n9448;
  assign n7228 = n4250 & ~n9448;
  assign n7229 = ~n1021 & n7228;
  assign n7230 = ~n7227 & ~n7229;
  assign n7231 = ~n9448 & ~n7226;
  assign n7232 = ~n7222 & ~n9449;
  assign n7233 = n7222 & n9449;
  assign n7234 = ~n7222 & ~n7232;
  assign n7235 = ~n9449 & ~n7232;
  assign n7236 = ~n7234 & ~n7235;
  assign n7237 = ~n7232 & ~n7233;
  assign n7238 = n7221 & ~n9450;
  assign n7239 = ~n7221 & n9450;
  assign n7240 = ~n9450 & ~n7238;
  assign n7241 = n7221 & ~n7238;
  assign n7242 = ~n7240 & ~n7241;
  assign n7243 = ~n7238 & ~n7239;
  assign n7244 = n7208 & ~n9451;
  assign n7245 = ~n7208 & ~n7241;
  assign n7246 = ~n7240 & n7245;
  assign n7247 = ~n7208 & n9451;
  assign n7248 = ~n7244 & ~n9452;
  assign n7249 = ~n7198 & n7248;
  assign n7250 = n7198 & ~n7248;
  assign n7251 = ~n7198 & ~n7249;
  assign n7252 = n7248 & ~n7249;
  assign n7253 = ~n7251 & ~n7252;
  assign n7254 = ~n7249 & ~n7250;
  assign n7255 = ~n7197 & ~n9453;
  assign n7256 = n7197 & ~n7252;
  assign n7257 = ~n7251 & n7256;
  assign n7258 = n7197 & n9453;
  assign n7259 = ~n7255 & ~n9454;
  assign n7260 = n7183 & n7259;
  assign n7261 = ~n7183 & ~n7259;
  assign n7262 = ~n7260 & ~n7261;
  assign n7263 = ~n7170 & n7262;
  assign n7264 = n7170 & ~n7262;
  assign n7265 = ~n7263 & ~n7264;
  assign n7266 = ~n7169 & n7265;
  assign n7267 = n7169 & ~n7265;
  assign n7268 = ~n7266 & ~n7267;
  assign n7269 = ~n641 & n1119;
  assign n7270 = n1023 & n7269;
  assign n7271 = n6307 & n7269;
  assign n7272 = n1023 & n7271;
  assign n7273 = n6307 & n7270;
  assign n7274 = n1643 & n3521;
  assign n7275 = n3604 & n7274;
  assign n7276 = n9070 & n7275;
  assign n7277 = n687 & n1643;
  assign n7278 = n1023 & n7277;
  assign n7279 = n9070 & n7278;
  assign n7280 = n3604 & n7279;
  assign n7281 = n1119 & n7280;
  assign n7282 = n3521 & n7281;
  assign n7283 = n602 & n7282;
  assign n7284 = ~n641 & n7283;
  assign n7285 = n9455 & n7276;
  assign n7286 = ~n164 & ~n443;
  assign n7287 = ~n362 & ~n636;
  assign n7288 = ~n362 & ~n443;
  assign n7289 = ~n164 & ~n636;
  assign n7290 = n7288 & n7289;
  assign n7291 = n7286 & n7287;
  assign n7292 = n657 & n3525;
  assign n7293 = n5378 & n7292;
  assign n7294 = n9457 & n7293;
  assign n7295 = n9076 & n7294;
  assign n7296 = n9456 & n7295;
  assign n7297 = n657 & n9304;
  assign n7298 = n9076 & n7297;
  assign n7299 = n5378 & n7298;
  assign n7300 = n9456 & n7299;
  assign n7301 = ~n295 & n7300;
  assign n7302 = ~n164 & n7301;
  assign n7303 = ~n443 & n7302;
  assign n7304 = ~n636 & n7303;
  assign n7305 = ~n8664 & n7304;
  assign n7306 = ~n362 & n7305;
  assign n7307 = n9304 & n7296;
  assign n7308 = ~n7268 & n9458;
  assign n7309 = n7268 & ~n9458;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = ~n7168 & n7310;
  assign n7312 = n7168 & ~n7310;
  assign n7313 = ~n7311 & ~n7312;
  assign n7314 = ~n7161 & ~n7313;
  assign n7315 = n7161 & n7313;
  assign n7316 = ~n7314 & ~n7315;
  assign n7317 = ~n7162 & n7163;
  assign n7318 = ~n9332 & ~n7317;
  assign n7319 = n7316 & ~n7318;
  assign n7320 = ~n7316 & n7318;
  assign n7321 = ~n7319 & ~n7320;
  assign n7322 = ~n7309 & ~n7311;
  assign n7323 = ~n7263 & ~n7266;
  assign n7324 = ~n7181 & ~n7260;
  assign n7325 = ~n7249 & ~n7255;
  assign n7326 = n4612 & n6341;
  assign n7327 = n4616 & ~n9337;
  assign n7328 = n4629 & n5875;
  assign n7329 = n4629 & ~n9283;
  assign n7330 = n9158 & ~n5437;
  assign n7331 = ~n9459 & ~n7330;
  assign n7332 = ~n7327 & n7331;
  assign n7333 = ~n6341 & n7332;
  assign n7334 = ~n4612 & n7332;
  assign n7335 = ~n7333 & ~n7334;
  assign n7336 = ~n7326 & n7332;
  assign n7337 = n854 & ~n9460;
  assign n7338 = ~n854 & n9460;
  assign n7339 = ~n7337 & ~n7338;
  assign n7340 = ~n7325 & n7339;
  assign n7341 = n7325 & ~n7339;
  assign n7342 = ~n7340 & ~n7341;
  assign n7343 = ~n7238 & ~n7244;
  assign n7344 = n4417 & n5466;
  assign n7345 = n4424 & n9246;
  assign n7346 = n4432 & ~n5405;
  assign n7347 = n9134 & n9233;
  assign n7348 = ~n7346 & ~n7347;
  assign n7349 = ~n7345 & n7348;
  assign n7350 = ~n4417 & n7349;
  assign n7351 = ~n5466 & n7349;
  assign n7352 = ~n7350 & ~n7351;
  assign n7353 = ~n7344 & n7349;
  assign n7354 = n8725 & ~n9461;
  assign n7355 = ~n8725 & n9461;
  assign n7356 = ~n7354 & ~n7355;
  assign n7357 = ~n9448 & ~n7232;
  assign n7358 = n4382 & n4462;
  assign n7359 = ~n4376 & n4472;
  assign n7360 = n4163 & n9151;
  assign n7361 = ~n9114 & n4470;
  assign n7362 = ~n7360 & ~n7361;
  assign n7363 = ~n7359 & n7362;
  assign n7364 = ~n7358 & n7363;
  assign n7365 = ~n1021 & ~n7364;
  assign n7366 = ~n7364 & ~n7365;
  assign n7367 = n1021 & ~n7364;
  assign n7368 = ~n1021 & ~n7365;
  assign n7369 = ~n1021 & n7364;
  assign n7370 = ~n9462 & ~n9463;
  assign n7371 = ~n1021 & ~n9115;
  assign n7372 = n8620 & n83;
  assign n7373 = ~n8620 & ~n83;
  assign n7374 = ~n7372 & ~n7373;
  assign n7375 = n7371 & n7374;
  assign n7376 = ~n7371 & ~n7374;
  assign n7377 = ~n7375 & ~n7376;
  assign n7378 = ~n7370 & n7377;
  assign n7379 = n7370 & ~n7377;
  assign n7380 = ~n7370 & ~n7378;
  assign n7381 = ~n7370 & ~n7377;
  assign n7382 = n7377 & ~n7378;
  assign n7383 = n7370 & n7377;
  assign n7384 = ~n9464 & ~n9465;
  assign n7385 = ~n7378 & ~n7379;
  assign n7386 = ~n7357 & ~n9466;
  assign n7387 = n7357 & n9466;
  assign n7388 = ~n7357 & n9466;
  assign n7389 = n7357 & ~n9466;
  assign n7390 = ~n7388 & ~n7389;
  assign n7391 = ~n7386 & ~n7387;
  assign n7392 = n7356 & ~n9467;
  assign n7393 = ~n7356 & n9467;
  assign n7394 = ~n9467 & ~n7392;
  assign n7395 = n7356 & ~n7392;
  assign n7396 = ~n7394 & ~n7395;
  assign n7397 = ~n7392 & ~n7393;
  assign n7398 = ~n7343 & ~n9468;
  assign n7399 = n7343 & n9468;
  assign n7400 = ~n7343 & ~n7398;
  assign n7401 = ~n9468 & ~n7398;
  assign n7402 = ~n7400 & ~n7401;
  assign n7403 = ~n7398 & ~n7399;
  assign n7404 = n7342 & ~n9469;
  assign n7405 = ~n7342 & n9469;
  assign n7406 = n7342 & ~n7404;
  assign n7407 = ~n9469 & ~n7404;
  assign n7408 = ~n7406 & ~n7407;
  assign n7409 = ~n7404 & ~n7405;
  assign n7410 = ~n7324 & ~n9470;
  assign n7411 = n7324 & n9470;
  assign n7412 = ~n7324 & n9470;
  assign n7413 = n7324 & ~n9470;
  assign n7414 = ~n7412 & ~n7413;
  assign n7415 = ~n7410 & ~n7411;
  assign n7416 = n7323 & n9471;
  assign n7417 = ~n7323 & ~n9471;
  assign n7418 = ~n7416 & ~n7417;
  assign n7419 = n763 & n1232;
  assign n7420 = ~n198 & ~n331;
  assign n7421 = n1602 & n7420;
  assign n7422 = n7419 & n7421;
  assign n7423 = ~n240 & ~n8663;
  assign n7424 = ~n220 & ~n398;
  assign n7425 = ~n220 & ~n8663;
  assign n7426 = ~n240 & ~n398;
  assign n7427 = n7425 & n7426;
  assign n7428 = n7423 & n7424;
  assign n7429 = n9441 & n9472;
  assign n7430 = n7422 & n7429;
  assign n7431 = n9456 & n7430;
  assign n7432 = n763 & n9032;
  assign n7433 = n9441 & n7432;
  assign n7434 = n1232 & n7433;
  assign n7435 = n9456 & n7434;
  assign n7436 = ~n240 & n7435;
  assign n7437 = ~n331 & n7436;
  assign n7438 = ~n220 & n7437;
  assign n7439 = ~n198 & n7438;
  assign n7440 = n1602 & n7439;
  assign n7441 = ~n8663 & n7440;
  assign n7442 = ~n398 & n7441;
  assign n7443 = n9032 & n7431;
  assign n7444 = n7418 & ~n9473;
  assign n7445 = ~n7418 & n9473;
  assign n7446 = ~n7444 & ~n7445;
  assign n7447 = ~n7322 & n7446;
  assign n7448 = n7322 & ~n7446;
  assign n7449 = ~n7447 & ~n7448;
  assign n7450 = n7315 & n7449;
  assign n7451 = ~n7315 & ~n7449;
  assign n7452 = ~n7450 & ~n7451;
  assign n7453 = ~n7316 & n7317;
  assign n7454 = ~n9332 & ~n7453;
  assign n7455 = n7452 & ~n7454;
  assign n7456 = ~n7452 & n7454;
  assign n7457 = ~n7455 & ~n7456;
  assign n7458 = ~n7444 & ~n7447;
  assign n7459 = ~n7410 & ~n7417;
  assign n7460 = ~n7340 & ~n7404;
  assign n7461 = n4612 & n9366;
  assign n7462 = n9158 & n5875;
  assign n7463 = n9158 & ~n9283;
  assign n7464 = n4629 & ~n9337;
  assign n7465 = ~n9474 & ~n7464;
  assign n7466 = ~n7461 & n7465;
  assign n7467 = ~n854 & ~n7466;
  assign n7468 = ~n7466 & ~n7467;
  assign n7469 = n854 & ~n7466;
  assign n7470 = ~n854 & ~n7467;
  assign n7471 = ~n854 & n7466;
  assign n7472 = ~n9475 & ~n9476;
  assign n7473 = ~n7392 & ~n7398;
  assign n7474 = n4417 & n5444;
  assign n7475 = n4424 & ~n5437;
  assign n7476 = n4432 & n9246;
  assign n7477 = n9134 & ~n5405;
  assign n7478 = ~n7476 & ~n7477;
  assign n7479 = ~n7475 & n7478;
  assign n7480 = ~n7474 & n7479;
  assign n7481 = ~n8725 & ~n7480;
  assign n7482 = n8725 & n7480;
  assign n7483 = ~n7481 & ~n7482;
  assign n7484 = ~n7378 & ~n7386;
  assign n7485 = n4462 & n5248;
  assign n7486 = n4472 & n9233;
  assign n7487 = ~n4376 & n4470;
  assign n7488 = ~n9114 & n9151;
  assign n7489 = ~n7487 & ~n7488;
  assign n7490 = ~n7486 & n7489;
  assign n7491 = ~n4462 & n7490;
  assign n7492 = ~n5248 & n7490;
  assign n7493 = ~n7491 & ~n7492;
  assign n7494 = ~n7485 & n7490;
  assign n7495 = n1021 & ~n9477;
  assign n7496 = ~n1021 & n9477;
  assign n7497 = ~n7495 & ~n7496;
  assign n7498 = ~n1021 & n4163;
  assign n7499 = ~n7372 & ~n7375;
  assign n7500 = ~n7498 & ~n7499;
  assign n7501 = n7498 & n7499;
  assign n7502 = ~n7498 & ~n7500;
  assign n7503 = ~n7498 & n7499;
  assign n7504 = ~n7499 & ~n7500;
  assign n7505 = n7498 & ~n7499;
  assign n7506 = ~n9478 & ~n9479;
  assign n7507 = ~n7500 & ~n7501;
  assign n7508 = n7497 & ~n9480;
  assign n7509 = ~n7497 & n9480;
  assign n7510 = ~n7508 & ~n7509;
  assign n7511 = ~n7484 & n7510;
  assign n7512 = n7484 & ~n7510;
  assign n7513 = ~n7484 & ~n7511;
  assign n7514 = n7510 & ~n7511;
  assign n7515 = ~n7513 & ~n7514;
  assign n7516 = ~n7511 & ~n7512;
  assign n7517 = n7483 & ~n9481;
  assign n7518 = ~n7483 & ~n7514;
  assign n7519 = ~n7513 & n7518;
  assign n7520 = ~n7483 & n9481;
  assign n7521 = ~n7517 & ~n9482;
  assign n7522 = ~n7473 & n7521;
  assign n7523 = n7473 & ~n7521;
  assign n7524 = ~n7522 & ~n7523;
  assign n7525 = ~n7472 & n7524;
  assign n7526 = n7472 & ~n7524;
  assign n7527 = ~n7525 & ~n7526;
  assign n7528 = ~n7460 & n7527;
  assign n7529 = n7460 & ~n7527;
  assign n7530 = ~n7528 & ~n7529;
  assign n7531 = ~n7459 & n7530;
  assign n7532 = n7459 & ~n7530;
  assign n7533 = ~n7531 & ~n7532;
  assign n7534 = ~n280 & ~n391;
  assign n7535 = ~n8631 & ~n280;
  assign n7536 = ~n391 & n7535;
  assign n7537 = ~n8631 & n7534;
  assign n7538 = n615 & n863;
  assign n7539 = n3384 & n7538;
  assign n7540 = n9483 & n7539;
  assign n7541 = n9085 & n7540;
  assign n7542 = n615 & n9085;
  assign n7543 = n8744 & n7542;
  assign n7544 = ~n8642 & n7543;
  assign n7545 = ~n8631 & n7544;
  assign n7546 = ~n280 & n7545;
  assign n7547 = ~n158 & n7546;
  assign n7548 = ~n658 & n7547;
  assign n7549 = ~n721 & n7548;
  assign n7550 = ~n391 & n7549;
  assign n7551 = n8744 & n7541;
  assign n7552 = ~n207 & ~n938;
  assign n7553 = ~n884 & n7552;
  assign n7554 = ~n222 & ~n271;
  assign n7555 = n3611 & n7554;
  assign n7556 = ~n271 & ~n938;
  assign n7557 = ~n884 & n7556;
  assign n7558 = ~n207 & ~n222;
  assign n7559 = n3611 & n7558;
  assign n7560 = n7557 & n7559;
  assign n7561 = n7553 & n7555;
  assign n7562 = n8679 & n9053;
  assign n7563 = n9485 & n7562;
  assign n7564 = n8675 & n7563;
  assign n7565 = n9317 & n7564;
  assign n7566 = n8675 & n7562;
  assign n7567 = n9317 & n7566;
  assign n7568 = n9484 & n7567;
  assign n7569 = ~n207 & n7568;
  assign n7570 = ~n222 & n7569;
  assign n7571 = ~n271 & n7570;
  assign n7572 = ~n938 & n7571;
  assign n7573 = ~n884 & n7572;
  assign n7574 = ~n1163 & n7573;
  assign n7575 = ~n656 & n7574;
  assign n7576 = n9484 & n7565;
  assign n7577 = ~n7533 & n9486;
  assign n7578 = n7533 & ~n9486;
  assign n7579 = ~n7577 & ~n7578;
  assign n7580 = ~n7458 & n7579;
  assign n7581 = n7458 & ~n7579;
  assign n7582 = ~n7580 & ~n7581;
  assign n7583 = ~n7450 & ~n7582;
  assign n7584 = n7450 & n7582;
  assign n7585 = ~n7583 & ~n7584;
  assign n7586 = ~n7452 & n7453;
  assign n7587 = ~n9332 & ~n7586;
  assign n7588 = n7585 & ~n7587;
  assign n7589 = ~n7585 & n7587;
  assign n7590 = ~n7588 & ~n7589;
  assign n7591 = ~n7578 & ~n7580;
  assign n7592 = ~n7528 & ~n7531;
  assign n7593 = ~n7522 & ~n7525;
  assign n7594 = ~n7511 & ~n7517;
  assign n7595 = n4612 & ~n9365;
  assign n7596 = ~n9158 & ~n7595;
  assign n7597 = n9158 & ~n9337;
  assign n7598 = n4612 & n6524;
  assign n7599 = ~n7597 & ~n7598;
  assign n7600 = ~n9337 & ~n7596;
  assign n7601 = ~n854 & n9487;
  assign n7602 = n854 & ~n9487;
  assign n7603 = ~n7601 & ~n7602;
  assign n7604 = ~n7594 & ~n7603;
  assign n7605 = n7594 & n7603;
  assign n7606 = ~n7604 & ~n7605;
  assign n7607 = n4417 & n5882;
  assign n7608 = n4424 & n5875;
  assign n7609 = n4424 & ~n9283;
  assign n7610 = n4432 & ~n5437;
  assign n7611 = n9134 & n9246;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = ~n9488 & n7612;
  assign n7614 = ~n7607 & n7613;
  assign n7615 = ~n8725 & ~n7614;
  assign n7616 = n8725 & n7614;
  assign n7617 = ~n7615 & ~n7616;
  assign n7618 = ~n7500 & ~n7508;
  assign n7619 = n4462 & n5484;
  assign n7620 = n4472 & ~n5405;
  assign n7621 = n4470 & n9233;
  assign n7622 = ~n4376 & n9151;
  assign n7623 = ~n7621 & ~n7622;
  assign n7624 = ~n7620 & n7623;
  assign n7625 = ~n7619 & n7624;
  assign n7626 = ~n1021 & ~n7625;
  assign n7627 = ~n7625 & ~n7626;
  assign n7628 = n1021 & ~n7625;
  assign n7629 = ~n1021 & ~n7626;
  assign n7630 = ~n1021 & n7625;
  assign n7631 = ~n9489 & ~n9490;
  assign n7632 = ~n1021 & n4332;
  assign n7633 = ~n7631 & ~n7632;
  assign n7634 = n7631 & n7632;
  assign n7635 = ~n7631 & ~n7633;
  assign n7636 = ~n7632 & ~n7633;
  assign n7637 = ~n7635 & ~n7636;
  assign n7638 = ~n7633 & ~n7634;
  assign n7639 = ~n7618 & ~n9491;
  assign n7640 = n7618 & n9491;
  assign n7641 = ~n7618 & n9491;
  assign n7642 = n7618 & ~n9491;
  assign n7643 = ~n7641 & ~n7642;
  assign n7644 = ~n7639 & ~n7640;
  assign n7645 = n7617 & ~n9492;
  assign n7646 = ~n7617 & n9492;
  assign n7647 = ~n9492 & ~n7645;
  assign n7648 = n7617 & ~n7645;
  assign n7649 = ~n7647 & ~n7648;
  assign n7650 = ~n7645 & ~n7646;
  assign n7651 = n7606 & ~n9493;
  assign n7652 = ~n7606 & n9493;
  assign n7653 = ~n9493 & ~n7651;
  assign n7654 = n7606 & ~n7651;
  assign n7655 = ~n7653 & ~n7654;
  assign n7656 = ~n7651 & ~n7652;
  assign n7657 = ~n7593 & ~n9494;
  assign n7658 = n7593 & n9494;
  assign n7659 = ~n7593 & n9494;
  assign n7660 = n7593 & ~n9494;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = ~n7657 & ~n7658;
  assign n7663 = n7592 & n9495;
  assign n7664 = ~n7592 & ~n9495;
  assign n7665 = ~n7663 & ~n7664;
  assign n7666 = ~n450 & ~n608;
  assign n7667 = ~n158 & ~n642;
  assign n7668 = n7666 & n7667;
  assign n7669 = ~n295 & ~n8647;
  assign n7670 = n1232 & n7669;
  assign n7671 = n5378 & n7670;
  assign n7672 = n7668 & n7671;
  assign n7673 = n8653 & n6477;
  assign n7674 = ~n295 & ~n450;
  assign n7675 = ~n158 & ~n8647;
  assign n7676 = n7674 & n7675;
  assign n7677 = n1232 & n5378;
  assign n7678 = n7676 & n7677;
  assign n7679 = ~n608 & ~n642;
  assign n7680 = ~n270 & n7679;
  assign n7681 = n9228 & n7680;
  assign n7682 = n7678 & n7681;
  assign n7683 = n8653 & n7682;
  assign n7684 = n7672 & n7673;
  assign n7685 = n9305 & n9496;
  assign n7686 = n8653 & n1232;
  assign n7687 = n9305 & n7686;
  assign n7688 = n9228 & n7687;
  assign n7689 = n9071 & n7688;
  assign n7690 = n5378 & n7689;
  assign n7691 = ~n295 & n7690;
  assign n7692 = ~n270 & n7691;
  assign n7693 = ~n158 & n7692;
  assign n7694 = ~n8647 & n7693;
  assign n7695 = ~n642 & n7694;
  assign n7696 = ~n608 & n7695;
  assign n7697 = ~n450 & n7696;
  assign n7698 = n9071 & n7685;
  assign n7699 = ~n7665 & n9497;
  assign n7700 = n7665 & ~n9497;
  assign n7701 = ~n7699 & ~n7700;
  assign n7702 = ~n7591 & n7701;
  assign n7703 = n7591 & ~n7701;
  assign n7704 = ~n7702 & ~n7703;
  assign n7705 = ~n7584 & ~n7704;
  assign n7706 = n7584 & n7704;
  assign n7707 = ~n7705 & ~n7706;
  assign n7708 = ~n7585 & n7586;
  assign n7709 = ~n9332 & ~n7708;
  assign n7710 = n7707 & ~n7709;
  assign n7711 = ~n7707 & n7709;
  assign n7712 = ~n7710 & ~n7711;
  assign n7713 = ~n7700 & ~n7702;
  assign n7714 = ~n7657 & ~n7664;
  assign n7715 = ~n7604 & ~n7651;
  assign n7716 = ~n7639 & ~n7645;
  assign n7717 = n4417 & n6341;
  assign n7718 = n4424 & ~n9337;
  assign n7719 = n4432 & n5875;
  assign n7720 = n4432 & ~n9283;
  assign n7721 = n9134 & ~n5437;
  assign n7722 = ~n9498 & ~n7721;
  assign n7723 = ~n7718 & n7722;
  assign n7724 = ~n4417 & n7723;
  assign n7725 = ~n6341 & n7723;
  assign n7726 = ~n7724 & ~n7725;
  assign n7727 = ~n7717 & n7723;
  assign n7728 = n8725 & ~n9499;
  assign n7729 = ~n8725 & n9499;
  assign n7730 = ~n7728 & ~n7729;
  assign n7731 = ~n7716 & n7730;
  assign n7732 = n7716 & ~n7730;
  assign n7733 = ~n7716 & ~n7731;
  assign n7734 = n7730 & ~n7731;
  assign n7735 = ~n7733 & ~n7734;
  assign n7736 = ~n7731 & ~n7732;
  assign n7737 = n4462 & n5466;
  assign n7738 = n4472 & n9246;
  assign n7739 = n4470 & ~n5405;
  assign n7740 = n9151 & n9233;
  assign n7741 = ~n7739 & ~n7740;
  assign n7742 = ~n7738 & n7741;
  assign n7743 = ~n7737 & n7742;
  assign n7744 = ~n1021 & ~n7743;
  assign n7745 = ~n1021 & ~n7744;
  assign n7746 = ~n1021 & n7743;
  assign n7747 = ~n7743 & ~n7744;
  assign n7748 = n1021 & ~n7743;
  assign n7749 = ~n9501 & ~n9502;
  assign n7750 = ~n1021 & ~n4376;
  assign n7751 = n854 & n7750;
  assign n7752 = ~n854 & ~n7750;
  assign n7753 = ~n7751 & ~n7752;
  assign n7754 = n7498 & ~n7751;
  assign n7755 = ~n7752 & n7754;
  assign n7756 = n7498 & ~n7755;
  assign n7757 = n7498 & ~n7753;
  assign n7758 = ~n7498 & ~n7751;
  assign n7759 = ~n7751 & ~n7755;
  assign n7760 = ~n7752 & ~n7758;
  assign n7761 = ~n7752 & n9504;
  assign n7762 = ~n7498 & n7753;
  assign n7763 = ~n9503 & ~n9505;
  assign n7764 = ~n1021 & ~n4163;
  assign n7765 = ~n9114 & ~n7498;
  assign n7766 = ~n1021 & n7765;
  assign n7767 = ~n9114 & n7764;
  assign n7768 = ~n7633 & ~n9506;
  assign n7769 = ~n7763 & ~n7768;
  assign n7770 = n7763 & n7768;
  assign n7771 = ~n7768 & ~n7769;
  assign n7772 = ~n7763 & ~n7769;
  assign n7773 = ~n7771 & ~n7772;
  assign n7774 = ~n7769 & ~n7770;
  assign n7775 = n7749 & n9507;
  assign n7776 = ~n7749 & ~n9507;
  assign n7777 = ~n9507 & ~n7776;
  assign n7778 = ~n7749 & ~n7776;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = ~n7775 & ~n7776;
  assign n7781 = ~n9500 & ~n9508;
  assign n7782 = ~n7734 & n9508;
  assign n7783 = ~n7733 & n7782;
  assign n7784 = n9500 & n9508;
  assign n7785 = ~n7781 & ~n9509;
  assign n7786 = ~n7715 & n7785;
  assign n7787 = n7715 & ~n7785;
  assign n7788 = ~n7786 & ~n7787;
  assign n7789 = ~n7714 & n7788;
  assign n7790 = n7714 & ~n7788;
  assign n7791 = ~n7789 & ~n7790;
  assign n7792 = n945 & n4166;
  assign n7793 = n5378 & n7792;
  assign n7794 = ~n309 & ~n511;
  assign n7795 = ~n511 & ~n8700;
  assign n7796 = ~n309 & n7795;
  assign n7797 = ~n8700 & n7794;
  assign n7798 = n447 & n9510;
  assign n7799 = n603 & n9230;
  assign n7800 = n7798 & n7799;
  assign n7801 = n7793 & n7800;
  assign n7802 = n8777 & n7801;
  assign n7803 = n8812 & n9321;
  assign n7804 = n8777 & n4166;
  assign n7805 = n447 & n7804;
  assign n7806 = n945 & n7805;
  assign n7807 = n9230 & n7806;
  assign n7808 = n9321 & n7807;
  assign n7809 = n8812 & n7808;
  assign n7810 = n5378 & n7809;
  assign n7811 = n603 & n7810;
  assign n7812 = ~n309 & n7811;
  assign n7813 = ~n8700 & n7812;
  assign n7814 = ~n511 & n7813;
  assign n7815 = n7802 & n7803;
  assign n7816 = ~n7791 & n9511;
  assign n7817 = n7791 & ~n9511;
  assign n7818 = ~n7816 & ~n7817;
  assign n7819 = ~n7713 & n7818;
  assign n7820 = n7713 & ~n7818;
  assign n7821 = ~n7819 & ~n7820;
  assign n7822 = ~n7706 & ~n7821;
  assign n7823 = n7706 & n7821;
  assign n7824 = ~n7822 & ~n7823;
  assign n7825 = ~n7707 & n7708;
  assign n7826 = ~n9332 & ~n7825;
  assign n7827 = n7824 & ~n7826;
  assign n7828 = ~n7824 & n7826;
  assign n7829 = ~n7827 & ~n7828;
  assign n7830 = ~n7817 & ~n7819;
  assign n7831 = ~n7786 & ~n7789;
  assign n7832 = ~n7731 & ~n7781;
  assign n7833 = n4417 & n9366;
  assign n7834 = n9134 & n5875;
  assign n7835 = n9134 & ~n9283;
  assign n7836 = n4432 & ~n9337;
  assign n7837 = ~n9512 & ~n7836;
  assign n7838 = ~n7833 & n7837;
  assign n7839 = ~n8725 & ~n7838;
  assign n7840 = n8725 & n7838;
  assign n7841 = ~n7839 & ~n7840;
  assign n7842 = n4462 & n5444;
  assign n7843 = n4472 & ~n5437;
  assign n7844 = n4470 & n9246;
  assign n7845 = n9151 & ~n5405;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = ~n7843 & n7846;
  assign n7848 = ~n4462 & n7847;
  assign n7849 = ~n5444 & n7847;
  assign n7850 = ~n7848 & ~n7849;
  assign n7851 = ~n7842 & n7847;
  assign n7852 = n1021 & ~n9513;
  assign n7853 = ~n1021 & n9513;
  assign n7854 = ~n7852 & ~n7853;
  assign n7855 = ~n1021 & n9233;
  assign n7856 = ~n9504 & ~n7855;
  assign n7857 = n9504 & n7855;
  assign n7858 = ~n9504 & n7855;
  assign n7859 = n9504 & ~n7855;
  assign n7860 = ~n7858 & ~n7859;
  assign n7861 = ~n7856 & ~n7857;
  assign n7862 = n7854 & ~n9514;
  assign n7863 = ~n7854 & n9514;
  assign n7864 = ~n7862 & ~n7863;
  assign n7865 = ~n7749 & ~n7770;
  assign n7866 = ~n7769 & ~n7776;
  assign n7867 = n7749 & ~n7769;
  assign n7868 = ~n7770 & ~n7867;
  assign n7869 = ~n7769 & ~n7865;
  assign n7870 = n7864 & ~n9515;
  assign n7871 = ~n7864 & n9515;
  assign n7872 = ~n9515 & ~n7870;
  assign n7873 = n7864 & ~n7870;
  assign n7874 = ~n7872 & ~n7873;
  assign n7875 = ~n7870 & ~n7871;
  assign n7876 = n7841 & ~n9516;
  assign n7877 = ~n7841 & ~n7873;
  assign n7878 = ~n7872 & n7877;
  assign n7879 = ~n7841 & n9516;
  assign n7880 = ~n7876 & ~n9517;
  assign n7881 = ~n7832 & n7880;
  assign n7882 = n7832 & ~n7880;
  assign n7883 = ~n7881 & ~n7882;
  assign n7884 = ~n7831 & n7883;
  assign n7885 = n7831 & ~n7883;
  assign n7886 = ~n7884 & ~n7885;
  assign n7887 = ~n223 & n712;
  assign n7888 = n655 & n7887;
  assign n7889 = n8708 & n7888;
  assign n7890 = n8721 & n7889;
  assign n7891 = n9281 & n7890;
  assign n7892 = n655 & n712;
  assign n7893 = n8721 & n7892;
  assign n7894 = n9281 & n7893;
  assign n7895 = n8775 & n7894;
  assign n7896 = n8708 & n7895;
  assign n7897 = ~n223 & n7896;
  assign n7898 = n8775 & n7891;
  assign n7899 = ~n7886 & n9518;
  assign n7900 = n7886 & ~n9518;
  assign n7901 = ~n7899 & ~n7900;
  assign n7902 = ~n7830 & n7901;
  assign n7903 = n7830 & ~n7901;
  assign n7904 = ~n7902 & ~n7903;
  assign n7905 = ~n7823 & ~n7904;
  assign n7906 = n7823 & n7904;
  assign n7907 = ~n7905 & ~n7906;
  assign n7908 = ~n7824 & n7825;
  assign n7909 = ~n9332 & ~n7908;
  assign n7910 = n7907 & ~n7909;
  assign n7911 = ~n7907 & n7909;
  assign n7912 = ~n7910 & ~n7911;
  assign n7913 = ~n7900 & ~n7902;
  assign n7914 = ~n7881 & ~n7884;
  assign n7915 = ~n7870 & ~n7876;
  assign n7916 = ~n7856 & ~n7862;
  assign n7917 = ~n1021 & ~n5405;
  assign n7918 = ~n7855 & n7917;
  assign n7919 = ~n9233 & n7917;
  assign n7920 = n7855 & ~n7917;
  assign n7921 = n5405 & n7855;
  assign n7922 = ~n9519 & ~n9520;
  assign n7923 = ~n7916 & ~n9520;
  assign n7924 = ~n9519 & n7923;
  assign n7925 = ~n7916 & n7922;
  assign n7926 = n7916 & ~n7922;
  assign n7927 = ~n7916 & ~n9521;
  assign n7928 = ~n9520 & ~n9521;
  assign n7929 = ~n9519 & n7928;
  assign n7930 = ~n7927 & ~n7929;
  assign n7931 = ~n9521 & ~n7926;
  assign n7932 = n4462 & n5882;
  assign n7933 = n4472 & n5875;
  assign n7934 = n4472 & ~n9283;
  assign n7935 = n4470 & ~n5437;
  assign n7936 = n9151 & n9246;
  assign n7937 = ~n7935 & ~n7936;
  assign n7938 = ~n9523 & n7937;
  assign n7939 = ~n7932 & n7938;
  assign n7940 = ~n1021 & ~n7939;
  assign n7941 = ~n1021 & ~n7940;
  assign n7942 = ~n1021 & n7939;
  assign n7943 = ~n7939 & ~n7940;
  assign n7944 = n1021 & ~n7939;
  assign n7945 = ~n9524 & ~n9525;
  assign n7946 = n4417 & ~n9365;
  assign n7947 = ~n9134 & ~n7946;
  assign n7948 = n9134 & ~n9337;
  assign n7949 = n4417 & n6524;
  assign n7950 = ~n7948 & ~n7949;
  assign n7951 = ~n9337 & ~n7947;
  assign n7952 = n8725 & ~n9526;
  assign n7953 = ~n8725 & n9526;
  assign n7954 = ~n8725 & ~n9526;
  assign n7955 = n8725 & n9526;
  assign n7956 = ~n7954 & ~n7955;
  assign n7957 = ~n7952 & ~n7953;
  assign n7958 = ~n7945 & n9527;
  assign n7959 = n7945 & ~n9527;
  assign n7960 = n9527 & ~n7958;
  assign n7961 = ~n7945 & ~n7958;
  assign n7962 = ~n7960 & ~n7961;
  assign n7963 = ~n7958 & ~n7959;
  assign n7964 = ~n9522 & ~n9528;
  assign n7965 = n9522 & n9528;
  assign n7966 = n9522 & ~n9528;
  assign n7967 = ~n9522 & n9528;
  assign n7968 = ~n7966 & ~n7967;
  assign n7969 = ~n7964 & ~n7965;
  assign n7970 = ~n7915 & ~n9529;
  assign n7971 = n7915 & n9529;
  assign n7972 = ~n7970 & ~n7971;
  assign n7973 = ~n7914 & n7972;
  assign n7974 = n7914 & ~n7972;
  assign n7975 = ~n7973 & ~n7974;
  assign n7976 = ~n271 & ~n820;
  assign n7977 = ~n177 & ~n392;
  assign n7978 = ~n642 & n7977;
  assign n7979 = ~n271 & n7977;
  assign n7980 = ~n642 & n7979;
  assign n7981 = ~n820 & n7980;
  assign n7982 = ~n271 & ~n642;
  assign n7983 = ~n820 & n7982;
  assign n7984 = n7977 & n7983;
  assign n7985 = n7976 & n7978;
  assign n7986 = ~n236 & ~n391;
  assign n7987 = n3691 & n7986;
  assign n7988 = n791 & n7987;
  assign n7989 = n9390 & n7988;
  assign n7990 = n9530 & n7989;
  assign n7991 = n9058 & n7990;
  assign n7992 = n3691 & n9530;
  assign n7993 = n791 & n7992;
  assign n7994 = n9390 & n7993;
  assign n7995 = n9022 & n7994;
  assign n7996 = n9058 & n7995;
  assign n7997 = ~n8643 & n7996;
  assign n7998 = ~n8637 & n7997;
  assign n7999 = ~n391 & n7998;
  assign n8000 = n9022 & n7990;
  assign n8001 = n9058 & n8000;
  assign n8002 = n9022 & n7991;
  assign n8003 = ~n7975 & n9531;
  assign n8004 = n7975 & ~n9531;
  assign n8005 = ~n8003 & ~n8004;
  assign n8006 = ~n7913 & n8005;
  assign n8007 = n7913 & ~n8005;
  assign n8008 = ~n8006 & ~n8007;
  assign n8009 = ~n7906 & ~n8008;
  assign n8010 = n7906 & n8008;
  assign n8011 = ~n8009 & ~n8010;
  assign n8012 = ~n7907 & n7908;
  assign n8013 = ~n9332 & ~n8012;
  assign n8014 = n8011 & ~n8013;
  assign n8015 = ~n8011 & n8013;
  assign n8016 = ~n8014 & ~n8015;
  assign n8017 = ~n8004 & ~n8006;
  assign n8018 = ~n7970 & ~n7973;
  assign n8019 = ~n7958 & ~n7964;
  assign n8020 = n4462 & n6341;
  assign n8021 = n4472 & ~n9337;
  assign n8022 = n4470 & n5875;
  assign n8023 = n4470 & ~n9283;
  assign n8024 = n9151 & ~n5437;
  assign n8025 = ~n9532 & ~n8024;
  assign n8026 = ~n8021 & n8025;
  assign n8027 = ~n8020 & n8026;
  assign n8028 = ~n1021 & ~n8027;
  assign n8029 = ~n8027 & ~n8028;
  assign n8030 = n1021 & ~n8027;
  assign n8031 = ~n1021 & ~n8028;
  assign n8032 = ~n1021 & n8027;
  assign n8033 = ~n9533 & ~n9534;
  assign n8034 = n8725 & n7917;
  assign n8035 = ~n8725 & ~n7917;
  assign n8036 = ~n8034 & ~n8035;
  assign n8037 = ~n1021 & n9246;
  assign n8038 = n8036 & n8037;
  assign n8039 = ~n8036 & ~n8037;
  assign n8040 = ~n8038 & ~n8039;
  assign n8041 = ~n8033 & n8040;
  assign n8042 = n8033 & ~n8040;
  assign n8043 = ~n8033 & ~n8041;
  assign n8044 = ~n8033 & ~n8040;
  assign n8045 = n8040 & ~n8041;
  assign n8046 = n8033 & n8040;
  assign n8047 = ~n9535 & ~n9536;
  assign n8048 = ~n8041 & ~n8042;
  assign n8049 = ~n7928 & ~n9537;
  assign n8050 = n7928 & n9537;
  assign n8051 = ~n7928 & n9537;
  assign n8052 = n7928 & ~n9537;
  assign n8053 = ~n8051 & ~n8052;
  assign n8054 = ~n8049 & ~n8050;
  assign n8055 = ~n8019 & ~n9538;
  assign n8056 = n8019 & n9538;
  assign n8057 = ~n8055 & ~n8056;
  assign n8058 = ~n8018 & n8057;
  assign n8059 = n8018 & ~n8057;
  assign n8060 = ~n8058 & ~n8059;
  assign n8061 = ~n251 & ~n8678;
  assign n8062 = ~n331 & ~n821;
  assign n8063 = ~n339 & n8062;
  assign n8064 = ~n331 & ~n339;
  assign n8065 = ~n251 & n8064;
  assign n8066 = ~n8678 & n8065;
  assign n8067 = ~n821 & n8066;
  assign n8068 = ~n339 & ~n821;
  assign n8069 = ~n331 & ~n8678;
  assign n8070 = ~n251 & n8069;
  assign n8071 = n8068 & n8070;
  assign n8072 = n8061 & n8063;
  assign n8073 = ~n222 & ~n8709;
  assign n8074 = n1119 & n8073;
  assign n8075 = n567 & n1728;
  assign n8076 = n8074 & n8075;
  assign n8077 = ~n412 & ~n486;
  assign n8078 = ~n386 & n8077;
  assign n8079 = n9361 & n8078;
  assign n8080 = n1119 & n8077;
  assign n8081 = n8075 & n8080;
  assign n8082 = ~n222 & ~n386;
  assign n8083 = ~n8709 & n8082;
  assign n8084 = n9361 & n8083;
  assign n8085 = n8081 & n8084;
  assign n8086 = n8076 & n8079;
  assign n8087 = n9539 & n9540;
  assign n8088 = n8816 & n8087;
  assign n8089 = n9102 & n9310;
  assign n8090 = n1119 & n9539;
  assign n8091 = n9361 & n8090;
  assign n8092 = n8816 & n8091;
  assign n8093 = n9102 & n8092;
  assign n8094 = n567 & n8093;
  assign n8095 = n9310 & n8094;
  assign n8096 = ~n341 & n8095;
  assign n8097 = ~n8709 & n8096;
  assign n8098 = ~n222 & n8097;
  assign n8099 = ~n636 & n8098;
  assign n8100 = ~n386 & n8099;
  assign n8101 = ~n486 & n8100;
  assign n8102 = ~n412 & n8101;
  assign n8103 = n8088 & n8089;
  assign n8104 = n8060 & ~n9541;
  assign n8105 = ~n8060 & n9541;
  assign n8106 = ~n8104 & ~n8105;
  assign n8107 = ~n8017 & ~n8105;
  assign n8108 = ~n8104 & n8107;
  assign n8109 = ~n8017 & n8106;
  assign n8110 = n8017 & ~n8106;
  assign n8111 = ~n8017 & ~n9542;
  assign n8112 = ~n8104 & ~n9542;
  assign n8113 = ~n8105 & n8112;
  assign n8114 = ~n8111 & ~n8113;
  assign n8115 = ~n9542 & ~n8110;
  assign n8116 = ~n8010 & n9543;
  assign n8117 = n8010 & ~n9543;
  assign n8118 = ~n8116 & ~n8117;
  assign n8119 = ~n8011 & n8012;
  assign n8120 = ~n9332 & ~n8119;
  assign n8121 = n8118 & ~n8120;
  assign n8122 = ~n8118 & n8120;
  assign n8123 = ~n8121 & ~n8122;
  assign n8124 = ~n8055 & ~n8058;
  assign n8125 = ~n8041 & ~n8049;
  assign n8126 = n4462 & n9366;
  assign n8127 = n9151 & n5875;
  assign n8128 = n9151 & ~n9283;
  assign n8129 = n4470 & ~n9337;
  assign n8130 = ~n9544 & ~n8129;
  assign n8131 = ~n4462 & n8130;
  assign n8132 = ~n9366 & n8130;
  assign n8133 = ~n8131 & ~n8132;
  assign n8134 = ~n8126 & n8130;
  assign n8135 = n1021 & ~n9545;
  assign n8136 = ~n1021 & n9545;
  assign n8137 = ~n8135 & ~n8136;
  assign n8138 = ~n1021 & ~n5437;
  assign n8139 = ~n8034 & ~n8038;
  assign n8140 = ~n8138 & ~n8139;
  assign n8141 = n8138 & n8139;
  assign n8142 = ~n8138 & ~n8140;
  assign n8143 = ~n8138 & n8139;
  assign n8144 = ~n8139 & ~n8140;
  assign n8145 = n8138 & ~n8139;
  assign n8146 = ~n9546 & ~n9547;
  assign n8147 = ~n8140 & ~n8141;
  assign n8148 = n8137 & ~n9548;
  assign n8149 = ~n8137 & n9548;
  assign n8150 = ~n8148 & ~n8149;
  assign n8151 = ~n8125 & n8150;
  assign n8152 = n8125 & ~n8150;
  assign n8153 = ~n8151 & ~n8152;
  assign n8154 = ~n8124 & n8153;
  assign n8155 = n8124 & ~n8153;
  assign n8156 = ~n8154 & ~n8155;
  assign n8157 = n1200 & n3691;
  assign n8158 = n3847 & n5378;
  assign n8159 = n8157 & n8158;
  assign n8160 = ~n212 & ~n256;
  assign n8161 = ~n417 & n8160;
  assign n8162 = ~n223 & ~n8709;
  assign n8163 = n903 & n8162;
  assign n8164 = n8161 & n8163;
  assign n8165 = n903 & n3691;
  assign n8166 = n8158 & n8165;
  assign n8167 = ~n223 & ~n256;
  assign n8168 = ~n8709 & n8167;
  assign n8169 = ~n212 & ~n417;
  assign n8170 = n1200 & n8169;
  assign n8171 = n8168 & n8170;
  assign n8172 = n8166 & n8171;
  assign n8173 = n8159 & n8164;
  assign n8174 = n8670 & n9549;
  assign n8175 = n8680 & n8892;
  assign n8176 = n8174 & n8175;
  assign n8177 = n3691 & n3847;
  assign n8178 = n903 & n8177;
  assign n8179 = n8680 & n8178;
  assign n8180 = n9087 & n8179;
  assign n8181 = n8892 & n8180;
  assign n8182 = n8670 & n8181;
  assign n8183 = n5378 & n8182;
  assign n8184 = ~n212 & n8183;
  assign n8185 = ~n256 & n8184;
  assign n8186 = ~n166 & n8185;
  assign n8187 = ~n8709 & n8186;
  assign n8188 = ~n545 & n8187;
  assign n8189 = ~n223 & n8188;
  assign n8190 = ~n417 & n8189;
  assign n8191 = n9087 & n8176;
  assign n8192 = ~n8156 & n9550;
  assign n8193 = n8156 & ~n9550;
  assign n8194 = ~n8192 & ~n8193;
  assign n8195 = ~n8112 & n8194;
  assign n8196 = n8112 & ~n8194;
  assign n8197 = ~n8195 & ~n8196;
  assign n8198 = ~n8117 & ~n8197;
  assign n8199 = n8117 & n8197;
  assign n8200 = ~n8198 & ~n8199;
  assign n8201 = ~n8118 & n8119;
  assign n8202 = ~n9332 & ~n8201;
  assign n8203 = n8200 & ~n8202;
  assign n8204 = ~n8200 & n8202;
  assign n8205 = ~n8203 & ~n8204;
  assign n8206 = ~n8193 & ~n8195;
  assign n8207 = ~n8140 & ~n8148;
  assign n8208 = n4462 & ~n9365;
  assign n8209 = ~n9151 & ~n8208;
  assign n8210 = n9151 & ~n9337;
  assign n8211 = n4462 & n6524;
  assign n8212 = ~n8210 & ~n8211;
  assign n8213 = ~n9337 & ~n8209;
  assign n8214 = ~n1021 & ~n9551;
  assign n8215 = n5879 & n8214;
  assign n8216 = ~n1021 & ~n5879;
  assign n8217 = n9551 & ~n8216;
  assign n8218 = ~n9551 & ~n8214;
  assign n8219 = n1021 & ~n9551;
  assign n8220 = ~n1021 & ~n8214;
  assign n8221 = ~n1021 & n9551;
  assign n8222 = ~n9552 & ~n9553;
  assign n8223 = ~n1021 & n5879;
  assign n8224 = ~n8222 & ~n8223;
  assign n8225 = ~n8214 & ~n8217;
  assign n8226 = ~n8223 & ~n9554;
  assign n8227 = n8222 & ~n8223;
  assign n8228 = ~n8222 & ~n9554;
  assign n8229 = n5879 & n9553;
  assign n8230 = ~n9555 & ~n9556;
  assign n8231 = ~n8215 & ~n9554;
  assign n8232 = n8207 & n9557;
  assign n8233 = ~n8207 & ~n9557;
  assign n8234 = ~n8232 & ~n8233;
  assign n8235 = ~n8151 & ~n8154;
  assign n8236 = ~n8234 & n8235;
  assign n8237 = n8234 & ~n8235;
  assign n8238 = ~n8236 & ~n8237;
  assign n8239 = ~n295 & ~n474;
  assign n8240 = ~n342 & n8239;
  assign n8241 = ~n474 & n3846;
  assign n8242 = ~n295 & n8820;
  assign n8243 = ~n342 & n8242;
  assign n8244 = ~n474 & n8243;
  assign n8245 = n8820 & n9558;
  assign n8246 = ~n8648 & ~n445;
  assign n8247 = ~n166 & ~n608;
  assign n8248 = ~n166 & ~n445;
  assign n8249 = ~n8648 & ~n608;
  assign n8250 = n8248 & n8249;
  assign n8251 = n8246 & n8247;
  assign n8252 = n657 & n1344;
  assign n8253 = n6192 & n8252;
  assign n8254 = n9560 & n8253;
  assign n8255 = n9530 & n8254;
  assign n8256 = n8817 & n8255;
  assign n8257 = n9061 & n8256;
  assign n8258 = n657 & n9559;
  assign n8259 = n1344 & n8258;
  assign n8260 = n9530 & n8259;
  assign n8261 = n9061 & n8260;
  assign n8262 = n8817 & n8261;
  assign n8263 = ~n166 & n8262;
  assign n8264 = ~n8648 & n8263;
  assign n8265 = ~n445 & n8264;
  assign n8266 = ~n608 & n8265;
  assign n8267 = ~n417 & n8266;
  assign n8268 = ~n448 & n8267;
  assign n8269 = n9559 & n8257;
  assign n8270 = n8238 & ~n9561;
  assign n8271 = ~n8238 & n9561;
  assign n8272 = ~n8270 & ~n8271;
  assign n8273 = ~n8206 & ~n8271;
  assign n8274 = ~n8270 & n8273;
  assign n8275 = ~n8206 & n8272;
  assign n8276 = n8206 & ~n8272;
  assign n8277 = ~n8206 & ~n9562;
  assign n8278 = ~n8270 & ~n9562;
  assign n8279 = ~n8271 & n8278;
  assign n8280 = ~n8277 & ~n8279;
  assign n8281 = ~n9562 & ~n8276;
  assign n8282 = ~n8199 & n9563;
  assign n8283 = n8199 & ~n9563;
  assign n8284 = ~n8282 & ~n8283;
  assign n8285 = ~n8200 & n8201;
  assign n8286 = ~n9332 & ~n8285;
  assign n8287 = n8284 & ~n8286;
  assign n8288 = ~n8284 & n8286;
  assign n8289 = ~n8287 & ~n8288;
  assign n8290 = ~n8640 & ~n904;
  assign n8291 = ~n8664 & ~n904;
  assign n8292 = ~n8640 & n8291;
  assign n8293 = ~n8664 & n8290;
  assign n8294 = n446 & n762;
  assign n8295 = n9564 & n8294;
  assign n8296 = n9028 & n8295;
  assign n8297 = n9301 & n9539;
  assign n8298 = n8296 & n8297;
  assign n8299 = n9311 & n8298;
  assign n8300 = n762 & n9041;
  assign n8301 = n9028 & n8300;
  assign n8302 = n9539 & n8301;
  assign n8303 = n9301 & n8302;
  assign n8304 = n446 & n8303;
  assign n8305 = n9311 & n8304;
  assign n8306 = ~n8640 & n8305;
  assign n8307 = ~n8664 & n8306;
  assign n8308 = ~n904 & n8307;
  assign n8309 = n9041 & n8299;
  assign n8310 = ~n1021 & ~n9283;
  assign n8311 = ~n9283 & ~n8138;
  assign n8312 = ~n1021 & n8311;
  assign n8313 = ~n8138 & n8310;
  assign n8314 = n5437 & n8310;
  assign n8315 = ~n9554 & ~n9566;
  assign n8316 = ~n8233 & ~n8237;
  assign n8317 = ~n5437 & n9337;
  assign n8318 = n5437 & ~n9337;
  assign n8319 = ~n1021 & ~n8318;
  assign n8320 = n9337 & n8138;
  assign n8321 = ~n9337 & ~n8138;
  assign n8322 = ~n8320 & ~n8321;
  assign n8323 = ~n1021 & n8322;
  assign n8324 = n8319 & ~n8320;
  assign n8325 = ~n8317 & n8319;
  assign n8326 = n8316 & ~n9567;
  assign n8327 = ~n8316 & n9567;
  assign n8328 = ~n8326 & ~n8327;
  assign n8329 = n8315 & n8328;
  assign n8330 = ~n8315 & ~n8328;
  assign n8331 = n8315 & ~n8316;
  assign n8332 = ~n8315 & n8316;
  assign n8333 = ~n8331 & ~n8332;
  assign n8334 = ~n9567 & n8333;
  assign n8335 = n9567 & ~n8333;
  assign n8336 = ~n8334 & ~n8335;
  assign n8337 = ~n8329 & ~n8330;
  assign n8338 = n9565 & n9568;
  assign n8339 = ~n9565 & ~n9568;
  assign n8340 = ~n8338 & ~n8339;
  assign n8341 = n8278 & ~n8340;
  assign n8342 = ~n8278 & ~n8338;
  assign n8343 = ~n8339 & n8342;
  assign n8344 = ~n8278 & n8340;
  assign n8345 = n8278 & ~n8339;
  assign n8346 = ~n8339 & ~n9569;
  assign n8347 = ~n8338 & ~n8345;
  assign n8348 = ~n8338 & n9570;
  assign n8349 = n8278 & n8340;
  assign n8350 = ~n8278 & ~n9569;
  assign n8351 = ~n8278 & ~n8340;
  assign n8352 = ~n9571 & ~n9572;
  assign n8353 = ~n8341 & ~n9569;
  assign n8354 = ~n8283 & n9573;
  assign n8355 = n8283 & ~n9573;
  assign n8356 = ~n8354 & ~n8355;
  assign n8357 = ~n8284 & n8285;
  assign n8358 = ~n9332 & ~n8357;
  assign n8359 = n8356 & ~n8358;
  assign n8360 = ~n8356 & n8358;
  assign n8361 = ~n8359 & ~n8360;
  assign n8362 = ~n8356 & n8357;
  assign n8363 = ~n9332 & ~n8362;
  assign n8364 = ~n271 & ~n430;
  assign n8365 = n4166 & n8364;
  assign n8366 = n567 & n701;
  assign n8367 = n8365 & n8366;
  assign n8368 = ~n393 & ~n493;
  assign n8369 = ~n8643 & n8368;
  assign n8370 = n8660 & n8369;
  assign n8371 = ~n8643 & ~n430;
  assign n8372 = n701 & n8371;
  assign n8373 = n567 & n4166;
  assign n8374 = n8372 & n8373;
  assign n8375 = ~n271 & n8368;
  assign n8376 = n8660 & n8375;
  assign n8377 = n8374 & n8376;
  assign n8378 = n8367 & n8370;
  assign n8379 = n8742 & n9574;
  assign n8380 = n8741 & n8379;
  assign n8381 = n8660 & n8742;
  assign n8382 = n701 & n8381;
  assign n8383 = n4166 & n8382;
  assign n8384 = n9229 & n8383;
  assign n8385 = n8741 & n8384;
  assign n8386 = n567 & n8385;
  assign n8387 = ~n8643 & n8386;
  assign n8388 = ~n271 & n8387;
  assign n8389 = ~n430 & n8388;
  assign n8390 = ~n493 & n8389;
  assign n8391 = ~n393 & n8390;
  assign n8392 = n9229 & n8380;
  assign n8393 = ~n9570 & ~n9575;
  assign n8394 = n9570 & n9575;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = n8355 & n8395;
  assign n8397 = ~n8355 & ~n8395;
  assign n8398 = ~n8396 & ~n8397;
  assign n8399 = ~n8355 & n8395;
  assign n8400 = n8355 & ~n8395;
  assign n8401 = ~n8399 & ~n8400;
  assign n8402 = n8363 & ~n8401;
  assign n8403 = n8363 & n8398;
  assign n8404 = ~n8363 & n8401;
  assign n8405 = ~n8363 & ~n8398;
  assign po17  = ~n9576 & ~n9577;
  assign n8407 = n8362 & ~n8398;
  assign n8408 = ~n9332 & ~n8407;
  assign n8409 = ~n271 & ~n641;
  assign n8410 = ~n256 & ~n8645;
  assign n8411 = ~n434 & n8410;
  assign n8412 = ~n256 & ~n434;
  assign n8413 = ~n8645 & ~n641;
  assign n8414 = ~n271 & n8413;
  assign n8415 = n8412 & n8414;
  assign n8416 = n8409 & n8411;
  assign n8417 = n8668 & n8773;
  assign n8418 = n9578 & n8417;
  assign n8419 = n8813 & n9100;
  assign n8420 = n8418 & n8419;
  assign n8421 = n8821 & n8420;
  assign n8422 = n8745 & n9316;
  assign n8423 = n8745 & n9100;
  assign n8424 = n8773 & n8423;
  assign n8425 = n8821 & n8424;
  assign n8426 = n8813 & n8425;
  assign n8427 = n8668 & n8426;
  assign n8428 = n9316 & n8427;
  assign n8429 = ~n256 & n8428;
  assign n8430 = ~n8645 & n8429;
  assign n8431 = ~n271 & n8430;
  assign n8432 = ~n641 & n8431;
  assign n8433 = ~n434 & n8432;
  assign n8434 = n9316 & n8421;
  assign n8435 = n8745 & n8434;
  assign n8436 = n8421 & n8422;
  assign n8437 = n8393 & ~n9579;
  assign n8438 = ~n8393 & n9579;
  assign n8439 = ~n8437 & ~n8438;
  assign n8440 = ~n8396 & ~n8439;
  assign n8441 = n8396 & ~n8438;
  assign n8442 = ~n8393 & ~n8396;
  assign n8443 = n9579 & ~n8442;
  assign n8444 = ~n9579 & n8442;
  assign n8445 = ~n8443 & ~n8444;
  assign n8446 = ~n8440 & ~n8441;
  assign n8447 = n8362 & n8401;
  assign n8448 = ~n9332 & ~n8447;
  assign n8449 = n9580 & n8448;
  assign n8450 = n8408 & n9580;
  assign n8451 = ~n9580 & ~n8448;
  assign n8452 = ~n8408 & ~n9580;
  assign n8453 = ~n9581 & ~n9582;
  assign n8454 = ~n287 & ~n382;
  assign n8455 = n1333 & n8454;
  assign n8456 = n5196 & n8455;
  assign n8457 = ~n8630 & ~n244;
  assign n8458 = ~n658 & n8457;
  assign n8459 = n9441 & n8458;
  assign n8460 = n5196 & n8457;
  assign n8461 = n1333 & n8460;
  assign n8462 = ~n658 & n8454;
  assign n8463 = n9441 & n8462;
  assign n8464 = n8461 & n8463;
  assign n8465 = n8456 & n8459;
  assign n8466 = n9126 & n9583;
  assign n8467 = n8696 & n8466;
  assign n8468 = n9441 & n9559;
  assign n8469 = n1333 & n8468;
  assign n8470 = n9126 & n8469;
  assign n8471 = n8696 & n8470;
  assign n8472 = ~n244 & n8471;
  assign n8473 = ~n8630 & n8472;
  assign n8474 = ~n8640 & n8473;
  assign n8475 = ~n287 & n8474;
  assign n8476 = ~n658 & n8475;
  assign n8477 = ~n382 & n8476;
  assign n8478 = ~n431 & n8477;
  assign n8479 = n9559 & n8467;
  assign n8480 = ~n8437 & n9584;
  assign n8481 = n8437 & ~n9584;
  assign n8482 = ~n8480 & ~n8481;
  assign n8483 = n8396 & ~n9579;
  assign n8484 = ~n8482 & ~n8483;
  assign n8485 = n8482 & n8483;
  assign n8486 = ~n8484 & ~n8485;
  assign n8487 = n8407 & n9580;
  assign n8488 = ~n9332 & ~n8487;
  assign n8489 = ~n8441 & ~n8482;
  assign n8490 = n8441 & n8482;
  assign n8491 = ~n8489 & ~n8490;
  assign n8492 = n9580 & n8447;
  assign n8493 = ~n9332 & ~n8492;
  assign n8494 = n8491 & ~n8493;
  assign n8495 = n8486 & ~n8488;
  assign n8496 = ~n8491 & n8493;
  assign n8497 = ~n8486 & n8488;
  assign n8498 = ~n9585 & ~n9586;
  assign n8499 = ~n8486 & n8487;
  assign n8500 = ~n9332 & ~n8499;
  assign n8501 = n866 & n6057;
  assign n8502 = n7420 & n8501;
  assign n8503 = n312 & ~n1073;
  assign n8504 = n7127 & n8503;
  assign n8505 = n8502 & n8504;
  assign n8506 = n8722 & n8505;
  assign n8507 = n8673 & n8506;
  assign n8508 = n178 & n866;
  assign n8509 = n8673 & n8508;
  assign n8510 = n8722 & n8509;
  assign n8511 = n9484 & n8510;
  assign n8512 = n3521 & n8511;
  assign n8513 = ~n331 & n8512;
  assign n8514 = ~n8645 & n8513;
  assign n8515 = ~n309 & n8514;
  assign n8516 = ~n198 & n8515;
  assign n8517 = ~n861 & n8516;
  assign n8518 = ~n377 & n8517;
  assign n8519 = ~n1073 & n8518;
  assign n8520 = n9484 & n8507;
  assign n8521 = n8481 & ~n9587;
  assign n8522 = ~n8481 & n9587;
  assign n8523 = ~n8521 & ~n8522;
  assign n8524 = ~n8490 & ~n8523;
  assign n8525 = n8490 & ~n8522;
  assign n8526 = ~n8481 & ~n8485;
  assign n8527 = n9587 & ~n8526;
  assign n8528 = ~n9587 & n8526;
  assign n8529 = ~n8527 & ~n8528;
  assign n8530 = ~n8524 & ~n8525;
  assign n8531 = ~n8491 & n8492;
  assign n8532 = ~n9332 & ~n8531;
  assign n8533 = n9588 & n8532;
  assign n8534 = n8500 & n9588;
  assign n8535 = ~n9588 & ~n8532;
  assign n8536 = ~n8500 & ~n9588;
  assign n8537 = ~n9589 & ~n9590;
  assign n8538 = ~n633 & n8714;
  assign n8539 = n9249 & n8538;
  assign n8540 = n8714 & n9249;
  assign n8541 = n8650 & n8540;
  assign n8542 = ~n8709 & n8541;
  assign n8543 = ~n8678 & n8542;
  assign n8544 = n8650 & n8539;
  assign n8545 = ~n8521 & n9591;
  assign n8546 = n8521 & ~n9591;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = n8485 & ~n9587;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = n8547 & n8548;
  assign n8551 = ~n8549 & ~n8550;
  assign n8552 = n8499 & n9588;
  assign n8553 = ~n9332 & ~n8552;
  assign n8554 = ~n8525 & ~n8547;
  assign n8555 = n8525 & n8547;
  assign n8556 = ~n8554 & ~n8555;
  assign n8557 = n9588 & n8531;
  assign n8558 = ~n9332 & ~n8557;
  assign n8559 = n8556 & ~n8558;
  assign n8560 = n8551 & ~n8553;
  assign n8561 = ~n8556 & n8558;
  assign n8562 = ~n8551 & n8553;
  assign n8563 = ~n9592 & ~n9593;
  assign n8564 = ~n8551 & n8552;
  assign n8565 = ~n9332 & ~n8564;
  assign n8566 = n8650 & n8719;
  assign n8567 = ~n8546 & ~n8550;
  assign n8568 = ~n8566 & ~n8567;
  assign n8569 = n8566 & n8567;
  assign n8570 = ~n8568 & ~n8569;
  assign n8571 = n8546 & ~n8566;
  assign n8572 = ~n8546 & n8566;
  assign n8573 = ~n8571 & ~n8572;
  assign n8574 = ~n8555 & ~n8573;
  assign n8575 = n8555 & ~n8572;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = ~n8556 & n8557;
  assign n8578 = ~n9332 & ~n8577;
  assign n8579 = n8576 & ~n8578;
  assign n8580 = n8566 & ~n8567;
  assign n8581 = ~n8566 & n8567;
  assign n8582 = ~n8580 & ~n8581;
  assign n8583 = ~n8565 & ~n8582;
  assign n8584 = ~n8565 & n8570;
  assign n8585 = ~n8576 & n8578;
  assign n8586 = n8565 & n8582;
  assign n8587 = n8565 & ~n8570;
  assign n8588 = ~n9594 & ~n9595;
  assign n8589 = n8564 & ~n8570;
  assign n8590 = ~n9332 & ~n8568;
  assign n8591 = ~n8571 & ~n8575;
  assign n8592 = ~n8576 & n8577;
  assign n8593 = ~n9332 & ~n8592;
  assign n8594 = n8591 & n8593;
  assign n8595 = n8564 & n8582;
  assign n8596 = ~n9332 & ~n8595;
  assign n8597 = ~n8568 & n8596;
  assign n8598 = ~n8589 & n8590;
  assign n8599 = n117 & n124;
  assign n8600 = ~n8565 & n8568;
  assign n8601 = ~n8599 & ~n8600;
  assign n8602 = ~pi22  & n127;
  assign n8603 = ~n8591 & ~n8593;
  assign n8604 = ~n9596 & ~n8603;
  assign n8605 = ~n8602 & n8604;
  assign n8606 = n8568 & ~n8596;
  assign n8607 = ~n9596 & ~n8602;
  assign n8608 = ~n8606 & n8607;
  assign n8609 = ~n9596 & n8601;
  assign n8610 = n8564 & n8568;
  assign n8611 = ~n8602 & ~n8610;
  assign n8612 = ~n8599 & ~n8610;
  assign n8613 = ~n8591 & n8592;
  assign n8614 = n8592 & ~n8613;
  assign n8615 = ~n8602 & n8614;
  assign n8616 = n8595 & n9598;
  assign n8617 = n8589 & n9598;
  assign po24  = ~n9332 & ~n9599;
  assign n8619 = n52 | n53;
  assign n8620 = n61 | ~n62;
  assign n8621 = n71 | ~n72;
  assign n8622 = n78 | ~n79;
  assign n8623 = n88 | ~n89;
  assign n8624 = n109 | n110;
  assign n8625 = n120 | n121;
  assign n8626 = n131 | n132;
  assign n8627 = n133 | n134;
  assign n8628 = n154 | ~n155;
  assign n8629 = n173 | n174;
  assign n8630 = n181 | n182;
  assign n8631 = n183 | n184;
  assign n8632 = n195 | n191 | n194;
  assign n8633 = n201 | n202;
  assign n8634 = n219 | n216 | n218;
  assign n8635 = n226 | n227;
  assign n8636 = n234 | n235;
  assign n8637 = n237 | n238;
  assign n8638 = n248 | n249;
  assign n8639 = n268 | n269;
  assign n8640 = n275 | n276;
  assign n8641 = n284 | n285;
  assign n8642 = n289 | n290;
  assign n8643 = n293 | n294;
  assign n8644 = n307 | n308;
  assign n8645 = n310 | n311;
  assign n8646 = n318 | n319;
  assign n8647 = n320 | n321;
  assign n8648 = n322 | n323;
  assign n8649 = n328 | n329;
  assign n8650 = n349 | n350;
  assign n8651 = n356 | ~n357;
  assign n8652 = n365 | n366;
  assign n8653 = n375 | n372 | n374;
  assign n8654 = n396 | n397;
  assign n8655 = n410 | n411;
  assign n8656 = n429 | n425 | n428;
  assign n8657 = n440 | n441;
  assign n8658 = n457 | n454 | n456;
  assign n8659 = n467 | n468;
  assign n8660 = n472 | n473;
  assign n8661 = n478 | n479;
  assign n8662 = n506 | n502 | n505;
  assign n8663 = n508 | n509;
  assign n8664 = n515 | n516;
  assign n8665 = n528 | n523 | n527;
  assign n8666 = n540 | n541;
  assign n8667 = n549 | n550;
  assign n8668 = n559 | n555 | n558;
  assign n8669 = n565 | n566;
  assign n8670 = n572 | n573;
  assign n8671 = n579 | n580;
  assign n8672 = n590 | n591;
  assign n8673 = n598 | n599;
  assign n8674 = n600 | n601;
  assign n8675 = n606 | n607;
  assign n8676 = n624 | n621 | n623;
  assign n8677 = n628 | n629;
  assign n8678 = n634 | n635;
  assign n8679 = n639 | n640;
  assign n8680 = n652 | n653;
  assign n8681 = n667 | n668;
  assign n8682 = n678 | n679;
  assign n8683 = n682 | n683;
  assign n8684 = n690 | n691;
  assign n8685 = n695 | n696;
  assign n8686 = n697 | n698;
  assign n8687 = n711 | n707 | n710;
  assign n8688 = n716 | n717;
  assign n8689 = n730 | n731;
  assign n8690 = n734 | n735;
  assign n8691 = n744 | n745;
  assign n8692 = n751 | n752;
  assign n8693 = n756 | n757;
  assign n8694 = n760 | n761;
  assign n8695 = n768 | n769;
  assign n8696 = n778 | n779;
  assign n8697 = n785 | n782 | n784;
  assign n8698 = n788 | n789;
  assign n8699 = n794 | n795;
  assign n8700 = n796 | n797;
  assign n8701 = n801 | n802;
  assign n8702 = n807 | n808;
  assign n8703 = n813 | n814;
  assign n8704 = n828 | n829;
  assign n8705 = n843 | n844;
  assign n8706 = n857 | n858;
  assign n8707 = n872 | n873;
  assign n8708 = n879 | n880;
  assign n8709 = n881 | n882;
  assign n8710 = n893 | n890 | n892;
  assign n8711 = n901 | n902;
  assign n8712 = n908 | n909;
  assign n8713 = n920 | n921;
  assign n8714 = n927 | n928;
  assign n8715 = n936 | n937;
  assign n8716 = n941 | n942;
  assign n8717 = n952 | n953;
  assign n8718 = n959 | n960;
  assign n8719 = n965 | n966;
  assign n8720 = n970 | n971;
  assign n8721 = n974 | n975;
  assign n8722 = n980 | n981;
  assign n8723 = n984 | n985;
  assign n8724 = n990 | ~n991;
  assign n8725 = n1004 | ~n1005;
  assign n8726 = n1009 | n1010;
  assign n8727 = n1013 | n1014;
  assign n8728 = n1019 | n1020;
  assign n8729 = n1032 | n1028 | n1031;
  assign n8730 = n1041 | n1042;
  assign n8731 = n1046 | n1047;
  assign n8732 = n1054 | n1051 | n1053;
  assign n8733 = n1056 | n1057;
  assign n8734 = n1067 | n1063 | n1066;
  assign n8735 = n1070 | n1071;
  assign n8736 = n1078 | n1079;
  assign n8737 = n1085 | n1082 | n1084;
  assign n8738 = n1088 | n1089;
  assign n8739 = n1104 | n1100 | n1103;
  assign n8740 = n1105 | ~n1106;
  assign n8741 = n1117 | n1118;
  assign n8742 = n1126 | n1123 | n1125;
  assign n8743 = n1137 | n1138;
  assign n8744 = n1145 | n1146;
  assign n8745 = n1149 | n1150;
  assign n8746 = n1162 | n1159 | n1161;
  assign n8747 = n1168 | n1169;
  assign n8748 = n1175 | n1176;
  assign n8749 = n1185 | n1186;
  assign n8750 = n1189 | n1190;
  assign n8751 = n1198 | n1199;
  assign n8752 = n1202 | n1203;
  assign n8753 = n1211 | n1207 | n1210;
  assign n8754 = n1215 | n1216;
  assign n8755 = n1219 | n1220;
  assign n8756 = n1223 | n1224;
  assign n8757 = n1230 | n1231;
  assign n8758 = n1244 | n1240 | n1243;
  assign n8759 = n1246 | n1247;
  assign n8760 = n1257 | n1258;
  assign n8761 = n1269 | n1270;
  assign n8762 = n1273 | n1274;
  assign n8763 = n1285 | n1286;
  assign n8764 = n1291 | ~n1292;
  assign n8765 = n1294 | n1295;
  assign n8766 = n1298 | n1299;
  assign n8767 = n1307 | ~n1308;
  assign n8768 = n1312 | n1313;
  assign n8769 = n1321 | n1317 | n1320;
  assign n8770 = n1330 | n1331;
  assign n8771 = n1341 | n1342;
  assign n8772 = n1349 | n1350;
  assign n8773 = n1353 | n1354;
  assign n8774 = n1358 | n1359;
  assign n8775 = n1370 | n1371;
  assign n8776 = n1380 | n1381;
  assign n8777 = n1384 | n1385;
  assign n8778 = n1390 | n1391;
  assign n8779 = n1397 | n1398;
  assign n8780 = n1416 | n1417;
  assign n8781 = n1422 | ~n1423;
  assign n8782 = n1425 | n1426;
  assign n8783 = n1429 | n1430;
  assign n8784 = n1436 | n1437;
  assign n8785 = n1441 | n1442;
  assign n8786 = n1447 | ~n1448;
  assign n8787 = n1453 | ~n1454;
  assign n8788 = n1460 | n1461;
  assign n8789 = n1464 | n1465;
  assign n8790 = n1471 | ~n1472;
  assign n8791 = n1487 | ~n1488;
  assign n8792 = n1501 | n1502;
  assign n8793 = n1510 | n1511;
  assign n8794 = n1514 | n1515;
  assign n8795 = n1523 | n1524;
  assign n8796 = n1535 | ~n1536;
  assign n8797 = n1547 | n1548;
  assign n8798 = n1551 | n1552;
  assign n8799 = n1560 | n1561;
  assign n8800 = n1562 | n1563;
  assign n8801 = n1564 | ~n1565;
  assign n8802 = n1568 | n1569;
  assign n8803 = n1570 | n1571;
  assign n8804 = n1572 | ~n1573;
  assign n8805 = n1579 | n1580;
  assign n8806 = n1583 | n1584;
  assign n8807 = n1592 | n1593;
  assign n8808 = n1600 | n1601;
  assign n8809 = n1606 | n1607;
  assign n8810 = n1613 | n1610 | n1612;
  assign n8811 = n1617 | n1618;
  assign n8812 = n1626 | n1627;
  assign n8813 = n1640 | n1641;
  assign n8814 = n1646 | n1647;
  assign n8815 = n1657 | n1658;
  assign n8816 = n1680 | n1672 | n1679;
  assign n8817 = n1699 | n1692 | n1698;
  assign n8818 = n1712 | n1713;
  assign n8819 = n1727 | n1724 | n1726;
  assign n8820 = n1753 | n1744 | n1752;
  assign n8821 = n1772 | n1764 | n1771;
  assign n8822 = n1788 | n1789;
  assign n8823 = n1799 | n1800;
  assign n8824 = n1805 | n1806;
  assign n8825 = n1814 | n1815;
  assign n8826 = n1819 | n1820;
  assign n8827 = n1823 | n1824;
  assign n8828 = n1837 | n1838;
  assign n8829 = n1841 | n1842;
  assign n8830 = n1852 | n1849 | n1851;
  assign n8831 = n1856 | n1857;
  assign n8832 = n1863 | ~n1864;
  assign n8833 = n1866 | n1867;
  assign n8834 = n1869 | ~n1870;
  assign n8835 = n1873 | n1874;
  assign n8836 = n1890 | n1886 | n1889;
  assign n8837 = n1898 | ~n1899;
  assign n8838 = n1901 | n1902;
  assign n8839 = n1903 | n1904;
  assign n8840 = n1905 | ~n1906;
  assign n8841 = n1917 | ~n1918;
  assign n8842 = n1927 | ~n1928;
  assign n8843 = n1933 | n1934;
  assign n8844 = n1937 | n1938;
  assign n8845 = n1946 | n1947;
  assign n8846 = n1952 | ~n1953;
  assign n8847 = n1954 | n1955;
  assign n8848 = n1964 | n1965;
  assign n8849 = n1976 | ~n1977;
  assign n8850 = n1981 | n1982;
  assign n8851 = n1983 | n1984;
  assign n8852 = n1985 | ~n1986;
  assign n8853 = n1990 | n1991;
  assign n8854 = n1992 | n1993;
  assign n8855 = n1994 | ~n1995;
  assign n8856 = n1999 | ~n2000;
  assign n8857 = n2002 | ~n2003;
  assign n8858 = n2006 | n2007;
  assign n8859 = n2008 | n2009;
  assign n8860 = n2022 | n2018 | n2021;
  assign n8861 = n2030 | ~n2031;
  assign n8862 = n2033 | n2034;
  assign n8863 = n2036 | ~n2037;
  assign n8864 = n2040 | n2041;
  assign n8865 = n2044 | n2045;
  assign n8866 = n2058 | n2059;
  assign n8867 = n2071 | n2067 | n2070;
  assign n8868 = n2076 | ~n2077;
  assign n8869 = n2085 | n2086;
  assign n8870 = n2096 | n2097;
  assign n8871 = n2106 | n2107;
  assign n8872 = n2109 | n2110;
  assign n8873 = n2116 | n2117;
  assign n8874 = n2120 | n2121;
  assign n8875 = n2136 | n2132 | n2135;
  assign n8876 = n2144 | n2145;
  assign n8877 = n2150 | ~n2151;
  assign n8878 = n2159 | n2160;
  assign n8879 = n2173 | ~n2174;
  assign n8880 = n2176 | n2177;
  assign n8881 = n2178 | n2179;
  assign n8882 = n2180 | ~n2181;
  assign n8883 = n2191 | ~n2192;
  assign n8884 = n2194 | n2195;
  assign n8885 = n2196 | n2197;
  assign n8886 = n2198 | ~n2199;
  assign n8887 = n2207 | n2208;
  assign n8888 = n2230 | n2221 | n2229;
  assign n8889 = n2242 | n2243;
  assign n8890 = n2267 | n2259 | n2266;
  assign n8891 = n2272 | n2273;
  assign n8892 = n2283 | n2284;
  assign n8893 = n2297 | n2298;
  assign n8894 = n2300 | n2301;
  assign n8895 = n2304 | ~n2305;
  assign n8896 = n2316 | n2317;
  assign n8897 = n2324 | n2325;
  assign n8898 = n2328 | n2329;
  assign n8899 = n2344 | n2340 | n2343;
  assign n8900 = n2352 | n2353;
  assign n8901 = n2358 | ~n2359;
  assign n8902 = n2367 | n2368;
  assign n8903 = n2374 | n2375;
  assign n8904 = n2376 | n2377;
  assign n8905 = n2378 | ~n2379;
  assign n8906 = n2392 | n2393;
  assign n8907 = n2394 | n2395;
  assign n8908 = n2396 | ~n2397;
  assign n8909 = n2408 | n2409;
  assign n8910 = n2415 | n2416;
  assign n8911 = n2419 | n2420;
  assign n8912 = n2433 | n2429 | n2432;
  assign n8913 = n2441 | n2442;
  assign n8914 = n2447 | ~n2448;
  assign n8915 = n2456 | n2457;
  assign n8916 = n2467 | ~n2468;
  assign n8917 = n2473 | ~n2474;
  assign n8918 = n2476 | n2477;
  assign n8919 = n2478 | n2479;
  assign n8920 = n2480 | ~n2481;
  assign n8921 = n2492 | ~n2493;
  assign n8922 = n2507 | n2508;
  assign n8923 = n2511 | n2512;
  assign n8924 = n2520 | n2521;
  assign n8925 = n2529 | n2530;
  assign n8926 = n2534 | n2535;
  assign n8927 = n2536 | n2537;
  assign n8928 = n2538 | ~n2539;
  assign n8929 = n2543 | n2544;
  assign n8930 = n2562 | n2563;
  assign n8931 = n2575 | n2571 | n2574;
  assign n8932 = n2582 | n2583;
  assign n8933 = n2593 | n2594;
  assign n8934 = n2599 | ~n2600;
  assign n8935 = n2612 | n2613;
  assign n8936 = n2621 | n2622;
  assign n8937 = n2627 | ~n2628;
  assign n8938 = n2636 | n2637;
  assign n8939 = n2642 | n2643;
  assign n8940 = n2644 | n2645;
  assign n8941 = n2646 | ~n2647;
  assign n8942 = n2649 | n2650;
  assign n8943 = n2651 | n2652;
  assign n8944 = n2653 | ~n2654;
  assign n8945 = n2665 | ~n2666;
  assign n8946 = n2682 | n2683;
  assign n8947 = n2695 | n2691 | n2694;
  assign n8948 = n2700 | ~n2701;
  assign n8949 = n2709 | n2710;
  assign n8950 = n2716 | n2717;
  assign n8951 = n2724 | ~n2725;
  assign n8952 = n2728 | n2729;
  assign n8953 = n2730 | n2731;
  assign n8954 = n2737 | ~n2738;
  assign n8955 = n2742 | ~n2743;
  assign n8956 = n2755 | ~n2756;
  assign n8957 = n2766 | n2767;
  assign n8958 = n2778 | n2779;
  assign n8959 = n2787 | n2788;
  assign n8960 = n2793 | ~n2794;
  assign n8961 = n2802 | n2803;
  assign n8962 = n2809 | ~n2810;
  assign n8963 = n2814 | n2815;
  assign n8964 = n2816 | n2817;
  assign n8965 = n2818 | ~n2819;
  assign n8966 = n2824 | ~n2825;
  assign n8967 = n2834 | n2835;
  assign n8968 = n2845 | n2846;
  assign n8969 = n2859 | n2855 | n2858;
  assign n8970 = n2864 | ~n2865;
  assign n8971 = n2887 | n2888;
  assign n8972 = n2896 | n2897;
  assign n8973 = n2902 | ~n2903;
  assign n8974 = n2915 | n2911 | n2914;
  assign n8975 = n2924 | ~n2925;
  assign n8976 = n2940 | n2941;
  assign n8977 = n2949 | n2950;
  assign n8978 = n2955 | ~n2956;
  assign n8979 = n2964 | n2965;
  assign n8980 = n2972 | n2973;
  assign n8981 = n2974 | n2975;
  assign n8982 = n2976 | ~n2977;
  assign n8983 = n2986 | n2987;
  assign n8984 = n2997 | n2998;
  assign n8985 = n3001 | n3002;
  assign n8986 = n3004 | n3005;
  assign n8987 = n3007 | n3008;
  assign n8988 = n3009 | ~n3010;
  assign n8989 = n3018 | n3019;
  assign n8990 = n3027 | n3028;
  assign n8991 = n3036 | n3037;
  assign n8992 = n3042 | ~n3043;
  assign n8993 = n3053 | n3054;
  assign n8994 = n3063 | n3064;
  assign n8995 = n3071 | n3072;
  assign n8996 = n3080 | n3081;
  assign n8997 = n3086 | ~n3087;
  assign n8998 = n3090 | n3091;
  assign n8999 = n3092 | n3093;
  assign n9000 = n3111 | n3112;
  assign n9001 = ~n3119 | n3115 | n3118;
  assign n9002 = n3122 | n3123;
  assign n9003 = ~n3129 | n3125 | ~n3128;
  assign n9004 = n3144 | ~n3145;
  assign n9005 = n3151 | n3152;
  assign n9006 = n3158 | n3159;
  assign n9007 = n3168 | n3165 | ~n3167;
  assign n9008 = n3179 | n3176 | ~n3178;
  assign n9009 = n3190 | n3187 | ~n3189;
  assign n9010 = n3202 | n3199 | ~n3201;
  assign n9011 = n3213 | n3210 | ~n3212;
  assign n9012 = n3225 | n3222 | ~n3224;
  assign n9013 = n3232 | n3229 | ~n3231;
  assign n9014 = n3246 | ~n3247;
  assign n9015 = n3257 | ~n3258;
  assign n9016 = n3268 | ~n3269;
  assign n9017 = n3279 | n3280;
  assign n9018 = n3283 | n3284;
  assign n9019 = n3319 | n3320;
  assign n9020 = n3335 | n3336;
  assign n9021 = n3354 | n3348 | n3353;
  assign n9022 = n3365 | n3366;
  assign n9023 = n3369 | n3370;
  assign n9024 = n3376 | n3377;
  assign n9025 = n3380 | n3381;
  assign n9026 = n3407 | n3398 | n3406;
  assign n9027 = n3410 | n3411;
  assign n9028 = n3414 | n3415;
  assign n9029 = n3419 | n3420;
  assign n9030 = n3436 | n3437;
  assign n9031 = n3443 | n3444;
  assign n9032 = n3447 | n3448;
  assign n9033 = n3453 | n3454;
  assign n9034 = n3459 | n3460;
  assign n9035 = n3466 | n3467;
  assign n9036 = n3475 | n3476;
  assign n9037 = n3482 | n3483;
  assign n9038 = n3488 | n3489;
  assign n9039 = n3497 | n3494 | n3496;
  assign n9040 = n3512 | n3513;
  assign n9041 = n3519 | n3520;
  assign n9042 = n3532 | n3533;
  assign n9043 = n3541 | n3542;
  assign n9044 = n3551 | n3548 | n3550;
  assign n9045 = n3565 | n3561 | n3564;
  assign n9046 = n3575 | n3576;
  assign n9047 = n3579 | n3580;
  assign n9048 = n3591 | n3592;
  assign n9049 = n3598 | n3599;
  assign n9050 = n3602 | n3603;
  assign n9051 = n3615 | n3616;
  assign n9052 = n3622 | n3623;
  assign n9053 = n3625 | n3626;
  assign n9054 = n3641 | n3642;
  assign n9055 = n3654 | n3655;
  assign n9056 = n3661 | n3662;
  assign n9057 = n3667 | n3668;
  assign n9058 = n3678 | n3679;
  assign n9059 = n3682 | n3683;
  assign n9060 = n3686 | n3687;
  assign n9061 = n3702 | n3703;
  assign n9062 = n3713 | n3714;
  assign n9063 = n3727 | n3728;
  assign n9064 = n3740 | n3741;
  assign n9065 = n3749 | n3750;
  assign n9066 = n3760 | n3761;
  assign n9067 = n3772 | n3773;
  assign n9068 = n3782 | n3783;
  assign n9069 = n3803 | n3804;
  assign n9070 = n3818 | n3815 | n3817;
  assign n9071 = n3845 | n3835 | n3844;
  assign n9072 = n3862 | n3863;
  assign n9073 = n3868 | n3869;
  assign n9074 = n3882 | n3883;
  assign n9075 = n3892 | n3893;
  assign n9076 = n3904 | n3900 | n3903;
  assign n9077 = n3910 | n3911;
  assign n9078 = n3921 | n3918 | n3920;
  assign n9079 = n3940 | n3941;
  assign n9080 = n3955 | n3956;
  assign n9081 = n3959 | n3960;
  assign n9082 = n3961 | n3962;
  assign n9083 = n3963 | ~n3964;
  assign n9084 = n3970 | n3971;
  assign n9085 = n3974 | n3975;
  assign n9086 = n3978 | n3979;
  assign n9087 = n3987 | n3988;
  assign n9088 = n4004 | n4005;
  assign n9089 = n4017 | n4018;
  assign n9090 = n4023 | n4024;
  assign n9091 = n4029 | n4030;
  assign n9092 = n4043 | n4044;
  assign n9093 = n4049 | ~n4050;
  assign n9094 = n4056 | n4057;
  assign n9095 = n4066 | n4067;
  assign n9096 = n4074 | ~n4075;
  assign n9097 = n4082 | n4083;
  assign n9098 = n4088 | ~n4089;
  assign n9099 = n4094 | ~n4095;
  assign n9100 = n4120 | n4115 | n4119;
  assign n9101 = n4132 | n4133;
  assign n9102 = n4141 | n4142;
  assign n9103 = n4156 | n4157;
  assign n9104 = n4174 | n4175;
  assign n9105 = n4178 | n4179;
  assign n9106 = n4183 | n4184;
  assign n9107 = n4187 | n4188;
  assign n9108 = n4191 | n4192;
  assign n9109 = n4207 | n4208;
  assign n9110 = n4213 | ~n4214;
  assign n9111 = n4219 | ~n4220;
  assign n9112 = n4221 | n4222;
  assign n9113 = n4234 | n4235;
  assign n9114 = n4240 | ~n4241;
  assign n9115 = n4246 | ~n4247;
  assign n9116 = n4255 | ~n4256;
  assign n9117 = n4261 | ~n4262;
  assign n9118 = n4267 | ~n4268;
  assign n9119 = n4279 | ~n4280;
  assign n9120 = n4290 | ~n4291;
  assign n9121 = n4295 | ~n4296;
  assign n9122 = n4298 | n4299;
  assign n9123 = n4304 | n4305;
  assign n9124 = n4341 | n4342;
  assign n9125 = n4352 | n4353;
  assign n9126 = n4358 | n4359;
  assign n9127 = n4372 | n4373;
  assign n9128 = n4390 | ~n4391;
  assign n9129 = n4394 | n4395;
  assign n9130 = n4409 | ~n4410;
  assign n9131 = n4415 | ~n4416;
  assign n9132 = n4421 | ~n4422;
  assign n9133 = n4430 | ~n4431;
  assign n9134 = n4436 | n4437;
  assign n9135 = n4441 | n4442;
  assign n9136 = n4445 | ~n4446;
  assign n9137 = n4454 | ~n4455;
  assign n9138 = n4459 | n4460;
  assign n9139 = n4468 | ~n4469;
  assign n9140 = n4485 | n4486;
  assign n9141 = n4488 | n4489;
  assign n9142 = n4501 | n4502;
  assign n9143 = n4507 | ~n4508;
  assign n9144 = n4517 | ~n4518;
  assign n9145 = n4522 | n4523;
  assign n9146 = n4528 | ~n4529;
  assign n9147 = n4536 | n4537;
  assign n9148 = n4543 | n4544;
  assign n9149 = n4545 | n4546;
  assign n9150 = n4547 | ~n4548;
  assign n9151 = n4573 | n4574;
  assign n9152 = n4580 | ~n4581;
  assign n9153 = n4590 | n4585 | n4589;
  assign n9154 = n4592 | n4593;
  assign n9155 = n4604 | ~n4605;
  assign n9156 = n4610 | ~n4611;
  assign n9157 = n4622 | ~n4623;
  assign n9158 = n4626 | n4627;
  assign n9159 = n4635 | ~n4636;
  assign n9160 = n4644 | ~n4645;
  assign n9161 = n4656 | n4657;
  assign n9162 = n4658 | n4659;
  assign n9163 = n4675 | ~n4676;
  assign n9164 = n4681 | n4682;
  assign n9165 = n4683 | n4684;
  assign n9166 = n4685 | ~n4686;
  assign n9167 = n4689 | n4690;
  assign n9168 = n4691 | n4692;
  assign n9169 = n4693 | ~n4694;
  assign n9170 = n4703 | n4704;
  assign n9171 = n4705 | n4706;
  assign n9172 = n4712 | n4713;
  assign n9173 = n4722 | n4723;
  assign n9174 = n4726 | ~n4727;
  assign n9175 = n4735 | n4736;
  assign n9176 = n4749 | n4750;
  assign n9177 = n4759 | ~n4760;
  assign n9178 = n4764 | n4765;
  assign n9179 = n4773 | n4774;
  assign n9180 = n4777 | n4778;
  assign n9181 = n4779 | n4780;
  assign n9182 = n4783 | n4784;
  assign n9183 = n4785 | n4786;
  assign n9184 = n4787 | ~n4788;
  assign n9185 = n4798 | ~n4799;
  assign n9186 = n4801 | ~n4802;
  assign n9187 = n4808 | ~n4809;
  assign n9188 = n4811 | ~n4812;
  assign n9189 = n4828 | n4826 | n4827;
  assign n9190 = n4838 | n4839;
  assign n9191 = n4844 | n4845;
  assign n9192 = n4846 | n4847;
  assign n9193 = n4850 | n4851;
  assign n9194 = n4853 | ~n4854;
  assign n9195 = ~n4859 | n4856 | ~n4858;
  assign n9196 = n4864 | ~n4865;
  assign n9197 = n4879 | ~n4880;
  assign n9198 = n4888 | ~n4889;
  assign n9199 = n4894 | ~n4895;
  assign n9200 = n4912 | ~n4913;
  assign n9201 = n4925 | ~n4926;
  assign n9202 = n4942 | ~n4943;
  assign n9203 = n4948 | n4949;
  assign n9204 = n4950 | n4951;
  assign n9205 = n4952 | ~n4953;
  assign n9206 = n4963 | ~n4964;
  assign n9207 = n4993 | ~n4994;
  assign n9208 = n5001 | ~n5002;
  assign n9209 = n5018 | n5019;
  assign n9210 = n5027 | n5028;
  assign n9211 = n5031 | ~n5032;
  assign n9212 = n5040 | n5041;
  assign n9213 = n5053 | n5054;
  assign n9214 = n5063 | ~n5064;
  assign n9215 = n5068 | n5069;
  assign n9216 = n5077 | n5078;
  assign n9217 = n5084 | n5085;
  assign n9218 = n5086 | n5087;
  assign n9219 = n5088 | ~n5089;
  assign n9220 = n5103 | ~n5104;
  assign n9221 = n5114 | ~n5115;
  assign n9222 = n5119 | n5120;
  assign n9223 = n5121 | n5122;
  assign n9224 = n5123 | ~n5124;
  assign n9225 = n5134 | ~n5135;
  assign n9226 = n5141 | ~n5142;
  assign n9227 = n5161 | n5156 | n5160;
  assign n9228 = n5171 | n5172;
  assign n9229 = n5195 | n5184 | n5194;
  assign n9230 = n5198 | n5199;
  assign n9231 = n5219 | n5220;
  assign n9232 = n5234 | n5235;
  assign n9233 = n5240 | ~n5241;
  assign n9234 = n5243 | n5244;
  assign n9235 = n5268 | ~n5269;
  assign n9236 = n5291 | n5292;
  assign n9237 = n5298 | n5299;
  assign n9238 = n5304 | ~n5305;
  assign n9239 = n5310 | ~n5311;
  assign n9240 = n5316 | ~n5317;
  assign n9241 = n5322 | ~n5323;
  assign n9242 = n5344 | ~n5345;
  assign n9243 = n5359 | n5360;
  assign n9244 = n5375 | n5376;
  assign n9245 = n5396 | n5397;
  assign n9246 = n5402 | ~n5403;
  assign n9247 = n5409 | n5410;
  assign n9248 = n5414 | n5415;
  assign n9249 = n5422 | n5423;
  assign n9250 = n5433 | n5434;
  assign n9251 = n5439 | n5440;
  assign n9252 = n5450 | n5451;
  assign n9253 = n5457 | ~n5458;
  assign n9254 = n5475 | ~n5476;
  assign n9255 = n5493 | ~n5494;
  assign n9256 = n5502 | ~n5503;
  assign n9257 = n5515 | ~n5516;
  assign n9258 = n5530 | ~n5531;
  assign n9259 = n5538 | ~n5539;
  assign n9260 = n5548 | n5549;
  assign n9261 = n5582 | n5575 | n5581;
  assign n9262 = n5599 | ~n5600;
  assign n9263 = n5610 | n5611;
  assign n9264 = n5620 | n5621;
  assign n9265 = n5633 | n5634;
  assign n9266 = n5635 | n5636;
  assign n9267 = n5644 | ~n5645;
  assign n9268 = ~n5670 | n5665 | n5669;
  assign n9269 = n5680 | n5681;
  assign n9270 = n5682 | n5683;
  assign n9271 = n5694 | ~n5695;
  assign n9272 = n5706 | n5707;
  assign n9273 = n5708 | n5709;
  assign n9274 = n5726 | n5727;
  assign n9275 = n5749 | n5750;
  assign n9276 = n5782 | ~n5783;
  assign n9277 = n5796 | n5797;
  assign n9278 = n5798 | n5799;
  assign n9279 = n5806 | ~n5807;
  assign n9280 = n5813 | ~n5814;
  assign n9281 = n5842 | n5834 | n5841;
  assign n9282 = n5857 | n5858;
  assign n9283 = n5873 | n5874;
  assign n9284 = n5876 | n5877;
  assign n9285 = n5884 | n5885;
  assign n9286 = n5892 | n5893;
  assign n9287 = n5894 | n5895;
  assign n9288 = n5907 | n5908;
  assign n9289 = n5909 | n5910;
  assign n9290 = n5936 | ~n5937;
  assign n9291 = n5945 | ~n5946;
  assign n9292 = n5951 | ~n5952;
  assign n9293 = n5957 | ~n5958;
  assign n9294 = n5970 | ~n5971;
  assign n9295 = n5979 | ~n5980;
  assign n9296 = n5985 | ~n5986;
  assign n9297 = n5991 | ~n5992;
  assign n9298 = n6000 | n6001;
  assign n9299 = n6016 | n6017;
  assign n9300 = n6027 | n6028;
  assign n9301 = n6033 | n6034;
  assign n9302 = n6039 | n6040;
  assign n9303 = n6055 | n6056;
  assign n9304 = n6063 | n6064;
  assign n9305 = n6071 | n6072;
  assign n9306 = n6076 | n6077;
  assign n9307 = n6095 | n6096;
  assign n9308 = n6100 | n6101;
  assign n9309 = n6109 | n6110;
  assign n9310 = n6117 | n6118;
  assign n9311 = n6126 | n6123 | n6125;
  assign n9312 = n6137 | n6138;
  assign n9313 = n6154 | n6155;
  assign n9314 = n6158 | n6159;
  assign n9315 = n6174 | n6175;
  assign n9316 = n6184 | n6185;
  assign n9317 = n6190 | n6191;
  assign n9318 = n6195 | n6196;
  assign n9319 = n6200 | n6201;
  assign n9320 = n6206 | n6207;
  assign n9321 = n6219 | n6220;
  assign n9322 = n6231 | n6232;
  assign n9323 = n6246 | n6247;
  assign n9324 = ~n6255 | n6250 | ~n6254;
  assign n9325 = n6259 | ~n6260;
  assign n9326 = n6262 | ~n6263;
  assign n9327 = n6267 | n6268;
  assign n9328 = n6269 | n6270;
  assign n9329 = n6274 | n6275;
  assign n9330 = n6276 | n6277;
  assign n9331 = n6278 | ~n6279;
  assign n9332 = n6284 | ~n6285;
  assign n9333 = n6297 | n6298;
  assign n9334 = n6305 | n6306;
  assign n9335 = n6314 | n6315;
  assign n9336 = n6318 | n6319;
  assign n9337 = n6329 | n6330;
  assign n9338 = n6331 | n6332;
  assign n9339 = n6333 | n6334;
  assign n9340 = n6337 | ~n6338;
  assign n9341 = n6344 | n6345;
  assign n9342 = n6351 | n6352;
  assign n9343 = n6353 | n6354;
  assign n9344 = n6366 | n6367;
  assign n9345 = n6368 | n6369;
  assign n9346 = n6380 | ~n6381;
  assign n9347 = n6401 | n6402;
  assign n9348 = n6403 | n6404;
  assign n9349 = n6405 | ~n6406;
  assign n9350 = n6409 | n6410;
  assign n9351 = n6411 | n6412;
  assign n9352 = n6413 | ~n6414;
  assign n9353 = n6417 | n6418;
  assign n9354 = n6419 | n6420;
  assign n9355 = n6421 | ~n6422;
  assign n9356 = n6427 | ~n6428;
  assign n9357 = n6440 | ~n6441;
  assign n9358 = n6449 | ~n6450;
  assign n9359 = n6455 | ~n6456;
  assign n9360 = n6461 | ~n6462;
  assign n9361 = n6472 | n6473;
  assign n9362 = n6488 | n6489;
  assign n9363 = n6502 | n6503;
  assign n9364 = n6513 | n6514;
  assign n9365 = n6520 | n6521;
  assign n9366 = n6526 | ~n6527;
  assign n9367 = n6529 | n6530;
  assign n9368 = n6535 | n6536;
  assign n9369 = n6537 | n6538;
  assign n9370 = n6550 | n6551;
  assign n9371 = n6552 | n6553;
  assign n9372 = n6564 | ~n6565;
  assign n9373 = n6582 | n6583;
  assign n9374 = n6587 | n6588;
  assign n9375 = n6589 | n6590;
  assign n9376 = n6591 | ~n6592;
  assign n9377 = n6595 | n6596;
  assign n9378 = n6597 | n6598;
  assign n9379 = n6599 | ~n6600;
  assign n9380 = n6603 | n6604;
  assign n9381 = n6605 | n6606;
  assign n9382 = n6607 | ~n6608;
  assign n9383 = n6613 | ~n6614;
  assign n9384 = n6626 | ~n6627;
  assign n9385 = n6635 | ~n6636;
  assign n9386 = n6641 | ~n6642;
  assign n9387 = n6647 | ~n6648;
  assign n9388 = n6653 | ~n6654;
  assign n9389 = n6657 | n6658;
  assign n9390 = n6664 | n6665;
  assign n9391 = n6677 | n6678;
  assign n9392 = n6691 | n6692;
  assign n9393 = n6697 | n6698;
  assign n9394 = n6703 | ~n6704;
  assign n9395 = n6721 | ~n6722;
  assign n9396 = n6724 | n6725;
  assign n9397 = n6726 | n6727;
  assign n9398 = n6738 | n6739;
  assign n9399 = n6740 | n6741;
  assign n9400 = n6752 | ~n6753;
  assign n9401 = n6770 | n6771;
  assign n9402 = n6775 | n6776;
  assign n9403 = n6777 | n6778;
  assign n9404 = n6779 | ~n6780;
  assign n9405 = n6791 | ~n6792;
  assign n9406 = n6797 | n6798;
  assign n9407 = n6805 | ~n6806;
  assign n9408 = n6837 | n6838;
  assign n9409 = n6853 | n6854;
  assign n9410 = n6859 | ~n6860;
  assign n9411 = n6863 | n6864;
  assign n9412 = n6870 | ~n6871;
  assign n9413 = n6887 | n6888;
  assign n9414 = n6889 | n6890;
  assign n9415 = n6911 | n6912;
  assign n9416 = n6913 | n6914;
  assign n9417 = n6918 | n6919;
  assign n9418 = n6924 | ~n6925;
  assign n9419 = n6930 | ~n6931;
  assign n9420 = n6939 | ~n6940;
  assign n9421 = n6943 | n6944;
  assign n9422 = n6945 | n6946;
  assign n9423 = n6947 | ~n6948;
  assign n9424 = n6953 | ~n6954;
  assign n9425 = n6963 | n6964;
  assign n9426 = n6993 | n6994;
  assign n9427 = n7006 | n7007;
  assign n9428 = n7026 | n7027;
  assign n9429 = n7043 | n7044;
  assign n9430 = n7045 | n7046;
  assign n9431 = n7067 | ~n7068;
  assign n9432 = n7074 | n7075;
  assign n9433 = n7080 | ~n7081;
  assign n9434 = n7086 | ~n7087;
  assign n9435 = n7092 | ~n7093;
  assign n9436 = n7096 | n7097;
  assign n9437 = n7103 | ~n7104;
  assign n9438 = n7107 | n7108;
  assign n9439 = n7114 | ~n7115;
  assign n9440 = n7118 | n7119;
  assign n9441 = n7129 | n7130;
  assign n9442 = n7152 | n7153;
  assign n9443 = n7176 | ~n7177;
  assign n9444 = n7185 | n7186;
  assign n9445 = n7193 | n7194;
  assign n9446 = n7195 | n7196;
  assign n9447 = n7217 | ~n7218;
  assign n9448 = n7224 | n7225;
  assign n9449 = n7230 | ~n7231;
  assign n9450 = n7236 | ~n7237;
  assign n9451 = n7242 | ~n7243;
  assign n9452 = n7246 | n7247;
  assign n9453 = n7253 | ~n7254;
  assign n9454 = n7257 | n7258;
  assign n9455 = n7272 | n7273;
  assign n9456 = n7284 | n7285;
  assign n9457 = n7290 | n7291;
  assign n9458 = n7306 | n7307;
  assign n9459 = n7328 | n7329;
  assign n9460 = n7335 | ~n7336;
  assign n9461 = n7352 | ~n7353;
  assign n9462 = n7366 | n7367;
  assign n9463 = n7368 | n7369;
  assign n9464 = n7380 | n7381;
  assign n9465 = n7382 | n7383;
  assign n9466 = n7384 | ~n7385;
  assign n9467 = n7390 | ~n7391;
  assign n9468 = n7396 | ~n7397;
  assign n9469 = n7402 | ~n7403;
  assign n9470 = n7408 | ~n7409;
  assign n9471 = n7414 | ~n7415;
  assign n9472 = n7427 | n7428;
  assign n9473 = n7442 | n7443;
  assign n9474 = n7462 | n7463;
  assign n9475 = n7468 | n7469;
  assign n9476 = n7470 | n7471;
  assign n9477 = n7493 | ~n7494;
  assign n9478 = n7502 | n7503;
  assign n9479 = n7504 | n7505;
  assign n9480 = n7506 | ~n7507;
  assign n9481 = n7515 | ~n7516;
  assign n9482 = n7519 | n7520;
  assign n9483 = n7536 | n7537;
  assign n9484 = n7550 | n7551;
  assign n9485 = n7560 | n7561;
  assign n9486 = n7575 | n7576;
  assign n9487 = n7599 | ~n7600;
  assign n9488 = n7608 | n7609;
  assign n9489 = n7627 | n7628;
  assign n9490 = n7629 | n7630;
  assign n9491 = n7637 | ~n7638;
  assign n9492 = n7643 | ~n7644;
  assign n9493 = n7649 | ~n7650;
  assign n9494 = n7655 | ~n7656;
  assign n9495 = n7661 | ~n7662;
  assign n9496 = n7683 | n7684;
  assign n9497 = n7697 | n7698;
  assign n9498 = n7719 | n7720;
  assign n9499 = n7726 | ~n7727;
  assign n9500 = n7735 | ~n7736;
  assign n9501 = n7745 | n7746;
  assign n9502 = n7747 | n7748;
  assign n9503 = n7756 | n7757;
  assign n9504 = n7759 | ~n7760;
  assign n9505 = n7761 | n7762;
  assign n9506 = n7766 | n7767;
  assign n9507 = n7773 | ~n7774;
  assign n9508 = n7779 | ~n7780;
  assign n9509 = n7783 | n7784;
  assign n9510 = n7796 | n7797;
  assign n9511 = n7814 | n7815;
  assign n9512 = n7834 | n7835;
  assign n9513 = n7850 | ~n7851;
  assign n9514 = n7860 | ~n7861;
  assign n9515 = n7869 | n7866 | ~n7868;
  assign n9516 = n7874 | ~n7875;
  assign n9517 = n7878 | n7879;
  assign n9518 = n7897 | n7898;
  assign n9519 = n7918 | n7919;
  assign n9520 = n7920 | n7921;
  assign n9521 = n7924 | n7925;
  assign n9522 = n7930 | ~n7931;
  assign n9523 = n7933 | n7934;
  assign n9524 = n7941 | n7942;
  assign n9525 = n7943 | n7944;
  assign n9526 = n7950 | ~n7951;
  assign n9527 = n7956 | ~n7957;
  assign n9528 = n7962 | ~n7963;
  assign n9529 = n7968 | ~n7969;
  assign n9530 = n7985 | n7981 | n7984;
  assign n9531 = n8002 | n7999 | n8001;
  assign n9532 = n8022 | n8023;
  assign n9533 = n8029 | n8030;
  assign n9534 = n8031 | n8032;
  assign n9535 = n8043 | n8044;
  assign n9536 = n8045 | n8046;
  assign n9537 = n8047 | ~n8048;
  assign n9538 = n8053 | ~n8054;
  assign n9539 = n8072 | n8067 | n8071;
  assign n9540 = n8085 | n8086;
  assign n9541 = n8102 | n8103;
  assign n9542 = n8108 | n8109;
  assign n9543 = n8114 | ~n8115;
  assign n9544 = n8127 | n8128;
  assign n9545 = n8133 | ~n8134;
  assign n9546 = n8142 | n8143;
  assign n9547 = n8144 | n8145;
  assign n9548 = n8146 | ~n8147;
  assign n9549 = n8172 | n8173;
  assign n9550 = n8190 | n8191;
  assign n9551 = n8212 | ~n8213;
  assign n9552 = n8218 | n8219;
  assign n9553 = n8220 | n8221;
  assign n9554 = n8224 | n8225;
  assign n9555 = n8226 | n8227;
  assign n9556 = n8228 | n8229;
  assign n9557 = n8230 | ~n8231;
  assign n9558 = n8240 | n8241;
  assign n9559 = n8244 | n8245;
  assign n9560 = n8250 | n8251;
  assign n9561 = n8268 | n8269;
  assign n9562 = n8274 | n8275;
  assign n9563 = n8280 | ~n8281;
  assign n9564 = n8292 | n8293;
  assign n9565 = n8308 | n8309;
  assign n9566 = n8314 | n8312 | n8313;
  assign n9567 = n8325 | n8323 | n8324;
  assign n9568 = n8336 | ~n8337;
  assign n9569 = n8343 | n8344;
  assign n9570 = n8346 | ~n8347;
  assign n9571 = n8348 | n8349;
  assign n9572 = n8350 | n8351;
  assign n9573 = n8352 | ~n8353;
  assign n9574 = n8377 | n8378;
  assign n9575 = n8391 | n8392;
  assign n9576 = n8402 | n8403;
  assign n9577 = n8404 | n8405;
  assign n9578 = n8415 | n8416;
  assign n9579 = n8436 | n8433 | n8435;
  assign n9580 = n8445 | ~n8446;
  assign n9581 = n8449 | n8450;
  assign n9582 = n8451 | n8452;
  assign n9583 = n8464 | n8465;
  assign n9584 = n8478 | n8479;
  assign n9585 = n8494 | n8495;
  assign n9586 = n8496 | n8497;
  assign n9587 = n8519 | n8520;
  assign n9588 = n8529 | ~n8530;
  assign n9589 = n8533 | n8534;
  assign n9590 = n8535 | n8536;
  assign n9591 = n8543 | n8544;
  assign n9592 = n8559 | n8560;
  assign n9593 = n8561 | n8562;
  assign n9594 = n8584 | n8579 | n8583;
  assign n9595 = n8587 | n8585 | n8586;
  assign n9596 = n8598 | n8594 | n8597;
  assign n9597 = n8609 | n8605 | n8608;
  assign n9598 = n8611 | n8612;
  assign n9599 = n8617 | n8615 | n8616;
  assign po0  = ~n9331;
  assign po1  = ~n6516;
  assign po2  = ~n6712;
  assign po4  = ~n7021;
  assign po5  = ~n7167;
  assign po6  = ~n7321;
  assign po7  = ~n7457;
  assign po8  = ~n7590;
  assign po9  = ~n7712;
  assign po10  = ~n7829;
  assign po11  = ~n7912;
  assign po12  = ~n8016;
  assign po13  = ~n8123;
  assign po14  = ~n8205;
  assign po15  = ~n8289;
  assign po16  = ~n8361;
  assign po18  = ~n8453;
  assign po19  = ~n8498;
  assign po20  = ~n8537;
  assign po21  = ~n8563;
  assign po22  = ~n8588;
  assign po23  = ~n9597;
endmodule
