module top ( 
    pi0 , pi1 , pi2 , pi3 ,
    pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 ,
    po0 , po1 , po2 , po3 ,
    po4 , po5 , po6 , po7 ,
    po8 , po9 , po10   );
  input  pi0 , pi1 , pi2 ,
    pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 ;
  output po0 , po1 , po2 ,
    po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 ;
  wire n22, n23, n24, n25, n26, n27, n28,
    n29, n30, n31, n32, n33, n34, n35, n36,
    n37, n38, n39, n40, n41, n42, n43, n44,
    n45, n46, n47, n48, n49, n50, n51, n52,
    n53, n54, n55, n56, n57, n58, n59, n60,
    n61, n62, n63, n64, n65, n66, n67, n68,
    n69, n70, n71, n72, n73, n74, n75, n76,
    n77, n78, n79, n80, n81, n82, n83, n84,
    n85, n86, n87, n88, n89, n90, n91, n92,
    n93, n94, n95, n96, n97, n98, n99,
    n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n109, n110, n111, n112, n113,
    n114, n115, n116, n117, n118, n119, n120,
    n121, n122, n123, n124, n125, n126, n127,
    n128, n129, n130, n131, n132, n133, n134,
    n135, n136, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n401, n402, n403, n404,
    n405, n406, n408, n409, n410, n412, n413,
    n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n486, n487, n488, n489, n490, n491,
    n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505,
    n506, n507, n508, n509, n510, n511, n512,
    n513, n514, n515, n516, n517, n518, n519,
    n520, n521, n522, n523, n524, n525, n526,
    n527, n528, n529, n530, n531, n532, n533,
    n534, n535, n536, n537, n538, n539, n540,
    n541, n542, n543, n544, n545, n546, n547,
    n548, n549, n550, n551, n552, n553, n554,
    n555, n556, n557, n558, n559, n560, n561,
    n562, n563, n564, n565, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626,
    n627, n628, n629, n630, n631, n632, n633,
    n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647,
    n648, n649, n651, n652, n653, n654, n655;
  assign n22 = pi7  & pi8 ;
  assign n23 = ~pi5  & n22;
  assign n24 = ~pi7  & pi9 ;
  assign n25 = ~n23 & ~n24;
  assign n26 = pi1  & ~n25;
  assign n27 = pi1  & ~pi7 ;
  assign n28 = ~pi5  & ~pi9 ;
  assign n29 = ~n27 & n28;
  assign n30 = ~n26 & ~n29;
  assign n31 = pi0  & ~pi2 ;
  assign n32 = ~n30 & n31;
  assign n33 = pi2  & ~pi9 ;
  assign n34 = ~pi0  & ~pi1 ;
  assign n35 = n33 & n34;
  assign n36 = n23 & n35;
  assign n37 = ~n32 & ~n36;
  assign n38 = ~pi3  & ~n37;
  assign n39 = ~pi3  & ~pi5 ;
  assign n40 = ~pi0  & pi9 ;
  assign n41 = pi1  & ~n40;
  assign n42 = ~pi1  & pi9 ;
  assign n43 = n39 & ~n42;
  assign n44 = ~n41 & n43;
  assign n45 = pi0  & ~pi9 ;
  assign n46 = ~pi1  & ~n45;
  assign n47 = pi1  & ~pi9 ;
  assign n48 = ~pi7  & ~n47;
  assign n49 = ~n46 & n48;
  assign n50 = ~n44 & ~n49;
  assign n51 = ~pi2  & ~n50;
  assign n52 = ~pi2  & ~pi3 ;
  assign n53 = pi9  & ~n52;
  assign n54 = pi0  & pi3 ;
  assign n55 = ~n53 & ~n54;
  assign n56 = ~pi1  & ~n55;
  assign n57 = pi1  & ~pi3 ;
  assign n58 = pi0  & ~n47;
  assign n59 = ~n40 & ~n45;
  assign n60 = ~pi2  & pi5 ;
  assign n61 = n59 & n60;
  assign n62 = ~n33 & ~n61;
  assign n63 = ~n58 & ~n62;
  assign n64 = ~n56 & ~n57;
  assign n65 = ~n63 & n64;
  assign n66 = ~pi7  & ~n65;
  assign n67 = ~n51 & ~n66;
  assign n68 = ~pi8  & ~n67;
  assign n69 = ~n38 & ~n68;
  assign n70 = ~pi6  & ~n69;
  assign n71 = ~pi2  & ~n45;
  assign n72 = pi6  & ~n71;
  assign n73 = pi1  & n59;
  assign n74 = n52 & n73;
  assign n75 = ~n72 & ~n74;
  assign n76 = pi5  & ~n75;
  assign n77 = pi2  & pi9 ;
  assign n78 = ~pi2  & n47;
  assign n79 = ~n77 & ~n78;
  assign n80 = ~pi0  & ~pi3 ;
  assign n81 = pi6  & n80;
  assign n82 = ~n79 & n81;
  assign n83 = ~n76 & ~n82;
  assign n84 = pi8  & ~n83;
  assign n85 = ~pi3  & ~pi8 ;
  assign n86 = ~pi1  & ~pi9 ;
  assign n87 = pi1  & pi9 ;
  assign n88 = ~n86 & ~n87;
  assign n89 = n85 & ~n88;
  assign n90 = ~pi1  & ~pi2 ;
  assign n91 = ~pi0  & n90;
  assign n92 = n89 & n91;
  assign n93 = pi1  & ~pi8 ;
  assign n94 = pi2  & ~pi3 ;
  assign n95 = n42 & n94;
  assign n96 = ~n93 & ~n95;
  assign n97 = ~pi0  & ~n96;
  assign n98 = pi3  & ~pi6 ;
  assign n99 = pi2  & pi3 ;
  assign n100 = n86 & ~n98;
  assign n101 = ~n99 & n100;
  assign n102 = ~n77 & ~n101;
  assign n103 = ~pi8  & ~n102;
  assign n104 = ~n97 & ~n103;
  assign n105 = ~pi5  & ~n104;
  assign n106 = ~pi1  & ~n40;
  assign n107 = ~pi8  & ~n106;
  assign n108 = ~pi1  & pi2 ;
  assign n109 = n45 & n108;
  assign n110 = ~n107 & ~n109;
  assign n111 = ~pi5  & ~n110;
  assign n112 = ~pi0  & ~pi2 ;
  assign n113 = ~pi6  & pi9 ;
  assign n114 = n112 & ~n113;
  assign n115 = n42 & n114;
  assign n116 = pi5  & pi6 ;
  assign n117 = pi2  & pi5 ;
  assign n118 = n73 & n117;
  assign n119 = ~n115 & ~n116;
  assign n120 = ~n118 & n119;
  assign n121 = pi8  & ~n120;
  assign n122 = ~n111 & ~n121;
  assign n123 = pi3  & ~n122;
  assign n124 = ~n92 & ~n105;
  assign n125 = ~n84 & n124;
  assign n126 = ~n123 & n125;
  assign n127 = ~pi7  & ~n126;
  assign n128 = ~n70 & ~n127;
  assign n129 = ~pi4  & ~n128;
  assign n130 = ~pi1  & ~pi3 ;
  assign n131 = pi6  & ~pi9 ;
  assign n132 = pi4  & pi9 ;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~pi8  & ~n116;
  assign n135 = ~n133 & n134;
  assign n136 = pi4  & pi8 ;
  assign n137 = ~pi6  & ~pi9 ;
  assign n138 = ~n136 & ~n137;
  assign n139 = ~pi6  & pi8 ;
  assign n140 = pi5  & ~n139;
  assign n141 = ~n138 & n140;
  assign n142 = ~n135 & ~n141;
  assign n143 = ~pi7  & n112;
  assign n144 = n130 & n143;
  assign n145 = ~n142 & n144;
  assign po0  = n129 | n145;
  assign n147 = pi2  & ~n34;
  assign n148 = pi0  & pi1 ;
  assign n149 = n71 & ~n148;
  assign n150 = ~pi8  & ~n147;
  assign n151 = ~n149 & n150;
  assign n152 = ~pi2  & pi8 ;
  assign n153 = n47 & n152;
  assign n154 = ~n151 & ~n153;
  assign n155 = pi7  & ~n154;
  assign n156 = ~n35 & ~n155;
  assign n157 = ~pi6  & n39;
  assign n158 = ~pi4  & n157;
  assign n159 = ~n156 & n158;
  assign n160 = pi1  & pi2 ;
  assign n161 = pi5  & ~pi8 ;
  assign n162 = ~pi6  & ~n161;
  assign n163 = pi3  & n160;
  assign n164 = ~n162 & n163;
  assign n165 = pi1  & pi5 ;
  assign n166 = pi3  & ~pi8 ;
  assign n167 = n90 & n166;
  assign n168 = ~n165 & ~n167;
  assign n169 = pi0  & ~n168;
  assign n170 = pi5  & ~n52;
  assign n171 = ~n169 & ~n170;
  assign n172 = pi6  & ~n171;
  assign n173 = ~n164 & ~n172;
  assign n174 = pi9  & ~n173;
  assign n175 = ~pi5  & pi8 ;
  assign n176 = ~n85 & ~n175;
  assign n177 = pi0  & n176;
  assign n178 = ~pi8  & n60;
  assign n179 = ~n177 & ~n178;
  assign n180 = ~pi1  & ~n179;
  assign n181 = ~pi0  & pi5 ;
  assign n182 = pi0  & n152;
  assign n183 = pi0  & ~pi5 ;
  assign n184 = ~n181 & ~n183;
  assign n185 = ~n182 & n184;
  assign n186 = pi1  & ~n185;
  assign n187 = ~pi2  & ~pi8 ;
  assign n188 = ~pi0  & ~n52;
  assign n189 = ~n187 & n188;
  assign n190 = ~n186 & ~n189;
  assign n191 = ~n180 & n190;
  assign n192 = ~pi6  & ~n191;
  assign n193 = ~pi1  & pi6 ;
  assign n194 = pi2  & ~n193;
  assign n195 = ~pi1  & ~pi8 ;
  assign n196 = pi3  & ~n195;
  assign n197 = ~n194 & n196;
  assign n198 = ~pi1  & ~pi6 ;
  assign n199 = ~pi0  & pi8 ;
  assign n200 = ~pi2  & ~n148;
  assign n201 = ~n198 & ~n199;
  assign n202 = n200 & n201;
  assign n203 = ~n197 & ~n202;
  assign n204 = ~pi5  & ~n203;
  assign n205 = ~n192 & ~n204;
  assign n206 = ~pi9  & ~n205;
  assign n207 = pi6  & pi9 ;
  assign n208 = ~n175 & ~n207;
  assign n209 = pi6  & pi8 ;
  assign n210 = pi0  & ~n209;
  assign n211 = ~n208 & n210;
  assign n212 = ~pi8  & pi9 ;
  assign n213 = n181 & n212;
  assign n214 = ~n211 & ~n213;
  assign n215 = ~pi2  & ~n214;
  assign n216 = ~pi6  & ~pi8 ;
  assign n217 = pi2  & ~pi5 ;
  assign n218 = ~pi6  & ~n217;
  assign n219 = ~n31 & n175;
  assign n220 = ~n218 & n219;
  assign n221 = ~n216 & ~n220;
  assign n222 = ~pi9  & ~n221;
  assign n223 = ~n215 & ~n222;
  assign n224 = pi1  & ~n223;
  assign n225 = n33 & n139;
  assign n226 = ~n224 & ~n225;
  assign n227 = ~pi3  & ~n226;
  assign n228 = ~n174 & ~n206;
  assign n229 = ~n227 & n228;
  assign n230 = ~pi4  & ~n229;
  assign n231 = ~n136 & ~n161;
  assign n232 = ~pi6  & ~n231;
  assign n233 = ~n132 & ~n232;
  assign n234 = n114 & ~n233;
  assign n235 = ~pi8  & n28;
  assign n236 = ~n45 & ~n208;
  assign n237 = ~n210 & n236;
  assign n238 = ~n235 & ~n237;
  assign n239 = pi2  & ~n238;
  assign n240 = ~pi8  & ~pi9 ;
  assign n241 = pi8  & pi9 ;
  assign n242 = pi0  & n241;
  assign n243 = ~n240 & ~n242;
  assign n244 = pi5  & ~n243;
  assign n245 = ~n31 & ~n33;
  assign n246 = n244 & n245;
  assign n247 = ~n239 & ~n246;
  assign n248 = ~pi4  & ~n247;
  assign n249 = ~n234 & ~n248;
  assign n250 = n130 & ~n249;
  assign n251 = ~n230 & ~n250;
  assign n252 = ~pi7  & ~n251;
  assign po1  = n159 | n252;
  assign n254 = pi6  & ~pi8 ;
  assign n255 = ~pi3  & pi9 ;
  assign n256 = pi1  & n255;
  assign n257 = n254 & n256;
  assign n258 = pi3  & ~n152;
  assign n259 = pi5  & ~n258;
  assign n260 = pi3  & ~n217;
  assign n261 = pi8  & ~n260;
  assign n262 = ~n259 & ~n261;
  assign n263 = pi1  & ~n262;
  assign n264 = ~pi5  & pi6 ;
  assign n265 = ~pi3  & n264;
  assign n266 = n195 & n265;
  assign n267 = ~n263 & ~n266;
  assign n268 = ~pi9  & ~n267;
  assign n269 = ~pi9  & ~n193;
  assign n270 = ~n254 & n269;
  assign n271 = ~pi2  & ~n270;
  assign n272 = ~pi8  & n42;
  assign n273 = ~n271 & ~n272;
  assign n274 = pi3  & ~n273;
  assign n275 = pi2  & ~n139;
  assign n276 = ~pi1  & pi8 ;
  assign n277 = ~n275 & ~n276;
  assign n278 = n170 & ~n277;
  assign n279 = ~n57 & ~n212;
  assign n280 = ~pi6  & ~n255;
  assign n281 = ~n279 & n280;
  assign n282 = ~n257 & ~n281;
  assign n283 = ~n278 & n282;
  assign n284 = ~n274 & n283;
  assign n285 = ~n268 & n284;
  assign n286 = ~pi4  & ~n285;
  assign n287 = ~n241 & ~n254;
  assign n288 = ~pi5  & ~n287;
  assign n289 = ~pi3  & pi4 ;
  assign n290 = n90 & n289;
  assign n291 = ~n288 & n290;
  assign n292 = ~n286 & ~n291;
  assign n293 = ~pi0  & ~n292;
  assign n294 = ~pi5  & n77;
  assign n295 = ~n244 & ~n294;
  assign n296 = pi1  & ~n295;
  assign n297 = ~n240 & ~n241;
  assign n298 = ~n86 & ~n297;
  assign n299 = pi2  & ~n298;
  assign n300 = ~n296 & ~n299;
  assign n301 = ~pi3  & ~n300;
  assign n302 = n53 & n276;
  assign n303 = ~pi2  & ~pi9 ;
  assign n304 = ~n167 & ~n235;
  assign n305 = n303 & ~n304;
  assign n306 = ~n302 & ~n305;
  assign n307 = pi0  & ~n306;
  assign n308 = ~n301 & ~n307;
  assign n309 = ~pi6  & ~n308;
  assign n310 = pi6  & ~n42;
  assign n311 = ~n47 & ~n310;
  assign n312 = pi8  & ~n311;
  assign n313 = ~n89 & ~n312;
  assign n314 = ~pi2  & ~n313;
  assign n315 = pi8  & ~n33;
  assign n316 = pi2  & n87;
  assign n317 = ~n276 & ~n316;
  assign n318 = pi6  & ~n317;
  assign n319 = pi2  & n240;
  assign n320 = ~n315 & ~n319;
  assign n321 = ~n318 & n320;
  assign n322 = pi3  & ~n321;
  assign n323 = ~n314 & ~n322;
  assign n324 = n183 & ~n323;
  assign n325 = ~n309 & ~n324;
  assign n326 = ~pi4  & ~n325;
  assign n327 = ~n293 & ~n326;
  assign n328 = ~pi7  & ~n327;
  assign n329 = n45 & n195;
  assign n330 = pi0  & ~n22;
  assign n331 = n73 & ~n330;
  assign n332 = ~n329 & ~n331;
  assign n333 = ~pi2  & n158;
  assign n334 = ~n332 & n333;
  assign po2  = n328 | n334;
  assign n336 = n264 & n270;
  assign n337 = ~n28 & ~n216;
  assign n338 = n60 & n86;
  assign n339 = ~n265 & ~n338;
  assign n340 = ~n337 & ~n339;
  assign n341 = pi2  & ~n176;
  assign n342 = pi8  & n60;
  assign n343 = ~n341 & ~n342;
  assign n344 = ~pi9  & ~n343;
  assign n345 = ~pi6  & ~n166;
  assign n346 = pi3  & ~pi5 ;
  assign n347 = ~n345 & ~n346;
  assign n348 = ~pi2  & pi3 ;
  assign n349 = pi5  & pi9 ;
  assign n350 = n187 & n349;
  assign n351 = ~n348 & ~n350;
  assign n352 = ~n347 & n351;
  assign n353 = ~n344 & n352;
  assign n354 = pi1  & ~n353;
  assign n355 = ~n340 & ~n354;
  assign n356 = pi0  & ~n355;
  assign n357 = ~pi8  & n264;
  assign n358 = pi5  & pi8 ;
  assign n359 = n113 & n358;
  assign n360 = ~n235 & ~n359;
  assign n361 = pi2  & ~n360;
  assign n362 = pi3  & ~n347;
  assign n363 = ~n357 & ~n361;
  assign n364 = ~n362 & n363;
  assign n365 = pi1  & ~n364;
  assign n366 = pi2  & n264;
  assign n367 = ~n365 & ~n366;
  assign n368 = ~pi0  & ~n367;
  assign n369 = pi2  & n98;
  assign n370 = ~n264 & ~n369;
  assign n371 = n53 & ~n370;
  assign n372 = ~pi5  & ~pi6 ;
  assign n373 = ~n116 & ~n372;
  assign n374 = ~pi6  & ~n241;
  assign n375 = ~n373 & ~n374;
  assign n376 = n208 & ~n345;
  assign n377 = ~n375 & n376;
  assign n378 = ~n371 & ~n377;
  assign n379 = ~pi1  & ~n378;
  assign n380 = ~pi2  & ~n337;
  assign n381 = ~pi6  & ~n349;
  assign n382 = ~n87 & ~n358;
  assign n383 = n381 & ~n382;
  assign n384 = ~n380 & ~n383;
  assign n385 = pi3  & ~n384;
  assign n386 = ~n336 & ~n385;
  assign n387 = ~n379 & n386;
  assign n388 = ~n356 & n387;
  assign n389 = ~n368 & n388;
  assign n390 = ~pi4  & ~n389;
  assign n391 = pi3  & ~pi9 ;
  assign n392 = pi6  & ~n52;
  assign n393 = ~n391 & ~n392;
  assign n394 = ~pi4  & ~n393;
  assign n395 = ~pi2  & n289;
  assign n396 = n375 & n395;
  assign n397 = ~n394 & ~n396;
  assign n398 = n34 & ~n397;
  assign n399 = ~n390 & ~n398;
  assign po3  = ~pi7  & ~n399;
  assign n401 = ~pi4  & n147;
  assign n402 = pi3  & ~pi4 ;
  assign n403 = ~n289 & ~n402;
  assign n404 = n91 & ~n403;
  assign n405 = ~n401 & ~n404;
  assign n406 = ~pi7  & n116;
  assign po4  = ~n405 & n406;
  assign n408 = ~n91 & n402;
  assign n409 = n34 & n395;
  assign n410 = ~n408 & ~n409;
  assign po5  = n406 & ~n410;
  assign n412 = ~n116 & ~n409;
  assign n413 = ~pi7  & ~n412;
  assign n414 = pi7  & ~pi9 ;
  assign n415 = pi8  & ~n414;
  assign n416 = n108 & ~n415;
  assign n417 = ~n78 & ~n416;
  assign n418 = ~pi0  & ~n417;
  assign n419 = ~pi2  & pi7 ;
  assign n420 = ~n276 & n419;
  assign n421 = ~n243 & n420;
  assign n422 = ~n418 & ~n421;
  assign n423 = n372 & ~n422;
  assign n424 = ~pi0  & pi2 ;
  assign n425 = pi9  & n424;
  assign n426 = ~pi9  & n195;
  assign n427 = ~n425 & ~n426;
  assign n428 = pi5  & ~n427;
  assign n429 = ~pi1  & ~pi5 ;
  assign n430 = pi2  & ~n429;
  assign n431 = n137 & ~n430;
  assign n432 = pi5  & n87;
  assign n433 = ~n431 & ~n432;
  assign n434 = pi0  & ~n433;
  assign n435 = ~n28 & n424;
  assign n436 = ~n434 & ~n435;
  assign n437 = pi8  & ~n436;
  assign n438 = pi6  & ~n297;
  assign n439 = pi2  & pi8 ;
  assign n440 = ~n187 & ~n439;
  assign n441 = n438 & ~n440;
  assign n442 = ~n428 & ~n441;
  assign n443 = ~n437 & n442;
  assign n444 = ~pi7  & ~n443;
  assign n445 = ~n423 & ~n444;
  assign n446 = ~pi3  & ~n445;
  assign n447 = n40 & n439;
  assign n448 = pi8  & ~n183;
  assign n449 = ~pi0  & ~pi6 ;
  assign n450 = n303 & ~n449;
  assign n451 = ~n448 & n450;
  assign n452 = ~n447 & ~n451;
  assign n453 = ~pi1  & ~n452;
  assign n454 = n40 & ~n218;
  assign n455 = ~n61 & ~n454;
  assign n456 = ~pi8  & ~n455;
  assign n457 = pi2  & ~n240;
  assign n458 = ~n242 & ~n457;
  assign n459 = pi6  & ~n458;
  assign n460 = ~n456 & ~n459;
  assign n461 = pi1  & ~n460;
  assign n462 = ~pi1  & ~n240;
  assign n463 = n58 & ~n462;
  assign n464 = ~n195 & n449;
  assign n465 = ~n160 & ~n464;
  assign n466 = n88 & ~n465;
  assign n467 = ~n463 & ~n466;
  assign n468 = ~pi5  & ~n467;
  assign n469 = n93 & ~n424;
  assign n470 = pi0  & n209;
  assign n471 = ~pi2  & n470;
  assign n472 = ~n469 & ~n471;
  assign n473 = pi9  & ~n472;
  assign n474 = ~pi0  & ~pi8 ;
  assign n475 = n47 & ~n183;
  assign n476 = ~n474 & n475;
  assign n477 = ~n473 & ~n476;
  assign n478 = ~n468 & n477;
  assign n479 = pi3  & ~n478;
  assign n480 = ~n453 & ~n461;
  assign n481 = ~n479 & n480;
  assign n482 = ~pi7  & ~n481;
  assign n483 = ~n446 & ~n482;
  assign n484 = ~pi4  & ~n483;
  assign po6  = ~n413 & ~n484;
  assign n486 = n98 & n199;
  assign n487 = ~n254 & ~n486;
  assign n488 = pi9  & ~n487;
  assign n489 = ~pi6  & ~n85;
  assign n490 = ~n80 & n489;
  assign n491 = ~n488 & n490;
  assign n492 = pi8  & n255;
  assign n493 = ~n491 & ~n492;
  assign n494 = pi2  & ~n493;
  assign n495 = ~pi3  & pi8 ;
  assign n496 = ~n207 & ~n495;
  assign n497 = pi0  & ~n496;
  assign n498 = ~pi9  & n209;
  assign n499 = ~n497 & ~n498;
  assign n500 = ~n488 & n499;
  assign n501 = ~pi2  & ~n500;
  assign n502 = n85 & n137;
  assign n503 = ~n501 & ~n502;
  assign n504 = ~n494 & n503;
  assign n505 = pi1  & ~n504;
  assign n506 = ~pi0  & n438;
  assign n507 = n71 & n374;
  assign n508 = ~n506 & ~n507;
  assign n509 = pi3  & ~n508;
  assign n510 = ~pi0  & n187;
  assign n511 = ~n470 & ~n510;
  assign n512 = ~pi9  & ~n511;
  assign n513 = n457 & ~n489;
  assign n514 = ~n512 & ~n513;
  assign n515 = ~n509 & n514;
  assign n516 = ~pi1  & ~n515;
  assign n517 = n348 & n441;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n505 & n518;
  assign n520 = ~pi5  & ~n519;
  assign n521 = ~pi9  & n181;
  assign n522 = pi0  & ~n77;
  assign n523 = ~n303 & n522;
  assign n524 = ~n521 & ~n523;
  assign n525 = pi8  & ~n524;
  assign n526 = n77 & n161;
  assign n527 = ~n525 & ~n526;
  assign n528 = ~pi3  & ~n527;
  assign n529 = pi3  & pi5 ;
  assign n530 = ~n33 & ~n529;
  assign n531 = ~pi0  & ~n530;
  assign n532 = pi3  & n60;
  assign n533 = ~n531 & ~n532;
  assign n534 = ~pi8  & ~n533;
  assign n535 = n303 & n529;
  assign n536 = ~n534 & ~n535;
  assign n537 = ~n528 & n536;
  assign n538 = pi1  & ~n537;
  assign n539 = n54 & n319;
  assign n540 = ~n112 & ~n297;
  assign n541 = ~n99 & ~n540;
  assign n542 = n170 & ~n541;
  assign n543 = ~n539 & ~n542;
  assign n544 = ~pi1  & ~n543;
  assign n545 = pi8  & n349;
  assign n546 = n99 & n545;
  assign n547 = ~n544 & ~n546;
  assign n548 = ~n538 & n547;
  assign n549 = ~pi6  & ~n548;
  assign n550 = ~n520 & ~n549;
  assign n551 = ~pi7  & ~n550;
  assign n552 = ~pi0  & ~n440;
  assign n553 = ~n182 & ~n552;
  assign n554 = ~pi9  & ~n553;
  assign n555 = ~pi8  & n425;
  assign n556 = ~n554 & ~n555;
  assign n557 = ~pi2  & ~n22;
  assign n558 = n130 & n372;
  assign n559 = ~n557 & n558;
  assign n560 = ~n556 & n559;
  assign n561 = ~n551 & ~n560;
  assign n562 = ~pi4  & ~n561;
  assign n563 = ~pi5  & ~pi7 ;
  assign n564 = n409 & n563;
  assign n565 = ~pi6  & n564;
  assign po7  = ~n562 & ~n565;
  assign n567 = n130 & n183;
  assign n568 = ~n165 & ~n346;
  assign n569 = ~pi2  & ~n80;
  assign n570 = n568 & n569;
  assign n571 = ~n567 & ~n570;
  assign n572 = pi8  & ~n571;
  assign n573 = pi2  & ~n183;
  assign n574 = n263 & n573;
  assign n575 = ~n572 & ~n574;
  assign n576 = ~pi9  & ~n575;
  assign n577 = ~n217 & ~n529;
  assign n578 = pi1  & ~n258;
  assign n579 = ~n577 & n578;
  assign n580 = n90 & ~n181;
  assign n581 = n196 & n580;
  assign n582 = ~n579 & ~n581;
  assign n583 = pi9  & ~n582;
  assign n584 = n88 & ~n429;
  assign n585 = n94 & ~n584;
  assign n586 = ~n256 & ~n338;
  assign n587 = ~pi0  & ~n586;
  assign n588 = ~pi2  & ~n86;
  assign n589 = ~n255 & n588;
  assign n590 = n568 & n589;
  assign n591 = ~n585 & ~n587;
  assign n592 = ~n590 & n591;
  assign n593 = ~pi8  & ~n592;
  assign n594 = ~n583 & ~n593;
  assign n595 = ~n576 & n594;
  assign n596 = ~pi6  & ~n595;
  assign n597 = ~pi8  & ~n46;
  assign n598 = ~pi6  & ~n148;
  assign n599 = ~n597 & n598;
  assign n600 = ~n47 & n199;
  assign n601 = n310 & ~n600;
  assign n602 = ~pi2  & ~n601;
  assign n603 = n346 & ~n599;
  assign n604 = ~n602 & n603;
  assign n605 = ~n596 & ~n604;
  assign n606 = ~pi7  & ~n605;
  assign n607 = ~pi1  & ~n556;
  assign n608 = n87 & n510;
  assign n609 = ~n607 & ~n608;
  assign n610 = n157 & ~n609;
  assign n611 = ~n606 & ~n610;
  assign n612 = ~pi4  & ~n611;
  assign po8  = ~n564 & ~n612;
  assign n614 = ~pi2  & n130;
  assign n615 = pi4  & ~n614;
  assign n616 = ~pi3  & ~n28;
  assign n617 = n199 & ~n496;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~pi2  & ~n618;
  assign n620 = ~pi6  & ~n545;
  assign n621 = ~pi3  & ~n620;
  assign n622 = ~pi5  & ~n241;
  assign n623 = n369 & n622;
  assign n624 = ~n621 & ~n623;
  assign n625 = ~n619 & n624;
  assign n626 = pi1  & ~n625;
  assign n627 = n289 & ~n372;
  assign n628 = n199 & ~n381;
  assign n629 = pi3  & ~n207;
  assign n630 = ~n628 & n629;
  assign n631 = ~pi2  & ~n627;
  assign n632 = ~n630 & n631;
  assign n633 = n457 & n616;
  assign n634 = ~n262 & n633;
  assign n635 = ~n632 & ~n634;
  assign n636 = ~pi1  & ~n635;
  assign n637 = n183 & n369;
  assign n638 = ~pi7  & ~n637;
  assign n639 = ~n462 & ~n638;
  assign n640 = pi7  & ~n94;
  assign n641 = ~pi7  & ~n614;
  assign n642 = pi0  & ~n641;
  assign n643 = ~pi5  & ~n94;
  assign n644 = pi6  & ~n643;
  assign n645 = ~n615 & ~n640;
  assign n646 = ~n644 & n645;
  assign n647 = ~n642 & n646;
  assign n648 = ~n639 & n647;
  assign n649 = ~n626 & n648;
  assign po9  = ~n636 & n649;
  assign n651 = ~n41 & ~n597;
  assign n652 = pi2  & n402;
  assign n653 = ~n651 & n652;
  assign n654 = ~n409 & ~n653;
  assign n655 = ~pi7  & n372;
  assign po10  = ~n654 & n655;
endmodule
