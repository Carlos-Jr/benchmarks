module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237,
    n238, n239, n240, n241, n242, n243, n244,
    n245, n246, n247, n248, n249, n250, n251,
    n252, n253, n254, n255, n256, n257, n258,
    n259, n260, n261, n262, n263, n264, n265,
    n266, n267, n268, n269, n270, n271, n272,
    n273, n274, n275, n276, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n300,
    n301, n302, n303, n304, n305, n306, n307,
    n308, n309, n310, n311, n312, n313, n314,
    n315, n316, n317, n318, n319, n320, n321,
    n322, n323, n324, n325, n326, n327, n328,
    n329, n330, n331, n332, n333, n334, n335,
    n336, n337, n338, n339, n340, n341, n342,
    n343, n344, n345, n346, n347, n348, n349,
    n350, n351, n352, n353, n354, n355, n356,
    n357, n358, n359, n360, n361, n362, n363,
    n364, n365, n366, n367, n368, n369, n370,
    n371, n372, n373, n374, n375, n376, n377,
    n378, n379, n380, n381, n382, n383, n384,
    n385, n386, n387, n388, n389, n390, n391,
    n392, n393, n394, n395, n396, n397, n398,
    n399, n400, n401, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n423, n424, n425, n426,
    n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440,
    n441, n442, n443, n444, n445, n446, n447,
    n448, n449, n450, n451, n452, n453, n454,
    n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468,
    n469, n470, n471, n472, n473, n474, n475,
    n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n546,
    n547, n548, n549, n550, n551, n552, n553,
    n554, n555, n556, n557, n558, n559, n560,
    n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574,
    n575;
  assign n91 = 1'b1;
  assign n92 = ~pi9  & ~pi10 ;
  assign n93 = pi11  & ~n92;
  assign n94 = ~pi12  & ~pi13 ;
  assign n95 = ~pi12  & ~n93;
  assign n96 = ~pi13  & n95;
  assign n97 = ~n93 & n94;
  assign n98 = pi14  & ~n556;
  assign n99 = pi15  & n98;
  assign n100 = ~pi16  & ~n99;
  assign n101 = pi17  & ~n100;
  assign n102 = ~pi18  & ~n101;
  assign n103 = pi19  & ~n102;
  assign n104 = pi20  & n103;
  assign n105 = ~pi21  & ~n104;
  assign n106 = ~pi22  & n105;
  assign n107 = pi23  & ~n106;
  assign n108 = pi24  & pi25 ;
  assign n109 = pi24  & n107;
  assign n110 = pi25  & n109;
  assign n111 = n107 & n108;
  assign n112 = ~pi26  & ~n557;
  assign n113 = pi28  & pi29 ;
  assign n114 = pi27  & n113;
  assign n115 = pi27  & ~n112;
  assign n116 = pi28  & n115;
  assign n117 = pi29  & n116;
  assign n118 = ~n112 & n114;
  assign n119 = pi26  & n557;
  assign n120 = pi22  & ~n105;
  assign n121 = pi18  & n101;
  assign n122 = ~pi17  & n100;
  assign n123 = ~n101 & ~n122;
  assign n124 = ~pi14  & n556;
  assign n125 = ~pi15  & n124;
  assign n126 = pi16  & ~n125;
  assign n127 = ~pi3  & ~pi4 ;
  assign n128 = ~pi5  & ~pi6 ;
  assign n129 = n127 & n128;
  assign n130 = ~pi1  & ~pi2 ;
  assign n131 = n94 & n130;
  assign n132 = n129 & n131;
  assign n133 = pi20  & ~pi21 ;
  assign n134 = ~pi20  & pi21 ;
  assign n135 = ~n133 & ~n134;
  assign n136 = pi11  & pi20 ;
  assign n137 = n108 & n136;
  assign n138 = ~pi7  & ~pi8 ;
  assign n139 = pi9  & ~pi10 ;
  assign n140 = n138 & n139;
  assign n141 = n137 & n140;
  assign n142 = ~n135 & n141;
  assign n143 = n132 & n142;
  assign n144 = ~n100 & n143;
  assign n145 = ~n126 & n144;
  assign n146 = ~n123 & n145;
  assign n147 = ~n121 & n146;
  assign n148 = n103 & n147;
  assign n149 = ~n120 & n148;
  assign n150 = pi25  & ~n109;
  assign n151 = ~pi25  & n109;
  assign n152 = ~n150 & ~n151;
  assign n153 = pi24  & ~n107;
  assign n154 = ~pi24  & n107;
  assign n155 = ~n153 & ~n154;
  assign n156 = ~pi23  & n106;
  assign n157 = ~n107 & ~n156;
  assign n158 = ~n106 & ~n120;
  assign n159 = pi21  & n104;
  assign n160 = ~n105 & ~n159;
  assign n161 = pi20  & ~n103;
  assign n162 = ~pi20  & n103;
  assign n163 = ~n161 & ~n162;
  assign n164 = ~pi19  & n102;
  assign n165 = ~n103 & ~n164;
  assign n166 = ~n102 & ~n121;
  assign n167 = pi16  & n99;
  assign n168 = ~n100 & ~n167;
  assign n169 = pi15  & ~n98;
  assign n170 = ~pi15  & n98;
  assign n171 = ~n169 & ~n170;
  assign n172 = ~n98 & ~n124;
  assign n173 = pi13  & ~n95;
  assign n174 = ~n556 & ~n173;
  assign n175 = pi12  & n93;
  assign n176 = ~n95 & ~n175;
  assign n177 = ~pi11  & n92;
  assign n178 = ~n93 & ~n177;
  assign n179 = ~pi3  & n130;
  assign n180 = ~pi4  & n179;
  assign n181 = ~pi5  & n180;
  assign n182 = ~pi6  & n181;
  assign n183 = n129 & n130;
  assign n184 = n140 & n559;
  assign n185 = ~n178 & n184;
  assign n186 = n176 & n185;
  assign n187 = n174 & n186;
  assign n188 = ~n172 & n187;
  assign n189 = n171 & n188;
  assign n190 = n168 & n189;
  assign n191 = ~n123 & n190;
  assign n192 = n166 & n191;
  assign n193 = ~n165 & n192;
  assign n194 = n163 & n193;
  assign n195 = n160 & n194;
  assign n196 = n158 & n195;
  assign n197 = ~n157 & n196;
  assign n198 = n155 & n197;
  assign n199 = n152 & n198;
  assign n200 = n107 & n149;
  assign n201 = ~n112 & ~n119;
  assign n202 = n560 & n201;
  assign n203 = ~n119 & n560;
  assign n204 = pi28  & ~n115;
  assign n205 = ~pi28  & n115;
  assign n206 = ~n204 & ~n205;
  assign n207 = ~pi27  & n112;
  assign n208 = ~n115 & ~n207;
  assign n209 = pi9  & pi10 ;
  assign n210 = ~n92 & ~n209;
  assign n211 = ~pi7  & n559;
  assign n212 = ~pi8  & n211;
  assign n213 = n210 & n212;
  assign n214 = ~n178 & n213;
  assign n215 = n176 & n214;
  assign n216 = n174 & n215;
  assign n217 = ~n172 & n216;
  assign n218 = n171 & n217;
  assign n219 = n168 & n218;
  assign n220 = ~n123 & n219;
  assign n221 = n166 & n220;
  assign n222 = ~n165 & n221;
  assign n223 = n163 & n222;
  assign n224 = n160 & n223;
  assign n225 = n158 & n224;
  assign n226 = ~n157 & n225;
  assign n227 = n155 & n226;
  assign n228 = n152 & n227;
  assign n229 = n201 & n228;
  assign n230 = ~n208 & n229;
  assign n231 = n206 & n230;
  assign n232 = pi9  & n231;
  assign n233 = n558 & ~n232;
  assign n234 = n561 & ~n208;
  assign n235 = n558 & ~n234;
  assign n236 = n558 & ~n561;
  assign n237 = ~pi39  & ~pi40 ;
  assign n238 = pi41  & ~n237;
  assign n239 = ~pi42  & ~n238;
  assign n240 = ~pi43  & n239;
  assign n241 = pi44  & ~n240;
  assign n242 = pi45  & n241;
  assign n243 = ~pi46  & ~n242;
  assign n244 = pi47  & ~n243;
  assign n245 = ~pi48  & ~n244;
  assign n246 = pi49  & ~n245;
  assign n247 = pi50  & n246;
  assign n248 = ~pi51  & ~n247;
  assign n249 = ~pi52  & n248;
  assign n250 = pi53  & ~n249;
  assign n251 = pi54  & n250;
  assign n252 = pi55  & n251;
  assign n253 = ~pi56  & ~n252;
  assign n254 = pi57  & ~n253;
  assign n255 = pi58  & pi59 ;
  assign n256 = pi58  & n254;
  assign n257 = pi59  & n256;
  assign n258 = n254 & n255;
  assign n259 = ~pi57  & n253;
  assign n260 = ~n254 & ~n259;
  assign n261 = pi56  & n252;
  assign n262 = ~n253 & ~n261;
  assign n263 = ~pi55  & ~n251;
  assign n264 = pi55  & ~n251;
  assign n265 = ~pi55  & n251;
  assign n266 = ~n264 & ~n265;
  assign n267 = ~n252 & ~n263;
  assign n268 = ~pi54  & ~n250;
  assign n269 = pi54  & ~n250;
  assign n270 = ~pi54  & n250;
  assign n271 = ~n269 & ~n270;
  assign n272 = ~n251 & ~n268;
  assign n273 = ~pi53  & n249;
  assign n274 = ~n250 & ~n273;
  assign n275 = pi43  & ~n239;
  assign n276 = ~pi31  & ~pi32 ;
  assign n277 = ~pi33  & ~pi34 ;
  assign n278 = ~pi35  & ~pi36 ;
  assign n279 = n277 & n278;
  assign n280 = ~pi33  & n276;
  assign n281 = ~pi34  & n280;
  assign n282 = ~pi35  & n281;
  assign n283 = ~pi36  & n282;
  assign n284 = n276 & n279;
  assign n285 = pi47  & ~pi48 ;
  assign n286 = pi49  & n285;
  assign n287 = pi41  & ~pi42 ;
  assign n288 = pi45  & ~pi46 ;
  assign n289 = n287 & n288;
  assign n290 = ~pi37  & ~pi38 ;
  assign n291 = pi39  & ~pi40 ;
  assign n292 = n290 & n291;
  assign n293 = n289 & n292;
  assign n294 = n286 & n293;
  assign n295 = n566 & n294;
  assign n296 = ~n275 & n295;
  assign n297 = ~pi49  & n245;
  assign n298 = ~n246 & ~n297;
  assign n299 = pi48  & n244;
  assign n300 = ~n245 & ~n299;
  assign n301 = ~pi47  & n243;
  assign n302 = ~n244 & ~n301;
  assign n303 = pi46  & n242;
  assign n304 = ~n243 & ~n303;
  assign n305 = pi45  & ~n241;
  assign n306 = ~pi45  & n241;
  assign n307 = ~n305 & ~n306;
  assign n308 = ~pi44  & n240;
  assign n309 = ~n241 & ~n308;
  assign n310 = ~n240 & ~n275;
  assign n311 = pi42  & n238;
  assign n312 = ~n239 & ~n311;
  assign n313 = ~pi41  & n237;
  assign n314 = ~n238 & ~n313;
  assign n315 = n566 & n292;
  assign n316 = ~n314 & n315;
  assign n317 = n312 & n316;
  assign n318 = n310 & n317;
  assign n319 = ~n309 & n318;
  assign n320 = n307 & n319;
  assign n321 = n304 & n320;
  assign n322 = ~n302 & n321;
  assign n323 = n300 & n322;
  assign n324 = ~n298 & n323;
  assign n325 = n241 & n296;
  assign n326 = ~n248 & n567;
  assign n327 = pi51  & n247;
  assign n328 = ~pi50  & ~n246;
  assign n329 = pi50  & ~n246;
  assign n330 = ~pi50  & n246;
  assign n331 = ~n329 & ~n330;
  assign n332 = ~n247 & ~n328;
  assign n333 = ~n327 & n568;
  assign n334 = ~n248 & ~n327;
  assign n335 = n567 & n568;
  assign n336 = n334 & n335;
  assign n337 = n326 & n333;
  assign n338 = pi52  & ~n248;
  assign n339 = ~n249 & ~n338;
  assign n340 = n569 & n339;
  assign n341 = ~n274 & n340;
  assign n342 = n565 & n341;
  assign n343 = n564 & n342;
  assign n344 = n262 & n343;
  assign n345 = ~n260 & n344;
  assign n346 = ~pi0  & ~pi30 ;
  assign n347 = n345 & n346;
  assign n348 = n563 & ~n347;
  assign n349 = pi47  & ~n241;
  assign n350 = ~pi47  & n241;
  assign n351 = ~n349 & ~n350;
  assign n352 = pi32  & pi33 ;
  assign n353 = pi34  & pi35 ;
  assign n354 = n352 & n353;
  assign n355 = pi30  & pi31 ;
  assign n356 = n237 & n355;
  assign n357 = n354 & n356;
  assign n358 = ~pi42  & ~pi43 ;
  assign n359 = pi44  & pi45 ;
  assign n360 = n358 & n359;
  assign n361 = pi36  & pi37 ;
  assign n362 = pi38  & pi41 ;
  assign n363 = n361 & n362;
  assign n364 = n360 & n363;
  assign n365 = ~pi52  & pi53 ;
  assign n366 = n255 & n365;
  assign n367 = ~pi46  & ~pi48 ;
  assign n368 = pi49  & ~pi51 ;
  assign n369 = n367 & n368;
  assign n370 = n366 & n369;
  assign n371 = n364 & n370;
  assign n372 = n357 & n371;
  assign n373 = ~n351 & n372;
  assign n374 = n352 & n355;
  assign n375 = n237 & n374;
  assign n376 = pi38  & pi58 ;
  assign n377 = pi59  & n376;
  assign n378 = n353 & n361;
  assign n379 = n377 & n378;
  assign n380 = n375 & n379;
  assign n381 = n314 & n380;
  assign n382 = ~n312 & n381;
  assign n383 = ~n310 & n382;
  assign n384 = n309 & n383;
  assign n385 = ~n307 & n384;
  assign n386 = ~n304 & n385;
  assign n387 = n302 & n386;
  assign n388 = ~n300 & n387;
  assign n389 = n298 & n388;
  assign n390 = ~n568 & n389;
  assign n391 = ~n334 & n390;
  assign n392 = ~n339 & n391;
  assign n393 = n274 & n392;
  assign n394 = ~n568 & n373;
  assign n395 = ~n565 & n570;
  assign n396 = ~n564 & n395;
  assign n397 = ~n262 & n396;
  assign n398 = pi39  & pi40 ;
  assign n399 = ~n237 & ~n398;
  assign n400 = pi58  & ~n254;
  assign n401 = ~pi58  & n254;
  assign n402 = ~n400 & ~n401;
  assign n403 = pi30  & ~pi39 ;
  assign n404 = pi59  & n403;
  assign n405 = ~n402 & n404;
  assign n406 = n260 & n405;
  assign n407 = ~n262 & n406;
  assign n408 = ~n564 & n407;
  assign n409 = ~n565 & n408;
  assign n410 = n274 & n409;
  assign n411 = ~n339 & n410;
  assign n412 = ~n334 & n411;
  assign n413 = ~n568 & n412;
  assign n414 = n298 & n413;
  assign n415 = ~n300 & n414;
  assign n416 = n302 & n415;
  assign n417 = ~n304 & n416;
  assign n418 = ~n307 & n417;
  assign n419 = n309 & n418;
  assign n420 = ~n310 & n419;
  assign n421 = ~n312 & n420;
  assign n422 = n314 & n421;
  assign n423 = ~n399 & n422;
  assign n424 = pi38  & n423;
  assign n425 = pi37  & n424;
  assign n426 = pi36  & n425;
  assign n427 = pi35  & n426;
  assign n428 = pi34  & n427;
  assign n429 = pi33  & n428;
  assign n430 = pi32  & n429;
  assign n431 = pi31  & n430;
  assign n432 = n260 & n397;
  assign n433 = n563 & ~n346;
  assign n434 = ~pi37  & n566;
  assign n435 = ~pi38  & n434;
  assign n436 = n399 & n435;
  assign n437 = ~n314 & n436;
  assign n438 = n312 & n437;
  assign n439 = n310 & n438;
  assign n440 = ~n309 & n439;
  assign n441 = n307 & n440;
  assign n442 = n304 & n441;
  assign n443 = ~n302 & n442;
  assign n444 = n300 & n443;
  assign n445 = ~n298 & n444;
  assign n446 = n568 & n445;
  assign n447 = n334 & n446;
  assign n448 = n339 & n447;
  assign n449 = ~n274 & n448;
  assign n450 = n565 & n449;
  assign n451 = n564 & n450;
  assign n452 = n262 & n451;
  assign n453 = ~n260 & n452;
  assign n454 = n402 & n453;
  assign n455 = pi39  & n454;
  assign n456 = n563 & ~n455;
  assign n457 = ~n571 & ~n456;
  assign n458 = ~n433 & n457;
  assign n459 = ~n348 & ~n571;
  assign n460 = ~pi23  & ~n120;
  assign n461 = ~pi12  & pi15 ;
  assign n462 = pi17  & ~pi18 ;
  assign n463 = n461 & n462;
  assign n464 = pi6  & pi7 ;
  assign n465 = pi8  & pi11 ;
  assign n466 = n464 & n465;
  assign n467 = n463 & n466;
  assign n468 = n114 & n467;
  assign n469 = pi19  & ~pi26 ;
  assign n470 = n108 & n469;
  assign n471 = n133 & n470;
  assign n472 = pi2  & pi3 ;
  assign n473 = pi4  & pi5 ;
  assign n474 = n472 & n473;
  assign n475 = pi0  & pi1 ;
  assign n476 = n92 & n475;
  assign n477 = n474 & n476;
  assign n478 = n471 & n477;
  assign n479 = n468 & n478;
  assign n480 = n172 & n479;
  assign n481 = ~n174 & n480;
  assign n482 = n100 & n481;
  assign n483 = ~n107 & n482;
  assign n484 = ~pi29  & n116;
  assign n485 = pi29  & ~n116;
  assign n486 = ~n484 & ~n485;
  assign n487 = ~pi9  & ~n486;
  assign n488 = ~n206 & n487;
  assign n489 = n208 & n488;
  assign n490 = ~n201 & n489;
  assign n491 = ~n152 & n490;
  assign n492 = ~n155 & n491;
  assign n493 = n157 & n492;
  assign n494 = ~n158 & n493;
  assign n495 = ~n160 & n494;
  assign n496 = ~n163 & n495;
  assign n497 = n165 & n496;
  assign n498 = ~n166 & n497;
  assign n499 = n123 & n498;
  assign n500 = ~n168 & n499;
  assign n501 = ~n171 & n500;
  assign n502 = n172 & n501;
  assign n503 = ~n174 & n502;
  assign n504 = ~n176 & n503;
  assign n505 = n178 & n504;
  assign n506 = ~n210 & n505;
  assign n507 = pi8  & n506;
  assign n508 = pi7  & n507;
  assign n509 = pi6  & n508;
  assign n510 = pi5  & n509;
  assign n511 = pi4  & n510;
  assign n512 = pi3  & n511;
  assign n513 = pi2  & n512;
  assign n514 = pi1  & n513;
  assign n515 = pi0  & n514;
  assign n516 = pi8  & pi29 ;
  assign n517 = n464 & n516;
  assign n518 = n477 & n517;
  assign n519 = n178 & n518;
  assign n520 = ~n176 & n519;
  assign n521 = ~n174 & n520;
  assign n522 = n172 & n521;
  assign n523 = ~n171 & n522;
  assign n524 = ~n168 & n523;
  assign n525 = n123 & n524;
  assign n526 = ~n166 & n525;
  assign n527 = n165 & n526;
  assign n528 = ~n163 & n527;
  assign n529 = ~n160 & n528;
  assign n530 = ~n158 & n529;
  assign n531 = n157 & n530;
  assign n532 = ~n155 & n531;
  assign n533 = ~n152 & n532;
  assign n534 = ~n201 & n533;
  assign n535 = ~pi28  & ~n115;
  assign n536 = n208 & ~n535;
  assign n537 = n534 & n536;
  assign n538 = ~n460 & n483;
  assign n539 = ~n558 & ~n573;
  assign n540 = pi0  & ~n563;
  assign n541 = ~n539 & ~n540;
  assign n542 = ~n572 & ~n539;
  assign n543 = ~n540 & n542;
  assign n544 = ~n572 & n541;
  assign po1  = ~n562 & ~n574;
  assign n546 = pi0  & pi30 ;
  assign n547 = n345 & ~n546;
  assign n548 = ~n562 & ~n539;
  assign n549 = n563 & n548;
  assign n550 = pi0  & n563;
  assign n551 = pi30  & n550;
  assign n552 = ~n456 & ~n551;
  assign n553 = n563 & ~n547;
  assign n554 = n548 & ~n575;
  assign n555 = ~n547 & n549;
  assign n556 = n96 | n97;
  assign n557 = n110 | n111;
  assign n558 = n117 | n118;
  assign n559 = n182 | n183;
  assign n560 = n199 | n200;
  assign n561 = n202 | n203;
  assign n562 = n236 | n233 | n235;
  assign n563 = n257 | n258;
  assign n564 = n266 | ~n267;
  assign n565 = n271 | ~n272;
  assign n566 = n283 | n284;
  assign n567 = n324 | n325;
  assign n568 = n331 | ~n332;
  assign n569 = n336 | n337;
  assign n570 = n393 | n394;
  assign n571 = n431 | n432;
  assign n572 = n458 | n459;
  assign n573 = n538 | n515 | n537;
  assign n574 = n543 | n544;
  assign n575 = n552 | ~n553;
  assign po2  = n554 | n555;
  assign po0  = ~n548;
  assign po3  = ~n91;
  assign po4  = ~n91;
  assign po5  = ~n91;
  assign po6  = ~n91;
  assign po7  = ~n91;
  assign po8  = ~n91;
  assign po9  = ~n91;
  assign po10  = ~n91;
  assign po11  = ~n91;
  assign po12  = ~n91;
  assign po13  = ~n91;
  assign po14  = ~n91;
  assign po15  = ~n91;
  assign po16  = ~n91;
  assign po17  = ~n91;
  assign po18  = ~n91;
  assign po19  = ~n91;
  assign po20  = ~n91;
  assign po21  = ~n91;
  assign po22  = ~n91;
  assign po23  = ~n91;
  assign po24  = ~n91;
  assign po25  = ~n91;
  assign po26  = ~n91;
  assign po27  = ~n91;
  assign po28  = ~n91;
  assign po29  = ~n91;
endmodule
