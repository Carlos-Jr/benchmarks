module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n175, n176,
    n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n264, n265, n267, n268,
    n269;
  assign n92 = pi28  & pi29 ;
  assign n93 = pi14  & pi15 ;
  assign n94 = ~pi9  & ~pi10 ;
  assign n95 = pi11  & ~n94;
  assign n96 = ~pi12  & ~pi13 ;
  assign n97 = ~n95 & n96;
  assign n98 = n93 & ~n97;
  assign n99 = ~pi16  & ~n98;
  assign n100 = pi17  & ~n99;
  assign n101 = ~pi18  & ~n100;
  assign n102 = pi19  & pi20 ;
  assign n103 = ~n101 & n102;
  assign n104 = ~pi21  & ~n103;
  assign n105 = ~pi22  & n104;
  assign n106 = pi23  & ~n105;
  assign n107 = pi24  & n106;
  assign n108 = pi25  & n107;
  assign n109 = ~pi26  & ~n108;
  assign n110 = pi27  & n92;
  assign n111 = ~n109 & n110;
  assign n112 = ~pi22  & pi23 ;
  assign n113 = ~pi24  & ~n106;
  assign n114 = ~pi17  & n99;
  assign n115 = pi16  & ~n98;
  assign n116 = ~pi16  & n98;
  assign n117 = ~n115 & ~n116;
  assign n118 = pi14  & ~n97;
  assign n119 = ~pi15  & ~n118;
  assign n120 = pi0  & pi1 ;
  assign n121 = pi2  & pi3 ;
  assign n122 = pi4  & pi5 ;
  assign n123 = pi6  & pi7 ;
  assign n124 = pi8  & pi11 ;
  assign n125 = pi14  & ~pi21 ;
  assign n126 = pi25  & ~pi26 ;
  assign n127 = n96 & n125;
  assign n128 = n123 & n124;
  assign n129 = n121 & n122;
  assign n130 = n120 & n126;
  assign n131 = n94 & n102;
  assign n132 = n112 & n131;
  assign n133 = n129 & n130;
  assign n134 = n127 & n128;
  assign n135 = n110 & n134;
  assign n136 = n132 & n133;
  assign n137 = n135 & n136;
  assign n138 = ~n98 & n137;
  assign n139 = ~n119 & n138;
  assign n140 = ~n114 & n117;
  assign n141 = n139 & n140;
  assign n142 = n101 & n141;
  assign n143 = ~n107 & n142;
  assign n144 = ~n113 & n143;
  assign n145 = ~n111 & ~n144;
  assign n146 = pi19  & ~n101;
  assign n147 = ~pi19  & n101;
  assign n148 = ~n146 & ~n147;
  assign n149 = ~pi20  & ~n103;
  assign n150 = ~n146 & n149;
  assign n151 = pi21  & ~n150;
  assign n152 = ~pi1  & ~pi2 ;
  assign n153 = ~pi3  & ~pi4 ;
  assign n154 = ~pi5  & ~pi6 ;
  assign n155 = ~pi7  & ~pi8 ;
  assign n156 = ~pi10  & ~pi12 ;
  assign n157 = ~pi13  & pi17 ;
  assign n158 = ~pi18  & pi24 ;
  assign n159 = n126 & n158;
  assign n160 = n156 & n157;
  assign n161 = n154 & n155;
  assign n162 = n152 & n153;
  assign n163 = n93 & n112;
  assign n164 = n162 & n163;
  assign n165 = n160 & n161;
  assign n166 = n95 & n159;
  assign n167 = n165 & n166;
  assign n168 = n164 & n167;
  assign n169 = ~n117 & n168;
  assign n170 = ~n104 & n169;
  assign n171 = ~n148 & n170;
  assign n172 = ~n151 & n171;
  assign n173 = n111 & ~n172;
  assign po0  = n145 | n173;
  assign n175 = ~pi39  & ~pi40 ;
  assign n176 = pi41  & ~n175;
  assign n177 = ~pi42  & ~n176;
  assign n178 = ~pi43  & n177;
  assign n179 = pi44  & ~n178;
  assign n180 = pi45  & n179;
  assign n181 = ~pi46  & ~n180;
  assign n182 = pi47  & ~n181;
  assign n183 = ~pi48  & ~n182;
  assign n184 = pi49  & pi50 ;
  assign n185 = ~n183 & n184;
  assign n186 = ~pi51  & ~n185;
  assign n187 = ~pi52  & n186;
  assign n188 = pi53  & ~n187;
  assign n189 = pi54  & pi55 ;
  assign n190 = n188 & n189;
  assign n191 = ~pi56  & ~n190;
  assign n192 = pi58  & pi59 ;
  assign n193 = ~n191 & n192;
  assign n194 = pi57  & n193;
  assign n195 = pi0  & ~n194;
  assign n196 = ~pi0  & ~pi30 ;
  assign n197 = n193 & ~n196;
  assign n198 = ~pi53  & n187;
  assign n199 = ~n188 & ~n198;
  assign n200 = pi52  & ~n186;
  assign n201 = ~n187 & ~n200;
  assign n202 = pi51  & n185;
  assign n203 = ~n186 & ~n202;
  assign n204 = ~pi46  & pi47 ;
  assign n205 = ~pi48  & n204;
  assign n206 = pi30  & pi31 ;
  assign n207 = pi32  & pi33 ;
  assign n208 = pi34  & pi35 ;
  assign n209 = pi36  & pi37 ;
  assign n210 = pi38  & pi41 ;
  assign n211 = pi44  & pi45 ;
  assign n212 = ~pi56  & pi58 ;
  assign n213 = pi59  & n212;
  assign n214 = n210 & n211;
  assign n215 = n208 & n209;
  assign n216 = n206 & n207;
  assign n217 = n184 & n189;
  assign n218 = n216 & n217;
  assign n219 = n214 & n215;
  assign n220 = n205 & n213;
  assign n221 = n219 & n220;
  assign n222 = n218 & n221;
  assign n223 = n178 & n222;
  assign n224 = ~n203 & n223;
  assign n225 = ~n201 & n224;
  assign n226 = n199 & n225;
  assign n227 = pi54  & n188;
  assign n228 = ~pi55  & ~n190;
  assign n229 = ~n227 & n228;
  assign n230 = pi56  & ~n229;
  assign n231 = pi49  & ~n183;
  assign n232 = ~pi50  & ~n231;
  assign n233 = ~n185 & ~n232;
  assign n234 = ~pi54  & ~n188;
  assign n235 = ~n227 & ~n234;
  assign n236 = pi43  & ~n177;
  assign n237 = ~pi31  & ~pi32 ;
  assign n238 = ~pi33  & ~pi34 ;
  assign n239 = ~pi35  & ~pi36 ;
  assign n240 = ~pi37  & ~pi38 ;
  assign n241 = pi39  & ~pi40 ;
  assign n242 = pi41  & ~pi42 ;
  assign n243 = pi45  & pi49 ;
  assign n244 = n242 & n243;
  assign n245 = n240 & n241;
  assign n246 = n238 & n239;
  assign n247 = n237 & n246;
  assign n248 = n244 & n245;
  assign n249 = n205 & n248;
  assign n250 = n247 & n249;
  assign n251 = ~n236 & n250;
  assign n252 = n179 & n251;
  assign n253 = n203 & n252;
  assign n254 = ~n233 & n253;
  assign n255 = n201 & n254;
  assign n256 = ~n199 & n255;
  assign n257 = ~n191 & ~n235;
  assign n258 = n256 & n257;
  assign n259 = ~n230 & n258;
  assign n260 = n193 & ~n259;
  assign n261 = ~n197 & ~n226;
  assign n262 = ~n260 & n261;
  assign n263 = pi57  & ~n145;
  assign n264 = ~n195 & n263;
  assign n265 = ~n262 & n264;
  assign po1  = ~n173 & ~n265;
  assign n267 = pi0  & pi30 ;
  assign n268 = n259 & ~n267;
  assign n269 = ~po0  & n194;
  assign po2  = ~n268 & n269;
  assign po3  = 1'b0;
  assign po4  = 1'b0;
  assign po5  = 1'b0;
  assign po6  = 1'b0;
  assign po7  = 1'b0;
  assign po8  = 1'b0;
  assign po9  = 1'b0;
  assign po10  = 1'b0;
  assign po11  = 1'b0;
  assign po12  = 1'b0;
  assign po13  = 1'b0;
  assign po14  = 1'b0;
  assign po15  = 1'b0;
  assign po16  = 1'b0;
  assign po17  = 1'b0;
  assign po18  = 1'b0;
  assign po19  = 1'b0;
  assign po20  = 1'b0;
  assign po21  = 1'b0;
  assign po22  = 1'b0;
  assign po23  = 1'b0;
  assign po24  = 1'b0;
  assign po25  = 1'b0;
  assign po26  = 1'b0;
  assign po27  = 1'b0;
  assign po28  = 1'b0;
  assign po29  = 1'b0;
endmodule
