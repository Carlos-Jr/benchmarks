module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ;
  wire n19, n20, n21, n22, n23, n24, n25,
    n26, n27, n28, n29, n30, n31, n32, n33,
    n34, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49,
    n50, n51, n52, n53, n54, n55, n56, n57,
    n58, n59, n60, n61, n62, n63, n64, n65,
    n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n78, n79, n80, n81,
    n82, n83, n84, n85, n86, n87, n88, n89,
    n90, n91, n92, n93, n94, n95, n96, n97,
    n98, n99, n100, n101, n102, n103, n104,
    n105, n106, n107, n108, n109, n110, n111,
    n112, n113, n114, n115, n116, n117, n118,
    n119, n120, n121, n122, n123, n124, n125,
    n126, n127, n128, n129, n130, n131, n132,
    n133, n134, n135, n136, n137, n138, n139,
    n140, n141, n142, n143, n144, n145, n146,
    n147, n148, n149, n150, n151, n152, n153,
    n154, n155, n156, n157, n158, n159, n160,
    n161, n162, n163, n164, n165, n166, n167,
    n168, n169, n170, n171, n172, n173, n174,
    n175, n176, n177, n178, n179, n180, n181,
    n182, n183, n184, n185, n186, n187, n188,
    n189, n190, n191, n192, n193, n194, n195,
    n196, n197, n198, n199, n200, n201, n202,
    n203, n204, n205, n206, n207, n208, n209,
    n210, n211, n212, n213, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n236, n237, n238,
    n239, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n276, n277, n278, n279, n280,
    n281, n282, n283, n284, n285, n286, n287,
    n288, n289, n290, n291, n292, n293, n294,
    n295, n296, n297, n298, n299, n300, n301,
    n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n329,
    n330, n331, n332, n333, n334, n335, n336,
    n337, n338, n339, n340, n341, n342, n343,
    n344, n345, n346, n347, n348, n349, n350,
    n351, n352, n353, n354, n355, n356, n357,
    n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371,
    n372, n373, n374, n375, n376, n377, n378,
    n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392,
    n393, n394, n395, n396, n397, n398, n399,
    n400, n401, n402, n403, n404, n405, n406,
    n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n433, n434,
    n435, n436, n437, n438, n439, n440, n441,
    n442, n443, n444, n445, n446, n447, n448,
    n449, n450, n451, n452, n453, n454, n455,
    n456, n457, n458, n459, n460, n461, n462,
    n463, n464, n465, n466, n467, n468, n469,
    n470, n471, n472, n473, n474, n475, n476,
    n477, n478, n479, n480, n481, n482, n483,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n492, n493, n494, n495, n496, n497,
    n498;
  assign n19 = ~pi4  & pi7 ;
  assign n20 = ~pi2  & ~pi7 ;
  assign n21 = pi1  & pi5 ;
  assign n22 = pi1  & ~pi2 ;
  assign n23 = pi5  & ~pi7 ;
  assign n24 = n22 & n23;
  assign n25 = n20 & n21;
  assign n26 = ~n19 & ~n435;
  assign n27 = pi3  & ~n26;
  assign n28 = ~pi3  & pi4 ;
  assign n29 = pi4  & pi7 ;
  assign n30 = ~pi3  & n29;
  assign n31 = pi7  & n28;
  assign n32 = ~n27 & ~n436;
  assign n33 = ~pi8  & ~n32;
  assign n34 = ~pi4  & pi8 ;
  assign n35 = pi5  & ~n34;
  assign n36 = pi1  & pi4 ;
  assign n37 = ~pi1  & pi4 ;
  assign n38 = ~pi4  & ~pi8 ;
  assign n39 = ~n37 & ~n38;
  assign n40 = ~n34 & ~n36;
  assign n41 = pi0  & n437;
  assign n42 = ~pi0  & ~n36;
  assign n43 = ~pi6  & ~pi7 ;
  assign n44 = ~n42 & n43;
  assign n45 = pi0  & ~n437;
  assign n46 = ~pi0  & pi1 ;
  assign n47 = ~pi0  & n36;
  assign n48 = pi4  & n46;
  assign n49 = ~n45 & ~n438;
  assign n50 = ~pi6  & ~n49;
  assign n51 = ~pi7  & n50;
  assign n52 = n43 & ~n49;
  assign n53 = ~n41 & n44;
  assign n54 = pi4  & pi8 ;
  assign n55 = ~pi5  & ~n54;
  assign n56 = ~n439 & n55;
  assign n57 = ~n439 & ~n54;
  assign n58 = ~pi5  & ~n57;
  assign n59 = ~pi4  & pi5 ;
  assign n60 = pi5  & pi8 ;
  assign n61 = ~pi4  & n60;
  assign n62 = pi5  & n34;
  assign n63 = pi8  & n59;
  assign n64 = ~n58 & ~n440;
  assign n65 = ~n35 & ~n56;
  assign n66 = ~n33 & ~n440;
  assign n67 = ~n58 & n66;
  assign n68 = ~n33 & n441;
  assign n69 = ~pi9  & ~n442;
  assign n70 = ~pi5  & pi6 ;
  assign n71 = pi6  & pi9 ;
  assign n72 = ~pi5  & n71;
  assign n73 = pi9  & n70;
  assign n74 = pi5  & ~pi6 ;
  assign n75 = ~n19 & n22;
  assign n76 = pi3  & pi4 ;
  assign n77 = ~n54 & ~n76;
  assign n78 = pi4  & ~pi8 ;
  assign n79 = ~pi3  & n78;
  assign n80 = ~pi4  & ~pi7 ;
  assign n81 = ~n79 & ~n80;
  assign n82 = ~pi2  & ~n81;
  assign n83 = pi1  & n82;
  assign n84 = n22 & ~n54;
  assign n85 = ~n19 & ~n76;
  assign n86 = n84 & n85;
  assign n87 = ~n19 & ~n54;
  assign n88 = n22 & ~n76;
  assign n89 = n87 & n88;
  assign n90 = n22 & ~n81;
  assign n91 = n75 & n77;
  assign n92 = ~pi7  & ~pi8 ;
  assign n93 = ~pi1  & pi2 ;
  assign n94 = n92 & n93;
  assign n95 = ~pi9  & ~n94;
  assign n96 = ~n444 & n95;
  assign n97 = ~pi6  & ~n96;
  assign n98 = pi5  & n97;
  assign n99 = n74 & ~n96;
  assign n100 = ~n443 & ~n445;
  assign n101 = ~n69 & n100;
  assign n102 = ~pi10  & ~n101;
  assign n103 = ~pi6  & pi7 ;
  assign n104 = ~pi6  & pi10 ;
  assign n105 = pi7  & n104;
  assign n106 = pi10  & n103;
  assign n107 = ~pi2  & pi3 ;
  assign n108 = pi2  & ~pi3 ;
  assign n109 = ~n107 & ~n108;
  assign n110 = ~pi8  & ~pi9 ;
  assign n111 = ~pi9  & ~n109;
  assign n112 = ~pi8  & n111;
  assign n113 = ~n109 & n110;
  assign n114 = ~pi10  & ~n447;
  assign n115 = ~pi7  & ~n114;
  assign n116 = pi8  & pi10 ;
  assign n117 = pi9  & pi10 ;
  assign n118 = pi8  & n117;
  assign n119 = pi8  & pi9 ;
  assign n120 = pi10  & n119;
  assign n121 = pi9  & n116;
  assign n122 = ~n115 & ~n448;
  assign n123 = pi6  & ~n122;
  assign n124 = ~n446 & ~n123;
  assign n125 = ~n102 & n124;
  assign n126 = pi1  & pi2 ;
  assign n127 = pi0  & ~n126;
  assign n128 = pi4  & ~pi7 ;
  assign n129 = ~pi0  & pi2 ;
  assign n130 = n128 & ~n129;
  assign n131 = pi0  & n126;
  assign n132 = ~pi0  & ~pi2 ;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~pi7  & ~n133;
  assign n135 = pi4  & n134;
  assign n136 = n128 & ~n133;
  assign n137 = ~n127 & n130;
  assign n138 = pi8  & ~pi9 ;
  assign n139 = ~pi4  & ~pi9 ;
  assign n140 = ~n20 & ~n139;
  assign n141 = ~pi1  & ~n140;
  assign n142 = ~n138 & ~n141;
  assign n143 = ~n449 & ~n138;
  assign n144 = ~n141 & n143;
  assign n145 = ~n449 & n142;
  assign n146 = ~pi6  & ~n450;
  assign n147 = ~pi7  & pi9 ;
  assign n148 = pi7  & ~n76;
  assign n149 = ~pi9  & n148;
  assign n150 = ~pi8  & n149;
  assign n151 = pi7  & ~pi8 ;
  assign n152 = ~pi9  & n151;
  assign n153 = ~n76 & n152;
  assign n154 = n110 & n148;
  assign n155 = ~n147 & ~n451;
  assign n156 = ~n146 & n155;
  assign n157 = ~pi5  & ~n156;
  assign n158 = ~pi7  & ~n126;
  assign n159 = pi3  & ~n158;
  assign n160 = pi4  & ~n110;
  assign n161 = ~pi4  & ~n43;
  assign n162 = pi4  & n110;
  assign n163 = ~pi9  & n78;
  assign n164 = ~pi4  & ~pi6 ;
  assign n165 = ~pi7  & n164;
  assign n166 = ~pi4  & n43;
  assign n167 = ~n452 & ~n453;
  assign n168 = ~n160 & ~n161;
  assign n169 = pi3  & ~n161;
  assign n170 = ~n158 & ~n160;
  assign n171 = n169 & n170;
  assign n172 = pi2  & ~n454;
  assign n173 = pi1  & n172;
  assign n174 = n126 & ~n454;
  assign n175 = pi7  & ~pi9 ;
  assign n176 = n78 & n175;
  assign n177 = ~n456 & ~n176;
  assign n178 = pi3  & ~n177;
  assign n179 = n159 & ~n454;
  assign n180 = pi6  & ~n110;
  assign n181 = ~n139 & ~n147;
  assign n182 = pi4  & n138;
  assign n183 = pi7  & pi9 ;
  assign n184 = ~n182 & ~n183;
  assign n185 = pi6  & ~n184;
  assign n186 = n180 & n181;
  assign n187 = ~n455 & ~n457;
  assign n188 = pi5  & ~n187;
  assign n189 = ~pi4  & n138;
  assign n190 = ~pi9  & n34;
  assign n191 = ~n147 & ~n458;
  assign n192 = ~pi6  & ~n191;
  assign n193 = ~n188 & ~n192;
  assign n194 = ~n157 & ~n192;
  assign n195 = ~n188 & n194;
  assign n196 = ~n157 & n193;
  assign n197 = ~pi10  & ~n459;
  assign n198 = pi6  & pi7 ;
  assign n199 = ~pi9  & n198;
  assign n200 = pi6  & pi10 ;
  assign n201 = pi7  & n200;
  assign n202 = pi10  & n198;
  assign n203 = n138 & n460;
  assign n204 = n116 & n199;
  assign n205 = pi6  & ~pi9 ;
  assign n206 = ~pi4  & n205;
  assign n207 = ~pi1  & n74;
  assign n208 = ~n206 & ~n207;
  assign n209 = ~pi3  & ~n208;
  assign n210 = pi2  & n76;
  assign n211 = pi2  & pi3 ;
  assign n212 = pi4  & n205;
  assign n213 = n211 & n212;
  assign n214 = n205 & n210;
  assign n215 = ~pi3  & pi5 ;
  assign n216 = ~pi3  & n74;
  assign n217 = ~pi6  & n215;
  assign n218 = ~n206 & ~n463;
  assign n219 = ~pi2  & ~n218;
  assign n220 = ~n462 & ~n219;
  assign n221 = ~n209 & n220;
  assign n222 = ~pi7  & ~n221;
  assign n223 = ~pi10  & ~n222;
  assign n224 = ~pi8  & ~n198;
  assign n225 = ~pi10  & ~n462;
  assign n226 = ~n219 & n225;
  assign n227 = ~n209 & n225;
  assign n228 = ~n219 & n227;
  assign n229 = ~n209 & n226;
  assign n230 = ~pi7  & ~n464;
  assign n231 = ~n104 & ~n230;
  assign n232 = ~pi8  & ~n231;
  assign n233 = ~n223 & n224;
  assign n234 = ~n461 & ~n465;
  assign po1  = ~n197 & n234;
  assign n236 = pi0  & ~pi6 ;
  assign n237 = pi0  & ~pi3 ;
  assign n238 = pi4  & ~pi6 ;
  assign n239 = n237 & n238;
  assign n240 = n28 & n236;
  assign n241 = pi3  & ~pi4 ;
  assign n242 = pi3  & n59;
  assign n243 = pi5  & n241;
  assign n244 = ~n466 & ~n467;
  assign n245 = pi1  & ~n244;
  assign n246 = pi0  & pi1 ;
  assign n247 = pi4  & ~n246;
  assign n248 = pi3  & n247;
  assign n249 = n76 & ~n246;
  assign n250 = ~n164 & ~n468;
  assign n251 = ~pi5  & ~n250;
  assign n252 = ~n245 & ~n251;
  assign n253 = pi2  & ~n252;
  assign n254 = pi3  & ~pi6 ;
  assign n255 = ~pi2  & n254;
  assign n256 = ~pi6  & n107;
  assign n257 = ~n215 & ~n469;
  assign n258 = pi4  & ~n257;
  assign n259 = ~n253 & ~n258;
  assign n260 = ~pi7  & ~n259;
  assign n261 = pi5  & pi6 ;
  assign n262 = pi5  & ~n76;
  assign n263 = pi6  & n262;
  assign n264 = ~n76 & n261;
  assign n265 = pi2  & n70;
  assign n266 = ~n207 & ~n265;
  assign n267 = pi4  & ~n266;
  assign n268 = pi3  & n267;
  assign n269 = n76 & ~n266;
  assign n270 = ~n470 & ~n471;
  assign n271 = ~n260 & n270;
  assign n272 = ~pi8  & ~n271;
  assign n273 = pi4  & pi5 ;
  assign n274 = ~n20 & ~n254;
  assign n275 = pi3  & n103;
  assign n276 = pi6  & ~pi7 ;
  assign n277 = ~pi2  & n276;
  assign n278 = ~n275 & ~n277;
  assign n279 = ~n43 & ~n274;
  assign n280 = n273 & n472;
  assign n281 = ~n198 & ~n273;
  assign n282 = pi5  & ~n472;
  assign n283 = pi4  & n282;
  assign n284 = n273 & ~n472;
  assign n285 = pi7  & ~n273;
  assign n286 = pi6  & n285;
  assign n287 = n198 & ~n273;
  assign n288 = ~n473 & ~n474;
  assign n289 = ~n280 & ~n281;
  assign n290 = ~n272 & n475;
  assign n291 = ~pi9  & ~n290;
  assign n292 = n273 & n276;
  assign n293 = pi4  & pi6 ;
  assign n294 = n23 & n293;
  assign n295 = n128 & n261;
  assign n296 = ~n103 & ~n476;
  assign n297 = pi8  & ~n296;
  assign n298 = ~n291 & ~n297;
  assign n299 = ~pi10  & ~n298;
  assign n300 = pi5  & ~pi8 ;
  assign n301 = ~pi8  & pi9 ;
  assign n302 = pi5  & n301;
  assign n303 = pi9  & n300;
  assign n304 = ~n116 & ~n477;
  assign n305 = pi7  & ~n304;
  assign n306 = pi6  & n305;
  assign n307 = n198 & ~n304;
  assign n308 = pi5  & pi7 ;
  assign n309 = pi8  & ~n308;
  assign n310 = ~pi10  & ~n309;
  assign n311 = pi9  & ~n310;
  assign n312 = ~n478 & ~n311;
  assign n313 = ~n299 & n312;
  assign n314 = ~pi5  & ~pi6 ;
  assign n315 = n246 & n314;
  assign n316 = ~n476 & ~n315;
  assign n317 = pi3  & ~n316;
  assign n318 = pi2  & n317;
  assign n319 = n211 & ~n316;
  assign n320 = pi7  & ~n261;
  assign n321 = ~pi6  & ~n126;
  assign n322 = pi5  & n321;
  assign n323 = n74 & ~n126;
  assign n324 = pi5  & ~n126;
  assign n325 = ~pi7  & ~n324;
  assign n326 = ~n261 & ~n325;
  assign n327 = ~n320 & ~n480;
  assign n328 = pi4  & ~n215;
  assign n329 = pi4  & ~pi5 ;
  assign n330 = ~pi6  & ~n76;
  assign n331 = ~n329 & n330;
  assign n332 = ~pi6  & ~n328;
  assign n333 = ~n148 & ~n482;
  assign n334 = ~n481 & n333;
  assign n335 = ~n479 & n334;
  assign n336 = ~pi8  & ~n335;
  assign n337 = pi3  & pi8 ;
  assign n338 = ~n108 & ~n337;
  assign n339 = n199 & n273;
  assign n340 = pi6  & ~n338;
  assign n341 = pi5  & n340;
  assign n342 = pi7  & n341;
  assign n343 = ~pi9  & n342;
  assign n344 = pi4  & n343;
  assign n345 = ~n338 & n339;
  assign n346 = pi6  & pi8 ;
  assign n347 = pi7  & n261;
  assign n348 = pi6  & n308;
  assign n349 = pi8  & n484;
  assign n350 = pi8  & n198;
  assign n351 = pi5  & n350;
  assign n352 = n308 & n346;
  assign n353 = pi9  & ~n485;
  assign n354 = ~n483 & ~n353;
  assign n355 = ~pi7  & ~n74;
  assign n356 = ~pi3  & ~n355;
  assign n357 = ~pi4  & ~n276;
  assign n358 = ~pi9  & ~n357;
  assign n359 = ~n481 & n358;
  assign n360 = ~pi9  & ~n480;
  assign n361 = ~n320 & n360;
  assign n362 = ~n356 & n361;
  assign n363 = ~n357 & n362;
  assign n364 = ~n356 & n358;
  assign n365 = ~n481 & n364;
  assign n366 = ~n356 & n359;
  assign n367 = ~n479 & n486;
  assign n368 = ~pi8  & ~n367;
  assign n369 = pi9  & ~n484;
  assign n370 = ~n483 & ~n369;
  assign n371 = ~n368 & n370;
  assign n372 = ~n336 & n354;
  assign n373 = ~pi10  & ~n487;
  assign n374 = ~pi5  & ~pi7 ;
  assign n375 = ~pi8  & n374;
  assign n376 = ~pi5  & n92;
  assign n377 = pi1  & pi3 ;
  assign n378 = pi0  & n377;
  assign n379 = pi3  & n246;
  assign n380 = pi3  & ~pi5 ;
  assign n381 = n92 & n380;
  assign n382 = n246 & n381;
  assign n383 = n488 & n489;
  assign n384 = ~n485 & ~n490;
  assign n385 = pi2  & ~n384;
  assign n386 = pi8  & n308;
  assign n387 = pi3  & pi6 ;
  assign n388 = n386 & n387;
  assign n389 = pi6  & n337;
  assign n390 = n308 & n389;
  assign n391 = n337 & n484;
  assign n392 = ~n385 & ~n491;
  assign n393 = pi4  & ~n392;
  assign n394 = ~pi9  & ~pi10 ;
  assign n395 = n210 & n261;
  assign n396 = n92 & ~n314;
  assign n397 = n211 & n293;
  assign n398 = pi5  & ~n397;
  assign n399 = ~n70 & ~n398;
  assign n400 = ~pi7  & ~n399;
  assign n401 = ~pi8  & n400;
  assign n402 = n92 & ~n399;
  assign n403 = ~n395 & n396;
  assign n404 = n394 & ~n492;
  assign n405 = ~n393 & n404;
  assign n406 = ~pi4  & n92;
  assign n407 = ~pi7  & n38;
  assign n408 = n314 & n493;
  assign n409 = ~pi5  & n38;
  assign n410 = n43 & n409;
  assign n411 = n164 & n488;
  assign n412 = ~pi2  & n54;
  assign n413 = ~pi2  & n198;
  assign n414 = pi5  & n54;
  assign n415 = n413 & n414;
  assign n416 = ~pi2  & n273;
  assign n417 = n350 & n416;
  assign n418 = ~pi2  & pi5 ;
  assign n419 = n198 & n418;
  assign n420 = n54 & n419;
  assign n421 = n484 & n412;
  assign n422 = ~n494 & ~n495;
  assign n423 = ~pi3  & ~pi9 ;
  assign n424 = ~pi10  & n423;
  assign n425 = ~pi3  & n394;
  assign n426 = ~pi9  & ~n422;
  assign n427 = ~pi10  & n426;
  assign n428 = ~pi3  & n427;
  assign n429 = ~n422 & n496;
  assign n430 = n92 & n394;
  assign n431 = ~pi9  & ~n395;
  assign n432 = ~pi10  & n431;
  assign n433 = n92 & n432;
  assign n434 = ~n395 & n430;
  assign n435 = n24 | n25;
  assign n436 = n30 | n31;
  assign n437 = n39 | ~n40;
  assign n438 = n47 | n48;
  assign n439 = n53 | n51 | n52;
  assign n440 = n63 | n61 | n62;
  assign n441 = n64 | ~n65;
  assign n442 = n67 | n68;
  assign n443 = n72 | n73;
  assign n444 = n89 | n83 | n86 | n90 | n91;
  assign n445 = n98 | n99;
  assign n446 = n105 | n106;
  assign n447 = n112 | n113;
  assign n448 = n121 | n118 | n120;
  assign n449 = n137 | n135 | n136;
  assign n450 = n144 | n145;
  assign n451 = n154 | n150 | n153;
  assign n452 = n162 | n163;
  assign n453 = n165 | n166;
  assign n454 = n167 | ~n168;
  assign n455 = n179 | n171 | n178;
  assign n456 = n173 | n174;
  assign n457 = n185 | n186;
  assign n458 = n189 | n190;
  assign n459 = n195 | n196;
  assign n460 = n201 | n202;
  assign n461 = n203 | n204;
  assign n462 = n213 | n214;
  assign n463 = n216 | n217;
  assign n464 = n228 | n229;
  assign n465 = n232 | n233;
  assign n466 = n239 | n240;
  assign n467 = n242 | n243;
  assign n468 = n248 | n249;
  assign n469 = n255 | n256;
  assign n470 = n263 | n264;
  assign n471 = n268 | n269;
  assign n472 = n278 | ~n279;
  assign n473 = n283 | n284;
  assign n474 = n286 | n287;
  assign n475 = n288 | ~n289;
  assign n476 = n295 | n292 | n294;
  assign n477 = n302 | n303;
  assign n478 = n306 | n307;
  assign n479 = n318 | n319;
  assign n480 = n322 | n323;
  assign n481 = n326 | ~n327;
  assign n482 = n331 | n332;
  assign n483 = n344 | n345;
  assign n484 = n347 | n348;
  assign n485 = n352 | n349 | n351;
  assign n486 = n366 | n363 | n365;
  assign n487 = n371 | n372;
  assign n488 = n375 | n376;
  assign n489 = n378 | n379;
  assign n490 = n382 | n383;
  assign n491 = n391 | n388 | n390;
  assign n492 = n403 | n401 | n402;
  assign n493 = n406 | n407;
  assign n494 = n411 | n408 | n410;
  assign n495 = n415 | n417 | n420 | n421;
  assign n496 = n424 | n425;
  assign n497 = n428 | n429;
  assign n498 = n433 | n434;
  assign po0  = ~n125;
  assign po2  = ~n313;
  assign po3  = ~n497;
  assign po4  = ~n373;
  assign po5  = ~n405;
  assign po6  = ~n498;
endmodule
