module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n402, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412,
    n414, n415, n416, n417, n418, n419, n420,
    n421, n422, n423, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435,
    n437, n438, n439, n440, n441, n442, n443,
    n444, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n456, n457, n458, n459,
    n460, n461, n462, n463, n465, n466, n467,
    n468, n469, n470, n471, n473, n474, n475,
    n476, n477, n478, n479, n480, n482, n483,
    n484, n485, n486, n487, n488, n489, n491,
    n492, n493, n494, n495, n497, n498, n499,
    n500, n501, n502, n503, n505, n506, n507,
    n508, n509, n510, n511, n512, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n538, n539, n540, n541, n542, n543, n544,
    n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n559, n560,
    n561, n562, n563, n565, n566, n567, n568,
    n569, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n591,
    n592, n593, n594, n595, n596, n597, n598,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n609, n610, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n677, n678, n679, n680,
    n681, n682, n683, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695,
    n696, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n766, n767, n768,
    n769, n770, n771, n773, n774, n775, n776,
    n777, n778, n780, n781, n782, n783, n784,
    n785, n787, n788, n789, n790, n791, n792,
    n794, n795, n796, n797, n798, n799, n801,
    n802, n803, n804, n805, n806, n808, n809,
    n810, n811, n812, n813, n815, n816, n817,
    n818, n819, n820, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n845, n846, n847,
    n848, n849, n850, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869,
    n870, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899,
    n900, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n920, n921, n922,
    n923, n924, n925, n926, n928, n929, n930,
    n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n944, n945,
    n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n958, n959, n960,
    n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n990,
    n991, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1018, n1019, n1020, n1022, n1023, n1024,
    n1026, n1027, n1028, n1029, n1030, n1031,
    n1032, n1033, n1034, n1036, n1037, n1038,
    n1041, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078,
    n1080, n1081, n1082, n1083, n1084, n1085,
    n1087, n1088, n1089, n1090, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1108, n1109, n1110, n1112,
    n1113, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1124, n1125, n1126,
    n1128, n1129, n1130, n1132, n1133, n1134,
    n1136, n1137, n1138, n1139, n1140, n1142,
    n1143, n1144, n1146, n1147, n1148, n1150,
    n1151, n1152, n1154, n1155, n1156, n1158,
    n1159, n1160, n1162, n1163, n1164, n1166,
    n1167, n1168, n1170, n1171, n1172, n1174,
    n1175, n1176, n1178, n1179, n1180, n1182,
    n1183, n1184, n1186, n1187, n1188, n1189,
    n1190, n1192, n1193, n1194, n1196, n1197,
    n1198, n1200, n1201, n1202, n1204, n1205,
    n1206, n1208, n1209, n1210, n1211, n1212,
    n1213, n1214, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1227, n1228, n1229, n1231, n1232,
    n1233, n1234, n1236, n1237, n1238, n1240,
    n1241, n1242, n1244, n1245, n1246, n1247,
    n1248, n1250, n1251, n1252, n1254, n1255,
    n1256, n1258, n1259, n1260, n1262, n1263,
    n1264, n1266, n1267, n1268, n1270, n1271,
    n1272, n1273, n1274, n1275, n1276, n1278,
    n1279, n1280, n1281, n1282, n1283, n1285,
    n1286, n1287, n1289, n1290, n1291, n1293,
    n1294, n1295, n1297, n1298, n1299, n1301,
    n1302, n1303, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314,
    n1315, n1316, n1317, n1318, n1319, n1320,
    n1321, n1323, n1324, n1325, n1326, n1327,
    n1328, n1329, n1330, n1331, n1332, n1333,
    n1334, n1335, n1336, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1368, n1369, n1370, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384,
    n1386, n1387, n1388, n1390, n1391, n1392,
    n1393, n1394, n1395, n1396, n1397, n1398,
    n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1408, n1409, n1410, n1411,
    n1412, n1413, n1414, n1415, n1416, n1417,
    n1418, n1419, n1420, n1421, n1422, n1423,
    n1424, n1426, n1427, n1428, n1430, n1431,
    n1433, n1434, n1435, n1436, n1438, n1439,
    n1440, n1442, n1443, n1444, n1445, n1447,
    n1448, n1449, n1451, n1452, n1453, n1454,
    n1457, n1458, n1459, n1460, n1463, n1464,
    n1466, n1471, n1472, n1474;
  assign n291 = ~pi9 & ~pi11;
  assign n292 = ~pi5 & ~pi22;
  assign n293 = ~pi6 & ~pi12;
  assign n294 = ~pi4 & ~pi19;
  assign n295 = ~pi18 & n294;
  assign n296 = ~pi16 & n295;
  assign n297 = ~pi8 & ~pi21;
  assign n298 = ~pi7 & ~pi13;
  assign n299 = n297 & n298;
  assign n300 = ~pi14 & ~pi17;
  assign n301 = n291 & n300;
  assign n302 = n292 & n293;
  assign n303 = n301 & n302;
  assign n304 = n299 & n303;
  assign n305 = n296 & n304;
  assign n306 = pi54 & ~n305;
  assign n307 = ~pi0 & ~n306;
  assign n308 = ~pi7 & n297;
  assign n309 = pi8 & pi21;
  assign n310 = ~pi13 & ~n309;
  assign n311 = ~n308 & ~n310;
  assign n312 = ~pi14 & ~n311;
  assign n313 = ~n299 & ~n312;
  assign n314 = pi7 & ~n297;
  assign n315 = ~n299 & ~n314;
  assign n316 = ~pi14 & ~n315;
  assign n317 = ~pi10 & ~n316;
  assign n318 = ~n313 & n317;
  assign n319 = ~pi14 & n297;
  assign n320 = pi10 & n298;
  assign n321 = n319 & n320;
  assign n322 = ~n318 & ~n321;
  assign n323 = ~pi17 & n293;
  assign n324 = n296 & n323;
  assign n325 = ~n322 & n324;
  assign n326 = n292 & ~n325;
  assign n327 = pi56 & ~n292;
  assign n328 = n291 & ~n327;
  assign n329 = ~n326 & n328;
  assign n330 = ~pi56 & ~n291;
  assign n331 = n292 & n330;
  assign n332 = ~n329 & ~n331;
  assign n333 = pi54 & ~n332;
  assign n334 = ~n307 & ~n333;
  assign n335 = ~pi3 & ~pi129;
  assign po15 = n334 | ~n335;
  assign n337 = ~pi17 & pi54;
  assign n338 = ~pi10 & ~pi22;
  assign n339 = ~pi11 & ~pi12;
  assign n340 = ~pi5 & ~pi6;
  assign n341 = n298 & n340;
  assign n342 = n338 & n339;
  assign n343 = n319 & n342;
  assign n344 = n341 & n343;
  assign n345 = n296 & n344;
  assign n346 = n337 & ~n345;
  assign n347 = ~pi1 & ~n346;
  assign n348 = ~pi17 & n297;
  assign n349 = ~pi11 & n348;
  assign n350 = ~pi14 & pi54;
  assign n351 = n338 & n350;
  assign n352 = ~pi5 & n293;
  assign n353 = ~pi7 & n352;
  assign n354 = pi5 & ~n293;
  assign n355 = pi6 & pi12;
  assign n356 = ~pi7 & ~n355;
  assign n357 = ~n352 & ~n356;
  assign n358 = ~pi13 & ~n354;
  assign n359 = ~n357 & n358;
  assign n360 = ~n353 & ~n359;
  assign n361 = ~pi9 & ~n360;
  assign n362 = n298 & n352;
  assign n363 = ~n361 & ~n362;
  assign n364 = ~pi9 & n362;
  assign n365 = n296 & n351;
  assign n366 = n349 & n365;
  assign n367 = ~n364 & n366;
  assign n368 = ~n363 & n367;
  assign n369 = ~n347 & ~n368;
  assign po16 = ~n335 | n369;
  assign n371 = pi122 & pi127;
  assign n372 = ~pi82 & n371;
  assign n373 = ~pi47 & ~pi48;
  assign n374 = ~pi41 & ~pi43;
  assign n375 = ~pi46 & ~pi50;
  assign n376 = ~pi42 & ~pi44;
  assign n377 = ~pi40 & n376;
  assign n378 = n375 & n377;
  assign n379 = ~pi38 & n378;
  assign n380 = n374 & n379;
  assign n381 = ~pi45 & n373;
  assign n382 = n380 & n381;
  assign n383 = ~pi15 & ~pi20;
  assign n384 = ~pi24 & ~pi49;
  assign n385 = n383 & n384;
  assign n386 = n382 & n385;
  assign n387 = pi82 & ~n386;
  assign n388 = ~n372 & ~n387;
  assign n389 = pi2 & ~n388;
  assign n390 = ~pi45 & ~pi48;
  assign n391 = ~pi47 & n374;
  assign n392 = n379 & n391;
  assign n393 = n390 & n392;
  assign n394 = ~pi2 & n383;
  assign n395 = n384 & n394;
  assign n396 = n393 & n395;
  assign n397 = pi82 & ~n396;
  assign n398 = ~pi65 & ~n371;
  assign n399 = ~n397 & n398;
  assign n400 = ~n389 & ~n399;
  assign po17 = ~pi129 & ~n400;
  assign n402 = pi0 & ~pi113;
  assign n403 = ~pi123 & n402;
  assign n404 = ~pi12 & n349;
  assign n405 = ~pi9 & ~pi14;
  assign n406 = n338 & n405;
  assign n407 = n341 & n406;
  assign n408 = n296 & n407;
  assign n409 = n404 & n408;
  assign n410 = ~pi61 & ~pi118;
  assign n411 = ~n409 & n410;
  assign n412 = ~n403 & ~n411;
  assign po18 = ~pi129 & ~n412;
  assign n414 = pi4 & ~pi54;
  assign n415 = ~pi16 & pi54;
  assign n416 = n294 & n415;
  assign n417 = ~pi18 & n416;
  assign n418 = n349 & n417;
  assign n419 = pi10 & ~pi22;
  assign n420 = n405 & n419;
  assign n421 = n362 & n420;
  assign n422 = n418 & n421;
  assign n423 = ~n414 & ~n422;
  assign po19 = n335 & ~n423;
  assign n425 = pi5 & ~pi54;
  assign n426 = ~pi13 & n406;
  assign n427 = ~pi59 & n349;
  assign n428 = n426 & n427;
  assign n429 = ~pi7 & ~pi25;
  assign n430 = ~pi29 & n429;
  assign n431 = pi28 & n352;
  assign n432 = n430 & n431;
  assign n433 = n417 & n432;
  assign n434 = n428 & n433;
  assign n435 = ~n425 & ~n434;
  assign po20 = n335 & ~n435;
  assign n437 = pi6 & ~pi54;
  assign n438 = n353 & n415;
  assign n439 = pi25 & ~pi28;
  assign n440 = ~pi29 & n439;
  assign n441 = n295 & n440;
  assign n442 = n438 & n441;
  assign n443 = n428 & n442;
  assign n444 = ~n437 & ~n443;
  assign po21 = n335 & ~n444;
  assign n446 = pi7 & ~pi54;
  assign n447 = ~pi7 & n339;
  assign n448 = n340 & n447;
  assign n449 = pi8 & ~pi17;
  assign n450 = ~pi21 & n449;
  assign n451 = n417 & n450;
  assign n452 = n426 & n448;
  assign n453 = n451 & n452;
  assign n454 = ~n446 & ~n453;
  assign po22 = n335 & ~n454;
  assign n456 = pi8 & ~pi54;
  assign n457 = n362 & n406;
  assign n458 = ~pi8 & ~pi11;
  assign n459 = ~pi17 & pi21;
  assign n460 = n458 & n459;
  assign n461 = n417 & n460;
  assign n462 = n457 & n461;
  assign n463 = ~n456 & ~n462;
  assign po23 = n335 & ~n463;
  assign n465 = pi9 & ~pi54;
  assign n466 = ~pi18 & n348;
  assign n467 = pi11 & n294;
  assign n468 = n426 & n467;
  assign n469 = n466 & n468;
  assign n470 = n438 & n469;
  assign n471 = ~n465 & ~n470;
  assign po24 = n335 & ~n471;
  assign n473 = pi10 & ~pi54;
  assign n474 = ~pi9 & n466;
  assign n475 = n338 & n474;
  assign n476 = ~pi13 & pi14;
  assign n477 = n416 & n476;
  assign n478 = n448 & n477;
  assign n479 = n475 & n478;
  assign n480 = ~n473 & ~n479;
  assign po25 = n335 & ~n480;
  assign n482 = pi11 & ~pi54;
  assign n483 = ~pi10 & ~pi11;
  assign n484 = pi22 & n483;
  assign n485 = n405 & n484;
  assign n486 = n416 & n485;
  assign n487 = n362 & n466;
  assign n488 = n486 & n487;
  assign n489 = ~n482 & ~n488;
  assign po26 = n335 & ~n489;
  assign n491 = pi12 & ~pi54;
  assign n492 = pi18 & n416;
  assign n493 = n407 & n492;
  assign n494 = n404 & n493;
  assign n495 = ~n491 & ~n494;
  assign po27 = n335 & ~n495;
  assign n497 = pi13 & ~pi54;
  assign n498 = ~pi25 & ~pi28;
  assign n499 = pi29 & n498;
  assign n500 = n417 & n499;
  assign n501 = n427 & n500;
  assign n502 = n457 & n501;
  assign n503 = ~n497 & ~n502;
  assign po28 = n335 & ~n503;
  assign n505 = pi14 & ~pi54;
  assign n506 = ~pi4 & ~pi16;
  assign n507 = pi13 & ~pi19;
  assign n508 = n506 & n507;
  assign n509 = n351 & n508;
  assign n510 = n448 & n509;
  assign n511 = n474 & n510;
  assign n512 = ~n505 & ~n511;
  assign po29 = n335 & ~n512;
  assign n514 = pi15 & n372;
  assign n515 = ~pi43 & ~pi47;
  assign n516 = ~pi41 & n375;
  assign n517 = ~pi38 & ~pi40;
  assign n518 = n376 & n517;
  assign n519 = n516 & n518;
  assign n520 = n384 & n390;
  assign n521 = n515 & n520;
  assign n522 = n519 & n521;
  assign n523 = pi15 & ~n522;
  assign n524 = ~pi2 & ~pi20;
  assign n525 = ~pi15 & n384;
  assign n526 = ~n524 & n525;
  assign n527 = n382 & n526;
  assign n528 = ~n523 & ~n527;
  assign n529 = pi82 & ~n528;
  assign n530 = ~pi15 & n520;
  assign n531 = n392 & n530;
  assign n532 = pi82 & ~n531;
  assign n533 = ~pi70 & ~n371;
  assign n534 = ~n532 & n533;
  assign n535 = ~n514 & ~n534;
  assign n536 = ~n529 & n535;
  assign po30 = ~pi129 & ~n536;
  assign n538 = pi16 & ~pi54;
  assign n539 = ~pi5 & pi6;
  assign n540 = ~pi12 & n539;
  assign n541 = n298 & n540;
  assign n542 = n406 & n541;
  assign n543 = n418 & n542;
  assign n544 = ~n538 & ~n543;
  assign po31 = n335 & ~n544;
  assign n546 = pi17 & ~pi54;
  assign n547 = ~pi11 & n297;
  assign n548 = n295 & n547;
  assign n549 = ~pi12 & ~pi16;
  assign n550 = ~pi28 & pi59;
  assign n551 = n549 & n550;
  assign n552 = n337 & n340;
  assign n553 = n551 & n552;
  assign n554 = n430 & n553;
  assign n555 = n426 & n548;
  assign n556 = n554 & n555;
  assign n557 = ~n546 & ~n556;
  assign po32 = n335 & ~n557;
  assign n559 = pi18 & ~pi54;
  assign n560 = pi16 & n337;
  assign n561 = n548 & n560;
  assign n562 = n457 & n561;
  assign n563 = ~n559 & ~n562;
  assign po33 = n335 & ~n563;
  assign n565 = pi19 & ~pi54;
  assign n566 = pi17 & n547;
  assign n567 = n417 & n566;
  assign n568 = n457 & n567;
  assign n569 = ~n565 & ~n568;
  assign po34 = n335 & ~n569;
  assign n571 = pi20 & n372;
  assign n572 = ~pi41 & ~pi46;
  assign n573 = n515 & n572;
  assign n574 = n390 & n573;
  assign n575 = ~pi50 & n376;
  assign n576 = n517 & n575;
  assign n577 = n574 & n576;
  assign n578 = n384 & n577;
  assign n579 = n383 & n578;
  assign n580 = pi2 & n579;
  assign n581 = ~pi15 & n578;
  assign n582 = pi20 & ~n581;
  assign n583 = ~n580 & ~n582;
  assign n584 = pi82 & ~n583;
  assign n585 = pi82 & ~n579;
  assign n586 = ~pi71 & ~n371;
  assign n587 = ~n585 & n586;
  assign n588 = ~n571 & ~n587;
  assign n589 = ~n584 & n588;
  assign po35 = ~pi129 & ~n589;
  assign n591 = pi21 & ~pi54;
  assign n592 = pi19 & ~pi21;
  assign n593 = ~pi18 & n592;
  assign n594 = n337 & n458;
  assign n595 = n506 & n594;
  assign n596 = n593 & n595;
  assign n597 = n457 & n596;
  assign n598 = ~n591 & ~n597;
  assign po36 = n335 & ~n598;
  assign n600 = pi22 & ~pi54;
  assign n601 = pi5 & ~pi6;
  assign n602 = ~pi14 & n601;
  assign n603 = n298 & n339;
  assign n604 = n602 & n603;
  assign n605 = n416 & n604;
  assign n606 = n475 & n605;
  assign n607 = ~n600 & ~n606;
  assign po37 = n335 & ~n607;
  assign n609 = ~pi23 & pi55;
  assign n610 = pi61 & ~pi129;
  assign po38 = ~n609 & n610;
  assign n612 = ~pi44 & pi82;
  assign n613 = ~pi42 & n517;
  assign n614 = ~pi50 & n613;
  assign n615 = pi24 & n612;
  assign n616 = n574 & n615;
  assign n617 = n614 & n616;
  assign n618 = pi82 & ~n393;
  assign n619 = ~pi49 & n394;
  assign n620 = pi82 & ~n619;
  assign n621 = n371 & ~n620;
  assign n622 = ~n618 & ~n621;
  assign n623 = ~pi24 & ~n622;
  assign n624 = n382 & n619;
  assign n625 = pi82 & ~n624;
  assign n626 = pi63 & ~n371;
  assign n627 = ~n625 & n626;
  assign n628 = ~pi129 & ~n617;
  assign n629 = ~n623 & n628;
  assign po39 = ~n627 & n629;
  assign n631 = pi85 & ~pi116;
  assign n632 = pi25 & n631;
  assign n633 = ~pi96 & ~pi110;
  assign n634 = ~pi85 & ~n633;
  assign n635 = pi100 & ~n631;
  assign n636 = ~n634 & n635;
  assign n637 = ~n632 & ~n636;
  assign n638 = ~pi26 & ~n637;
  assign n639 = pi25 & ~pi116;
  assign n640 = pi26 & n639;
  assign n641 = ~pi95 & ~pi100;
  assign n642 = ~pi97 & n641;
  assign n643 = ~pi110 & ~n642;
  assign n644 = pi25 & ~n643;
  assign n645 = pi26 & pi116;
  assign n646 = ~n644 & ~n645;
  assign n647 = ~pi51 & ~pi52;
  assign n648 = ~pi39 & n647;
  assign n649 = ~n646 & ~n648;
  assign n650 = ~n640 & ~n649;
  assign n651 = ~pi85 & ~n650;
  assign n652 = ~n638 & ~n651;
  assign n653 = ~pi27 & ~n652;
  assign n654 = ~pi39 & ~pi52;
  assign n655 = ~pi51 & n654;
  assign n656 = pi116 & n655;
  assign n657 = ~n639 & ~n656;
  assign n658 = pi27 & ~n657;
  assign n659 = n644 & n648;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~pi26 & ~pi85;
  assign n662 = ~n660 & n661;
  assign n663 = ~n653 & ~n662;
  assign n664 = ~pi53 & ~n663;
  assign n665 = ~pi26 & n639;
  assign n666 = pi53 & ~pi85;
  assign n667 = ~pi27 & n666;
  assign n668 = n665 & n667;
  assign n669 = ~n664 & ~n668;
  assign n670 = ~pi58 & ~n669;
  assign n671 = ~pi27 & ~pi85;
  assign n672 = ~pi53 & pi58;
  assign n673 = n671 & n672;
  assign n674 = n665 & n673;
  assign n675 = ~n670 & ~n674;
  assign po40 = n335 & ~n675;
  assign n677 = ~pi27 & ~pi53;
  assign n678 = ~pi58 & n677;
  assign n679 = ~pi85 & ~n656;
  assign n680 = pi26 & n679;
  assign n681 = n636 & ~n645;
  assign n682 = ~n680 & ~n681;
  assign n683 = n335 & n678;
  assign po41 = ~n682 & n683;
  assign n685 = ~pi53 & ~pi58;
  assign n686 = ~pi26 & n335;
  assign n687 = pi27 & n679;
  assign n688 = pi27 & pi116;
  assign n689 = pi85 & pi116;
  assign n690 = pi95 & ~n631;
  assign n691 = n633 & n690;
  assign n692 = ~n689 & ~n691;
  assign n693 = ~pi100 & ~n688;
  assign n694 = ~n692 & n693;
  assign n695 = ~n687 & ~n694;
  assign n696 = n685 & n686;
  assign po42 = ~n695 & n696;
  assign n698 = ~pi26 & ~pi27;
  assign n699 = ~pi28 & ~pi116;
  assign n700 = pi100 & pi116;
  assign n701 = n698 & ~n699;
  assign n702 = ~n700 & n701;
  assign n703 = pi85 & ~n702;
  assign n704 = ~pi26 & ~n648;
  assign n705 = n688 & n704;
  assign n706 = ~pi27 & n655;
  assign n707 = ~n704 & ~n706;
  assign n708 = ~n643 & ~n707;
  assign n709 = pi26 & ~pi27;
  assign n710 = ~pi26 & pi27;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~pi116 & ~n711;
  assign n713 = ~n708 & ~n712;
  assign n714 = pi28 & ~n713;
  assign n715 = ~pi26 & pi95;
  assign n716 = ~pi100 & n715;
  assign n717 = n633 & n716;
  assign n718 = pi26 & n656;
  assign n719 = ~n717 & ~n718;
  assign n720 = ~pi27 & ~n719;
  assign n721 = ~pi85 & ~n705;
  assign n722 = ~n720 & n721;
  assign n723 = ~n714 & n722;
  assign n724 = ~pi53 & ~n703;
  assign n725 = ~n723 & n724;
  assign n726 = ~pi27 & pi28;
  assign n727 = ~pi116 & n726;
  assign n728 = ~pi26 & n666;
  assign n729 = n727 & n728;
  assign n730 = ~n725 & ~n729;
  assign n731 = ~pi58 & ~n730;
  assign n732 = n661 & n672;
  assign n733 = n727 & n732;
  assign n734 = ~n731 & ~n733;
  assign po43 = n335 & ~n734;
  assign n736 = pi97 & pi116;
  assign n737 = pi29 & ~pi116;
  assign n738 = pi58 & ~n736;
  assign n739 = ~n737 & n738;
  assign n740 = pi29 & pi110;
  assign n741 = ~pi29 & ~pi97;
  assign n742 = pi97 & ~n633;
  assign n743 = n641 & ~n741;
  assign n744 = ~n742 & n743;
  assign n745 = ~pi58 & ~n740;
  assign n746 = ~n744 & n745;
  assign n747 = ~pi53 & ~n739;
  assign n748 = ~n746 & n747;
  assign n749 = pi53 & ~pi58;
  assign n750 = n737 & n749;
  assign n751 = ~n748 & ~n750;
  assign n752 = ~pi27 & ~n751;
  assign n753 = pi27 & n685;
  assign n754 = n737 & n753;
  assign n755 = ~n752 & ~n754;
  assign n756 = ~pi85 & ~n755;
  assign n757 = pi85 & n737;
  assign n758 = n678 & n757;
  assign n759 = ~n756 & ~n758;
  assign n760 = ~pi26 & ~n759;
  assign n761 = ~pi85 & n685;
  assign n762 = n709 & n761;
  assign n763 = n737 & n762;
  assign n764 = ~n760 & ~n763;
  assign po44 = n335 & ~n764;
  assign n766 = ~pi88 & pi106;
  assign n767 = pi30 & ~pi109;
  assign n768 = pi60 & pi109;
  assign n769 = ~pi106 & ~n767;
  assign n770 = ~n768 & n769;
  assign n771 = ~pi129 & ~n766;
  assign po45 = ~n770 & n771;
  assign n773 = ~pi89 & pi106;
  assign n774 = pi31 & ~pi109;
  assign n775 = pi30 & pi109;
  assign n776 = ~pi106 & ~n774;
  assign n777 = ~n775 & n776;
  assign n778 = ~pi129 & ~n773;
  assign po46 = ~n777 & n778;
  assign n780 = ~pi99 & pi106;
  assign n781 = pi32 & ~pi109;
  assign n782 = pi31 & pi109;
  assign n783 = ~pi106 & ~n781;
  assign n784 = ~n782 & n783;
  assign n785 = ~pi129 & ~n780;
  assign po47 = ~n784 & n785;
  assign n787 = ~pi90 & pi106;
  assign n788 = pi33 & ~pi109;
  assign n789 = pi32 & pi109;
  assign n790 = ~pi106 & ~n788;
  assign n791 = ~n789 & n790;
  assign n792 = ~pi129 & ~n787;
  assign po48 = ~n791 & n792;
  assign n794 = ~pi91 & pi106;
  assign n795 = pi34 & ~pi109;
  assign n796 = pi33 & pi109;
  assign n797 = ~pi106 & ~n795;
  assign n798 = ~n796 & n797;
  assign n799 = ~pi129 & ~n794;
  assign po49 = ~n798 & n799;
  assign n801 = ~pi92 & pi106;
  assign n802 = pi35 & ~pi109;
  assign n803 = pi34 & pi109;
  assign n804 = ~pi106 & ~n802;
  assign n805 = ~n803 & n804;
  assign n806 = ~pi129 & ~n801;
  assign po50 = ~n805 & n806;
  assign n808 = ~pi98 & pi106;
  assign n809 = pi36 & ~pi109;
  assign n810 = pi35 & pi109;
  assign n811 = ~pi106 & ~n809;
  assign n812 = ~n810 & n811;
  assign n813 = ~pi129 & ~n808;
  assign po51 = ~n812 & n813;
  assign n815 = ~pi93 & pi106;
  assign n816 = pi37 & ~pi109;
  assign n817 = pi36 & pi109;
  assign n818 = ~pi106 & ~n816;
  assign n819 = ~n817 & n818;
  assign n820 = ~pi129 & ~n815;
  assign po52 = ~n819 & n820;
  assign n822 = pi82 & ~n377;
  assign n823 = ~pi43 & n373;
  assign n824 = n572 & n823;
  assign n825 = ~pi50 & n824;
  assign n826 = ~pi2 & ~pi45;
  assign n827 = n385 & n826;
  assign n828 = n825 & n827;
  assign n829 = pi82 & ~n828;
  assign n830 = n371 & ~n829;
  assign n831 = ~n822 & ~n830;
  assign n832 = ~pi38 & ~n831;
  assign n833 = ~pi42 & n612;
  assign n834 = ~pi40 & n833;
  assign n835 = pi38 & n834;
  assign n836 = n390 & n395;
  assign n837 = n391 & n836;
  assign n838 = n378 & n837;
  assign n839 = pi82 & ~n838;
  assign n840 = pi74 & ~n371;
  assign n841 = ~n839 & n840;
  assign n842 = ~pi129 & ~n835;
  assign n843 = ~n841 & n842;
  assign po53 = ~n832 & n843;
  assign n845 = pi109 & n647;
  assign n846 = pi39 & ~n845;
  assign n847 = ~pi51 & pi109;
  assign n848 = n654 & n847;
  assign n849 = ~pi106 & ~n848;
  assign n850 = ~n846 & n849;
  assign po54 = ~pi129 & ~n850;
  assign n852 = pi82 & ~n376;
  assign n853 = ~pi48 & n515;
  assign n854 = n827 & n853;
  assign n855 = ~pi38 & n516;
  assign n856 = n854 & n855;
  assign n857 = pi82 & ~n856;
  assign n858 = n371 & ~n857;
  assign n859 = ~n852 & ~n858;
  assign n860 = ~pi40 & ~n859;
  assign n861 = pi40 & n833;
  assign n862 = ~pi38 & ~pi46;
  assign n863 = ~pi50 & n862;
  assign n864 = n376 & n863;
  assign n865 = n837 & n864;
  assign n866 = pi82 & ~n865;
  assign n867 = pi73 & ~n371;
  assign n868 = ~n866 & n867;
  assign n869 = ~pi129 & ~n861;
  assign n870 = ~n868 & n869;
  assign po55 = ~n860 & n870;
  assign n872 = pi82 & ~n379;
  assign n873 = pi82 & ~n854;
  assign n874 = n371 & ~n873;
  assign n875 = ~n872 & ~n874;
  assign n876 = ~pi41 & ~n875;
  assign n877 = n375 & n517;
  assign n878 = pi41 & n833;
  assign n879 = n877 & n878;
  assign n880 = n379 & n515;
  assign n881 = n836 & n880;
  assign n882 = pi82 & ~n881;
  assign n883 = pi76 & ~n371;
  assign n884 = ~n882 & n883;
  assign n885 = ~pi129 & ~n879;
  assign n886 = ~n876 & n885;
  assign po56 = ~n884 & n886;
  assign n888 = pi44 & pi82;
  assign n889 = n837 & n877;
  assign n890 = pi82 & ~n889;
  assign n891 = n371 & ~n890;
  assign n892 = ~n888 & ~n891;
  assign n893 = ~pi42 & ~n892;
  assign n894 = pi42 & n612;
  assign n895 = ~pi44 & n889;
  assign n896 = pi82 & ~n895;
  assign n897 = pi72 & ~n371;
  assign n898 = ~n896 & n897;
  assign n899 = ~pi129 & ~n894;
  assign n900 = ~n898 & n899;
  assign po57 = ~n893 & n900;
  assign n902 = pi82 & ~n519;
  assign n903 = ~pi2 & n373;
  assign n904 = n385 & n903;
  assign n905 = ~pi45 & n904;
  assign n906 = pi82 & ~n905;
  assign n907 = n371 & ~n906;
  assign n908 = ~n902 & ~n907;
  assign n909 = ~pi43 & ~n908;
  assign n910 = pi43 & n834;
  assign n911 = n855 & n910;
  assign n912 = ~pi47 & n519;
  assign n913 = n836 & n912;
  assign n914 = pi82 & ~n913;
  assign n915 = pi77 & ~n371;
  assign n916 = ~n914 & n915;
  assign n917 = ~pi129 & ~n911;
  assign n918 = ~n916 & n917;
  assign po58 = ~n909 & n918;
  assign n920 = ~pi42 & n889;
  assign n921 = pi82 & ~n920;
  assign n922 = ~pi67 & ~n371;
  assign n923 = pi44 & n371;
  assign n924 = ~n922 & ~n923;
  assign n925 = ~n921 & n924;
  assign n926 = ~pi129 & ~n888;
  assign po59 = ~n925 & n926;
  assign n928 = pi45 & pi82;
  assign n929 = n518 & n928;
  assign n930 = n825 & n929;
  assign n931 = pi82 & ~n395;
  assign n932 = n371 & ~n931;
  assign n933 = n518 & n825;
  assign n934 = pi82 & ~n933;
  assign n935 = ~n932 & ~n934;
  assign n936 = ~pi45 & ~n935;
  assign n937 = n380 & n904;
  assign n938 = pi82 & ~n937;
  assign n939 = pi68 & ~n371;
  assign n940 = ~n938 & n939;
  assign n941 = ~pi129 & ~n930;
  assign n942 = ~n936 & n941;
  assign po60 = ~n940 & n942;
  assign n944 = pi82 & ~n576;
  assign n945 = pi82 & ~n837;
  assign n946 = n371 & ~n945;
  assign n947 = ~n944 & ~n946;
  assign n948 = ~pi46 & ~n947;
  assign n949 = pi46 & n612;
  assign n950 = n614 & n949;
  assign n951 = n576 & n837;
  assign n952 = pi82 & ~n951;
  assign n953 = pi75 & ~n371;
  assign n954 = ~n952 & n953;
  assign n955 = ~pi129 & ~n950;
  assign n956 = ~n954 & n955;
  assign po61 = ~n948 & n956;
  assign n958 = pi47 & n374;
  assign n959 = n863 & n958;
  assign n960 = n834 & n959;
  assign n961 = pi82 & ~n380;
  assign n962 = pi82 & ~n836;
  assign n963 = n371 & ~n962;
  assign n964 = ~n961 & ~n963;
  assign n965 = ~pi47 & ~n964;
  assign n966 = n380 & n836;
  assign n967 = pi82 & ~n966;
  assign n968 = pi64 & ~n371;
  assign n969 = ~n967 & n968;
  assign n970 = ~pi129 & ~n960;
  assign n971 = ~n965 & n970;
  assign po62 = ~n969 & n971;
  assign n973 = pi48 & n515;
  assign n974 = n612 & n973;
  assign n975 = n516 & n613;
  assign n976 = n974 & n975;
  assign n977 = pi82 & ~n827;
  assign n978 = n371 & ~n977;
  assign n979 = n573 & n576;
  assign n980 = pi82 & ~n979;
  assign n981 = ~n978 & ~n980;
  assign n982 = ~pi48 & ~n981;
  assign n983 = n392 & n827;
  assign n984 = pi82 & ~n983;
  assign n985 = pi62 & ~n371;
  assign n986 = ~n984 & n985;
  assign n987 = ~pi129 & ~n976;
  assign n988 = ~n982 & n987;
  assign po63 = ~n986 & n988;
  assign n990 = pi49 & n372;
  assign n991 = ~pi24 & n577;
  assign n992 = pi49 & ~n991;
  assign n993 = ~n394 & n578;
  assign n994 = ~n992 & ~n993;
  assign n995 = pi82 & ~n994;
  assign n996 = pi82 & ~n578;
  assign n997 = ~pi69 & ~n371;
  assign n998 = ~n996 & n997;
  assign n999 = ~n990 & ~n998;
  assign n1000 = ~n995 & n999;
  assign po64 = ~pi129 & ~n1000;
  assign n1002 = pi50 & pi82;
  assign n1003 = n518 & n1002;
  assign n1004 = pi82 & ~n518;
  assign n1005 = n824 & n827;
  assign n1006 = pi82 & ~n1005;
  assign n1007 = n371 & ~n1006;
  assign n1008 = ~n1004 & ~n1007;
  assign n1009 = ~pi50 & ~n1008;
  assign n1010 = n377 & n862;
  assign n1011 = n837 & n1010;
  assign n1012 = pi82 & ~n1011;
  assign n1013 = pi66 & ~n371;
  assign n1014 = ~n1012 & n1013;
  assign n1015 = ~pi129 & ~n1003;
  assign n1016 = ~n1009 & n1015;
  assign po65 = ~n1014 & n1016;
  assign n1018 = pi51 & ~pi109;
  assign n1019 = ~pi106 & ~n847;
  assign n1020 = ~n1018 & n1019;
  assign po66 = ~pi129 & ~n1020;
  assign n1022 = pi52 & ~n847;
  assign n1023 = ~pi106 & ~n845;
  assign n1024 = ~n1022 & n1023;
  assign po67 = ~pi129 & ~n1024;
  assign n1026 = ~pi116 & n749;
  assign n1027 = pi58 & pi116;
  assign n1028 = ~pi58 & n633;
  assign n1029 = n641 & n1028;
  assign n1030 = ~n1027 & ~n1029;
  assign n1031 = ~pi53 & pi97;
  assign n1032 = ~n1030 & n1031;
  assign n1033 = ~n1026 & ~n1032;
  assign n1034 = n671 & n686;
  assign po68 = ~n1033 & n1034;
  assign n1036 = n380 & n905;
  assign n1037 = pi82 & ~n1036;
  assign n1038 = ~n371 & ~n1037;
  assign po69 = pi129 | n1038;
  assign po129 = pi123 | pi129;
  assign n1041 = pi114 & ~pi122;
  assign po70 = ~po129 & n1041;
  assign n1043 = ~pi26 & pi58;
  assign n1044 = ~pi58 & n645;
  assign n1045 = ~n1043 & ~n1044;
  assign n1046 = pi94 & ~n1045;
  assign n1047 = pi58 & ~pi116;
  assign n1048 = pi37 & ~pi116;
  assign n1049 = ~n1043 & ~n1048;
  assign n1050 = ~n1047 & ~n1049;
  assign n1051 = ~n1046 & ~n1050;
  assign n1052 = ~pi53 & ~n1051;
  assign n1053 = ~pi26 & pi37;
  assign n1054 = ~pi58 & n1053;
  assign n1055 = ~n1052 & ~n1054;
  assign n1056 = ~pi85 & ~n1055;
  assign n1057 = n685 & n1053;
  assign n1058 = ~n1056 & ~n1057;
  assign n1059 = ~pi27 & ~n1058;
  assign n1060 = n761 & n1053;
  assign n1061 = ~n1059 & ~n1060;
  assign po71 = n335 & ~n1061;
  assign n1063 = ~pi26 & ~pi53;
  assign n1064 = ~pi85 & n1063;
  assign n1065 = ~pi116 & n1064;
  assign n1066 = pi26 & pi53;
  assign n1067 = pi85 & ~n1063;
  assign n1068 = ~pi58 & ~n1066;
  assign n1069 = ~n1067 & n1068;
  assign n1070 = ~n1065 & ~n1069;
  assign n1071 = pi57 & ~n1070;
  assign n1072 = pi60 & n1027;
  assign n1073 = n1064 & n1072;
  assign n1074 = ~n1071 & ~n1073;
  assign n1075 = ~pi27 & ~n1074;
  assign n1076 = pi57 & ~pi58;
  assign n1077 = n1064 & n1076;
  assign n1078 = ~n1075 & ~n1077;
  assign po72 = n335 & ~n1078;
  assign n1080 = n698 & n1047;
  assign n1081 = ~pi58 & ~n711;
  assign n1082 = n656 & n1081;
  assign n1083 = ~n1080 & ~n1082;
  assign n1084 = ~pi53 & ~pi85;
  assign n1085 = n335 & n1084;
  assign po73 = ~n1083 & n1085;
  assign n1087 = ~n672 & ~n749;
  assign n1088 = ~pi116 & ~n1087;
  assign n1089 = ~n643 & n685;
  assign n1090 = ~n1088 & ~n1089;
  assign n1091 = pi59 & ~n1090;
  assign n1092 = pi96 & n685;
  assign n1093 = n643 & n1092;
  assign n1094 = ~n1091 & ~n1093;
  assign n1095 = ~pi85 & ~n1094;
  assign n1096 = pi59 & ~pi116;
  assign n1097 = pi85 & n685;
  assign n1098 = n1096 & n1097;
  assign n1099 = ~n1095 & ~n1098;
  assign n1100 = ~pi27 & ~n1099;
  assign n1101 = pi27 & n1096;
  assign n1102 = n761 & n1101;
  assign n1103 = ~n1100 & ~n1102;
  assign n1104 = ~pi26 & ~n1103;
  assign n1105 = n762 & n1096;
  assign n1106 = ~n1104 & ~n1105;
  assign po74 = n335 & ~n1106;
  assign n1108 = ~pi117 & ~pi122;
  assign n1109 = pi60 & ~n1108;
  assign n1110 = pi123 & n1108;
  assign po75 = n1109 | n1110;
  assign n1112 = ~pi114 & ~pi122;
  assign n1113 = pi123 & ~pi129;
  assign po76 = n1112 & n1113;
  assign n1115 = pi136 & ~pi137;
  assign n1116 = pi131 & pi132;
  assign n1117 = pi133 & n1116;
  assign n1118 = ~pi138 & n1117;
  assign n1119 = n1115 & n1118;
  assign n1120 = ~pi62 & ~n1119;
  assign n1121 = pi140 & n1119;
  assign n1122 = ~pi129 & ~n1120;
  assign po77 = n1121 | ~n1122;
  assign n1124 = ~pi63 & ~n1119;
  assign n1125 = pi142 & n1119;
  assign n1126 = ~pi129 & ~n1124;
  assign po78 = n1125 | ~n1126;
  assign n1128 = ~pi64 & ~n1119;
  assign n1129 = pi139 & n1119;
  assign n1130 = ~pi129 & ~n1128;
  assign po79 = n1129 | ~n1130;
  assign n1132 = ~pi65 & ~n1119;
  assign n1133 = pi146 & n1119;
  assign n1134 = ~pi129 & ~n1132;
  assign po80 = n1133 | ~n1134;
  assign n1136 = ~pi136 & ~pi137;
  assign n1137 = n1118 & n1136;
  assign n1138 = ~pi66 & ~n1137;
  assign n1139 = pi143 & n1137;
  assign n1140 = ~pi129 & ~n1138;
  assign po81 = n1139 | ~n1140;
  assign n1142 = ~pi67 & ~n1137;
  assign n1143 = pi139 & n1137;
  assign n1144 = ~pi129 & ~n1142;
  assign po82 = n1143 | ~n1144;
  assign n1146 = ~pi68 & ~n1119;
  assign n1147 = pi141 & n1119;
  assign n1148 = ~pi129 & ~n1146;
  assign po83 = n1147 | ~n1148;
  assign n1150 = ~pi69 & ~n1119;
  assign n1151 = pi143 & n1119;
  assign n1152 = ~pi129 & ~n1150;
  assign po84 = n1151 | ~n1152;
  assign n1154 = ~pi70 & ~n1119;
  assign n1155 = pi144 & n1119;
  assign n1156 = ~pi129 & ~n1154;
  assign po85 = n1155 | ~n1156;
  assign n1158 = ~pi71 & ~n1119;
  assign n1159 = pi145 & n1119;
  assign n1160 = ~pi129 & ~n1158;
  assign po86 = n1159 | ~n1160;
  assign n1162 = ~pi72 & ~n1137;
  assign n1163 = pi140 & n1137;
  assign n1164 = ~pi129 & ~n1162;
  assign po87 = n1163 | ~n1164;
  assign n1166 = ~pi73 & ~n1137;
  assign n1167 = pi141 & n1137;
  assign n1168 = ~pi129 & ~n1166;
  assign po88 = n1167 | ~n1168;
  assign n1170 = ~pi74 & ~n1137;
  assign n1171 = pi142 & n1137;
  assign n1172 = ~pi129 & ~n1170;
  assign po89 = n1171 | ~n1172;
  assign n1174 = ~pi75 & ~n1137;
  assign n1175 = pi144 & n1137;
  assign n1176 = ~pi129 & ~n1174;
  assign po90 = n1175 | ~n1176;
  assign n1178 = ~pi76 & ~n1137;
  assign n1179 = pi145 & n1137;
  assign n1180 = ~pi129 & ~n1178;
  assign po91 = n1179 | ~n1180;
  assign n1182 = ~pi77 & ~n1137;
  assign n1183 = pi146 & n1137;
  assign n1184 = ~pi129 & ~n1182;
  assign po92 = n1183 | ~n1184;
  assign n1186 = ~pi136 & pi137;
  assign n1187 = n1118 & n1186;
  assign n1188 = ~pi78 & ~n1187;
  assign n1189 = ~pi142 & n1187;
  assign n1190 = ~pi129 & ~n1188;
  assign po93 = ~n1189 & n1190;
  assign n1192 = ~pi79 & ~n1187;
  assign n1193 = ~pi143 & n1187;
  assign n1194 = ~pi129 & ~n1192;
  assign po94 = ~n1193 & n1194;
  assign n1196 = ~pi80 & ~n1187;
  assign n1197 = ~pi144 & n1187;
  assign n1198 = ~pi129 & ~n1196;
  assign po95 = ~n1197 & n1198;
  assign n1200 = ~pi81 & ~n1187;
  assign n1201 = ~pi145 & n1187;
  assign n1202 = ~pi129 & ~n1200;
  assign po96 = ~n1201 & n1202;
  assign n1204 = ~pi82 & ~n1187;
  assign n1205 = ~pi146 & n1187;
  assign n1206 = ~pi129 & ~n1204;
  assign po97 = ~n1205 & n1206;
  assign n1208 = ~pi89 & pi138;
  assign n1209 = pi62 & ~pi138;
  assign n1210 = pi136 & ~n1208;
  assign n1211 = ~n1209 & n1210;
  assign n1212 = ~pi119 & pi138;
  assign n1213 = pi72 & ~pi138;
  assign n1214 = ~pi136 & ~n1212;
  assign n1215 = ~n1213 & n1214;
  assign n1216 = ~n1211 & ~n1215;
  assign n1217 = ~pi137 & ~n1216;
  assign n1218 = pi136 & ~pi138;
  assign n1219 = pi31 & n1218;
  assign n1220 = ~pi87 & ~pi138;
  assign n1221 = pi115 & pi138;
  assign n1222 = ~pi136 & ~n1220;
  assign n1223 = ~n1221 & n1222;
  assign n1224 = ~n1219 & ~n1223;
  assign n1225 = pi137 & ~n1224;
  assign po98 = n1217 | n1225;
  assign n1227 = ~pi84 & ~n1187;
  assign n1228 = ~pi141 & n1187;
  assign n1229 = ~pi129 & ~n1227;
  assign po99 = ~n1228 & n1229;
  assign n1231 = ~pi85 & n643;
  assign n1232 = pi96 & n1231;
  assign n1233 = ~n631 & ~n1232;
  assign n1234 = n678 & n686;
  assign po100 = ~n1233 & n1234;
  assign n1236 = ~pi86 & ~n1187;
  assign n1237 = ~pi139 & n1187;
  assign n1238 = ~pi129 & ~n1236;
  assign po101 = ~n1237 & n1238;
  assign n1240 = ~pi87 & ~n1187;
  assign n1241 = ~pi140 & n1187;
  assign n1242 = ~pi129 & ~n1240;
  assign po102 = ~n1241 & n1242;
  assign n1244 = pi137 & n1218;
  assign n1245 = n1117 & n1244;
  assign n1246 = ~pi88 & ~n1245;
  assign n1247 = ~pi139 & n1245;
  assign n1248 = ~pi129 & ~n1246;
  assign po103 = ~n1247 & n1248;
  assign n1250 = ~pi89 & ~n1245;
  assign n1251 = ~pi140 & n1245;
  assign n1252 = ~pi129 & ~n1250;
  assign po104 = ~n1251 & n1252;
  assign n1254 = ~pi90 & ~n1245;
  assign n1255 = ~pi142 & n1245;
  assign n1256 = ~pi129 & ~n1254;
  assign po105 = ~n1255 & n1256;
  assign n1258 = ~pi91 & ~n1245;
  assign n1259 = ~pi143 & n1245;
  assign n1260 = ~pi129 & ~n1258;
  assign po106 = ~n1259 & n1260;
  assign n1262 = ~pi92 & ~n1245;
  assign n1263 = ~pi144 & n1245;
  assign n1264 = ~pi129 & ~n1262;
  assign po107 = ~n1263 & n1264;
  assign n1266 = ~pi93 & ~n1245;
  assign n1267 = ~pi146 & n1245;
  assign n1268 = ~pi129 & ~n1266;
  assign po108 = ~n1267 & n1268;
  assign n1270 = pi82 & ~pi136;
  assign n1271 = ~pi137 & pi138;
  assign n1272 = n1270 & n1271;
  assign n1273 = n1117 & n1272;
  assign n1274 = ~pi94 & ~n1273;
  assign n1275 = ~pi142 & n1273;
  assign n1276 = ~pi129 & ~n1274;
  assign po109 = ~n1275 & n1276;
  assign n1278 = ~pi3 & ~pi110;
  assign n1279 = ~n1117 & ~n1278;
  assign n1280 = ~n1273 & ~n1279;
  assign n1281 = pi95 & n1280;
  assign n1282 = pi143 & n1273;
  assign n1283 = ~n1281 & ~n1282;
  assign po110 = ~pi129 & ~n1283;
  assign n1285 = pi96 & n1280;
  assign n1286 = pi146 & n1273;
  assign n1287 = ~n1285 & ~n1286;
  assign po111 = ~pi129 & ~n1287;
  assign n1289 = pi97 & n1280;
  assign n1290 = pi145 & n1273;
  assign n1291 = ~n1289 & ~n1290;
  assign po112 = ~pi129 & ~n1291;
  assign n1293 = ~pi98 & ~n1245;
  assign n1294 = ~pi145 & n1245;
  assign n1295 = ~pi129 & ~n1293;
  assign po113 = ~n1294 & n1295;
  assign n1297 = ~pi99 & ~n1245;
  assign n1298 = ~pi141 & n1245;
  assign n1299 = ~pi129 & ~n1297;
  assign po114 = ~n1298 & n1299;
  assign n1301 = pi100 & n1280;
  assign n1302 = pi144 & n1273;
  assign n1303 = ~n1301 & ~n1302;
  assign po115 = ~pi129 & ~n1303;
  assign n1305 = ~pi124 & pi138;
  assign n1306 = pi77 & ~pi138;
  assign n1307 = ~pi136 & ~n1305;
  assign n1308 = ~n1306 & n1307;
  assign n1309 = ~pi93 & pi138;
  assign n1310 = pi65 & ~pi138;
  assign n1311 = pi136 & ~n1309;
  assign n1312 = ~n1310 & n1311;
  assign n1313 = ~n1308 & ~n1312;
  assign n1314 = ~pi137 & ~n1313;
  assign n1315 = pi37 & n1218;
  assign n1316 = ~pi82 & ~pi138;
  assign n1317 = ~pi96 & pi138;
  assign n1318 = ~pi136 & ~n1316;
  assign n1319 = ~n1317 & n1318;
  assign n1320 = ~n1315 & ~n1319;
  assign n1321 = pi137 & ~n1320;
  assign po116 = n1314 | n1321;
  assign n1323 = pi91 & n1115;
  assign n1324 = pi95 & n1186;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = pi138 & ~n1325;
  assign n1327 = ~pi79 & ~pi136;
  assign n1328 = ~pi34 & pi136;
  assign n1329 = pi137 & ~n1327;
  assign n1330 = ~n1328 & n1329;
  assign n1331 = pi66 & ~pi136;
  assign n1332 = pi69 & pi136;
  assign n1333 = ~pi137 & ~n1331;
  assign n1334 = ~n1332 & n1333;
  assign n1335 = ~n1330 & ~n1334;
  assign n1336 = ~pi138 & ~n1335;
  assign po117 = n1326 | n1336;
  assign n1338 = pi90 & n1115;
  assign n1339 = pi94 & n1186;
  assign n1340 = ~n1338 & ~n1339;
  assign n1341 = pi138 & ~n1340;
  assign n1342 = ~pi78 & ~pi136;
  assign n1343 = ~pi33 & pi136;
  assign n1344 = pi137 & ~n1342;
  assign n1345 = ~n1343 & n1344;
  assign n1346 = pi74 & ~pi136;
  assign n1347 = pi63 & pi136;
  assign n1348 = ~pi137 & ~n1346;
  assign n1349 = ~n1347 & n1348;
  assign n1350 = ~n1345 & ~n1349;
  assign n1351 = ~pi138 & ~n1350;
  assign po118 = n1341 | n1351;
  assign n1353 = pi99 & n1115;
  assign n1354 = ~pi112 & n1186;
  assign n1355 = ~n1353 & ~n1354;
  assign n1356 = pi138 & ~n1355;
  assign n1357 = pi73 & ~pi136;
  assign n1358 = pi68 & pi136;
  assign n1359 = ~pi137 & ~n1357;
  assign n1360 = ~n1358 & n1359;
  assign n1361 = ~pi84 & ~pi136;
  assign n1362 = ~pi32 & pi136;
  assign n1363 = pi137 & ~n1361;
  assign n1364 = ~n1362 & n1363;
  assign n1365 = ~n1360 & ~n1364;
  assign n1366 = ~pi138 & ~n1365;
  assign po119 = n1356 | n1366;
  assign n1368 = ~pi92 & pi138;
  assign n1369 = pi70 & ~pi138;
  assign n1370 = pi136 & ~n1368;
  assign n1371 = ~n1369 & n1370;
  assign n1372 = ~pi125 & pi138;
  assign n1373 = pi75 & ~pi138;
  assign n1374 = ~pi136 & ~n1372;
  assign n1375 = ~n1373 & n1374;
  assign n1376 = ~n1371 & ~n1375;
  assign n1377 = ~pi137 & ~n1376;
  assign n1378 = pi35 & n1218;
  assign n1379 = ~pi80 & ~pi138;
  assign n1380 = ~pi100 & pi138;
  assign n1381 = ~pi136 & ~n1379;
  assign n1382 = ~n1380 & n1381;
  assign n1383 = ~n1378 & ~n1382;
  assign n1384 = pi137 & ~n1383;
  assign po120 = n1377 | n1384;
  assign n1386 = ~pi26 & n678;
  assign n1387 = n1231 & n1386;
  assign n1388 = ~n689 & ~n1387;
  assign po121 = n335 & ~n1388;
  assign n1390 = ~pi98 & pi138;
  assign n1391 = pi71 & ~pi138;
  assign n1392 = pi136 & ~n1390;
  assign n1393 = ~n1391 & n1392;
  assign n1394 = ~pi23 & pi138;
  assign n1395 = pi76 & ~pi138;
  assign n1396 = ~pi136 & ~n1394;
  assign n1397 = ~n1395 & n1396;
  assign n1398 = ~n1393 & ~n1397;
  assign n1399 = ~pi137 & ~n1398;
  assign n1400 = pi36 & n1218;
  assign n1401 = ~pi81 & ~pi138;
  assign n1402 = ~pi97 & pi138;
  assign n1403 = ~pi136 & ~n1401;
  assign n1404 = ~n1402 & n1403;
  assign n1405 = ~n1400 & ~n1404;
  assign n1406 = pi137 & ~n1405;
  assign po122 = n1399 | n1406;
  assign n1408 = ~pi88 & pi138;
  assign n1409 = pi64 & ~pi138;
  assign n1410 = pi136 & ~n1408;
  assign n1411 = ~n1409 & n1410;
  assign n1412 = ~pi120 & pi138;
  assign n1413 = pi67 & ~pi138;
  assign n1414 = ~pi136 & ~n1412;
  assign n1415 = ~n1413 & n1414;
  assign n1416 = ~n1411 & ~n1415;
  assign n1417 = ~pi137 & ~n1416;
  assign n1418 = pi30 & n1218;
  assign n1419 = ~pi86 & ~pi138;
  assign n1420 = ~pi111 & pi138;
  assign n1421 = ~pi136 & ~n1419;
  assign n1422 = ~n1420 & n1421;
  assign n1423 = ~n1418 & ~n1422;
  assign n1424 = pi137 & ~n1423;
  assign po123 = n1417 | n1424;
  assign n1426 = ~pi26 & n648;
  assign n1427 = pi116 & n335;
  assign n1428 = ~n711 & n1427;
  assign po124 = ~n1426 & n1428;
  assign n1430 = ~pi97 & n672;
  assign n1431 = ~n749 & ~n1430;
  assign po125 = n1427 & ~n1431;
  assign n1433 = ~pi111 & ~n1272;
  assign n1434 = ~pi129 & n1117;
  assign n1435 = ~pi139 & n1272;
  assign n1436 = ~n1433 & n1434;
  assign po126 = ~n1435 & n1436;
  assign n1438 = ~pi141 & n1272;
  assign n1439 = pi112 & ~n1272;
  assign n1440 = n1434 & ~n1438;
  assign po127 = ~n1439 & n1440;
  assign n1442 = ~pi54 & pi113;
  assign n1443 = ~pi11 & ~pi22;
  assign n1444 = pi54 & n1443;
  assign n1445 = n335 & ~n1442;
  assign po128 = ~n1444 & n1445;
  assign n1447 = ~pi140 & n1272;
  assign n1448 = pi115 & ~n1272;
  assign n1449 = n1434 & ~n1447;
  assign po130 = ~n1448 & n1449;
  assign n1451 = ~pi4 & ~pi7;
  assign n1452 = ~pi9 & ~pi12;
  assign n1453 = n1451 & n1452;
  assign n1454 = pi54 & n335;
  assign po131 = ~n1453 & n1454;
  assign po132 = ~pi122 | pi129;
  assign n1457 = ~pi54 & pi118;
  assign n1458 = pi54 & ~pi59;
  assign n1459 = n499 & n1458;
  assign n1460 = ~n1457 & ~n1459;
  assign po133 = ~pi129 & ~n1460;
  assign po134 = ~pi129 & ~n641;
  assign n1463 = ~pi120 & n1278;
  assign n1464 = ~pi111 & ~pi129;
  assign po135 = ~n1463 & n1464;
  assign n1466 = pi81 & pi120;
  assign po136 = ~pi129 & n1466;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi57 & ~pi129;
  assign n1471 = ~pi96 & pi125;
  assign n1472 = ~pi3 & ~n1471;
  assign po140 = ~pi129 & ~n1472;
  assign n1474 = ~pi126 & pi132;
  assign po141 = pi133 & n1474;
  assign po12 = 1'b1;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
endmodule
