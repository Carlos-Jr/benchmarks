module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7  );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7;
  wire n137, n138, n139, n140, n141, n142, n143,
    n144, n145, n146, n147, n148, n149, n150,
    n151, n152, n153, n154, n155, n156, n157,
    n158, n159, n160, n161, n162, n163, n164,
    n165, n166, n167, n168, n169, n170, n171,
    n172, n173, n174, n175, n176, n177, n178,
    n179, n180, n181, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n340, n341, n342, n343, n344, n345, n346,
    n347, n348, n349, n350, n351, n352, n353,
    n354, n355, n356, n357, n358, n359, n360,
    n361, n362, n363, n364, n365, n366, n367,
    n368, n369, n370, n371, n372, n373, n374,
    n375, n376, n377, n378, n379, n380, n381,
    n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465,
    n466, n467, n468, n469, n470, n471, n472,
    n473, n474, n475, n476, n477, n478, n479,
    n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493,
    n494, n495, n496, n497, n498, n499, n500,
    n501, n502, n503, n504, n505, n506, n507,
    n508, n509, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n887, n888,
    n889, n890, n891, n892, n893, n894, n895,
    n896, n897, n898, n899, n900, n901, n902,
    n903, n904, n905, n906, n907, n908, n909,
    n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923,
    n924, n926, n927, n928, n929, n930, n931,
    n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n941, n942, n943, n944, n945,
    n946, n947, n948, n950, n951, n952, n953,
    n956, n957, n958, n959, n960, n961;
  assign n137 = pi126  & ~pi127 ;
  assign n138 = ~pi124  & ~n137;
  assign n139 = ~pi125  & pi127 ;
  assign n140 = pi125  & ~n137;
  assign n141 = ~n139 & ~n140;
  assign n142 = pi124  & ~n141;
  assign n143 = ~n138 & ~n142;
  assign n144 = ~pi122  & ~n143;
  assign n145 = ~pi123  & ~n141;
  assign n146 = pi123  & ~n143;
  assign n147 = ~n145 & ~n146;
  assign n148 = pi122  & ~n147;
  assign n149 = ~n144 & ~n148;
  assign n150 = ~pi120  & ~n149;
  assign n151 = ~pi121  & ~n147;
  assign n152 = pi121  & ~n149;
  assign n153 = ~n151 & ~n152;
  assign n154 = pi120  & ~n153;
  assign n155 = ~n150 & ~n154;
  assign n156 = ~pi118  & ~n155;
  assign n157 = ~pi119  & ~n153;
  assign n158 = pi119  & ~n155;
  assign n159 = ~n157 & ~n158;
  assign n160 = pi118  & ~n159;
  assign n161 = ~n156 & ~n160;
  assign n162 = ~pi116  & ~n161;
  assign n163 = ~pi117  & ~n159;
  assign n164 = pi117  & ~n161;
  assign n165 = ~n163 & ~n164;
  assign n166 = pi116  & ~n165;
  assign n167 = ~n162 & ~n166;
  assign n168 = ~pi114  & ~n167;
  assign n169 = ~pi115  & ~n165;
  assign n170 = pi115  & ~n167;
  assign n171 = ~n169 & ~n170;
  assign n172 = pi114  & ~n171;
  assign n173 = ~n168 & ~n172;
  assign n174 = ~pi112  & ~n173;
  assign n175 = ~pi113  & ~n171;
  assign n176 = pi113  & ~n173;
  assign n177 = ~n175 & ~n176;
  assign n178 = pi112  & ~n177;
  assign n179 = ~n174 & ~n178;
  assign n180 = ~pi110  & ~n179;
  assign n181 = ~pi111  & ~n177;
  assign n182 = pi111  & ~n179;
  assign n183 = ~n181 & ~n182;
  assign n184 = pi110  & ~n183;
  assign n185 = ~n180 & ~n184;
  assign n186 = ~pi108  & ~n185;
  assign n187 = ~pi109  & ~n183;
  assign n188 = pi109  & ~n185;
  assign n189 = ~n187 & ~n188;
  assign n190 = pi108  & ~n189;
  assign n191 = ~n186 & ~n190;
  assign n192 = ~pi106  & ~n191;
  assign n193 = ~pi107  & ~n189;
  assign n194 = pi107  & ~n191;
  assign n195 = ~n193 & ~n194;
  assign n196 = pi106  & ~n195;
  assign n197 = ~n192 & ~n196;
  assign n198 = ~pi104  & ~n197;
  assign n199 = ~pi105  & ~n195;
  assign n200 = pi105  & ~n197;
  assign n201 = ~n199 & ~n200;
  assign n202 = pi104  & ~n201;
  assign n203 = ~n198 & ~n202;
  assign n204 = ~pi102  & ~n203;
  assign n205 = ~pi103  & ~n201;
  assign n206 = pi103  & ~n203;
  assign n207 = ~n205 & ~n206;
  assign n208 = pi102  & ~n207;
  assign n209 = ~n204 & ~n208;
  assign n210 = ~pi100  & ~n209;
  assign n211 = ~pi101  & ~n207;
  assign n212 = pi101  & ~n209;
  assign n213 = ~n211 & ~n212;
  assign n214 = pi100  & ~n213;
  assign n215 = ~n210 & ~n214;
  assign n216 = ~pi98  & ~n215;
  assign n217 = ~pi99  & ~n213;
  assign n218 = pi99  & ~n215;
  assign n219 = ~n217 & ~n218;
  assign n220 = pi98  & ~n219;
  assign n221 = ~n216 & ~n220;
  assign n222 = ~pi96  & ~n221;
  assign n223 = ~pi97  & ~n219;
  assign n224 = pi97  & ~n221;
  assign n225 = ~n223 & ~n224;
  assign n226 = pi96  & ~n225;
  assign n227 = ~n222 & ~n226;
  assign n228 = ~pi94  & ~n227;
  assign n229 = ~pi95  & ~n225;
  assign n230 = pi95  & ~n227;
  assign n231 = ~n229 & ~n230;
  assign n232 = pi94  & ~n231;
  assign n233 = ~n228 & ~n232;
  assign n234 = ~pi92  & ~n233;
  assign n235 = ~pi93  & ~n231;
  assign n236 = pi93  & ~n233;
  assign n237 = ~n235 & ~n236;
  assign n238 = pi92  & ~n237;
  assign n239 = ~n234 & ~n238;
  assign n240 = ~pi90  & ~n239;
  assign n241 = ~pi91  & ~n237;
  assign n242 = pi91  & ~n239;
  assign n243 = ~n241 & ~n242;
  assign n244 = pi90  & ~n243;
  assign n245 = ~n240 & ~n244;
  assign n246 = ~pi88  & ~n245;
  assign n247 = ~pi89  & ~n243;
  assign n248 = pi89  & ~n245;
  assign n249 = ~n247 & ~n248;
  assign n250 = pi88  & ~n249;
  assign n251 = ~n246 & ~n250;
  assign n252 = ~pi86  & ~n251;
  assign n253 = ~pi87  & ~n249;
  assign n254 = pi87  & ~n251;
  assign n255 = ~n253 & ~n254;
  assign n256 = pi86  & ~n255;
  assign n257 = ~n252 & ~n256;
  assign n258 = ~pi84  & ~n257;
  assign n259 = ~pi85  & ~n255;
  assign n260 = pi85  & ~n257;
  assign n261 = ~n259 & ~n260;
  assign n262 = pi84  & ~n261;
  assign n263 = ~n258 & ~n262;
  assign n264 = ~pi82  & ~n263;
  assign n265 = ~pi83  & ~n261;
  assign n266 = pi83  & ~n263;
  assign n267 = ~n265 & ~n266;
  assign n268 = pi82  & ~n267;
  assign n269 = ~n264 & ~n268;
  assign n270 = ~pi80  & ~n269;
  assign n271 = ~pi81  & ~n267;
  assign n272 = pi81  & ~n269;
  assign n273 = ~n271 & ~n272;
  assign n274 = pi80  & ~n273;
  assign n275 = ~n270 & ~n274;
  assign n276 = ~pi78  & ~n275;
  assign n277 = ~pi79  & ~n273;
  assign n278 = pi79  & ~n275;
  assign n279 = ~n277 & ~n278;
  assign n280 = pi78  & ~n279;
  assign n281 = ~n276 & ~n280;
  assign n282 = ~pi76  & ~n281;
  assign n283 = ~pi77  & ~n279;
  assign n284 = pi77  & ~n281;
  assign n285 = ~n283 & ~n284;
  assign n286 = pi76  & ~n285;
  assign n287 = ~n282 & ~n286;
  assign n288 = ~pi74  & ~n287;
  assign n289 = ~pi75  & ~n285;
  assign n290 = pi75  & ~n287;
  assign n291 = ~n289 & ~n290;
  assign n292 = pi74  & ~n291;
  assign n293 = ~n288 & ~n292;
  assign n294 = ~pi72  & ~n293;
  assign n295 = ~pi73  & ~n291;
  assign n296 = pi73  & ~n293;
  assign n297 = ~n295 & ~n296;
  assign n298 = pi72  & ~n297;
  assign n299 = ~n294 & ~n298;
  assign n300 = ~pi70  & ~n299;
  assign n301 = ~pi71  & ~n297;
  assign n302 = pi71  & ~n299;
  assign n303 = ~n301 & ~n302;
  assign n304 = pi70  & ~n303;
  assign n305 = ~n300 & ~n304;
  assign n306 = ~pi68  & ~n305;
  assign n307 = ~pi69  & ~n303;
  assign n308 = pi69  & ~n305;
  assign n309 = ~n307 & ~n308;
  assign n310 = pi68  & ~n309;
  assign n311 = ~n306 & ~n310;
  assign n312 = ~pi66  & ~n311;
  assign n313 = ~pi67  & ~n309;
  assign n314 = pi67  & ~n311;
  assign n315 = ~n313 & ~n314;
  assign n316 = pi66  & ~n315;
  assign n317 = ~n312 & ~n316;
  assign n318 = ~pi64  & ~n317;
  assign n319 = ~pi65  & ~n315;
  assign n320 = pi65  & ~n317;
  assign n321 = ~n319 & ~n320;
  assign n322 = pi64  & ~n321;
  assign n323 = ~n318 & ~n322;
  assign n324 = ~pi62  & ~n323;
  assign n325 = ~pi63  & ~n321;
  assign n326 = pi63  & ~n323;
  assign n327 = ~n325 & ~n326;
  assign n328 = pi62  & ~n327;
  assign n329 = ~n324 & ~n328;
  assign n330 = ~pi60  & ~n329;
  assign n331 = ~pi61  & ~n327;
  assign n332 = pi61  & ~n329;
  assign n333 = ~n331 & ~n332;
  assign n334 = pi60  & ~n333;
  assign n335 = ~n330 & ~n334;
  assign n336 = ~pi58  & ~n335;
  assign n337 = ~pi59  & ~n333;
  assign n338 = pi59  & ~n335;
  assign n339 = ~n337 & ~n338;
  assign n340 = pi58  & ~n339;
  assign n341 = ~n336 & ~n340;
  assign n342 = ~pi56  & ~n341;
  assign n343 = ~pi57  & ~n339;
  assign n344 = pi57  & ~n341;
  assign n345 = ~n343 & ~n344;
  assign n346 = pi56  & ~n345;
  assign n347 = ~n342 & ~n346;
  assign n348 = ~pi54  & ~n347;
  assign n349 = ~pi55  & ~n345;
  assign n350 = pi55  & ~n347;
  assign n351 = ~n349 & ~n350;
  assign n352 = pi54  & ~n351;
  assign n353 = ~n348 & ~n352;
  assign n354 = ~pi52  & ~n353;
  assign n355 = ~pi53  & ~n351;
  assign n356 = pi53  & ~n353;
  assign n357 = ~n355 & ~n356;
  assign n358 = pi52  & ~n357;
  assign n359 = ~n354 & ~n358;
  assign n360 = ~pi50  & ~n359;
  assign n361 = ~pi51  & ~n357;
  assign n362 = pi51  & ~n359;
  assign n363 = ~n361 & ~n362;
  assign n364 = pi50  & ~n363;
  assign n365 = ~n360 & ~n364;
  assign n366 = ~pi48  & ~n365;
  assign n367 = ~pi49  & ~n363;
  assign n368 = pi49  & ~n365;
  assign n369 = ~n367 & ~n368;
  assign n370 = pi48  & ~n369;
  assign n371 = ~n366 & ~n370;
  assign n372 = ~pi46  & ~n371;
  assign n373 = ~pi47  & ~n369;
  assign n374 = pi47  & ~n371;
  assign n375 = ~n373 & ~n374;
  assign n376 = pi46  & ~n375;
  assign n377 = ~n372 & ~n376;
  assign n378 = ~pi44  & ~n377;
  assign n379 = ~pi45  & ~n375;
  assign n380 = pi45  & ~n377;
  assign n381 = ~n379 & ~n380;
  assign n382 = pi44  & ~n381;
  assign n383 = ~n378 & ~n382;
  assign n384 = ~pi42  & ~n383;
  assign n385 = ~pi43  & ~n381;
  assign n386 = pi43  & ~n383;
  assign n387 = ~n385 & ~n386;
  assign n388 = pi42  & ~n387;
  assign n389 = ~n384 & ~n388;
  assign n390 = ~pi40  & ~n389;
  assign n391 = ~pi41  & ~n387;
  assign n392 = pi41  & ~n389;
  assign n393 = ~n391 & ~n392;
  assign n394 = pi40  & ~n393;
  assign n395 = ~n390 & ~n394;
  assign n396 = ~pi38  & ~n395;
  assign n397 = ~pi39  & ~n393;
  assign n398 = pi39  & ~n395;
  assign n399 = ~n397 & ~n398;
  assign n400 = pi38  & ~n399;
  assign n401 = ~n396 & ~n400;
  assign n402 = ~pi36  & ~n401;
  assign n403 = ~pi37  & ~n399;
  assign n404 = pi37  & ~n401;
  assign n405 = ~n403 & ~n404;
  assign n406 = pi36  & ~n405;
  assign n407 = ~n402 & ~n406;
  assign n408 = ~pi34  & ~n407;
  assign n409 = ~pi35  & ~n405;
  assign n410 = pi35  & ~n407;
  assign n411 = ~n409 & ~n410;
  assign n412 = pi34  & ~n411;
  assign n413 = ~n408 & ~n412;
  assign n414 = ~pi32  & ~n413;
  assign n415 = ~pi33  & ~n411;
  assign n416 = pi33  & ~n413;
  assign n417 = ~n415 & ~n416;
  assign n418 = pi32  & ~n417;
  assign n419 = ~n414 & ~n418;
  assign n420 = ~pi30  & ~n419;
  assign n421 = ~pi31  & ~n417;
  assign n422 = pi31  & ~n419;
  assign n423 = ~n421 & ~n422;
  assign n424 = pi30  & ~n423;
  assign n425 = ~n420 & ~n424;
  assign n426 = ~pi28  & ~n425;
  assign n427 = ~pi29  & ~n423;
  assign n428 = pi29  & ~n425;
  assign n429 = ~n427 & ~n428;
  assign n430 = pi28  & ~n429;
  assign n431 = ~n426 & ~n430;
  assign n432 = ~pi26  & ~n431;
  assign n433 = ~pi27  & ~n429;
  assign n434 = pi27  & ~n431;
  assign n435 = ~n433 & ~n434;
  assign n436 = pi26  & ~n435;
  assign n437 = ~n432 & ~n436;
  assign n438 = ~pi24  & ~n437;
  assign n439 = ~pi25  & ~n435;
  assign n440 = pi25  & ~n437;
  assign n441 = ~n439 & ~n440;
  assign n442 = pi24  & ~n441;
  assign n443 = ~n438 & ~n442;
  assign n444 = ~pi22  & ~n443;
  assign n445 = ~pi23  & ~n441;
  assign n446 = pi23  & ~n443;
  assign n447 = ~n445 & ~n446;
  assign n448 = pi22  & ~n447;
  assign n449 = ~n444 & ~n448;
  assign n450 = ~pi20  & ~n449;
  assign n451 = ~pi21  & ~n447;
  assign n452 = pi21  & ~n449;
  assign n453 = ~n451 & ~n452;
  assign n454 = pi20  & ~n453;
  assign n455 = ~n450 & ~n454;
  assign n456 = ~pi18  & ~n455;
  assign n457 = ~pi19  & ~n453;
  assign n458 = pi19  & ~n455;
  assign n459 = ~n457 & ~n458;
  assign n460 = pi18  & ~n459;
  assign n461 = ~n456 & ~n460;
  assign n462 = ~pi16  & ~n461;
  assign n463 = ~pi17  & ~n459;
  assign n464 = pi17  & ~n461;
  assign n465 = ~n463 & ~n464;
  assign n466 = pi16  & ~n465;
  assign n467 = ~n462 & ~n466;
  assign n468 = ~pi14  & ~n467;
  assign n469 = ~pi15  & ~n465;
  assign n470 = pi15  & ~n467;
  assign n471 = ~n469 & ~n470;
  assign n472 = pi14  & ~n471;
  assign n473 = ~n468 & ~n472;
  assign n474 = ~pi12  & ~n473;
  assign n475 = ~pi13  & ~n471;
  assign n476 = pi13  & ~n473;
  assign n477 = ~n475 & ~n476;
  assign n478 = pi12  & ~n477;
  assign n479 = ~n474 & ~n478;
  assign n480 = ~pi10  & ~n479;
  assign n481 = ~pi11  & ~n477;
  assign n482 = pi11  & ~n479;
  assign n483 = ~n481 & ~n482;
  assign n484 = pi10  & ~n483;
  assign n485 = ~n480 & ~n484;
  assign n486 = ~pi8  & ~n485;
  assign n487 = ~pi9  & ~n483;
  assign n488 = pi9  & ~n485;
  assign n489 = ~n487 & ~n488;
  assign n490 = pi8  & ~n489;
  assign n491 = ~n486 & ~n490;
  assign n492 = ~pi6  & ~n491;
  assign n493 = ~pi7  & ~n489;
  assign n494 = pi7  & ~n491;
  assign n495 = ~n493 & ~n494;
  assign n496 = pi6  & ~n495;
  assign n497 = ~n492 & ~n496;
  assign n498 = ~pi4  & ~n497;
  assign n499 = ~pi5  & ~n495;
  assign n500 = pi5  & ~n497;
  assign n501 = ~n499 & ~n500;
  assign n502 = pi4  & ~n501;
  assign n503 = ~n498 & ~n502;
  assign n504 = pi3  & ~n503;
  assign n505 = ~pi3  & ~n501;
  assign n506 = pi1  & ~pi2 ;
  assign n507 = ~n505 & ~n506;
  assign n508 = ~n504 & n507;
  assign n509 = n503 & n506;
  assign po0  = ~n508 & ~n509;
  assign n511 = ~pi110  & ~pi111 ;
  assign n512 = ~pi118  & ~pi119 ;
  assign n513 = ~pi126  & ~pi127 ;
  assign n514 = ~pi124  & ~pi125 ;
  assign n515 = ~pi122  & ~pi123 ;
  assign n516 = n514 & ~n515;
  assign n517 = n513 & ~n516;
  assign n518 = n513 & n514;
  assign n519 = ~pi120  & ~pi121 ;
  assign n520 = n515 & n519;
  assign n521 = n518 & n520;
  assign n522 = n517 & ~n521;
  assign n523 = ~n512 & n522;
  assign n524 = n512 & n517;
  assign n525 = ~n523 & ~n524;
  assign n526 = ~pi116  & ~pi117 ;
  assign n527 = n525 & ~n526;
  assign n528 = ~n522 & n526;
  assign n529 = ~pi114  & ~pi115 ;
  assign n530 = ~n528 & ~n529;
  assign n531 = ~n527 & n530;
  assign n532 = ~n525 & n529;
  assign n533 = ~n531 & ~n532;
  assign n534 = n512 & n526;
  assign n535 = ~pi112  & ~pi113 ;
  assign n536 = n529 & n535;
  assign n537 = n534 & n536;
  assign n538 = n521 & n537;
  assign n539 = ~n533 & ~n538;
  assign n540 = ~n511 & n539;
  assign n541 = n511 & ~n533;
  assign n542 = ~n540 & ~n541;
  assign n543 = ~pi108  & ~pi109 ;
  assign n544 = n542 & ~n543;
  assign n545 = ~n539 & n543;
  assign n546 = ~n544 & ~n545;
  assign n547 = ~pi106  & ~pi107 ;
  assign n548 = n546 & ~n547;
  assign n549 = ~n542 & n547;
  assign n550 = ~n548 & ~n549;
  assign n551 = ~pi104  & ~pi105 ;
  assign n552 = n550 & ~n551;
  assign n553 = ~n546 & n551;
  assign n554 = ~n552 & ~n553;
  assign n555 = ~pi102  & ~pi103 ;
  assign n556 = n554 & ~n555;
  assign n557 = ~n550 & n555;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~pi100  & ~pi101 ;
  assign n560 = n558 & ~n559;
  assign n561 = ~n554 & n559;
  assign n562 = ~n560 & ~n561;
  assign n563 = ~pi98  & ~pi99 ;
  assign n564 = n562 & ~n563;
  assign n565 = ~n558 & n563;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~pi96  & ~pi97 ;
  assign n568 = n566 & ~n567;
  assign n569 = ~n562 & n567;
  assign n570 = ~n568 & ~n569;
  assign n571 = ~pi94  & ~pi95 ;
  assign n572 = n570 & ~n571;
  assign n573 = ~n566 & n571;
  assign n574 = ~n572 & ~n573;
  assign n575 = ~pi92  & ~pi93 ;
  assign n576 = n574 & ~n575;
  assign n577 = ~n570 & n575;
  assign n578 = ~n576 & ~n577;
  assign n579 = ~pi90  & ~pi91 ;
  assign n580 = n578 & ~n579;
  assign n581 = ~n574 & n579;
  assign n582 = ~n580 & ~n581;
  assign n583 = ~pi88  & ~pi89 ;
  assign n584 = n582 & ~n583;
  assign n585 = ~n578 & n583;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~pi86  & ~pi87 ;
  assign n588 = n586 & ~n587;
  assign n589 = ~n582 & n587;
  assign n590 = ~n588 & ~n589;
  assign n591 = ~pi84  & ~pi85 ;
  assign n592 = n590 & ~n591;
  assign n593 = ~n586 & n591;
  assign n594 = ~n592 & ~n593;
  assign n595 = ~pi82  & ~pi83 ;
  assign n596 = n594 & ~n595;
  assign n597 = ~n590 & n595;
  assign n598 = ~n596 & ~n597;
  assign n599 = ~pi80  & ~pi81 ;
  assign n600 = n598 & ~n599;
  assign n601 = ~n594 & n599;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~pi78  & ~pi79 ;
  assign n604 = n602 & ~n603;
  assign n605 = ~n598 & n603;
  assign n606 = ~n604 & ~n605;
  assign n607 = ~pi76  & ~pi77 ;
  assign n608 = n606 & ~n607;
  assign n609 = ~n602 & n607;
  assign n610 = ~n608 & ~n609;
  assign n611 = ~pi74  & ~pi75 ;
  assign n612 = n610 & ~n611;
  assign n613 = ~n606 & n611;
  assign n614 = ~n612 & ~n613;
  assign n615 = ~pi72  & ~pi73 ;
  assign n616 = n614 & ~n615;
  assign n617 = ~n610 & n615;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~pi70  & ~pi71 ;
  assign n620 = n618 & ~n619;
  assign n621 = ~n614 & n619;
  assign n622 = ~n620 & ~n621;
  assign n623 = ~pi68  & ~pi69 ;
  assign n624 = n622 & ~n623;
  assign n625 = ~n618 & n623;
  assign n626 = ~n624 & ~n625;
  assign n627 = ~pi66  & ~pi67 ;
  assign n628 = n626 & ~n627;
  assign n629 = ~n622 & n627;
  assign n630 = ~n628 & ~n629;
  assign n631 = ~pi64  & ~pi65 ;
  assign n632 = n630 & ~n631;
  assign n633 = ~n626 & n631;
  assign n634 = ~n632 & ~n633;
  assign n635 = ~pi62  & ~pi63 ;
  assign n636 = n634 & ~n635;
  assign n637 = ~n630 & n635;
  assign n638 = ~n636 & ~n637;
  assign n639 = ~pi60  & ~pi61 ;
  assign n640 = n638 & ~n639;
  assign n641 = ~n634 & n639;
  assign n642 = ~n640 & ~n641;
  assign n643 = ~pi58  & ~pi59 ;
  assign n644 = n642 & ~n643;
  assign n645 = ~n638 & n643;
  assign n646 = ~n644 & ~n645;
  assign n647 = ~pi56  & ~pi57 ;
  assign n648 = n646 & ~n647;
  assign n649 = ~n642 & n647;
  assign n650 = ~n648 & ~n649;
  assign n651 = ~pi54  & ~pi55 ;
  assign n652 = n650 & ~n651;
  assign n653 = ~n646 & n651;
  assign n654 = ~n652 & ~n653;
  assign n655 = ~pi52  & ~pi53 ;
  assign n656 = n654 & ~n655;
  assign n657 = ~n650 & n655;
  assign n658 = ~n656 & ~n657;
  assign n659 = ~pi50  & ~pi51 ;
  assign n660 = n658 & ~n659;
  assign n661 = ~n654 & n659;
  assign n662 = ~n660 & ~n661;
  assign n663 = ~pi48  & ~pi49 ;
  assign n664 = n662 & ~n663;
  assign n665 = ~n658 & n663;
  assign n666 = ~n664 & ~n665;
  assign n667 = ~pi46  & ~pi47 ;
  assign n668 = n666 & ~n667;
  assign n669 = ~n662 & n667;
  assign n670 = ~n668 & ~n669;
  assign n671 = ~pi44  & ~pi45 ;
  assign n672 = n670 & ~n671;
  assign n673 = ~n666 & n671;
  assign n674 = ~n672 & ~n673;
  assign n675 = ~pi42  & ~pi43 ;
  assign n676 = n674 & ~n675;
  assign n677 = ~n670 & n675;
  assign n678 = ~n676 & ~n677;
  assign n679 = ~pi40  & ~pi41 ;
  assign n680 = n678 & ~n679;
  assign n681 = ~n674 & n679;
  assign n682 = ~n680 & ~n681;
  assign n683 = ~pi38  & ~pi39 ;
  assign n684 = n682 & ~n683;
  assign n685 = ~n678 & n683;
  assign n686 = ~n684 & ~n685;
  assign n687 = ~pi36  & ~pi37 ;
  assign n688 = n686 & ~n687;
  assign n689 = ~n682 & n687;
  assign n690 = ~n688 & ~n689;
  assign n691 = ~pi34  & ~pi35 ;
  assign n692 = n690 & ~n691;
  assign n693 = ~n686 & n691;
  assign n694 = ~n692 & ~n693;
  assign n695 = ~pi32  & ~pi33 ;
  assign n696 = n694 & ~n695;
  assign n697 = ~n690 & n695;
  assign n698 = ~n696 & ~n697;
  assign n699 = ~pi30  & ~pi31 ;
  assign n700 = n698 & ~n699;
  assign n701 = ~n694 & n699;
  assign n702 = ~n700 & ~n701;
  assign n703 = ~pi28  & ~pi29 ;
  assign n704 = n702 & ~n703;
  assign n705 = ~n698 & n703;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~pi26  & ~pi27 ;
  assign n708 = n706 & ~n707;
  assign n709 = ~n702 & n707;
  assign n710 = ~n708 & ~n709;
  assign n711 = ~pi24  & ~pi25 ;
  assign n712 = n710 & ~n711;
  assign n713 = ~n706 & n711;
  assign n714 = ~n712 & ~n713;
  assign n715 = ~pi22  & ~pi23 ;
  assign n716 = n714 & ~n715;
  assign n717 = ~n710 & n715;
  assign n718 = ~n716 & ~n717;
  assign n719 = ~pi20  & ~pi21 ;
  assign n720 = n718 & ~n719;
  assign n721 = ~n714 & n719;
  assign n722 = ~n720 & ~n721;
  assign n723 = ~pi18  & ~pi19 ;
  assign n724 = n722 & ~n723;
  assign n725 = ~n718 & n723;
  assign n726 = ~n724 & ~n725;
  assign n727 = ~pi16  & ~pi17 ;
  assign n728 = n726 & ~n727;
  assign n729 = ~n722 & n727;
  assign n730 = ~n728 & ~n729;
  assign n731 = ~pi14  & ~pi15 ;
  assign n732 = n730 & ~n731;
  assign n733 = ~n726 & n731;
  assign n734 = ~n732 & ~n733;
  assign n735 = ~pi12  & ~pi13 ;
  assign n736 = n734 & ~n735;
  assign n737 = ~n730 & n735;
  assign n738 = ~n736 & ~n737;
  assign n739 = ~pi10  & ~pi11 ;
  assign n740 = n738 & ~n739;
  assign n741 = ~n734 & n739;
  assign n742 = ~n740 & ~n741;
  assign n743 = ~pi8  & ~pi9 ;
  assign n744 = n742 & ~n743;
  assign n745 = ~n738 & n743;
  assign n746 = ~n744 & ~n745;
  assign n747 = ~pi6  & ~pi7 ;
  assign n748 = n746 & ~n747;
  assign n749 = ~n742 & n747;
  assign n750 = ~n748 & ~n749;
  assign n751 = ~pi4  & ~pi5 ;
  assign n752 = n750 & ~n751;
  assign n753 = ~n746 & n751;
  assign n754 = ~pi2  & ~pi3 ;
  assign n755 = ~n753 & ~n754;
  assign n756 = ~n752 & n755;
  assign n757 = ~n750 & n754;
  assign po1  = ~n756 & ~n757;
  assign n759 = n571 & n575;
  assign n760 = n511 & n543;
  assign n761 = n520 & ~n534;
  assign n762 = n518 & ~n761;
  assign n763 = ~n538 & n762;
  assign n764 = ~n760 & ~n763;
  assign n765 = n760 & ~n762;
  assign n766 = ~n764 & ~n765;
  assign n767 = n547 & n551;
  assign n768 = n766 & ~n767;
  assign n769 = n763 & n767;
  assign n770 = n555 & n559;
  assign n771 = ~n769 & ~n770;
  assign n772 = ~n768 & n771;
  assign n773 = ~n766 & n770;
  assign n774 = ~n772 & ~n773;
  assign n775 = n760 & n767;
  assign n776 = n563 & n567;
  assign n777 = n770 & n776;
  assign n778 = n775 & n777;
  assign n779 = n538 & n778;
  assign n780 = n774 & ~n779;
  assign n781 = ~n759 & ~n780;
  assign n782 = n759 & ~n774;
  assign n783 = ~n781 & ~n782;
  assign n784 = n579 & n583;
  assign n785 = n783 & ~n784;
  assign n786 = n780 & n784;
  assign n787 = ~n785 & ~n786;
  assign n788 = n587 & n591;
  assign n789 = n787 & ~n788;
  assign n790 = ~n783 & n788;
  assign n791 = ~n789 & ~n790;
  assign n792 = n595 & n599;
  assign n793 = n791 & ~n792;
  assign n794 = ~n787 & n792;
  assign n795 = ~n793 & ~n794;
  assign n796 = n603 & n607;
  assign n797 = n795 & ~n796;
  assign n798 = ~n791 & n796;
  assign n799 = ~n797 & ~n798;
  assign n800 = n611 & n615;
  assign n801 = n799 & ~n800;
  assign n802 = ~n795 & n800;
  assign n803 = ~n801 & ~n802;
  assign n804 = n619 & n623;
  assign n805 = n803 & ~n804;
  assign n806 = ~n799 & n804;
  assign n807 = ~n805 & ~n806;
  assign n808 = n627 & n631;
  assign n809 = n807 & ~n808;
  assign n810 = ~n803 & n808;
  assign n811 = ~n809 & ~n810;
  assign n812 = n635 & n639;
  assign n813 = n811 & ~n812;
  assign n814 = ~n807 & n812;
  assign n815 = ~n813 & ~n814;
  assign n816 = n643 & n647;
  assign n817 = n815 & ~n816;
  assign n818 = ~n811 & n816;
  assign n819 = ~n817 & ~n818;
  assign n820 = n651 & n655;
  assign n821 = n819 & ~n820;
  assign n822 = ~n815 & n820;
  assign n823 = ~n821 & ~n822;
  assign n824 = n659 & n663;
  assign n825 = n823 & ~n824;
  assign n826 = ~n819 & n824;
  assign n827 = ~n825 & ~n826;
  assign n828 = n667 & n671;
  assign n829 = n827 & ~n828;
  assign n830 = ~n823 & n828;
  assign n831 = ~n829 & ~n830;
  assign n832 = n675 & n679;
  assign n833 = n831 & ~n832;
  assign n834 = ~n827 & n832;
  assign n835 = ~n833 & ~n834;
  assign n836 = n683 & n687;
  assign n837 = n835 & ~n836;
  assign n838 = ~n831 & n836;
  assign n839 = ~n837 & ~n838;
  assign n840 = n691 & n695;
  assign n841 = n839 & ~n840;
  assign n842 = ~n835 & n840;
  assign n843 = ~n841 & ~n842;
  assign n844 = n699 & n703;
  assign n845 = n843 & ~n844;
  assign n846 = ~n839 & n844;
  assign n847 = ~n845 & ~n846;
  assign n848 = n707 & n711;
  assign n849 = n847 & ~n848;
  assign n850 = ~n843 & n848;
  assign n851 = ~n849 & ~n850;
  assign n852 = n715 & n719;
  assign n853 = n851 & ~n852;
  assign n854 = ~n847 & n852;
  assign n855 = ~n853 & ~n854;
  assign n856 = n723 & n727;
  assign n857 = n855 & ~n856;
  assign n858 = ~n851 & n856;
  assign n859 = ~n857 & ~n858;
  assign n860 = n731 & n735;
  assign n861 = n859 & ~n860;
  assign n862 = ~n855 & n860;
  assign n863 = ~n861 & ~n862;
  assign n864 = n739 & n743;
  assign n865 = n863 & ~n864;
  assign n866 = ~n859 & n864;
  assign n867 = n747 & n751;
  assign n868 = ~n866 & ~n867;
  assign n869 = ~n865 & n868;
  assign n870 = ~n863 & n867;
  assign po2  = n869 | n870;
  assign n872 = n537 & ~n775;
  assign n873 = n521 & ~n872;
  assign n874 = ~pi102  & n559;
  assign n875 = n776 & n874;
  assign n876 = n873 & ~n875;
  assign n877 = pi103  & n775;
  assign n878 = n537 & ~n877;
  assign n879 = n521 & n875;
  assign n880 = ~n878 & n879;
  assign n881 = ~n876 & ~n880;
  assign n882 = n759 & n784;
  assign n883 = n881 & ~n882;
  assign n884 = ~n873 & n882;
  assign n885 = ~n883 & ~n884;
  assign n886 = n788 & n792;
  assign n887 = n885 & ~n886;
  assign n888 = ~n881 & n886;
  assign n889 = ~n887 & ~n888;
  assign n890 = n796 & n800;
  assign n891 = n889 & ~n890;
  assign n892 = ~n885 & n890;
  assign n893 = ~n891 & ~n892;
  assign n894 = n804 & n808;
  assign n895 = n893 & ~n894;
  assign n896 = ~n889 & n894;
  assign n897 = ~n895 & ~n896;
  assign n898 = n812 & n816;
  assign n899 = n897 & ~n898;
  assign n900 = ~n893 & n898;
  assign n901 = ~n899 & ~n900;
  assign n902 = n820 & n824;
  assign n903 = n901 & ~n902;
  assign n904 = ~n897 & n902;
  assign n905 = ~n903 & ~n904;
  assign n906 = n828 & n832;
  assign n907 = n905 & ~n906;
  assign n908 = ~n901 & n906;
  assign n909 = ~n907 & ~n908;
  assign n910 = n836 & n840;
  assign n911 = n909 & ~n910;
  assign n912 = ~n905 & n910;
  assign n913 = ~n911 & ~n912;
  assign n914 = n844 & n848;
  assign n915 = n913 & ~n914;
  assign n916 = ~n909 & n914;
  assign n917 = ~n915 & ~n916;
  assign n918 = n852 & n856;
  assign n919 = n917 & ~n918;
  assign n920 = ~n913 & n918;
  assign n921 = n860 & n864;
  assign n922 = ~n920 & ~n921;
  assign n923 = ~n919 & n922;
  assign n924 = ~n917 & n921;
  assign po3  = n923 | n924;
  assign n926 = n882 & n886;
  assign n927 = n778 & ~n926;
  assign n928 = n538 & ~n927;
  assign n929 = ~pi78  & n607;
  assign n930 = n800 & n929;
  assign n931 = n894 & n930;
  assign n932 = n928 & ~n931;
  assign n933 = pi79  & n926;
  assign n934 = n778 & ~n933;
  assign n935 = n538 & n931;
  assign n936 = ~n934 & n935;
  assign n937 = ~n932 & ~n936;
  assign n938 = n898 & n902;
  assign n939 = n937 & ~n938;
  assign n940 = ~n928 & n938;
  assign n941 = ~n939 & ~n940;
  assign n942 = n906 & n910;
  assign n943 = n941 & ~n942;
  assign n944 = ~n937 & n942;
  assign n945 = n914 & n918;
  assign n946 = ~n944 & ~n945;
  assign n947 = ~n943 & n946;
  assign n948 = ~n941 & n945;
  assign po4  = n947 | n948;
  assign n950 = n890 & n894;
  assign n951 = n926 & n950;
  assign n952 = n938 & n942;
  assign n953 = n951 & ~n952;
  assign po5  = ~n779 | n953;
  assign po6  = ~n779 | ~n951;
  assign n956 = ~pi0  & ~pi1 ;
  assign n957 = n754 & n956;
  assign n958 = n867 & n957;
  assign n959 = n921 & n958;
  assign n960 = n945 & n959;
  assign n961 = n952 & n960;
  assign po7 = po6  | ~n961;
endmodule
