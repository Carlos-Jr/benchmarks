module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 , pi73 ,
    pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 , pi81 ,
    pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 , pi89 ,
    pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 , pi97 ,
    pi98 , pi99 , pi100 , pi101 , pi102 , pi103 , pi104 , pi105 ,
    pi106 , pi107 , pi108 , pi109 , pi110 , pi111 , pi112 , pi113 ,
    pi114 , pi115 , pi116 , pi117 , pi118 , pi119 , pi120 , pi121 ,
    pi122 , pi123 , pi124 , pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 , po8 ,
    po9 , po10 , po11 , po12 , po13 , po14 , po15 , po16 ,
    po17 , po18 , po19 , po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 , po30 , po31 , po32 ,
    po33 , po34 , po35 , po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 , po46 , po47 , po48 ,
    po49 , po50 , po51 , po52 , po53 , po54 , po55 , po56 ,
    po57 , po58 , po59 , po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 , po70 , po71 , po72 ,
    po73 , po74 , po75 , po76 , po77 , po78 , po79 , po80 ,
    po81 , po82 , po83 , po84 , po85 , po86 , po87 , po88 ,
    po89 , po90 , po91 , po92 , po93 , po94 , po95 , po96 ,
    po97 , po98 , po99 , po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 , po108 , po109 , po110 ,
    po111 , po112 , po113 , po114 , po115 , po116 , po117 ,
    po118 , po119 , po120 , po121 , po122 , po123 , po124 ,
    po125 , po126 , po127   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 , pi104 ,
    pi105 , pi106 , pi107 , pi108 , pi109 , pi110 , pi111 , pi112 ,
    pi113 , pi114 , pi115 , pi116 , pi117 , pi118 , pi119 , pi120 ,
    pi121 , pi122 , pi123 , pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 , po7 ,
    po8 , po9 , po10 , po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 , po21 , po22 , po23 ,
    po24 , po25 , po26 , po27 , po28 , po29 , po30 , po31 ,
    po32 , po33 , po34 , po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 , po45 , po46 , po47 ,
    po48 , po49 , po50 , po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 , po61 , po62 , po63 ,
    po64 , po65 , po66 , po67 , po68 , po69 , po70 , po71 ,
    po72 , po73 , po74 , po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 , po85 , po86 , po87 ,
    po88 , po89 , po90 , po91 , po92 , po93 , po94 , po95 ,
    po96 , po97 , po98 , po99 , po100 , po101 , po102 ,
    po103 , po104 , po105 , po106 , po107 , po108 , po109 ,
    po110 , po111 , po112 , po113 , po114 , po115 , po116 ,
    po117 , po118 , po119 , po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ;
  wire n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278,
    n280, n281, n282, n283, n284, n285, n286,
    n287, n288, n289, n290, n291, n292, n293,
    n294, n295, n296, n297, n298, n299, n301,
    n302, n303, n304, n305, n306, n307, n308,
    n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322,
    n323, n324, n325, n326, n327, n328, n330,
    n331, n332, n333, n334, n335, n336, n337,
    n338, n339, n340, n341, n342, n343, n344,
    n345, n346, n347, n348, n349, n350, n351,
    n352, n353, n354, n355, n356, n357, n358,
    n359, n360, n361, n362, n363, n364, n365,
    n366, n367, n368, n369, n370, n371, n372,
    n373, n374, n375, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415,
    n416, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686,
    n687, n688, n689, n690, n691, n692, n693,
    n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707,
    n708, n709, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n735, n736,
    n737, n738, n739, n740, n741, n742, n743,
    n744, n745, n746, n747, n748, n749, n750,
    n751, n752, n753, n754, n755, n756, n757,
    n758, n759, n760, n761, n762, n763, n764,
    n765, n766, n767, n768, n769, n770, n771,
    n772, n773, n774, n775, n776, n777, n778,
    n779, n780, n781, n782, n783, n784, n785,
    n786, n787, n788, n789, n790, n791, n792,
    n793, n794, n795, n796, n797, n798, n799,
    n800, n801, n802, n803, n804, n805, n806,
    n807, n808, n809, n810, n812, n813, n814,
    n815, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n834, n835,
    n836, n837, n838, n839, n840, n841, n842,
    n843, n844, n845, n846, n847, n848, n849,
    n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863,
    n864, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877,
    n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n889, n890, n891,
    n892, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n994, n995, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1312, n1313,
    n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325,
    n1326, n1327, n1328, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1336, n1337,
    n1338, n1339, n1340, n1341, n1342, n1343,
    n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355,
    n1356, n1357, n1358, n1359, n1360, n1361,
    n1362, n1363, n1364, n1365, n1366, n1367,
    n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385,
    n1386, n1387, n1388, n1389, n1390, n1391,
    n1392, n1393, n1394, n1395, n1396, n1397,
    n1398, n1399, n1400, n1401, n1402, n1403,
    n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415,
    n1416, n1417, n1418, n1419, n1420, n1421,
    n1422, n1423, n1424, n1425, n1426, n1427,
    n1429, n1430, n1431, n1432, n1433, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446,
    n1447, n1448, n1449, n1450, n1451, n1452,
    n1453, n1454, n1455, n1456, n1457, n1458,
    n1459, n1460, n1461, n1462, n1463, n1464,
    n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476,
    n1477, n1478, n1479, n1480, n1481, n1482,
    n1483, n1484, n1485, n1486, n1487, n1488,
    n1489, n1490, n1491, n1492, n1493, n1494,
    n1495, n1496, n1497, n1498, n1499, n1500,
    n1501, n1502, n1503, n1504, n1505, n1506,
    n1507, n1508, n1509, n1510, n1511, n1512,
    n1513, n1514, n1515, n1516, n1517, n1518,
    n1519, n1520, n1521, n1522, n1523, n1524,
    n1525, n1526, n1527, n1528, n1529, n1530,
    n1531, n1532, n1533, n1534, n1535, n1536,
    n1537, n1538, n1539, n1540, n1541, n1542,
    n1543, n1544, n1545, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561,
    n1562, n1563, n1564, n1565, n1566, n1567,
    n1568, n1569, n1570, n1571, n1572, n1573,
    n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591,
    n1592, n1593, n1594, n1595, n1596, n1597,
    n1598, n1599, n1600, n1601, n1602, n1603,
    n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615,
    n1616, n1617, n1618, n1619, n1620, n1621,
    n1622, n1623, n1624, n1625, n1626, n1627,
    n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645,
    n1646, n1647, n1648, n1649, n1650, n1651,
    n1652, n1653, n1654, n1655, n1656, n1657,
    n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675,
    n1676, n1677, n1678, n1679, n1680, n1681,
    n1682, n1683, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1956, n1957, n1958, n1959, n1960,
    n1961, n1962, n1963, n1964, n1965, n1966,
    n1967, n1968, n1969, n1970, n1971, n1972,
    n1973, n1974, n1975, n1976, n1977, n1978,
    n1979, n1980, n1981, n1982, n1983, n1984,
    n1985, n1986, n1987, n1988, n1989, n1990,
    n1991, n1992, n1993, n1994, n1995, n1996,
    n1997, n1998, n1999, n2000, n2001, n2002,
    n2003, n2004, n2005, n2006, n2007, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026,
    n2027, n2028, n2029, n2030, n2031, n2032,
    n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056,
    n2057, n2058, n2059, n2060, n2061, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2080,
    n2081, n2082, n2083, n2084, n2085, n2086,
    n2087, n2088, n2089, n2090, n2091, n2092,
    n2093, n2094, n2095, n2096, n2097, n2098,
    n2099, n2100, n2101, n2102, n2103, n2104,
    n2105, n2106, n2107, n2108, n2109, n2110,
    n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2153,
    n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165,
    n2166, n2167, n2168, n2169, n2170, n2171,
    n2172, n2173, n2174, n2175, n2176, n2177,
    n2178, n2179, n2180, n2181, n2182, n2183,
    n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195,
    n2196, n2197, n2198, n2199, n2200, n2201,
    n2202, n2203, n2204, n2205, n2206, n2207,
    n2208, n2209, n2210, n2211, n2212, n2213,
    n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225,
    n2226, n2227, n2228, n2229, n2230, n2231,
    n2232, n2233, n2234, n2235, n2236, n2237,
    n2238, n2239, n2240, n2241, n2242, n2243,
    n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255,
    n2256, n2257, n2258, n2259, n2260, n2261,
    n2262, n2263, n2265, n2266, n2267, n2268,
    n2269, n2270, n2271, n2272, n2273, n2274,
    n2275, n2276, n2277, n2278, n2279, n2280,
    n2281, n2282, n2283, n2284, n2285, n2286,
    n2287, n2288, n2289, n2290, n2291, n2292,
    n2293, n2294, n2295, n2296, n2297, n2298,
    n2299, n2300, n2301, n2302, n2303, n2304,
    n2305, n2306, n2307, n2308, n2309, n2310,
    n2311, n2312, n2313, n2314, n2315, n2316,
    n2317, n2318, n2319, n2320, n2321, n2322,
    n2323, n2324, n2325, n2326, n2327, n2328,
    n2329, n2330, n2331, n2332, n2333, n2334,
    n2335, n2336, n2337, n2338, n2339, n2340,
    n2341, n2342, n2343, n2344, n2345, n2346,
    n2347, n2348, n2349, n2350, n2351, n2352,
    n2353, n2354, n2355, n2356, n2357, n2358,
    n2359, n2360, n2361, n2362, n2363, n2364,
    n2365, n2366, n2367, n2368, n2369, n2370,
    n2371, n2372, n2373, n2374, n2375, n2376,
    n2377, n2378, n2379, n2380, n2381, n2382,
    n2383, n2384, n2385, n2386, n2387, n2388,
    n2389, n2390, n2391, n2392, n2393, n2394,
    n2395, n2396, n2397, n2398, n2399, n2400,
    n2401, n2402, n2403, n2404, n2405, n2406,
    n2407, n2408, n2409, n2410, n2411, n2412,
    n2413, n2414, n2415, n2416, n2417, n2418,
    n2420, n2421, n2422, n2423, n2424, n2425,
    n2426, n2427, n2428, n2429, n2430, n2431,
    n2432, n2433, n2434, n2435, n2436, n2437,
    n2438, n2439, n2440, n2441, n2442, n2443,
    n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455,
    n2456, n2457, n2458, n2459, n2460, n2461,
    n2462, n2463, n2464, n2465, n2466, n2467,
    n2468, n2469, n2470, n2471, n2472, n2473,
    n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485,
    n2486, n2487, n2488, n2489, n2490, n2491,
    n2492, n2493, n2494, n2495, n2496, n2497,
    n2498, n2499, n2500, n2501, n2502, n2503,
    n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515,
    n2516, n2517, n2518, n2519, n2520, n2521,
    n2522, n2523, n2524, n2525, n2526, n2527,
    n2528, n2529, n2530, n2531, n2532, n2533,
    n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545,
    n2546, n2547, n2548, n2549, n2550, n2551,
    n2552, n2553, n2554, n2555, n2556, n2557,
    n2558, n2559, n2560, n2561, n2562, n2563,
    n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575,
    n2576, n2577, n2578, n2579, n2580, n2581,
    n2582, n2583, n2584, n2585, n2586, n2587,
    n2588, n2589, n2590, n2591, n2592, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2939, n2940, n2941, n2942, n2943, n2944,
    n2945, n2946, n2947, n2948, n2949, n2950,
    n2951, n2952, n2953, n2954, n2955, n2956,
    n2957, n2958, n2959, n2960, n2961, n2962,
    n2963, n2964, n2965, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2982, n2983, n2984, n2985, n2986,
    n2987, n2988, n2989, n2990, n2991, n2992,
    n2993, n2994, n2995, n2996, n2997, n2998,
    n2999, n3000, n3001, n3002, n3003, n3004,
    n3005, n3006, n3007, n3008, n3009, n3010,
    n3011, n3012, n3013, n3014, n3015, n3016,
    n3017, n3018, n3019, n3020, n3021, n3022,
    n3023, n3024, n3025, n3026, n3027, n3028,
    n3029, n3030, n3031, n3032, n3033, n3034,
    n3035, n3036, n3037, n3038, n3039, n3040,
    n3041, n3042, n3043, n3044, n3045, n3046,
    n3047, n3048, n3049, n3050, n3051, n3052,
    n3053, n3054, n3055, n3056, n3057, n3058,
    n3059, n3060, n3061, n3062, n3063, n3064,
    n3065, n3066, n3067, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3079, n3080, n3081, n3082,
    n3083, n3084, n3085, n3086, n3087, n3088,
    n3089, n3090, n3091, n3092, n3093, n3094,
    n3095, n3096, n3097, n3098, n3099, n3100,
    n3101, n3102, n3103, n3104, n3105, n3106,
    n3107, n3108, n3109, n3110, n3111, n3112,
    n3113, n3114, n3115, n3116, n3117, n3118,
    n3119, n3120, n3121, n3122, n3123, n3124,
    n3125, n3126, n3127, n3128, n3129, n3130,
    n3132, n3133, n3134, n3135, n3136, n3137,
    n3138, n3139, n3140, n3141, n3142, n3143,
    n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3151, n3152, n3153, n3154, n3155,
    n3156, n3157, n3158, n3159, n3160, n3161,
    n3162, n3163, n3164, n3165, n3166, n3167,
    n3168, n3169, n3170, n3171, n3172, n3173,
    n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3184, n3185,
    n3186, n3187, n3188, n3189, n3190, n3191,
    n3192, n3193, n3194, n3195, n3196, n3197,
    n3198, n3199, n3200, n3201, n3202, n3203,
    n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215,
    n3216, n3217, n3218, n3219, n3220, n3221,
    n3222, n3223, n3224, n3225, n3226, n3227,
    n3228, n3229, n3230, n3231, n3232, n3233,
    n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245,
    n3246, n3247, n3248, n3249, n3250, n3251,
    n3252, n3253, n3254, n3255, n3256, n3257,
    n3258, n3259, n3260, n3261, n3262, n3263,
    n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275,
    n3276, n3277, n3278, n3279, n3280, n3281,
    n3282, n3283, n3284, n3285, n3286, n3287,
    n3288, n3289, n3290, n3291, n3292, n3293,
    n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305,
    n3306, n3307, n3308, n3309, n3310, n3311,
    n3312, n3313, n3314, n3315, n3316, n3317,
    n3318, n3319, n3320, n3322, n3323, n3324,
    n3325, n3326, n3327, n3328, n3329, n3330,
    n3331, n3332, n3333, n3334, n3335, n3336,
    n3337, n3338, n3339, n3340, n3341, n3342,
    n3343, n3344, n3345, n3346, n3347, n3348,
    n3349, n3350, n3351, n3352, n3353, n3354,
    n3355, n3356, n3357, n3358, n3359, n3360,
    n3361, n3362, n3363, n3364, n3365, n3366,
    n3367, n3368, n3369, n3370, n3371, n3372,
    n3373, n3374, n3375, n3376, n3377, n3378,
    n3379, n3380, n3381, n3382, n3383, n3384,
    n3385, n3386, n3387, n3388, n3389, n3390,
    n3391, n3392, n3393, n3394, n3395, n3396,
    n3397, n3398, n3399, n3400, n3401, n3402,
    n3403, n3404, n3405, n3406, n3407, n3408,
    n3409, n3410, n3411, n3412, n3413, n3414,
    n3415, n3416, n3417, n3418, n3419, n3420,
    n3421, n3422, n3423, n3424, n3425, n3426,
    n3427, n3428, n3429, n3430, n3431, n3432,
    n3433, n3434, n3435, n3436, n3437, n3438,
    n3439, n3440, n3441, n3442, n3443, n3444,
    n3445, n3446, n3447, n3448, n3449, n3450,
    n3451, n3452, n3453, n3454, n3455, n3456,
    n3457, n3458, n3459, n3460, n3461, n3462,
    n3463, n3464, n3465, n3466, n3467, n3468,
    n3469, n3470, n3471, n3472, n3473, n3474,
    n3475, n3476, n3477, n3478, n3479, n3480,
    n3481, n3482, n3483, n3484, n3485, n3486,
    n3487, n3488, n3489, n3490, n3491, n3492,
    n3493, n3494, n3495, n3496, n3497, n3498,
    n3499, n3500, n3501, n3502, n3503, n3504,
    n3505, n3506, n3507, n3508, n3509, n3510,
    n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3523,
    n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535,
    n3536, n3537, n3538, n3539, n3540, n3541,
    n3542, n3543, n3544, n3545, n3546, n3547,
    n3548, n3549, n3550, n3551, n3552, n3553,
    n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565,
    n3566, n3567, n3568, n3569, n3570, n3571,
    n3572, n3573, n3574, n3575, n3576, n3577,
    n3578, n3579, n3580, n3581, n3582, n3583,
    n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595,
    n3596, n3597, n3598, n3599, n3600, n3601,
    n3602, n3603, n3604, n3605, n3606, n3607,
    n3608, n3609, n3610, n3611, n3612, n3613,
    n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625,
    n3626, n3627, n3628, n3629, n3630, n3631,
    n3632, n3633, n3634, n3635, n3636, n3637,
    n3638, n3639, n3640, n3641, n3642, n3643,
    n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655,
    n3656, n3657, n3658, n3659, n3660, n3661,
    n3662, n3663, n3664, n3665, n3666, n3667,
    n3668, n3669, n3670, n3671, n3672, n3673,
    n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685,
    n3686, n3687, n3688, n3689, n3690, n3691,
    n3692, n3693, n3694, n3695, n3696, n3697,
    n3698, n3699, n3700, n3701, n3702, n3703,
    n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715,
    n3716, n3717, n3718, n3719, n3720, n3721,
    n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782,
    n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932,
    n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951,
    n3952, n3953, n3954, n3955, n3956, n3957,
    n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987,
    n3988, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4017,
    n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047,
    n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077,
    n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101,
    n4102, n4103, n4104, n4105, n4106, n4107,
    n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131,
    n4132, n4133, n4134, n4135, n4136, n4137,
    n4138, n4140, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156,
    n4157, n4158, n4159, n4160, n4161, n4162,
    n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174,
    n4175, n4176, n4177, n4178, n4179, n4180,
    n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192,
    n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204,
    n4205, n4206, n4207, n4208, n4209, n4210,
    n4211, n4212, n4213, n4214, n4215, n4216,
    n4217, n4218, n4219, n4220, n4221, n4222,
    n4223, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234,
    n4235, n4236, n4237, n4238, n4239, n4240,
    n4241, n4242, n4243, n4244, n4245, n4246,
    n4247, n4248, n4249, n4250, n4251, n4252,
    n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4267, n4268, n4269, n4270,
    n4271, n4272, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4280, n4281, n4282,
    n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294,
    n4295, n4296, n4297, n4298, n4299, n4300,
    n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4322, n4323, n4324,
    n4325, n4326, n4327, n4328, n4329, n4330,
    n4331, n4332, n4333, n4334, n4335, n4336,
    n4337, n4338, n4339, n4340, n4341, n4342,
    n4343, n4344, n4345, n4346, n4347, n4348,
    n4349, n4350, n4351, n4352, n4353, n4354,
    n4355, n4356, n4357, n4358, n4359, n4360,
    n4361, n4362, n4363, n4364, n4365, n4366,
    n4367, n4368, n4369, n4370, n4371, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385,
    n4386, n4387, n4388, n4389, n4390, n4391,
    n4392, n4393, n4394, n4395, n4396, n4397,
    n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4421,
    n4422, n4423, n4424, n4425, n4426, n4427,
    n4428, n4429, n4430, n4431, n4432, n4433,
    n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451,
    n4452, n4453, n4454, n4455, n4456, n4457,
    n4458, n4459, n4460, n4461, n4462, n4463,
    n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481,
    n4482, n4483, n4484, n4485, n4486, n4487,
    n4488, n4489, n4490, n4491, n4492, n4493,
    n4494, n4495, n4496, n4497, n4498, n4499,
    n4500, n4501, n4502, n4503, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511,
    n4512, n4513, n4514, n4515, n4516, n4517,
    n4518, n4519, n4520, n4521, n4522, n4523,
    n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535,
    n4536, n4537, n4538, n4539, n4540, n4541,
    n4542, n4543, n4544, n4545, n4546, n4547,
    n4548, n4549, n4550, n4551, n4552, n4553,
    n4554, n4555, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571,
    n4572, n4573, n4574, n4575, n4576, n4577,
    n4578, n4579, n4580, n4581, n4582, n4583,
    n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595,
    n4597, n4598, n4599, n4600, n4601, n4602,
    n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662,
    n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686,
    n4687, n4688, n4689, n4690, n4691, n4692,
    n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710,
    n4711, n4712, n4713, n4714, n4715, n4716,
    n4717, n4718, n4719, n4720, n4721, n4722,
    n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734,
    n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752,
    n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764,
    n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776,
    n4777, n4778, n4779, n4780, n4781, n4782,
    n4783, n4784, n4785, n4786, n4787, n4788,
    n4789, n4790, n4791, n4792, n4793, n4794,
    n4795, n4796, n4797, n4798, n4799, n4800,
    n4801, n4802, n4803, n4804, n4805, n4806,
    n4807, n4808, n4809, n4810, n4811, n4812,
    n4813, n4814, n4815, n4816, n4817, n4818,
    n4819, n4821, n4822, n4823, n4824, n4825,
    n4826, n4827, n4828, n4829, n4830, n4831,
    n4832, n4833, n4834, n4835, n4836, n4837,
    n4838, n4839, n4840, n4841, n4842, n4843,
    n4844, n4845, n4846, n4847, n4848, n4849,
    n4850, n4851, n4852, n4853, n4854, n4855,
    n4856, n4857, n4858, n4859, n4860, n4861,
    n4862, n4863, n4864, n4865, n4866, n4867,
    n4868, n4869, n4870, n4871, n4872, n4873,
    n4874, n4875, n4876, n4877, n4878, n4879,
    n4880, n4881, n4882, n4883, n4884, n4885,
    n4886, n4887, n4888, n4889, n4890, n4891,
    n4892, n4893, n4894, n4895, n4896, n4897,
    n4898, n4899, n4900, n4901, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5069, n5070, n5071, n5072,
    n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5309, n5310, n5311, n5312, n5313,
    n5314, n5315, n5316, n5317, n5318, n5319,
    n5320, n5321, n5322, n5323, n5324, n5325,
    n5326, n5327, n5328, n5329, n5330, n5331,
    n5332, n5333, n5334, n5335, n5336, n5337,
    n5338, n5339, n5340, n5341, n5342, n5343,
    n5344, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5352, n5353, n5354, n5355,
    n5356, n5357, n5358, n5359, n5360, n5361,
    n5362, n5363, n5364, n5365, n5366, n5367,
    n5368, n5369, n5370, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391,
    n5392, n5393, n5394, n5395, n5396, n5397,
    n5398, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409,
    n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421,
    n5422, n5423, n5424, n5425, n5426, n5427,
    n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451,
    n5452, n5453, n5454, n5455, n5456, n5457,
    n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481,
    n5482, n5483, n5484, n5485, n5486, n5487,
    n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499,
    n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511,
    n5512, n5513, n5514, n5515, n5516, n5517,
    n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541,
    n5542, n5543, n5544, n5545, n5546, n5547,
    n5548, n5549, n5550, n5551, n5553, n5554,
    n5555, n5556, n5557, n5558, n5559, n5560,
    n5561, n5562, n5563, n5564, n5565, n5566,
    n5567, n5568, n5569, n5570, n5571, n5572,
    n5573, n5574, n5575, n5576, n5577, n5578,
    n5579, n5580, n5581, n5582, n5583, n5584,
    n5585, n5586, n5587, n5588, n5589, n5590,
    n5591, n5592, n5593, n5594, n5595, n5596,
    n5597, n5598, n5599, n5600, n5601, n5602,
    n5603, n5604, n5605, n5606, n5607, n5608,
    n5609, n5610, n5611, n5612, n5613, n5614,
    n5615, n5616, n5617, n5618, n5619, n5620,
    n5621, n5622, n5623, n5624, n5625, n5626,
    n5627, n5628, n5629, n5630, n5631, n5632,
    n5633, n5634, n5635, n5636, n5637, n5638,
    n5639, n5640, n5641, n5642, n5643, n5644,
    n5645, n5646, n5647, n5648, n5649, n5650,
    n5651, n5652, n5653, n5654, n5655, n5656,
    n5657, n5658, n5659, n5660, n5661, n5662,
    n5663, n5664, n5665, n5666, n5667, n5668,
    n5669, n5670, n5671, n5672, n5673, n5674,
    n5675, n5676, n5677, n5678, n5679, n5680,
    n5681, n5682, n5683, n5684, n5685, n5686,
    n5687, n5688, n5689, n5690, n5691, n5692,
    n5693, n5694, n5695, n5696, n5697, n5698,
    n5699, n5700, n5701, n5702, n5703, n5704,
    n5705, n5706, n5707, n5708, n5709, n5710,
    n5711, n5712, n5713, n5714, n5715, n5716,
    n5717, n5718, n5719, n5720, n5721, n5722,
    n5723, n5724, n5725, n5726, n5727, n5728,
    n5729, n5730, n5731, n5732, n5733, n5734,
    n5735, n5736, n5737, n5738, n5739, n5740,
    n5741, n5742, n5743, n5744, n5745, n5746,
    n5747, n5748, n5749, n5750, n5751, n5752,
    n5753, n5754, n5755, n5756, n5757, n5758,
    n5759, n5760, n5761, n5762, n5763, n5764,
    n5765, n5766, n5767, n5768, n5769, n5770,
    n5771, n5772, n5773, n5774, n5775, n5776,
    n5777, n5778, n5779, n5780, n5781, n5782,
    n5783, n5784, n5785, n5786, n5787, n5788,
    n5789, n5790, n5791, n5792, n5793, n5794,
    n5795, n5796, n5797, n5798, n5799, n5800,
    n5801, n5802, n5803, n5804, n5805, n5806,
    n5807, n5808, n5809, n5810, n5811, n5812,
    n5813, n5814, n5815, n5816, n5817, n5819,
    n5820, n5821, n5822, n5823, n5824, n5825,
    n5826, n5827, n5828, n5829, n5830, n5831,
    n5832, n5833, n5834, n5835, n5836, n5837,
    n5838, n5839, n5840, n5841, n5842, n5843,
    n5844, n5845, n5846, n5847, n5848, n5849,
    n5850, n5851, n5852, n5853, n5854, n5855,
    n5856, n5857, n5858, n5859, n5860, n5861,
    n5862, n5863, n5864, n5865, n5866, n5867,
    n5868, n5869, n5870, n5871, n5872, n5873,
    n5874, n5875, n5876, n5877, n5878, n5879,
    n5880, n5881, n5882, n5883, n5884, n5885,
    n5886, n5887, n5888, n5889, n5890, n5891,
    n5892, n5893, n5894, n5895, n5896, n5897,
    n5898, n5899, n5900, n5901, n5902, n5903,
    n5904, n5905, n5906, n5907, n5908, n5909,
    n5910, n5911, n5912, n5913, n5914, n5915,
    n5916, n5917, n5918, n5919, n5920, n5921,
    n5922, n5923, n5924, n5925, n5926, n5927,
    n5928, n5929, n5930, n5931, n5932, n5933,
    n5934, n5935, n5936, n5937, n5938, n5939,
    n5940, n5941, n5942, n5943, n5944, n5945,
    n5946, n5947, n5948, n5949, n5950, n5951,
    n5952, n5953, n5954, n5955, n5956, n5957,
    n5958, n5959, n5960, n5961, n5962, n5963,
    n5964, n5965, n5966, n5967, n5968, n5969,
    n5970, n5971, n5972, n5973, n5974, n5975,
    n5976, n5977, n5978, n5979, n5980, n5981,
    n5982, n5983, n5984, n5985, n5986, n5987,
    n5988, n5989, n5990, n5991, n5992, n5993,
    n5994, n5995, n5996, n5997, n5998, n5999,
    n6000, n6001, n6002, n6003, n6004, n6005,
    n6006, n6007, n6008, n6009, n6010, n6011,
    n6012, n6013, n6014, n6015, n6016, n6017,
    n6018, n6019, n6020, n6021, n6022, n6023,
    n6024, n6025, n6026, n6027, n6028, n6029,
    n6030, n6031, n6032, n6033, n6034, n6035,
    n6036, n6037, n6038, n6039, n6040, n6041,
    n6042, n6043, n6044, n6045, n6046, n6047,
    n6048, n6049, n6050, n6051, n6052, n6053,
    n6054, n6055, n6056, n6057, n6058, n6059,
    n6060, n6061, n6062, n6063, n6064, n6065,
    n6066, n6067, n6068, n6069, n6070, n6071,
    n6072, n6073, n6074, n6075, n6076, n6078,
    n6079, n6080, n6081, n6082, n6083, n6084,
    n6085, n6086, n6087, n6088, n6089, n6090,
    n6091, n6092, n6093, n6094, n6095, n6096,
    n6097, n6098, n6099, n6100, n6101, n6102,
    n6103, n6104, n6105, n6106, n6107, n6108,
    n6109, n6110, n6111, n6112, n6113, n6114,
    n6115, n6116, n6117, n6118, n6119, n6120,
    n6121, n6122, n6123, n6124, n6125, n6126,
    n6127, n6128, n6129, n6130, n6131, n6132,
    n6133, n6134, n6135, n6136, n6137, n6138,
    n6139, n6140, n6141, n6142, n6143, n6144,
    n6145, n6146, n6147, n6148, n6149, n6150,
    n6151, n6152, n6153, n6154, n6155, n6156,
    n6157, n6158, n6159, n6160, n6161, n6162,
    n6163, n6164, n6165, n6166, n6167, n6168,
    n6169, n6170, n6171, n6172, n6173, n6174,
    n6175, n6176, n6177, n6178, n6179, n6180,
    n6181, n6182, n6183, n6184, n6185, n6186,
    n6187, n6188, n6189, n6190, n6191, n6192,
    n6193, n6194, n6195, n6196, n6197, n6198,
    n6199, n6200, n6201, n6202, n6203, n6204,
    n6205, n6206, n6207, n6208, n6209, n6210,
    n6211, n6212, n6213, n6214, n6215, n6216,
    n6217, n6218, n6219, n6220, n6221, n6222,
    n6223, n6224, n6225, n6226, n6227, n6228,
    n6229, n6230, n6231, n6232, n6233, n6234,
    n6235, n6236, n6237, n6238, n6239, n6240,
    n6241, n6242, n6243, n6244, n6245, n6246,
    n6247, n6248, n6249, n6250, n6251, n6252,
    n6253, n6254, n6255, n6256, n6257, n6258,
    n6259, n6260, n6261, n6262, n6263, n6264,
    n6265, n6266, n6267, n6268, n6269, n6270,
    n6271, n6272, n6273, n6274, n6275, n6276,
    n6277, n6278, n6279, n6280, n6281, n6282,
    n6283, n6284, n6285, n6286, n6287, n6288,
    n6289, n6290, n6291, n6292, n6293, n6294,
    n6295, n6296, n6297, n6298, n6299, n6300,
    n6301, n6302, n6303, n6304, n6305, n6306,
    n6307, n6308, n6309, n6310, n6311, n6312,
    n6313, n6314, n6315, n6316, n6317, n6318,
    n6319, n6320, n6321, n6322, n6323, n6324,
    n6325, n6326, n6327, n6328, n6329, n6330,
    n6331, n6332, n6333, n6334, n6335, n6336,
    n6337, n6338, n6339, n6341, n6342, n6343,
    n6344, n6345, n6346, n6347, n6348, n6349,
    n6350, n6351, n6352, n6353, n6354, n6355,
    n6356, n6357, n6358, n6359, n6360, n6361,
    n6362, n6363, n6364, n6365, n6366, n6367,
    n6368, n6369, n6370, n6371, n6372, n6373,
    n6374, n6375, n6376, n6377, n6378, n6379,
    n6380, n6381, n6382, n6383, n6384, n6385,
    n6386, n6387, n6388, n6389, n6390, n6391,
    n6392, n6393, n6394, n6395, n6396, n6397,
    n6398, n6399, n6400, n6401, n6402, n6403,
    n6404, n6405, n6406, n6407, n6408, n6409,
    n6410, n6411, n6412, n6413, n6414, n6415,
    n6416, n6417, n6418, n6419, n6420, n6421,
    n6422, n6423, n6424, n6425, n6426, n6427,
    n6428, n6429, n6430, n6431, n6432, n6433,
    n6434, n6435, n6436, n6437, n6438, n6439,
    n6440, n6441, n6442, n6443, n6444, n6445,
    n6446, n6447, n6448, n6449, n6450, n6451,
    n6452, n6453, n6454, n6455, n6456, n6457,
    n6458, n6459, n6460, n6461, n6462, n6463,
    n6464, n6465, n6466, n6467, n6468, n6469,
    n6470, n6471, n6472, n6473, n6474, n6475,
    n6476, n6477, n6478, n6479, n6480, n6481,
    n6482, n6483, n6484, n6485, n6486, n6487,
    n6488, n6489, n6490, n6491, n6492, n6493,
    n6494, n6495, n6496, n6497, n6498, n6499,
    n6500, n6501, n6502, n6503, n6504, n6505,
    n6506, n6507, n6508, n6509, n6510, n6511,
    n6512, n6513, n6514, n6515, n6516, n6517,
    n6518, n6519, n6520, n6521, n6522, n6523,
    n6524, n6525, n6526, n6527, n6528, n6529,
    n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541,
    n6542, n6543, n6544, n6545, n6546, n6547,
    n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571,
    n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601,
    n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625,
    n6627, n6628, n6629, n6630, n6631, n6632,
    n6633, n6634, n6635, n6636, n6637, n6638,
    n6639, n6640, n6641, n6642, n6643, n6644,
    n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6903,
    n6904, n6905, n6906, n6907, n6908, n6909,
    n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921,
    n6922, n6923, n6924, n6925, n6926, n6927,
    n6928, n6929, n6930, n6931, n6932, n6933,
    n6934, n6935, n6936, n6937, n6938, n6939,
    n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951,
    n6952, n6953, n6954, n6955, n6956, n6957,
    n6958, n6959, n6960, n6961, n6962, n6963,
    n6964, n6965, n6966, n6967, n6968, n6969,
    n6970, n6971, n6972, n6973, n6974, n6975,
    n6976, n6977, n6978, n6979, n6980, n6981,
    n6982, n6983, n6984, n6985, n6986, n6987,
    n6988, n6989, n6990, n6991, n6992, n6993,
    n6994, n6995, n6996, n6997, n6998, n6999,
    n7000, n7001, n7002, n7003, n7004, n7005,
    n7006, n7007, n7008, n7009, n7010, n7011,
    n7012, n7013, n7014, n7015, n7016, n7017,
    n7018, n7019, n7020, n7021, n7022, n7023,
    n7024, n7025, n7026, n7027, n7028, n7029,
    n7030, n7031, n7032, n7033, n7034, n7035,
    n7036, n7037, n7038, n7039, n7040, n7041,
    n7042, n7043, n7044, n7045, n7046, n7047,
    n7048, n7049, n7050, n7051, n7052, n7053,
    n7054, n7055, n7056, n7057, n7058, n7059,
    n7060, n7061, n7062, n7063, n7064, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071,
    n7072, n7073, n7074, n7075, n7076, n7077,
    n7078, n7079, n7080, n7081, n7082, n7083,
    n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101,
    n7102, n7103, n7104, n7105, n7106, n7107,
    n7108, n7109, n7110, n7111, n7112, n7113,
    n7114, n7115, n7116, n7117, n7118, n7119,
    n7120, n7121, n7122, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131,
    n7132, n7133, n7134, n7135, n7136, n7137,
    n7138, n7139, n7140, n7141, n7142, n7143,
    n7144, n7145, n7146, n7147, n7148, n7149,
    n7150, n7151, n7152, n7153, n7154, n7155,
    n7156, n7157, n7158, n7159, n7160, n7161,
    n7162, n7163, n7164, n7165, n7166, n7167,
    n7168, n7169, n7170, n7171, n7172, n7173,
    n7174, n7175, n7176, n7177, n7178, n7179,
    n7180, n7181, n7183, n7184, n7185, n7186,
    n7187, n7188, n7189, n7190, n7191, n7192,
    n7193, n7194, n7195, n7196, n7197, n7198,
    n7199, n7200, n7201, n7202, n7203, n7204,
    n7205, n7206, n7207, n7208, n7209, n7210,
    n7211, n7212, n7213, n7214, n7215, n7216,
    n7217, n7218, n7219, n7220, n7221, n7222,
    n7223, n7224, n7225, n7226, n7227, n7228,
    n7229, n7230, n7231, n7232, n7233, n7234,
    n7235, n7236, n7237, n7238, n7239, n7240,
    n7241, n7242, n7243, n7244, n7245, n7246,
    n7247, n7248, n7249, n7250, n7251, n7252,
    n7253, n7254, n7255, n7256, n7257, n7258,
    n7259, n7260, n7261, n7262, n7263, n7264,
    n7265, n7266, n7267, n7268, n7269, n7270,
    n7271, n7272, n7273, n7274, n7275, n7276,
    n7277, n7278, n7279, n7280, n7281, n7282,
    n7283, n7284, n7285, n7286, n7287, n7288,
    n7289, n7290, n7291, n7292, n7293, n7294,
    n7295, n7296, n7297, n7298, n7299, n7300,
    n7301, n7302, n7303, n7304, n7305, n7306,
    n7307, n7308, n7309, n7310, n7311, n7312,
    n7313, n7314, n7315, n7316, n7317, n7318,
    n7319, n7320, n7321, n7322, n7323, n7324,
    n7325, n7326, n7327, n7328, n7329, n7330,
    n7331, n7332, n7333, n7334, n7335, n7336,
    n7337, n7338, n7339, n7340, n7341, n7342,
    n7343, n7344, n7345, n7346, n7347, n7348,
    n7349, n7350, n7351, n7352, n7353, n7354,
    n7355, n7356, n7357, n7358, n7359, n7360,
    n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7370, n7371, n7372,
    n7373, n7374, n7375, n7376, n7377, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390,
    n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7398, n7399, n7400, n7401, n7402,
    n7403, n7404, n7405, n7406, n7407, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414,
    n7415, n7416, n7417, n7418, n7419, n7420,
    n7421, n7422, n7423, n7424, n7425, n7426,
    n7427, n7428, n7429, n7430, n7431, n7432,
    n7433, n7434, n7435, n7436, n7437, n7438,
    n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7448, n7449, n7450,
    n7451, n7452, n7453, n7454, n7455, n7456,
    n7457, n7458, n7459, n7460, n7461, n7462,
    n7463, n7464, n7465, n7466, n7467, n7468,
    n7469, n7470, n7471, n7472, n7473, n7474,
    n7475, n7476, n7477, n7478, n7479, n7480,
    n7481, n7482, n7483, n7484, n7485, n7487,
    n7488, n7489, n7490, n7491, n7492, n7493,
    n7494, n7495, n7496, n7497, n7498, n7499,
    n7500, n7501, n7502, n7503, n7504, n7505,
    n7506, n7507, n7508, n7509, n7510, n7511,
    n7512, n7513, n7514, n7515, n7516, n7517,
    n7518, n7519, n7520, n7521, n7522, n7523,
    n7524, n7525, n7526, n7527, n7528, n7529,
    n7530, n7531, n7532, n7533, n7534, n7535,
    n7536, n7537, n7538, n7539, n7540, n7541,
    n7542, n7543, n7544, n7545, n7546, n7547,
    n7548, n7549, n7550, n7551, n7552, n7553,
    n7554, n7555, n7556, n7557, n7558, n7559,
    n7560, n7561, n7562, n7563, n7564, n7565,
    n7566, n7567, n7568, n7569, n7570, n7571,
    n7572, n7573, n7574, n7575, n7576, n7577,
    n7578, n7579, n7580, n7581, n7582, n7583,
    n7584, n7585, n7586, n7587, n7588, n7589,
    n7590, n7591, n7592, n7593, n7594, n7595,
    n7596, n7597, n7598, n7599, n7600, n7601,
    n7602, n7603, n7604, n7605, n7606, n7607,
    n7608, n7609, n7610, n7611, n7612, n7613,
    n7614, n7615, n7616, n7617, n7618, n7619,
    n7620, n7621, n7622, n7623, n7624, n7625,
    n7626, n7627, n7628, n7629, n7630, n7631,
    n7632, n7633, n7634, n7635, n7636, n7637,
    n7638, n7639, n7640, n7641, n7642, n7643,
    n7644, n7645, n7646, n7647, n7648, n7649,
    n7650, n7651, n7652, n7653, n7654, n7655,
    n7656, n7657, n7658, n7659, n7660, n7661,
    n7662, n7663, n7664, n7665, n7666, n7667,
    n7668, n7669, n7670, n7671, n7672, n7673,
    n7674, n7675, n7676, n7677, n7678, n7679,
    n7680, n7681, n7682, n7683, n7684, n7685,
    n7686, n7687, n7688, n7689, n7690, n7691,
    n7692, n7693, n7694, n7695, n7696, n7697,
    n7698, n7699, n7700, n7701, n7702, n7703,
    n7704, n7705, n7706, n7707, n7708, n7709,
    n7710, n7711, n7712, n7713, n7714, n7715,
    n7716, n7717, n7718, n7719, n7720, n7721,
    n7722, n7723, n7724, n7725, n7726, n7727,
    n7728, n7729, n7730, n7731, n7732, n7733,
    n7734, n7735, n7736, n7737, n7738, n7739,
    n7740, n7741, n7742, n7743, n7744, n7745,
    n7746, n7747, n7748, n7749, n7750, n7751,
    n7752, n7753, n7754, n7755, n7756, n7757,
    n7758, n7759, n7760, n7761, n7762, n7763,
    n7764, n7765, n7766, n7767, n7768, n7769,
    n7770, n7771, n7772, n7773, n7774, n7775,
    n7776, n7777, n7778, n7779, n7780, n7781,
    n7783, n7784, n7785, n7786, n7787, n7788,
    n7789, n7790, n7791, n7792, n7793, n7794,
    n7795, n7796, n7797, n7798, n7799, n7800,
    n7801, n7802, n7803, n7804, n7805, n7806,
    n7807, n7808, n7809, n7810, n7811, n7812,
    n7813, n7814, n7815, n7816, n7817, n7818,
    n7819, n7820, n7821, n7822, n7823, n7824,
    n7825, n7826, n7827, n7828, n7829, n7830,
    n7831, n7832, n7833, n7834, n7835, n7836,
    n7837, n7838, n7839, n7840, n7841, n7842,
    n7843, n7844, n7845, n7846, n7847, n7848,
    n7849, n7850, n7851, n7852, n7853, n7854,
    n7855, n7856, n7857, n7858, n7859, n7860,
    n7861, n7862, n7863, n7864, n7865, n7866,
    n7867, n7868, n7869, n7870, n7871, n7872,
    n7873, n7874, n7875, n7876, n7877, n7878,
    n7879, n7880, n7881, n7882, n7883, n7884,
    n7885, n7886, n7887, n7888, n7889, n7890,
    n7891, n7892, n7893, n7894, n7895, n7896,
    n7897, n7898, n7899, n7900, n7901, n7902,
    n7903, n7904, n7905, n7906, n7907, n7908,
    n7909, n7910, n7911, n7912, n7913, n7914,
    n7915, n7916, n7917, n7918, n7919, n7920,
    n7921, n7922, n7923, n7924, n7925, n7926,
    n7927, n7928, n7929, n7930, n7931, n7932,
    n7933, n7934, n7935, n7936, n7937, n7938,
    n7939, n7940, n7941, n7942, n7943, n7944,
    n7945, n7946, n7947, n7948, n7949, n7950,
    n7951, n7952, n7953, n7954, n7955, n7956,
    n7957, n7958, n7959, n7960, n7961, n7962,
    n7963, n7964, n7965, n7966, n7967, n7968,
    n7969, n7970, n7971, n7972, n7973, n7974,
    n7975, n7976, n7977, n7978, n7979, n7980,
    n7981, n7982, n7983, n7984, n7985, n7986,
    n7987, n7988, n7989, n7990, n7991, n7992,
    n7993, n7994, n7995, n7996, n7997, n7998,
    n7999, n8000, n8001, n8002, n8003, n8004,
    n8005, n8006, n8007, n8008, n8009, n8010,
    n8011, n8012, n8013, n8014, n8015, n8016,
    n8017, n8018, n8019, n8020, n8021, n8022,
    n8023, n8024, n8025, n8026, n8027, n8028,
    n8029, n8030, n8031, n8032, n8033, n8034,
    n8035, n8036, n8037, n8038, n8039, n8040,
    n8041, n8042, n8043, n8044, n8045, n8046,
    n8047, n8048, n8049, n8050, n8051, n8052,
    n8053, n8054, n8055, n8056, n8057, n8058,
    n8059, n8060, n8061, n8062, n8063, n8064,
    n8065, n8066, n8067, n8068, n8069, n8070,
    n8071, n8072, n8073, n8074, n8075, n8076,
    n8077, n8078, n8080, n8081, n8082, n8083,
    n8084, n8085, n8086, n8087, n8088, n8089,
    n8090, n8091, n8092, n8093, n8094, n8095,
    n8096, n8097, n8098, n8099, n8100, n8101,
    n8102, n8103, n8104, n8105, n8106, n8107,
    n8108, n8109, n8110, n8111, n8112, n8113,
    n8114, n8115, n8116, n8117, n8118, n8119,
    n8120, n8121, n8122, n8123, n8124, n8125,
    n8126, n8127, n8128, n8129, n8130, n8131,
    n8132, n8133, n8134, n8135, n8136, n8137,
    n8138, n8139, n8140, n8141, n8142, n8143,
    n8144, n8145, n8146, n8147, n8148, n8149,
    n8150, n8151, n8152, n8153, n8154, n8155,
    n8156, n8157, n8158, n8159, n8160, n8161,
    n8162, n8163, n8164, n8165, n8166, n8167,
    n8168, n8169, n8170, n8171, n8172, n8173,
    n8174, n8175, n8176, n8177, n8178, n8179,
    n8180, n8181, n8182, n8183, n8184, n8185,
    n8186, n8187, n8188, n8189, n8190, n8191,
    n8192, n8193, n8194, n8195, n8196, n8197,
    n8198, n8199, n8200, n8201, n8202, n8203,
    n8204, n8205, n8206, n8207, n8208, n8209,
    n8210, n8211, n8212, n8213, n8214, n8215,
    n8216, n8217, n8218, n8219, n8220, n8221,
    n8222, n8223, n8224, n8225, n8226, n8227,
    n8228, n8229, n8230, n8231, n8232, n8233,
    n8234, n8235, n8236, n8237, n8238, n8239,
    n8240, n8241, n8242, n8243, n8244, n8245,
    n8246, n8247, n8248, n8249, n8250, n8251,
    n8252, n8253, n8254, n8255, n8256, n8257,
    n8258, n8259, n8260, n8261, n8262, n8263,
    n8264, n8265, n8266, n8267, n8268, n8269,
    n8270, n8271, n8272, n8273, n8274, n8275,
    n8276, n8277, n8278, n8279, n8280, n8281,
    n8282, n8283, n8284, n8285, n8286, n8287,
    n8288, n8289, n8290, n8291, n8292, n8293,
    n8294, n8295, n8296, n8297, n8298, n8299,
    n8300, n8301, n8302, n8303, n8304, n8305,
    n8306, n8307, n8308, n8309, n8310, n8311,
    n8312, n8313, n8314, n8315, n8316, n8317,
    n8318, n8319, n8320, n8321, n8322, n8323,
    n8324, n8325, n8326, n8327, n8328, n8329,
    n8330, n8331, n8332, n8333, n8334, n8335,
    n8336, n8337, n8338, n8339, n8340, n8341,
    n8342, n8343, n8344, n8345, n8346, n8347,
    n8348, n8349, n8350, n8351, n8352, n8353,
    n8354, n8355, n8356, n8357, n8358, n8359,
    n8360, n8361, n8362, n8363, n8364, n8365,
    n8366, n8367, n8368, n8369, n8370, n8371,
    n8372, n8373, n8374, n8375, n8376, n8377,
    n8378, n8379, n8380, n8381, n8382, n8383,
    n8384, n8385, n8386, n8387, n8388, n8389,
    n8390, n8391, n8392, n8393, n8394, n8395,
    n8396, n8397, n8398, n8400, n8401, n8402,
    n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456,
    n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486,
    n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564,
    n8565, n8566, n8567, n8568, n8569, n8570,
    n8571, n8572, n8573, n8574, n8575, n8576,
    n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8593, n8594,
    n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606,
    n8607, n8608, n8609, n8610, n8611, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618,
    n8619, n8620, n8621, n8622, n8623, n8624,
    n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648,
    n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678,
    n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708,
    n8709, n8710, n8711, n8712, n8713, n8715,
    n8716, n8717, n8718, n8719, n8720, n8721,
    n8722, n8723, n8724, n8725, n8726, n8727,
    n8728, n8729, n8730, n8731, n8732, n8733,
    n8734, n8735, n8736, n8737, n8738, n8739,
    n8740, n8741, n8742, n8743, n8744, n8745,
    n8746, n8747, n8748, n8749, n8750, n8751,
    n8752, n8753, n8754, n8755, n8756, n8757,
    n8758, n8759, n8760, n8761, n8762, n8763,
    n8764, n8765, n8766, n8767, n8768, n8769,
    n8770, n8771, n8772, n8773, n8774, n8775,
    n8776, n8777, n8778, n8779, n8780, n8781,
    n8782, n8783, n8784, n8785, n8786, n8787,
    n8788, n8789, n8790, n8791, n8792, n8793,
    n8794, n8795, n8796, n8797, n8798, n8799,
    n8800, n8801, n8802, n8803, n8804, n8805,
    n8806, n8807, n8808, n8809, n8810, n8811,
    n8812, n8813, n8814, n8815, n8816, n8817,
    n8818, n8819, n8820, n8821, n8822, n8823,
    n8824, n8825, n8826, n8827, n8828, n8829,
    n8830, n8831, n8832, n8833, n8834, n8835,
    n8836, n8837, n8838, n8839, n8840, n8841,
    n8842, n8843, n8844, n8845, n8846, n8847,
    n8848, n8849, n8850, n8851, n8852, n8853,
    n8854, n8855, n8856, n8857, n8858, n8859,
    n8860, n8861, n8862, n8863, n8864, n8865,
    n8866, n8867, n8868, n8869, n8870, n8871,
    n8872, n8873, n8874, n8875, n8876, n8877,
    n8878, n8879, n8880, n8881, n8882, n8883,
    n8884, n8885, n8886, n8887, n8888, n8889,
    n8890, n8891, n8892, n8893, n8894, n8895,
    n8896, n8897, n8898, n8899, n8900, n8901,
    n8902, n8903, n8904, n8905, n8906, n8907,
    n8908, n8909, n8910, n8911, n8912, n8913,
    n8914, n8915, n8916, n8917, n8918, n8919,
    n8920, n8921, n8922, n8923, n8924, n8925,
    n8926, n8927, n8928, n8929, n8930, n8931,
    n8932, n8933, n8934, n8935, n8936, n8937,
    n8938, n8939, n8940, n8941, n8942, n8943,
    n8944, n8945, n8946, n8947, n8948, n8949,
    n8950, n8951, n8952, n8953, n8954, n8955,
    n8956, n8957, n8958, n8959, n8960, n8961,
    n8962, n8963, n8964, n8965, n8966, n8967,
    n8968, n8969, n8970, n8971, n8972, n8973,
    n8974, n8975, n8976, n8977, n8978, n8979,
    n8980, n8981, n8982, n8983, n8984, n8985,
    n8986, n8987, n8988, n8989, n8990, n8991,
    n8992, n8993, n8994, n8995, n8996, n8997,
    n8998, n8999, n9000, n9001, n9002, n9003,
    n9004, n9005, n9006, n9007, n9008, n9009,
    n9010, n9011, n9012, n9013, n9014, n9015,
    n9016, n9017, n9018, n9019, n9020, n9021,
    n9022, n9023, n9024, n9025, n9026, n9027,
    n9028, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040,
    n9041, n9042, n9043, n9044, n9045, n9046,
    n9047, n9048, n9049, n9050, n9051, n9052,
    n9053, n9054, n9055, n9056, n9057, n9058,
    n9059, n9060, n9061, n9062, n9063, n9064,
    n9065, n9066, n9067, n9068, n9069, n9070,
    n9071, n9072, n9073, n9074, n9075, n9076,
    n9077, n9078, n9079, n9080, n9081, n9082,
    n9083, n9084, n9085, n9086, n9087, n9088,
    n9089, n9090, n9091, n9092, n9093, n9094,
    n9095, n9096, n9097, n9098, n9099, n9100,
    n9101, n9102, n9103, n9104, n9105, n9106,
    n9107, n9108, n9109, n9110, n9111, n9112,
    n9113, n9114, n9115, n9116, n9117, n9118,
    n9119, n9120, n9121, n9122, n9123, n9124,
    n9125, n9126, n9127, n9128, n9129, n9130,
    n9131, n9132, n9133, n9134, n9135, n9136,
    n9137, n9138, n9139, n9140, n9141, n9142,
    n9143, n9144, n9145, n9146, n9147, n9148,
    n9149, n9150, n9151, n9152, n9153, n9154,
    n9155, n9156, n9157, n9158, n9159, n9160,
    n9161, n9162, n9163, n9164, n9165, n9166,
    n9167, n9168, n9169, n9170, n9171, n9172,
    n9173, n9174, n9175, n9176, n9177, n9178,
    n9179, n9180, n9181, n9182, n9183, n9184,
    n9185, n9186, n9187, n9188, n9189, n9190,
    n9191, n9192, n9193, n9194, n9195, n9196,
    n9197, n9198, n9199, n9200, n9201, n9202,
    n9203, n9204, n9205, n9206, n9207, n9208,
    n9209, n9210, n9211, n9212, n9213, n9214,
    n9215, n9216, n9217, n9218, n9219, n9220,
    n9221, n9222, n9223, n9224, n9225, n9226,
    n9227, n9228, n9229, n9230, n9231, n9232,
    n9233, n9234, n9235, n9236, n9237, n9238,
    n9239, n9240, n9241, n9242, n9243, n9244,
    n9245, n9246, n9247, n9248, n9249, n9250,
    n9251, n9252, n9253, n9254, n9255, n9256,
    n9257, n9258, n9259, n9260, n9261, n9262,
    n9263, n9264, n9265, n9266, n9267, n9268,
    n9269, n9270, n9271, n9272, n9273, n9274,
    n9275, n9276, n9277, n9278, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9286,
    n9287, n9288, n9289, n9290, n9291, n9292,
    n9293, n9294, n9295, n9296, n9297, n9298,
    n9299, n9300, n9301, n9302, n9303, n9304,
    n9305, n9306, n9307, n9308, n9309, n9310,
    n9311, n9312, n9313, n9314, n9315, n9316,
    n9317, n9318, n9319, n9320, n9321, n9322,
    n9323, n9324, n9325, n9326, n9327, n9328,
    n9329, n9330, n9331, n9332, n9333, n9334,
    n9335, n9336, n9337, n9338, n9339, n9340,
    n9341, n9342, n9343, n9344, n9345, n9346,
    n9347, n9348, n9349, n9350, n9351, n9352,
    n9353, n9354, n9355, n9356, n9357, n9358,
    n9359, n9360, n9361, n9362, n9363, n9364,
    n9365, n9366, n9367, n9368, n9369, n9371,
    n9372, n9373, n9374, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9382, n9383,
    n9384, n9385, n9386, n9387, n9388, n9389,
    n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401,
    n9402, n9403, n9404, n9405, n9406, n9407,
    n9408, n9409, n9410, n9411, n9412, n9413,
    n9414, n9415, n9416, n9417, n9418, n9419,
    n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431,
    n9432, n9433, n9434, n9435, n9436, n9437,
    n9438, n9439, n9440, n9441, n9442, n9443,
    n9444, n9445, n9446, n9447, n9448, n9449,
    n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461,
    n9462, n9463, n9464, n9465, n9466, n9467,
    n9468, n9469, n9470, n9471, n9472, n9473,
    n9474, n9475, n9476, n9477, n9478, n9479,
    n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491,
    n9492, n9493, n9494, n9495, n9496, n9497,
    n9498, n9499, n9500, n9501, n9502, n9503,
    n9504, n9505, n9506, n9507, n9508, n9509,
    n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521,
    n9522, n9523, n9524, n9525, n9526, n9527,
    n9528, n9529, n9530, n9531, n9532, n9533,
    n9534, n9535, n9536, n9537, n9538, n9539,
    n9540, n9541, n9542, n9543, n9544, n9545,
    n9546, n9547, n9548, n9549, n9550, n9551,
    n9552, n9553, n9554, n9555, n9556, n9557,
    n9558, n9559, n9560, n9561, n9562, n9563,
    n9564, n9565, n9566, n9567, n9568, n9569,
    n9570, n9571, n9572, n9573, n9574, n9575,
    n9576, n9577, n9578, n9579, n9580, n9581,
    n9582, n9583, n9584, n9585, n9586, n9587,
    n9588, n9589, n9590, n9591, n9592, n9593,
    n9594, n9595, n9596, n9597, n9598, n9599,
    n9600, n9601, n9602, n9603, n9604, n9605,
    n9606, n9607, n9608, n9609, n9610, n9611,
    n9612, n9613, n9614, n9615, n9616, n9617,
    n9618, n9619, n9620, n9621, n9622, n9623,
    n9624, n9625, n9626, n9627, n9628, n9629,
    n9630, n9631, n9632, n9633, n9634, n9635,
    n9636, n9637, n9638, n9639, n9640, n9641,
    n9642, n9643, n9644, n9645, n9646, n9647,
    n9648, n9649, n9650, n9651, n9652, n9653,
    n9654, n9655, n9656, n9657, n9658, n9659,
    n9660, n9661, n9662, n9663, n9664, n9665,
    n9666, n9667, n9668, n9669, n9670, n9671,
    n9672, n9673, n9674, n9675, n9676, n9677,
    n9678, n9679, n9680, n9681, n9682, n9683,
    n9684, n9685, n9686, n9687, n9688, n9689,
    n9690, n9691, n9692, n9693, n9694, n9695,
    n9696, n9697, n9698, n9699, n9700, n9701,
    n9702, n9704, n9705, n9706, n9707, n9708,
    n9709, n9710, n9711, n9712, n9713, n9714,
    n9715, n9716, n9717, n9718, n9719, n9720,
    n9721, n9722, n9723, n9724, n9725, n9726,
    n9727, n9728, n9729, n9730, n9731, n9732,
    n9733, n9734, n9735, n9736, n9737, n9738,
    n9739, n9740, n9741, n9742, n9743, n9744,
    n9745, n9746, n9747, n9748, n9749, n9750,
    n9751, n9752, n9753, n9754, n9755, n9756,
    n9757, n9758, n9759, n9760, n9761, n9762,
    n9763, n9764, n9765, n9766, n9767, n9768,
    n9769, n9770, n9771, n9772, n9773, n9774,
    n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786,
    n9787, n9788, n9789, n9790, n9791, n9792,
    n9793, n9794, n9795, n9796, n9797, n9798,
    n9799, n9800, n9801, n9802, n9803, n9804,
    n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9813, n9814, n9815, n9816,
    n9817, n9818, n9819, n9820, n9821, n9822,
    n9823, n9824, n9825, n9826, n9827, n9828,
    n9829, n9830, n9831, n9832, n9833, n9834,
    n9835, n9836, n9837, n9838, n9839, n9840,
    n9841, n9842, n9843, n9844, n9845, n9846,
    n9847, n9848, n9849, n9850, n9851, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858,
    n9859, n9860, n9861, n9862, n9863, n9864,
    n9865, n9866, n9867, n9868, n9869, n9870,
    n9871, n9872, n9873, n9874, n9875, n9876,
    n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888,
    n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900,
    n9901, n9902, n9903, n9904, n9905, n9906,
    n9907, n9908, n9909, n9910, n9911, n9912,
    n9913, n9914, n9915, n9916, n9917, n9918,
    n9919, n9920, n9921, n9922, n9923, n9924,
    n9925, n9926, n9927, n9928, n9929, n9930,
    n9931, n9932, n9933, n9934, n9935, n9936,
    n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948,
    n9949, n9950, n9951, n9952, n9953, n9954,
    n9955, n9956, n9957, n9958, n9959, n9960,
    n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990,
    n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10036, n10037, n10038, n10039,
    n10040, n10041, n10042, n10043, n10044, n10045,
    n10046, n10047, n10048, n10049, n10050, n10051,
    n10052, n10053, n10054, n10055, n10056, n10057,
    n10058, n10059, n10060, n10061, n10062, n10063,
    n10064, n10065, n10066, n10067, n10068, n10069,
    n10070, n10071, n10072, n10073, n10074, n10075,
    n10076, n10077, n10078, n10079, n10080, n10081,
    n10082, n10083, n10084, n10085, n10086, n10087,
    n10088, n10089, n10090, n10091, n10092, n10093,
    n10094, n10095, n10096, n10097, n10098, n10099,
    n10100, n10101, n10102, n10103, n10104, n10105,
    n10106, n10107, n10108, n10109, n10110, n10111,
    n10112, n10113, n10114, n10115, n10116, n10117,
    n10118, n10119, n10120, n10121, n10122, n10123,
    n10124, n10125, n10126, n10127, n10128, n10129,
    n10130, n10131, n10132, n10133, n10134, n10135,
    n10136, n10137, n10138, n10139, n10140, n10141,
    n10142, n10143, n10144, n10145, n10146, n10147,
    n10148, n10149, n10150, n10151, n10152, n10153,
    n10154, n10155, n10156, n10157, n10158, n10159,
    n10160, n10161, n10162, n10163, n10164, n10165,
    n10166, n10167, n10168, n10169, n10170, n10171,
    n10172, n10173, n10174, n10175, n10176, n10177,
    n10178, n10179, n10180, n10181, n10182, n10183,
    n10184, n10185, n10186, n10187, n10188, n10189,
    n10190, n10191, n10192, n10193, n10194, n10195,
    n10196, n10197, n10198, n10199, n10200, n10201,
    n10202, n10203, n10204, n10205, n10206, n10207,
    n10208, n10209, n10210, n10211, n10212, n10213,
    n10214, n10215, n10216, n10217, n10218, n10219,
    n10220, n10221, n10222, n10223, n10224, n10225,
    n10226, n10227, n10228, n10229, n10230, n10231,
    n10232, n10233, n10234, n10235, n10236, n10237,
    n10238, n10239, n10240, n10241, n10242, n10243,
    n10244, n10245, n10246, n10247, n10248, n10249,
    n10250, n10251, n10252, n10253, n10254, n10255,
    n10256, n10257, n10258, n10259, n10260, n10261,
    n10262, n10263, n10264, n10265, n10266, n10267,
    n10268, n10269, n10270, n10271, n10272, n10273,
    n10274, n10275, n10276, n10277, n10278, n10279,
    n10280, n10281, n10282, n10283, n10284, n10285,
    n10286, n10287, n10288, n10289, n10290, n10291,
    n10292, n10293, n10294, n10295, n10296, n10297,
    n10298, n10299, n10300, n10301, n10302, n10303,
    n10304, n10305, n10306, n10307, n10308, n10309,
    n10310, n10311, n10312, n10313, n10314, n10315,
    n10316, n10317, n10318, n10319, n10320, n10321,
    n10322, n10323, n10324, n10325, n10326, n10327,
    n10328, n10329, n10330, n10331, n10332, n10333,
    n10334, n10335, n10336, n10337, n10338, n10339,
    n10340, n10341, n10342, n10343, n10344, n10345,
    n10346, n10347, n10348, n10349, n10350, n10351,
    n10352, n10353, n10354, n10355, n10356, n10357,
    n10358, n10359, n10360, n10361, n10362, n10363,
    n10364, n10365, n10366, n10367, n10368, n10369,
    n10370, n10371, n10372, n10373, n10374, n10375,
    n10376, n10377, n10378, n10379, n10380, n10381,
    n10382, n10383, n10384, n10385, n10386, n10387,
    n10388, n10389, n10390, n10391, n10392, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406,
    n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424,
    n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442,
    n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460,
    n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472,
    n10473, n10474, n10475, n10476, n10477, n10478,
    n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490,
    n10491, n10492, n10493, n10494, n10495, n10496,
    n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514,
    n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532,
    n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10546, n10547, n10548, n10549, n10550,
    n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562,
    n10563, n10564, n10565, n10566, n10567, n10568,
    n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580,
    n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598,
    n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10651, n10652,
    n10653, n10654, n10655, n10656, n10657, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664,
    n10665, n10666, n10667, n10668, n10669, n10670,
    n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706,
    n10707, n10708, n10709, n10710, n10711, n10712,
    n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724,
    n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742,
    n10743, n10744, n10745, n10747, n10748, n10749,
    n10750, n10751, n10752, n10753, n10754, n10755,
    n10756, n10757, n10758, n10759, n10760, n10761,
    n10762, n10763, n10764, n10765, n10766, n10767,
    n10768, n10769, n10770, n10771, n10772, n10773,
    n10774, n10775, n10776, n10777, n10778, n10779,
    n10780, n10781, n10782, n10783, n10784, n10785,
    n10786, n10787, n10788, n10789, n10790, n10791,
    n10792, n10793, n10794, n10795, n10796, n10797,
    n10798, n10799, n10800, n10801, n10802, n10803,
    n10804, n10805, n10806, n10807, n10808, n10809,
    n10810, n10811, n10812, n10813, n10814, n10815,
    n10816, n10817, n10818, n10819, n10820, n10821,
    n10822, n10823, n10824, n10825, n10826, n10827,
    n10828, n10829, n10830, n10831, n10832, n10833,
    n10834, n10835, n10836, n10837, n10838, n10839,
    n10840, n10841, n10842, n10843, n10844, n10845,
    n10846, n10847, n10848, n10849, n10850, n10851,
    n10852, n10853, n10854, n10855, n10856, n10857,
    n10858, n10859, n10860, n10861, n10862, n10863,
    n10864, n10865, n10866, n10867, n10868, n10869,
    n10870, n10871, n10872, n10873, n10874, n10875,
    n10876, n10877, n10878, n10879, n10880, n10881,
    n10882, n10883, n10884, n10885, n10886, n10887,
    n10888, n10889, n10890, n10891, n10892, n10893,
    n10894, n10895, n10896, n10897, n10898, n10899,
    n10900, n10901, n10902, n10903, n10904, n10905,
    n10906, n10907, n10908, n10909, n10910, n10911,
    n10912, n10913, n10914, n10915, n10916, n10917,
    n10918, n10919, n10920, n10921, n10922, n10923,
    n10924, n10925, n10926, n10927, n10928, n10929,
    n10930, n10931, n10932, n10933, n10934, n10935,
    n10936, n10937, n10938, n10939, n10940, n10941,
    n10942, n10943, n10944, n10945, n10946, n10947,
    n10948, n10949, n10950, n10951, n10952, n10953,
    n10954, n10955, n10956, n10957, n10958, n10959,
    n10960, n10961, n10962, n10963, n10964, n10965,
    n10966, n10967, n10968, n10969, n10970, n10971,
    n10972, n10973, n10974, n10975, n10976, n10977,
    n10978, n10979, n10980, n10981, n10982, n10983,
    n10984, n10985, n10986, n10987, n10988, n10989,
    n10990, n10991, n10992, n10993, n10994, n10995,
    n10996, n10997, n10998, n10999, n11000, n11001,
    n11002, n11003, n11004, n11005, n11006, n11007,
    n11008, n11009, n11010, n11011, n11012, n11013,
    n11014, n11015, n11016, n11017, n11018, n11019,
    n11020, n11021, n11022, n11023, n11024, n11025,
    n11026, n11027, n11028, n11029, n11030, n11031,
    n11032, n11033, n11034, n11035, n11036, n11037,
    n11038, n11039, n11040, n11041, n11042, n11043,
    n11044, n11045, n11046, n11047, n11048, n11049,
    n11050, n11051, n11052, n11053, n11054, n11055,
    n11056, n11057, n11058, n11059, n11060, n11061,
    n11062, n11063, n11064, n11065, n11066, n11067,
    n11068, n11069, n11070, n11071, n11072, n11073,
    n11074, n11075, n11076, n11077, n11078, n11079,
    n11080, n11081, n11082, n11083, n11084, n11085,
    n11086, n11087, n11088, n11089, n11090, n11091,
    n11092, n11093, n11094, n11095, n11096, n11097,
    n11099, n11100, n11101, n11102, n11103, n11104,
    n11105, n11106, n11107, n11108, n11109, n11110,
    n11111, n11112, n11113, n11114, n11115, n11116,
    n11117, n11118, n11119, n11120, n11121, n11122,
    n11123, n11124, n11125, n11126, n11127, n11128,
    n11129, n11130, n11131, n11132, n11133, n11134,
    n11135, n11136, n11137, n11138, n11139, n11140,
    n11141, n11142, n11143, n11144, n11145, n11146,
    n11147, n11148, n11149, n11150, n11151, n11152,
    n11153, n11154, n11155, n11156, n11157, n11158,
    n11159, n11160, n11161, n11162, n11163, n11164,
    n11165, n11166, n11167, n11168, n11169, n11170,
    n11171, n11172, n11173, n11174, n11175, n11176,
    n11177, n11178, n11179, n11180, n11181, n11182,
    n11183, n11184, n11185, n11186, n11187, n11188,
    n11189, n11190, n11191, n11192, n11193, n11194,
    n11195, n11196, n11197, n11198, n11199, n11200,
    n11201, n11202, n11203, n11204, n11205, n11206,
    n11207, n11208, n11209, n11210, n11211, n11212,
    n11213, n11214, n11215, n11216, n11217, n11218,
    n11219, n11220, n11221, n11222, n11223, n11224,
    n11225, n11226, n11227, n11228, n11229, n11230,
    n11231, n11232, n11233, n11234, n11235, n11236,
    n11237, n11238, n11239, n11240, n11241, n11242,
    n11243, n11244, n11245, n11246, n11247, n11248,
    n11249, n11250, n11251, n11252, n11253, n11254,
    n11255, n11256, n11257, n11258, n11259, n11260,
    n11261, n11262, n11263, n11264, n11265, n11266,
    n11267, n11268, n11269, n11270, n11271, n11272,
    n11273, n11274, n11275, n11276, n11277, n11278,
    n11279, n11280, n11281, n11282, n11283, n11284,
    n11285, n11286, n11287, n11288, n11289, n11290,
    n11291, n11292, n11293, n11294, n11295, n11296,
    n11297, n11298, n11299, n11300, n11301, n11302,
    n11303, n11304, n11305, n11306, n11307, n11308,
    n11309, n11310, n11311, n11312, n11313, n11314,
    n11315, n11316, n11317, n11318, n11319, n11320,
    n11321, n11322, n11323, n11324, n11325, n11326,
    n11327, n11328, n11329, n11330, n11331, n11332,
    n11333, n11334, n11335, n11336, n11337, n11338,
    n11339, n11340, n11341, n11342, n11343, n11344,
    n11345, n11346, n11347, n11348, n11349, n11350,
    n11351, n11352, n11353, n11354, n11355, n11356,
    n11357, n11358, n11359, n11360, n11361, n11362,
    n11363, n11364, n11365, n11366, n11367, n11368,
    n11369, n11370, n11371, n11372, n11373, n11374,
    n11375, n11376, n11377, n11378, n11379, n11380,
    n11381, n11382, n11383, n11384, n11385, n11386,
    n11387, n11388, n11389, n11390, n11391, n11392,
    n11393, n11394, n11395, n11396, n11397, n11398,
    n11399, n11400, n11401, n11402, n11403, n11404,
    n11405, n11406, n11407, n11408, n11409, n11410,
    n11411, n11412, n11413, n11414, n11415, n11416,
    n11417, n11418, n11419, n11420, n11421, n11422,
    n11423, n11424, n11425, n11426, n11427, n11428,
    n11429, n11430, n11431, n11432, n11433, n11434,
    n11435, n11436, n11437, n11438, n11439, n11440,
    n11441, n11442, n11443, n11444, n11445, n11446,
    n11447, n11448, n11449, n11450, n11451, n11452,
    n11453, n11454, n11455, n11456, n11457, n11458,
    n11459, n11460, n11461, n11462, n11463, n11464,
    n11465, n11466, n11467, n11468, n11469, n11470,
    n11471, n11472, n11473, n11474, n11476, n11477,
    n11478, n11479, n11480, n11481, n11482, n11483,
    n11484, n11485, n11486, n11487, n11488, n11489,
    n11490, n11491, n11492, n11493, n11494, n11495,
    n11496, n11497, n11498, n11499, n11500, n11501,
    n11502, n11503, n11504, n11505, n11506, n11507,
    n11508, n11509, n11510, n11511, n11512, n11513,
    n11514, n11515, n11516, n11517, n11518, n11519,
    n11520, n11521, n11522, n11523, n11524, n11525,
    n11526, n11527, n11528, n11529, n11530, n11531,
    n11532, n11533, n11534, n11535, n11536, n11537,
    n11538, n11539, n11540, n11541, n11542, n11543,
    n11544, n11545, n11546, n11547, n11548, n11549,
    n11550, n11551, n11552, n11553, n11554, n11555,
    n11556, n11557, n11558, n11559, n11560, n11561,
    n11562, n11563, n11564, n11565, n11566, n11567,
    n11568, n11569, n11570, n11571, n11572, n11573,
    n11574, n11575, n11576, n11577, n11578, n11579,
    n11580, n11581, n11582, n11583, n11584, n11585,
    n11586, n11587, n11588, n11589, n11590, n11591,
    n11592, n11593, n11594, n11595, n11596, n11597,
    n11598, n11599, n11600, n11601, n11602, n11603,
    n11604, n11605, n11606, n11607, n11608, n11609,
    n11610, n11611, n11612, n11613, n11614, n11615,
    n11616, n11617, n11618, n11619, n11620, n11621,
    n11622, n11623, n11624, n11625, n11626, n11627,
    n11628, n11629, n11630, n11631, n11632, n11633,
    n11634, n11635, n11636, n11637, n11638, n11639,
    n11640, n11641, n11642, n11643, n11644, n11645,
    n11646, n11647, n11648, n11649, n11650, n11651,
    n11652, n11653, n11654, n11655, n11656, n11657,
    n11658, n11659, n11660, n11661, n11662, n11663,
    n11664, n11665, n11666, n11667, n11668, n11669,
    n11670, n11671, n11672, n11673, n11674, n11675,
    n11676, n11677, n11678, n11679, n11680, n11681,
    n11682, n11683, n11684, n11685, n11686, n11687,
    n11688, n11689, n11690, n11691, n11692, n11693,
    n11694, n11695, n11696, n11697, n11698, n11699,
    n11700, n11701, n11702, n11703, n11704, n11705,
    n11706, n11707, n11708, n11709, n11710, n11711,
    n11712, n11713, n11714, n11715, n11716, n11717,
    n11718, n11719, n11720, n11721, n11722, n11723,
    n11724, n11725, n11726, n11727, n11728, n11729,
    n11730, n11731, n11732, n11733, n11734, n11735,
    n11736, n11737, n11738, n11739, n11740, n11741,
    n11742, n11743, n11744, n11745, n11746, n11747,
    n11748, n11749, n11750, n11751, n11752, n11753,
    n11754, n11755, n11756, n11757, n11758, n11759,
    n11760, n11761, n11762, n11763, n11764, n11765,
    n11766, n11767, n11768, n11769, n11770, n11771,
    n11772, n11773, n11774, n11775, n11776, n11777,
    n11778, n11779, n11780, n11781, n11782, n11783,
    n11784, n11785, n11786, n11787, n11788, n11789,
    n11790, n11791, n11792, n11793, n11794, n11795,
    n11796, n11797, n11798, n11799, n11800, n11801,
    n11802, n11803, n11804, n11805, n11806, n11807,
    n11808, n11809, n11810, n11811, n11812, n11813,
    n11814, n11815, n11816, n11817, n11818, n11819,
    n11820, n11821, n11822, n11823, n11824, n11825,
    n11826, n11827, n11828, n11829, n11830, n11831,
    n11832, n11833, n11834, n11835, n11836, n11837,
    n11838, n11839, n11840, n11841, n11842, n11843,
    n11845, n11846, n11847, n11848, n11849, n11850,
    n11851, n11852, n11853, n11854, n11855, n11856,
    n11857, n11858, n11859, n11860, n11861, n11862,
    n11863, n11864, n11865, n11866, n11867, n11868,
    n11869, n11870, n11871, n11872, n11873, n11874,
    n11875, n11876, n11877, n11878, n11879, n11880,
    n11881, n11882, n11883, n11884, n11885, n11886,
    n11887, n11888, n11889, n11890, n11891, n11892,
    n11893, n11894, n11895, n11896, n11897, n11898,
    n11899, n11900, n11901, n11902, n11903, n11904,
    n11905, n11906, n11907, n11908, n11909, n11910,
    n11911, n11912, n11913, n11914, n11915, n11916,
    n11917, n11918, n11919, n11920, n11921, n11922,
    n11923, n11924, n11925, n11926, n11927, n11928,
    n11929, n11930, n11931, n11932, n11933, n11934,
    n11935, n11936, n11937, n11938, n11939, n11940,
    n11941, n11942, n11943, n11944, n11945, n11946,
    n11947, n11948, n11949, n11950, n11951, n11952,
    n11953, n11954, n11955, n11956, n11957, n11958,
    n11959, n11960, n11961, n11962, n11963, n11964,
    n11965, n11966, n11967, n11968, n11969, n11970,
    n11971, n11972, n11973, n11974, n11975, n11976,
    n11977, n11978, n11979, n11980, n11981, n11982,
    n11983, n11984, n11985, n11986, n11987, n11988,
    n11989, n11990, n11991, n11992, n11993, n11994,
    n11995, n11996, n11997, n11998, n11999, n12000,
    n12001, n12002, n12003, n12004, n12005, n12006,
    n12007, n12008, n12009, n12010, n12011, n12012,
    n12013, n12014, n12015, n12016, n12017, n12018,
    n12019, n12020, n12021, n12022, n12023, n12024,
    n12025, n12026, n12027, n12028, n12029, n12030,
    n12031, n12032, n12033, n12034, n12035, n12036,
    n12037, n12038, n12039, n12040, n12041, n12042,
    n12043, n12044, n12045, n12046, n12047, n12048,
    n12049, n12050, n12051, n12052, n12053, n12054,
    n12055, n12056, n12057, n12058, n12059, n12060,
    n12061, n12062, n12063, n12064, n12065, n12066,
    n12067, n12068, n12069, n12070, n12071, n12072,
    n12073, n12074, n12075, n12076, n12077, n12078,
    n12079, n12080, n12081, n12082, n12083, n12084,
    n12085, n12086, n12087, n12088, n12089, n12090,
    n12091, n12092, n12093, n12094, n12095, n12096,
    n12097, n12098, n12099, n12100, n12101, n12102,
    n12103, n12104, n12105, n12106, n12107, n12108,
    n12109, n12110, n12111, n12112, n12113, n12114,
    n12115, n12116, n12117, n12118, n12119, n12120,
    n12121, n12122, n12123, n12124, n12125, n12126,
    n12127, n12128, n12129, n12130, n12131, n12132,
    n12133, n12134, n12135, n12136, n12137, n12138,
    n12139, n12140, n12141, n12142, n12143, n12144,
    n12145, n12146, n12147, n12148, n12149, n12150,
    n12151, n12152, n12153, n12154, n12155, n12156,
    n12157, n12158, n12159, n12160, n12161, n12162,
    n12163, n12164, n12165, n12166, n12167, n12168,
    n12169, n12170, n12171, n12172, n12173, n12174,
    n12175, n12176, n12177, n12178, n12179, n12180,
    n12181, n12182, n12183, n12184, n12185, n12186,
    n12187, n12188, n12189, n12190, n12191, n12192,
    n12193, n12194, n12195, n12196, n12197, n12198,
    n12199, n12200, n12201, n12202, n12203, n12204,
    n12205, n12206, n12207, n12208, n12209, n12210,
    n12211, n12213, n12214, n12215, n12216, n12217,
    n12218, n12219, n12220, n12221, n12222, n12223,
    n12224, n12225, n12226, n12227, n12228, n12229,
    n12230, n12231, n12232, n12233, n12234, n12235,
    n12236, n12237, n12238, n12239, n12240, n12241,
    n12242, n12243, n12244, n12245, n12246, n12247,
    n12248, n12249, n12250, n12251, n12252, n12253,
    n12254, n12255, n12256, n12257, n12258, n12259,
    n12260, n12261, n12262, n12263, n12264, n12265,
    n12266, n12267, n12268, n12269, n12270, n12271,
    n12272, n12273, n12274, n12275, n12276, n12277,
    n12278, n12279, n12280, n12281, n12282, n12283,
    n12284, n12285, n12286, n12287, n12288, n12289,
    n12290, n12291, n12292, n12293, n12294, n12295,
    n12296, n12297, n12298, n12299, n12300, n12301,
    n12302, n12303, n12304, n12305, n12306, n12307,
    n12308, n12309, n12310, n12311, n12312, n12313,
    n12314, n12315, n12316, n12317, n12318, n12319,
    n12320, n12321, n12322, n12323, n12324, n12325,
    n12326, n12327, n12328, n12329, n12330, n12331,
    n12332, n12333, n12334, n12335, n12336, n12337,
    n12338, n12339, n12340, n12341, n12342, n12343,
    n12344, n12345, n12346, n12347, n12348, n12349,
    n12350, n12351, n12352, n12353, n12354, n12355,
    n12356, n12357, n12358, n12359, n12360, n12361,
    n12362, n12363, n12364, n12365, n12366, n12367,
    n12368, n12369, n12370, n12371, n12372, n12373,
    n12374, n12375, n12376, n12377, n12378, n12379,
    n12380, n12381, n12382, n12383, n12384, n12385,
    n12386, n12387, n12388, n12389, n12390, n12391,
    n12392, n12393, n12394, n12395, n12396, n12397,
    n12398, n12399, n12400, n12401, n12402, n12403,
    n12404, n12405, n12406, n12407, n12408, n12409,
    n12410, n12411, n12412, n12413, n12414, n12415,
    n12416, n12417, n12418, n12419, n12420, n12421,
    n12422, n12423, n12424, n12425, n12426, n12427,
    n12428, n12429, n12430, n12431, n12432, n12433,
    n12434, n12435, n12436, n12437, n12438, n12439,
    n12440, n12441, n12442, n12443, n12444, n12445,
    n12446, n12447, n12448, n12449, n12450, n12451,
    n12452, n12453, n12454, n12455, n12456, n12457,
    n12458, n12459, n12460, n12461, n12462, n12463,
    n12464, n12465, n12466, n12467, n12468, n12469,
    n12470, n12471, n12472, n12473, n12474, n12475,
    n12476, n12477, n12478, n12479, n12480, n12481,
    n12482, n12483, n12484, n12485, n12486, n12487,
    n12488, n12489, n12490, n12491, n12492, n12493,
    n12494, n12495, n12496, n12497, n12498, n12499,
    n12500, n12501, n12502, n12503, n12504, n12505,
    n12506, n12507, n12508, n12509, n12510, n12511,
    n12512, n12513, n12514, n12515, n12516, n12517,
    n12518, n12519, n12520, n12521, n12522, n12523,
    n12524, n12525, n12526, n12527, n12528, n12529,
    n12530, n12531, n12532, n12533, n12534, n12535,
    n12536, n12537, n12538, n12539, n12540, n12541,
    n12542, n12543, n12544, n12545, n12546, n12547,
    n12548, n12549, n12550, n12551, n12552, n12553,
    n12554, n12555, n12556, n12557, n12558, n12559,
    n12560, n12561, n12562, n12563, n12564, n12565,
    n12566, n12567, n12568, n12569, n12570, n12571,
    n12572, n12573, n12574, n12575, n12576, n12577,
    n12578, n12579, n12580, n12581, n12582, n12583,
    n12584, n12585, n12586, n12587, n12588, n12589,
    n12590, n12591, n12592, n12593, n12594, n12595,
    n12596, n12597, n12598, n12599, n12600, n12601,
    n12602, n12603, n12604, n12605, n12606, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614,
    n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632,
    n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650,
    n12651, n12652, n12653, n12654, n12655, n12656,
    n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668,
    n12669, n12670, n12671, n12672, n12673, n12674,
    n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12691, n12692,
    n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704,
    n12705, n12706, n12707, n12708, n12709, n12710,
    n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722,
    n12723, n12724, n12725, n12726, n12727, n12728,
    n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740,
    n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758,
    n12759, n12760, n12761, n12762, n12763, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776,
    n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794,
    n12795, n12796, n12797, n12798, n12799, n12800,
    n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812,
    n12813, n12814, n12815, n12816, n12817, n12818,
    n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12830,
    n12831, n12832, n12833, n12834, n12835, n12836,
    n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848,
    n12849, n12850, n12851, n12852, n12853, n12854,
    n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866,
    n12867, n12868, n12869, n12870, n12871, n12872,
    n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884,
    n12885, n12886, n12887, n12888, n12889, n12890,
    n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902,
    n12903, n12904, n12905, n12906, n12907, n12908,
    n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920,
    n12921, n12922, n12923, n12924, n12925, n12926,
    n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938,
    n12939, n12940, n12941, n12942, n12943, n12944,
    n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956,
    n12957, n12958, n12959, n12960, n12961, n12962,
    n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974,
    n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12995, n12996, n12997, n12998, n12999,
    n13000, n13001, n13002, n13003, n13004, n13005,
    n13006, n13007, n13008, n13009, n13010, n13011,
    n13012, n13013, n13014, n13015, n13016, n13017,
    n13018, n13019, n13020, n13021, n13022, n13023,
    n13024, n13025, n13026, n13027, n13028, n13029,
    n13030, n13031, n13032, n13033, n13034, n13035,
    n13036, n13037, n13038, n13039, n13040, n13041,
    n13042, n13043, n13044, n13045, n13046, n13047,
    n13048, n13049, n13050, n13051, n13052, n13053,
    n13054, n13055, n13056, n13057, n13058, n13059,
    n13060, n13061, n13062, n13063, n13064, n13065,
    n13066, n13067, n13068, n13069, n13070, n13071,
    n13072, n13073, n13074, n13075, n13076, n13077,
    n13078, n13079, n13080, n13081, n13082, n13083,
    n13084, n13085, n13086, n13087, n13088, n13089,
    n13090, n13091, n13092, n13093, n13094, n13095,
    n13096, n13097, n13098, n13099, n13100, n13101,
    n13102, n13103, n13104, n13105, n13106, n13107,
    n13108, n13109, n13110, n13111, n13112, n13113,
    n13114, n13115, n13116, n13117, n13118, n13119,
    n13120, n13121, n13122, n13123, n13124, n13125,
    n13126, n13127, n13128, n13129, n13130, n13131,
    n13132, n13133, n13134, n13135, n13136, n13137,
    n13138, n13139, n13140, n13141, n13142, n13143,
    n13144, n13145, n13146, n13147, n13148, n13149,
    n13150, n13151, n13152, n13153, n13154, n13155,
    n13156, n13157, n13158, n13159, n13160, n13161,
    n13162, n13163, n13164, n13165, n13166, n13167,
    n13168, n13169, n13170, n13171, n13172, n13173,
    n13174, n13175, n13176, n13177, n13178, n13179,
    n13180, n13181, n13182, n13183, n13184, n13185,
    n13186, n13187, n13188, n13189, n13190, n13191,
    n13192, n13193, n13194, n13195, n13196, n13197,
    n13198, n13199, n13200, n13201, n13202, n13203,
    n13204, n13205, n13206, n13207, n13208, n13209,
    n13210, n13211, n13212, n13213, n13214, n13215,
    n13216, n13217, n13218, n13219, n13220, n13221,
    n13222, n13223, n13224, n13225, n13226, n13227,
    n13228, n13229, n13230, n13231, n13232, n13233,
    n13234, n13235, n13236, n13237, n13238, n13239,
    n13240, n13241, n13242, n13243, n13244, n13245,
    n13246, n13247, n13248, n13249, n13250, n13251,
    n13252, n13253, n13254, n13255, n13256, n13257,
    n13258, n13259, n13260, n13261, n13262, n13263,
    n13264, n13265, n13266, n13267, n13268, n13269,
    n13270, n13271, n13272, n13273, n13274, n13275,
    n13276, n13277, n13278, n13279, n13280, n13281,
    n13282, n13283, n13284, n13285, n13286, n13287,
    n13288, n13289, n13290, n13291, n13292, n13293,
    n13294, n13295, n13296, n13297, n13298, n13299,
    n13300, n13301, n13302, n13303, n13304, n13305,
    n13306, n13307, n13308, n13309, n13310, n13311,
    n13312, n13313, n13314, n13315, n13316, n13317,
    n13318, n13319, n13320, n13321, n13322, n13323,
    n13324, n13325, n13326, n13327, n13328, n13329,
    n13330, n13331, n13332, n13333, n13334, n13335,
    n13336, n13337, n13338, n13339, n13340, n13341,
    n13342, n13343, n13344, n13345, n13346, n13347,
    n13348, n13349, n13350, n13351, n13352, n13353,
    n13354, n13355, n13356, n13357, n13358, n13359,
    n13360, n13361, n13362, n13363, n13364, n13365,
    n13366, n13367, n13368, n13369, n13370, n13371,
    n13372, n13373, n13374, n13375, n13376, n13377,
    n13378, n13379, n13381, n13382, n13383, n13384,
    n13385, n13386, n13387, n13388, n13389, n13390,
    n13391, n13392, n13393, n13394, n13395, n13396,
    n13397, n13398, n13399, n13400, n13401, n13402,
    n13403, n13404, n13405, n13406, n13407, n13408,
    n13409, n13410, n13411, n13412, n13413, n13414,
    n13415, n13416, n13417, n13418, n13419, n13420,
    n13421, n13422, n13423, n13424, n13425, n13426,
    n13427, n13428, n13429, n13430, n13431, n13432,
    n13433, n13434, n13435, n13436, n13437, n13438,
    n13439, n13440, n13441, n13442, n13443, n13444,
    n13445, n13446, n13447, n13448, n13449, n13450,
    n13451, n13452, n13453, n13454, n13455, n13456,
    n13457, n13458, n13459, n13460, n13461, n13462,
    n13463, n13464, n13465, n13466, n13467, n13468,
    n13469, n13470, n13471, n13472, n13473, n13474,
    n13475, n13476, n13477, n13478, n13479, n13480,
    n13481, n13482, n13483, n13484, n13485, n13486,
    n13487, n13488, n13489, n13490, n13491, n13492,
    n13493, n13494, n13495, n13496, n13497, n13498,
    n13499, n13500, n13501, n13502, n13503, n13504,
    n13505, n13506, n13507, n13508, n13509, n13510,
    n13511, n13512, n13513, n13514, n13515, n13516,
    n13517, n13518, n13519, n13520, n13521, n13522,
    n13523, n13524, n13525, n13526, n13527, n13528,
    n13529, n13530, n13531, n13532, n13533, n13534,
    n13535, n13536, n13537, n13538, n13539, n13540,
    n13541, n13542, n13543, n13544, n13545, n13546,
    n13547, n13548, n13549, n13550, n13551, n13552,
    n13553, n13554, n13555, n13556, n13557, n13558,
    n13559, n13560, n13561, n13562, n13563, n13564,
    n13565, n13566, n13567, n13568, n13569, n13570,
    n13571, n13572, n13573, n13574, n13575, n13576,
    n13577, n13578, n13579, n13580, n13581, n13582,
    n13583, n13584, n13585, n13586, n13587, n13588,
    n13589, n13590, n13591, n13592, n13593, n13594,
    n13595, n13596, n13597, n13598, n13599, n13600,
    n13601, n13602, n13603, n13604, n13605, n13606,
    n13607, n13608, n13609, n13610, n13611, n13612,
    n13613, n13614, n13615, n13616, n13617, n13618,
    n13619, n13620, n13621, n13622, n13623, n13624,
    n13625, n13626, n13627, n13628, n13629, n13630,
    n13631, n13632, n13633, n13634, n13635, n13636,
    n13637, n13638, n13639, n13640, n13641, n13642,
    n13643, n13644, n13645, n13646, n13647, n13648,
    n13649, n13650, n13651, n13652, n13653, n13654,
    n13655, n13656, n13657, n13658, n13659, n13660,
    n13661, n13662, n13663, n13664, n13665, n13666,
    n13667, n13668, n13669, n13670, n13671, n13672,
    n13673, n13674, n13675, n13676, n13677, n13678,
    n13679, n13680, n13681, n13682, n13683, n13684,
    n13685, n13686, n13687, n13688, n13689, n13690,
    n13691, n13692, n13693, n13694, n13695, n13696,
    n13697, n13698, n13699, n13700, n13701, n13702,
    n13703, n13704, n13705, n13706, n13707, n13708,
    n13709, n13710, n13711, n13712, n13713, n13714,
    n13715, n13716, n13717, n13718, n13719, n13720,
    n13721, n13722, n13723, n13724, n13725, n13726,
    n13727, n13728, n13729, n13730, n13731, n13732,
    n13733, n13734, n13735, n13736, n13737, n13738,
    n13739, n13740, n13741, n13742, n13743, n13744,
    n13745, n13746, n13747, n13748, n13749, n13750,
    n13751, n13752, n13753, n13754, n13755, n13756,
    n13757, n13758, n13759, n13760, n13761, n13762,
    n13763, n13764, n13766, n13767, n13768, n13769,
    n13770, n13771, n13772, n13773, n13774, n13775,
    n13776, n13777, n13778, n13779, n13780, n13781,
    n13782, n13783, n13784, n13785, n13786, n13787,
    n13788, n13789, n13790, n13791, n13792, n13793,
    n13794, n13795, n13796, n13797, n13798, n13799,
    n13800, n13801, n13802, n13803, n13804, n13805,
    n13806, n13807, n13808, n13809, n13810, n13811,
    n13812, n13813, n13814, n13815, n13816, n13817,
    n13818, n13819, n13820, n13821, n13822, n13823,
    n13824, n13825, n13826, n13827, n13828, n13829,
    n13830, n13831, n13832, n13833, n13834, n13835,
    n13836, n13837, n13838, n13839, n13840, n13841,
    n13842, n13843, n13844, n13845, n13846, n13847,
    n13848, n13849, n13850, n13851, n13852, n13853,
    n13854, n13855, n13856, n13857, n13858, n13859,
    n13860, n13861, n13862, n13863, n13864, n13865,
    n13866, n13867, n13868, n13869, n13870, n13871,
    n13872, n13873, n13874, n13875, n13876, n13877,
    n13878, n13879, n13880, n13881, n13882, n13883,
    n13884, n13885, n13886, n13887, n13888, n13889,
    n13890, n13891, n13892, n13893, n13894, n13895,
    n13896, n13897, n13898, n13899, n13900, n13901,
    n13902, n13903, n13904, n13905, n13906, n13907,
    n13908, n13909, n13910, n13911, n13912, n13913,
    n13914, n13915, n13916, n13917, n13918, n13919,
    n13920, n13921, n13922, n13923, n13924, n13925,
    n13926, n13927, n13928, n13929, n13930, n13931,
    n13932, n13933, n13934, n13935, n13936, n13937,
    n13938, n13939, n13940, n13941, n13942, n13943,
    n13944, n13945, n13946, n13947, n13948, n13949,
    n13950, n13951, n13952, n13953, n13954, n13955,
    n13956, n13957, n13958, n13959, n13960, n13961,
    n13962, n13963, n13964, n13965, n13966, n13967,
    n13968, n13969, n13970, n13971, n13972, n13973,
    n13974, n13975, n13976, n13977, n13978, n13979,
    n13980, n13981, n13982, n13983, n13984, n13985,
    n13986, n13987, n13988, n13989, n13990, n13991,
    n13992, n13993, n13994, n13995, n13996, n13997,
    n13998, n13999, n14000, n14001, n14002, n14003,
    n14004, n14005, n14006, n14007, n14008, n14009,
    n14010, n14011, n14012, n14013, n14014, n14015,
    n14016, n14017, n14018, n14019, n14020, n14021,
    n14022, n14023, n14024, n14025, n14026, n14027,
    n14028, n14029, n14030, n14031, n14032, n14033,
    n14034, n14035, n14036, n14037, n14038, n14039,
    n14040, n14041, n14042, n14043, n14044, n14045,
    n14046, n14047, n14048, n14049, n14050, n14051,
    n14052, n14053, n14054, n14055, n14056, n14057,
    n14058, n14059, n14060, n14061, n14062, n14063,
    n14064, n14065, n14066, n14067, n14068, n14069,
    n14070, n14071, n14072, n14073, n14074, n14075,
    n14076, n14077, n14078, n14079, n14080, n14081,
    n14082, n14083, n14084, n14085, n14086, n14087,
    n14088, n14089, n14090, n14091, n14092, n14093,
    n14094, n14095, n14096, n14097, n14098, n14099,
    n14100, n14101, n14102, n14103, n14104, n14105,
    n14106, n14107, n14108, n14109, n14110, n14111,
    n14112, n14113, n14114, n14115, n14116, n14117,
    n14118, n14119, n14120, n14121, n14122, n14123,
    n14124, n14125, n14126, n14127, n14128, n14129,
    n14130, n14131, n14132, n14133, n14134, n14135,
    n14136, n14137, n14138, n14139, n14140, n14141,
    n14142, n14143, n14144, n14145, n14146, n14147,
    n14149, n14150, n14151, n14152, n14153, n14154,
    n14155, n14156, n14157, n14158, n14159, n14160,
    n14161, n14162, n14163, n14164, n14165, n14166,
    n14167, n14168, n14169, n14170, n14171, n14172,
    n14173, n14174, n14175, n14176, n14177, n14178,
    n14179, n14180, n14181, n14182, n14183, n14184,
    n14185, n14186, n14187, n14188, n14189, n14190,
    n14191, n14192, n14193, n14194, n14195, n14196,
    n14197, n14198, n14199, n14200, n14201, n14202,
    n14203, n14204, n14205, n14206, n14207, n14208,
    n14209, n14210, n14211, n14212, n14213, n14214,
    n14215, n14216, n14217, n14218, n14219, n14220,
    n14221, n14222, n14223, n14224, n14225, n14226,
    n14227, n14228, n14229, n14230, n14231, n14232,
    n14233, n14234, n14235, n14236, n14237, n14238,
    n14239, n14240, n14241, n14242, n14243, n14244,
    n14245, n14246, n14247, n14248, n14249, n14250,
    n14251, n14252, n14253, n14254, n14255, n14256,
    n14257, n14258, n14259, n14260, n14261, n14262,
    n14263, n14264, n14265, n14266, n14267, n14268,
    n14269, n14270, n14271, n14272, n14273, n14274,
    n14275, n14276, n14277, n14278, n14279, n14280,
    n14281, n14282, n14283, n14284, n14285, n14286,
    n14287, n14288, n14289, n14290, n14291, n14292,
    n14293, n14294, n14295, n14296, n14297, n14298,
    n14299, n14300, n14301, n14302, n14303, n14304,
    n14305, n14306, n14307, n14308, n14309, n14310,
    n14311, n14312, n14313, n14314, n14315, n14316,
    n14317, n14318, n14319, n14320, n14321, n14322,
    n14323, n14324, n14325, n14326, n14327, n14328,
    n14329, n14330, n14331, n14332, n14333, n14334,
    n14335, n14336, n14337, n14338, n14339, n14340,
    n14341, n14342, n14343, n14344, n14345, n14346,
    n14347, n14348, n14349, n14350, n14351, n14352,
    n14353, n14354, n14355, n14356, n14357, n14358,
    n14359, n14360, n14361, n14362, n14363, n14364,
    n14365, n14366, n14367, n14368, n14369, n14370,
    n14371, n14372, n14373, n14374, n14375, n14376,
    n14377, n14378, n14379, n14380, n14381, n14382,
    n14383, n14384, n14385, n14386, n14387, n14388,
    n14389, n14390, n14391, n14392, n14393, n14394,
    n14395, n14396, n14397, n14398, n14399, n14400,
    n14401, n14402, n14403, n14404, n14405, n14406,
    n14407, n14408, n14409, n14410, n14411, n14412,
    n14413, n14414, n14415, n14416, n14417, n14418,
    n14419, n14420, n14421, n14422, n14423, n14424,
    n14425, n14426, n14427, n14428, n14429, n14430,
    n14431, n14432, n14433, n14434, n14435, n14436,
    n14437, n14438, n14439, n14440, n14441, n14442,
    n14443, n14444, n14445, n14446, n14447, n14448,
    n14449, n14450, n14451, n14452, n14453, n14454,
    n14455, n14456, n14457, n14458, n14459, n14460,
    n14461, n14462, n14463, n14464, n14465, n14466,
    n14467, n14468, n14469, n14470, n14471, n14472,
    n14473, n14474, n14475, n14476, n14477, n14478,
    n14479, n14480, n14481, n14482, n14483, n14484,
    n14485, n14486, n14487, n14488, n14489, n14490,
    n14491, n14492, n14493, n14494, n14495, n14496,
    n14497, n14498, n14499, n14500, n14501, n14502,
    n14503, n14504, n14505, n14506, n14507, n14508,
    n14509, n14510, n14511, n14512, n14513, n14514,
    n14515, n14516, n14517, n14518, n14519, n14521,
    n14522, n14523, n14524, n14525, n14526, n14527,
    n14528, n14529, n14530, n14531, n14532, n14533,
    n14534, n14535, n14536, n14537, n14538, n14539,
    n14540, n14541, n14542, n14543, n14544, n14545,
    n14546, n14547, n14548, n14549, n14550, n14551,
    n14552, n14553, n14554, n14555, n14556, n14557,
    n14558, n14559, n14560, n14561, n14562, n14563,
    n14564, n14565, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14573, n14574, n14575,
    n14576, n14577, n14578, n14579, n14580, n14581,
    n14582, n14583, n14584, n14585, n14586, n14587,
    n14588, n14589, n14590, n14591, n14592, n14593,
    n14594, n14595, n14596, n14597, n14598, n14599,
    n14600, n14601, n14602, n14603, n14604, n14605,
    n14606, n14607, n14608, n14609, n14610, n14611,
    n14612, n14613, n14614, n14615, n14616, n14617,
    n14618, n14619, n14620, n14621, n14622, n14623,
    n14624, n14625, n14626, n14627, n14628, n14629,
    n14630, n14631, n14632, n14633, n14634, n14635,
    n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647,
    n14648, n14649, n14650, n14651, n14652, n14653,
    n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665,
    n14666, n14667, n14668, n14669, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683,
    n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701,
    n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719,
    n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731,
    n14732, n14733, n14734, n14735, n14736, n14737,
    n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749,
    n14750, n14751, n14752, n14753, n14754, n14755,
    n14756, n14757, n14758, n14759, n14760, n14761,
    n14762, n14763, n14764, n14765, n14766, n14767,
    n14768, n14769, n14770, n14771, n14772, n14773,
    n14774, n14775, n14776, n14777, n14778, n14779,
    n14780, n14781, n14782, n14783, n14784, n14785,
    n14786, n14787, n14788, n14789, n14790, n14791,
    n14792, n14793, n14794, n14795, n14796, n14797,
    n14798, n14799, n14800, n14801, n14802, n14803,
    n14804, n14805, n14806, n14807, n14808, n14809,
    n14810, n14811, n14812, n14813, n14814, n14815,
    n14816, n14817, n14818, n14819, n14820, n14821,
    n14822, n14823, n14824, n14825, n14826, n14827,
    n14828, n14829, n14830, n14831, n14832, n14833,
    n14834, n14835, n14836, n14837, n14838, n14839,
    n14840, n14841, n14842, n14843, n14844, n14845,
    n14846, n14847, n14848, n14849, n14850, n14851,
    n14852, n14853, n14854, n14855, n14856, n14857,
    n14858, n14859, n14860, n14861, n14862, n14863,
    n14864, n14865, n14866, n14867, n14868, n14869,
    n14870, n14871, n14872, n14873, n14874, n14875,
    n14876, n14877, n14878, n14879, n14880, n14881,
    n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906,
    n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924,
    n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942,
    n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978,
    n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996,
    n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014,
    n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032,
    n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050,
    n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068,
    n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086,
    n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122,
    n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194,
    n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230,
    n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248,
    n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15258, n15259, n15260, n15261,
    n15262, n15263, n15264, n15265, n15266, n15267,
    n15268, n15269, n15270, n15271, n15272, n15273,
    n15274, n15275, n15276, n15277, n15278, n15279,
    n15280, n15281, n15282, n15283, n15284, n15285,
    n15286, n15287, n15288, n15289, n15290, n15291,
    n15292, n15293, n15294, n15295, n15296, n15297,
    n15298, n15299, n15300, n15301, n15302, n15303,
    n15304, n15305, n15306, n15307, n15308, n15309,
    n15310, n15311, n15312, n15313, n15314, n15315,
    n15316, n15317, n15318, n15319, n15320, n15321,
    n15322, n15323, n15324, n15325, n15326, n15327,
    n15328, n15329, n15330, n15331, n15332, n15333,
    n15334, n15335, n15336, n15337, n15338, n15339,
    n15340, n15341, n15342, n15343, n15344, n15345,
    n15346, n15347, n15348, n15349, n15350, n15351,
    n15352, n15353, n15354, n15355, n15356, n15357,
    n15358, n15359, n15360, n15361, n15362, n15363,
    n15364, n15365, n15366, n15367, n15368, n15369,
    n15370, n15371, n15372, n15373, n15374, n15375,
    n15376, n15377, n15378, n15379, n15380, n15381,
    n15382, n15383, n15384, n15385, n15386, n15387,
    n15388, n15389, n15390, n15391, n15392, n15393,
    n15394, n15395, n15396, n15397, n15398, n15399,
    n15400, n15401, n15402, n15403, n15404, n15405,
    n15406, n15407, n15408, n15409, n15410, n15411,
    n15412, n15413, n15414, n15415, n15416, n15417,
    n15418, n15419, n15420, n15421, n15422, n15423,
    n15424, n15425, n15426, n15427, n15428, n15429,
    n15430, n15431, n15432, n15433, n15434, n15435,
    n15436, n15437, n15438, n15439, n15440, n15441,
    n15442, n15443, n15444, n15445, n15446, n15447,
    n15448, n15449, n15450, n15451, n15452, n15453,
    n15454, n15455, n15456, n15457, n15458, n15459,
    n15460, n15461, n15462, n15463, n15464, n15465,
    n15466, n15467, n15468, n15469, n15470, n15471,
    n15472, n15473, n15474, n15475, n15476, n15477,
    n15478, n15479, n15480, n15481, n15482, n15483,
    n15484, n15485, n15486, n15487, n15488, n15489,
    n15490, n15491, n15492, n15493, n15494, n15495,
    n15496, n15497, n15498, n15499, n15500, n15501,
    n15502, n15503, n15504, n15505, n15506, n15507,
    n15508, n15509, n15510, n15511, n15512, n15513,
    n15514, n15515, n15516, n15517, n15518, n15519,
    n15520, n15521, n15522, n15523, n15524, n15525,
    n15526, n15527, n15528, n15529, n15530, n15531,
    n15532, n15533, n15534, n15535, n15536, n15537,
    n15538, n15539, n15540, n15541, n15542, n15543,
    n15544, n15545, n15546, n15547, n15548, n15549,
    n15550, n15551, n15552, n15553, n15554, n15555,
    n15556, n15557, n15558, n15559, n15560, n15561,
    n15562, n15563, n15564, n15565, n15566, n15567,
    n15568, n15569, n15570, n15571, n15572, n15573,
    n15574, n15575, n15576, n15577, n15578, n15579,
    n15580, n15581, n15582, n15583, n15584, n15585,
    n15586, n15587, n15588, n15589, n15590, n15591,
    n15592, n15593, n15594, n15595, n15596, n15597,
    n15598, n15599, n15600, n15601, n15602, n15603,
    n15604, n15605, n15606, n15607, n15608, n15609,
    n15610, n15611, n15612, n15613, n15614, n15615,
    n15616, n15617, n15618, n15619, n15621, n15622,
    n15623, n15624, n15625, n15626, n15627, n15628,
    n15629, n15630, n15631, n15632, n15633, n15634,
    n15635, n15636, n15637, n15638, n15639, n15640,
    n15641, n15642, n15643, n15644, n15645, n15646,
    n15647, n15648, n15649, n15650, n15651, n15652,
    n15653, n15654, n15655, n15656, n15657, n15658,
    n15659, n15660, n15661, n15662, n15663, n15664,
    n15665, n15666, n15667, n15668, n15669, n15670,
    n15671, n15672, n15673, n15674, n15675, n15676,
    n15677, n15678, n15679, n15680, n15681, n15682,
    n15683, n15684, n15685, n15686, n15687, n15688,
    n15689, n15690, n15691, n15692, n15693, n15694,
    n15695, n15696, n15697, n15698, n15699, n15700,
    n15701, n15702, n15703, n15704, n15705, n15706,
    n15707, n15708, n15709, n15710, n15711, n15712,
    n15713, n15714, n15715, n15716, n15717, n15718,
    n15719, n15720, n15721, n15722, n15723, n15724,
    n15725, n15726, n15727, n15728, n15729, n15730,
    n15731, n15732, n15733, n15734, n15735, n15736,
    n15737, n15738, n15739, n15740, n15741, n15742,
    n15743, n15744, n15745, n15746, n15747, n15748,
    n15749, n15750, n15751, n15752, n15753, n15754,
    n15755, n15756, n15757, n15758, n15759, n15760,
    n15761, n15762, n15763, n15764, n15765, n15766,
    n15767, n15768, n15769, n15770, n15771, n15772,
    n15773, n15774, n15775, n15776, n15777, n15778,
    n15779, n15780, n15781, n15782, n15783, n15784,
    n15785, n15786, n15787, n15788, n15789, n15790,
    n15791, n15792, n15793, n15794, n15795, n15796,
    n15797, n15798, n15799, n15800, n15801, n15802,
    n15803, n15804, n15805, n15806, n15807, n15808,
    n15809, n15810, n15811, n15812, n15813, n15814,
    n15815, n15816, n15817, n15818, n15819, n15820,
    n15821, n15822, n15823, n15824, n15825, n15826,
    n15827, n15828, n15829, n15830, n15831, n15832,
    n15833, n15834, n15835, n15836, n15837, n15838,
    n15839, n15840, n15841, n15842, n15843, n15844,
    n15845, n15846, n15847, n15848, n15849, n15850,
    n15851, n15852, n15853, n15854, n15855, n15856,
    n15857, n15858, n15859, n15860, n15861, n15862,
    n15863, n15864, n15865, n15866, n15867, n15868,
    n15869, n15870, n15871, n15872, n15873, n15874,
    n15875, n15876, n15877, n15878, n15879, n15880,
    n15881, n15882, n15883, n15884, n15885, n15886,
    n15887, n15888, n15889, n15890, n15891, n15892,
    n15893, n15894, n15895, n15896, n15897, n15898,
    n15899, n15900, n15901, n15902, n15903, n15904,
    n15905, n15906, n15907, n15908, n15909, n15910,
    n15911, n15912, n15913, n15914, n15915, n15916,
    n15917, n15918, n15919, n15920, n15921, n15922,
    n15923, n15924, n15925, n15926, n15927, n15928,
    n15929, n15930, n15931, n15932, n15933, n15934,
    n15935, n15936, n15937, n15938, n15939, n15940,
    n15941, n15942, n15943, n15944, n15945, n15946,
    n15947, n15948, n15949, n15950, n15951, n15952,
    n15953, n15954, n15955, n15956, n15957, n15958,
    n15959, n15960, n15961, n15962, n15963, n15964,
    n15965, n15966, n15967, n15968, n15969, n15970,
    n15971, n15972, n15973, n15974, n15975, n15977,
    n15978, n15979, n15980, n15981, n15982, n15983,
    n15984, n15985, n15986, n15987, n15988, n15989,
    n15990, n15991, n15992, n15993, n15994, n15995,
    n15996, n15997, n15998, n15999, n16000, n16001,
    n16002, n16003, n16004, n16005, n16006, n16007,
    n16008, n16009, n16010, n16011, n16012, n16013,
    n16014, n16015, n16016, n16017, n16018, n16019,
    n16020, n16021, n16022, n16023, n16024, n16025,
    n16026, n16027, n16028, n16029, n16030, n16031,
    n16032, n16033, n16034, n16035, n16036, n16037,
    n16038, n16039, n16040, n16041, n16042, n16043,
    n16044, n16045, n16046, n16047, n16048, n16049,
    n16050, n16051, n16052, n16053, n16054, n16055,
    n16056, n16057, n16058, n16059, n16060, n16061,
    n16062, n16063, n16064, n16065, n16066, n16067,
    n16068, n16069, n16070, n16071, n16072, n16073,
    n16074, n16075, n16076, n16077, n16078, n16079,
    n16080, n16081, n16082, n16083, n16084, n16085,
    n16086, n16087, n16088, n16089, n16090, n16091,
    n16092, n16093, n16094, n16095, n16096, n16097,
    n16098, n16099, n16100, n16101, n16102, n16103,
    n16104, n16105, n16106, n16107, n16108, n16109,
    n16110, n16111, n16112, n16113, n16114, n16115,
    n16116, n16117, n16118, n16119, n16120, n16121,
    n16122, n16123, n16124, n16125, n16126, n16127,
    n16128, n16129, n16130, n16131, n16132, n16133,
    n16134, n16135, n16136, n16137, n16138, n16139,
    n16140, n16141, n16142, n16143, n16144, n16145,
    n16146, n16147, n16148, n16149, n16150, n16151,
    n16152, n16153, n16154, n16155, n16156, n16157,
    n16158, n16159, n16160, n16161, n16162, n16163,
    n16164, n16165, n16166, n16167, n16168, n16169,
    n16170, n16171, n16172, n16173, n16174, n16175,
    n16176, n16177, n16178, n16179, n16180, n16181,
    n16182, n16183, n16184, n16185, n16186, n16187,
    n16188, n16189, n16190, n16191, n16192, n16193,
    n16194, n16195, n16196, n16197, n16198, n16199,
    n16200, n16201, n16202, n16203, n16204, n16205,
    n16206, n16207, n16208, n16209, n16210, n16211,
    n16212, n16213, n16214, n16215, n16216, n16217,
    n16218, n16219, n16220, n16221, n16222, n16223,
    n16224, n16225, n16226, n16227, n16228, n16229,
    n16230, n16231, n16232, n16233, n16234, n16235,
    n16236, n16237, n16238, n16239, n16240, n16241,
    n16242, n16243, n16244, n16245, n16246, n16247,
    n16248, n16249, n16250, n16251, n16252, n16253,
    n16254, n16255, n16256, n16257, n16258, n16259,
    n16260, n16261, n16262, n16263, n16264, n16265,
    n16266, n16267, n16268, n16269, n16270, n16271,
    n16272, n16273, n16274, n16275, n16276, n16277,
    n16278, n16279, n16280, n16281, n16282, n16283,
    n16284, n16285, n16286, n16287, n16288, n16289,
    n16290, n16291, n16292, n16293, n16294, n16295,
    n16296, n16297, n16298, n16299, n16300, n16301,
    n16302, n16303, n16304, n16305, n16306, n16307,
    n16308, n16309, n16310, n16311, n16312, n16313,
    n16314, n16315, n16316, n16317, n16318, n16319,
    n16320, n16321, n16322, n16323, n16324, n16325,
    n16326, n16327, n16328, n16329, n16330, n16331,
    n16333, n16334, n16335, n16336, n16337, n16338,
    n16339, n16340, n16341, n16342, n16343, n16344,
    n16345, n16346, n16347, n16348, n16349, n16350,
    n16351, n16352, n16353, n16354, n16355, n16356,
    n16357, n16358, n16359, n16360, n16361, n16362,
    n16363, n16364, n16365, n16366, n16367, n16368,
    n16369, n16370, n16371, n16372, n16373, n16374,
    n16375, n16376, n16377, n16378, n16379, n16380,
    n16381, n16382, n16383, n16384, n16385, n16386,
    n16387, n16388, n16389, n16390, n16391, n16392,
    n16393, n16394, n16395, n16396, n16397, n16398,
    n16399, n16400, n16401, n16402, n16403, n16404,
    n16405, n16406, n16407, n16408, n16409, n16410,
    n16411, n16412, n16413, n16414, n16415, n16416,
    n16417, n16418, n16419, n16420, n16421, n16422,
    n16423, n16424, n16425, n16426, n16427, n16428,
    n16429, n16430, n16431, n16432, n16433, n16434,
    n16435, n16436, n16437, n16438, n16439, n16440,
    n16441, n16442, n16443, n16444, n16445, n16446,
    n16447, n16448, n16449, n16450, n16451, n16452,
    n16453, n16454, n16455, n16456, n16457, n16458,
    n16459, n16460, n16461, n16462, n16463, n16464,
    n16465, n16466, n16467, n16468, n16469, n16470,
    n16471, n16472, n16473, n16474, n16475, n16476,
    n16477, n16478, n16479, n16480, n16481, n16482,
    n16483, n16484, n16485, n16486, n16487, n16488,
    n16489, n16490, n16491, n16492, n16493, n16494,
    n16495, n16496, n16497, n16498, n16499, n16500,
    n16501, n16502, n16503, n16504, n16505, n16506,
    n16507, n16508, n16509, n16510, n16511, n16512,
    n16513, n16514, n16515, n16516, n16517, n16518,
    n16519, n16520, n16521, n16522, n16523, n16524,
    n16525, n16526, n16527, n16528, n16529, n16530,
    n16531, n16532, n16533, n16534, n16535, n16536,
    n16537, n16538, n16539, n16540, n16541, n16542,
    n16543, n16544, n16545, n16546, n16547, n16548,
    n16549, n16550, n16551, n16552, n16553, n16554,
    n16555, n16556, n16557, n16558, n16559, n16560,
    n16561, n16562, n16563, n16564, n16565, n16566,
    n16567, n16568, n16569, n16570, n16571, n16572,
    n16573, n16574, n16575, n16576, n16577, n16578,
    n16579, n16580, n16581, n16582, n16583, n16584,
    n16585, n16586, n16587, n16588, n16589, n16590,
    n16591, n16592, n16593, n16594, n16595, n16596,
    n16597, n16598, n16599, n16600, n16601, n16602,
    n16603, n16604, n16605, n16606, n16607, n16608,
    n16609, n16610, n16611, n16612, n16613, n16614,
    n16615, n16616, n16617, n16618, n16619, n16620,
    n16621, n16622, n16623, n16624, n16625, n16626,
    n16627, n16628, n16629, n16630, n16631, n16632,
    n16633, n16634, n16635, n16636, n16637, n16638,
    n16639, n16640, n16641, n16642, n16643, n16644,
    n16645, n16646, n16647, n16648, n16649, n16650,
    n16651, n16652, n16653, n16654, n16655, n16656,
    n16657, n16658, n16659, n16660, n16661, n16662,
    n16663, n16664, n16665, n16666, n16667, n16668,
    n16669, n16670, n16671, n16672, n16673, n16674,
    n16675, n16676, n16677, n16679, n16680, n16681,
    n16682, n16683, n16684, n16685, n16686, n16687,
    n16688, n16689, n16690, n16691, n16692, n16693,
    n16694, n16695, n16696, n16697, n16698, n16699,
    n16700, n16701, n16702, n16703, n16704, n16705,
    n16706, n16707, n16708, n16709, n16710, n16711,
    n16712, n16713, n16714, n16715, n16716, n16717,
    n16718, n16719, n16720, n16721, n16722, n16723,
    n16724, n16725, n16726, n16727, n16728, n16729,
    n16730, n16731, n16732, n16733, n16734, n16735,
    n16736, n16737, n16738, n16739, n16740, n16741,
    n16742, n16743, n16744, n16745, n16746, n16747,
    n16748, n16749, n16750, n16751, n16752, n16753,
    n16754, n16755, n16756, n16757, n16758, n16759,
    n16760, n16761, n16762, n16763, n16764, n16765,
    n16766, n16767, n16768, n16769, n16770, n16771,
    n16772, n16773, n16774, n16775, n16776, n16777,
    n16778, n16779, n16780, n16781, n16782, n16783,
    n16784, n16785, n16786, n16787, n16788, n16789,
    n16790, n16791, n16792, n16793, n16794, n16795,
    n16796, n16797, n16798, n16799, n16800, n16801,
    n16802, n16803, n16804, n16805, n16806, n16807,
    n16808, n16809, n16810, n16811, n16812, n16813,
    n16814, n16815, n16816, n16817, n16818, n16819,
    n16820, n16821, n16822, n16823, n16824, n16825,
    n16826, n16827, n16828, n16829, n16830, n16831,
    n16832, n16833, n16834, n16835, n16836, n16837,
    n16838, n16839, n16840, n16841, n16842, n16843,
    n16844, n16845, n16846, n16847, n16848, n16849,
    n16850, n16851, n16852, n16853, n16854, n16855,
    n16856, n16857, n16858, n16859, n16860, n16861,
    n16862, n16863, n16864, n16865, n16866, n16867,
    n16868, n16869, n16870, n16871, n16872, n16873,
    n16874, n16875, n16876, n16877, n16878, n16879,
    n16880, n16881, n16882, n16883, n16884, n16885,
    n16886, n16887, n16888, n16889, n16890, n16891,
    n16892, n16893, n16894, n16895, n16896, n16897,
    n16898, n16899, n16900, n16901, n16902, n16903,
    n16904, n16905, n16906, n16907, n16908, n16909,
    n16910, n16911, n16912, n16913, n16914, n16915,
    n16916, n16917, n16918, n16919, n16920, n16921,
    n16922, n16923, n16924, n16925, n16926, n16927,
    n16928, n16929, n16930, n16931, n16932, n16933,
    n16934, n16935, n16936, n16937, n16938, n16939,
    n16940, n16941, n16942, n16943, n16944, n16945,
    n16946, n16947, n16948, n16949, n16950, n16951,
    n16952, n16953, n16954, n16955, n16956, n16957,
    n16958, n16959, n16960, n16961, n16962, n16963,
    n16964, n16965, n16966, n16967, n16968, n16969,
    n16970, n16971, n16972, n16973, n16974, n16975,
    n16976, n16977, n16978, n16979, n16980, n16981,
    n16982, n16983, n16984, n16985, n16986, n16987,
    n16988, n16989, n16990, n16991, n16992, n16993,
    n16994, n16995, n16996, n16997, n16998, n16999,
    n17000, n17001, n17002, n17003, n17004, n17005,
    n17006, n17007, n17008, n17009, n17010, n17011,
    n17012, n17013, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024,
    n17025, n17026, n17027, n17028, n17029, n17030,
    n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042,
    n17043, n17044, n17045, n17046, n17047, n17048,
    n17049, n17050, n17051, n17052, n17053, n17054,
    n17055, n17056, n17057, n17058, n17059, n17060,
    n17061, n17062, n17063, n17064, n17065, n17066,
    n17067, n17068, n17069, n17070, n17071, n17072,
    n17073, n17074, n17075, n17076, n17077, n17078,
    n17079, n17080, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090,
    n17091, n17092, n17093, n17094, n17095, n17096,
    n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17114,
    n17115, n17116, n17117, n17118, n17119, n17120,
    n17121, n17122, n17123, n17124, n17125, n17126,
    n17127, n17128, n17129, n17130, n17131, n17132,
    n17133, n17134, n17135, n17136, n17137, n17138,
    n17139, n17140, n17141, n17142, n17143, n17144,
    n17145, n17146, n17147, n17148, n17149, n17150,
    n17151, n17152, n17153, n17154, n17155, n17156,
    n17157, n17158, n17159, n17160, n17161, n17162,
    n17163, n17164, n17165, n17166, n17167, n17168,
    n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180,
    n17181, n17182, n17183, n17184, n17185, n17186,
    n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204,
    n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222,
    n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240,
    n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258,
    n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276,
    n17277, n17278, n17279, n17280, n17281, n17282,
    n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294,
    n17295, n17296, n17297, n17298, n17299, n17300,
    n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312,
    n17313, n17314, n17315, n17316, n17317, n17318,
    n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330,
    n17331, n17332, n17333, n17334, n17335, n17336,
    n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348,
    n17349, n17351, n17352, n17353, n17354, n17355,
    n17356, n17357, n17358, n17359, n17360, n17361,
    n17362, n17363, n17364, n17365, n17366, n17367,
    n17368, n17369, n17370, n17371, n17372, n17373,
    n17374, n17375, n17376, n17377, n17378, n17379,
    n17380, n17381, n17382, n17383, n17384, n17385,
    n17386, n17387, n17388, n17389, n17390, n17391,
    n17392, n17393, n17394, n17395, n17396, n17397,
    n17398, n17399, n17400, n17401, n17402, n17403,
    n17404, n17405, n17406, n17407, n17408, n17409,
    n17410, n17411, n17412, n17413, n17414, n17415,
    n17416, n17417, n17418, n17419, n17420, n17421,
    n17422, n17423, n17424, n17425, n17426, n17427,
    n17428, n17429, n17430, n17431, n17432, n17433,
    n17434, n17435, n17436, n17437, n17438, n17439,
    n17440, n17441, n17442, n17443, n17444, n17445,
    n17446, n17447, n17448, n17449, n17450, n17451,
    n17452, n17453, n17454, n17455, n17456, n17457,
    n17458, n17459, n17460, n17461, n17462, n17463,
    n17464, n17465, n17466, n17467, n17468, n17469,
    n17470, n17471, n17472, n17473, n17474, n17475,
    n17476, n17477, n17478, n17479, n17480, n17481,
    n17482, n17483, n17484, n17485, n17486, n17487,
    n17488, n17489, n17490, n17491, n17492, n17493,
    n17494, n17495, n17496, n17497, n17498, n17499,
    n17500, n17501, n17502, n17503, n17504, n17505,
    n17506, n17507, n17508, n17509, n17510, n17511,
    n17512, n17513, n17514, n17515, n17516, n17517,
    n17518, n17519, n17520, n17521, n17522, n17523,
    n17524, n17525, n17526, n17527, n17528, n17529,
    n17530, n17531, n17532, n17533, n17534, n17535,
    n17536, n17537, n17538, n17539, n17540, n17541,
    n17542, n17543, n17544, n17545, n17546, n17547,
    n17548, n17549, n17550, n17551, n17552, n17553,
    n17554, n17555, n17556, n17557, n17558, n17559,
    n17560, n17561, n17562, n17563, n17564, n17565,
    n17566, n17567, n17568, n17569, n17570, n17571,
    n17572, n17573, n17574, n17575, n17576, n17577,
    n17578, n17579, n17580, n17581, n17582, n17583,
    n17584, n17585, n17586, n17587, n17588, n17589,
    n17590, n17591, n17592, n17593, n17594, n17595,
    n17596, n17597, n17598, n17599, n17600, n17601,
    n17602, n17603, n17604, n17605, n17606, n17607,
    n17608, n17609, n17610, n17611, n17612, n17613,
    n17614, n17615, n17616, n17617, n17618, n17619,
    n17620, n17621, n17622, n17623, n17624, n17625,
    n17626, n17627, n17628, n17629, n17630, n17631,
    n17632, n17633, n17634, n17635, n17636, n17637,
    n17638, n17639, n17640, n17641, n17642, n17643,
    n17644, n17645, n17646, n17647, n17648, n17649,
    n17650, n17651, n17652, n17653, n17654, n17655,
    n17656, n17657, n17658, n17659, n17660, n17661,
    n17662, n17663, n17664, n17665, n17666, n17667,
    n17668, n17669, n17670, n17671, n17672, n17673,
    n17674, n17675, n17676, n17677, n17678, n17679,
    n17680, n17681, n17682, n17683, n17684, n17686,
    n17687, n17688, n17689, n17690, n17691, n17692,
    n17693, n17694, n17695, n17696, n17697, n17698,
    n17699, n17700, n17701, n17702, n17703, n17704,
    n17705, n17706, n17707, n17708, n17709, n17710,
    n17711, n17712, n17713, n17714, n17715, n17716,
    n17717, n17718, n17719, n17720, n17721, n17722,
    n17723, n17724, n17725, n17726, n17727, n17728,
    n17729, n17730, n17731, n17732, n17733, n17734,
    n17735, n17736, n17737, n17738, n17739, n17740,
    n17741, n17742, n17743, n17744, n17745, n17746,
    n17747, n17748, n17749, n17750, n17751, n17752,
    n17753, n17754, n17755, n17756, n17757, n17758,
    n17759, n17760, n17761, n17762, n17763, n17764,
    n17765, n17766, n17767, n17768, n17769, n17770,
    n17771, n17772, n17773, n17774, n17775, n17776,
    n17777, n17778, n17779, n17780, n17781, n17782,
    n17783, n17784, n17785, n17786, n17787, n17788,
    n17789, n17790, n17791, n17792, n17793, n17794,
    n17795, n17796, n17797, n17798, n17799, n17800,
    n17801, n17802, n17803, n17804, n17805, n17806,
    n17807, n17808, n17809, n17810, n17811, n17812,
    n17813, n17814, n17815, n17816, n17817, n17818,
    n17819, n17820, n17821, n17822, n17823, n17824,
    n17825, n17826, n17827, n17828, n17829, n17830,
    n17831, n17832, n17833, n17834, n17835, n17836,
    n17837, n17838, n17839, n17840, n17841, n17842,
    n17843, n17844, n17845, n17846, n17847, n17848,
    n17849, n17850, n17851, n17852, n17853, n17854,
    n17855, n17856, n17857, n17858, n17859, n17860,
    n17861, n17862, n17863, n17864, n17865, n17866,
    n17867, n17868, n17869, n17870, n17871, n17872,
    n17873, n17874, n17875, n17876, n17877, n17878,
    n17879, n17880, n17881, n17882, n17883, n17884,
    n17885, n17886, n17887, n17888, n17889, n17890,
    n17891, n17892, n17893, n17894, n17895, n17896,
    n17897, n17898, n17899, n17900, n17901, n17902,
    n17903, n17904, n17905, n17906, n17907, n17908,
    n17909, n17910, n17911, n17912, n17913, n17914,
    n17915, n17916, n17917, n17918, n17919, n17920,
    n17921, n17922, n17923, n17924, n17925, n17926,
    n17927, n17928, n17929, n17930, n17931, n17932,
    n17933, n17934, n17935, n17936, n17937, n17938,
    n17939, n17940, n17941, n17942, n17943, n17944,
    n17945, n17946, n17947, n17948, n17949, n17950,
    n17951, n17952, n17953, n17954, n17955, n17956,
    n17957, n17958, n17959, n17960, n17961, n17962,
    n17963, n17964, n17965, n17966, n17967, n17968,
    n17969, n17970, n17971, n17972, n17973, n17974,
    n17975, n17976, n17977, n17978, n17979, n17980,
    n17981, n17982, n17983, n17984, n17985, n17986,
    n17987, n17988, n17989, n17990, n17991, n17992,
    n17993, n17994, n17995, n17996, n17997, n17998,
    n17999, n18000, n18002, n18003, n18004, n18005,
    n18006, n18007, n18008, n18009, n18010, n18011,
    n18012, n18013, n18014, n18015, n18016, n18017,
    n18018, n18019, n18020, n18021, n18022, n18023,
    n18024, n18025, n18026, n18027, n18028, n18029,
    n18030, n18031, n18032, n18033, n18034, n18035,
    n18036, n18037, n18038, n18039, n18040, n18041,
    n18042, n18043, n18044, n18045, n18046, n18047,
    n18048, n18049, n18050, n18051, n18052, n18053,
    n18054, n18055, n18056, n18057, n18058, n18059,
    n18060, n18061, n18062, n18063, n18064, n18065,
    n18066, n18067, n18068, n18069, n18070, n18071,
    n18072, n18073, n18074, n18075, n18076, n18077,
    n18078, n18079, n18080, n18081, n18082, n18083,
    n18084, n18085, n18086, n18087, n18088, n18089,
    n18090, n18091, n18092, n18093, n18094, n18095,
    n18096, n18097, n18098, n18099, n18100, n18101,
    n18102, n18103, n18104, n18105, n18106, n18107,
    n18108, n18109, n18110, n18111, n18112, n18113,
    n18114, n18115, n18116, n18117, n18118, n18119,
    n18120, n18121, n18122, n18123, n18124, n18125,
    n18126, n18127, n18128, n18129, n18130, n18131,
    n18132, n18133, n18134, n18135, n18136, n18137,
    n18138, n18139, n18140, n18141, n18142, n18143,
    n18144, n18145, n18146, n18147, n18148, n18149,
    n18150, n18151, n18152, n18153, n18154, n18155,
    n18156, n18157, n18158, n18159, n18160, n18161,
    n18162, n18163, n18164, n18165, n18166, n18167,
    n18168, n18169, n18170, n18171, n18172, n18173,
    n18174, n18175, n18176, n18177, n18178, n18179,
    n18180, n18181, n18182, n18183, n18184, n18185,
    n18186, n18187, n18188, n18189, n18190, n18191,
    n18192, n18193, n18194, n18195, n18196, n18197,
    n18198, n18199, n18200, n18201, n18202, n18203,
    n18204, n18205, n18206, n18207, n18208, n18209,
    n18210, n18211, n18212, n18213, n18214, n18215,
    n18216, n18217, n18218, n18219, n18220, n18221,
    n18222, n18223, n18224, n18225, n18226, n18227,
    n18228, n18229, n18230, n18231, n18232, n18233,
    n18234, n18235, n18236, n18237, n18238, n18239,
    n18240, n18241, n18242, n18243, n18244, n18245,
    n18246, n18247, n18248, n18249, n18250, n18251,
    n18252, n18253, n18254, n18255, n18256, n18257,
    n18258, n18259, n18260, n18261, n18262, n18263,
    n18264, n18265, n18266, n18267, n18268, n18269,
    n18270, n18271, n18272, n18273, n18274, n18275,
    n18276, n18277, n18278, n18279, n18280, n18281,
    n18282, n18283, n18284, n18285, n18286, n18287,
    n18288, n18289, n18290, n18291, n18292, n18293,
    n18294, n18295, n18296, n18297, n18298, n18299,
    n18300, n18301, n18302, n18303, n18304, n18305,
    n18306, n18307, n18308, n18309, n18310, n18311,
    n18312, n18313, n18314, n18315, n18316, n18317,
    n18318, n18320, n18321, n18322, n18323, n18324,
    n18325, n18326, n18327, n18328, n18329, n18330,
    n18331, n18332, n18333, n18334, n18335, n18336,
    n18337, n18338, n18339, n18340, n18341, n18342,
    n18343, n18344, n18345, n18346, n18347, n18348,
    n18349, n18350, n18351, n18352, n18353, n18354,
    n18355, n18356, n18357, n18358, n18359, n18360,
    n18361, n18362, n18363, n18364, n18365, n18366,
    n18367, n18368, n18369, n18370, n18371, n18372,
    n18373, n18374, n18375, n18376, n18377, n18378,
    n18379, n18380, n18381, n18382, n18383, n18384,
    n18385, n18386, n18387, n18388, n18389, n18390,
    n18391, n18392, n18393, n18394, n18395, n18396,
    n18397, n18398, n18399, n18400, n18401, n18402,
    n18403, n18404, n18405, n18406, n18407, n18408,
    n18409, n18410, n18411, n18412, n18413, n18414,
    n18415, n18416, n18417, n18418, n18419, n18420,
    n18421, n18422, n18423, n18424, n18425, n18426,
    n18427, n18428, n18429, n18430, n18431, n18432,
    n18433, n18434, n18435, n18436, n18437, n18438,
    n18439, n18440, n18441, n18442, n18443, n18444,
    n18445, n18446, n18447, n18448, n18449, n18450,
    n18451, n18452, n18453, n18454, n18455, n18456,
    n18457, n18458, n18459, n18460, n18461, n18462,
    n18463, n18464, n18465, n18466, n18467, n18468,
    n18469, n18470, n18471, n18472, n18473, n18474,
    n18475, n18476, n18477, n18478, n18479, n18480,
    n18481, n18482, n18483, n18484, n18485, n18486,
    n18487, n18488, n18489, n18490, n18491, n18492,
    n18493, n18494, n18495, n18496, n18497, n18498,
    n18499, n18500, n18501, n18502, n18503, n18504,
    n18505, n18506, n18507, n18508, n18509, n18510,
    n18511, n18512, n18513, n18514, n18515, n18516,
    n18517, n18518, n18519, n18520, n18521, n18522,
    n18523, n18524, n18525, n18526, n18527, n18528,
    n18529, n18530, n18531, n18532, n18533, n18534,
    n18535, n18536, n18537, n18538, n18539, n18540,
    n18541, n18542, n18543, n18544, n18545, n18546,
    n18547, n18548, n18549, n18550, n18551, n18552,
    n18553, n18554, n18555, n18556, n18557, n18558,
    n18559, n18560, n18561, n18562, n18563, n18564,
    n18565, n18566, n18567, n18568, n18569, n18570,
    n18571, n18572, n18573, n18574, n18575, n18576,
    n18577, n18578, n18579, n18580, n18581, n18582,
    n18583, n18584, n18585, n18586, n18587, n18588,
    n18589, n18590, n18591, n18592, n18593, n18594,
    n18595, n18596, n18597, n18598, n18599, n18600,
    n18601, n18602, n18603, n18604, n18605, n18606,
    n18607, n18608, n18609, n18610, n18611, n18612,
    n18613, n18614, n18615, n18616, n18617, n18618,
    n18619, n18620, n18621, n18622, n18623, n18624,
    n18625, n18626, n18627, n18628, n18629, n18630,
    n18631, n18632, n18633, n18635, n18636, n18637,
    n18638, n18639, n18640, n18641, n18642, n18643,
    n18644, n18645, n18646, n18647, n18648, n18649,
    n18650, n18651, n18652, n18653, n18654, n18655,
    n18656, n18657, n18658, n18659, n18660, n18661,
    n18662, n18663, n18664, n18665, n18666, n18667,
    n18668, n18669, n18670, n18671, n18672, n18673,
    n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685,
    n18686, n18687, n18688, n18689, n18690, n18691,
    n18692, n18693, n18694, n18695, n18696, n18697,
    n18698, n18699, n18700, n18701, n18702, n18703,
    n18704, n18705, n18706, n18707, n18708, n18709,
    n18710, n18711, n18712, n18713, n18714, n18715,
    n18716, n18717, n18718, n18719, n18720, n18721,
    n18722, n18723, n18724, n18725, n18726, n18727,
    n18728, n18729, n18730, n18731, n18732, n18733,
    n18734, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18742, n18743, n18744, n18745,
    n18746, n18747, n18748, n18749, n18750, n18751,
    n18752, n18753, n18754, n18755, n18756, n18757,
    n18758, n18759, n18760, n18761, n18762, n18763,
    n18764, n18765, n18766, n18767, n18768, n18769,
    n18770, n18771, n18772, n18773, n18774, n18775,
    n18776, n18777, n18778, n18779, n18780, n18781,
    n18782, n18783, n18784, n18785, n18786, n18787,
    n18788, n18789, n18790, n18791, n18792, n18793,
    n18794, n18795, n18796, n18797, n18798, n18799,
    n18800, n18801, n18802, n18803, n18804, n18805,
    n18806, n18807, n18808, n18809, n18810, n18811,
    n18812, n18813, n18814, n18815, n18816, n18817,
    n18818, n18819, n18820, n18821, n18822, n18823,
    n18824, n18825, n18826, n18827, n18828, n18829,
    n18830, n18831, n18832, n18833, n18834, n18835,
    n18836, n18837, n18838, n18839, n18840, n18841,
    n18842, n18843, n18844, n18845, n18846, n18847,
    n18848, n18849, n18850, n18851, n18852, n18853,
    n18854, n18855, n18856, n18857, n18858, n18859,
    n18860, n18861, n18862, n18863, n18864, n18865,
    n18866, n18867, n18868, n18869, n18870, n18871,
    n18872, n18873, n18874, n18875, n18876, n18877,
    n18878, n18879, n18880, n18881, n18882, n18883,
    n18884, n18885, n18886, n18887, n18888, n18889,
    n18890, n18891, n18892, n18893, n18894, n18895,
    n18896, n18897, n18898, n18899, n18900, n18901,
    n18902, n18903, n18904, n18905, n18906, n18907,
    n18908, n18909, n18910, n18911, n18912, n18913,
    n18914, n18915, n18916, n18917, n18918, n18919,
    n18920, n18921, n18922, n18923, n18924, n18925,
    n18926, n18927, n18928, n18929, n18930, n18931,
    n18932, n18933, n18934, n18935, n18936, n18938,
    n18939, n18940, n18941, n18942, n18943, n18944,
    n18945, n18946, n18947, n18948, n18949, n18950,
    n18951, n18952, n18953, n18954, n18955, n18956,
    n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968,
    n18969, n18970, n18971, n18972, n18973, n18974,
    n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986,
    n18987, n18988, n18989, n18990, n18991, n18992,
    n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004,
    n19005, n19006, n19007, n19008, n19009, n19010,
    n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022,
    n19023, n19024, n19025, n19026, n19027, n19028,
    n19029, n19030, n19031, n19032, n19033, n19034,
    n19035, n19036, n19037, n19038, n19039, n19040,
    n19041, n19042, n19043, n19044, n19045, n19046,
    n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058,
    n19059, n19060, n19061, n19062, n19063, n19064,
    n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076,
    n19077, n19078, n19079, n19080, n19081, n19082,
    n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094,
    n19095, n19096, n19097, n19098, n19099, n19100,
    n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112,
    n19113, n19114, n19115, n19116, n19117, n19118,
    n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130,
    n19131, n19132, n19133, n19134, n19135, n19136,
    n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148,
    n19149, n19150, n19151, n19152, n19153, n19154,
    n19155, n19156, n19157, n19158, n19159, n19160,
    n19161, n19162, n19163, n19164, n19165, n19166,
    n19167, n19168, n19169, n19170, n19171, n19172,
    n19173, n19174, n19175, n19176, n19177, n19178,
    n19179, n19180, n19181, n19182, n19183, n19184,
    n19185, n19186, n19187, n19188, n19189, n19190,
    n19191, n19192, n19193, n19194, n19195, n19196,
    n19197, n19198, n19199, n19200, n19201, n19202,
    n19203, n19204, n19205, n19206, n19207, n19208,
    n19209, n19210, n19211, n19212, n19213, n19214,
    n19215, n19216, n19217, n19218, n19219, n19220,
    n19221, n19222, n19223, n19224, n19225, n19226,
    n19227, n19228, n19229, n19230, n19231, n19232,
    n19233, n19234, n19235, n19236, n19237, n19239,
    n19240, n19241, n19242, n19243, n19244, n19245,
    n19246, n19247, n19248, n19249, n19250, n19251,
    n19252, n19253, n19254, n19255, n19256, n19257,
    n19258, n19259, n19260, n19261, n19262, n19263,
    n19264, n19265, n19266, n19267, n19268, n19269,
    n19270, n19271, n19272, n19273, n19274, n19275,
    n19276, n19277, n19278, n19279, n19280, n19281,
    n19282, n19283, n19284, n19285, n19286, n19287,
    n19288, n19289, n19290, n19291, n19292, n19293,
    n19294, n19295, n19296, n19297, n19298, n19299,
    n19300, n19301, n19302, n19303, n19304, n19305,
    n19306, n19307, n19308, n19309, n19310, n19311,
    n19312, n19313, n19314, n19315, n19316, n19317,
    n19318, n19319, n19320, n19321, n19322, n19323,
    n19324, n19325, n19326, n19327, n19328, n19329,
    n19330, n19331, n19332, n19333, n19334, n19335,
    n19336, n19337, n19338, n19339, n19340, n19341,
    n19342, n19343, n19344, n19345, n19346, n19347,
    n19348, n19349, n19350, n19351, n19352, n19353,
    n19354, n19355, n19356, n19357, n19358, n19359,
    n19360, n19361, n19362, n19363, n19364, n19365,
    n19366, n19367, n19368, n19369, n19370, n19371,
    n19372, n19373, n19374, n19375, n19376, n19377,
    n19378, n19379, n19380, n19381, n19382, n19383,
    n19384, n19385, n19386, n19387, n19388, n19389,
    n19390, n19391, n19392, n19393, n19394, n19395,
    n19396, n19397, n19398, n19399, n19400, n19401,
    n19402, n19403, n19404, n19405, n19406, n19407,
    n19408, n19409, n19410, n19411, n19412, n19413,
    n19414, n19415, n19416, n19417, n19418, n19419,
    n19420, n19421, n19422, n19423, n19424, n19425,
    n19426, n19427, n19428, n19429, n19430, n19431,
    n19432, n19433, n19434, n19435, n19436, n19437,
    n19438, n19439, n19440, n19441, n19442, n19443,
    n19444, n19445, n19446, n19447, n19448, n19449,
    n19450, n19451, n19452, n19453, n19454, n19455,
    n19456, n19457, n19458, n19459, n19460, n19461,
    n19462, n19463, n19464, n19465, n19466, n19467,
    n19468, n19469, n19470, n19471, n19472, n19473,
    n19474, n19475, n19476, n19477, n19478, n19479,
    n19480, n19481, n19482, n19483, n19484, n19485,
    n19486, n19487, n19488, n19489, n19490, n19491,
    n19492, n19493, n19494, n19495, n19496, n19497,
    n19498, n19499, n19500, n19501, n19502, n19503,
    n19504, n19505, n19506, n19507, n19508, n19509,
    n19510, n19511, n19512, n19513, n19514, n19515,
    n19516, n19517, n19518, n19519, n19520, n19521,
    n19522, n19523, n19524, n19525, n19527, n19528,
    n19529, n19530, n19531, n19532, n19533, n19534,
    n19535, n19536, n19537, n19538, n19539, n19540,
    n19541, n19542, n19543, n19544, n19545, n19546,
    n19547, n19548, n19549, n19550, n19551, n19552,
    n19553, n19554, n19555, n19556, n19557, n19558,
    n19559, n19560, n19561, n19562, n19563, n19564,
    n19565, n19566, n19567, n19568, n19569, n19570,
    n19571, n19572, n19573, n19574, n19575, n19576,
    n19577, n19578, n19579, n19580, n19581, n19582,
    n19583, n19584, n19585, n19586, n19587, n19588,
    n19589, n19590, n19591, n19592, n19593, n19594,
    n19595, n19596, n19597, n19598, n19599, n19600,
    n19601, n19602, n19603, n19604, n19605, n19606,
    n19607, n19608, n19609, n19610, n19611, n19612,
    n19613, n19614, n19615, n19616, n19617, n19618,
    n19619, n19620, n19621, n19622, n19623, n19624,
    n19625, n19626, n19627, n19628, n19629, n19630,
    n19631, n19632, n19633, n19634, n19635, n19636,
    n19637, n19638, n19639, n19640, n19641, n19642,
    n19643, n19644, n19645, n19646, n19647, n19648,
    n19649, n19650, n19651, n19652, n19653, n19654,
    n19655, n19656, n19657, n19658, n19659, n19660,
    n19661, n19662, n19663, n19664, n19665, n19666,
    n19667, n19668, n19669, n19670, n19671, n19672,
    n19673, n19674, n19675, n19676, n19677, n19678,
    n19679, n19680, n19681, n19682, n19683, n19684,
    n19685, n19686, n19687, n19688, n19689, n19690,
    n19691, n19692, n19693, n19694, n19695, n19696,
    n19697, n19698, n19699, n19700, n19701, n19702,
    n19703, n19704, n19705, n19706, n19707, n19708,
    n19709, n19710, n19711, n19712, n19713, n19714,
    n19715, n19716, n19717, n19718, n19719, n19720,
    n19721, n19722, n19723, n19724, n19725, n19726,
    n19727, n19728, n19729, n19730, n19731, n19732,
    n19733, n19734, n19735, n19736, n19737, n19738,
    n19739, n19740, n19741, n19742, n19743, n19744,
    n19745, n19746, n19747, n19748, n19749, n19750,
    n19751, n19752, n19753, n19754, n19755, n19756,
    n19757, n19758, n19759, n19760, n19761, n19762,
    n19763, n19764, n19765, n19766, n19767, n19768,
    n19769, n19770, n19771, n19772, n19773, n19774,
    n19775, n19776, n19777, n19778, n19779, n19780,
    n19781, n19782, n19783, n19784, n19785, n19786,
    n19787, n19788, n19789, n19790, n19791, n19792,
    n19793, n19794, n19795, n19796, n19797, n19798,
    n19799, n19800, n19801, n19802, n19803, n19804,
    n19805, n19806, n19807, n19808, n19810, n19811,
    n19812, n19813, n19814, n19815, n19816, n19817,
    n19818, n19819, n19820, n19821, n19822, n19823,
    n19824, n19825, n19826, n19827, n19828, n19829,
    n19830, n19831, n19832, n19833, n19834, n19835,
    n19836, n19837, n19838, n19839, n19840, n19841,
    n19842, n19843, n19844, n19845, n19846, n19847,
    n19848, n19849, n19850, n19851, n19852, n19853,
    n19854, n19855, n19856, n19857, n19858, n19859,
    n19860, n19861, n19862, n19863, n19864, n19865,
    n19866, n19867, n19868, n19869, n19870, n19871,
    n19872, n19873, n19874, n19875, n19876, n19877,
    n19878, n19879, n19880, n19881, n19882, n19883,
    n19884, n19885, n19886, n19887, n19888, n19889,
    n19890, n19891, n19892, n19893, n19894, n19895,
    n19896, n19897, n19898, n19899, n19900, n19901,
    n19902, n19903, n19904, n19905, n19906, n19907,
    n19908, n19909, n19910, n19911, n19912, n19913,
    n19914, n19915, n19916, n19917, n19918, n19919,
    n19920, n19921, n19922, n19923, n19924, n19925,
    n19926, n19927, n19928, n19929, n19930, n19931,
    n19932, n19933, n19934, n19935, n19936, n19937,
    n19938, n19939, n19940, n19941, n19942, n19943,
    n19944, n19945, n19946, n19947, n19948, n19949,
    n19950, n19951, n19952, n19953, n19954, n19955,
    n19956, n19957, n19958, n19959, n19960, n19961,
    n19962, n19963, n19964, n19965, n19966, n19967,
    n19968, n19969, n19970, n19971, n19972, n19973,
    n19974, n19975, n19976, n19977, n19978, n19979,
    n19980, n19981, n19982, n19983, n19984, n19985,
    n19986, n19987, n19988, n19989, n19990, n19991,
    n19992, n19993, n19994, n19995, n19996, n19997,
    n19998, n19999, n20000, n20001, n20002, n20003,
    n20004, n20005, n20006, n20007, n20008, n20009,
    n20010, n20011, n20012, n20013, n20014, n20015,
    n20016, n20017, n20018, n20019, n20020, n20021,
    n20022, n20023, n20024, n20025, n20026, n20027,
    n20028, n20029, n20030, n20031, n20032, n20033,
    n20034, n20035, n20036, n20037, n20038, n20039,
    n20040, n20041, n20042, n20043, n20044, n20045,
    n20046, n20047, n20048, n20049, n20050, n20051,
    n20052, n20053, n20054, n20055, n20056, n20057,
    n20058, n20059, n20060, n20061, n20062, n20063,
    n20064, n20065, n20066, n20067, n20068, n20069,
    n20070, n20071, n20072, n20073, n20074, n20075,
    n20076, n20077, n20078, n20079, n20080, n20081,
    n20082, n20083, n20084, n20085, n20086, n20087,
    n20088, n20090, n20091, n20092, n20093, n20094,
    n20095, n20096, n20097, n20098, n20099, n20100,
    n20101, n20102, n20103, n20104, n20105, n20106,
    n20107, n20108, n20109, n20110, n20111, n20112,
    n20113, n20114, n20115, n20116, n20117, n20118,
    n20119, n20120, n20121, n20122, n20123, n20124,
    n20125, n20126, n20127, n20128, n20129, n20130,
    n20131, n20132, n20133, n20134, n20135, n20136,
    n20137, n20138, n20139, n20140, n20141, n20142,
    n20143, n20144, n20145, n20146, n20147, n20148,
    n20149, n20150, n20151, n20152, n20153, n20154,
    n20155, n20156, n20157, n20158, n20159, n20160,
    n20161, n20162, n20163, n20164, n20165, n20166,
    n20167, n20168, n20169, n20170, n20171, n20172,
    n20173, n20174, n20175, n20176, n20177, n20178,
    n20179, n20180, n20181, n20182, n20183, n20184,
    n20185, n20186, n20187, n20188, n20189, n20190,
    n20191, n20192, n20193, n20194, n20195, n20196,
    n20197, n20198, n20199, n20200, n20201, n20202,
    n20203, n20204, n20205, n20206, n20207, n20208,
    n20209, n20210, n20211, n20212, n20213, n20214,
    n20215, n20216, n20217, n20218, n20219, n20220,
    n20221, n20222, n20223, n20224, n20225, n20226,
    n20227, n20228, n20229, n20230, n20231, n20232,
    n20233, n20234, n20235, n20236, n20237, n20238,
    n20239, n20240, n20241, n20242, n20243, n20244,
    n20245, n20246, n20247, n20248, n20249, n20250,
    n20251, n20252, n20253, n20254, n20255, n20256,
    n20257, n20258, n20259, n20260, n20261, n20262,
    n20263, n20264, n20265, n20266, n20267, n20268,
    n20269, n20270, n20271, n20272, n20273, n20274,
    n20275, n20276, n20277, n20278, n20279, n20280,
    n20281, n20282, n20283, n20284, n20285, n20286,
    n20287, n20288, n20289, n20290, n20291, n20292,
    n20293, n20294, n20295, n20296, n20297, n20298,
    n20299, n20300, n20301, n20302, n20303, n20304,
    n20305, n20306, n20307, n20308, n20309, n20310,
    n20311, n20312, n20313, n20314, n20315, n20316,
    n20317, n20318, n20319, n20320, n20321, n20322,
    n20323, n20324, n20325, n20326, n20327, n20328,
    n20329, n20330, n20331, n20332, n20333, n20334,
    n20335, n20336, n20337, n20338, n20339, n20340,
    n20341, n20342, n20343, n20344, n20345, n20346,
    n20347, n20348, n20349, n20350, n20351, n20352,
    n20353, n20354, n20355, n20356, n20357, n20358,
    n20359, n20360, n20361, n20362, n20363, n20364,
    n20365, n20366, n20368, n20369, n20370, n20371,
    n20372, n20373, n20374, n20375, n20376, n20377,
    n20378, n20379, n20380, n20381, n20382, n20383,
    n20384, n20385, n20386, n20387, n20388, n20389,
    n20390, n20391, n20392, n20393, n20394, n20395,
    n20396, n20397, n20398, n20399, n20400, n20401,
    n20402, n20403, n20404, n20405, n20406, n20407,
    n20408, n20409, n20410, n20411, n20412, n20413,
    n20414, n20415, n20416, n20417, n20418, n20419,
    n20420, n20421, n20422, n20423, n20424, n20425,
    n20426, n20427, n20428, n20429, n20430, n20431,
    n20432, n20433, n20434, n20435, n20436, n20437,
    n20438, n20439, n20440, n20441, n20442, n20443,
    n20444, n20445, n20446, n20447, n20448, n20449,
    n20450, n20451, n20452, n20453, n20454, n20455,
    n20456, n20457, n20458, n20459, n20460, n20461,
    n20462, n20463, n20464, n20465, n20466, n20467,
    n20468, n20469, n20470, n20471, n20472, n20473,
    n20474, n20475, n20476, n20477, n20478, n20479,
    n20480, n20481, n20482, n20483, n20484, n20485,
    n20486, n20487, n20488, n20489, n20490, n20491,
    n20492, n20493, n20494, n20495, n20496, n20497,
    n20498, n20499, n20500, n20501, n20502, n20503,
    n20504, n20505, n20506, n20507, n20508, n20509,
    n20510, n20511, n20512, n20513, n20514, n20515,
    n20516, n20517, n20518, n20519, n20520, n20521,
    n20522, n20523, n20524, n20525, n20526, n20527,
    n20528, n20529, n20530, n20531, n20532, n20533,
    n20534, n20535, n20536, n20537, n20538, n20539,
    n20540, n20541, n20542, n20543, n20544, n20545,
    n20546, n20547, n20548, n20549, n20550, n20551,
    n20552, n20553, n20554, n20555, n20556, n20557,
    n20558, n20559, n20560, n20561, n20562, n20563,
    n20564, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581,
    n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599,
    n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617,
    n20618, n20619, n20620, n20621, n20622, n20623,
    n20624, n20625, n20626, n20627, n20628, n20629,
    n20630, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20645, n20646, n20647, n20648,
    n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660,
    n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20675, n20676, n20677, n20678,
    n20679, n20680, n20681, n20682, n20683, n20684,
    n20685, n20686, n20687, n20688, n20689, n20690,
    n20691, n20692, n20693, n20694, n20695, n20696,
    n20697, n20698, n20699, n20700, n20701, n20702,
    n20703, n20704, n20705, n20706, n20707, n20708,
    n20709, n20710, n20711, n20712, n20713, n20714,
    n20715, n20716, n20717, n20718, n20719, n20720,
    n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732,
    n20733, n20734, n20735, n20736, n20737, n20738,
    n20739, n20740, n20741, n20742, n20743, n20744,
    n20745, n20746, n20747, n20748, n20749, n20750,
    n20751, n20752, n20753, n20754, n20755, n20756,
    n20757, n20758, n20759, n20760, n20761, n20762,
    n20763, n20764, n20765, n20766, n20767, n20768,
    n20769, n20770, n20771, n20772, n20773, n20774,
    n20775, n20776, n20777, n20778, n20779, n20780,
    n20781, n20782, n20783, n20784, n20785, n20786,
    n20787, n20788, n20789, n20790, n20791, n20792,
    n20793, n20794, n20795, n20796, n20797, n20798,
    n20799, n20800, n20801, n20802, n20803, n20804,
    n20805, n20806, n20807, n20808, n20809, n20810,
    n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822,
    n20823, n20824, n20825, n20826, n20827, n20828,
    n20829, n20830, n20831, n20832, n20833, n20834,
    n20835, n20836, n20837, n20838, n20839, n20840,
    n20841, n20842, n20843, n20844, n20845, n20846,
    n20847, n20848, n20849, n20850, n20851, n20852,
    n20853, n20854, n20855, n20856, n20857, n20858,
    n20859, n20860, n20861, n20862, n20863, n20864,
    n20865, n20866, n20867, n20868, n20869, n20870,
    n20871, n20872, n20873, n20874, n20875, n20876,
    n20877, n20878, n20879, n20880, n20881, n20882,
    n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20893, n20894, n20895,
    n20896, n20897, n20898, n20899, n20900, n20901,
    n20902, n20903, n20904, n20905, n20906, n20907,
    n20908, n20909, n20910, n20911, n20912, n20913,
    n20914, n20915, n20916, n20917, n20918, n20919,
    n20920, n20921, n20922, n20923, n20924, n20925,
    n20926, n20927, n20928, n20929, n20930, n20931,
    n20932, n20933, n20934, n20935, n20936, n20937,
    n20938, n20939, n20940, n20941, n20942, n20943,
    n20944, n20945, n20946, n20947, n20948, n20949,
    n20950, n20951, n20952, n20953, n20954, n20955,
    n20956, n20957, n20958, n20959, n20960, n20961,
    n20962, n20963, n20964, n20965, n20966, n20967,
    n20968, n20969, n20970, n20971, n20972, n20973,
    n20974, n20975, n20976, n20977, n20978, n20979,
    n20980, n20981, n20982, n20983, n20984, n20985,
    n20986, n20987, n20988, n20989, n20990, n20991,
    n20992, n20993, n20994, n20995, n20996, n20997,
    n20998, n20999, n21000, n21001, n21002, n21003,
    n21004, n21005, n21006, n21007, n21008, n21009,
    n21010, n21011, n21012, n21013, n21014, n21015,
    n21016, n21017, n21018, n21019, n21020, n21021,
    n21022, n21023, n21024, n21025, n21026, n21027,
    n21028, n21029, n21030, n21031, n21032, n21033,
    n21034, n21035, n21036, n21037, n21038, n21039,
    n21040, n21041, n21042, n21043, n21044, n21045,
    n21046, n21047, n21048, n21049, n21050, n21051,
    n21052, n21053, n21054, n21055, n21056, n21057,
    n21058, n21059, n21060, n21061, n21062, n21063,
    n21064, n21065, n21066, n21067, n21068, n21069,
    n21070, n21071, n21072, n21073, n21074, n21075,
    n21076, n21077, n21078, n21079, n21080, n21081,
    n21082, n21083, n21084, n21085, n21086, n21087,
    n21088, n21089, n21090, n21091, n21092, n21093,
    n21094, n21095, n21096, n21097, n21098, n21099,
    n21100, n21101, n21102, n21103, n21104, n21105,
    n21106, n21107, n21108, n21109, n21110, n21111,
    n21112, n21113, n21114, n21115, n21116, n21117,
    n21118, n21119, n21120, n21121, n21122, n21123,
    n21124, n21125, n21126, n21127, n21128, n21129,
    n21130, n21131, n21132, n21133, n21134, n21135,
    n21136, n21137, n21138, n21139, n21140, n21141,
    n21142, n21143, n21144, n21145, n21146, n21147,
    n21149, n21150, n21151, n21152, n21153, n21154,
    n21155, n21156, n21157, n21158, n21159, n21160,
    n21161, n21162, n21163, n21164, n21165, n21166,
    n21167, n21168, n21169, n21170, n21171, n21172,
    n21173, n21174, n21175, n21176, n21177, n21178,
    n21179, n21180, n21181, n21182, n21183, n21184,
    n21185, n21186, n21187, n21188, n21189, n21190,
    n21191, n21192, n21193, n21194, n21195, n21196,
    n21197, n21198, n21199, n21200, n21201, n21202,
    n21203, n21204, n21205, n21206, n21207, n21208,
    n21209, n21210, n21211, n21212, n21213, n21214,
    n21215, n21216, n21217, n21218, n21219, n21220,
    n21221, n21222, n21223, n21224, n21225, n21226,
    n21227, n21228, n21229, n21230, n21231, n21232,
    n21233, n21234, n21235, n21236, n21237, n21238,
    n21239, n21240, n21241, n21242, n21243, n21244,
    n21245, n21246, n21247, n21248, n21249, n21250,
    n21251, n21252, n21253, n21254, n21255, n21256,
    n21257, n21258, n21259, n21260, n21261, n21262,
    n21263, n21264, n21265, n21266, n21267, n21268,
    n21269, n21270, n21271, n21272, n21273, n21274,
    n21275, n21276, n21277, n21278, n21279, n21280,
    n21281, n21282, n21283, n21284, n21285, n21286,
    n21287, n21288, n21289, n21290, n21291, n21292,
    n21293, n21294, n21295, n21296, n21297, n21298,
    n21299, n21300, n21301, n21302, n21303, n21304,
    n21305, n21306, n21307, n21308, n21309, n21310,
    n21311, n21312, n21313, n21314, n21315, n21316,
    n21317, n21318, n21319, n21320, n21321, n21322,
    n21323, n21324, n21325, n21326, n21327, n21328,
    n21329, n21330, n21331, n21332, n21333, n21334,
    n21335, n21336, n21337, n21338, n21339, n21340,
    n21341, n21342, n21343, n21344, n21345, n21346,
    n21347, n21348, n21349, n21350, n21351, n21352,
    n21353, n21354, n21355, n21356, n21357, n21358,
    n21359, n21360, n21361, n21362, n21363, n21364,
    n21365, n21366, n21367, n21368, n21369, n21370,
    n21371, n21372, n21373, n21374, n21375, n21376,
    n21377, n21378, n21379, n21380, n21381, n21382,
    n21383, n21384, n21385, n21386, n21387, n21388,
    n21389, n21390, n21392, n21393, n21394, n21395,
    n21396, n21397, n21398, n21399, n21400, n21401,
    n21402, n21403, n21404, n21405, n21406, n21407,
    n21408, n21409, n21410, n21411, n21412, n21413,
    n21414, n21415, n21416, n21417, n21418, n21419,
    n21420, n21421, n21422, n21423, n21424, n21425,
    n21426, n21427, n21428, n21429, n21430, n21431,
    n21432, n21433, n21434, n21435, n21436, n21437,
    n21438, n21439, n21440, n21441, n21442, n21443,
    n21444, n21445, n21446, n21447, n21448, n21449,
    n21450, n21451, n21452, n21453, n21454, n21455,
    n21456, n21457, n21458, n21459, n21460, n21461,
    n21462, n21463, n21464, n21465, n21466, n21467,
    n21468, n21469, n21470, n21471, n21472, n21473,
    n21474, n21475, n21476, n21477, n21478, n21479,
    n21480, n21481, n21482, n21483, n21484, n21485,
    n21486, n21487, n21488, n21489, n21490, n21491,
    n21492, n21493, n21494, n21495, n21496, n21497,
    n21498, n21499, n21500, n21501, n21502, n21503,
    n21504, n21505, n21506, n21507, n21508, n21509,
    n21510, n21511, n21512, n21513, n21514, n21515,
    n21516, n21517, n21518, n21519, n21520, n21521,
    n21522, n21523, n21524, n21525, n21526, n21527,
    n21528, n21529, n21530, n21531, n21532, n21533,
    n21534, n21535, n21536, n21537, n21538, n21539,
    n21540, n21541, n21542, n21543, n21544, n21545,
    n21546, n21547, n21548, n21549, n21550, n21551,
    n21552, n21553, n21554, n21555, n21556, n21557,
    n21558, n21559, n21560, n21561, n21562, n21563,
    n21564, n21565, n21566, n21567, n21568, n21569,
    n21570, n21571, n21572, n21573, n21574, n21575,
    n21576, n21577, n21578, n21579, n21580, n21581,
    n21582, n21583, n21584, n21585, n21586, n21587,
    n21588, n21589, n21590, n21591, n21592, n21593,
    n21594, n21595, n21596, n21597, n21598, n21599,
    n21600, n21601, n21602, n21603, n21604, n21605,
    n21606, n21607, n21608, n21609, n21610, n21611,
    n21612, n21613, n21614, n21615, n21616, n21617,
    n21618, n21619, n21620, n21621, n21622, n21623,
    n21624, n21625, n21626, n21627, n21628, n21629,
    n21630, n21631, n21632, n21634, n21635, n21636,
    n21637, n21638, n21639, n21640, n21641, n21642,
    n21643, n21644, n21645, n21646, n21647, n21648,
    n21649, n21650, n21651, n21652, n21653, n21654,
    n21655, n21656, n21657, n21658, n21659, n21660,
    n21661, n21662, n21663, n21664, n21665, n21666,
    n21667, n21668, n21669, n21670, n21671, n21672,
    n21673, n21674, n21675, n21676, n21677, n21678,
    n21679, n21680, n21681, n21682, n21683, n21684,
    n21685, n21686, n21687, n21688, n21689, n21690,
    n21691, n21692, n21693, n21694, n21695, n21696,
    n21697, n21698, n21699, n21700, n21701, n21702,
    n21703, n21704, n21705, n21706, n21707, n21708,
    n21709, n21710, n21711, n21712, n21713, n21714,
    n21715, n21716, n21717, n21718, n21719, n21720,
    n21721, n21722, n21723, n21724, n21725, n21726,
    n21727, n21728, n21729, n21730, n21731, n21732,
    n21733, n21734, n21735, n21736, n21737, n21738,
    n21739, n21740, n21741, n21742, n21743, n21744,
    n21745, n21746, n21747, n21748, n21749, n21750,
    n21751, n21752, n21753, n21754, n21755, n21756,
    n21757, n21758, n21759, n21760, n21761, n21762,
    n21763, n21764, n21765, n21766, n21767, n21768,
    n21769, n21770, n21771, n21772, n21773, n21774,
    n21775, n21776, n21777, n21778, n21779, n21780,
    n21781, n21782, n21783, n21784, n21785, n21786,
    n21787, n21788, n21789, n21790, n21791, n21792,
    n21793, n21794, n21795, n21796, n21797, n21798,
    n21799, n21800, n21801, n21802, n21803, n21804,
    n21805, n21806, n21807, n21808, n21809, n21810,
    n21811, n21812, n21813, n21814, n21815, n21816,
    n21817, n21818, n21819, n21820, n21821, n21822,
    n21823, n21824, n21825, n21826, n21827, n21828,
    n21829, n21830, n21831, n21832, n21833, n21834,
    n21835, n21836, n21837, n21838, n21839, n21840,
    n21841, n21842, n21843, n21844, n21845, n21846,
    n21847, n21848, n21849, n21850, n21851, n21852,
    n21853, n21854, n21855, n21856, n21857, n21858,
    n21859, n21860, n21861, n21862, n21863, n21864,
    n21865, n21866, n21867, n21868, n21869, n21870,
    n21872, n21873, n21874, n21875, n21876, n21877,
    n21878, n21879, n21880, n21881, n21882, n21883,
    n21884, n21885, n21886, n21887, n21888, n21889,
    n21890, n21891, n21892, n21893, n21894, n21895,
    n21896, n21897, n21898, n21899, n21900, n21901,
    n21902, n21903, n21904, n21905, n21906, n21907,
    n21908, n21909, n21910, n21911, n21912, n21913,
    n21914, n21915, n21916, n21917, n21918, n21919,
    n21920, n21921, n21922, n21923, n21924, n21925,
    n21926, n21927, n21928, n21929, n21930, n21931,
    n21932, n21933, n21934, n21935, n21936, n21937,
    n21938, n21939, n21940, n21941, n21942, n21943,
    n21944, n21945, n21946, n21947, n21948, n21949,
    n21950, n21951, n21952, n21953, n21954, n21955,
    n21956, n21957, n21958, n21959, n21960, n21961,
    n21962, n21963, n21964, n21965, n21966, n21967,
    n21968, n21969, n21970, n21971, n21972, n21973,
    n21974, n21975, n21976, n21977, n21978, n21979,
    n21980, n21981, n21982, n21983, n21984, n21985,
    n21986, n21987, n21988, n21989, n21990, n21991,
    n21992, n21993, n21994, n21995, n21996, n21997,
    n21998, n21999, n22000, n22001, n22002, n22003,
    n22004, n22005, n22006, n22007, n22008, n22009,
    n22010, n22011, n22012, n22013, n22014, n22015,
    n22016, n22017, n22018, n22019, n22020, n22021,
    n22022, n22023, n22024, n22025, n22026, n22027,
    n22028, n22029, n22030, n22031, n22032, n22033,
    n22034, n22035, n22036, n22037, n22038, n22039,
    n22040, n22041, n22042, n22043, n22044, n22045,
    n22046, n22047, n22048, n22049, n22050, n22051,
    n22052, n22053, n22054, n22055, n22056, n22057,
    n22058, n22059, n22060, n22061, n22062, n22063,
    n22064, n22065, n22066, n22067, n22068, n22069,
    n22070, n22071, n22072, n22073, n22074, n22075,
    n22076, n22077, n22078, n22079, n22080, n22081,
    n22082, n22083, n22084, n22085, n22086, n22087,
    n22088, n22089, n22090, n22091, n22092, n22093,
    n22094, n22095, n22096, n22097, n22098, n22100,
    n22101, n22102, n22103, n22104, n22105, n22106,
    n22107, n22108, n22109, n22110, n22111, n22112,
    n22113, n22114, n22115, n22116, n22117, n22118,
    n22119, n22120, n22121, n22122, n22123, n22124,
    n22125, n22126, n22127, n22128, n22129, n22130,
    n22131, n22132, n22133, n22134, n22135, n22136,
    n22137, n22138, n22139, n22140, n22141, n22142,
    n22143, n22144, n22145, n22146, n22147, n22148,
    n22149, n22150, n22151, n22152, n22153, n22154,
    n22155, n22156, n22157, n22158, n22159, n22160,
    n22161, n22162, n22163, n22164, n22165, n22166,
    n22167, n22168, n22169, n22170, n22171, n22172,
    n22173, n22174, n22175, n22176, n22177, n22178,
    n22179, n22180, n22181, n22182, n22183, n22184,
    n22185, n22186, n22187, n22188, n22189, n22190,
    n22191, n22192, n22193, n22194, n22195, n22196,
    n22197, n22198, n22199, n22200, n22201, n22202,
    n22203, n22204, n22205, n22206, n22207, n22208,
    n22209, n22210, n22211, n22212, n22213, n22214,
    n22215, n22216, n22217, n22218, n22219, n22220,
    n22221, n22222, n22223, n22224, n22225, n22226,
    n22227, n22228, n22229, n22230, n22231, n22232,
    n22233, n22234, n22235, n22236, n22237, n22238,
    n22239, n22240, n22241, n22242, n22243, n22244,
    n22245, n22246, n22247, n22248, n22249, n22250,
    n22251, n22252, n22253, n22254, n22255, n22256,
    n22257, n22258, n22259, n22260, n22261, n22262,
    n22263, n22264, n22265, n22266, n22267, n22268,
    n22269, n22270, n22271, n22272, n22273, n22274,
    n22275, n22276, n22277, n22278, n22279, n22280,
    n22281, n22282, n22283, n22284, n22285, n22286,
    n22287, n22288, n22289, n22290, n22291, n22292,
    n22293, n22294, n22295, n22296, n22297, n22298,
    n22299, n22300, n22301, n22302, n22303, n22304,
    n22305, n22306, n22307, n22308, n22309, n22310,
    n22311, n22312, n22313, n22314, n22315, n22316,
    n22317, n22318, n22319, n22320, n22321, n22322,
    n22323, n22324, n22325, n22327, n22328, n22329,
    n22330, n22331, n22332, n22333, n22334, n22335,
    n22336, n22337, n22338, n22339, n22340, n22341,
    n22342, n22343, n22344, n22345, n22346, n22347,
    n22348, n22349, n22350, n22351, n22352, n22353,
    n22354, n22355, n22356, n22357, n22358, n22359,
    n22360, n22361, n22362, n22363, n22364, n22365,
    n22366, n22367, n22368, n22369, n22370, n22371,
    n22372, n22373, n22374, n22375, n22376, n22377,
    n22378, n22379, n22380, n22381, n22382, n22383,
    n22384, n22385, n22386, n22387, n22388, n22389,
    n22390, n22391, n22392, n22393, n22394, n22395,
    n22396, n22397, n22398, n22399, n22400, n22401,
    n22402, n22403, n22404, n22405, n22406, n22407,
    n22408, n22409, n22410, n22411, n22412, n22413,
    n22414, n22415, n22416, n22417, n22418, n22419,
    n22420, n22421, n22422, n22423, n22424, n22425,
    n22426, n22427, n22428, n22429, n22430, n22431,
    n22432, n22433, n22434, n22435, n22436, n22437,
    n22438, n22439, n22440, n22441, n22442, n22443,
    n22444, n22445, n22446, n22447, n22448, n22449,
    n22450, n22451, n22452, n22453, n22454, n22455,
    n22456, n22457, n22458, n22459, n22460, n22461,
    n22462, n22463, n22464, n22465, n22466, n22467,
    n22468, n22469, n22470, n22471, n22472, n22473,
    n22474, n22475, n22476, n22477, n22478, n22479,
    n22480, n22481, n22482, n22483, n22484, n22485,
    n22486, n22487, n22488, n22489, n22490, n22491,
    n22492, n22493, n22494, n22495, n22496, n22497,
    n22498, n22499, n22500, n22501, n22502, n22503,
    n22504, n22505, n22506, n22507, n22508, n22509,
    n22510, n22511, n22512, n22513, n22514, n22515,
    n22516, n22517, n22518, n22519, n22520, n22521,
    n22522, n22523, n22524, n22525, n22526, n22527,
    n22528, n22529, n22530, n22531, n22532, n22533,
    n22534, n22535, n22536, n22537, n22538, n22539,
    n22540, n22541, n22542, n22543, n22545, n22546,
    n22547, n22548, n22549, n22550, n22551, n22552,
    n22553, n22554, n22555, n22556, n22557, n22558,
    n22559, n22560, n22561, n22562, n22563, n22564,
    n22565, n22566, n22567, n22568, n22569, n22570,
    n22571, n22572, n22573, n22574, n22575, n22576,
    n22577, n22578, n22579, n22580, n22581, n22582,
    n22583, n22584, n22585, n22586, n22587, n22588,
    n22589, n22590, n22591, n22592, n22593, n22594,
    n22595, n22596, n22597, n22598, n22599, n22600,
    n22601, n22602, n22603, n22604, n22605, n22606,
    n22607, n22608, n22609, n22610, n22611, n22612,
    n22613, n22614, n22615, n22616, n22617, n22618,
    n22619, n22620, n22621, n22622, n22623, n22624,
    n22625, n22626, n22627, n22628, n22629, n22630,
    n22631, n22632, n22633, n22634, n22635, n22636,
    n22637, n22638, n22639, n22640, n22641, n22642,
    n22643, n22644, n22645, n22646, n22647, n22648,
    n22649, n22650, n22651, n22652, n22653, n22654,
    n22655, n22656, n22657, n22658, n22659, n22660,
    n22661, n22662, n22663, n22664, n22665, n22666,
    n22667, n22668, n22669, n22670, n22671, n22672,
    n22673, n22674, n22675, n22676, n22677, n22678,
    n22679, n22680, n22681, n22682, n22683, n22684,
    n22685, n22686, n22687, n22688, n22689, n22690,
    n22691, n22692, n22693, n22694, n22695, n22696,
    n22697, n22698, n22699, n22700, n22701, n22702,
    n22703, n22704, n22705, n22706, n22707, n22708,
    n22709, n22710, n22711, n22712, n22713, n22714,
    n22715, n22716, n22717, n22718, n22719, n22720,
    n22721, n22722, n22723, n22724, n22725, n22726,
    n22727, n22728, n22729, n22730, n22731, n22732,
    n22733, n22734, n22735, n22736, n22737, n22738,
    n22739, n22740, n22741, n22742, n22743, n22744,
    n22745, n22746, n22747, n22748, n22749, n22750,
    n22751, n22752, n22754, n22755, n22756, n22757,
    n22758, n22759, n22760, n22761, n22762, n22763,
    n22764, n22765, n22766, n22767, n22768, n22769,
    n22770, n22771, n22772, n22773, n22774, n22775,
    n22776, n22777, n22778, n22779, n22780, n22781,
    n22782, n22783, n22784, n22785, n22786, n22787,
    n22788, n22789, n22790, n22791, n22792, n22793,
    n22794, n22795, n22796, n22797, n22798, n22799,
    n22800, n22801, n22802, n22803, n22804, n22805,
    n22806, n22807, n22808, n22809, n22810, n22811,
    n22812, n22813, n22814, n22815, n22816, n22817,
    n22818, n22819, n22820, n22821, n22822, n22823,
    n22824, n22825, n22826, n22827, n22828, n22829,
    n22830, n22831, n22832, n22833, n22834, n22835,
    n22836, n22837, n22838, n22839, n22840, n22841,
    n22842, n22843, n22844, n22845, n22846, n22847,
    n22848, n22849, n22850, n22851, n22852, n22853,
    n22854, n22855, n22856, n22857, n22858, n22859,
    n22860, n22861, n22862, n22863, n22864, n22865,
    n22866, n22867, n22868, n22869, n22870, n22871,
    n22872, n22873, n22874, n22875, n22876, n22877,
    n22878, n22879, n22880, n22881, n22882, n22883,
    n22884, n22885, n22886, n22887, n22888, n22889,
    n22890, n22891, n22892, n22893, n22894, n22895,
    n22896, n22897, n22898, n22899, n22900, n22901,
    n22902, n22903, n22904, n22905, n22906, n22907,
    n22908, n22909, n22910, n22911, n22912, n22913,
    n22914, n22915, n22916, n22917, n22918, n22919,
    n22920, n22921, n22922, n22923, n22924, n22925,
    n22926, n22927, n22928, n22929, n22930, n22931,
    n22932, n22933, n22934, n22935, n22936, n22937,
    n22938, n22939, n22940, n22941, n22942, n22943,
    n22944, n22945, n22946, n22947, n22948, n22949,
    n22950, n22951, n22952, n22953, n22954, n22955,
    n22956, n22957, n22958, n22959, n22960, n22961,
    n22963, n22964, n22965, n22966, n22967, n22968,
    n22969, n22970, n22971, n22972, n22973, n22974,
    n22975, n22976, n22977, n22978, n22979, n22980,
    n22981, n22982, n22983, n22984, n22985, n22986,
    n22987, n22988, n22989, n22990, n22991, n22992,
    n22993, n22994, n22995, n22996, n22997, n22998,
    n22999, n23000, n23001, n23002, n23003, n23004,
    n23005, n23006, n23007, n23008, n23009, n23010,
    n23011, n23012, n23013, n23014, n23015, n23016,
    n23017, n23018, n23019, n23020, n23021, n23022,
    n23023, n23024, n23025, n23026, n23027, n23028,
    n23029, n23030, n23031, n23032, n23033, n23034,
    n23035, n23036, n23037, n23038, n23039, n23040,
    n23041, n23042, n23043, n23044, n23045, n23046,
    n23047, n23048, n23049, n23050, n23051, n23052,
    n23053, n23054, n23055, n23056, n23057, n23058,
    n23059, n23060, n23061, n23062, n23063, n23064,
    n23065, n23066, n23067, n23068, n23069, n23070,
    n23071, n23072, n23073, n23074, n23075, n23076,
    n23077, n23078, n23079, n23080, n23081, n23082,
    n23083, n23084, n23085, n23086, n23087, n23088,
    n23089, n23090, n23091, n23092, n23093, n23094,
    n23095, n23096, n23097, n23098, n23099, n23100,
    n23101, n23102, n23103, n23104, n23105, n23106,
    n23107, n23108, n23109, n23110, n23111, n23112,
    n23113, n23114, n23115, n23116, n23117, n23118,
    n23119, n23120, n23121, n23122, n23123, n23124,
    n23125, n23126, n23127, n23128, n23129, n23130,
    n23131, n23132, n23133, n23134, n23135, n23136,
    n23137, n23138, n23139, n23140, n23141, n23142,
    n23143, n23144, n23145, n23146, n23147, n23148,
    n23149, n23150, n23151, n23152, n23153, n23154,
    n23155, n23156, n23157, n23158, n23159, n23160,
    n23161, n23163, n23164, n23165, n23166, n23167,
    n23168, n23169, n23170, n23171, n23172, n23173,
    n23174, n23175, n23176, n23177, n23178, n23179,
    n23180, n23181, n23182, n23183, n23184, n23185,
    n23186, n23187, n23188, n23189, n23190, n23191,
    n23192, n23193, n23194, n23195, n23196, n23197,
    n23198, n23199, n23200, n23201, n23202, n23203,
    n23204, n23205, n23206, n23207, n23208, n23209,
    n23210, n23211, n23212, n23213, n23214, n23215,
    n23216, n23217, n23218, n23219, n23220, n23221,
    n23222, n23223, n23224, n23225, n23226, n23227,
    n23228, n23229, n23230, n23231, n23232, n23233,
    n23234, n23235, n23236, n23237, n23238, n23239,
    n23240, n23241, n23242, n23243, n23244, n23245,
    n23246, n23247, n23248, n23249, n23250, n23251,
    n23252, n23253, n23254, n23255, n23256, n23257,
    n23258, n23259, n23260, n23261, n23262, n23263,
    n23264, n23265, n23266, n23267, n23268, n23269,
    n23270, n23271, n23272, n23273, n23274, n23275,
    n23276, n23277, n23278, n23279, n23280, n23281,
    n23282, n23283, n23284, n23285, n23286, n23287,
    n23288, n23289, n23290, n23291, n23292, n23293,
    n23294, n23295, n23296, n23297, n23298, n23299,
    n23300, n23301, n23302, n23303, n23304, n23305,
    n23306, n23307, n23308, n23309, n23310, n23311,
    n23312, n23313, n23314, n23315, n23316, n23317,
    n23318, n23319, n23320, n23321, n23322, n23323,
    n23324, n23325, n23326, n23327, n23328, n23329,
    n23330, n23331, n23332, n23333, n23334, n23335,
    n23336, n23337, n23338, n23339, n23340, n23341,
    n23342, n23343, n23344, n23345, n23346, n23347,
    n23348, n23349, n23350, n23351, n23352, n23354,
    n23355, n23356, n23357, n23358, n23359, n23360,
    n23361, n23362, n23363, n23364, n23365, n23366,
    n23367, n23368, n23369, n23370, n23371, n23372,
    n23373, n23374, n23375, n23376, n23377, n23378,
    n23379, n23380, n23381, n23382, n23383, n23384,
    n23385, n23386, n23387, n23388, n23389, n23390,
    n23391, n23392, n23393, n23394, n23395, n23396,
    n23397, n23398, n23399, n23400, n23401, n23402,
    n23403, n23404, n23405, n23406, n23407, n23408,
    n23409, n23410, n23411, n23412, n23413, n23414,
    n23415, n23416, n23417, n23418, n23419, n23420,
    n23421, n23422, n23423, n23424, n23425, n23426,
    n23427, n23428, n23429, n23430, n23431, n23432,
    n23433, n23434, n23435, n23436, n23437, n23438,
    n23439, n23440, n23441, n23442, n23443, n23444,
    n23445, n23446, n23447, n23448, n23449, n23450,
    n23451, n23452, n23453, n23454, n23455, n23456,
    n23457, n23458, n23459, n23460, n23461, n23462,
    n23463, n23464, n23465, n23466, n23467, n23468,
    n23469, n23470, n23471, n23472, n23473, n23474,
    n23475, n23476, n23477, n23478, n23479, n23480,
    n23481, n23482, n23483, n23484, n23485, n23486,
    n23487, n23488, n23489, n23490, n23491, n23492,
    n23493, n23494, n23495, n23496, n23497, n23498,
    n23499, n23500, n23501, n23502, n23503, n23504,
    n23505, n23506, n23507, n23508, n23509, n23510,
    n23511, n23512, n23513, n23514, n23515, n23516,
    n23517, n23518, n23519, n23520, n23521, n23522,
    n23523, n23524, n23525, n23526, n23527, n23528,
    n23529, n23530, n23531, n23532, n23533, n23534,
    n23535, n23536, n23537, n23538, n23539, n23540,
    n23541, n23543, n23544, n23545, n23546, n23547,
    n23548, n23549, n23550, n23551, n23552, n23553,
    n23554, n23555, n23556, n23557, n23558, n23559,
    n23560, n23561, n23562, n23563, n23564, n23565,
    n23566, n23567, n23568, n23569, n23570, n23571,
    n23572, n23573, n23574, n23575, n23576, n23577,
    n23578, n23579, n23580, n23581, n23582, n23583,
    n23584, n23585, n23586, n23587, n23588, n23589,
    n23590, n23591, n23592, n23593, n23594, n23595,
    n23596, n23597, n23598, n23599, n23600, n23601,
    n23602, n23603, n23604, n23605, n23606, n23607,
    n23608, n23609, n23610, n23611, n23612, n23613,
    n23614, n23615, n23616, n23617, n23618, n23619,
    n23620, n23621, n23622, n23623, n23624, n23625,
    n23626, n23627, n23628, n23629, n23630, n23631,
    n23632, n23633, n23634, n23635, n23636, n23637,
    n23638, n23639, n23640, n23641, n23642, n23643,
    n23644, n23645, n23646, n23647, n23648, n23649,
    n23650, n23651, n23652, n23653, n23654, n23655,
    n23656, n23657, n23658, n23659, n23660, n23661,
    n23662, n23663, n23664, n23665, n23666, n23667,
    n23668, n23669, n23670, n23671, n23672, n23673,
    n23674, n23675, n23676, n23677, n23678, n23679,
    n23680, n23681, n23682, n23683, n23684, n23685,
    n23686, n23687, n23688, n23689, n23690, n23691,
    n23692, n23693, n23694, n23695, n23696, n23697,
    n23698, n23699, n23700, n23701, n23702, n23703,
    n23704, n23705, n23706, n23707, n23708, n23709,
    n23710, n23711, n23712, n23713, n23714, n23715,
    n23716, n23717, n23718, n23719, n23720, n23722,
    n23723, n23724, n23725, n23726, n23727, n23728,
    n23729, n23730, n23731, n23732, n23733, n23734,
    n23735, n23736, n23737, n23738, n23739, n23740,
    n23741, n23742, n23743, n23744, n23745, n23746,
    n23747, n23748, n23749, n23750, n23751, n23752,
    n23753, n23754, n23755, n23756, n23757, n23758,
    n23759, n23760, n23761, n23762, n23763, n23764,
    n23765, n23766, n23767, n23768, n23769, n23770,
    n23771, n23772, n23773, n23774, n23775, n23776,
    n23777, n23778, n23779, n23780, n23781, n23782,
    n23783, n23784, n23785, n23786, n23787, n23788,
    n23789, n23790, n23791, n23792, n23793, n23794,
    n23795, n23796, n23797, n23798, n23799, n23800,
    n23801, n23802, n23803, n23804, n23805, n23806,
    n23807, n23808, n23809, n23810, n23811, n23812,
    n23813, n23814, n23815, n23816, n23817, n23818,
    n23819, n23820, n23821, n23822, n23823, n23824,
    n23825, n23826, n23827, n23828, n23829, n23830,
    n23831, n23832, n23833, n23834, n23835, n23836,
    n23837, n23838, n23839, n23840, n23841, n23842,
    n23843, n23844, n23845, n23846, n23847, n23848,
    n23849, n23850, n23851, n23852, n23853, n23854,
    n23855, n23856, n23857, n23858, n23859, n23860,
    n23861, n23862, n23863, n23864, n23865, n23866,
    n23867, n23868, n23869, n23870, n23871, n23872,
    n23873, n23874, n23875, n23876, n23877, n23878,
    n23879, n23880, n23881, n23882, n23883, n23884,
    n23885, n23886, n23887, n23888, n23889, n23890,
    n23891, n23892, n23893, n23894, n23896, n23897,
    n23898, n23899, n23900, n23901, n23902, n23903,
    n23904, n23905, n23906, n23907, n23908, n23909,
    n23910, n23911, n23912, n23913, n23914, n23915,
    n23916, n23917, n23918, n23919, n23920, n23921,
    n23922, n23923, n23924, n23925, n23926, n23927,
    n23928, n23929, n23930, n23931, n23932, n23933,
    n23934, n23935, n23936, n23937, n23938, n23939,
    n23940, n23941, n23942, n23943, n23944, n23945,
    n23946, n23947, n23948, n23949, n23950, n23951,
    n23952, n23953, n23954, n23955, n23956, n23957,
    n23958, n23959, n23960, n23961, n23962, n23963,
    n23964, n23965, n23966, n23967, n23968, n23969,
    n23970, n23971, n23972, n23973, n23974, n23975,
    n23976, n23977, n23978, n23979, n23980, n23981,
    n23982, n23983, n23984, n23985, n23986, n23987,
    n23988, n23989, n23990, n23991, n23992, n23993,
    n23994, n23995, n23996, n23997, n23998, n23999,
    n24000, n24001, n24002, n24003, n24004, n24005,
    n24006, n24007, n24008, n24009, n24010, n24011,
    n24012, n24013, n24014, n24015, n24016, n24017,
    n24018, n24019, n24020, n24021, n24022, n24023,
    n24024, n24025, n24026, n24027, n24028, n24029,
    n24030, n24031, n24032, n24033, n24034, n24035,
    n24036, n24037, n24038, n24039, n24040, n24041,
    n24042, n24043, n24044, n24045, n24046, n24047,
    n24048, n24049, n24050, n24051, n24052, n24053,
    n24054, n24055, n24056, n24057, n24058, n24059,
    n24060, n24061, n24062, n24063, n24064, n24065,
    n24067, n24068, n24069, n24070, n24071, n24072,
    n24073, n24074, n24075, n24076, n24077, n24078,
    n24079, n24080, n24081, n24082, n24083, n24084,
    n24085, n24086, n24087, n24088, n24089, n24090,
    n24091, n24092, n24093, n24094, n24095, n24096,
    n24097, n24098, n24099, n24100, n24101, n24102,
    n24103, n24104, n24105, n24106, n24107, n24108,
    n24109, n24110, n24111, n24112, n24113, n24114,
    n24115, n24116, n24117, n24118, n24119, n24120,
    n24121, n24122, n24123, n24124, n24125, n24126,
    n24127, n24128, n24129, n24130, n24131, n24132,
    n24133, n24134, n24135, n24136, n24137, n24138,
    n24139, n24140, n24141, n24142, n24143, n24144,
    n24145, n24146, n24147, n24148, n24149, n24150,
    n24151, n24152, n24153, n24154, n24155, n24156,
    n24157, n24158, n24159, n24160, n24161, n24162,
    n24163, n24164, n24165, n24166, n24167, n24168,
    n24169, n24170, n24171, n24172, n24173, n24174,
    n24175, n24176, n24177, n24178, n24179, n24180,
    n24181, n24182, n24183, n24184, n24185, n24186,
    n24187, n24188, n24189, n24190, n24191, n24192,
    n24193, n24194, n24195, n24196, n24197, n24198,
    n24199, n24200, n24201, n24202, n24203, n24204,
    n24205, n24206, n24207, n24208, n24209, n24210,
    n24211, n24212, n24213, n24214, n24215, n24216,
    n24217, n24218, n24219, n24220, n24221, n24222,
    n24223, n24224, n24225, n24226, n24227, n24228,
    n24230, n24231, n24232, n24233, n24234, n24235,
    n24236, n24237, n24238, n24239, n24240, n24241,
    n24242, n24243, n24244, n24245, n24246, n24247,
    n24248, n24249, n24250, n24251, n24252, n24253,
    n24254, n24255, n24256, n24257, n24258, n24259,
    n24260, n24261, n24262, n24263, n24264, n24265,
    n24266, n24267, n24268, n24269, n24270, n24271,
    n24272, n24273, n24274, n24275, n24276, n24277,
    n24278, n24279, n24280, n24281, n24282, n24283,
    n24284, n24285, n24286, n24287, n24288, n24289,
    n24290, n24291, n24292, n24293, n24294, n24295,
    n24296, n24297, n24298, n24299, n24300, n24301,
    n24302, n24303, n24304, n24305, n24306, n24307,
    n24308, n24309, n24310, n24311, n24312, n24313,
    n24314, n24315, n24316, n24317, n24318, n24319,
    n24320, n24321, n24322, n24323, n24324, n24325,
    n24326, n24327, n24328, n24329, n24330, n24331,
    n24332, n24333, n24334, n24335, n24336, n24337,
    n24338, n24339, n24340, n24341, n24342, n24343,
    n24344, n24345, n24346, n24347, n24348, n24349,
    n24350, n24351, n24352, n24353, n24354, n24355,
    n24356, n24357, n24358, n24359, n24360, n24361,
    n24362, n24363, n24364, n24365, n24366, n24367,
    n24368, n24369, n24370, n24371, n24372, n24373,
    n24374, n24375, n24376, n24377, n24378, n24379,
    n24380, n24381, n24382, n24383, n24384, n24386,
    n24387, n24388, n24389, n24390, n24391, n24392,
    n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404,
    n24405, n24406, n24407, n24408, n24409, n24410,
    n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422,
    n24423, n24424, n24425, n24426, n24427, n24428,
    n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440,
    n24441, n24442, n24443, n24444, n24445, n24446,
    n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24458,
    n24459, n24460, n24461, n24462, n24463, n24464,
    n24465, n24466, n24467, n24468, n24469, n24470,
    n24471, n24472, n24473, n24474, n24475, n24476,
    n24477, n24478, n24479, n24480, n24481, n24482,
    n24483, n24484, n24485, n24486, n24487, n24488,
    n24489, n24490, n24491, n24492, n24493, n24494,
    n24495, n24496, n24497, n24498, n24499, n24500,
    n24501, n24502, n24503, n24504, n24505, n24506,
    n24507, n24508, n24509, n24510, n24511, n24512,
    n24513, n24514, n24515, n24516, n24517, n24518,
    n24519, n24520, n24521, n24522, n24523, n24524,
    n24525, n24526, n24527, n24528, n24529, n24530,
    n24531, n24532, n24533, n24534, n24536, n24537,
    n24538, n24539, n24540, n24541, n24542, n24543,
    n24544, n24545, n24546, n24547, n24548, n24549,
    n24550, n24551, n24552, n24553, n24554, n24555,
    n24556, n24557, n24558, n24559, n24560, n24561,
    n24562, n24563, n24564, n24565, n24566, n24567,
    n24568, n24569, n24570, n24571, n24572, n24573,
    n24574, n24575, n24576, n24577, n24578, n24579,
    n24580, n24581, n24582, n24583, n24584, n24585,
    n24586, n24587, n24588, n24589, n24590, n24591,
    n24592, n24593, n24594, n24595, n24596, n24597,
    n24598, n24599, n24600, n24601, n24602, n24603,
    n24604, n24605, n24606, n24607, n24608, n24609,
    n24610, n24611, n24612, n24613, n24614, n24615,
    n24616, n24617, n24618, n24619, n24620, n24621,
    n24622, n24623, n24624, n24625, n24626, n24627,
    n24628, n24629, n24630, n24631, n24632, n24633,
    n24634, n24635, n24636, n24637, n24638, n24639,
    n24640, n24641, n24642, n24643, n24644, n24645,
    n24646, n24647, n24648, n24649, n24650, n24651,
    n24652, n24653, n24654, n24655, n24656, n24657,
    n24658, n24659, n24660, n24661, n24662, n24663,
    n24664, n24665, n24666, n24667, n24668, n24669,
    n24670, n24671, n24672, n24673, n24674, n24675,
    n24676, n24677, n24678, n24679, n24681, n24682,
    n24683, n24684, n24685, n24686, n24687, n24688,
    n24689, n24690, n24691, n24692, n24693, n24694,
    n24695, n24696, n24697, n24698, n24699, n24700,
    n24701, n24702, n24703, n24704, n24705, n24706,
    n24707, n24708, n24709, n24710, n24711, n24712,
    n24713, n24714, n24715, n24716, n24717, n24718,
    n24719, n24720, n24721, n24722, n24723, n24724,
    n24725, n24726, n24727, n24728, n24729, n24730,
    n24731, n24732, n24733, n24734, n24735, n24736,
    n24737, n24738, n24739, n24740, n24741, n24742,
    n24743, n24744, n24745, n24746, n24747, n24748,
    n24749, n24750, n24751, n24752, n24753, n24754,
    n24755, n24756, n24757, n24758, n24759, n24760,
    n24761, n24762, n24763, n24764, n24765, n24766,
    n24767, n24768, n24769, n24770, n24771, n24772,
    n24773, n24774, n24775, n24776, n24777, n24778,
    n24779, n24780, n24781, n24782, n24783, n24784,
    n24785, n24786, n24787, n24788, n24789, n24790,
    n24791, n24792, n24793, n24794, n24795, n24796,
    n24797, n24798, n24799, n24800, n24801, n24802,
    n24803, n24804, n24805, n24806, n24807, n24808,
    n24809, n24810, n24811, n24812, n24813, n24814,
    n24815, n24817, n24818, n24819, n24820, n24821,
    n24822, n24823, n24824, n24825, n24826, n24827,
    n24828, n24829, n24830, n24831, n24832, n24833,
    n24834, n24835, n24836, n24837, n24838, n24839,
    n24840, n24841, n24842, n24843, n24844, n24845,
    n24846, n24847, n24848, n24849, n24850, n24851,
    n24852, n24853, n24854, n24855, n24856, n24857,
    n24858, n24859, n24860, n24861, n24862, n24863,
    n24864, n24865, n24866, n24867, n24868, n24869,
    n24870, n24871, n24872, n24873, n24874, n24875,
    n24876, n24877, n24878, n24879, n24880, n24881,
    n24882, n24883, n24884, n24885, n24886, n24887,
    n24888, n24889, n24890, n24891, n24892, n24893,
    n24894, n24895, n24896, n24897, n24898, n24899,
    n24900, n24901, n24902, n24903, n24904, n24905,
    n24906, n24907, n24908, n24909, n24910, n24911,
    n24912, n24913, n24914, n24915, n24916, n24917,
    n24918, n24919, n24920, n24921, n24922, n24923,
    n24924, n24925, n24926, n24927, n24928, n24929,
    n24930, n24931, n24932, n24933, n24934, n24935,
    n24936, n24937, n24938, n24939, n24940, n24941,
    n24942, n24943, n24944, n24945, n24946, n24947,
    n24948, n24949, n24951, n24952, n24953, n24954,
    n24955, n24956, n24957, n24958, n24959, n24960,
    n24961, n24962, n24963, n24964, n24965, n24966,
    n24967, n24968, n24969, n24970, n24971, n24972,
    n24973, n24974, n24975, n24976, n24977, n24978,
    n24979, n24980, n24981, n24982, n24983, n24984,
    n24985, n24986, n24987, n24988, n24989, n24990,
    n24991, n24992, n24993, n24994, n24995, n24996,
    n24997, n24998, n24999, n25000, n25001, n25002,
    n25003, n25004, n25005, n25006, n25007, n25008,
    n25009, n25010, n25011, n25012, n25013, n25014,
    n25015, n25016, n25017, n25018, n25019, n25020,
    n25021, n25022, n25023, n25024, n25025, n25026,
    n25027, n25028, n25029, n25030, n25031, n25032,
    n25033, n25034, n25035, n25036, n25037, n25038,
    n25039, n25040, n25041, n25042, n25043, n25044,
    n25045, n25046, n25047, n25048, n25049, n25050,
    n25051, n25052, n25053, n25054, n25055, n25056,
    n25057, n25058, n25059, n25060, n25061, n25062,
    n25063, n25064, n25065, n25066, n25067, n25068,
    n25069, n25070, n25071, n25072, n25073, n25074,
    n25075, n25076, n25078, n25079, n25080, n25081,
    n25082, n25083, n25084, n25085, n25086, n25087,
    n25088, n25089, n25090, n25091, n25092, n25093,
    n25094, n25095, n25096, n25097, n25098, n25099,
    n25100, n25101, n25102, n25103, n25104, n25105,
    n25106, n25107, n25108, n25109, n25110, n25111,
    n25112, n25113, n25114, n25115, n25116, n25117,
    n25118, n25119, n25120, n25121, n25122, n25123,
    n25124, n25125, n25126, n25127, n25128, n25129,
    n25130, n25131, n25132, n25133, n25134, n25135,
    n25136, n25137, n25138, n25139, n25140, n25141,
    n25142, n25143, n25144, n25145, n25146, n25147,
    n25148, n25149, n25150, n25151, n25152, n25153,
    n25154, n25155, n25156, n25157, n25158, n25159,
    n25160, n25161, n25162, n25163, n25164, n25165,
    n25166, n25167, n25168, n25169, n25170, n25171,
    n25172, n25173, n25174, n25175, n25176, n25177,
    n25178, n25179, n25180, n25181, n25182, n25183,
    n25184, n25185, n25186, n25187, n25188, n25189,
    n25190, n25191, n25192, n25193, n25194, n25196,
    n25197, n25198, n25199, n25200, n25201, n25202,
    n25203, n25204, n25205, n25206, n25207, n25208,
    n25209, n25210, n25211, n25212, n25213, n25214,
    n25215, n25216, n25217, n25218, n25219, n25220,
    n25221, n25222, n25223, n25224, n25225, n25226,
    n25227, n25228, n25229, n25230, n25231, n25232,
    n25233, n25234, n25235, n25236, n25237, n25238,
    n25239, n25240, n25241, n25242, n25243, n25244,
    n25245, n25246, n25247, n25248, n25249, n25250,
    n25251, n25252, n25253, n25254, n25255, n25256,
    n25257, n25258, n25259, n25260, n25261, n25262,
    n25263, n25264, n25265, n25266, n25267, n25268,
    n25269, n25270, n25271, n25272, n25273, n25274,
    n25275, n25276, n25277, n25278, n25279, n25280,
    n25281, n25282, n25283, n25284, n25285, n25286,
    n25287, n25288, n25289, n25290, n25291, n25292,
    n25293, n25294, n25295, n25296, n25297, n25298,
    n25299, n25300, n25301, n25302, n25303, n25304,
    n25305, n25306, n25307, n25308, n25309, n25310,
    n25311, n25313, n25314, n25315, n25316, n25317,
    n25318, n25319, n25320, n25321, n25322, n25323,
    n25324, n25325, n25326, n25327, n25328, n25329,
    n25330, n25331, n25332, n25333, n25334, n25335,
    n25336, n25337, n25338, n25339, n25340, n25341,
    n25342, n25343, n25344, n25345, n25346, n25347,
    n25348, n25349, n25350, n25351, n25352, n25353,
    n25354, n25355, n25356, n25357, n25358, n25359,
    n25360, n25361, n25362, n25363, n25364, n25365,
    n25366, n25367, n25368, n25369, n25370, n25371,
    n25372, n25373, n25374, n25375, n25376, n25377,
    n25378, n25379, n25380, n25381, n25382, n25383,
    n25384, n25385, n25386, n25387, n25388, n25389,
    n25390, n25391, n25392, n25393, n25394, n25395,
    n25396, n25397, n25398, n25399, n25400, n25401,
    n25402, n25403, n25404, n25405, n25406, n25407,
    n25408, n25409, n25410, n25411, n25412, n25413,
    n25414, n25415, n25416, n25417, n25418, n25420,
    n25421, n25422, n25423, n25424, n25425, n25426,
    n25427, n25428, n25429, n25430, n25431, n25432,
    n25433, n25434, n25435, n25436, n25437, n25438,
    n25439, n25440, n25441, n25442, n25443, n25444,
    n25445, n25446, n25447, n25448, n25449, n25450,
    n25451, n25452, n25453, n25454, n25455, n25456,
    n25457, n25458, n25459, n25460, n25461, n25462,
    n25463, n25464, n25465, n25466, n25467, n25468,
    n25469, n25470, n25471, n25472, n25473, n25474,
    n25475, n25476, n25477, n25478, n25479, n25480,
    n25481, n25482, n25483, n25484, n25485, n25486,
    n25487, n25488, n25489, n25490, n25491, n25492,
    n25493, n25494, n25495, n25496, n25497, n25498,
    n25499, n25500, n25501, n25502, n25503, n25504,
    n25505, n25506, n25507, n25508, n25509, n25510,
    n25511, n25512, n25513, n25514, n25515, n25516,
    n25517, n25518, n25520, n25521, n25522, n25523,
    n25524, n25525, n25526, n25527, n25528, n25529,
    n25530, n25531, n25532, n25533, n25534, n25535,
    n25536, n25537, n25538, n25539, n25540, n25541,
    n25542, n25543, n25544, n25545, n25546, n25547,
    n25548, n25549, n25550, n25551, n25552, n25553,
    n25554, n25555, n25556, n25557, n25558, n25559,
    n25560, n25561, n25562, n25563, n25564, n25565,
    n25566, n25567, n25568, n25569, n25570, n25571,
    n25572, n25573, n25574, n25575, n25576, n25577,
    n25578, n25579, n25580, n25581, n25582, n25583,
    n25584, n25585, n25586, n25587, n25588, n25589,
    n25590, n25591, n25592, n25593, n25594, n25595,
    n25596, n25597, n25598, n25599, n25600, n25601,
    n25602, n25603, n25604, n25605, n25606, n25607,
    n25608, n25609, n25610, n25611, n25612, n25613,
    n25614, n25615, n25617, n25618, n25619, n25620,
    n25621, n25622, n25623, n25624, n25625, n25626,
    n25627, n25628, n25629, n25630, n25631, n25632,
    n25633, n25634, n25635, n25636, n25637, n25638,
    n25639, n25640, n25641, n25642, n25643, n25644,
    n25645, n25646, n25647, n25648, n25649, n25650,
    n25651, n25652, n25653, n25654, n25655, n25656,
    n25657, n25658, n25659, n25660, n25661, n25662,
    n25663, n25664, n25665, n25666, n25667, n25668,
    n25669, n25670, n25671, n25672, n25673, n25674,
    n25675, n25676, n25677, n25678, n25679, n25680,
    n25681, n25682, n25683, n25684, n25685, n25686,
    n25687, n25688, n25689, n25690, n25691, n25692,
    n25693, n25694, n25695, n25696, n25697, n25698,
    n25699, n25700, n25701, n25702, n25703, n25704,
    n25706, n25707, n25708, n25709, n25710, n25711,
    n25712, n25713, n25714, n25715, n25716, n25717,
    n25718, n25719, n25720, n25721, n25722, n25723,
    n25724, n25725, n25726, n25727, n25728, n25729,
    n25730, n25731, n25732, n25733, n25734, n25735,
    n25736, n25737, n25738, n25739, n25740, n25741,
    n25742, n25743, n25744, n25745, n25746, n25747,
    n25748, n25749, n25750, n25751, n25752, n25753,
    n25754, n25755, n25756, n25757, n25758, n25759,
    n25760, n25761, n25762, n25763, n25764, n25765,
    n25766, n25767, n25768, n25769, n25770, n25771,
    n25772, n25773, n25774, n25775, n25776, n25777,
    n25778, n25779, n25780, n25781, n25782, n25783,
    n25784, n25785, n25786, n25788, n25789, n25790,
    n25791, n25792, n25793, n25794, n25795, n25796,
    n25797, n25798, n25799, n25800, n25801, n25802,
    n25803, n25804, n25805, n25806, n25807, n25808,
    n25809, n25810, n25811, n25812, n25813, n25814,
    n25815, n25816, n25817, n25818, n25819, n25820,
    n25821, n25822, n25823, n25824, n25825, n25826,
    n25827, n25828, n25829, n25830, n25831, n25832,
    n25833, n25834, n25835, n25836, n25837, n25838,
    n25839, n25840, n25841, n25842, n25843, n25844,
    n25845, n25846, n25847, n25848, n25849, n25850,
    n25851, n25852, n25853, n25854, n25855, n25856,
    n25857, n25858, n25859, n25860, n25861, n25862,
    n25863, n25864, n25865, n25866, n25868, n25869,
    n25870, n25871, n25872, n25873, n25874, n25875,
    n25876, n25877, n25878, n25879, n25880, n25881,
    n25882, n25883, n25884, n25885, n25886, n25887,
    n25888, n25889, n25890, n25891, n25892, n25893,
    n25894, n25895, n25896, n25897, n25898, n25899,
    n25900, n25901, n25902, n25903, n25904, n25905,
    n25906, n25907, n25908, n25909, n25910, n25911,
    n25912, n25913, n25914, n25915, n25916, n25917,
    n25918, n25919, n25920, n25921, n25922, n25923,
    n25924, n25925, n25926, n25927, n25928, n25929,
    n25930, n25931, n25932, n25933, n25934, n25935,
    n25936, n25937, n25939, n25940, n25941, n25942,
    n25943, n25944, n25945, n25946, n25947, n25948,
    n25949, n25950, n25951, n25952, n25953, n25954,
    n25955, n25956, n25957, n25958, n25959, n25960,
    n25961, n25962, n25963, n25964, n25965, n25966,
    n25967, n25968, n25969, n25970, n25971, n25972,
    n25973, n25974, n25975, n25976, n25977, n25978,
    n25979, n25980, n25981, n25982, n25983, n25984,
    n25985, n25986, n25987, n25988, n25989, n25990,
    n25991, n25992, n25993, n25994, n25995, n25996,
    n25997, n25998, n25999, n26000, n26002, n26003,
    n26004, n26005, n26006, n26007, n26008, n26009,
    n26010, n26011, n26012, n26013, n26014, n26015,
    n26016, n26017, n26018, n26019, n26020, n26021,
    n26022, n26023, n26024, n26025, n26026, n26027,
    n26028, n26029, n26030, n26031, n26032, n26033,
    n26034, n26035, n26036, n26037, n26038, n26039,
    n26040, n26041, n26042, n26043, n26044, n26045,
    n26046, n26047, n26048, n26049, n26050, n26051,
    n26052, n26053, n26054, n26055, n26056, n26057,
    n26058, n26059, n26060, n26062, n26063, n26064,
    n26065, n26066, n26067, n26068, n26069, n26070,
    n26071, n26072, n26073, n26074, n26075, n26076,
    n26077, n26078, n26079, n26080, n26081, n26082,
    n26083, n26084, n26085, n26086, n26087, n26088,
    n26089, n26090, n26091, n26092, n26093, n26094,
    n26095, n26096, n26097, n26098, n26099, n26100,
    n26101, n26102, n26103, n26104, n26105, n26106,
    n26107, n26108, n26109, n26110, n26111, n26112,
    n26113, n26114, n26115, n26116, n26118, n26119,
    n26120, n26121, n26122, n26123, n26124, n26125,
    n26126, n26127, n26128, n26129, n26130, n26131,
    n26132, n26133, n26134, n26135, n26136, n26137,
    n26138, n26139, n26140, n26141, n26142, n26143,
    n26144, n26145, n26146, n26147, n26148, n26149,
    n26150, n26151, n26152, n26153, n26154, n26155,
    n26156, n26157, n26158, n26159, n26160, n26161,
    n26162, n26164, n26165, n26166, n26167, n26168,
    n26169, n26170, n26171, n26172, n26173, n26174,
    n26175, n26176, n26177, n26178, n26179, n26180,
    n26181, n26182, n26183, n26184, n26185, n26186,
    n26187, n26188, n26189, n26190, n26191, n26192,
    n26193, n26194, n26195, n26196, n26197, n26198,
    n26199, n26200, n26201, n26202, n26203, n26204,
    n26205, n26206, n26208, n26209, n26210, n26211,
    n26212, n26213, n26214, n26215, n26216, n26217,
    n26218, n26219, n26220, n26221, n26222, n26223,
    n26224, n26225, n26226, n26227, n26228, n26229,
    n26230, n26231, n26232, n26233, n26234, n26235,
    n26236, n26237, n26238, n26239, n26240, n26241,
    n26243, n26244, n26245, n26246, n26247, n26248,
    n26249, n26250, n26251, n26252, n26253, n26254,
    n26255, n26256, n26257, n26258, n26259, n26260,
    n26261, n26262, n26263, n26264, n26265, n26266,
    n26267, n26268, n26270, n26271, n26272, n26273,
    n26274, n26275, n26276, n26277, n26278, n26279,
    n26280, n26281, n26282, n26283, n26284, n26285,
    n26286, n26287, n26288, n26289, n26290, n26291,
    n26292, n26294, n26295, n26296, n26297, n26298,
    n26299, n26300, n26301, n26302, n26303, n26304,
    n26305, n26306, n26307, n26308, n26309, n26311,
    n26312, n26313, n26314, n26315, n26316, n26317,
    n26318;
  assign po0  = pi0  & pi64 ;
  assign n258 = pi2  & ~po0 ;
  assign n259 = ~pi0  & pi1 ;
  assign n260 = pi64  & n259;
  assign n261 = ~pi1  & pi2 ;
  assign n262 = pi1  & ~pi2 ;
  assign n263 = ~n261 & ~n262;
  assign n264 = pi0  & n263;
  assign n265 = pi65  & n264;
  assign n266 = ~n260 & ~n265;
  assign n267 = pi0  & ~n263;
  assign n268 = pi64  & pi65 ;
  assign n269 = ~pi64  & ~pi65 ;
  assign n270 = ~n268 & ~n269;
  assign n271 = n267 & n270;
  assign n272 = n266 & ~n271;
  assign n273 = pi2  & ~n272;
  assign n274 = pi2  & ~n273;
  assign n275 = ~n272 & ~n273;
  assign n276 = ~n274 & ~n275;
  assign n277 = n258 & ~n276;
  assign n278 = ~n258 & n276;
  assign po1  = ~n277 & ~n278;
  assign n280 = pi66  & n264;
  assign n281 = n261 & ~n267;
  assign n282 = pi64  & n281;
  assign n283 = pi65  & n259;
  assign n284 = ~n282 & ~n283;
  assign n285 = ~n280 & n284;
  assign n286 = pi65  & ~pi66 ;
  assign n287 = ~pi65  & pi66 ;
  assign n288 = ~n286 & ~n287;
  assign n289 = ~n268 & n288;
  assign n290 = pi64  & n286;
  assign n291 = ~n289 & ~n290;
  assign n292 = n267 & n291;
  assign n293 = n285 & ~n292;
  assign n294 = pi2  & ~n293;
  assign n295 = pi2  & ~n294;
  assign n296 = ~n293 & ~n294;
  assign n297 = ~n295 & ~n296;
  assign n298 = n277 & ~n297;
  assign n299 = ~n277 & n297;
  assign po2  = ~n298 & ~n299;
  assign n301 = pi67  & n264;
  assign n302 = pi65  & n281;
  assign n303 = pi66  & n259;
  assign n304 = ~n302 & ~n303;
  assign n305 = ~n301 & n304;
  assign n306 = pi65  & pi66 ;
  assign n307 = ~n290 & ~n306;
  assign n308 = ~pi66  & ~pi67 ;
  assign n309 = pi66  & pi67 ;
  assign n310 = ~n308 & ~n309;
  assign n311 = ~n307 & n310;
  assign n312 = n307 & ~n310;
  assign n313 = ~n311 & ~n312;
  assign n314 = n267 & n313;
  assign n315 = n305 & ~n314;
  assign n316 = pi2  & ~n315;
  assign n317 = pi2  & ~n316;
  assign n318 = ~n315 & ~n316;
  assign n319 = ~n317 & ~n318;
  assign n320 = pi2  & ~pi3 ;
  assign n321 = ~pi2  & pi3 ;
  assign n322 = ~n320 & ~n321;
  assign n323 = pi64  & ~n322;
  assign n324 = ~n319 & n323;
  assign n325 = n319 & ~n323;
  assign n326 = ~n324 & ~n325;
  assign n327 = n298 & n326;
  assign n328 = ~n298 & ~n326;
  assign po3  = ~n327 & ~n328;
  assign n330 = ~n324 & ~n327;
  assign n331 = pi5  & ~n323;
  assign n332 = ~pi3  & pi4 ;
  assign n333 = pi3  & ~pi4 ;
  assign n334 = ~n332 & ~n333;
  assign n335 = n322 & ~n334;
  assign n336 = pi64  & n335;
  assign n337 = ~pi4  & pi5 ;
  assign n338 = pi4  & ~pi5 ;
  assign n339 = ~n337 & ~n338;
  assign n340 = ~n322 & n339;
  assign n341 = pi65  & n340;
  assign n342 = ~n336 & ~n341;
  assign n343 = ~n322 & ~n339;
  assign n344 = n270 & n343;
  assign n345 = n342 & ~n344;
  assign n346 = pi5  & ~n345;
  assign n347 = pi5  & ~n346;
  assign n348 = ~n345 & ~n346;
  assign n349 = ~n347 & ~n348;
  assign n350 = n331 & ~n349;
  assign n351 = ~n331 & n349;
  assign n352 = ~n350 & ~n351;
  assign n353 = pi68  & n264;
  assign n354 = pi66  & n281;
  assign n355 = pi67  & n259;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n353 & n356;
  assign n358 = ~n309 & ~n311;
  assign n359 = ~pi67  & ~pi68 ;
  assign n360 = pi67  & pi68 ;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~n358 & n361;
  assign n363 = n358 & ~n361;
  assign n364 = ~n362 & ~n363;
  assign n365 = n267 & n364;
  assign n366 = n357 & ~n365;
  assign n367 = pi2  & ~n366;
  assign n368 = pi2  & ~n367;
  assign n369 = ~n366 & ~n367;
  assign n370 = ~n368 & ~n369;
  assign n371 = n352 & ~n370;
  assign n372 = ~n352 & n370;
  assign n373 = ~n371 & ~n372;
  assign n374 = ~n330 & n373;
  assign n375 = n330 & ~n373;
  assign po4  = ~n374 & ~n375;
  assign n377 = ~n371 & ~n374;
  assign n378 = pi66  & n340;
  assign n379 = n322 & ~n339;
  assign n380 = n334 & n379;
  assign n381 = pi64  & n380;
  assign n382 = pi65  & n335;
  assign n383 = ~n381 & ~n382;
  assign n384 = ~n378 & n383;
  assign n385 = ~n343 & n384;
  assign n386 = ~n291 & n384;
  assign n387 = ~n385 & ~n386;
  assign n388 = pi5  & ~n387;
  assign n389 = ~pi5  & n387;
  assign n390 = ~n388 & ~n389;
  assign n391 = n350 & ~n390;
  assign n392 = ~n350 & n390;
  assign n393 = ~n391 & ~n392;
  assign n394 = pi69  & n264;
  assign n395 = pi67  & n281;
  assign n396 = pi68  & n259;
  assign n397 = ~n395 & ~n396;
  assign n398 = ~n394 & n397;
  assign n399 = ~n360 & ~n362;
  assign n400 = ~pi68  & ~pi69 ;
  assign n401 = pi68  & pi69 ;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~n399 & n402;
  assign n404 = n399 & ~n402;
  assign n405 = ~n403 & ~n404;
  assign n406 = n267 & n405;
  assign n407 = n398 & ~n406;
  assign n408 = pi2  & ~n407;
  assign n409 = pi2  & ~n408;
  assign n410 = ~n407 & ~n408;
  assign n411 = ~n409 & ~n410;
  assign n412 = n393 & ~n411;
  assign n413 = ~n393 & n411;
  assign n414 = ~n412 & ~n413;
  assign n415 = ~n377 & n414;
  assign n416 = n377 & ~n414;
  assign po5  = ~n415 & ~n416;
  assign n418 = ~n412 & ~n415;
  assign n419 = pi70  & n264;
  assign n420 = pi68  & n281;
  assign n421 = pi69  & n259;
  assign n422 = ~n420 & ~n421;
  assign n423 = ~n419 & n422;
  assign n424 = ~n401 & ~n403;
  assign n425 = ~pi69  & ~pi70 ;
  assign n426 = pi69  & pi70 ;
  assign n427 = ~n425 & ~n426;
  assign n428 = ~n424 & n427;
  assign n429 = n424 & ~n427;
  assign n430 = ~n428 & ~n429;
  assign n431 = n267 & n430;
  assign n432 = n423 & ~n431;
  assign n433 = pi2  & ~n432;
  assign n434 = pi2  & ~n433;
  assign n435 = ~n432 & ~n433;
  assign n436 = ~n434 & ~n435;
  assign n437 = pi67  & n340;
  assign n438 = pi65  & n380;
  assign n439 = pi66  & n335;
  assign n440 = ~n438 & ~n439;
  assign n441 = ~n437 & n440;
  assign n442 = n313 & n343;
  assign n443 = n441 & ~n442;
  assign n444 = pi5  & ~n443;
  assign n445 = pi5  & ~n444;
  assign n446 = ~n443 & ~n444;
  assign n447 = ~n445 & ~n446;
  assign n448 = pi5  & ~pi6 ;
  assign n449 = ~pi5  & pi6 ;
  assign n450 = ~n448 & ~n449;
  assign n451 = pi64  & ~n450;
  assign n452 = n391 & n451;
  assign n453 = ~n391 & ~n451;
  assign n454 = ~n452 & ~n453;
  assign n455 = ~n447 & n454;
  assign n456 = n447 & ~n454;
  assign n457 = ~n455 & ~n456;
  assign n458 = ~n436 & n457;
  assign n459 = n436 & ~n457;
  assign n460 = ~n458 & ~n459;
  assign n461 = ~n418 & n460;
  assign n462 = n418 & ~n460;
  assign po6  = ~n461 & ~n462;
  assign n464 = ~n458 & ~n461;
  assign n465 = pi71  & n264;
  assign n466 = pi69  & n281;
  assign n467 = pi70  & n259;
  assign n468 = ~n466 & ~n467;
  assign n469 = ~n465 & n468;
  assign n470 = ~n426 & ~n428;
  assign n471 = ~pi70  & ~pi71 ;
  assign n472 = pi70  & pi71 ;
  assign n473 = ~n471 & ~n472;
  assign n474 = ~n470 & n473;
  assign n475 = n470 & ~n473;
  assign n476 = ~n474 & ~n475;
  assign n477 = n267 & n476;
  assign n478 = n469 & ~n477;
  assign n479 = pi2  & ~n478;
  assign n480 = pi2  & ~n479;
  assign n481 = ~n478 & ~n479;
  assign n482 = ~n480 & ~n481;
  assign n483 = ~n452 & ~n455;
  assign n484 = pi8  & ~n451;
  assign n485 = ~pi6  & pi7 ;
  assign n486 = pi6  & ~pi7 ;
  assign n487 = ~n485 & ~n486;
  assign n488 = n450 & ~n487;
  assign n489 = pi64  & n488;
  assign n490 = ~pi7  & pi8 ;
  assign n491 = pi7  & ~pi8 ;
  assign n492 = ~n490 & ~n491;
  assign n493 = ~n450 & n492;
  assign n494 = pi65  & n493;
  assign n495 = ~n489 & ~n494;
  assign n496 = ~n450 & ~n492;
  assign n497 = n270 & n496;
  assign n498 = n495 & ~n497;
  assign n499 = pi8  & ~n498;
  assign n500 = pi8  & ~n499;
  assign n501 = ~n498 & ~n499;
  assign n502 = ~n500 & ~n501;
  assign n503 = n484 & ~n502;
  assign n504 = ~n484 & n502;
  assign n505 = ~n503 & ~n504;
  assign n506 = pi68  & n340;
  assign n507 = pi66  & n380;
  assign n508 = pi67  & n335;
  assign n509 = ~n507 & ~n508;
  assign n510 = ~n506 & n509;
  assign n511 = n343 & n364;
  assign n512 = n510 & ~n511;
  assign n513 = pi5  & ~n512;
  assign n514 = pi5  & ~n513;
  assign n515 = ~n512 & ~n513;
  assign n516 = ~n514 & ~n515;
  assign n517 = n505 & ~n516;
  assign n518 = ~n505 & n516;
  assign n519 = ~n517 & ~n518;
  assign n520 = ~n483 & n519;
  assign n521 = n483 & ~n519;
  assign n522 = ~n520 & ~n521;
  assign n523 = ~n482 & n522;
  assign n524 = n482 & ~n522;
  assign n525 = ~n523 & ~n524;
  assign n526 = ~n464 & n525;
  assign n527 = n464 & ~n525;
  assign po7  = ~n526 & ~n527;
  assign n529 = ~n523 & ~n526;
  assign n530 = ~n517 & ~n520;
  assign n531 = pi66  & n493;
  assign n532 = n450 & ~n492;
  assign n533 = n487 & n532;
  assign n534 = pi64  & n533;
  assign n535 = pi65  & n488;
  assign n536 = ~n534 & ~n535;
  assign n537 = ~n531 & n536;
  assign n538 = n291 & n496;
  assign n539 = n537 & ~n538;
  assign n540 = pi8  & ~n539;
  assign n541 = pi8  & ~n540;
  assign n542 = ~n539 & ~n540;
  assign n543 = ~n541 & ~n542;
  assign n544 = ~n503 & n543;
  assign n545 = n503 & ~n543;
  assign n546 = ~n544 & ~n545;
  assign n547 = pi69  & n340;
  assign n548 = pi67  & n380;
  assign n549 = pi68  & n335;
  assign n550 = ~n548 & ~n549;
  assign n551 = ~n547 & n550;
  assign n552 = n343 & n405;
  assign n553 = n551 & ~n552;
  assign n554 = pi5  & ~n553;
  assign n555 = pi5  & ~n554;
  assign n556 = ~n553 & ~n554;
  assign n557 = ~n555 & ~n556;
  assign n558 = n546 & ~n557;
  assign n559 = ~n546 & n557;
  assign n560 = ~n558 & ~n559;
  assign n561 = n530 & ~n560;
  assign n562 = ~n530 & n560;
  assign n563 = ~n561 & ~n562;
  assign n564 = pi72  & n264;
  assign n565 = pi70  & n281;
  assign n566 = pi71  & n259;
  assign n567 = ~n565 & ~n566;
  assign n568 = ~n564 & n567;
  assign n569 = ~n472 & ~n474;
  assign n570 = ~pi71  & ~pi72 ;
  assign n571 = pi71  & pi72 ;
  assign n572 = ~n570 & ~n571;
  assign n573 = ~n569 & n572;
  assign n574 = n569 & ~n572;
  assign n575 = ~n573 & ~n574;
  assign n576 = n267 & n575;
  assign n577 = n568 & ~n576;
  assign n578 = pi2  & ~n577;
  assign n579 = pi2  & ~n578;
  assign n580 = ~n577 & ~n578;
  assign n581 = ~n579 & ~n580;
  assign n582 = n563 & ~n581;
  assign n583 = ~n563 & n581;
  assign n584 = ~n582 & ~n583;
  assign n585 = ~n529 & n584;
  assign n586 = n529 & ~n584;
  assign po8  = ~n585 & ~n586;
  assign n588 = ~n582 & ~n585;
  assign n589 = ~n558 & ~n562;
  assign n590 = pi67  & n493;
  assign n591 = pi65  & n533;
  assign n592 = pi66  & n488;
  assign n593 = ~n591 & ~n592;
  assign n594 = ~n590 & n593;
  assign n595 = n313 & n496;
  assign n596 = n594 & ~n595;
  assign n597 = pi8  & ~n596;
  assign n598 = pi8  & ~n597;
  assign n599 = ~n596 & ~n597;
  assign n600 = ~n598 & ~n599;
  assign n601 = pi8  & ~pi9 ;
  assign n602 = ~pi8  & pi9 ;
  assign n603 = ~n601 & ~n602;
  assign n604 = pi64  & ~n603;
  assign n605 = n545 & n604;
  assign n606 = ~n545 & ~n604;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~n600 & n607;
  assign n609 = n600 & ~n607;
  assign n610 = ~n608 & ~n609;
  assign n611 = pi70  & n340;
  assign n612 = pi68  & n380;
  assign n613 = pi69  & n335;
  assign n614 = ~n612 & ~n613;
  assign n615 = ~n611 & n614;
  assign n616 = n343 & n430;
  assign n617 = n615 & ~n616;
  assign n618 = pi5  & ~n617;
  assign n619 = pi5  & ~n618;
  assign n620 = ~n617 & ~n618;
  assign n621 = ~n619 & ~n620;
  assign n622 = n610 & ~n621;
  assign n623 = ~n610 & n621;
  assign n624 = ~n622 & ~n623;
  assign n625 = n589 & ~n624;
  assign n626 = ~n589 & n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = pi73  & n264;
  assign n629 = pi71  & n281;
  assign n630 = pi72  & n259;
  assign n631 = ~n629 & ~n630;
  assign n632 = ~n628 & n631;
  assign n633 = ~n571 & ~n573;
  assign n634 = ~pi72  & ~pi73 ;
  assign n635 = pi72  & pi73 ;
  assign n636 = ~n634 & ~n635;
  assign n637 = ~n633 & n636;
  assign n638 = n633 & ~n636;
  assign n639 = ~n637 & ~n638;
  assign n640 = n267 & n639;
  assign n641 = n632 & ~n640;
  assign n642 = pi2  & ~n641;
  assign n643 = pi2  & ~n642;
  assign n644 = ~n641 & ~n642;
  assign n645 = ~n643 & ~n644;
  assign n646 = n627 & ~n645;
  assign n647 = ~n627 & n645;
  assign n648 = ~n646 & ~n647;
  assign n649 = ~n588 & n648;
  assign n650 = n588 & ~n648;
  assign po9  = ~n649 & ~n650;
  assign n652 = ~n646 & ~n649;
  assign n653 = ~n622 & ~n626;
  assign n654 = ~n605 & ~n608;
  assign n655 = pi68  & n493;
  assign n656 = pi66  & n533;
  assign n657 = pi67  & n488;
  assign n658 = ~n656 & ~n657;
  assign n659 = ~n655 & n658;
  assign n660 = n364 & n496;
  assign n661 = n659 & ~n660;
  assign n662 = pi8  & ~n661;
  assign n663 = pi8  & ~n662;
  assign n664 = ~n661 & ~n662;
  assign n665 = ~n663 & ~n664;
  assign n666 = pi11  & ~n604;
  assign n667 = ~pi9  & pi10 ;
  assign n668 = pi9  & ~pi10 ;
  assign n669 = ~n667 & ~n668;
  assign n670 = n603 & ~n669;
  assign n671 = pi64  & n670;
  assign n672 = ~pi10  & pi11 ;
  assign n673 = pi10  & ~pi11 ;
  assign n674 = ~n672 & ~n673;
  assign n675 = ~n603 & n674;
  assign n676 = pi65  & n675;
  assign n677 = ~n671 & ~n676;
  assign n678 = ~n603 & ~n674;
  assign n679 = n270 & n678;
  assign n680 = n677 & ~n679;
  assign n681 = pi11  & ~n680;
  assign n682 = pi11  & ~n681;
  assign n683 = ~n680 & ~n681;
  assign n684 = ~n682 & ~n683;
  assign n685 = n666 & ~n684;
  assign n686 = ~n666 & n684;
  assign n687 = ~n685 & ~n686;
  assign n688 = n665 & ~n687;
  assign n689 = ~n665 & n687;
  assign n690 = ~n688 & ~n689;
  assign n691 = ~n654 & n690;
  assign n692 = n654 & ~n690;
  assign n693 = ~n691 & ~n692;
  assign n694 = pi71  & n340;
  assign n695 = pi69  & n380;
  assign n696 = pi70  & n335;
  assign n697 = ~n695 & ~n696;
  assign n698 = ~n694 & n697;
  assign n699 = n343 & n476;
  assign n700 = n698 & ~n699;
  assign n701 = pi5  & ~n700;
  assign n702 = pi5  & ~n701;
  assign n703 = ~n700 & ~n701;
  assign n704 = ~n702 & ~n703;
  assign n705 = n693 & ~n704;
  assign n706 = ~n693 & n704;
  assign n707 = ~n705 & ~n706;
  assign n708 = n653 & ~n707;
  assign n709 = ~n653 & n707;
  assign n710 = ~n708 & ~n709;
  assign n711 = pi74  & n264;
  assign n712 = pi72  & n281;
  assign n713 = pi73  & n259;
  assign n714 = ~n712 & ~n713;
  assign n715 = ~n711 & n714;
  assign n716 = ~n635 & ~n637;
  assign n717 = ~pi73  & ~pi74 ;
  assign n718 = pi73  & pi74 ;
  assign n719 = ~n717 & ~n718;
  assign n720 = ~n716 & n719;
  assign n721 = n716 & ~n719;
  assign n722 = ~n720 & ~n721;
  assign n723 = n267 & n722;
  assign n724 = n715 & ~n723;
  assign n725 = pi2  & ~n724;
  assign n726 = pi2  & ~n725;
  assign n727 = ~n724 & ~n725;
  assign n728 = ~n726 & ~n727;
  assign n729 = ~n710 & n728;
  assign n730 = n710 & ~n728;
  assign n731 = ~n729 & ~n730;
  assign n732 = ~n652 & n731;
  assign n733 = n652 & ~n731;
  assign po10  = ~n732 & ~n733;
  assign n735 = ~n730 & ~n732;
  assign n736 = pi75  & n264;
  assign n737 = pi73  & n281;
  assign n738 = pi74  & n259;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~n736 & n739;
  assign n741 = ~n718 & ~n720;
  assign n742 = ~pi74  & ~pi75 ;
  assign n743 = pi74  & pi75 ;
  assign n744 = ~n742 & ~n743;
  assign n745 = ~n741 & n744;
  assign n746 = n741 & ~n744;
  assign n747 = ~n745 & ~n746;
  assign n748 = n267 & n747;
  assign n749 = n740 & ~n748;
  assign n750 = pi2  & ~n749;
  assign n751 = pi2  & ~n750;
  assign n752 = ~n749 & ~n750;
  assign n753 = ~n751 & ~n752;
  assign n754 = ~n705 & ~n709;
  assign n755 = pi72  & n340;
  assign n756 = pi70  & n380;
  assign n757 = pi71  & n335;
  assign n758 = ~n756 & ~n757;
  assign n759 = ~n755 & n758;
  assign n760 = n343 & n575;
  assign n761 = n759 & ~n760;
  assign n762 = pi5  & ~n761;
  assign n763 = pi5  & ~n762;
  assign n764 = ~n761 & ~n762;
  assign n765 = ~n763 & ~n764;
  assign n766 = ~n689 & ~n691;
  assign n767 = pi66  & n675;
  assign n768 = n603 & ~n674;
  assign n769 = n669 & n768;
  assign n770 = pi64  & n769;
  assign n771 = pi65  & n670;
  assign n772 = ~n770 & ~n771;
  assign n773 = ~n767 & n772;
  assign n774 = n291 & n678;
  assign n775 = n773 & ~n774;
  assign n776 = pi11  & ~n775;
  assign n777 = pi11  & ~n776;
  assign n778 = ~n775 & ~n776;
  assign n779 = ~n777 & ~n778;
  assign n780 = ~n685 & n779;
  assign n781 = n685 & ~n779;
  assign n782 = ~n780 & ~n781;
  assign n783 = pi69  & n493;
  assign n784 = pi67  & n533;
  assign n785 = pi68  & n488;
  assign n786 = ~n784 & ~n785;
  assign n787 = ~n783 & n786;
  assign n788 = n405 & n496;
  assign n789 = n787 & ~n788;
  assign n790 = pi8  & ~n789;
  assign n791 = pi8  & ~n790;
  assign n792 = ~n789 & ~n790;
  assign n793 = ~n791 & ~n792;
  assign n794 = n782 & ~n793;
  assign n795 = ~n782 & n793;
  assign n796 = ~n794 & ~n795;
  assign n797 = ~n766 & n796;
  assign n798 = n766 & ~n796;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~n765 & n799;
  assign n801 = n765 & ~n799;
  assign n802 = ~n800 & ~n801;
  assign n803 = ~n754 & n802;
  assign n804 = n754 & ~n802;
  assign n805 = ~n803 & ~n804;
  assign n806 = ~n753 & n805;
  assign n807 = n753 & ~n805;
  assign n808 = ~n806 & ~n807;
  assign n809 = ~n735 & n808;
  assign n810 = n735 & ~n808;
  assign po11  = ~n809 & ~n810;
  assign n812 = ~n806 & ~n809;
  assign n813 = ~n794 & ~n797;
  assign n814 = pi67  & n675;
  assign n815 = pi65  & n769;
  assign n816 = pi66  & n670;
  assign n817 = ~n815 & ~n816;
  assign n818 = ~n814 & n817;
  assign n819 = n313 & n678;
  assign n820 = n818 & ~n819;
  assign n821 = pi11  & ~n820;
  assign n822 = pi11  & ~n821;
  assign n823 = ~n820 & ~n821;
  assign n824 = ~n822 & ~n823;
  assign n825 = pi11  & ~pi12 ;
  assign n826 = ~pi11  & pi12 ;
  assign n827 = ~n825 & ~n826;
  assign n828 = pi64  & ~n827;
  assign n829 = n781 & n828;
  assign n830 = ~n781 & ~n828;
  assign n831 = ~n829 & ~n830;
  assign n832 = ~n824 & n831;
  assign n833 = n824 & ~n831;
  assign n834 = ~n832 & ~n833;
  assign n835 = pi70  & n493;
  assign n836 = pi68  & n533;
  assign n837 = pi69  & n488;
  assign n838 = ~n836 & ~n837;
  assign n839 = ~n835 & n838;
  assign n840 = n430 & n496;
  assign n841 = n839 & ~n840;
  assign n842 = pi8  & ~n841;
  assign n843 = pi8  & ~n842;
  assign n844 = ~n841 & ~n842;
  assign n845 = ~n843 & ~n844;
  assign n846 = n834 & ~n845;
  assign n847 = ~n834 & n845;
  assign n848 = ~n846 & ~n847;
  assign n849 = n813 & ~n848;
  assign n850 = ~n813 & n848;
  assign n851 = ~n849 & ~n850;
  assign n852 = pi73  & n340;
  assign n853 = pi71  & n380;
  assign n854 = pi72  & n335;
  assign n855 = ~n853 & ~n854;
  assign n856 = ~n852 & n855;
  assign n857 = n343 & n639;
  assign n858 = n856 & ~n857;
  assign n859 = pi5  & ~n858;
  assign n860 = pi5  & ~n859;
  assign n861 = ~n858 & ~n859;
  assign n862 = ~n860 & ~n861;
  assign n863 = ~n851 & n862;
  assign n864 = n851 & ~n862;
  assign n865 = ~n863 & ~n864;
  assign n866 = ~n800 & ~n803;
  assign n867 = n865 & ~n866;
  assign n868 = ~n865 & n866;
  assign n869 = ~n867 & ~n868;
  assign n870 = pi76  & n264;
  assign n871 = pi74  & n281;
  assign n872 = pi75  & n259;
  assign n873 = ~n871 & ~n872;
  assign n874 = ~n870 & n873;
  assign n875 = ~n743 & ~n745;
  assign n876 = ~pi75  & ~pi76 ;
  assign n877 = pi75  & pi76 ;
  assign n878 = ~n876 & ~n877;
  assign n879 = ~n875 & n878;
  assign n880 = n875 & ~n878;
  assign n881 = ~n879 & ~n880;
  assign n882 = n267 & n881;
  assign n883 = n874 & ~n882;
  assign n884 = pi2  & ~n883;
  assign n885 = pi2  & ~n884;
  assign n886 = ~n883 & ~n884;
  assign n887 = ~n885 & ~n886;
  assign n888 = n869 & ~n887;
  assign n889 = ~n869 & n887;
  assign n890 = ~n888 & ~n889;
  assign n891 = ~n812 & n890;
  assign n892 = n812 & ~n890;
  assign po12  = ~n891 & ~n892;
  assign n894 = ~n888 & ~n891;
  assign n895 = ~n864 & ~n867;
  assign n896 = ~n846 & ~n850;
  assign n897 = ~n829 & ~n832;
  assign n898 = pi68  & n675;
  assign n899 = pi66  & n769;
  assign n900 = pi67  & n670;
  assign n901 = ~n899 & ~n900;
  assign n902 = ~n898 & n901;
  assign n903 = n364 & n678;
  assign n904 = n902 & ~n903;
  assign n905 = pi11  & ~n904;
  assign n906 = pi11  & ~n905;
  assign n907 = ~n904 & ~n905;
  assign n908 = ~n906 & ~n907;
  assign n909 = pi14  & ~n828;
  assign n910 = ~pi12  & pi13 ;
  assign n911 = pi12  & ~pi13 ;
  assign n912 = ~n910 & ~n911;
  assign n913 = n827 & ~n912;
  assign n914 = pi64  & n913;
  assign n915 = ~pi13  & pi14 ;
  assign n916 = pi13  & ~pi14 ;
  assign n917 = ~n915 & ~n916;
  assign n918 = ~n827 & n917;
  assign n919 = pi65  & n918;
  assign n920 = ~n914 & ~n919;
  assign n921 = ~n827 & ~n917;
  assign n922 = n270 & n921;
  assign n923 = n920 & ~n922;
  assign n924 = pi14  & ~n923;
  assign n925 = pi14  & ~n924;
  assign n926 = ~n923 & ~n924;
  assign n927 = ~n925 & ~n926;
  assign n928 = n909 & ~n927;
  assign n929 = ~n909 & n927;
  assign n930 = ~n928 & ~n929;
  assign n931 = n908 & ~n930;
  assign n932 = ~n908 & n930;
  assign n933 = ~n931 & ~n932;
  assign n934 = ~n897 & n933;
  assign n935 = n897 & ~n933;
  assign n936 = ~n934 & ~n935;
  assign n937 = pi71  & n493;
  assign n938 = pi69  & n533;
  assign n939 = pi70  & n488;
  assign n940 = ~n938 & ~n939;
  assign n941 = ~n937 & n940;
  assign n942 = n476 & n496;
  assign n943 = n941 & ~n942;
  assign n944 = pi8  & ~n943;
  assign n945 = pi8  & ~n944;
  assign n946 = ~n943 & ~n944;
  assign n947 = ~n945 & ~n946;
  assign n948 = n936 & ~n947;
  assign n949 = ~n936 & n947;
  assign n950 = ~n948 & ~n949;
  assign n951 = n896 & ~n950;
  assign n952 = ~n896 & n950;
  assign n953 = ~n951 & ~n952;
  assign n954 = pi74  & n340;
  assign n955 = pi72  & n380;
  assign n956 = pi73  & n335;
  assign n957 = ~n955 & ~n956;
  assign n958 = ~n954 & n957;
  assign n959 = n343 & n722;
  assign n960 = n958 & ~n959;
  assign n961 = pi5  & ~n960;
  assign n962 = pi5  & ~n961;
  assign n963 = ~n960 & ~n961;
  assign n964 = ~n962 & ~n963;
  assign n965 = n953 & ~n964;
  assign n966 = ~n953 & n964;
  assign n967 = ~n895 & ~n966;
  assign n968 = ~n965 & n967;
  assign n969 = ~n895 & ~n968;
  assign n970 = ~n965 & ~n968;
  assign n971 = ~n966 & n970;
  assign n972 = ~n969 & ~n971;
  assign n973 = pi77  & n264;
  assign n974 = pi75  & n281;
  assign n975 = pi76  & n259;
  assign n976 = ~n974 & ~n975;
  assign n977 = ~n973 & n976;
  assign n978 = ~n877 & ~n879;
  assign n979 = ~pi76  & ~pi77 ;
  assign n980 = pi76  & pi77 ;
  assign n981 = ~n979 & ~n980;
  assign n982 = ~n978 & n981;
  assign n983 = n978 & ~n981;
  assign n984 = ~n982 & ~n983;
  assign n985 = n267 & n984;
  assign n986 = n977 & ~n985;
  assign n987 = pi2  & ~n986;
  assign n988 = pi2  & ~n987;
  assign n989 = ~n986 & ~n987;
  assign n990 = ~n988 & ~n989;
  assign n991 = ~n972 & ~n990;
  assign n992 = n972 & n990;
  assign n993 = ~n991 & ~n992;
  assign n994 = ~n894 & n993;
  assign n995 = n894 & ~n993;
  assign po13  = ~n994 & ~n995;
  assign n997 = ~n991 & ~n994;
  assign n998 = pi78  & n264;
  assign n999 = pi76  & n281;
  assign n1000 = pi77  & n259;
  assign n1001 = ~n999 & ~n1000;
  assign n1002 = ~n998 & n1001;
  assign n1003 = ~n980 & ~n982;
  assign n1004 = ~pi77  & ~pi78 ;
  assign n1005 = pi77  & pi78 ;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~n1003 & n1006;
  assign n1008 = n1003 & ~n1006;
  assign n1009 = ~n1007 & ~n1008;
  assign n1010 = n267 & n1009;
  assign n1011 = n1002 & ~n1010;
  assign n1012 = pi2  & ~n1011;
  assign n1013 = pi2  & ~n1012;
  assign n1014 = ~n1011 & ~n1012;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = pi75  & n340;
  assign n1017 = pi73  & n380;
  assign n1018 = pi74  & n335;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = ~n1016 & n1019;
  assign n1021 = n343 & n747;
  assign n1022 = n1020 & ~n1021;
  assign n1023 = pi5  & ~n1022;
  assign n1024 = pi5  & ~n1023;
  assign n1025 = ~n1022 & ~n1023;
  assign n1026 = ~n1024 & ~n1025;
  assign n1027 = ~n948 & ~n952;
  assign n1028 = ~n932 & ~n934;
  assign n1029 = pi66  & n918;
  assign n1030 = n827 & ~n917;
  assign n1031 = n912 & n1030;
  assign n1032 = pi64  & n1031;
  assign n1033 = pi65  & n913;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = ~n1029 & n1034;
  assign n1036 = n291 & n921;
  assign n1037 = n1035 & ~n1036;
  assign n1038 = pi14  & ~n1037;
  assign n1039 = pi14  & ~n1038;
  assign n1040 = ~n1037 & ~n1038;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = ~n928 & n1041;
  assign n1043 = n928 & ~n1041;
  assign n1044 = ~n1042 & ~n1043;
  assign n1045 = pi69  & n675;
  assign n1046 = pi67  & n769;
  assign n1047 = pi68  & n670;
  assign n1048 = ~n1046 & ~n1047;
  assign n1049 = ~n1045 & n1048;
  assign n1050 = n405 & n678;
  assign n1051 = n1049 & ~n1050;
  assign n1052 = pi11  & ~n1051;
  assign n1053 = pi11  & ~n1052;
  assign n1054 = ~n1051 & ~n1052;
  assign n1055 = ~n1053 & ~n1054;
  assign n1056 = n1044 & ~n1055;
  assign n1057 = ~n1044 & n1055;
  assign n1058 = ~n1028 & ~n1057;
  assign n1059 = ~n1056 & n1058;
  assign n1060 = ~n1028 & ~n1059;
  assign n1061 = ~n1056 & ~n1059;
  assign n1062 = ~n1057 & n1061;
  assign n1063 = ~n1060 & ~n1062;
  assign n1064 = pi72  & n493;
  assign n1065 = pi70  & n533;
  assign n1066 = pi71  & n488;
  assign n1067 = ~n1065 & ~n1066;
  assign n1068 = ~n1064 & n1067;
  assign n1069 = n496 & n575;
  assign n1070 = n1068 & ~n1069;
  assign n1071 = pi8  & ~n1070;
  assign n1072 = pi8  & ~n1071;
  assign n1073 = ~n1070 & ~n1071;
  assign n1074 = ~n1072 & ~n1073;
  assign n1075 = n1063 & n1074;
  assign n1076 = ~n1063 & ~n1074;
  assign n1077 = ~n1075 & ~n1076;
  assign n1078 = ~n1027 & n1077;
  assign n1079 = n1027 & ~n1077;
  assign n1080 = ~n1078 & ~n1079;
  assign n1081 = n1026 & ~n1080;
  assign n1082 = ~n1026 & n1080;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~n970 & n1083;
  assign n1085 = n970 & ~n1083;
  assign n1086 = ~n1084 & ~n1085;
  assign n1087 = ~n1015 & n1086;
  assign n1088 = n1015 & ~n1086;
  assign n1089 = ~n1087 & ~n1088;
  assign n1090 = ~n997 & n1089;
  assign n1091 = n997 & ~n1089;
  assign po14  = ~n1090 & ~n1091;
  assign n1093 = ~n1087 & ~n1090;
  assign n1094 = pi79  & n264;
  assign n1095 = pi77  & n281;
  assign n1096 = pi78  & n259;
  assign n1097 = ~n1095 & ~n1096;
  assign n1098 = ~n1094 & n1097;
  assign n1099 = ~n1005 & ~n1007;
  assign n1100 = ~pi78  & ~pi79 ;
  assign n1101 = pi78  & pi79 ;
  assign n1102 = ~n1100 & ~n1101;
  assign n1103 = ~n1099 & n1102;
  assign n1104 = n1099 & ~n1102;
  assign n1105 = ~n1103 & ~n1104;
  assign n1106 = n267 & n1105;
  assign n1107 = n1098 & ~n1106;
  assign n1108 = pi2  & ~n1107;
  assign n1109 = pi2  & ~n1108;
  assign n1110 = ~n1107 & ~n1108;
  assign n1111 = ~n1109 & ~n1110;
  assign n1112 = ~n1082 & ~n1084;
  assign n1113 = pi76  & n340;
  assign n1114 = pi74  & n380;
  assign n1115 = pi75  & n335;
  assign n1116 = ~n1114 & ~n1115;
  assign n1117 = ~n1113 & n1116;
  assign n1118 = n343 & n881;
  assign n1119 = n1117 & ~n1118;
  assign n1120 = pi5  & ~n1119;
  assign n1121 = pi5  & ~n1120;
  assign n1122 = ~n1119 & ~n1120;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = ~n1076 & ~n1078;
  assign n1125 = pi73  & n493;
  assign n1126 = pi71  & n533;
  assign n1127 = pi72  & n488;
  assign n1128 = ~n1126 & ~n1127;
  assign n1129 = ~n1125 & n1128;
  assign n1130 = n496 & n639;
  assign n1131 = n1129 & ~n1130;
  assign n1132 = pi8  & ~n1131;
  assign n1133 = pi8  & ~n1132;
  assign n1134 = ~n1131 & ~n1132;
  assign n1135 = ~n1133 & ~n1134;
  assign n1136 = pi67  & n918;
  assign n1137 = pi65  & n1031;
  assign n1138 = pi66  & n913;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = ~n1136 & n1139;
  assign n1141 = n313 & n921;
  assign n1142 = n1140 & ~n1141;
  assign n1143 = pi14  & ~n1142;
  assign n1144 = pi14  & ~n1143;
  assign n1145 = ~n1142 & ~n1143;
  assign n1146 = ~n1144 & ~n1145;
  assign n1147 = pi14  & ~pi15 ;
  assign n1148 = ~pi14  & pi15 ;
  assign n1149 = ~n1147 & ~n1148;
  assign n1150 = pi64  & ~n1149;
  assign n1151 = n1043 & n1150;
  assign n1152 = ~n1043 & ~n1150;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~n1146 & n1153;
  assign n1155 = n1146 & ~n1153;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = pi70  & n675;
  assign n1158 = pi68  & n769;
  assign n1159 = pi69  & n670;
  assign n1160 = ~n1158 & ~n1159;
  assign n1161 = ~n1157 & n1160;
  assign n1162 = n430 & n678;
  assign n1163 = n1161 & ~n1162;
  assign n1164 = pi11  & ~n1163;
  assign n1165 = pi11  & ~n1164;
  assign n1166 = ~n1163 & ~n1164;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = n1156 & ~n1167;
  assign n1169 = ~n1156 & n1167;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = ~n1061 & n1170;
  assign n1172 = n1061 & ~n1170;
  assign n1173 = ~n1171 & ~n1172;
  assign n1174 = ~n1135 & n1173;
  assign n1175 = n1135 & ~n1173;
  assign n1176 = ~n1174 & ~n1175;
  assign n1177 = ~n1124 & n1176;
  assign n1178 = n1124 & ~n1176;
  assign n1179 = ~n1177 & ~n1178;
  assign n1180 = ~n1123 & n1179;
  assign n1181 = n1123 & ~n1179;
  assign n1182 = ~n1180 & ~n1181;
  assign n1183 = ~n1112 & n1182;
  assign n1184 = n1112 & ~n1182;
  assign n1185 = ~n1183 & ~n1184;
  assign n1186 = ~n1111 & n1185;
  assign n1187 = ~n1111 & ~n1186;
  assign n1188 = n1185 & ~n1186;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1093 & ~n1189;
  assign n1191 = n1093 & n1189;
  assign po15  = ~n1190 & ~n1191;
  assign n1193 = ~n1186 & ~n1190;
  assign n1194 = pi80  & n264;
  assign n1195 = pi78  & n281;
  assign n1196 = pi79  & n259;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = ~n1194 & n1197;
  assign n1199 = ~n1101 & ~n1103;
  assign n1200 = ~pi79  & ~pi80 ;
  assign n1201 = pi79  & pi80 ;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = ~n1199 & n1202;
  assign n1204 = n1199 & ~n1202;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = n267 & n1205;
  assign n1207 = n1198 & ~n1206;
  assign n1208 = pi2  & ~n1207;
  assign n1209 = pi2  & ~n1208;
  assign n1210 = ~n1207 & ~n1208;
  assign n1211 = ~n1209 & ~n1210;
  assign n1212 = ~n1180 & ~n1183;
  assign n1213 = pi77  & n340;
  assign n1214 = pi75  & n380;
  assign n1215 = pi76  & n335;
  assign n1216 = ~n1214 & ~n1215;
  assign n1217 = ~n1213 & n1216;
  assign n1218 = n343 & n984;
  assign n1219 = n1217 & ~n1218;
  assign n1220 = pi5  & ~n1219;
  assign n1221 = pi5  & ~n1220;
  assign n1222 = ~n1219 & ~n1220;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~n1174 & ~n1177;
  assign n1225 = pi74  & n493;
  assign n1226 = pi72  & n533;
  assign n1227 = pi73  & n488;
  assign n1228 = ~n1226 & ~n1227;
  assign n1229 = ~n1225 & n1228;
  assign n1230 = n496 & n722;
  assign n1231 = n1229 & ~n1230;
  assign n1232 = pi8  & ~n1231;
  assign n1233 = pi8  & ~n1232;
  assign n1234 = ~n1231 & ~n1232;
  assign n1235 = ~n1233 & ~n1234;
  assign n1236 = ~n1168 & ~n1171;
  assign n1237 = pi71  & n675;
  assign n1238 = pi69  & n769;
  assign n1239 = pi70  & n670;
  assign n1240 = ~n1238 & ~n1239;
  assign n1241 = ~n1237 & n1240;
  assign n1242 = n476 & n678;
  assign n1243 = n1241 & ~n1242;
  assign n1244 = pi11  & ~n1243;
  assign n1245 = pi11  & ~n1244;
  assign n1246 = ~n1243 & ~n1244;
  assign n1247 = ~n1245 & ~n1246;
  assign n1248 = ~n1151 & ~n1154;
  assign n1249 = pi68  & n918;
  assign n1250 = pi66  & n1031;
  assign n1251 = pi67  & n913;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = ~n1249 & n1252;
  assign n1254 = n364 & n921;
  assign n1255 = n1253 & ~n1254;
  assign n1256 = pi14  & ~n1255;
  assign n1257 = pi14  & ~n1256;
  assign n1258 = ~n1255 & ~n1256;
  assign n1259 = ~n1257 & ~n1258;
  assign n1260 = pi17  & ~n1150;
  assign n1261 = ~pi15  & pi16 ;
  assign n1262 = pi15  & ~pi16 ;
  assign n1263 = ~n1261 & ~n1262;
  assign n1264 = n1149 & ~n1263;
  assign n1265 = pi64  & n1264;
  assign n1266 = ~pi16  & pi17 ;
  assign n1267 = pi16  & ~pi17 ;
  assign n1268 = ~n1266 & ~n1267;
  assign n1269 = ~n1149 & n1268;
  assign n1270 = pi65  & n1269;
  assign n1271 = ~n1265 & ~n1270;
  assign n1272 = ~n1149 & ~n1268;
  assign n1273 = n270 & n1272;
  assign n1274 = n1271 & ~n1273;
  assign n1275 = pi17  & ~n1274;
  assign n1276 = pi17  & ~n1275;
  assign n1277 = ~n1274 & ~n1275;
  assign n1278 = ~n1276 & ~n1277;
  assign n1279 = n1260 & ~n1278;
  assign n1280 = ~n1260 & n1278;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = n1259 & ~n1281;
  assign n1283 = ~n1259 & n1281;
  assign n1284 = ~n1282 & ~n1283;
  assign n1285 = ~n1248 & n1284;
  assign n1286 = n1248 & ~n1284;
  assign n1287 = ~n1285 & ~n1286;
  assign n1288 = n1247 & ~n1287;
  assign n1289 = ~n1247 & n1287;
  assign n1290 = ~n1288 & ~n1289;
  assign n1291 = ~n1236 & n1290;
  assign n1292 = n1236 & ~n1290;
  assign n1293 = ~n1291 & ~n1292;
  assign n1294 = n1235 & ~n1293;
  assign n1295 = ~n1235 & n1293;
  assign n1296 = ~n1294 & ~n1295;
  assign n1297 = ~n1224 & n1296;
  assign n1298 = n1224 & ~n1296;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = n1223 & ~n1299;
  assign n1301 = ~n1223 & n1299;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = ~n1212 & n1302;
  assign n1304 = n1212 & ~n1302;
  assign n1305 = ~n1303 & ~n1304;
  assign n1306 = n1211 & n1305;
  assign n1307 = ~n1211 & ~n1305;
  assign n1308 = ~n1306 & ~n1307;
  assign n1309 = ~n1193 & ~n1308;
  assign n1310 = n1193 & n1308;
  assign po16  = ~n1309 & ~n1310;
  assign n1312 = ~n1301 & ~n1303;
  assign n1313 = pi78  & n340;
  assign n1314 = pi76  & n380;
  assign n1315 = pi77  & n335;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317 = ~n1313 & n1316;
  assign n1318 = n343 & n1009;
  assign n1319 = n1317 & ~n1318;
  assign n1320 = pi5  & ~n1319;
  assign n1321 = pi5  & ~n1320;
  assign n1322 = ~n1319 & ~n1320;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = ~n1295 & ~n1297;
  assign n1325 = pi75  & n493;
  assign n1326 = pi73  & n533;
  assign n1327 = pi74  & n488;
  assign n1328 = ~n1326 & ~n1327;
  assign n1329 = ~n1325 & n1328;
  assign n1330 = n496 & n747;
  assign n1331 = n1329 & ~n1330;
  assign n1332 = pi8  & ~n1331;
  assign n1333 = pi8  & ~n1332;
  assign n1334 = ~n1331 & ~n1332;
  assign n1335 = ~n1333 & ~n1334;
  assign n1336 = ~n1289 & ~n1291;
  assign n1337 = ~n1283 & ~n1285;
  assign n1338 = pi66  & n1269;
  assign n1339 = n1149 & ~n1268;
  assign n1340 = n1263 & n1339;
  assign n1341 = pi64  & n1340;
  assign n1342 = pi65  & n1264;
  assign n1343 = ~n1341 & ~n1342;
  assign n1344 = ~n1338 & n1343;
  assign n1345 = n291 & n1272;
  assign n1346 = n1344 & ~n1345;
  assign n1347 = pi17  & ~n1346;
  assign n1348 = pi17  & ~n1347;
  assign n1349 = ~n1346 & ~n1347;
  assign n1350 = ~n1348 & ~n1349;
  assign n1351 = ~n1279 & n1350;
  assign n1352 = n1279 & ~n1350;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = pi69  & n918;
  assign n1355 = pi67  & n1031;
  assign n1356 = pi68  & n913;
  assign n1357 = ~n1355 & ~n1356;
  assign n1358 = ~n1354 & n1357;
  assign n1359 = n405 & n921;
  assign n1360 = n1358 & ~n1359;
  assign n1361 = pi14  & ~n1360;
  assign n1362 = pi14  & ~n1361;
  assign n1363 = ~n1360 & ~n1361;
  assign n1364 = ~n1362 & ~n1363;
  assign n1365 = n1353 & ~n1364;
  assign n1366 = ~n1353 & n1364;
  assign n1367 = ~n1337 & ~n1366;
  assign n1368 = ~n1365 & n1367;
  assign n1369 = ~n1337 & ~n1368;
  assign n1370 = ~n1365 & ~n1368;
  assign n1371 = ~n1366 & n1370;
  assign n1372 = ~n1369 & ~n1371;
  assign n1373 = pi72  & n675;
  assign n1374 = pi70  & n769;
  assign n1375 = pi71  & n670;
  assign n1376 = ~n1374 & ~n1375;
  assign n1377 = ~n1373 & n1376;
  assign n1378 = n575 & n678;
  assign n1379 = n1377 & ~n1378;
  assign n1380 = pi11  & ~n1379;
  assign n1381 = pi11  & ~n1380;
  assign n1382 = ~n1379 & ~n1380;
  assign n1383 = ~n1381 & ~n1382;
  assign n1384 = n1372 & n1383;
  assign n1385 = ~n1372 & ~n1383;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = ~n1336 & n1386;
  assign n1388 = n1336 & ~n1386;
  assign n1389 = ~n1387 & ~n1388;
  assign n1390 = n1335 & ~n1389;
  assign n1391 = ~n1335 & n1389;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = ~n1324 & n1392;
  assign n1394 = n1324 & ~n1392;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = n1323 & ~n1395;
  assign n1397 = ~n1323 & n1395;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = ~n1312 & n1398;
  assign n1400 = n1312 & ~n1398;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = pi81  & n264;
  assign n1403 = pi79  & n281;
  assign n1404 = pi80  & n259;
  assign n1405 = ~n1403 & ~n1404;
  assign n1406 = ~n1402 & n1405;
  assign n1407 = ~n1201 & ~n1203;
  assign n1408 = ~pi80  & ~pi81 ;
  assign n1409 = pi80  & pi81 ;
  assign n1410 = ~n1408 & ~n1409;
  assign n1411 = ~n1407 & n1410;
  assign n1412 = n1407 & ~n1410;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = n267 & n1413;
  assign n1415 = n1406 & ~n1414;
  assign n1416 = pi2  & ~n1415;
  assign n1417 = pi2  & ~n1416;
  assign n1418 = ~n1415 & ~n1416;
  assign n1419 = ~n1417 & ~n1418;
  assign n1420 = n1401 & ~n1419;
  assign n1421 = n1401 & ~n1420;
  assign n1422 = ~n1419 & ~n1420;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = ~n1211 & n1305;
  assign n1425 = ~n1309 & ~n1424;
  assign n1426 = ~n1423 & ~n1425;
  assign n1427 = n1423 & n1425;
  assign po17  = ~n1426 & ~n1427;
  assign n1429 = ~n1397 & ~n1399;
  assign n1430 = pi79  & n340;
  assign n1431 = pi77  & n380;
  assign n1432 = pi78  & n335;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = ~n1430 & n1433;
  assign n1435 = n343 & n1105;
  assign n1436 = n1434 & ~n1435;
  assign n1437 = pi5  & ~n1436;
  assign n1438 = pi5  & ~n1437;
  assign n1439 = ~n1436 & ~n1437;
  assign n1440 = ~n1438 & ~n1439;
  assign n1441 = ~n1391 & ~n1393;
  assign n1442 = pi76  & n493;
  assign n1443 = pi74  & n533;
  assign n1444 = pi75  & n488;
  assign n1445 = ~n1443 & ~n1444;
  assign n1446 = ~n1442 & n1445;
  assign n1447 = n496 & n881;
  assign n1448 = n1446 & ~n1447;
  assign n1449 = pi8  & ~n1448;
  assign n1450 = pi8  & ~n1449;
  assign n1451 = ~n1448 & ~n1449;
  assign n1452 = ~n1450 & ~n1451;
  assign n1453 = ~n1385 & ~n1387;
  assign n1454 = pi73  & n675;
  assign n1455 = pi71  & n769;
  assign n1456 = pi72  & n670;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = ~n1454 & n1457;
  assign n1459 = n639 & n678;
  assign n1460 = n1458 & ~n1459;
  assign n1461 = pi11  & ~n1460;
  assign n1462 = pi11  & ~n1461;
  assign n1463 = ~n1460 & ~n1461;
  assign n1464 = ~n1462 & ~n1463;
  assign n1465 = pi67  & n1269;
  assign n1466 = pi65  & n1340;
  assign n1467 = pi66  & n1264;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = ~n1465 & n1468;
  assign n1470 = n313 & n1272;
  assign n1471 = n1469 & ~n1470;
  assign n1472 = pi17  & ~n1471;
  assign n1473 = pi17  & ~n1472;
  assign n1474 = ~n1471 & ~n1472;
  assign n1475 = ~n1473 & ~n1474;
  assign n1476 = pi17  & ~pi18 ;
  assign n1477 = ~pi17  & pi18 ;
  assign n1478 = ~n1476 & ~n1477;
  assign n1479 = pi64  & ~n1478;
  assign n1480 = n1352 & n1479;
  assign n1481 = ~n1352 & ~n1479;
  assign n1482 = ~n1480 & ~n1481;
  assign n1483 = ~n1475 & n1482;
  assign n1484 = n1475 & ~n1482;
  assign n1485 = ~n1483 & ~n1484;
  assign n1486 = pi70  & n918;
  assign n1487 = pi68  & n1031;
  assign n1488 = pi69  & n913;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = ~n1486 & n1489;
  assign n1491 = n430 & n921;
  assign n1492 = n1490 & ~n1491;
  assign n1493 = pi14  & ~n1492;
  assign n1494 = pi14  & ~n1493;
  assign n1495 = ~n1492 & ~n1493;
  assign n1496 = ~n1494 & ~n1495;
  assign n1497 = n1485 & ~n1496;
  assign n1498 = ~n1485 & n1496;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = ~n1370 & n1499;
  assign n1501 = n1370 & ~n1499;
  assign n1502 = ~n1500 & ~n1501;
  assign n1503 = ~n1464 & n1502;
  assign n1504 = n1464 & ~n1502;
  assign n1505 = ~n1503 & ~n1504;
  assign n1506 = ~n1453 & n1505;
  assign n1507 = n1453 & ~n1505;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = n1452 & ~n1508;
  assign n1510 = ~n1452 & n1508;
  assign n1511 = ~n1509 & ~n1510;
  assign n1512 = ~n1441 & n1511;
  assign n1513 = n1441 & ~n1511;
  assign n1514 = ~n1512 & ~n1513;
  assign n1515 = ~n1440 & n1514;
  assign n1516 = n1440 & ~n1514;
  assign n1517 = ~n1515 & ~n1516;
  assign n1518 = ~n1429 & n1517;
  assign n1519 = n1429 & ~n1517;
  assign n1520 = ~n1518 & ~n1519;
  assign n1521 = pi82  & n264;
  assign n1522 = pi80  & n281;
  assign n1523 = pi81  & n259;
  assign n1524 = ~n1522 & ~n1523;
  assign n1525 = ~n1521 & n1524;
  assign n1526 = ~n1409 & ~n1411;
  assign n1527 = ~pi81  & ~pi82 ;
  assign n1528 = pi81  & pi82 ;
  assign n1529 = ~n1527 & ~n1528;
  assign n1530 = ~n1526 & n1529;
  assign n1531 = n1526 & ~n1529;
  assign n1532 = ~n1530 & ~n1531;
  assign n1533 = n267 & n1532;
  assign n1534 = n1525 & ~n1533;
  assign n1535 = pi2  & ~n1534;
  assign n1536 = pi2  & ~n1535;
  assign n1537 = ~n1534 & ~n1535;
  assign n1538 = ~n1536 & ~n1537;
  assign n1539 = n1520 & ~n1538;
  assign n1540 = n1520 & ~n1539;
  assign n1541 = ~n1538 & ~n1539;
  assign n1542 = ~n1540 & ~n1541;
  assign n1543 = ~n1420 & ~n1426;
  assign n1544 = ~n1542 & ~n1543;
  assign n1545 = n1542 & n1543;
  assign po18  = ~n1544 & ~n1545;
  assign n1547 = ~n1539 & ~n1544;
  assign n1548 = ~n1503 & ~n1506;
  assign n1549 = ~n1497 & ~n1500;
  assign n1550 = pi71  & n918;
  assign n1551 = pi69  & n1031;
  assign n1552 = pi70  & n913;
  assign n1553 = ~n1551 & ~n1552;
  assign n1554 = ~n1550 & n1553;
  assign n1555 = n476 & n921;
  assign n1556 = n1554 & ~n1555;
  assign n1557 = pi14  & ~n1556;
  assign n1558 = pi14  & ~n1557;
  assign n1559 = ~n1556 & ~n1557;
  assign n1560 = ~n1558 & ~n1559;
  assign n1561 = ~n1480 & ~n1483;
  assign n1562 = pi68  & n1269;
  assign n1563 = pi66  & n1340;
  assign n1564 = pi67  & n1264;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = ~n1562 & n1565;
  assign n1567 = n364 & n1272;
  assign n1568 = n1566 & ~n1567;
  assign n1569 = pi17  & ~n1568;
  assign n1570 = pi17  & ~n1569;
  assign n1571 = ~n1568 & ~n1569;
  assign n1572 = ~n1570 & ~n1571;
  assign n1573 = pi20  & ~n1479;
  assign n1574 = ~pi18  & pi19 ;
  assign n1575 = pi18  & ~pi19 ;
  assign n1576 = ~n1574 & ~n1575;
  assign n1577 = n1478 & ~n1576;
  assign n1578 = pi64  & n1577;
  assign n1579 = ~pi19  & pi20 ;
  assign n1580 = pi19  & ~pi20 ;
  assign n1581 = ~n1579 & ~n1580;
  assign n1582 = ~n1478 & n1581;
  assign n1583 = pi65  & n1582;
  assign n1584 = ~n1578 & ~n1583;
  assign n1585 = ~n1478 & ~n1581;
  assign n1586 = n270 & n1585;
  assign n1587 = n1584 & ~n1586;
  assign n1588 = pi20  & ~n1587;
  assign n1589 = pi20  & ~n1588;
  assign n1590 = ~n1587 & ~n1588;
  assign n1591 = ~n1589 & ~n1590;
  assign n1592 = n1573 & ~n1591;
  assign n1593 = ~n1573 & n1591;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = ~n1572 & n1594;
  assign n1596 = n1572 & ~n1594;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n1561 & n1597;
  assign n1599 = n1561 & ~n1597;
  assign n1600 = ~n1598 & ~n1599;
  assign n1601 = ~n1560 & n1600;
  assign n1602 = n1560 & ~n1600;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = ~n1549 & n1603;
  assign n1605 = n1549 & ~n1603;
  assign n1606 = ~n1604 & ~n1605;
  assign n1607 = pi74  & n675;
  assign n1608 = pi72  & n769;
  assign n1609 = pi73  & n670;
  assign n1610 = ~n1608 & ~n1609;
  assign n1611 = ~n1607 & n1610;
  assign n1612 = n678 & n722;
  assign n1613 = n1611 & ~n1612;
  assign n1614 = pi11  & ~n1613;
  assign n1615 = pi11  & ~n1614;
  assign n1616 = ~n1613 & ~n1614;
  assign n1617 = ~n1615 & ~n1616;
  assign n1618 = n1606 & ~n1617;
  assign n1619 = ~n1606 & n1617;
  assign n1620 = ~n1618 & ~n1619;
  assign n1621 = n1548 & ~n1620;
  assign n1622 = ~n1548 & n1620;
  assign n1623 = ~n1621 & ~n1622;
  assign n1624 = pi77  & n493;
  assign n1625 = pi75  & n533;
  assign n1626 = pi76  & n488;
  assign n1627 = ~n1625 & ~n1626;
  assign n1628 = ~n1624 & n1627;
  assign n1629 = n496 & n984;
  assign n1630 = n1628 & ~n1629;
  assign n1631 = pi8  & ~n1630;
  assign n1632 = pi8  & ~n1631;
  assign n1633 = ~n1630 & ~n1631;
  assign n1634 = ~n1632 & ~n1633;
  assign n1635 = ~n1623 & n1634;
  assign n1636 = n1623 & ~n1634;
  assign n1637 = ~n1635 & ~n1636;
  assign n1638 = ~n1510 & ~n1512;
  assign n1639 = n1637 & ~n1638;
  assign n1640 = ~n1637 & n1638;
  assign n1641 = ~n1639 & ~n1640;
  assign n1642 = pi80  & n340;
  assign n1643 = pi78  & n380;
  assign n1644 = pi79  & n335;
  assign n1645 = ~n1643 & ~n1644;
  assign n1646 = ~n1642 & n1645;
  assign n1647 = n343 & n1205;
  assign n1648 = n1646 & ~n1647;
  assign n1649 = pi5  & ~n1648;
  assign n1650 = pi5  & ~n1649;
  assign n1651 = ~n1648 & ~n1649;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = n1641 & ~n1652;
  assign n1654 = n1641 & ~n1653;
  assign n1655 = ~n1652 & ~n1653;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = ~n1515 & ~n1518;
  assign n1658 = n1656 & n1657;
  assign n1659 = ~n1656 & ~n1657;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = pi83  & n264;
  assign n1662 = pi81  & n281;
  assign n1663 = pi82  & n259;
  assign n1664 = ~n1662 & ~n1663;
  assign n1665 = ~n1661 & n1664;
  assign n1666 = ~n1528 & ~n1530;
  assign n1667 = ~pi82  & ~pi83 ;
  assign n1668 = pi82  & pi83 ;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = ~n1666 & n1669;
  assign n1671 = n1666 & ~n1669;
  assign n1672 = ~n1670 & ~n1671;
  assign n1673 = n267 & n1672;
  assign n1674 = n1665 & ~n1673;
  assign n1675 = pi2  & ~n1674;
  assign n1676 = pi2  & ~n1675;
  assign n1677 = ~n1674 & ~n1675;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = n1660 & ~n1678;
  assign n1680 = ~n1660 & n1678;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = ~n1547 & n1681;
  assign n1683 = n1547 & ~n1681;
  assign po19  = ~n1682 & ~n1683;
  assign n1685 = ~n1653 & ~n1659;
  assign n1686 = pi81  & n340;
  assign n1687 = pi79  & n380;
  assign n1688 = pi80  & n335;
  assign n1689 = ~n1687 & ~n1688;
  assign n1690 = ~n1686 & n1689;
  assign n1691 = n343 & n1413;
  assign n1692 = n1690 & ~n1691;
  assign n1693 = pi5  & ~n1692;
  assign n1694 = pi5  & ~n1693;
  assign n1695 = ~n1692 & ~n1693;
  assign n1696 = ~n1694 & ~n1695;
  assign n1697 = ~n1618 & ~n1622;
  assign n1698 = pi75  & n675;
  assign n1699 = pi73  & n769;
  assign n1700 = pi74  & n670;
  assign n1701 = ~n1699 & ~n1700;
  assign n1702 = ~n1698 & n1701;
  assign n1703 = n678 & n747;
  assign n1704 = n1702 & ~n1703;
  assign n1705 = pi11  & ~n1704;
  assign n1706 = pi11  & ~n1705;
  assign n1707 = ~n1704 & ~n1705;
  assign n1708 = ~n1706 & ~n1707;
  assign n1709 = ~n1601 & ~n1604;
  assign n1710 = ~n1595 & ~n1598;
  assign n1711 = pi66  & n1582;
  assign n1712 = n1478 & ~n1581;
  assign n1713 = n1576 & n1712;
  assign n1714 = pi64  & n1713;
  assign n1715 = pi65  & n1577;
  assign n1716 = ~n1714 & ~n1715;
  assign n1717 = ~n1711 & n1716;
  assign n1718 = n291 & n1585;
  assign n1719 = n1717 & ~n1718;
  assign n1720 = pi20  & ~n1719;
  assign n1721 = pi20  & ~n1720;
  assign n1722 = ~n1719 & ~n1720;
  assign n1723 = ~n1721 & ~n1722;
  assign n1724 = ~n1592 & n1723;
  assign n1725 = n1592 & ~n1723;
  assign n1726 = ~n1724 & ~n1725;
  assign n1727 = pi69  & n1269;
  assign n1728 = pi67  & n1340;
  assign n1729 = pi68  & n1264;
  assign n1730 = ~n1728 & ~n1729;
  assign n1731 = ~n1727 & n1730;
  assign n1732 = n405 & n1272;
  assign n1733 = n1731 & ~n1732;
  assign n1734 = pi17  & ~n1733;
  assign n1735 = pi17  & ~n1734;
  assign n1736 = ~n1733 & ~n1734;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = n1726 & ~n1737;
  assign n1739 = ~n1726 & n1737;
  assign n1740 = ~n1710 & ~n1739;
  assign n1741 = ~n1738 & n1740;
  assign n1742 = ~n1710 & ~n1741;
  assign n1743 = ~n1738 & ~n1741;
  assign n1744 = ~n1739 & n1743;
  assign n1745 = ~n1742 & ~n1744;
  assign n1746 = pi72  & n918;
  assign n1747 = pi70  & n1031;
  assign n1748 = pi71  & n913;
  assign n1749 = ~n1747 & ~n1748;
  assign n1750 = ~n1746 & n1749;
  assign n1751 = n575 & n921;
  assign n1752 = n1750 & ~n1751;
  assign n1753 = pi14  & ~n1752;
  assign n1754 = pi14  & ~n1753;
  assign n1755 = ~n1752 & ~n1753;
  assign n1756 = ~n1754 & ~n1755;
  assign n1757 = n1745 & n1756;
  assign n1758 = ~n1745 & ~n1756;
  assign n1759 = ~n1757 & ~n1758;
  assign n1760 = ~n1709 & n1759;
  assign n1761 = n1709 & ~n1759;
  assign n1762 = ~n1760 & ~n1761;
  assign n1763 = n1708 & ~n1762;
  assign n1764 = ~n1708 & n1762;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = ~n1697 & n1765;
  assign n1767 = n1697 & ~n1765;
  assign n1768 = ~n1766 & ~n1767;
  assign n1769 = pi78  & n493;
  assign n1770 = pi76  & n533;
  assign n1771 = pi77  & n488;
  assign n1772 = ~n1770 & ~n1771;
  assign n1773 = ~n1769 & n1772;
  assign n1774 = n496 & n1009;
  assign n1775 = n1773 & ~n1774;
  assign n1776 = pi8  & ~n1775;
  assign n1777 = pi8  & ~n1776;
  assign n1778 = ~n1775 & ~n1776;
  assign n1779 = ~n1777 & ~n1778;
  assign n1780 = n1768 & ~n1779;
  assign n1781 = n1768 & ~n1780;
  assign n1782 = ~n1779 & ~n1780;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = ~n1636 & ~n1639;
  assign n1785 = ~n1783 & ~n1784;
  assign n1786 = n1783 & n1784;
  assign n1787 = ~n1785 & ~n1786;
  assign n1788 = ~n1696 & n1787;
  assign n1789 = n1696 & ~n1787;
  assign n1790 = ~n1788 & ~n1789;
  assign n1791 = ~n1685 & n1790;
  assign n1792 = n1685 & ~n1790;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = pi84  & n264;
  assign n1795 = pi82  & n281;
  assign n1796 = pi83  & n259;
  assign n1797 = ~n1795 & ~n1796;
  assign n1798 = ~n1794 & n1797;
  assign n1799 = ~n1668 & ~n1670;
  assign n1800 = ~pi83  & ~pi84 ;
  assign n1801 = pi83  & pi84 ;
  assign n1802 = ~n1800 & ~n1801;
  assign n1803 = ~n1799 & n1802;
  assign n1804 = n1799 & ~n1802;
  assign n1805 = ~n1803 & ~n1804;
  assign n1806 = n267 & n1805;
  assign n1807 = n1798 & ~n1806;
  assign n1808 = pi2  & ~n1807;
  assign n1809 = pi2  & ~n1808;
  assign n1810 = ~n1807 & ~n1808;
  assign n1811 = ~n1809 & ~n1810;
  assign n1812 = n1793 & ~n1811;
  assign n1813 = n1793 & ~n1812;
  assign n1814 = ~n1811 & ~n1812;
  assign n1815 = ~n1813 & ~n1814;
  assign n1816 = ~n1679 & ~n1682;
  assign n1817 = ~n1815 & ~n1816;
  assign n1818 = n1815 & n1816;
  assign po20  = ~n1817 & ~n1818;
  assign n1820 = ~n1812 & ~n1817;
  assign n1821 = ~n1780 & ~n1785;
  assign n1822 = pi79  & n493;
  assign n1823 = pi77  & n533;
  assign n1824 = pi78  & n488;
  assign n1825 = ~n1823 & ~n1824;
  assign n1826 = ~n1822 & n1825;
  assign n1827 = n496 & n1105;
  assign n1828 = n1826 & ~n1827;
  assign n1829 = pi8  & ~n1828;
  assign n1830 = pi8  & ~n1829;
  assign n1831 = ~n1828 & ~n1829;
  assign n1832 = ~n1830 & ~n1831;
  assign n1833 = ~n1764 & ~n1766;
  assign n1834 = pi76  & n675;
  assign n1835 = pi74  & n769;
  assign n1836 = pi75  & n670;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = ~n1834 & n1837;
  assign n1839 = n678 & n881;
  assign n1840 = n1838 & ~n1839;
  assign n1841 = pi11  & ~n1840;
  assign n1842 = pi11  & ~n1841;
  assign n1843 = ~n1840 & ~n1841;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = ~n1758 & ~n1760;
  assign n1846 = pi73  & n918;
  assign n1847 = pi71  & n1031;
  assign n1848 = pi72  & n913;
  assign n1849 = ~n1847 & ~n1848;
  assign n1850 = ~n1846 & n1849;
  assign n1851 = n639 & n921;
  assign n1852 = n1850 & ~n1851;
  assign n1853 = pi14  & ~n1852;
  assign n1854 = pi14  & ~n1853;
  assign n1855 = ~n1852 & ~n1853;
  assign n1856 = ~n1854 & ~n1855;
  assign n1857 = pi67  & n1582;
  assign n1858 = pi65  & n1713;
  assign n1859 = pi66  & n1577;
  assign n1860 = ~n1858 & ~n1859;
  assign n1861 = ~n1857 & n1860;
  assign n1862 = n313 & n1585;
  assign n1863 = n1861 & ~n1862;
  assign n1864 = pi20  & ~n1863;
  assign n1865 = pi20  & ~n1864;
  assign n1866 = ~n1863 & ~n1864;
  assign n1867 = ~n1865 & ~n1866;
  assign n1868 = pi20  & ~pi21 ;
  assign n1869 = ~pi20  & pi21 ;
  assign n1870 = ~n1868 & ~n1869;
  assign n1871 = pi64  & ~n1870;
  assign n1872 = n1725 & n1871;
  assign n1873 = ~n1725 & ~n1871;
  assign n1874 = ~n1872 & ~n1873;
  assign n1875 = ~n1867 & n1874;
  assign n1876 = n1867 & ~n1874;
  assign n1877 = ~n1875 & ~n1876;
  assign n1878 = pi70  & n1269;
  assign n1879 = pi68  & n1340;
  assign n1880 = pi69  & n1264;
  assign n1881 = ~n1879 & ~n1880;
  assign n1882 = ~n1878 & n1881;
  assign n1883 = n430 & n1272;
  assign n1884 = n1882 & ~n1883;
  assign n1885 = pi17  & ~n1884;
  assign n1886 = pi17  & ~n1885;
  assign n1887 = ~n1884 & ~n1885;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = n1877 & ~n1888;
  assign n1890 = ~n1877 & n1888;
  assign n1891 = ~n1889 & ~n1890;
  assign n1892 = ~n1743 & n1891;
  assign n1893 = n1743 & ~n1891;
  assign n1894 = ~n1892 & ~n1893;
  assign n1895 = ~n1856 & n1894;
  assign n1896 = n1856 & ~n1894;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = ~n1845 & n1897;
  assign n1899 = n1845 & ~n1897;
  assign n1900 = ~n1898 & ~n1899;
  assign n1901 = n1844 & ~n1900;
  assign n1902 = ~n1844 & n1900;
  assign n1903 = ~n1901 & ~n1902;
  assign n1904 = ~n1833 & n1903;
  assign n1905 = n1833 & ~n1903;
  assign n1906 = ~n1904 & ~n1905;
  assign n1907 = ~n1832 & n1906;
  assign n1908 = n1832 & ~n1906;
  assign n1909 = ~n1907 & ~n1908;
  assign n1910 = ~n1821 & n1909;
  assign n1911 = n1821 & ~n1909;
  assign n1912 = ~n1910 & ~n1911;
  assign n1913 = pi82  & n340;
  assign n1914 = pi80  & n380;
  assign n1915 = pi81  & n335;
  assign n1916 = ~n1914 & ~n1915;
  assign n1917 = ~n1913 & n1916;
  assign n1918 = n343 & n1532;
  assign n1919 = n1917 & ~n1918;
  assign n1920 = pi5  & ~n1919;
  assign n1921 = pi5  & ~n1920;
  assign n1922 = ~n1919 & ~n1920;
  assign n1923 = ~n1921 & ~n1922;
  assign n1924 = n1912 & ~n1923;
  assign n1925 = n1912 & ~n1924;
  assign n1926 = ~n1923 & ~n1924;
  assign n1927 = ~n1925 & ~n1926;
  assign n1928 = ~n1788 & ~n1791;
  assign n1929 = n1927 & n1928;
  assign n1930 = ~n1927 & ~n1928;
  assign n1931 = ~n1929 & ~n1930;
  assign n1932 = pi85  & n264;
  assign n1933 = pi83  & n281;
  assign n1934 = pi84  & n259;
  assign n1935 = ~n1933 & ~n1934;
  assign n1936 = ~n1932 & n1935;
  assign n1937 = ~n1801 & ~n1803;
  assign n1938 = ~pi84  & ~pi85 ;
  assign n1939 = pi84  & pi85 ;
  assign n1940 = ~n1938 & ~n1939;
  assign n1941 = ~n1937 & n1940;
  assign n1942 = n1937 & ~n1940;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = n267 & n1943;
  assign n1945 = n1936 & ~n1944;
  assign n1946 = pi2  & ~n1945;
  assign n1947 = pi2  & ~n1946;
  assign n1948 = ~n1945 & ~n1946;
  assign n1949 = ~n1947 & ~n1948;
  assign n1950 = n1931 & ~n1949;
  assign n1951 = ~n1931 & n1949;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = ~n1820 & n1952;
  assign n1954 = n1820 & ~n1952;
  assign po21  = ~n1953 & ~n1954;
  assign n1956 = ~n1950 & ~n1953;
  assign n1957 = ~n1907 & ~n1910;
  assign n1958 = pi80  & n493;
  assign n1959 = pi78  & n533;
  assign n1960 = pi79  & n488;
  assign n1961 = ~n1959 & ~n1960;
  assign n1962 = ~n1958 & n1961;
  assign n1963 = n496 & n1205;
  assign n1964 = n1962 & ~n1963;
  assign n1965 = pi8  & ~n1964;
  assign n1966 = pi8  & ~n1965;
  assign n1967 = ~n1964 & ~n1965;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = ~n1902 & ~n1904;
  assign n1970 = ~n1895 & ~n1898;
  assign n1971 = ~n1889 & ~n1892;
  assign n1972 = pi71  & n1269;
  assign n1973 = pi69  & n1340;
  assign n1974 = pi70  & n1264;
  assign n1975 = ~n1973 & ~n1974;
  assign n1976 = ~n1972 & n1975;
  assign n1977 = n476 & n1272;
  assign n1978 = n1976 & ~n1977;
  assign n1979 = pi17  & ~n1978;
  assign n1980 = pi17  & ~n1979;
  assign n1981 = ~n1978 & ~n1979;
  assign n1982 = ~n1980 & ~n1981;
  assign n1983 = ~n1872 & ~n1875;
  assign n1984 = pi68  & n1582;
  assign n1985 = pi66  & n1713;
  assign n1986 = pi67  & n1577;
  assign n1987 = ~n1985 & ~n1986;
  assign n1988 = ~n1984 & n1987;
  assign n1989 = n364 & n1585;
  assign n1990 = n1988 & ~n1989;
  assign n1991 = pi20  & ~n1990;
  assign n1992 = pi20  & ~n1991;
  assign n1993 = ~n1990 & ~n1991;
  assign n1994 = ~n1992 & ~n1993;
  assign n1995 = pi23  & ~n1871;
  assign n1996 = ~pi21  & pi22 ;
  assign n1997 = pi21  & ~pi22 ;
  assign n1998 = ~n1996 & ~n1997;
  assign n1999 = n1870 & ~n1998;
  assign n2000 = pi64  & n1999;
  assign n2001 = ~pi22  & pi23 ;
  assign n2002 = pi22  & ~pi23 ;
  assign n2003 = ~n2001 & ~n2002;
  assign n2004 = ~n1870 & n2003;
  assign n2005 = pi65  & n2004;
  assign n2006 = ~n2000 & ~n2005;
  assign n2007 = ~n1870 & ~n2003;
  assign n2008 = n270 & n2007;
  assign n2009 = n2006 & ~n2008;
  assign n2010 = pi23  & ~n2009;
  assign n2011 = pi23  & ~n2010;
  assign n2012 = ~n2009 & ~n2010;
  assign n2013 = ~n2011 & ~n2012;
  assign n2014 = n1995 & ~n2013;
  assign n2015 = ~n1995 & n2013;
  assign n2016 = ~n2014 & ~n2015;
  assign n2017 = ~n1994 & n2016;
  assign n2018 = n1994 & ~n2016;
  assign n2019 = ~n2017 & ~n2018;
  assign n2020 = ~n1983 & n2019;
  assign n2021 = n1983 & ~n2019;
  assign n2022 = ~n2020 & ~n2021;
  assign n2023 = ~n1982 & n2022;
  assign n2024 = n1982 & ~n2022;
  assign n2025 = ~n2023 & ~n2024;
  assign n2026 = ~n1971 & n2025;
  assign n2027 = n1971 & ~n2025;
  assign n2028 = ~n2026 & ~n2027;
  assign n2029 = pi74  & n918;
  assign n2030 = pi72  & n1031;
  assign n2031 = pi73  & n913;
  assign n2032 = ~n2030 & ~n2031;
  assign n2033 = ~n2029 & n2032;
  assign n2034 = n722 & n921;
  assign n2035 = n2033 & ~n2034;
  assign n2036 = pi14  & ~n2035;
  assign n2037 = pi14  & ~n2036;
  assign n2038 = ~n2035 & ~n2036;
  assign n2039 = ~n2037 & ~n2038;
  assign n2040 = n2028 & ~n2039;
  assign n2041 = ~n2028 & n2039;
  assign n2042 = ~n2040 & ~n2041;
  assign n2043 = n1970 & ~n2042;
  assign n2044 = ~n1970 & n2042;
  assign n2045 = ~n2043 & ~n2044;
  assign n2046 = pi77  & n675;
  assign n2047 = pi75  & n769;
  assign n2048 = pi76  & n670;
  assign n2049 = ~n2047 & ~n2048;
  assign n2050 = ~n2046 & n2049;
  assign n2051 = n678 & n984;
  assign n2052 = n2050 & ~n2051;
  assign n2053 = pi11  & ~n2052;
  assign n2054 = pi11  & ~n2053;
  assign n2055 = ~n2052 & ~n2053;
  assign n2056 = ~n2054 & ~n2055;
  assign n2057 = ~n2045 & n2056;
  assign n2058 = n2045 & ~n2056;
  assign n2059 = ~n2057 & ~n2058;
  assign n2060 = ~n1969 & n2059;
  assign n2061 = n1969 & ~n2059;
  assign n2062 = ~n2060 & ~n2061;
  assign n2063 = ~n1968 & n2062;
  assign n2064 = n1968 & ~n2062;
  assign n2065 = ~n2063 & ~n2064;
  assign n2066 = ~n1957 & n2065;
  assign n2067 = n1957 & ~n2065;
  assign n2068 = ~n2066 & ~n2067;
  assign n2069 = pi83  & n340;
  assign n2070 = pi81  & n380;
  assign n2071 = pi82  & n335;
  assign n2072 = ~n2070 & ~n2071;
  assign n2073 = ~n2069 & n2072;
  assign n2074 = n343 & n1672;
  assign n2075 = n2073 & ~n2074;
  assign n2076 = pi5  & ~n2075;
  assign n2077 = pi5  & ~n2076;
  assign n2078 = ~n2075 & ~n2076;
  assign n2079 = ~n2077 & ~n2078;
  assign n2080 = n2068 & ~n2079;
  assign n2081 = n2068 & ~n2080;
  assign n2082 = ~n2079 & ~n2080;
  assign n2083 = ~n2081 & ~n2082;
  assign n2084 = ~n1924 & ~n1930;
  assign n2085 = n2083 & n2084;
  assign n2086 = ~n2083 & ~n2084;
  assign n2087 = ~n2085 & ~n2086;
  assign n2088 = pi86  & n264;
  assign n2089 = pi84  & n281;
  assign n2090 = pi85  & n259;
  assign n2091 = ~n2089 & ~n2090;
  assign n2092 = ~n2088 & n2091;
  assign n2093 = ~n1939 & ~n1941;
  assign n2094 = ~pi85  & ~pi86 ;
  assign n2095 = pi85  & pi86 ;
  assign n2096 = ~n2094 & ~n2095;
  assign n2097 = ~n2093 & n2096;
  assign n2098 = n2093 & ~n2096;
  assign n2099 = ~n2097 & ~n2098;
  assign n2100 = n267 & n2099;
  assign n2101 = n2092 & ~n2100;
  assign n2102 = pi2  & ~n2101;
  assign n2103 = pi2  & ~n2102;
  assign n2104 = ~n2101 & ~n2102;
  assign n2105 = ~n2103 & ~n2104;
  assign n2106 = ~n2087 & n2105;
  assign n2107 = n2087 & ~n2105;
  assign n2108 = ~n2106 & ~n2107;
  assign n2109 = ~n1956 & n2108;
  assign n2110 = n1956 & ~n2108;
  assign po22  = ~n2109 & ~n2110;
  assign n2112 = ~n2107 & ~n2109;
  assign n2113 = ~n2063 & ~n2066;
  assign n2114 = pi81  & n493;
  assign n2115 = pi79  & n533;
  assign n2116 = pi80  & n488;
  assign n2117 = ~n2115 & ~n2116;
  assign n2118 = ~n2114 & n2117;
  assign n2119 = n496 & n1413;
  assign n2120 = n2118 & ~n2119;
  assign n2121 = pi8  & ~n2120;
  assign n2122 = pi8  & ~n2121;
  assign n2123 = ~n2120 & ~n2121;
  assign n2124 = ~n2122 & ~n2123;
  assign n2125 = ~n2040 & ~n2044;
  assign n2126 = pi75  & n918;
  assign n2127 = pi73  & n1031;
  assign n2128 = pi74  & n913;
  assign n2129 = ~n2127 & ~n2128;
  assign n2130 = ~n2126 & n2129;
  assign n2131 = n747 & n921;
  assign n2132 = n2130 & ~n2131;
  assign n2133 = pi14  & ~n2132;
  assign n2134 = pi14  & ~n2133;
  assign n2135 = ~n2132 & ~n2133;
  assign n2136 = ~n2134 & ~n2135;
  assign n2137 = ~n2023 & ~n2026;
  assign n2138 = ~n2017 & ~n2020;
  assign n2139 = pi66  & n2004;
  assign n2140 = n1870 & ~n2003;
  assign n2141 = n1998 & n2140;
  assign n2142 = pi64  & n2141;
  assign n2143 = pi65  & n1999;
  assign n2144 = ~n2142 & ~n2143;
  assign n2145 = ~n2139 & n2144;
  assign n2146 = n291 & n2007;
  assign n2147 = n2145 & ~n2146;
  assign n2148 = pi23  & ~n2147;
  assign n2149 = pi23  & ~n2148;
  assign n2150 = ~n2147 & ~n2148;
  assign n2151 = ~n2149 & ~n2150;
  assign n2152 = ~n2014 & n2151;
  assign n2153 = n2014 & ~n2151;
  assign n2154 = ~n2152 & ~n2153;
  assign n2155 = pi69  & n1582;
  assign n2156 = pi67  & n1713;
  assign n2157 = pi68  & n1577;
  assign n2158 = ~n2156 & ~n2157;
  assign n2159 = ~n2155 & n2158;
  assign n2160 = n405 & n1585;
  assign n2161 = n2159 & ~n2160;
  assign n2162 = pi20  & ~n2161;
  assign n2163 = pi20  & ~n2162;
  assign n2164 = ~n2161 & ~n2162;
  assign n2165 = ~n2163 & ~n2164;
  assign n2166 = n2154 & ~n2165;
  assign n2167 = ~n2154 & n2165;
  assign n2168 = ~n2138 & ~n2167;
  assign n2169 = ~n2166 & n2168;
  assign n2170 = ~n2138 & ~n2169;
  assign n2171 = ~n2166 & ~n2169;
  assign n2172 = ~n2167 & n2171;
  assign n2173 = ~n2170 & ~n2172;
  assign n2174 = pi72  & n1269;
  assign n2175 = pi70  & n1340;
  assign n2176 = pi71  & n1264;
  assign n2177 = ~n2175 & ~n2176;
  assign n2178 = ~n2174 & n2177;
  assign n2179 = n575 & n1272;
  assign n2180 = n2178 & ~n2179;
  assign n2181 = pi17  & ~n2180;
  assign n2182 = pi17  & ~n2181;
  assign n2183 = ~n2180 & ~n2181;
  assign n2184 = ~n2182 & ~n2183;
  assign n2185 = n2173 & n2184;
  assign n2186 = ~n2173 & ~n2184;
  assign n2187 = ~n2185 & ~n2186;
  assign n2188 = ~n2137 & n2187;
  assign n2189 = n2137 & ~n2187;
  assign n2190 = ~n2188 & ~n2189;
  assign n2191 = n2136 & ~n2190;
  assign n2192 = ~n2136 & n2190;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = ~n2125 & n2193;
  assign n2195 = n2125 & ~n2193;
  assign n2196 = ~n2194 & ~n2195;
  assign n2197 = pi78  & n675;
  assign n2198 = pi76  & n769;
  assign n2199 = pi77  & n670;
  assign n2200 = ~n2198 & ~n2199;
  assign n2201 = ~n2197 & n2200;
  assign n2202 = n678 & n1009;
  assign n2203 = n2201 & ~n2202;
  assign n2204 = pi11  & ~n2203;
  assign n2205 = pi11  & ~n2204;
  assign n2206 = ~n2203 & ~n2204;
  assign n2207 = ~n2205 & ~n2206;
  assign n2208 = n2196 & ~n2207;
  assign n2209 = n2196 & ~n2208;
  assign n2210 = ~n2207 & ~n2208;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = ~n2058 & ~n2060;
  assign n2213 = ~n2211 & ~n2212;
  assign n2214 = n2211 & n2212;
  assign n2215 = ~n2213 & ~n2214;
  assign n2216 = ~n2124 & n2215;
  assign n2217 = n2124 & ~n2215;
  assign n2218 = ~n2216 & ~n2217;
  assign n2219 = ~n2113 & n2218;
  assign n2220 = n2113 & ~n2218;
  assign n2221 = ~n2219 & ~n2220;
  assign n2222 = pi84  & n340;
  assign n2223 = pi82  & n380;
  assign n2224 = pi83  & n335;
  assign n2225 = ~n2223 & ~n2224;
  assign n2226 = ~n2222 & n2225;
  assign n2227 = n343 & n1805;
  assign n2228 = n2226 & ~n2227;
  assign n2229 = pi5  & ~n2228;
  assign n2230 = pi5  & ~n2229;
  assign n2231 = ~n2228 & ~n2229;
  assign n2232 = ~n2230 & ~n2231;
  assign n2233 = n2221 & ~n2232;
  assign n2234 = n2221 & ~n2233;
  assign n2235 = ~n2232 & ~n2233;
  assign n2236 = ~n2234 & ~n2235;
  assign n2237 = ~n2080 & ~n2086;
  assign n2238 = n2236 & n2237;
  assign n2239 = ~n2236 & ~n2237;
  assign n2240 = ~n2238 & ~n2239;
  assign n2241 = pi87  & n264;
  assign n2242 = pi85  & n281;
  assign n2243 = pi86  & n259;
  assign n2244 = ~n2242 & ~n2243;
  assign n2245 = ~n2241 & n2244;
  assign n2246 = ~n2095 & ~n2097;
  assign n2247 = ~pi86  & ~pi87 ;
  assign n2248 = pi86  & pi87 ;
  assign n2249 = ~n2247 & ~n2248;
  assign n2250 = ~n2246 & n2249;
  assign n2251 = n2246 & ~n2249;
  assign n2252 = ~n2250 & ~n2251;
  assign n2253 = n267 & n2252;
  assign n2254 = n2245 & ~n2253;
  assign n2255 = pi2  & ~n2254;
  assign n2256 = pi2  & ~n2255;
  assign n2257 = ~n2254 & ~n2255;
  assign n2258 = ~n2256 & ~n2257;
  assign n2259 = n2240 & ~n2258;
  assign n2260 = ~n2240 & n2258;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = ~n2112 & n2261;
  assign n2263 = n2112 & ~n2261;
  assign po23  = ~n2262 & ~n2263;
  assign n2265 = ~n2259 & ~n2262;
  assign n2266 = pi88  & n264;
  assign n2267 = pi86  & n281;
  assign n2268 = pi87  & n259;
  assign n2269 = ~n2267 & ~n2268;
  assign n2270 = ~n2266 & n2269;
  assign n2271 = ~n2248 & ~n2250;
  assign n2272 = ~pi87  & ~pi88 ;
  assign n2273 = pi87  & pi88 ;
  assign n2274 = ~n2272 & ~n2273;
  assign n2275 = ~n2271 & n2274;
  assign n2276 = n2271 & ~n2274;
  assign n2277 = ~n2275 & ~n2276;
  assign n2278 = n267 & n2277;
  assign n2279 = n2270 & ~n2278;
  assign n2280 = pi2  & ~n2279;
  assign n2281 = pi2  & ~n2280;
  assign n2282 = ~n2279 & ~n2280;
  assign n2283 = ~n2281 & ~n2282;
  assign n2284 = ~n2233 & ~n2239;
  assign n2285 = pi85  & n340;
  assign n2286 = pi83  & n380;
  assign n2287 = pi84  & n335;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = ~n2285 & n2288;
  assign n2290 = n343 & n1943;
  assign n2291 = n2289 & ~n2290;
  assign n2292 = pi5  & ~n2291;
  assign n2293 = pi5  & ~n2292;
  assign n2294 = ~n2291 & ~n2292;
  assign n2295 = ~n2293 & ~n2294;
  assign n2296 = ~n2216 & ~n2219;
  assign n2297 = ~n2192 & ~n2194;
  assign n2298 = pi76  & n918;
  assign n2299 = pi74  & n1031;
  assign n2300 = pi75  & n913;
  assign n2301 = ~n2299 & ~n2300;
  assign n2302 = ~n2298 & n2301;
  assign n2303 = n881 & n921;
  assign n2304 = n2302 & ~n2303;
  assign n2305 = pi14  & ~n2304;
  assign n2306 = pi14  & ~n2305;
  assign n2307 = ~n2304 & ~n2305;
  assign n2308 = ~n2306 & ~n2307;
  assign n2309 = ~n2186 & ~n2188;
  assign n2310 = pi73  & n1269;
  assign n2311 = pi71  & n1340;
  assign n2312 = pi72  & n1264;
  assign n2313 = ~n2311 & ~n2312;
  assign n2314 = ~n2310 & n2313;
  assign n2315 = n639 & n1272;
  assign n2316 = n2314 & ~n2315;
  assign n2317 = pi17  & ~n2316;
  assign n2318 = pi17  & ~n2317;
  assign n2319 = ~n2316 & ~n2317;
  assign n2320 = ~n2318 & ~n2319;
  assign n2321 = pi67  & n2004;
  assign n2322 = pi65  & n2141;
  assign n2323 = pi66  & n1999;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~n2321 & n2324;
  assign n2326 = n313 & n2007;
  assign n2327 = n2325 & ~n2326;
  assign n2328 = pi23  & ~n2327;
  assign n2329 = pi23  & ~n2328;
  assign n2330 = ~n2327 & ~n2328;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = pi23  & ~pi24 ;
  assign n2333 = ~pi23  & pi24 ;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = pi64  & ~n2334;
  assign n2336 = n2153 & n2335;
  assign n2337 = ~n2153 & ~n2335;
  assign n2338 = ~n2336 & ~n2337;
  assign n2339 = ~n2331 & n2338;
  assign n2340 = n2331 & ~n2338;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = pi70  & n1582;
  assign n2343 = pi68  & n1713;
  assign n2344 = pi69  & n1577;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = ~n2342 & n2345;
  assign n2347 = n430 & n1585;
  assign n2348 = n2346 & ~n2347;
  assign n2349 = pi20  & ~n2348;
  assign n2350 = pi20  & ~n2349;
  assign n2351 = ~n2348 & ~n2349;
  assign n2352 = ~n2350 & ~n2351;
  assign n2353 = n2341 & ~n2352;
  assign n2354 = ~n2341 & n2352;
  assign n2355 = ~n2353 & ~n2354;
  assign n2356 = ~n2171 & n2355;
  assign n2357 = n2171 & ~n2355;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = ~n2320 & n2358;
  assign n2360 = n2320 & ~n2358;
  assign n2361 = ~n2359 & ~n2360;
  assign n2362 = ~n2309 & n2361;
  assign n2363 = n2309 & ~n2361;
  assign n2364 = ~n2362 & ~n2363;
  assign n2365 = n2308 & ~n2364;
  assign n2366 = ~n2308 & n2364;
  assign n2367 = ~n2365 & ~n2366;
  assign n2368 = ~n2297 & n2367;
  assign n2369 = n2297 & ~n2367;
  assign n2370 = ~n2368 & ~n2369;
  assign n2371 = pi79  & n675;
  assign n2372 = pi77  & n769;
  assign n2373 = pi78  & n670;
  assign n2374 = ~n2372 & ~n2373;
  assign n2375 = ~n2371 & n2374;
  assign n2376 = n678 & n1105;
  assign n2377 = n2375 & ~n2376;
  assign n2378 = pi11  & ~n2377;
  assign n2379 = pi11  & ~n2378;
  assign n2380 = ~n2377 & ~n2378;
  assign n2381 = ~n2379 & ~n2380;
  assign n2382 = n2370 & ~n2381;
  assign n2383 = n2370 & ~n2382;
  assign n2384 = ~n2381 & ~n2382;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = ~n2208 & ~n2213;
  assign n2387 = n2385 & n2386;
  assign n2388 = ~n2385 & ~n2386;
  assign n2389 = ~n2387 & ~n2388;
  assign n2390 = pi82  & n493;
  assign n2391 = pi80  & n533;
  assign n2392 = pi81  & n488;
  assign n2393 = ~n2391 & ~n2392;
  assign n2394 = ~n2390 & n2393;
  assign n2395 = n496 & n1532;
  assign n2396 = n2394 & ~n2395;
  assign n2397 = pi8  & ~n2396;
  assign n2398 = pi8  & ~n2397;
  assign n2399 = ~n2396 & ~n2397;
  assign n2400 = ~n2398 & ~n2399;
  assign n2401 = ~n2389 & n2400;
  assign n2402 = n2389 & ~n2400;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = ~n2296 & n2403;
  assign n2405 = n2296 & ~n2403;
  assign n2406 = ~n2404 & ~n2405;
  assign n2407 = ~n2295 & n2406;
  assign n2408 = ~n2295 & ~n2407;
  assign n2409 = n2406 & ~n2407;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = ~n2284 & ~n2410;
  assign n2412 = n2284 & n2410;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = ~n2283 & n2413;
  assign n2415 = n2283 & ~n2413;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = ~n2265 & n2416;
  assign n2418 = n2265 & ~n2416;
  assign po24  = ~n2417 & ~n2418;
  assign n2420 = ~n2414 & ~n2417;
  assign n2421 = pi89  & n264;
  assign n2422 = pi87  & n281;
  assign n2423 = pi88  & n259;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = ~n2421 & n2424;
  assign n2426 = ~n2273 & ~n2275;
  assign n2427 = ~pi88  & ~pi89 ;
  assign n2428 = pi88  & pi89 ;
  assign n2429 = ~n2427 & ~n2428;
  assign n2430 = ~n2426 & n2429;
  assign n2431 = n2426 & ~n2429;
  assign n2432 = ~n2430 & ~n2431;
  assign n2433 = n267 & n2432;
  assign n2434 = n2425 & ~n2433;
  assign n2435 = pi2  & ~n2434;
  assign n2436 = pi2  & ~n2435;
  assign n2437 = ~n2434 & ~n2435;
  assign n2438 = ~n2436 & ~n2437;
  assign n2439 = ~n2407 & ~n2411;
  assign n2440 = pi86  & n340;
  assign n2441 = pi84  & n380;
  assign n2442 = pi85  & n335;
  assign n2443 = ~n2441 & ~n2442;
  assign n2444 = ~n2440 & n2443;
  assign n2445 = n343 & n2099;
  assign n2446 = n2444 & ~n2445;
  assign n2447 = pi5  & ~n2446;
  assign n2448 = pi5  & ~n2447;
  assign n2449 = ~n2446 & ~n2447;
  assign n2450 = ~n2448 & ~n2449;
  assign n2451 = ~n2402 & ~n2404;
  assign n2452 = ~n2359 & ~n2362;
  assign n2453 = ~n2353 & ~n2356;
  assign n2454 = pi71  & n1582;
  assign n2455 = pi69  & n1713;
  assign n2456 = pi70  & n1577;
  assign n2457 = ~n2455 & ~n2456;
  assign n2458 = ~n2454 & n2457;
  assign n2459 = n476 & n1585;
  assign n2460 = n2458 & ~n2459;
  assign n2461 = pi20  & ~n2460;
  assign n2462 = pi20  & ~n2461;
  assign n2463 = ~n2460 & ~n2461;
  assign n2464 = ~n2462 & ~n2463;
  assign n2465 = ~n2336 & ~n2339;
  assign n2466 = pi68  & n2004;
  assign n2467 = pi66  & n2141;
  assign n2468 = pi67  & n1999;
  assign n2469 = ~n2467 & ~n2468;
  assign n2470 = ~n2466 & n2469;
  assign n2471 = n364 & n2007;
  assign n2472 = n2470 & ~n2471;
  assign n2473 = pi23  & ~n2472;
  assign n2474 = pi23  & ~n2473;
  assign n2475 = ~n2472 & ~n2473;
  assign n2476 = ~n2474 & ~n2475;
  assign n2477 = pi26  & ~n2335;
  assign n2478 = ~pi24  & pi25 ;
  assign n2479 = pi24  & ~pi25 ;
  assign n2480 = ~n2478 & ~n2479;
  assign n2481 = n2334 & ~n2480;
  assign n2482 = pi64  & n2481;
  assign n2483 = ~pi25  & pi26 ;
  assign n2484 = pi25  & ~pi26 ;
  assign n2485 = ~n2483 & ~n2484;
  assign n2486 = ~n2334 & n2485;
  assign n2487 = pi65  & n2486;
  assign n2488 = ~n2482 & ~n2487;
  assign n2489 = ~n2334 & ~n2485;
  assign n2490 = n270 & n2489;
  assign n2491 = n2488 & ~n2490;
  assign n2492 = pi26  & ~n2491;
  assign n2493 = pi26  & ~n2492;
  assign n2494 = ~n2491 & ~n2492;
  assign n2495 = ~n2493 & ~n2494;
  assign n2496 = n2477 & ~n2495;
  assign n2497 = ~n2477 & n2495;
  assign n2498 = ~n2496 & ~n2497;
  assign n2499 = ~n2476 & n2498;
  assign n2500 = n2476 & ~n2498;
  assign n2501 = ~n2499 & ~n2500;
  assign n2502 = ~n2465 & n2501;
  assign n2503 = n2465 & ~n2501;
  assign n2504 = ~n2502 & ~n2503;
  assign n2505 = ~n2464 & n2504;
  assign n2506 = n2464 & ~n2504;
  assign n2507 = ~n2505 & ~n2506;
  assign n2508 = ~n2453 & n2507;
  assign n2509 = n2453 & ~n2507;
  assign n2510 = ~n2508 & ~n2509;
  assign n2511 = pi74  & n1269;
  assign n2512 = pi72  & n1340;
  assign n2513 = pi73  & n1264;
  assign n2514 = ~n2512 & ~n2513;
  assign n2515 = ~n2511 & n2514;
  assign n2516 = n722 & n1272;
  assign n2517 = n2515 & ~n2516;
  assign n2518 = pi17  & ~n2517;
  assign n2519 = pi17  & ~n2518;
  assign n2520 = ~n2517 & ~n2518;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = n2510 & ~n2521;
  assign n2523 = ~n2510 & n2521;
  assign n2524 = ~n2522 & ~n2523;
  assign n2525 = n2452 & ~n2524;
  assign n2526 = ~n2452 & n2524;
  assign n2527 = ~n2525 & ~n2526;
  assign n2528 = pi77  & n918;
  assign n2529 = pi75  & n1031;
  assign n2530 = pi76  & n913;
  assign n2531 = ~n2529 & ~n2530;
  assign n2532 = ~n2528 & n2531;
  assign n2533 = n921 & n984;
  assign n2534 = n2532 & ~n2533;
  assign n2535 = pi14  & ~n2534;
  assign n2536 = pi14  & ~n2535;
  assign n2537 = ~n2534 & ~n2535;
  assign n2538 = ~n2536 & ~n2537;
  assign n2539 = ~n2527 & n2538;
  assign n2540 = n2527 & ~n2538;
  assign n2541 = ~n2539 & ~n2540;
  assign n2542 = ~n2366 & ~n2368;
  assign n2543 = n2541 & ~n2542;
  assign n2544 = ~n2541 & n2542;
  assign n2545 = ~n2543 & ~n2544;
  assign n2546 = pi80  & n675;
  assign n2547 = pi78  & n769;
  assign n2548 = pi79  & n670;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = ~n2546 & n2549;
  assign n2551 = n678 & n1205;
  assign n2552 = n2550 & ~n2551;
  assign n2553 = pi11  & ~n2552;
  assign n2554 = pi11  & ~n2553;
  assign n2555 = ~n2552 & ~n2553;
  assign n2556 = ~n2554 & ~n2555;
  assign n2557 = n2545 & ~n2556;
  assign n2558 = n2545 & ~n2557;
  assign n2559 = ~n2556 & ~n2557;
  assign n2560 = ~n2558 & ~n2559;
  assign n2561 = ~n2382 & ~n2388;
  assign n2562 = n2560 & n2561;
  assign n2563 = ~n2560 & ~n2561;
  assign n2564 = ~n2562 & ~n2563;
  assign n2565 = pi83  & n493;
  assign n2566 = pi81  & n533;
  assign n2567 = pi82  & n488;
  assign n2568 = ~n2566 & ~n2567;
  assign n2569 = ~n2565 & n2568;
  assign n2570 = n496 & n1672;
  assign n2571 = n2569 & ~n2570;
  assign n2572 = pi8  & ~n2571;
  assign n2573 = pi8  & ~n2572;
  assign n2574 = ~n2571 & ~n2572;
  assign n2575 = ~n2573 & ~n2574;
  assign n2576 = n2564 & ~n2575;
  assign n2577 = ~n2564 & n2575;
  assign n2578 = ~n2576 & ~n2577;
  assign n2579 = ~n2451 & n2578;
  assign n2580 = n2451 & ~n2578;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = n2450 & n2581;
  assign n2583 = ~n2450 & ~n2581;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = ~n2439 & ~n2584;
  assign n2586 = n2439 & n2584;
  assign n2587 = ~n2585 & ~n2586;
  assign n2588 = ~n2438 & n2587;
  assign n2589 = n2438 & ~n2587;
  assign n2590 = ~n2588 & ~n2589;
  assign n2591 = ~n2420 & n2590;
  assign n2592 = n2420 & ~n2590;
  assign po25  = ~n2591 & ~n2592;
  assign n2594 = ~n2588 & ~n2591;
  assign n2595 = pi90  & n264;
  assign n2596 = pi88  & n281;
  assign n2597 = pi89  & n259;
  assign n2598 = ~n2596 & ~n2597;
  assign n2599 = ~n2595 & n2598;
  assign n2600 = ~n2428 & ~n2430;
  assign n2601 = ~pi89  & ~pi90 ;
  assign n2602 = pi89  & pi90 ;
  assign n2603 = ~n2601 & ~n2602;
  assign n2604 = ~n2600 & n2603;
  assign n2605 = n2600 & ~n2603;
  assign n2606 = ~n2604 & ~n2605;
  assign n2607 = n267 & n2606;
  assign n2608 = n2599 & ~n2607;
  assign n2609 = pi2  & ~n2608;
  assign n2610 = pi2  & ~n2609;
  assign n2611 = ~n2608 & ~n2609;
  assign n2612 = ~n2610 & ~n2611;
  assign n2613 = ~n2450 & n2581;
  assign n2614 = ~n2585 & ~n2613;
  assign n2615 = ~n2557 & ~n2563;
  assign n2616 = pi81  & n675;
  assign n2617 = pi79  & n769;
  assign n2618 = pi80  & n670;
  assign n2619 = ~n2617 & ~n2618;
  assign n2620 = ~n2616 & n2619;
  assign n2621 = n678 & n1413;
  assign n2622 = n2620 & ~n2621;
  assign n2623 = pi11  & ~n2622;
  assign n2624 = pi11  & ~n2623;
  assign n2625 = ~n2622 & ~n2623;
  assign n2626 = ~n2624 & ~n2625;
  assign n2627 = ~n2540 & ~n2543;
  assign n2628 = ~n2522 & ~n2526;
  assign n2629 = pi75  & n1269;
  assign n2630 = pi73  & n1340;
  assign n2631 = pi74  & n1264;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = ~n2629 & n2632;
  assign n2634 = n747 & n1272;
  assign n2635 = n2633 & ~n2634;
  assign n2636 = pi17  & ~n2635;
  assign n2637 = pi17  & ~n2636;
  assign n2638 = ~n2635 & ~n2636;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = ~n2505 & ~n2508;
  assign n2641 = ~n2499 & ~n2502;
  assign n2642 = pi66  & n2486;
  assign n2643 = n2334 & ~n2485;
  assign n2644 = n2480 & n2643;
  assign n2645 = pi64  & n2644;
  assign n2646 = pi65  & n2481;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = ~n2642 & n2647;
  assign n2649 = n291 & n2489;
  assign n2650 = n2648 & ~n2649;
  assign n2651 = pi26  & ~n2650;
  assign n2652 = pi26  & ~n2651;
  assign n2653 = ~n2650 & ~n2651;
  assign n2654 = ~n2652 & ~n2653;
  assign n2655 = ~n2496 & n2654;
  assign n2656 = n2496 & ~n2654;
  assign n2657 = ~n2655 & ~n2656;
  assign n2658 = pi69  & n2004;
  assign n2659 = pi67  & n2141;
  assign n2660 = pi68  & n1999;
  assign n2661 = ~n2659 & ~n2660;
  assign n2662 = ~n2658 & n2661;
  assign n2663 = n405 & n2007;
  assign n2664 = n2662 & ~n2663;
  assign n2665 = pi23  & ~n2664;
  assign n2666 = pi23  & ~n2665;
  assign n2667 = ~n2664 & ~n2665;
  assign n2668 = ~n2666 & ~n2667;
  assign n2669 = n2657 & ~n2668;
  assign n2670 = ~n2657 & n2668;
  assign n2671 = ~n2641 & ~n2670;
  assign n2672 = ~n2669 & n2671;
  assign n2673 = ~n2641 & ~n2672;
  assign n2674 = ~n2669 & ~n2672;
  assign n2675 = ~n2670 & n2674;
  assign n2676 = ~n2673 & ~n2675;
  assign n2677 = pi72  & n1582;
  assign n2678 = pi70  & n1713;
  assign n2679 = pi71  & n1577;
  assign n2680 = ~n2678 & ~n2679;
  assign n2681 = ~n2677 & n2680;
  assign n2682 = n575 & n1585;
  assign n2683 = n2681 & ~n2682;
  assign n2684 = pi20  & ~n2683;
  assign n2685 = pi20  & ~n2684;
  assign n2686 = ~n2683 & ~n2684;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = n2676 & n2687;
  assign n2689 = ~n2676 & ~n2687;
  assign n2690 = ~n2688 & ~n2689;
  assign n2691 = ~n2640 & n2690;
  assign n2692 = n2640 & ~n2690;
  assign n2693 = ~n2691 & ~n2692;
  assign n2694 = n2639 & ~n2693;
  assign n2695 = ~n2639 & n2693;
  assign n2696 = ~n2694 & ~n2695;
  assign n2697 = ~n2628 & n2696;
  assign n2698 = n2628 & ~n2696;
  assign n2699 = ~n2697 & ~n2698;
  assign n2700 = pi78  & n918;
  assign n2701 = pi76  & n1031;
  assign n2702 = pi77  & n913;
  assign n2703 = ~n2701 & ~n2702;
  assign n2704 = ~n2700 & n2703;
  assign n2705 = n921 & n1009;
  assign n2706 = n2704 & ~n2705;
  assign n2707 = pi14  & ~n2706;
  assign n2708 = pi14  & ~n2707;
  assign n2709 = ~n2706 & ~n2707;
  assign n2710 = ~n2708 & ~n2709;
  assign n2711 = n2699 & ~n2710;
  assign n2712 = n2699 & ~n2711;
  assign n2713 = ~n2710 & ~n2711;
  assign n2714 = ~n2712 & ~n2713;
  assign n2715 = ~n2627 & ~n2714;
  assign n2716 = n2627 & n2714;
  assign n2717 = ~n2715 & ~n2716;
  assign n2718 = ~n2626 & n2717;
  assign n2719 = n2626 & ~n2717;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = n2615 & ~n2720;
  assign n2722 = ~n2615 & n2720;
  assign n2723 = ~n2721 & ~n2722;
  assign n2724 = pi84  & n493;
  assign n2725 = pi82  & n533;
  assign n2726 = pi83  & n488;
  assign n2727 = ~n2725 & ~n2726;
  assign n2728 = ~n2724 & n2727;
  assign n2729 = n496 & n1805;
  assign n2730 = n2728 & ~n2729;
  assign n2731 = pi8  & ~n2730;
  assign n2732 = pi8  & ~n2731;
  assign n2733 = ~n2730 & ~n2731;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = n2723 & ~n2734;
  assign n2736 = n2723 & ~n2735;
  assign n2737 = ~n2734 & ~n2735;
  assign n2738 = ~n2736 & ~n2737;
  assign n2739 = ~n2576 & ~n2579;
  assign n2740 = n2738 & n2739;
  assign n2741 = ~n2738 & ~n2739;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = pi87  & n340;
  assign n2744 = pi85  & n380;
  assign n2745 = pi86  & n335;
  assign n2746 = ~n2744 & ~n2745;
  assign n2747 = ~n2743 & n2746;
  assign n2748 = n343 & n2252;
  assign n2749 = n2747 & ~n2748;
  assign n2750 = pi5  & ~n2749;
  assign n2751 = pi5  & ~n2750;
  assign n2752 = ~n2749 & ~n2750;
  assign n2753 = ~n2751 & ~n2752;
  assign n2754 = n2742 & ~n2753;
  assign n2755 = ~n2742 & n2753;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = ~n2614 & n2756;
  assign n2758 = n2614 & ~n2756;
  assign n2759 = ~n2757 & ~n2758;
  assign n2760 = ~n2612 & n2759;
  assign n2761 = n2612 & ~n2759;
  assign n2762 = ~n2760 & ~n2761;
  assign n2763 = ~n2594 & n2762;
  assign n2764 = n2594 & ~n2762;
  assign po26  = ~n2763 & ~n2764;
  assign n2766 = ~n2760 & ~n2763;
  assign n2767 = ~n2718 & ~n2722;
  assign n2768 = ~n2695 & ~n2697;
  assign n2769 = pi76  & n1269;
  assign n2770 = pi74  & n1340;
  assign n2771 = pi75  & n1264;
  assign n2772 = ~n2770 & ~n2771;
  assign n2773 = ~n2769 & n2772;
  assign n2774 = n881 & n1272;
  assign n2775 = n2773 & ~n2774;
  assign n2776 = pi17  & ~n2775;
  assign n2777 = pi17  & ~n2776;
  assign n2778 = ~n2775 & ~n2776;
  assign n2779 = ~n2777 & ~n2778;
  assign n2780 = ~n2689 & ~n2691;
  assign n2781 = pi73  & n1582;
  assign n2782 = pi71  & n1713;
  assign n2783 = pi72  & n1577;
  assign n2784 = ~n2782 & ~n2783;
  assign n2785 = ~n2781 & n2784;
  assign n2786 = n639 & n1585;
  assign n2787 = n2785 & ~n2786;
  assign n2788 = pi20  & ~n2787;
  assign n2789 = pi20  & ~n2788;
  assign n2790 = ~n2787 & ~n2788;
  assign n2791 = ~n2789 & ~n2790;
  assign n2792 = pi67  & n2486;
  assign n2793 = pi65  & n2644;
  assign n2794 = pi66  & n2481;
  assign n2795 = ~n2793 & ~n2794;
  assign n2796 = ~n2792 & n2795;
  assign n2797 = n313 & n2489;
  assign n2798 = n2796 & ~n2797;
  assign n2799 = pi26  & ~n2798;
  assign n2800 = pi26  & ~n2799;
  assign n2801 = ~n2798 & ~n2799;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = pi26  & ~pi27 ;
  assign n2804 = ~pi26  & pi27 ;
  assign n2805 = ~n2803 & ~n2804;
  assign n2806 = pi64  & ~n2805;
  assign n2807 = n2656 & n2806;
  assign n2808 = ~n2656 & ~n2806;
  assign n2809 = ~n2807 & ~n2808;
  assign n2810 = ~n2802 & n2809;
  assign n2811 = n2802 & ~n2809;
  assign n2812 = ~n2810 & ~n2811;
  assign n2813 = pi70  & n2004;
  assign n2814 = pi68  & n2141;
  assign n2815 = pi69  & n1999;
  assign n2816 = ~n2814 & ~n2815;
  assign n2817 = ~n2813 & n2816;
  assign n2818 = n430 & n2007;
  assign n2819 = n2817 & ~n2818;
  assign n2820 = pi23  & ~n2819;
  assign n2821 = pi23  & ~n2820;
  assign n2822 = ~n2819 & ~n2820;
  assign n2823 = ~n2821 & ~n2822;
  assign n2824 = n2812 & ~n2823;
  assign n2825 = ~n2812 & n2823;
  assign n2826 = ~n2824 & ~n2825;
  assign n2827 = ~n2674 & n2826;
  assign n2828 = n2674 & ~n2826;
  assign n2829 = ~n2827 & ~n2828;
  assign n2830 = ~n2791 & n2829;
  assign n2831 = n2791 & ~n2829;
  assign n2832 = ~n2830 & ~n2831;
  assign n2833 = ~n2780 & n2832;
  assign n2834 = n2780 & ~n2832;
  assign n2835 = ~n2833 & ~n2834;
  assign n2836 = n2779 & ~n2835;
  assign n2837 = ~n2779 & n2835;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = ~n2768 & n2838;
  assign n2840 = n2768 & ~n2838;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = pi79  & n918;
  assign n2843 = pi77  & n1031;
  assign n2844 = pi78  & n913;
  assign n2845 = ~n2843 & ~n2844;
  assign n2846 = ~n2842 & n2845;
  assign n2847 = n921 & n1105;
  assign n2848 = n2846 & ~n2847;
  assign n2849 = pi14  & ~n2848;
  assign n2850 = pi14  & ~n2849;
  assign n2851 = ~n2848 & ~n2849;
  assign n2852 = ~n2850 & ~n2851;
  assign n2853 = n2841 & ~n2852;
  assign n2854 = n2841 & ~n2853;
  assign n2855 = ~n2852 & ~n2853;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857 = ~n2711 & ~n2715;
  assign n2858 = n2856 & n2857;
  assign n2859 = ~n2856 & ~n2857;
  assign n2860 = ~n2858 & ~n2859;
  assign n2861 = pi82  & n675;
  assign n2862 = pi80  & n769;
  assign n2863 = pi81  & n670;
  assign n2864 = ~n2862 & ~n2863;
  assign n2865 = ~n2861 & n2864;
  assign n2866 = n678 & n1532;
  assign n2867 = n2865 & ~n2866;
  assign n2868 = pi11  & ~n2867;
  assign n2869 = pi11  & ~n2868;
  assign n2870 = ~n2867 & ~n2868;
  assign n2871 = ~n2869 & ~n2870;
  assign n2872 = n2860 & ~n2871;
  assign n2873 = ~n2860 & n2871;
  assign n2874 = ~n2872 & ~n2873;
  assign n2875 = n2767 & ~n2874;
  assign n2876 = ~n2767 & n2874;
  assign n2877 = ~n2875 & ~n2876;
  assign n2878 = pi85  & n493;
  assign n2879 = pi83  & n533;
  assign n2880 = pi84  & n488;
  assign n2881 = ~n2879 & ~n2880;
  assign n2882 = ~n2878 & n2881;
  assign n2883 = n496 & n1943;
  assign n2884 = n2882 & ~n2883;
  assign n2885 = pi8  & ~n2884;
  assign n2886 = pi8  & ~n2885;
  assign n2887 = ~n2884 & ~n2885;
  assign n2888 = ~n2886 & ~n2887;
  assign n2889 = ~n2877 & n2888;
  assign n2890 = n2877 & ~n2888;
  assign n2891 = ~n2889 & ~n2890;
  assign n2892 = ~n2735 & ~n2741;
  assign n2893 = n2891 & ~n2892;
  assign n2894 = ~n2891 & n2892;
  assign n2895 = ~n2893 & ~n2894;
  assign n2896 = pi88  & n340;
  assign n2897 = pi86  & n380;
  assign n2898 = pi87  & n335;
  assign n2899 = ~n2897 & ~n2898;
  assign n2900 = ~n2896 & n2899;
  assign n2901 = n343 & n2277;
  assign n2902 = n2900 & ~n2901;
  assign n2903 = pi5  & ~n2902;
  assign n2904 = pi5  & ~n2903;
  assign n2905 = ~n2902 & ~n2903;
  assign n2906 = ~n2904 & ~n2905;
  assign n2907 = n2895 & ~n2906;
  assign n2908 = n2895 & ~n2907;
  assign n2909 = ~n2906 & ~n2907;
  assign n2910 = ~n2908 & ~n2909;
  assign n2911 = ~n2754 & ~n2757;
  assign n2912 = n2910 & n2911;
  assign n2913 = ~n2910 & ~n2911;
  assign n2914 = ~n2912 & ~n2913;
  assign n2915 = pi91  & n264;
  assign n2916 = pi89  & n281;
  assign n2917 = pi90  & n259;
  assign n2918 = ~n2916 & ~n2917;
  assign n2919 = ~n2915 & n2918;
  assign n2920 = ~n2602 & ~n2604;
  assign n2921 = ~pi90  & ~pi91 ;
  assign n2922 = pi90  & pi91 ;
  assign n2923 = ~n2921 & ~n2922;
  assign n2924 = ~n2920 & n2923;
  assign n2925 = n2920 & ~n2923;
  assign n2926 = ~n2924 & ~n2925;
  assign n2927 = n267 & n2926;
  assign n2928 = n2919 & ~n2927;
  assign n2929 = pi2  & ~n2928;
  assign n2930 = pi2  & ~n2929;
  assign n2931 = ~n2928 & ~n2929;
  assign n2932 = ~n2930 & ~n2931;
  assign n2933 = ~n2914 & n2932;
  assign n2934 = n2914 & ~n2932;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = ~n2766 & n2935;
  assign n2937 = n2766 & ~n2935;
  assign po27  = ~n2936 & ~n2937;
  assign n2939 = ~n2934 & ~n2936;
  assign n2940 = ~n2872 & ~n2876;
  assign n2941 = ~n2837 & ~n2839;
  assign n2942 = ~n2830 & ~n2833;
  assign n2943 = ~n2824 & ~n2827;
  assign n2944 = pi71  & n2004;
  assign n2945 = pi69  & n2141;
  assign n2946 = pi70  & n1999;
  assign n2947 = ~n2945 & ~n2946;
  assign n2948 = ~n2944 & n2947;
  assign n2949 = n476 & n2007;
  assign n2950 = n2948 & ~n2949;
  assign n2951 = pi23  & ~n2950;
  assign n2952 = pi23  & ~n2951;
  assign n2953 = ~n2950 & ~n2951;
  assign n2954 = ~n2952 & ~n2953;
  assign n2955 = ~n2807 & ~n2810;
  assign n2956 = pi68  & n2486;
  assign n2957 = pi66  & n2644;
  assign n2958 = pi67  & n2481;
  assign n2959 = ~n2957 & ~n2958;
  assign n2960 = ~n2956 & n2959;
  assign n2961 = n364 & n2489;
  assign n2962 = n2960 & ~n2961;
  assign n2963 = pi26  & ~n2962;
  assign n2964 = pi26  & ~n2963;
  assign n2965 = ~n2962 & ~n2963;
  assign n2966 = ~n2964 & ~n2965;
  assign n2967 = pi29  & ~n2806;
  assign n2968 = ~pi27  & pi28 ;
  assign n2969 = pi27  & ~pi28 ;
  assign n2970 = ~n2968 & ~n2969;
  assign n2971 = n2805 & ~n2970;
  assign n2972 = pi64  & n2971;
  assign n2973 = ~pi28  & pi29 ;
  assign n2974 = pi28  & ~pi29 ;
  assign n2975 = ~n2973 & ~n2974;
  assign n2976 = ~n2805 & n2975;
  assign n2977 = pi65  & n2976;
  assign n2978 = ~n2972 & ~n2977;
  assign n2979 = ~n2805 & ~n2975;
  assign n2980 = n270 & n2979;
  assign n2981 = n2978 & ~n2980;
  assign n2982 = pi29  & ~n2981;
  assign n2983 = pi29  & ~n2982;
  assign n2984 = ~n2981 & ~n2982;
  assign n2985 = ~n2983 & ~n2984;
  assign n2986 = n2967 & ~n2985;
  assign n2987 = ~n2967 & n2985;
  assign n2988 = ~n2986 & ~n2987;
  assign n2989 = ~n2966 & n2988;
  assign n2990 = n2966 & ~n2988;
  assign n2991 = ~n2989 & ~n2990;
  assign n2992 = ~n2955 & n2991;
  assign n2993 = n2955 & ~n2991;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = ~n2954 & n2994;
  assign n2996 = n2954 & ~n2994;
  assign n2997 = ~n2995 & ~n2996;
  assign n2998 = ~n2943 & n2997;
  assign n2999 = n2943 & ~n2997;
  assign n3000 = ~n2998 & ~n2999;
  assign n3001 = pi74  & n1582;
  assign n3002 = pi72  & n1713;
  assign n3003 = pi73  & n1577;
  assign n3004 = ~n3002 & ~n3003;
  assign n3005 = ~n3001 & n3004;
  assign n3006 = n722 & n1585;
  assign n3007 = n3005 & ~n3006;
  assign n3008 = pi20  & ~n3007;
  assign n3009 = pi20  & ~n3008;
  assign n3010 = ~n3007 & ~n3008;
  assign n3011 = ~n3009 & ~n3010;
  assign n3012 = n3000 & ~n3011;
  assign n3013 = ~n3000 & n3011;
  assign n3014 = ~n3012 & ~n3013;
  assign n3015 = n2942 & ~n3014;
  assign n3016 = ~n2942 & n3014;
  assign n3017 = ~n3015 & ~n3016;
  assign n3018 = pi77  & n1269;
  assign n3019 = pi75  & n1340;
  assign n3020 = pi76  & n1264;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = ~n3018 & n3021;
  assign n3023 = n984 & n1272;
  assign n3024 = n3022 & ~n3023;
  assign n3025 = pi17  & ~n3024;
  assign n3026 = pi17  & ~n3025;
  assign n3027 = ~n3024 & ~n3025;
  assign n3028 = ~n3026 & ~n3027;
  assign n3029 = n3017 & ~n3028;
  assign n3030 = ~n3017 & n3028;
  assign n3031 = ~n3029 & ~n3030;
  assign n3032 = ~n2941 & n3031;
  assign n3033 = n2941 & ~n3031;
  assign n3034 = ~n3032 & ~n3033;
  assign n3035 = pi80  & n918;
  assign n3036 = pi78  & n1031;
  assign n3037 = pi79  & n913;
  assign n3038 = ~n3036 & ~n3037;
  assign n3039 = ~n3035 & n3038;
  assign n3040 = n921 & n1205;
  assign n3041 = n3039 & ~n3040;
  assign n3042 = pi14  & ~n3041;
  assign n3043 = pi14  & ~n3042;
  assign n3044 = ~n3041 & ~n3042;
  assign n3045 = ~n3043 & ~n3044;
  assign n3046 = n3034 & ~n3045;
  assign n3047 = n3034 & ~n3046;
  assign n3048 = ~n3045 & ~n3046;
  assign n3049 = ~n3047 & ~n3048;
  assign n3050 = ~n2853 & ~n2859;
  assign n3051 = n3049 & n3050;
  assign n3052 = ~n3049 & ~n3050;
  assign n3053 = ~n3051 & ~n3052;
  assign n3054 = pi83  & n675;
  assign n3055 = pi81  & n769;
  assign n3056 = pi82  & n670;
  assign n3057 = ~n3055 & ~n3056;
  assign n3058 = ~n3054 & n3057;
  assign n3059 = n678 & n1672;
  assign n3060 = n3058 & ~n3059;
  assign n3061 = pi11  & ~n3060;
  assign n3062 = pi11  & ~n3061;
  assign n3063 = ~n3060 & ~n3061;
  assign n3064 = ~n3062 & ~n3063;
  assign n3065 = n3053 & ~n3064;
  assign n3066 = ~n3053 & n3064;
  assign n3067 = ~n3065 & ~n3066;
  assign n3068 = n2940 & ~n3067;
  assign n3069 = ~n2940 & n3067;
  assign n3070 = ~n3068 & ~n3069;
  assign n3071 = pi86  & n493;
  assign n3072 = pi84  & n533;
  assign n3073 = pi85  & n488;
  assign n3074 = ~n3072 & ~n3073;
  assign n3075 = ~n3071 & n3074;
  assign n3076 = n496 & n2099;
  assign n3077 = n3075 & ~n3076;
  assign n3078 = pi8  & ~n3077;
  assign n3079 = pi8  & ~n3078;
  assign n3080 = ~n3077 & ~n3078;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = ~n3070 & n3081;
  assign n3083 = n3070 & ~n3081;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = ~n2890 & ~n2893;
  assign n3086 = n3084 & ~n3085;
  assign n3087 = ~n3084 & n3085;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = pi89  & n340;
  assign n3090 = pi87  & n380;
  assign n3091 = pi88  & n335;
  assign n3092 = ~n3090 & ~n3091;
  assign n3093 = ~n3089 & n3092;
  assign n3094 = n343 & n2432;
  assign n3095 = n3093 & ~n3094;
  assign n3096 = pi5  & ~n3095;
  assign n3097 = pi5  & ~n3096;
  assign n3098 = ~n3095 & ~n3096;
  assign n3099 = ~n3097 & ~n3098;
  assign n3100 = n3088 & ~n3099;
  assign n3101 = n3088 & ~n3100;
  assign n3102 = ~n3099 & ~n3100;
  assign n3103 = ~n3101 & ~n3102;
  assign n3104 = ~n2907 & ~n2913;
  assign n3105 = n3103 & n3104;
  assign n3106 = ~n3103 & ~n3104;
  assign n3107 = ~n3105 & ~n3106;
  assign n3108 = pi92  & n264;
  assign n3109 = pi90  & n281;
  assign n3110 = pi91  & n259;
  assign n3111 = ~n3109 & ~n3110;
  assign n3112 = ~n3108 & n3111;
  assign n3113 = ~n2922 & ~n2924;
  assign n3114 = ~pi91  & ~pi92 ;
  assign n3115 = pi91  & pi92 ;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = ~n3113 & n3116;
  assign n3118 = n3113 & ~n3116;
  assign n3119 = ~n3117 & ~n3118;
  assign n3120 = n267 & n3119;
  assign n3121 = n3112 & ~n3120;
  assign n3122 = pi2  & ~n3121;
  assign n3123 = pi2  & ~n3122;
  assign n3124 = ~n3121 & ~n3122;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = ~n3107 & n3125;
  assign n3127 = n3107 & ~n3125;
  assign n3128 = ~n3126 & ~n3127;
  assign n3129 = ~n2939 & n3128;
  assign n3130 = n2939 & ~n3128;
  assign po28  = ~n3129 & ~n3130;
  assign n3132 = ~n3127 & ~n3129;
  assign n3133 = pi93  & n264;
  assign n3134 = pi91  & n281;
  assign n3135 = pi92  & n259;
  assign n3136 = ~n3134 & ~n3135;
  assign n3137 = ~n3133 & n3136;
  assign n3138 = ~n3115 & ~n3117;
  assign n3139 = ~pi92  & ~pi93 ;
  assign n3140 = pi92  & pi93 ;
  assign n3141 = ~n3139 & ~n3140;
  assign n3142 = ~n3138 & n3141;
  assign n3143 = n3138 & ~n3141;
  assign n3144 = ~n3142 & ~n3143;
  assign n3145 = n267 & n3144;
  assign n3146 = n3137 & ~n3145;
  assign n3147 = pi2  & ~n3146;
  assign n3148 = pi2  & ~n3147;
  assign n3149 = ~n3146 & ~n3147;
  assign n3150 = ~n3148 & ~n3149;
  assign n3151 = ~n3100 & ~n3106;
  assign n3152 = pi90  & n340;
  assign n3153 = pi88  & n380;
  assign n3154 = pi89  & n335;
  assign n3155 = ~n3153 & ~n3154;
  assign n3156 = ~n3152 & n3155;
  assign n3157 = n343 & n2606;
  assign n3158 = n3156 & ~n3157;
  assign n3159 = pi5  & ~n3158;
  assign n3160 = pi5  & ~n3159;
  assign n3161 = ~n3158 & ~n3159;
  assign n3162 = ~n3160 & ~n3161;
  assign n3163 = ~n3083 & ~n3086;
  assign n3164 = ~n3065 & ~n3069;
  assign n3165 = ~n3046 & ~n3052;
  assign n3166 = ~n3012 & ~n3016;
  assign n3167 = pi75  & n1582;
  assign n3168 = pi73  & n1713;
  assign n3169 = pi74  & n1577;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = ~n3167 & n3170;
  assign n3172 = n747 & n1585;
  assign n3173 = n3171 & ~n3172;
  assign n3174 = pi20  & ~n3173;
  assign n3175 = pi20  & ~n3174;
  assign n3176 = ~n3173 & ~n3174;
  assign n3177 = ~n3175 & ~n3176;
  assign n3178 = ~n2995 & ~n2998;
  assign n3179 = ~n2989 & ~n2992;
  assign n3180 = pi66  & n2976;
  assign n3181 = n2805 & ~n2975;
  assign n3182 = n2970 & n3181;
  assign n3183 = pi64  & n3182;
  assign n3184 = pi65  & n2971;
  assign n3185 = ~n3183 & ~n3184;
  assign n3186 = ~n3180 & n3185;
  assign n3187 = n291 & n2979;
  assign n3188 = n3186 & ~n3187;
  assign n3189 = pi29  & ~n3188;
  assign n3190 = pi29  & ~n3189;
  assign n3191 = ~n3188 & ~n3189;
  assign n3192 = ~n3190 & ~n3191;
  assign n3193 = ~n2986 & n3192;
  assign n3194 = n2986 & ~n3192;
  assign n3195 = ~n3193 & ~n3194;
  assign n3196 = pi69  & n2486;
  assign n3197 = pi67  & n2644;
  assign n3198 = pi68  & n2481;
  assign n3199 = ~n3197 & ~n3198;
  assign n3200 = ~n3196 & n3199;
  assign n3201 = n405 & n2489;
  assign n3202 = n3200 & ~n3201;
  assign n3203 = pi26  & ~n3202;
  assign n3204 = pi26  & ~n3203;
  assign n3205 = ~n3202 & ~n3203;
  assign n3206 = ~n3204 & ~n3205;
  assign n3207 = n3195 & ~n3206;
  assign n3208 = ~n3195 & n3206;
  assign n3209 = ~n3179 & ~n3208;
  assign n3210 = ~n3207 & n3209;
  assign n3211 = ~n3179 & ~n3210;
  assign n3212 = ~n3207 & ~n3210;
  assign n3213 = ~n3208 & n3212;
  assign n3214 = ~n3211 & ~n3213;
  assign n3215 = pi72  & n2004;
  assign n3216 = pi70  & n2141;
  assign n3217 = pi71  & n1999;
  assign n3218 = ~n3216 & ~n3217;
  assign n3219 = ~n3215 & n3218;
  assign n3220 = n575 & n2007;
  assign n3221 = n3219 & ~n3220;
  assign n3222 = pi23  & ~n3221;
  assign n3223 = pi23  & ~n3222;
  assign n3224 = ~n3221 & ~n3222;
  assign n3225 = ~n3223 & ~n3224;
  assign n3226 = n3214 & n3225;
  assign n3227 = ~n3214 & ~n3225;
  assign n3228 = ~n3226 & ~n3227;
  assign n3229 = ~n3178 & n3228;
  assign n3230 = n3178 & ~n3228;
  assign n3231 = ~n3229 & ~n3230;
  assign n3232 = n3177 & ~n3231;
  assign n3233 = ~n3177 & n3231;
  assign n3234 = ~n3232 & ~n3233;
  assign n3235 = ~n3166 & n3234;
  assign n3236 = n3166 & ~n3234;
  assign n3237 = ~n3235 & ~n3236;
  assign n3238 = pi78  & n1269;
  assign n3239 = pi76  & n1340;
  assign n3240 = pi77  & n1264;
  assign n3241 = ~n3239 & ~n3240;
  assign n3242 = ~n3238 & n3241;
  assign n3243 = n1009 & n1272;
  assign n3244 = n3242 & ~n3243;
  assign n3245 = pi17  & ~n3244;
  assign n3246 = pi17  & ~n3245;
  assign n3247 = ~n3244 & ~n3245;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = n3237 & ~n3248;
  assign n3250 = n3237 & ~n3249;
  assign n3251 = ~n3248 & ~n3249;
  assign n3252 = ~n3250 & ~n3251;
  assign n3253 = ~n3029 & ~n3032;
  assign n3254 = n3252 & n3253;
  assign n3255 = ~n3252 & ~n3253;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = pi81  & n918;
  assign n3258 = pi79  & n1031;
  assign n3259 = pi80  & n913;
  assign n3260 = ~n3258 & ~n3259;
  assign n3261 = ~n3257 & n3260;
  assign n3262 = n921 & n1413;
  assign n3263 = n3261 & ~n3262;
  assign n3264 = pi14  & ~n3263;
  assign n3265 = pi14  & ~n3264;
  assign n3266 = ~n3263 & ~n3264;
  assign n3267 = ~n3265 & ~n3266;
  assign n3268 = n3256 & ~n3267;
  assign n3269 = ~n3256 & n3267;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = n3165 & ~n3270;
  assign n3272 = ~n3165 & n3270;
  assign n3273 = ~n3271 & ~n3272;
  assign n3274 = pi84  & n675;
  assign n3275 = pi82  & n769;
  assign n3276 = pi83  & n670;
  assign n3277 = ~n3275 & ~n3276;
  assign n3278 = ~n3274 & n3277;
  assign n3279 = n678 & n1805;
  assign n3280 = n3278 & ~n3279;
  assign n3281 = pi11  & ~n3280;
  assign n3282 = pi11  & ~n3281;
  assign n3283 = ~n3280 & ~n3281;
  assign n3284 = ~n3282 & ~n3283;
  assign n3285 = n3273 & ~n3284;
  assign n3286 = ~n3273 & n3284;
  assign n3287 = ~n3164 & ~n3286;
  assign n3288 = ~n3285 & n3287;
  assign n3289 = ~n3164 & ~n3288;
  assign n3290 = ~n3285 & ~n3288;
  assign n3291 = ~n3286 & n3290;
  assign n3292 = ~n3289 & ~n3291;
  assign n3293 = pi87  & n493;
  assign n3294 = pi85  & n533;
  assign n3295 = pi86  & n488;
  assign n3296 = ~n3294 & ~n3295;
  assign n3297 = ~n3293 & n3296;
  assign n3298 = n496 & n2252;
  assign n3299 = n3297 & ~n3298;
  assign n3300 = pi8  & ~n3299;
  assign n3301 = pi8  & ~n3300;
  assign n3302 = ~n3299 & ~n3300;
  assign n3303 = ~n3301 & ~n3302;
  assign n3304 = ~n3292 & ~n3303;
  assign n3305 = n3292 & n3303;
  assign n3306 = ~n3304 & ~n3305;
  assign n3307 = ~n3163 & n3306;
  assign n3308 = n3163 & ~n3306;
  assign n3309 = ~n3307 & ~n3308;
  assign n3310 = ~n3162 & n3309;
  assign n3311 = n3162 & ~n3309;
  assign n3312 = ~n3310 & ~n3311;
  assign n3313 = ~n3151 & n3312;
  assign n3314 = n3151 & ~n3312;
  assign n3315 = ~n3313 & ~n3314;
  assign n3316 = ~n3150 & n3315;
  assign n3317 = n3150 & ~n3315;
  assign n3318 = ~n3316 & ~n3317;
  assign n3319 = ~n3132 & n3318;
  assign n3320 = n3132 & ~n3318;
  assign po29  = ~n3319 & ~n3320;
  assign n3322 = ~n3316 & ~n3319;
  assign n3323 = ~n3310 & ~n3313;
  assign n3324 = ~n3304 & ~n3307;
  assign n3325 = pi88  & n493;
  assign n3326 = pi86  & n533;
  assign n3327 = pi87  & n488;
  assign n3328 = ~n3326 & ~n3327;
  assign n3329 = ~n3325 & n3328;
  assign n3330 = n496 & n2277;
  assign n3331 = n3329 & ~n3330;
  assign n3332 = pi8  & ~n3331;
  assign n3333 = pi8  & ~n3332;
  assign n3334 = ~n3331 & ~n3332;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = ~n3268 & ~n3272;
  assign n3337 = ~n3233 & ~n3235;
  assign n3338 = pi76  & n1582;
  assign n3339 = pi74  & n1713;
  assign n3340 = pi75  & n1577;
  assign n3341 = ~n3339 & ~n3340;
  assign n3342 = ~n3338 & n3341;
  assign n3343 = n881 & n1585;
  assign n3344 = n3342 & ~n3343;
  assign n3345 = pi20  & ~n3344;
  assign n3346 = pi20  & ~n3345;
  assign n3347 = ~n3344 & ~n3345;
  assign n3348 = ~n3346 & ~n3347;
  assign n3349 = ~n3227 & ~n3229;
  assign n3350 = pi73  & n2004;
  assign n3351 = pi71  & n2141;
  assign n3352 = pi72  & n1999;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = ~n3350 & n3353;
  assign n3355 = n639 & n2007;
  assign n3356 = n3354 & ~n3355;
  assign n3357 = pi23  & ~n3356;
  assign n3358 = pi23  & ~n3357;
  assign n3359 = ~n3356 & ~n3357;
  assign n3360 = ~n3358 & ~n3359;
  assign n3361 = pi67  & n2976;
  assign n3362 = pi65  & n3182;
  assign n3363 = pi66  & n2971;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = ~n3361 & n3364;
  assign n3366 = n313 & n2979;
  assign n3367 = n3365 & ~n3366;
  assign n3368 = pi29  & ~n3367;
  assign n3369 = pi29  & ~n3368;
  assign n3370 = ~n3367 & ~n3368;
  assign n3371 = ~n3369 & ~n3370;
  assign n3372 = pi29  & ~pi30 ;
  assign n3373 = ~pi29  & pi30 ;
  assign n3374 = ~n3372 & ~n3373;
  assign n3375 = pi64  & ~n3374;
  assign n3376 = n3194 & n3375;
  assign n3377 = ~n3194 & ~n3375;
  assign n3378 = ~n3376 & ~n3377;
  assign n3379 = ~n3371 & n3378;
  assign n3380 = n3371 & ~n3378;
  assign n3381 = ~n3379 & ~n3380;
  assign n3382 = pi70  & n2486;
  assign n3383 = pi68  & n2644;
  assign n3384 = pi69  & n2481;
  assign n3385 = ~n3383 & ~n3384;
  assign n3386 = ~n3382 & n3385;
  assign n3387 = n430 & n2489;
  assign n3388 = n3386 & ~n3387;
  assign n3389 = pi26  & ~n3388;
  assign n3390 = pi26  & ~n3389;
  assign n3391 = ~n3388 & ~n3389;
  assign n3392 = ~n3390 & ~n3391;
  assign n3393 = n3381 & ~n3392;
  assign n3394 = ~n3381 & n3392;
  assign n3395 = ~n3393 & ~n3394;
  assign n3396 = ~n3212 & n3395;
  assign n3397 = n3212 & ~n3395;
  assign n3398 = ~n3396 & ~n3397;
  assign n3399 = ~n3360 & n3398;
  assign n3400 = n3360 & ~n3398;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = ~n3349 & n3401;
  assign n3403 = n3349 & ~n3401;
  assign n3404 = ~n3402 & ~n3403;
  assign n3405 = n3348 & ~n3404;
  assign n3406 = ~n3348 & n3404;
  assign n3407 = ~n3405 & ~n3406;
  assign n3408 = ~n3337 & n3407;
  assign n3409 = n3337 & ~n3407;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = pi79  & n1269;
  assign n3412 = pi77  & n1340;
  assign n3413 = pi78  & n1264;
  assign n3414 = ~n3412 & ~n3413;
  assign n3415 = ~n3411 & n3414;
  assign n3416 = n1105 & n1272;
  assign n3417 = n3415 & ~n3416;
  assign n3418 = pi17  & ~n3417;
  assign n3419 = pi17  & ~n3418;
  assign n3420 = ~n3417 & ~n3418;
  assign n3421 = ~n3419 & ~n3420;
  assign n3422 = n3410 & ~n3421;
  assign n3423 = n3410 & ~n3422;
  assign n3424 = ~n3421 & ~n3422;
  assign n3425 = ~n3423 & ~n3424;
  assign n3426 = ~n3249 & ~n3255;
  assign n3427 = n3425 & n3426;
  assign n3428 = ~n3425 & ~n3426;
  assign n3429 = ~n3427 & ~n3428;
  assign n3430 = pi82  & n918;
  assign n3431 = pi80  & n1031;
  assign n3432 = pi81  & n913;
  assign n3433 = ~n3431 & ~n3432;
  assign n3434 = ~n3430 & n3433;
  assign n3435 = n921 & n1532;
  assign n3436 = n3434 & ~n3435;
  assign n3437 = pi14  & ~n3436;
  assign n3438 = pi14  & ~n3437;
  assign n3439 = ~n3436 & ~n3437;
  assign n3440 = ~n3438 & ~n3439;
  assign n3441 = n3429 & ~n3440;
  assign n3442 = ~n3429 & n3440;
  assign n3443 = ~n3441 & ~n3442;
  assign n3444 = n3336 & ~n3443;
  assign n3445 = ~n3336 & n3443;
  assign n3446 = ~n3444 & ~n3445;
  assign n3447 = pi85  & n675;
  assign n3448 = pi83  & n769;
  assign n3449 = pi84  & n670;
  assign n3450 = ~n3448 & ~n3449;
  assign n3451 = ~n3447 & n3450;
  assign n3452 = n678 & n1943;
  assign n3453 = n3451 & ~n3452;
  assign n3454 = pi11  & ~n3453;
  assign n3455 = pi11  & ~n3454;
  assign n3456 = ~n3453 & ~n3454;
  assign n3457 = ~n3455 & ~n3456;
  assign n3458 = n3446 & ~n3457;
  assign n3459 = n3446 & ~n3458;
  assign n3460 = ~n3457 & ~n3458;
  assign n3461 = ~n3459 & ~n3460;
  assign n3462 = ~n3290 & ~n3461;
  assign n3463 = n3290 & n3461;
  assign n3464 = ~n3462 & ~n3463;
  assign n3465 = ~n3335 & n3464;
  assign n3466 = n3335 & ~n3464;
  assign n3467 = ~n3465 & ~n3466;
  assign n3468 = n3324 & ~n3467;
  assign n3469 = ~n3324 & n3467;
  assign n3470 = ~n3468 & ~n3469;
  assign n3471 = pi91  & n340;
  assign n3472 = pi89  & n380;
  assign n3473 = pi90  & n335;
  assign n3474 = ~n3472 & ~n3473;
  assign n3475 = ~n3471 & n3474;
  assign n3476 = n343 & n2926;
  assign n3477 = n3475 & ~n3476;
  assign n3478 = pi5  & ~n3477;
  assign n3479 = pi5  & ~n3478;
  assign n3480 = ~n3477 & ~n3478;
  assign n3481 = ~n3479 & ~n3480;
  assign n3482 = n3470 & ~n3481;
  assign n3483 = ~n3470 & n3481;
  assign n3484 = ~n3482 & ~n3483;
  assign n3485 = n3323 & ~n3484;
  assign n3486 = ~n3323 & n3484;
  assign n3487 = ~n3485 & ~n3486;
  assign n3488 = pi94  & n264;
  assign n3489 = pi92  & n281;
  assign n3490 = pi93  & n259;
  assign n3491 = ~n3489 & ~n3490;
  assign n3492 = ~n3488 & n3491;
  assign n3493 = ~n3140 & ~n3142;
  assign n3494 = ~pi93  & ~pi94 ;
  assign n3495 = pi93  & pi94 ;
  assign n3496 = ~n3494 & ~n3495;
  assign n3497 = ~n3493 & n3496;
  assign n3498 = n3493 & ~n3496;
  assign n3499 = ~n3497 & ~n3498;
  assign n3500 = n267 & n3499;
  assign n3501 = n3492 & ~n3500;
  assign n3502 = pi2  & ~n3501;
  assign n3503 = pi2  & ~n3502;
  assign n3504 = ~n3501 & ~n3502;
  assign n3505 = ~n3503 & ~n3504;
  assign n3506 = n3487 & ~n3505;
  assign n3507 = ~n3487 & n3505;
  assign n3508 = ~n3506 & ~n3507;
  assign n3509 = ~n3322 & n3508;
  assign n3510 = n3322 & ~n3508;
  assign po30  = ~n3509 & ~n3510;
  assign n3512 = ~n3506 & ~n3509;
  assign n3513 = ~n3482 & ~n3486;
  assign n3514 = ~n3465 & ~n3469;
  assign n3515 = ~n3441 & ~n3445;
  assign n3516 = ~n3399 & ~n3402;
  assign n3517 = ~n3393 & ~n3396;
  assign n3518 = pi71  & n2486;
  assign n3519 = pi69  & n2644;
  assign n3520 = pi70  & n2481;
  assign n3521 = ~n3519 & ~n3520;
  assign n3522 = ~n3518 & n3521;
  assign n3523 = n476 & n2489;
  assign n3524 = n3522 & ~n3523;
  assign n3525 = pi26  & ~n3524;
  assign n3526 = pi26  & ~n3525;
  assign n3527 = ~n3524 & ~n3525;
  assign n3528 = ~n3526 & ~n3527;
  assign n3529 = ~n3376 & ~n3379;
  assign n3530 = pi68  & n2976;
  assign n3531 = pi66  & n3182;
  assign n3532 = pi67  & n2971;
  assign n3533 = ~n3531 & ~n3532;
  assign n3534 = ~n3530 & n3533;
  assign n3535 = n364 & n2979;
  assign n3536 = n3534 & ~n3535;
  assign n3537 = pi29  & ~n3536;
  assign n3538 = pi29  & ~n3537;
  assign n3539 = ~n3536 & ~n3537;
  assign n3540 = ~n3538 & ~n3539;
  assign n3541 = pi32  & ~n3375;
  assign n3542 = ~pi30  & pi31 ;
  assign n3543 = pi30  & ~pi31 ;
  assign n3544 = ~n3542 & ~n3543;
  assign n3545 = n3374 & ~n3544;
  assign n3546 = pi64  & n3545;
  assign n3547 = ~pi31  & pi32 ;
  assign n3548 = pi31  & ~pi32 ;
  assign n3549 = ~n3547 & ~n3548;
  assign n3550 = ~n3374 & n3549;
  assign n3551 = pi65  & n3550;
  assign n3552 = ~n3546 & ~n3551;
  assign n3553 = ~n3374 & ~n3549;
  assign n3554 = n270 & n3553;
  assign n3555 = n3552 & ~n3554;
  assign n3556 = pi32  & ~n3555;
  assign n3557 = pi32  & ~n3556;
  assign n3558 = ~n3555 & ~n3556;
  assign n3559 = ~n3557 & ~n3558;
  assign n3560 = n3541 & ~n3559;
  assign n3561 = ~n3541 & n3559;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = ~n3540 & n3562;
  assign n3564 = n3540 & ~n3562;
  assign n3565 = ~n3563 & ~n3564;
  assign n3566 = ~n3529 & n3565;
  assign n3567 = n3529 & ~n3565;
  assign n3568 = ~n3566 & ~n3567;
  assign n3569 = ~n3528 & n3568;
  assign n3570 = n3528 & ~n3568;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = ~n3517 & n3571;
  assign n3573 = n3517 & ~n3571;
  assign n3574 = ~n3572 & ~n3573;
  assign n3575 = pi74  & n2004;
  assign n3576 = pi72  & n2141;
  assign n3577 = pi73  & n1999;
  assign n3578 = ~n3576 & ~n3577;
  assign n3579 = ~n3575 & n3578;
  assign n3580 = n722 & n2007;
  assign n3581 = n3579 & ~n3580;
  assign n3582 = pi23  & ~n3581;
  assign n3583 = pi23  & ~n3582;
  assign n3584 = ~n3581 & ~n3582;
  assign n3585 = ~n3583 & ~n3584;
  assign n3586 = n3574 & ~n3585;
  assign n3587 = ~n3574 & n3585;
  assign n3588 = ~n3586 & ~n3587;
  assign n3589 = n3516 & ~n3588;
  assign n3590 = ~n3516 & n3588;
  assign n3591 = ~n3589 & ~n3590;
  assign n3592 = pi77  & n1582;
  assign n3593 = pi75  & n1713;
  assign n3594 = pi76  & n1577;
  assign n3595 = ~n3593 & ~n3594;
  assign n3596 = ~n3592 & n3595;
  assign n3597 = n984 & n1585;
  assign n3598 = n3596 & ~n3597;
  assign n3599 = pi20  & ~n3598;
  assign n3600 = pi20  & ~n3599;
  assign n3601 = ~n3598 & ~n3599;
  assign n3602 = ~n3600 & ~n3601;
  assign n3603 = ~n3591 & n3602;
  assign n3604 = n3591 & ~n3602;
  assign n3605 = ~n3603 & ~n3604;
  assign n3606 = ~n3406 & ~n3408;
  assign n3607 = n3605 & ~n3606;
  assign n3608 = ~n3605 & n3606;
  assign n3609 = ~n3607 & ~n3608;
  assign n3610 = pi80  & n1269;
  assign n3611 = pi78  & n1340;
  assign n3612 = pi79  & n1264;
  assign n3613 = ~n3611 & ~n3612;
  assign n3614 = ~n3610 & n3613;
  assign n3615 = n1205 & n1272;
  assign n3616 = n3614 & ~n3615;
  assign n3617 = pi17  & ~n3616;
  assign n3618 = pi17  & ~n3617;
  assign n3619 = ~n3616 & ~n3617;
  assign n3620 = ~n3618 & ~n3619;
  assign n3621 = n3609 & ~n3620;
  assign n3622 = n3609 & ~n3621;
  assign n3623 = ~n3620 & ~n3621;
  assign n3624 = ~n3622 & ~n3623;
  assign n3625 = ~n3422 & ~n3428;
  assign n3626 = n3624 & n3625;
  assign n3627 = ~n3624 & ~n3625;
  assign n3628 = ~n3626 & ~n3627;
  assign n3629 = pi83  & n918;
  assign n3630 = pi81  & n1031;
  assign n3631 = pi82  & n913;
  assign n3632 = ~n3630 & ~n3631;
  assign n3633 = ~n3629 & n3632;
  assign n3634 = n921 & n1672;
  assign n3635 = n3633 & ~n3634;
  assign n3636 = pi14  & ~n3635;
  assign n3637 = pi14  & ~n3636;
  assign n3638 = ~n3635 & ~n3636;
  assign n3639 = ~n3637 & ~n3638;
  assign n3640 = n3628 & ~n3639;
  assign n3641 = ~n3628 & n3639;
  assign n3642 = ~n3640 & ~n3641;
  assign n3643 = n3515 & ~n3642;
  assign n3644 = ~n3515 & n3642;
  assign n3645 = ~n3643 & ~n3644;
  assign n3646 = pi86  & n675;
  assign n3647 = pi84  & n769;
  assign n3648 = pi85  & n670;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = ~n3646 & n3649;
  assign n3651 = n678 & n2099;
  assign n3652 = n3650 & ~n3651;
  assign n3653 = pi11  & ~n3652;
  assign n3654 = pi11  & ~n3653;
  assign n3655 = ~n3652 & ~n3653;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = n3645 & ~n3656;
  assign n3658 = n3645 & ~n3657;
  assign n3659 = ~n3656 & ~n3657;
  assign n3660 = ~n3658 & ~n3659;
  assign n3661 = ~n3458 & ~n3462;
  assign n3662 = n3660 & n3661;
  assign n3663 = ~n3660 & ~n3661;
  assign n3664 = ~n3662 & ~n3663;
  assign n3665 = pi89  & n493;
  assign n3666 = pi87  & n533;
  assign n3667 = pi88  & n488;
  assign n3668 = ~n3666 & ~n3667;
  assign n3669 = ~n3665 & n3668;
  assign n3670 = n496 & n2432;
  assign n3671 = n3669 & ~n3670;
  assign n3672 = pi8  & ~n3671;
  assign n3673 = pi8  & ~n3672;
  assign n3674 = ~n3671 & ~n3672;
  assign n3675 = ~n3673 & ~n3674;
  assign n3676 = n3664 & ~n3675;
  assign n3677 = ~n3664 & n3675;
  assign n3678 = ~n3676 & ~n3677;
  assign n3679 = n3514 & ~n3678;
  assign n3680 = ~n3514 & n3678;
  assign n3681 = ~n3679 & ~n3680;
  assign n3682 = pi92  & n340;
  assign n3683 = pi90  & n380;
  assign n3684 = pi91  & n335;
  assign n3685 = ~n3683 & ~n3684;
  assign n3686 = ~n3682 & n3685;
  assign n3687 = n343 & n3119;
  assign n3688 = n3686 & ~n3687;
  assign n3689 = pi5  & ~n3688;
  assign n3690 = pi5  & ~n3689;
  assign n3691 = ~n3688 & ~n3689;
  assign n3692 = ~n3690 & ~n3691;
  assign n3693 = n3681 & ~n3692;
  assign n3694 = ~n3681 & n3692;
  assign n3695 = ~n3693 & ~n3694;
  assign n3696 = n3513 & ~n3695;
  assign n3697 = ~n3513 & n3695;
  assign n3698 = ~n3696 & ~n3697;
  assign n3699 = pi95  & n264;
  assign n3700 = pi93  & n281;
  assign n3701 = pi94  & n259;
  assign n3702 = ~n3700 & ~n3701;
  assign n3703 = ~n3699 & n3702;
  assign n3704 = ~n3495 & ~n3497;
  assign n3705 = ~pi94  & ~pi95 ;
  assign n3706 = pi94  & pi95 ;
  assign n3707 = ~n3705 & ~n3706;
  assign n3708 = ~n3704 & n3707;
  assign n3709 = n3704 & ~n3707;
  assign n3710 = ~n3708 & ~n3709;
  assign n3711 = n267 & n3710;
  assign n3712 = n3703 & ~n3711;
  assign n3713 = pi2  & ~n3712;
  assign n3714 = pi2  & ~n3713;
  assign n3715 = ~n3712 & ~n3713;
  assign n3716 = ~n3714 & ~n3715;
  assign n3717 = n3698 & ~n3716;
  assign n3718 = ~n3698 & n3716;
  assign n3719 = ~n3717 & ~n3718;
  assign n3720 = ~n3512 & n3719;
  assign n3721 = n3512 & ~n3719;
  assign po31  = ~n3720 & ~n3721;
  assign n3723 = ~n3717 & ~n3720;
  assign n3724 = ~n3693 & ~n3697;
  assign n3725 = ~n3676 & ~n3680;
  assign n3726 = ~n3657 & ~n3663;
  assign n3727 = ~n3640 & ~n3644;
  assign n3728 = ~n3621 & ~n3627;
  assign n3729 = ~n3604 & ~n3607;
  assign n3730 = ~n3586 & ~n3590;
  assign n3731 = ~n3569 & ~n3572;
  assign n3732 = ~n3563 & ~n3566;
  assign n3733 = pi66  & n3550;
  assign n3734 = n3374 & ~n3549;
  assign n3735 = n3544 & n3734;
  assign n3736 = pi64  & n3735;
  assign n3737 = pi65  & n3545;
  assign n3738 = ~n3736 & ~n3737;
  assign n3739 = ~n3733 & n3738;
  assign n3740 = n291 & n3553;
  assign n3741 = n3739 & ~n3740;
  assign n3742 = pi32  & ~n3741;
  assign n3743 = pi32  & ~n3742;
  assign n3744 = ~n3741 & ~n3742;
  assign n3745 = ~n3743 & ~n3744;
  assign n3746 = ~n3560 & n3745;
  assign n3747 = n3560 & ~n3745;
  assign n3748 = ~n3746 & ~n3747;
  assign n3749 = pi69  & n2976;
  assign n3750 = pi67  & n3182;
  assign n3751 = pi68  & n2971;
  assign n3752 = ~n3750 & ~n3751;
  assign n3753 = ~n3749 & n3752;
  assign n3754 = n405 & n2979;
  assign n3755 = n3753 & ~n3754;
  assign n3756 = pi29  & ~n3755;
  assign n3757 = pi29  & ~n3756;
  assign n3758 = ~n3755 & ~n3756;
  assign n3759 = ~n3757 & ~n3758;
  assign n3760 = n3748 & ~n3759;
  assign n3761 = ~n3748 & n3759;
  assign n3762 = ~n3732 & ~n3761;
  assign n3763 = ~n3760 & n3762;
  assign n3764 = ~n3732 & ~n3763;
  assign n3765 = ~n3760 & ~n3763;
  assign n3766 = ~n3761 & n3765;
  assign n3767 = ~n3764 & ~n3766;
  assign n3768 = pi72  & n2486;
  assign n3769 = pi70  & n2644;
  assign n3770 = pi71  & n2481;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = ~n3768 & n3771;
  assign n3773 = n575 & n2489;
  assign n3774 = n3772 & ~n3773;
  assign n3775 = pi26  & ~n3774;
  assign n3776 = pi26  & ~n3775;
  assign n3777 = ~n3774 & ~n3775;
  assign n3778 = ~n3776 & ~n3777;
  assign n3779 = ~n3767 & ~n3778;
  assign n3780 = n3767 & n3778;
  assign n3781 = ~n3779 & ~n3780;
  assign n3782 = n3731 & ~n3781;
  assign n3783 = ~n3731 & n3781;
  assign n3784 = ~n3782 & ~n3783;
  assign n3785 = pi75  & n2004;
  assign n3786 = pi73  & n2141;
  assign n3787 = pi74  & n1999;
  assign n3788 = ~n3786 & ~n3787;
  assign n3789 = ~n3785 & n3788;
  assign n3790 = n747 & n2007;
  assign n3791 = n3789 & ~n3790;
  assign n3792 = pi23  & ~n3791;
  assign n3793 = pi23  & ~n3792;
  assign n3794 = ~n3791 & ~n3792;
  assign n3795 = ~n3793 & ~n3794;
  assign n3796 = n3784 & ~n3795;
  assign n3797 = ~n3784 & n3795;
  assign n3798 = ~n3730 & ~n3797;
  assign n3799 = ~n3796 & n3798;
  assign n3800 = ~n3730 & ~n3799;
  assign n3801 = ~n3796 & ~n3799;
  assign n3802 = ~n3797 & n3801;
  assign n3803 = ~n3800 & ~n3802;
  assign n3804 = pi78  & n1582;
  assign n3805 = pi76  & n1713;
  assign n3806 = pi77  & n1577;
  assign n3807 = ~n3805 & ~n3806;
  assign n3808 = ~n3804 & n3807;
  assign n3809 = n1009 & n1585;
  assign n3810 = n3808 & ~n3809;
  assign n3811 = pi20  & ~n3810;
  assign n3812 = pi20  & ~n3811;
  assign n3813 = ~n3810 & ~n3811;
  assign n3814 = ~n3812 & ~n3813;
  assign n3815 = n3803 & n3814;
  assign n3816 = ~n3803 & ~n3814;
  assign n3817 = ~n3815 & ~n3816;
  assign n3818 = ~n3729 & n3817;
  assign n3819 = n3729 & ~n3817;
  assign n3820 = ~n3818 & ~n3819;
  assign n3821 = pi81  & n1269;
  assign n3822 = pi79  & n1340;
  assign n3823 = pi80  & n1264;
  assign n3824 = ~n3822 & ~n3823;
  assign n3825 = ~n3821 & n3824;
  assign n3826 = n1272 & n1413;
  assign n3827 = n3825 & ~n3826;
  assign n3828 = pi17  & ~n3827;
  assign n3829 = pi17  & ~n3828;
  assign n3830 = ~n3827 & ~n3828;
  assign n3831 = ~n3829 & ~n3830;
  assign n3832 = n3820 & ~n3831;
  assign n3833 = ~n3820 & n3831;
  assign n3834 = ~n3832 & ~n3833;
  assign n3835 = n3728 & ~n3834;
  assign n3836 = ~n3728 & n3834;
  assign n3837 = ~n3835 & ~n3836;
  assign n3838 = pi84  & n918;
  assign n3839 = pi82  & n1031;
  assign n3840 = pi83  & n913;
  assign n3841 = ~n3839 & ~n3840;
  assign n3842 = ~n3838 & n3841;
  assign n3843 = n921 & n1805;
  assign n3844 = n3842 & ~n3843;
  assign n3845 = pi14  & ~n3844;
  assign n3846 = pi14  & ~n3845;
  assign n3847 = ~n3844 & ~n3845;
  assign n3848 = ~n3846 & ~n3847;
  assign n3849 = n3837 & ~n3848;
  assign n3850 = ~n3837 & n3848;
  assign n3851 = ~n3727 & ~n3850;
  assign n3852 = ~n3849 & n3851;
  assign n3853 = ~n3727 & ~n3852;
  assign n3854 = ~n3849 & ~n3852;
  assign n3855 = ~n3850 & n3854;
  assign n3856 = ~n3853 & ~n3855;
  assign n3857 = pi87  & n675;
  assign n3858 = pi85  & n769;
  assign n3859 = pi86  & n670;
  assign n3860 = ~n3858 & ~n3859;
  assign n3861 = ~n3857 & n3860;
  assign n3862 = n678 & n2252;
  assign n3863 = n3861 & ~n3862;
  assign n3864 = pi11  & ~n3863;
  assign n3865 = pi11  & ~n3864;
  assign n3866 = ~n3863 & ~n3864;
  assign n3867 = ~n3865 & ~n3866;
  assign n3868 = n3856 & n3867;
  assign n3869 = ~n3856 & ~n3867;
  assign n3870 = ~n3868 & ~n3869;
  assign n3871 = ~n3726 & n3870;
  assign n3872 = n3726 & ~n3870;
  assign n3873 = ~n3871 & ~n3872;
  assign n3874 = pi90  & n493;
  assign n3875 = pi88  & n533;
  assign n3876 = pi89  & n488;
  assign n3877 = ~n3875 & ~n3876;
  assign n3878 = ~n3874 & n3877;
  assign n3879 = n496 & n2606;
  assign n3880 = n3878 & ~n3879;
  assign n3881 = pi8  & ~n3880;
  assign n3882 = pi8  & ~n3881;
  assign n3883 = ~n3880 & ~n3881;
  assign n3884 = ~n3882 & ~n3883;
  assign n3885 = n3873 & ~n3884;
  assign n3886 = ~n3873 & n3884;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = n3725 & ~n3887;
  assign n3889 = ~n3725 & n3887;
  assign n3890 = ~n3888 & ~n3889;
  assign n3891 = pi93  & n340;
  assign n3892 = pi91  & n380;
  assign n3893 = pi92  & n335;
  assign n3894 = ~n3892 & ~n3893;
  assign n3895 = ~n3891 & n3894;
  assign n3896 = n343 & n3144;
  assign n3897 = n3895 & ~n3896;
  assign n3898 = pi5  & ~n3897;
  assign n3899 = pi5  & ~n3898;
  assign n3900 = ~n3897 & ~n3898;
  assign n3901 = ~n3899 & ~n3900;
  assign n3902 = n3890 & ~n3901;
  assign n3903 = ~n3890 & n3901;
  assign n3904 = ~n3724 & ~n3903;
  assign n3905 = ~n3902 & n3904;
  assign n3906 = ~n3724 & ~n3905;
  assign n3907 = ~n3902 & ~n3905;
  assign n3908 = ~n3903 & n3907;
  assign n3909 = ~n3906 & ~n3908;
  assign n3910 = pi96  & n264;
  assign n3911 = pi94  & n281;
  assign n3912 = pi95  & n259;
  assign n3913 = ~n3911 & ~n3912;
  assign n3914 = ~n3910 & n3913;
  assign n3915 = ~n3706 & ~n3708;
  assign n3916 = ~pi95  & ~pi96 ;
  assign n3917 = pi95  & pi96 ;
  assign n3918 = ~n3916 & ~n3917;
  assign n3919 = ~n3915 & n3918;
  assign n3920 = n3915 & ~n3918;
  assign n3921 = ~n3919 & ~n3920;
  assign n3922 = n267 & n3921;
  assign n3923 = n3914 & ~n3922;
  assign n3924 = pi2  & ~n3923;
  assign n3925 = pi2  & ~n3924;
  assign n3926 = ~n3923 & ~n3924;
  assign n3927 = ~n3925 & ~n3926;
  assign n3928 = ~n3909 & ~n3927;
  assign n3929 = n3909 & n3927;
  assign n3930 = ~n3928 & ~n3929;
  assign n3931 = ~n3723 & n3930;
  assign n3932 = n3723 & ~n3930;
  assign po32  = ~n3931 & ~n3932;
  assign n3934 = ~n3928 & ~n3931;
  assign n3935 = pi97  & n264;
  assign n3936 = pi95  & n281;
  assign n3937 = pi96  & n259;
  assign n3938 = ~n3936 & ~n3937;
  assign n3939 = ~n3935 & n3938;
  assign n3940 = ~n3917 & ~n3919;
  assign n3941 = ~pi96  & ~pi97 ;
  assign n3942 = pi96  & pi97 ;
  assign n3943 = ~n3941 & ~n3942;
  assign n3944 = ~n3940 & n3943;
  assign n3945 = n3940 & ~n3943;
  assign n3946 = ~n3944 & ~n3945;
  assign n3947 = n267 & n3946;
  assign n3948 = n3939 & ~n3947;
  assign n3949 = pi2  & ~n3948;
  assign n3950 = pi2  & ~n3949;
  assign n3951 = ~n3948 & ~n3949;
  assign n3952 = ~n3950 & ~n3951;
  assign n3953 = ~n3885 & ~n3889;
  assign n3954 = ~n3869 & ~n3871;
  assign n3955 = pi88  & n675;
  assign n3956 = pi86  & n769;
  assign n3957 = pi87  & n670;
  assign n3958 = ~n3956 & ~n3957;
  assign n3959 = ~n3955 & n3958;
  assign n3960 = n678 & n2277;
  assign n3961 = n3959 & ~n3960;
  assign n3962 = pi11  & ~n3961;
  assign n3963 = pi11  & ~n3962;
  assign n3964 = ~n3961 & ~n3962;
  assign n3965 = ~n3963 & ~n3964;
  assign n3966 = ~n3832 & ~n3836;
  assign n3967 = pi82  & n1269;
  assign n3968 = pi80  & n1340;
  assign n3969 = pi81  & n1264;
  assign n3970 = ~n3968 & ~n3969;
  assign n3971 = ~n3967 & n3970;
  assign n3972 = n1272 & n1532;
  assign n3973 = n3971 & ~n3972;
  assign n3974 = pi17  & ~n3973;
  assign n3975 = pi17  & ~n3974;
  assign n3976 = ~n3973 & ~n3974;
  assign n3977 = ~n3975 & ~n3976;
  assign n3978 = ~n3816 & ~n3818;
  assign n3979 = ~n3779 & ~n3783;
  assign n3980 = pi73  & n2486;
  assign n3981 = pi71  & n2644;
  assign n3982 = pi72  & n2481;
  assign n3983 = ~n3981 & ~n3982;
  assign n3984 = ~n3980 & n3983;
  assign n3985 = n639 & n2489;
  assign n3986 = n3984 & ~n3985;
  assign n3987 = pi26  & ~n3986;
  assign n3988 = pi26  & ~n3987;
  assign n3989 = ~n3986 & ~n3987;
  assign n3990 = ~n3988 & ~n3989;
  assign n3991 = pi67  & n3550;
  assign n3992 = pi65  & n3735;
  assign n3993 = pi66  & n3545;
  assign n3994 = ~n3992 & ~n3993;
  assign n3995 = ~n3991 & n3994;
  assign n3996 = n313 & n3553;
  assign n3997 = n3995 & ~n3996;
  assign n3998 = pi32  & ~n3997;
  assign n3999 = pi32  & ~n3998;
  assign n4000 = ~n3997 & ~n3998;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = pi32  & ~pi33 ;
  assign n4003 = ~pi32  & pi33 ;
  assign n4004 = ~n4002 & ~n4003;
  assign n4005 = pi64  & ~n4004;
  assign n4006 = n3747 & n4005;
  assign n4007 = ~n3747 & ~n4005;
  assign n4008 = ~n4006 & ~n4007;
  assign n4009 = ~n4001 & n4008;
  assign n4010 = n4001 & ~n4008;
  assign n4011 = ~n4009 & ~n4010;
  assign n4012 = pi70  & n2976;
  assign n4013 = pi68  & n3182;
  assign n4014 = pi69  & n2971;
  assign n4015 = ~n4013 & ~n4014;
  assign n4016 = ~n4012 & n4015;
  assign n4017 = n430 & n2979;
  assign n4018 = n4016 & ~n4017;
  assign n4019 = pi29  & ~n4018;
  assign n4020 = pi29  & ~n4019;
  assign n4021 = ~n4018 & ~n4019;
  assign n4022 = ~n4020 & ~n4021;
  assign n4023 = n4011 & ~n4022;
  assign n4024 = ~n4011 & n4022;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = ~n3765 & n4025;
  assign n4027 = n3765 & ~n4025;
  assign n4028 = ~n4026 & ~n4027;
  assign n4029 = ~n3990 & n4028;
  assign n4030 = n3990 & ~n4028;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = n3979 & ~n4031;
  assign n4033 = ~n3979 & n4031;
  assign n4034 = ~n4032 & ~n4033;
  assign n4035 = pi76  & n2004;
  assign n4036 = pi74  & n2141;
  assign n4037 = pi75  & n1999;
  assign n4038 = ~n4036 & ~n4037;
  assign n4039 = ~n4035 & n4038;
  assign n4040 = n881 & n2007;
  assign n4041 = n4039 & ~n4040;
  assign n4042 = pi23  & ~n4041;
  assign n4043 = pi23  & ~n4042;
  assign n4044 = ~n4041 & ~n4042;
  assign n4045 = ~n4043 & ~n4044;
  assign n4046 = ~n4034 & n4045;
  assign n4047 = n4034 & ~n4045;
  assign n4048 = ~n4046 & ~n4047;
  assign n4049 = ~n3801 & n4048;
  assign n4050 = n3801 & ~n4048;
  assign n4051 = ~n4049 & ~n4050;
  assign n4052 = pi79  & n1582;
  assign n4053 = pi77  & n1713;
  assign n4054 = pi78  & n1577;
  assign n4055 = ~n4053 & ~n4054;
  assign n4056 = ~n4052 & n4055;
  assign n4057 = n1105 & n1585;
  assign n4058 = n4056 & ~n4057;
  assign n4059 = pi20  & ~n4058;
  assign n4060 = pi20  & ~n4059;
  assign n4061 = ~n4058 & ~n4059;
  assign n4062 = ~n4060 & ~n4061;
  assign n4063 = n4051 & ~n4062;
  assign n4064 = n4051 & ~n4063;
  assign n4065 = ~n4062 & ~n4063;
  assign n4066 = ~n4064 & ~n4065;
  assign n4067 = ~n3978 & ~n4066;
  assign n4068 = n3978 & n4066;
  assign n4069 = ~n4067 & ~n4068;
  assign n4070 = ~n3977 & n4069;
  assign n4071 = n3977 & ~n4069;
  assign n4072 = ~n4070 & ~n4071;
  assign n4073 = n3966 & ~n4072;
  assign n4074 = ~n3966 & n4072;
  assign n4075 = ~n4073 & ~n4074;
  assign n4076 = pi85  & n918;
  assign n4077 = pi83  & n1031;
  assign n4078 = pi84  & n913;
  assign n4079 = ~n4077 & ~n4078;
  assign n4080 = ~n4076 & n4079;
  assign n4081 = n921 & n1943;
  assign n4082 = n4080 & ~n4081;
  assign n4083 = pi14  & ~n4082;
  assign n4084 = pi14  & ~n4083;
  assign n4085 = ~n4082 & ~n4083;
  assign n4086 = ~n4084 & ~n4085;
  assign n4087 = n4075 & ~n4086;
  assign n4088 = n4075 & ~n4087;
  assign n4089 = ~n4086 & ~n4087;
  assign n4090 = ~n4088 & ~n4089;
  assign n4091 = ~n3854 & ~n4090;
  assign n4092 = n3854 & n4090;
  assign n4093 = ~n4091 & ~n4092;
  assign n4094 = n3965 & ~n4093;
  assign n4095 = ~n3965 & n4093;
  assign n4096 = ~n4094 & ~n4095;
  assign n4097 = ~n3954 & n4096;
  assign n4098 = n3954 & ~n4096;
  assign n4099 = ~n4097 & ~n4098;
  assign n4100 = pi91  & n493;
  assign n4101 = pi89  & n533;
  assign n4102 = pi90  & n488;
  assign n4103 = ~n4101 & ~n4102;
  assign n4104 = ~n4100 & n4103;
  assign n4105 = n496 & n2926;
  assign n4106 = n4104 & ~n4105;
  assign n4107 = pi8  & ~n4106;
  assign n4108 = pi8  & ~n4107;
  assign n4109 = ~n4106 & ~n4107;
  assign n4110 = ~n4108 & ~n4109;
  assign n4111 = n4099 & ~n4110;
  assign n4112 = ~n4099 & n4110;
  assign n4113 = ~n4111 & ~n4112;
  assign n4114 = n3953 & ~n4113;
  assign n4115 = ~n3953 & n4113;
  assign n4116 = ~n4114 & ~n4115;
  assign n4117 = pi94  & n340;
  assign n4118 = pi92  & n380;
  assign n4119 = pi93  & n335;
  assign n4120 = ~n4118 & ~n4119;
  assign n4121 = ~n4117 & n4120;
  assign n4122 = n343 & n3499;
  assign n4123 = n4121 & ~n4122;
  assign n4124 = pi5  & ~n4123;
  assign n4125 = pi5  & ~n4124;
  assign n4126 = ~n4123 & ~n4124;
  assign n4127 = ~n4125 & ~n4126;
  assign n4128 = n4116 & ~n4127;
  assign n4129 = ~n4116 & n4127;
  assign n4130 = ~n4128 & ~n4129;
  assign n4131 = ~n3907 & n4130;
  assign n4132 = n3907 & ~n4130;
  assign n4133 = ~n4131 & ~n4132;
  assign n4134 = ~n3952 & n4133;
  assign n4135 = n3952 & ~n4133;
  assign n4136 = ~n4134 & ~n4135;
  assign n4137 = ~n3934 & n4136;
  assign n4138 = n3934 & ~n4136;
  assign po33  = ~n4137 & ~n4138;
  assign n4140 = ~n4134 & ~n4137;
  assign n4141 = ~n4128 & ~n4131;
  assign n4142 = ~n4111 & ~n4115;
  assign n4143 = ~n4095 & ~n4097;
  assign n4144 = ~n4087 & ~n4091;
  assign n4145 = ~n4070 & ~n4074;
  assign n4146 = ~n4063 & ~n4067;
  assign n4147 = ~n4047 & ~n4049;
  assign n4148 = ~n4029 & ~n4033;
  assign n4149 = ~n4023 & ~n4026;
  assign n4150 = pi71  & n2976;
  assign n4151 = pi69  & n3182;
  assign n4152 = pi70  & n2971;
  assign n4153 = ~n4151 & ~n4152;
  assign n4154 = ~n4150 & n4153;
  assign n4155 = n476 & n2979;
  assign n4156 = n4154 & ~n4155;
  assign n4157 = pi29  & ~n4156;
  assign n4158 = pi29  & ~n4157;
  assign n4159 = ~n4156 & ~n4157;
  assign n4160 = ~n4158 & ~n4159;
  assign n4161 = ~n4006 & ~n4009;
  assign n4162 = pi68  & n3550;
  assign n4163 = pi66  & n3735;
  assign n4164 = pi67  & n3545;
  assign n4165 = ~n4163 & ~n4164;
  assign n4166 = ~n4162 & n4165;
  assign n4167 = n364 & n3553;
  assign n4168 = n4166 & ~n4167;
  assign n4169 = pi32  & ~n4168;
  assign n4170 = pi32  & ~n4169;
  assign n4171 = ~n4168 & ~n4169;
  assign n4172 = ~n4170 & ~n4171;
  assign n4173 = pi35  & ~n4005;
  assign n4174 = ~pi33  & pi34 ;
  assign n4175 = pi33  & ~pi34 ;
  assign n4176 = ~n4174 & ~n4175;
  assign n4177 = n4004 & ~n4176;
  assign n4178 = pi64  & n4177;
  assign n4179 = ~pi34  & pi35 ;
  assign n4180 = pi34  & ~pi35 ;
  assign n4181 = ~n4179 & ~n4180;
  assign n4182 = ~n4004 & n4181;
  assign n4183 = pi65  & n4182;
  assign n4184 = ~n4178 & ~n4183;
  assign n4185 = ~n4004 & ~n4181;
  assign n4186 = n270 & n4185;
  assign n4187 = n4184 & ~n4186;
  assign n4188 = pi35  & ~n4187;
  assign n4189 = pi35  & ~n4188;
  assign n4190 = ~n4187 & ~n4188;
  assign n4191 = ~n4189 & ~n4190;
  assign n4192 = n4173 & ~n4191;
  assign n4193 = ~n4173 & n4191;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = n4172 & ~n4194;
  assign n4196 = ~n4172 & n4194;
  assign n4197 = ~n4195 & ~n4196;
  assign n4198 = ~n4161 & n4197;
  assign n4199 = n4161 & ~n4197;
  assign n4200 = ~n4198 & ~n4199;
  assign n4201 = n4160 & ~n4200;
  assign n4202 = ~n4160 & n4200;
  assign n4203 = ~n4201 & ~n4202;
  assign n4204 = ~n4149 & n4203;
  assign n4205 = n4149 & ~n4203;
  assign n4206 = ~n4204 & ~n4205;
  assign n4207 = pi74  & n2486;
  assign n4208 = pi72  & n2644;
  assign n4209 = pi73  & n2481;
  assign n4210 = ~n4208 & ~n4209;
  assign n4211 = ~n4207 & n4210;
  assign n4212 = n722 & n2489;
  assign n4213 = n4211 & ~n4212;
  assign n4214 = pi26  & ~n4213;
  assign n4215 = pi26  & ~n4214;
  assign n4216 = ~n4213 & ~n4214;
  assign n4217 = ~n4215 & ~n4216;
  assign n4218 = n4206 & ~n4217;
  assign n4219 = ~n4206 & n4217;
  assign n4220 = ~n4218 & ~n4219;
  assign n4221 = n4148 & ~n4220;
  assign n4222 = ~n4148 & n4220;
  assign n4223 = ~n4221 & ~n4222;
  assign n4224 = pi77  & n2004;
  assign n4225 = pi75  & n2141;
  assign n4226 = pi76  & n1999;
  assign n4227 = ~n4225 & ~n4226;
  assign n4228 = ~n4224 & n4227;
  assign n4229 = n984 & n2007;
  assign n4230 = n4228 & ~n4229;
  assign n4231 = pi23  & ~n4230;
  assign n4232 = pi23  & ~n4231;
  assign n4233 = ~n4230 & ~n4231;
  assign n4234 = ~n4232 & ~n4233;
  assign n4235 = n4223 & ~n4234;
  assign n4236 = ~n4223 & n4234;
  assign n4237 = ~n4147 & ~n4236;
  assign n4238 = ~n4235 & n4237;
  assign n4239 = ~n4147 & ~n4238;
  assign n4240 = ~n4235 & ~n4238;
  assign n4241 = ~n4236 & n4240;
  assign n4242 = ~n4239 & ~n4241;
  assign n4243 = pi80  & n1582;
  assign n4244 = pi78  & n1713;
  assign n4245 = pi79  & n1577;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = ~n4243 & n4246;
  assign n4248 = n1205 & n1585;
  assign n4249 = n4247 & ~n4248;
  assign n4250 = pi20  & ~n4249;
  assign n4251 = pi20  & ~n4250;
  assign n4252 = ~n4249 & ~n4250;
  assign n4253 = ~n4251 & ~n4252;
  assign n4254 = ~n4242 & ~n4253;
  assign n4255 = n4242 & n4253;
  assign n4256 = ~n4254 & ~n4255;
  assign n4257 = n4146 & ~n4256;
  assign n4258 = ~n4146 & n4256;
  assign n4259 = ~n4257 & ~n4258;
  assign n4260 = pi83  & n1269;
  assign n4261 = pi81  & n1340;
  assign n4262 = pi82  & n1264;
  assign n4263 = ~n4261 & ~n4262;
  assign n4264 = ~n4260 & n4263;
  assign n4265 = n1272 & n1672;
  assign n4266 = n4264 & ~n4265;
  assign n4267 = pi17  & ~n4266;
  assign n4268 = pi17  & ~n4267;
  assign n4269 = ~n4266 & ~n4267;
  assign n4270 = ~n4268 & ~n4269;
  assign n4271 = n4259 & ~n4270;
  assign n4272 = ~n4259 & n4270;
  assign n4273 = ~n4271 & ~n4272;
  assign n4274 = n4145 & ~n4273;
  assign n4275 = ~n4145 & n4273;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = pi86  & n918;
  assign n4278 = pi84  & n1031;
  assign n4279 = pi85  & n913;
  assign n4280 = ~n4278 & ~n4279;
  assign n4281 = ~n4277 & n4280;
  assign n4282 = n921 & n2099;
  assign n4283 = n4281 & ~n4282;
  assign n4284 = pi14  & ~n4283;
  assign n4285 = pi14  & ~n4284;
  assign n4286 = ~n4283 & ~n4284;
  assign n4287 = ~n4285 & ~n4286;
  assign n4288 = n4276 & ~n4287;
  assign n4289 = ~n4276 & n4287;
  assign n4290 = ~n4288 & ~n4289;
  assign n4291 = n4144 & ~n4290;
  assign n4292 = ~n4144 & n4290;
  assign n4293 = ~n4291 & ~n4292;
  assign n4294 = pi89  & n675;
  assign n4295 = pi87  & n769;
  assign n4296 = pi88  & n670;
  assign n4297 = ~n4295 & ~n4296;
  assign n4298 = ~n4294 & n4297;
  assign n4299 = n678 & n2432;
  assign n4300 = n4298 & ~n4299;
  assign n4301 = pi11  & ~n4300;
  assign n4302 = pi11  & ~n4301;
  assign n4303 = ~n4300 & ~n4301;
  assign n4304 = ~n4302 & ~n4303;
  assign n4305 = n4293 & ~n4304;
  assign n4306 = ~n4293 & n4304;
  assign n4307 = ~n4143 & ~n4306;
  assign n4308 = ~n4305 & n4307;
  assign n4309 = ~n4143 & ~n4308;
  assign n4310 = ~n4305 & ~n4308;
  assign n4311 = ~n4306 & n4310;
  assign n4312 = ~n4309 & ~n4311;
  assign n4313 = pi92  & n493;
  assign n4314 = pi90  & n533;
  assign n4315 = pi91  & n488;
  assign n4316 = ~n4314 & ~n4315;
  assign n4317 = ~n4313 & n4316;
  assign n4318 = n496 & n3119;
  assign n4319 = n4317 & ~n4318;
  assign n4320 = pi8  & ~n4319;
  assign n4321 = pi8  & ~n4320;
  assign n4322 = ~n4319 & ~n4320;
  assign n4323 = ~n4321 & ~n4322;
  assign n4324 = ~n4312 & ~n4323;
  assign n4325 = n4312 & n4323;
  assign n4326 = ~n4324 & ~n4325;
  assign n4327 = n4142 & ~n4326;
  assign n4328 = ~n4142 & n4326;
  assign n4329 = ~n4327 & ~n4328;
  assign n4330 = pi95  & n340;
  assign n4331 = pi93  & n380;
  assign n4332 = pi94  & n335;
  assign n4333 = ~n4331 & ~n4332;
  assign n4334 = ~n4330 & n4333;
  assign n4335 = n343 & n3710;
  assign n4336 = n4334 & ~n4335;
  assign n4337 = pi5  & ~n4336;
  assign n4338 = pi5  & ~n4337;
  assign n4339 = ~n4336 & ~n4337;
  assign n4340 = ~n4338 & ~n4339;
  assign n4341 = n4329 & ~n4340;
  assign n4342 = ~n4329 & n4340;
  assign n4343 = ~n4141 & ~n4342;
  assign n4344 = ~n4341 & n4343;
  assign n4345 = ~n4141 & ~n4344;
  assign n4346 = ~n4341 & ~n4344;
  assign n4347 = ~n4342 & n4346;
  assign n4348 = ~n4345 & ~n4347;
  assign n4349 = pi98  & n264;
  assign n4350 = pi96  & n281;
  assign n4351 = pi97  & n259;
  assign n4352 = ~n4350 & ~n4351;
  assign n4353 = ~n4349 & n4352;
  assign n4354 = ~n3942 & ~n3944;
  assign n4355 = ~pi97  & ~pi98 ;
  assign n4356 = pi97  & pi98 ;
  assign n4357 = ~n4355 & ~n4356;
  assign n4358 = ~n4354 & n4357;
  assign n4359 = n4354 & ~n4357;
  assign n4360 = ~n4358 & ~n4359;
  assign n4361 = n267 & n4360;
  assign n4362 = n4353 & ~n4361;
  assign n4363 = pi2  & ~n4362;
  assign n4364 = pi2  & ~n4363;
  assign n4365 = ~n4362 & ~n4363;
  assign n4366 = ~n4364 & ~n4365;
  assign n4367 = ~n4348 & ~n4366;
  assign n4368 = n4348 & n4366;
  assign n4369 = ~n4367 & ~n4368;
  assign n4370 = ~n4140 & n4369;
  assign n4371 = n4140 & ~n4369;
  assign po34  = ~n4370 & ~n4371;
  assign n4373 = ~n4367 & ~n4370;
  assign n4374 = ~n4324 & ~n4328;
  assign n4375 = pi90  & n675;
  assign n4376 = pi88  & n769;
  assign n4377 = pi89  & n670;
  assign n4378 = ~n4376 & ~n4377;
  assign n4379 = ~n4375 & n4378;
  assign n4380 = n678 & n2606;
  assign n4381 = n4379 & ~n4380;
  assign n4382 = pi11  & ~n4381;
  assign n4383 = pi11  & ~n4382;
  assign n4384 = ~n4381 & ~n4382;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = ~n4288 & ~n4292;
  assign n4387 = ~n4271 & ~n4275;
  assign n4388 = ~n4254 & ~n4258;
  assign n4389 = pi78  & n2004;
  assign n4390 = pi76  & n2141;
  assign n4391 = pi77  & n1999;
  assign n4392 = ~n4390 & ~n4391;
  assign n4393 = ~n4389 & n4392;
  assign n4394 = n1009 & n2007;
  assign n4395 = n4393 & ~n4394;
  assign n4396 = pi23  & ~n4395;
  assign n4397 = pi23  & ~n4396;
  assign n4398 = ~n4395 & ~n4396;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n4218 & ~n4222;
  assign n4401 = pi75  & n2486;
  assign n4402 = pi73  & n2644;
  assign n4403 = pi74  & n2481;
  assign n4404 = ~n4402 & ~n4403;
  assign n4405 = ~n4401 & n4404;
  assign n4406 = n747 & n2489;
  assign n4407 = n4405 & ~n4406;
  assign n4408 = pi26  & ~n4407;
  assign n4409 = pi26  & ~n4408;
  assign n4410 = ~n4407 & ~n4408;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = ~n4202 & ~n4204;
  assign n4413 = ~n4196 & ~n4198;
  assign n4414 = pi66  & n4182;
  assign n4415 = n4004 & ~n4181;
  assign n4416 = n4176 & n4415;
  assign n4417 = pi64  & n4416;
  assign n4418 = pi65  & n4177;
  assign n4419 = ~n4417 & ~n4418;
  assign n4420 = ~n4414 & n4419;
  assign n4421 = n291 & n4185;
  assign n4422 = n4420 & ~n4421;
  assign n4423 = pi35  & ~n4422;
  assign n4424 = pi35  & ~n4423;
  assign n4425 = ~n4422 & ~n4423;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = ~n4192 & n4426;
  assign n4428 = n4192 & ~n4426;
  assign n4429 = ~n4427 & ~n4428;
  assign n4430 = pi69  & n3550;
  assign n4431 = pi67  & n3735;
  assign n4432 = pi68  & n3545;
  assign n4433 = ~n4431 & ~n4432;
  assign n4434 = ~n4430 & n4433;
  assign n4435 = n405 & n3553;
  assign n4436 = n4434 & ~n4435;
  assign n4437 = pi32  & ~n4436;
  assign n4438 = pi32  & ~n4437;
  assign n4439 = ~n4436 & ~n4437;
  assign n4440 = ~n4438 & ~n4439;
  assign n4441 = n4429 & ~n4440;
  assign n4442 = ~n4429 & n4440;
  assign n4443 = ~n4413 & ~n4442;
  assign n4444 = ~n4441 & n4443;
  assign n4445 = ~n4413 & ~n4444;
  assign n4446 = ~n4441 & ~n4444;
  assign n4447 = ~n4442 & n4446;
  assign n4448 = ~n4445 & ~n4447;
  assign n4449 = pi72  & n2976;
  assign n4450 = pi70  & n3182;
  assign n4451 = pi71  & n2971;
  assign n4452 = ~n4450 & ~n4451;
  assign n4453 = ~n4449 & n4452;
  assign n4454 = n575 & n2979;
  assign n4455 = n4453 & ~n4454;
  assign n4456 = pi29  & ~n4455;
  assign n4457 = pi29  & ~n4456;
  assign n4458 = ~n4455 & ~n4456;
  assign n4459 = ~n4457 & ~n4458;
  assign n4460 = ~n4448 & ~n4459;
  assign n4461 = n4448 & n4459;
  assign n4462 = ~n4460 & ~n4461;
  assign n4463 = ~n4412 & n4462;
  assign n4464 = n4412 & ~n4462;
  assign n4465 = ~n4463 & ~n4464;
  assign n4466 = ~n4411 & n4465;
  assign n4467 = n4411 & ~n4465;
  assign n4468 = ~n4466 & ~n4467;
  assign n4469 = ~n4400 & n4468;
  assign n4470 = n4400 & ~n4468;
  assign n4471 = ~n4469 & ~n4470;
  assign n4472 = n4399 & ~n4471;
  assign n4473 = ~n4399 & n4471;
  assign n4474 = ~n4472 & ~n4473;
  assign n4475 = ~n4240 & n4474;
  assign n4476 = n4240 & ~n4474;
  assign n4477 = ~n4475 & ~n4476;
  assign n4478 = pi81  & n1582;
  assign n4479 = pi79  & n1713;
  assign n4480 = pi80  & n1577;
  assign n4481 = ~n4479 & ~n4480;
  assign n4482 = ~n4478 & n4481;
  assign n4483 = n1413 & n1585;
  assign n4484 = n4482 & ~n4483;
  assign n4485 = pi20  & ~n4484;
  assign n4486 = pi20  & ~n4485;
  assign n4487 = ~n4484 & ~n4485;
  assign n4488 = ~n4486 & ~n4487;
  assign n4489 = n4477 & ~n4488;
  assign n4490 = ~n4477 & n4488;
  assign n4491 = ~n4489 & ~n4490;
  assign n4492 = n4388 & ~n4491;
  assign n4493 = ~n4388 & n4491;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495 = pi84  & n1269;
  assign n4496 = pi82  & n1340;
  assign n4497 = pi83  & n1264;
  assign n4498 = ~n4496 & ~n4497;
  assign n4499 = ~n4495 & n4498;
  assign n4500 = n1272 & n1805;
  assign n4501 = n4499 & ~n4500;
  assign n4502 = pi17  & ~n4501;
  assign n4503 = pi17  & ~n4502;
  assign n4504 = ~n4501 & ~n4502;
  assign n4505 = ~n4503 & ~n4504;
  assign n4506 = n4494 & ~n4505;
  assign n4507 = ~n4494 & n4505;
  assign n4508 = ~n4387 & ~n4507;
  assign n4509 = ~n4506 & n4508;
  assign n4510 = ~n4387 & ~n4509;
  assign n4511 = ~n4506 & ~n4509;
  assign n4512 = ~n4507 & n4511;
  assign n4513 = ~n4510 & ~n4512;
  assign n4514 = pi87  & n918;
  assign n4515 = pi85  & n1031;
  assign n4516 = pi86  & n913;
  assign n4517 = ~n4515 & ~n4516;
  assign n4518 = ~n4514 & n4517;
  assign n4519 = n921 & n2252;
  assign n4520 = n4518 & ~n4519;
  assign n4521 = pi14  & ~n4520;
  assign n4522 = pi14  & ~n4521;
  assign n4523 = ~n4520 & ~n4521;
  assign n4524 = ~n4522 & ~n4523;
  assign n4525 = n4513 & n4524;
  assign n4526 = ~n4513 & ~n4524;
  assign n4527 = ~n4525 & ~n4526;
  assign n4528 = ~n4386 & n4527;
  assign n4529 = n4386 & ~n4527;
  assign n4530 = ~n4528 & ~n4529;
  assign n4531 = n4385 & ~n4530;
  assign n4532 = ~n4385 & n4530;
  assign n4533 = ~n4531 & ~n4532;
  assign n4534 = ~n4310 & n4533;
  assign n4535 = n4310 & ~n4533;
  assign n4536 = ~n4534 & ~n4535;
  assign n4537 = pi93  & n493;
  assign n4538 = pi91  & n533;
  assign n4539 = pi92  & n488;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = ~n4537 & n4540;
  assign n4542 = n496 & n3144;
  assign n4543 = n4541 & ~n4542;
  assign n4544 = pi8  & ~n4543;
  assign n4545 = pi8  & ~n4544;
  assign n4546 = ~n4543 & ~n4544;
  assign n4547 = ~n4545 & ~n4546;
  assign n4548 = n4536 & ~n4547;
  assign n4549 = ~n4536 & n4547;
  assign n4550 = ~n4548 & ~n4549;
  assign n4551 = n4374 & ~n4550;
  assign n4552 = ~n4374 & n4550;
  assign n4553 = ~n4551 & ~n4552;
  assign n4554 = pi96  & n340;
  assign n4555 = pi94  & n380;
  assign n4556 = pi95  & n335;
  assign n4557 = ~n4555 & ~n4556;
  assign n4558 = ~n4554 & n4557;
  assign n4559 = n343 & n3921;
  assign n4560 = n4558 & ~n4559;
  assign n4561 = pi5  & ~n4560;
  assign n4562 = pi5  & ~n4561;
  assign n4563 = ~n4560 & ~n4561;
  assign n4564 = ~n4562 & ~n4563;
  assign n4565 = n4553 & ~n4564;
  assign n4566 = ~n4553 & n4564;
  assign n4567 = ~n4346 & ~n4566;
  assign n4568 = ~n4565 & n4567;
  assign n4569 = ~n4346 & ~n4568;
  assign n4570 = ~n4565 & ~n4568;
  assign n4571 = ~n4566 & n4570;
  assign n4572 = ~n4569 & ~n4571;
  assign n4573 = pi99  & n264;
  assign n4574 = pi97  & n281;
  assign n4575 = pi98  & n259;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = ~n4573 & n4576;
  assign n4578 = ~n4356 & ~n4358;
  assign n4579 = ~pi98  & ~pi99 ;
  assign n4580 = pi98  & pi99 ;
  assign n4581 = ~n4579 & ~n4580;
  assign n4582 = ~n4578 & n4581;
  assign n4583 = n4578 & ~n4581;
  assign n4584 = ~n4582 & ~n4583;
  assign n4585 = n267 & n4584;
  assign n4586 = n4577 & ~n4585;
  assign n4587 = pi2  & ~n4586;
  assign n4588 = pi2  & ~n4587;
  assign n4589 = ~n4586 & ~n4587;
  assign n4590 = ~n4588 & ~n4589;
  assign n4591 = ~n4572 & ~n4590;
  assign n4592 = n4572 & n4590;
  assign n4593 = ~n4591 & ~n4592;
  assign n4594 = ~n4373 & n4593;
  assign n4595 = n4373 & ~n4593;
  assign po35  = ~n4594 & ~n4595;
  assign n4597 = ~n4591 & ~n4594;
  assign n4598 = pi97  & n340;
  assign n4599 = pi95  & n380;
  assign n4600 = pi96  & n335;
  assign n4601 = ~n4599 & ~n4600;
  assign n4602 = ~n4598 & n4601;
  assign n4603 = n343 & n3946;
  assign n4604 = n4602 & ~n4603;
  assign n4605 = pi5  & ~n4604;
  assign n4606 = pi5  & ~n4605;
  assign n4607 = ~n4604 & ~n4605;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = ~n4548 & ~n4552;
  assign n4610 = pi94  & n493;
  assign n4611 = pi92  & n533;
  assign n4612 = pi93  & n488;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 = ~n4610 & n4613;
  assign n4615 = n496 & n3499;
  assign n4616 = n4614 & ~n4615;
  assign n4617 = pi8  & ~n4616;
  assign n4618 = pi8  & ~n4617;
  assign n4619 = ~n4616 & ~n4617;
  assign n4620 = ~n4618 & ~n4619;
  assign n4621 = ~n4532 & ~n4534;
  assign n4622 = ~n4526 & ~n4528;
  assign n4623 = pi88  & n918;
  assign n4624 = pi86  & n1031;
  assign n4625 = pi87  & n913;
  assign n4626 = ~n4624 & ~n4625;
  assign n4627 = ~n4623 & n4626;
  assign n4628 = n921 & n2277;
  assign n4629 = n4627 & ~n4628;
  assign n4630 = pi14  & ~n4629;
  assign n4631 = pi14  & ~n4630;
  assign n4632 = ~n4629 & ~n4630;
  assign n4633 = ~n4631 & ~n4632;
  assign n4634 = ~n4489 & ~n4493;
  assign n4635 = pi82  & n1582;
  assign n4636 = pi80  & n1713;
  assign n4637 = pi81  & n1577;
  assign n4638 = ~n4636 & ~n4637;
  assign n4639 = ~n4635 & n4638;
  assign n4640 = n1532 & n1585;
  assign n4641 = n4639 & ~n4640;
  assign n4642 = pi20  & ~n4641;
  assign n4643 = pi20  & ~n4642;
  assign n4644 = ~n4641 & ~n4642;
  assign n4645 = ~n4643 & ~n4644;
  assign n4646 = ~n4473 & ~n4475;
  assign n4647 = ~n4460 & ~n4463;
  assign n4648 = pi73  & n2976;
  assign n4649 = pi71  & n3182;
  assign n4650 = pi72  & n2971;
  assign n4651 = ~n4649 & ~n4650;
  assign n4652 = ~n4648 & n4651;
  assign n4653 = n639 & n2979;
  assign n4654 = n4652 & ~n4653;
  assign n4655 = pi29  & ~n4654;
  assign n4656 = pi29  & ~n4655;
  assign n4657 = ~n4654 & ~n4655;
  assign n4658 = ~n4656 & ~n4657;
  assign n4659 = pi67  & n4182;
  assign n4660 = pi65  & n4416;
  assign n4661 = pi66  & n4177;
  assign n4662 = ~n4660 & ~n4661;
  assign n4663 = ~n4659 & n4662;
  assign n4664 = n313 & n4185;
  assign n4665 = n4663 & ~n4664;
  assign n4666 = pi35  & ~n4665;
  assign n4667 = pi35  & ~n4666;
  assign n4668 = ~n4665 & ~n4666;
  assign n4669 = ~n4667 & ~n4668;
  assign n4670 = pi35  & ~pi36 ;
  assign n4671 = ~pi35  & pi36 ;
  assign n4672 = ~n4670 & ~n4671;
  assign n4673 = pi64  & ~n4672;
  assign n4674 = n4428 & n4673;
  assign n4675 = ~n4428 & ~n4673;
  assign n4676 = ~n4674 & ~n4675;
  assign n4677 = ~n4669 & n4676;
  assign n4678 = n4669 & ~n4676;
  assign n4679 = ~n4677 & ~n4678;
  assign n4680 = pi70  & n3550;
  assign n4681 = pi68  & n3735;
  assign n4682 = pi69  & n3545;
  assign n4683 = ~n4681 & ~n4682;
  assign n4684 = ~n4680 & n4683;
  assign n4685 = n430 & n3553;
  assign n4686 = n4684 & ~n4685;
  assign n4687 = pi32  & ~n4686;
  assign n4688 = pi32  & ~n4687;
  assign n4689 = ~n4686 & ~n4687;
  assign n4690 = ~n4688 & ~n4689;
  assign n4691 = n4679 & ~n4690;
  assign n4692 = ~n4679 & n4690;
  assign n4693 = ~n4691 & ~n4692;
  assign n4694 = ~n4446 & n4693;
  assign n4695 = n4446 & ~n4693;
  assign n4696 = ~n4694 & ~n4695;
  assign n4697 = ~n4658 & n4696;
  assign n4698 = n4658 & ~n4696;
  assign n4699 = ~n4697 & ~n4698;
  assign n4700 = n4647 & ~n4699;
  assign n4701 = ~n4647 & n4699;
  assign n4702 = ~n4700 & ~n4701;
  assign n4703 = pi76  & n2486;
  assign n4704 = pi74  & n2644;
  assign n4705 = pi75  & n2481;
  assign n4706 = ~n4704 & ~n4705;
  assign n4707 = ~n4703 & n4706;
  assign n4708 = n881 & n2489;
  assign n4709 = n4707 & ~n4708;
  assign n4710 = pi26  & ~n4709;
  assign n4711 = pi26  & ~n4710;
  assign n4712 = ~n4709 & ~n4710;
  assign n4713 = ~n4711 & ~n4712;
  assign n4714 = ~n4702 & n4713;
  assign n4715 = n4702 & ~n4713;
  assign n4716 = ~n4714 & ~n4715;
  assign n4717 = ~n4466 & ~n4469;
  assign n4718 = n4716 & ~n4717;
  assign n4719 = ~n4716 & n4717;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = pi79  & n2004;
  assign n4722 = pi77  & n2141;
  assign n4723 = pi78  & n1999;
  assign n4724 = ~n4722 & ~n4723;
  assign n4725 = ~n4721 & n4724;
  assign n4726 = n1105 & n2007;
  assign n4727 = n4725 & ~n4726;
  assign n4728 = pi23  & ~n4727;
  assign n4729 = pi23  & ~n4728;
  assign n4730 = ~n4727 & ~n4728;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = n4720 & ~n4731;
  assign n4733 = n4720 & ~n4732;
  assign n4734 = ~n4731 & ~n4732;
  assign n4735 = ~n4733 & ~n4734;
  assign n4736 = ~n4646 & ~n4735;
  assign n4737 = n4646 & n4735;
  assign n4738 = ~n4736 & ~n4737;
  assign n4739 = ~n4645 & n4738;
  assign n4740 = n4645 & ~n4738;
  assign n4741 = ~n4739 & ~n4740;
  assign n4742 = n4634 & ~n4741;
  assign n4743 = ~n4634 & n4741;
  assign n4744 = ~n4742 & ~n4743;
  assign n4745 = pi85  & n1269;
  assign n4746 = pi83  & n1340;
  assign n4747 = pi84  & n1264;
  assign n4748 = ~n4746 & ~n4747;
  assign n4749 = ~n4745 & n4748;
  assign n4750 = n1272 & n1943;
  assign n4751 = n4749 & ~n4750;
  assign n4752 = pi17  & ~n4751;
  assign n4753 = pi17  & ~n4752;
  assign n4754 = ~n4751 & ~n4752;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = n4744 & ~n4755;
  assign n4757 = ~n4744 & n4755;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = ~n4511 & n4758;
  assign n4760 = n4511 & ~n4758;
  assign n4761 = ~n4759 & ~n4760;
  assign n4762 = n4633 & ~n4761;
  assign n4763 = ~n4633 & n4761;
  assign n4764 = ~n4762 & ~n4763;
  assign n4765 = ~n4622 & n4764;
  assign n4766 = n4622 & ~n4764;
  assign n4767 = ~n4765 & ~n4766;
  assign n4768 = pi91  & n675;
  assign n4769 = pi89  & n769;
  assign n4770 = pi90  & n670;
  assign n4771 = ~n4769 & ~n4770;
  assign n4772 = ~n4768 & n4771;
  assign n4773 = n678 & n2926;
  assign n4774 = n4772 & ~n4773;
  assign n4775 = pi11  & ~n4774;
  assign n4776 = pi11  & ~n4775;
  assign n4777 = ~n4774 & ~n4775;
  assign n4778 = ~n4776 & ~n4777;
  assign n4779 = n4767 & ~n4778;
  assign n4780 = ~n4767 & n4778;
  assign n4781 = ~n4779 & ~n4780;
  assign n4782 = ~n4621 & n4781;
  assign n4783 = n4621 & ~n4781;
  assign n4784 = ~n4782 & ~n4783;
  assign n4785 = n4620 & ~n4784;
  assign n4786 = ~n4620 & n4784;
  assign n4787 = ~n4785 & ~n4786;
  assign n4788 = ~n4609 & n4787;
  assign n4789 = n4609 & ~n4787;
  assign n4790 = ~n4788 & ~n4789;
  assign n4791 = ~n4608 & n4790;
  assign n4792 = n4608 & ~n4790;
  assign n4793 = ~n4791 & ~n4792;
  assign n4794 = ~n4570 & n4793;
  assign n4795 = n4570 & ~n4793;
  assign n4796 = ~n4794 & ~n4795;
  assign n4797 = pi100  & n264;
  assign n4798 = pi98  & n281;
  assign n4799 = pi99  & n259;
  assign n4800 = ~n4798 & ~n4799;
  assign n4801 = ~n4797 & n4800;
  assign n4802 = ~n4580 & ~n4582;
  assign n4803 = ~pi99  & ~pi100 ;
  assign n4804 = pi99  & pi100 ;
  assign n4805 = ~n4803 & ~n4804;
  assign n4806 = ~n4802 & n4805;
  assign n4807 = n4802 & ~n4805;
  assign n4808 = ~n4806 & ~n4807;
  assign n4809 = n267 & n4808;
  assign n4810 = n4801 & ~n4809;
  assign n4811 = pi2  & ~n4810;
  assign n4812 = pi2  & ~n4811;
  assign n4813 = ~n4810 & ~n4811;
  assign n4814 = ~n4812 & ~n4813;
  assign n4815 = n4796 & ~n4814;
  assign n4816 = ~n4796 & n4814;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = ~n4597 & n4817;
  assign n4819 = n4597 & ~n4817;
  assign po36  = ~n4818 & ~n4819;
  assign n4821 = ~n4815 & ~n4818;
  assign n4822 = ~n4791 & ~n4794;
  assign n4823 = ~n4786 & ~n4788;
  assign n4824 = pi95  & n493;
  assign n4825 = pi93  & n533;
  assign n4826 = pi94  & n488;
  assign n4827 = ~n4825 & ~n4826;
  assign n4828 = ~n4824 & n4827;
  assign n4829 = n496 & n3710;
  assign n4830 = n4828 & ~n4829;
  assign n4831 = pi8  & ~n4830;
  assign n4832 = pi8  & ~n4831;
  assign n4833 = ~n4830 & ~n4831;
  assign n4834 = ~n4832 & ~n4833;
  assign n4835 = ~n4779 & ~n4782;
  assign n4836 = ~n4763 & ~n4765;
  assign n4837 = ~n4756 & ~n4759;
  assign n4838 = ~n4739 & ~n4743;
  assign n4839 = ~n4715 & ~n4718;
  assign n4840 = pi77  & n2486;
  assign n4841 = pi75  & n2644;
  assign n4842 = pi76  & n2481;
  assign n4843 = ~n4841 & ~n4842;
  assign n4844 = ~n4840 & n4843;
  assign n4845 = n984 & n2489;
  assign n4846 = n4844 & ~n4845;
  assign n4847 = pi26  & ~n4846;
  assign n4848 = pi26  & ~n4847;
  assign n4849 = ~n4846 & ~n4847;
  assign n4850 = ~n4848 & ~n4849;
  assign n4851 = ~n4697 & ~n4701;
  assign n4852 = pi74  & n2976;
  assign n4853 = pi72  & n3182;
  assign n4854 = pi73  & n2971;
  assign n4855 = ~n4853 & ~n4854;
  assign n4856 = ~n4852 & n4855;
  assign n4857 = n722 & n2979;
  assign n4858 = n4856 & ~n4857;
  assign n4859 = pi29  & ~n4858;
  assign n4860 = pi29  & ~n4859;
  assign n4861 = ~n4858 & ~n4859;
  assign n4862 = ~n4860 & ~n4861;
  assign n4863 = ~n4691 & ~n4694;
  assign n4864 = pi71  & n3550;
  assign n4865 = pi69  & n3735;
  assign n4866 = pi70  & n3545;
  assign n4867 = ~n4865 & ~n4866;
  assign n4868 = ~n4864 & n4867;
  assign n4869 = n476 & n3553;
  assign n4870 = n4868 & ~n4869;
  assign n4871 = pi32  & ~n4870;
  assign n4872 = pi32  & ~n4871;
  assign n4873 = ~n4870 & ~n4871;
  assign n4874 = ~n4872 & ~n4873;
  assign n4875 = ~n4674 & ~n4677;
  assign n4876 = pi68  & n4182;
  assign n4877 = pi66  & n4416;
  assign n4878 = pi67  & n4177;
  assign n4879 = ~n4877 & ~n4878;
  assign n4880 = ~n4876 & n4879;
  assign n4881 = n364 & n4185;
  assign n4882 = n4880 & ~n4881;
  assign n4883 = pi35  & ~n4882;
  assign n4884 = pi35  & ~n4883;
  assign n4885 = ~n4882 & ~n4883;
  assign n4886 = ~n4884 & ~n4885;
  assign n4887 = pi38  & ~n4673;
  assign n4888 = ~pi36  & pi37 ;
  assign n4889 = pi36  & ~pi37 ;
  assign n4890 = ~n4888 & ~n4889;
  assign n4891 = n4672 & ~n4890;
  assign n4892 = pi64  & n4891;
  assign n4893 = ~pi37  & pi38 ;
  assign n4894 = pi37  & ~pi38 ;
  assign n4895 = ~n4893 & ~n4894;
  assign n4896 = ~n4672 & n4895;
  assign n4897 = pi65  & n4896;
  assign n4898 = ~n4892 & ~n4897;
  assign n4899 = ~n4672 & ~n4895;
  assign n4900 = n270 & n4899;
  assign n4901 = n4898 & ~n4900;
  assign n4902 = pi38  & ~n4901;
  assign n4903 = pi38  & ~n4902;
  assign n4904 = ~n4901 & ~n4902;
  assign n4905 = ~n4903 & ~n4904;
  assign n4906 = n4887 & ~n4905;
  assign n4907 = ~n4887 & n4905;
  assign n4908 = ~n4906 & ~n4907;
  assign n4909 = n4886 & ~n4908;
  assign n4910 = ~n4886 & n4908;
  assign n4911 = ~n4909 & ~n4910;
  assign n4912 = ~n4875 & n4911;
  assign n4913 = n4875 & ~n4911;
  assign n4914 = ~n4912 & ~n4913;
  assign n4915 = n4874 & ~n4914;
  assign n4916 = ~n4874 & n4914;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = ~n4863 & n4917;
  assign n4919 = n4863 & ~n4917;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = n4862 & ~n4920;
  assign n4922 = ~n4862 & n4920;
  assign n4923 = ~n4921 & ~n4922;
  assign n4924 = ~n4851 & n4923;
  assign n4925 = n4851 & ~n4923;
  assign n4926 = ~n4924 & ~n4925;
  assign n4927 = n4850 & ~n4926;
  assign n4928 = ~n4850 & n4926;
  assign n4929 = ~n4927 & ~n4928;
  assign n4930 = ~n4839 & n4929;
  assign n4931 = n4839 & ~n4929;
  assign n4932 = ~n4930 & ~n4931;
  assign n4933 = pi80  & n2004;
  assign n4934 = pi78  & n2141;
  assign n4935 = pi79  & n1999;
  assign n4936 = ~n4934 & ~n4935;
  assign n4937 = ~n4933 & n4936;
  assign n4938 = n1205 & n2007;
  assign n4939 = n4937 & ~n4938;
  assign n4940 = pi23  & ~n4939;
  assign n4941 = pi23  & ~n4940;
  assign n4942 = ~n4939 & ~n4940;
  assign n4943 = ~n4941 & ~n4942;
  assign n4944 = n4932 & ~n4943;
  assign n4945 = n4932 & ~n4944;
  assign n4946 = ~n4943 & ~n4944;
  assign n4947 = ~n4945 & ~n4946;
  assign n4948 = ~n4732 & ~n4736;
  assign n4949 = n4947 & n4948;
  assign n4950 = ~n4947 & ~n4948;
  assign n4951 = ~n4949 & ~n4950;
  assign n4952 = pi83  & n1582;
  assign n4953 = pi81  & n1713;
  assign n4954 = pi82  & n1577;
  assign n4955 = ~n4953 & ~n4954;
  assign n4956 = ~n4952 & n4955;
  assign n4957 = n1585 & n1672;
  assign n4958 = n4956 & ~n4957;
  assign n4959 = pi20  & ~n4958;
  assign n4960 = pi20  & ~n4959;
  assign n4961 = ~n4958 & ~n4959;
  assign n4962 = ~n4960 & ~n4961;
  assign n4963 = n4951 & ~n4962;
  assign n4964 = ~n4951 & n4962;
  assign n4965 = ~n4963 & ~n4964;
  assign n4966 = n4838 & ~n4965;
  assign n4967 = ~n4838 & n4965;
  assign n4968 = ~n4966 & ~n4967;
  assign n4969 = pi86  & n1269;
  assign n4970 = pi84  & n1340;
  assign n4971 = pi85  & n1264;
  assign n4972 = ~n4970 & ~n4971;
  assign n4973 = ~n4969 & n4972;
  assign n4974 = n1272 & n2099;
  assign n4975 = n4973 & ~n4974;
  assign n4976 = pi17  & ~n4975;
  assign n4977 = pi17  & ~n4976;
  assign n4978 = ~n4975 & ~n4976;
  assign n4979 = ~n4977 & ~n4978;
  assign n4980 = n4968 & ~n4979;
  assign n4981 = ~n4968 & n4979;
  assign n4982 = ~n4980 & ~n4981;
  assign n4983 = n4837 & ~n4982;
  assign n4984 = ~n4837 & n4982;
  assign n4985 = ~n4983 & ~n4984;
  assign n4986 = pi89  & n918;
  assign n4987 = pi87  & n1031;
  assign n4988 = pi88  & n913;
  assign n4989 = ~n4987 & ~n4988;
  assign n4990 = ~n4986 & n4989;
  assign n4991 = n921 & n2432;
  assign n4992 = n4990 & ~n4991;
  assign n4993 = pi14  & ~n4992;
  assign n4994 = pi14  & ~n4993;
  assign n4995 = ~n4992 & ~n4993;
  assign n4996 = ~n4994 & ~n4995;
  assign n4997 = n4985 & ~n4996;
  assign n4998 = ~n4985 & n4996;
  assign n4999 = ~n4836 & ~n4998;
  assign n5000 = ~n4997 & n4999;
  assign n5001 = ~n4836 & ~n5000;
  assign n5002 = ~n4997 & ~n5000;
  assign n5003 = ~n4998 & n5002;
  assign n5004 = ~n5001 & ~n5003;
  assign n5005 = pi92  & n675;
  assign n5006 = pi90  & n769;
  assign n5007 = pi91  & n670;
  assign n5008 = ~n5006 & ~n5007;
  assign n5009 = ~n5005 & n5008;
  assign n5010 = n678 & n3119;
  assign n5011 = n5009 & ~n5010;
  assign n5012 = pi11  & ~n5011;
  assign n5013 = pi11  & ~n5012;
  assign n5014 = ~n5011 & ~n5012;
  assign n5015 = ~n5013 & ~n5014;
  assign n5016 = n5004 & n5015;
  assign n5017 = ~n5004 & ~n5015;
  assign n5018 = ~n5016 & ~n5017;
  assign n5019 = ~n4835 & n5018;
  assign n5020 = n4835 & ~n5018;
  assign n5021 = ~n5019 & ~n5020;
  assign n5022 = n4834 & ~n5021;
  assign n5023 = ~n4834 & n5021;
  assign n5024 = ~n5022 & ~n5023;
  assign n5025 = ~n4823 & n5024;
  assign n5026 = n4823 & ~n5024;
  assign n5027 = ~n5025 & ~n5026;
  assign n5028 = pi98  & n340;
  assign n5029 = pi96  & n380;
  assign n5030 = pi97  & n335;
  assign n5031 = ~n5029 & ~n5030;
  assign n5032 = ~n5028 & n5031;
  assign n5033 = n343 & n4360;
  assign n5034 = n5032 & ~n5033;
  assign n5035 = pi5  & ~n5034;
  assign n5036 = pi5  & ~n5035;
  assign n5037 = ~n5034 & ~n5035;
  assign n5038 = ~n5036 & ~n5037;
  assign n5039 = n5027 & ~n5038;
  assign n5040 = ~n5027 & n5038;
  assign n5041 = ~n5039 & ~n5040;
  assign n5042 = n4822 & ~n5041;
  assign n5043 = ~n4822 & n5041;
  assign n5044 = ~n5042 & ~n5043;
  assign n5045 = pi101  & n264;
  assign n5046 = pi99  & n281;
  assign n5047 = pi100  & n259;
  assign n5048 = ~n5046 & ~n5047;
  assign n5049 = ~n5045 & n5048;
  assign n5050 = ~n4804 & ~n4806;
  assign n5051 = ~pi100  & ~pi101 ;
  assign n5052 = pi100  & pi101 ;
  assign n5053 = ~n5051 & ~n5052;
  assign n5054 = ~n5050 & n5053;
  assign n5055 = n5050 & ~n5053;
  assign n5056 = ~n5054 & ~n5055;
  assign n5057 = n267 & n5056;
  assign n5058 = n5049 & ~n5057;
  assign n5059 = pi2  & ~n5058;
  assign n5060 = pi2  & ~n5059;
  assign n5061 = ~n5058 & ~n5059;
  assign n5062 = ~n5060 & ~n5061;
  assign n5063 = ~n5044 & n5062;
  assign n5064 = n5044 & ~n5062;
  assign n5065 = ~n5063 & ~n5064;
  assign n5066 = ~n4821 & n5065;
  assign n5067 = n4821 & ~n5065;
  assign po37  = ~n5066 & ~n5067;
  assign n5069 = ~n5064 & ~n5066;
  assign n5070 = ~n5039 & ~n5043;
  assign n5071 = pi99  & n340;
  assign n5072 = pi97  & n380;
  assign n5073 = pi98  & n335;
  assign n5074 = ~n5072 & ~n5073;
  assign n5075 = ~n5071 & n5074;
  assign n5076 = n343 & n4584;
  assign n5077 = n5075 & ~n5076;
  assign n5078 = pi5  & ~n5077;
  assign n5079 = pi5  & ~n5078;
  assign n5080 = ~n5077 & ~n5078;
  assign n5081 = ~n5079 & ~n5080;
  assign n5082 = ~n5023 & ~n5025;
  assign n5083 = pi96  & n493;
  assign n5084 = pi94  & n533;
  assign n5085 = pi95  & n488;
  assign n5086 = ~n5084 & ~n5085;
  assign n5087 = ~n5083 & n5086;
  assign n5088 = n496 & n3921;
  assign n5089 = n5087 & ~n5088;
  assign n5090 = pi8  & ~n5089;
  assign n5091 = pi8  & ~n5090;
  assign n5092 = ~n5089 & ~n5090;
  assign n5093 = ~n5091 & ~n5092;
  assign n5094 = ~n5017 & ~n5019;
  assign n5095 = pi93  & n675;
  assign n5096 = pi91  & n769;
  assign n5097 = pi92  & n670;
  assign n5098 = ~n5096 & ~n5097;
  assign n5099 = ~n5095 & n5098;
  assign n5100 = n678 & n3144;
  assign n5101 = n5099 & ~n5100;
  assign n5102 = pi11  & ~n5101;
  assign n5103 = pi11  & ~n5102;
  assign n5104 = ~n5101 & ~n5102;
  assign n5105 = ~n5103 & ~n5104;
  assign n5106 = ~n4980 & ~n4984;
  assign n5107 = ~n4963 & ~n4967;
  assign n5108 = ~n4944 & ~n4950;
  assign n5109 = ~n4928 & ~n4930;
  assign n5110 = pi78  & n2486;
  assign n5111 = pi76  & n2644;
  assign n5112 = pi77  & n2481;
  assign n5113 = ~n5111 & ~n5112;
  assign n5114 = ~n5110 & n5113;
  assign n5115 = n1009 & n2489;
  assign n5116 = n5114 & ~n5115;
  assign n5117 = pi26  & ~n5116;
  assign n5118 = pi26  & ~n5117;
  assign n5119 = ~n5116 & ~n5117;
  assign n5120 = ~n5118 & ~n5119;
  assign n5121 = ~n4922 & ~n4924;
  assign n5122 = pi75  & n2976;
  assign n5123 = pi73  & n3182;
  assign n5124 = pi74  & n2971;
  assign n5125 = ~n5123 & ~n5124;
  assign n5126 = ~n5122 & n5125;
  assign n5127 = n747 & n2979;
  assign n5128 = n5126 & ~n5127;
  assign n5129 = pi29  & ~n5128;
  assign n5130 = pi29  & ~n5129;
  assign n5131 = ~n5128 & ~n5129;
  assign n5132 = ~n5130 & ~n5131;
  assign n5133 = ~n4916 & ~n4918;
  assign n5134 = pi72  & n3550;
  assign n5135 = pi70  & n3735;
  assign n5136 = pi71  & n3545;
  assign n5137 = ~n5135 & ~n5136;
  assign n5138 = ~n5134 & n5137;
  assign n5139 = n575 & n3553;
  assign n5140 = n5138 & ~n5139;
  assign n5141 = pi32  & ~n5140;
  assign n5142 = pi32  & ~n5141;
  assign n5143 = ~n5140 & ~n5141;
  assign n5144 = ~n5142 & ~n5143;
  assign n5145 = ~n4910 & ~n4912;
  assign n5146 = pi66  & n4896;
  assign n5147 = n4672 & ~n4895;
  assign n5148 = n4890 & n5147;
  assign n5149 = pi64  & n5148;
  assign n5150 = pi65  & n4891;
  assign n5151 = ~n5149 & ~n5150;
  assign n5152 = ~n5146 & n5151;
  assign n5153 = n291 & n4899;
  assign n5154 = n5152 & ~n5153;
  assign n5155 = pi38  & ~n5154;
  assign n5156 = pi38  & ~n5155;
  assign n5157 = ~n5154 & ~n5155;
  assign n5158 = ~n5156 & ~n5157;
  assign n5159 = ~n4906 & n5158;
  assign n5160 = n4906 & ~n5158;
  assign n5161 = ~n5159 & ~n5160;
  assign n5162 = pi69  & n4182;
  assign n5163 = pi67  & n4416;
  assign n5164 = pi68  & n4177;
  assign n5165 = ~n5163 & ~n5164;
  assign n5166 = ~n5162 & n5165;
  assign n5167 = n405 & n4185;
  assign n5168 = n5166 & ~n5167;
  assign n5169 = pi35  & ~n5168;
  assign n5170 = pi35  & ~n5169;
  assign n5171 = ~n5168 & ~n5169;
  assign n5172 = ~n5170 & ~n5171;
  assign n5173 = n5161 & ~n5172;
  assign n5174 = ~n5161 & n5172;
  assign n5175 = ~n5173 & ~n5174;
  assign n5176 = ~n5145 & n5175;
  assign n5177 = n5145 & ~n5175;
  assign n5178 = ~n5176 & ~n5177;
  assign n5179 = ~n5144 & n5178;
  assign n5180 = n5144 & ~n5178;
  assign n5181 = ~n5179 & ~n5180;
  assign n5182 = ~n5133 & n5181;
  assign n5183 = n5133 & ~n5181;
  assign n5184 = ~n5182 & ~n5183;
  assign n5185 = ~n5132 & n5184;
  assign n5186 = n5132 & ~n5184;
  assign n5187 = ~n5185 & ~n5186;
  assign n5188 = ~n5121 & n5187;
  assign n5189 = n5121 & ~n5187;
  assign n5190 = ~n5188 & ~n5189;
  assign n5191 = n5120 & ~n5190;
  assign n5192 = ~n5120 & n5190;
  assign n5193 = ~n5191 & ~n5192;
  assign n5194 = ~n5109 & n5193;
  assign n5195 = n5109 & ~n5193;
  assign n5196 = ~n5194 & ~n5195;
  assign n5197 = pi81  & n2004;
  assign n5198 = pi79  & n2141;
  assign n5199 = pi80  & n1999;
  assign n5200 = ~n5198 & ~n5199;
  assign n5201 = ~n5197 & n5200;
  assign n5202 = n1413 & n2007;
  assign n5203 = n5201 & ~n5202;
  assign n5204 = pi23  & ~n5203;
  assign n5205 = pi23  & ~n5204;
  assign n5206 = ~n5203 & ~n5204;
  assign n5207 = ~n5205 & ~n5206;
  assign n5208 = n5196 & ~n5207;
  assign n5209 = ~n5196 & n5207;
  assign n5210 = ~n5208 & ~n5209;
  assign n5211 = n5108 & ~n5210;
  assign n5212 = ~n5108 & n5210;
  assign n5213 = ~n5211 & ~n5212;
  assign n5214 = pi84  & n1582;
  assign n5215 = pi82  & n1713;
  assign n5216 = pi83  & n1577;
  assign n5217 = ~n5215 & ~n5216;
  assign n5218 = ~n5214 & n5217;
  assign n5219 = n1585 & n1805;
  assign n5220 = n5218 & ~n5219;
  assign n5221 = pi20  & ~n5220;
  assign n5222 = pi20  & ~n5221;
  assign n5223 = ~n5220 & ~n5221;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = n5213 & ~n5224;
  assign n5226 = ~n5213 & n5224;
  assign n5227 = ~n5225 & ~n5226;
  assign n5228 = n5107 & ~n5227;
  assign n5229 = ~n5107 & n5227;
  assign n5230 = ~n5228 & ~n5229;
  assign n5231 = pi87  & n1269;
  assign n5232 = pi85  & n1340;
  assign n5233 = pi86  & n1264;
  assign n5234 = ~n5232 & ~n5233;
  assign n5235 = ~n5231 & n5234;
  assign n5236 = n1272 & n2252;
  assign n5237 = n5235 & ~n5236;
  assign n5238 = pi17  & ~n5237;
  assign n5239 = pi17  & ~n5238;
  assign n5240 = ~n5237 & ~n5238;
  assign n5241 = ~n5239 & ~n5240;
  assign n5242 = n5230 & ~n5241;
  assign n5243 = ~n5230 & n5241;
  assign n5244 = ~n5106 & ~n5243;
  assign n5245 = ~n5242 & n5244;
  assign n5246 = ~n5106 & ~n5245;
  assign n5247 = ~n5242 & ~n5245;
  assign n5248 = ~n5243 & n5247;
  assign n5249 = ~n5246 & ~n5248;
  assign n5250 = pi90  & n918;
  assign n5251 = pi88  & n1031;
  assign n5252 = pi89  & n913;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = ~n5250 & n5253;
  assign n5255 = n921 & n2606;
  assign n5256 = n5254 & ~n5255;
  assign n5257 = pi14  & ~n5256;
  assign n5258 = pi14  & ~n5257;
  assign n5259 = ~n5256 & ~n5257;
  assign n5260 = ~n5258 & ~n5259;
  assign n5261 = n5249 & n5260;
  assign n5262 = ~n5249 & ~n5260;
  assign n5263 = ~n5261 & ~n5262;
  assign n5264 = ~n5002 & n5263;
  assign n5265 = n5002 & ~n5263;
  assign n5266 = ~n5264 & ~n5265;
  assign n5267 = n5105 & ~n5266;
  assign n5268 = ~n5105 & n5266;
  assign n5269 = ~n5267 & ~n5268;
  assign n5270 = ~n5094 & n5269;
  assign n5271 = n5094 & ~n5269;
  assign n5272 = ~n5270 & ~n5271;
  assign n5273 = n5093 & ~n5272;
  assign n5274 = ~n5093 & n5272;
  assign n5275 = ~n5273 & ~n5274;
  assign n5276 = ~n5082 & n5275;
  assign n5277 = n5082 & ~n5275;
  assign n5278 = ~n5276 & ~n5277;
  assign n5279 = n5081 & ~n5278;
  assign n5280 = ~n5081 & n5278;
  assign n5281 = ~n5279 & ~n5280;
  assign n5282 = ~n5070 & n5281;
  assign n5283 = n5070 & ~n5281;
  assign n5284 = ~n5282 & ~n5283;
  assign n5285 = pi102  & n264;
  assign n5286 = pi100  & n281;
  assign n5287 = pi101  & n259;
  assign n5288 = ~n5286 & ~n5287;
  assign n5289 = ~n5285 & n5288;
  assign n5290 = ~n5052 & ~n5054;
  assign n5291 = ~pi101  & ~pi102 ;
  assign n5292 = pi101  & pi102 ;
  assign n5293 = ~n5291 & ~n5292;
  assign n5294 = ~n5290 & n5293;
  assign n5295 = n5290 & ~n5293;
  assign n5296 = ~n5294 & ~n5295;
  assign n5297 = n267 & n5296;
  assign n5298 = n5289 & ~n5297;
  assign n5299 = pi2  & ~n5298;
  assign n5300 = pi2  & ~n5299;
  assign n5301 = ~n5298 & ~n5299;
  assign n5302 = ~n5300 & ~n5301;
  assign n5303 = n5284 & ~n5302;
  assign n5304 = ~n5284 & n5302;
  assign n5305 = ~n5303 & ~n5304;
  assign n5306 = ~n5069 & n5305;
  assign n5307 = n5069 & ~n5305;
  assign po38  = ~n5306 & ~n5307;
  assign n5309 = ~n5303 & ~n5306;
  assign n5310 = ~n5280 & ~n5282;
  assign n5311 = pi100  & n340;
  assign n5312 = pi98  & n380;
  assign n5313 = pi99  & n335;
  assign n5314 = ~n5312 & ~n5313;
  assign n5315 = ~n5311 & n5314;
  assign n5316 = n343 & n4808;
  assign n5317 = n5315 & ~n5316;
  assign n5318 = pi5  & ~n5317;
  assign n5319 = pi5  & ~n5318;
  assign n5320 = ~n5317 & ~n5318;
  assign n5321 = ~n5319 & ~n5320;
  assign n5322 = ~n5274 & ~n5276;
  assign n5323 = ~n5268 & ~n5270;
  assign n5324 = pi94  & n675;
  assign n5325 = pi92  & n769;
  assign n5326 = pi93  & n670;
  assign n5327 = ~n5325 & ~n5326;
  assign n5328 = ~n5324 & n5327;
  assign n5329 = n678 & n3499;
  assign n5330 = n5328 & ~n5329;
  assign n5331 = pi11  & ~n5330;
  assign n5332 = pi11  & ~n5331;
  assign n5333 = ~n5330 & ~n5331;
  assign n5334 = ~n5332 & ~n5333;
  assign n5335 = ~n5262 & ~n5264;
  assign n5336 = ~n5225 & ~n5229;
  assign n5337 = ~n5208 & ~n5212;
  assign n5338 = pi82  & n2004;
  assign n5339 = pi80  & n2141;
  assign n5340 = pi81  & n1999;
  assign n5341 = ~n5339 & ~n5340;
  assign n5342 = ~n5338 & n5341;
  assign n5343 = n1532 & n2007;
  assign n5344 = n5342 & ~n5343;
  assign n5345 = pi23  & ~n5344;
  assign n5346 = pi23  & ~n5345;
  assign n5347 = ~n5344 & ~n5345;
  assign n5348 = ~n5346 & ~n5347;
  assign n5349 = ~n5192 & ~n5194;
  assign n5350 = ~n5179 & ~n5182;
  assign n5351 = ~n5173 & ~n5176;
  assign n5352 = pi67  & n4896;
  assign n5353 = pi65  & n5148;
  assign n5354 = pi66  & n4891;
  assign n5355 = ~n5353 & ~n5354;
  assign n5356 = ~n5352 & n5355;
  assign n5357 = n313 & n4899;
  assign n5358 = n5356 & ~n5357;
  assign n5359 = pi38  & ~n5358;
  assign n5360 = pi38  & ~n5359;
  assign n5361 = ~n5358 & ~n5359;
  assign n5362 = ~n5360 & ~n5361;
  assign n5363 = pi38  & ~pi39 ;
  assign n5364 = ~pi38  & pi39 ;
  assign n5365 = ~n5363 & ~n5364;
  assign n5366 = pi64  & ~n5365;
  assign n5367 = n5160 & n5366;
  assign n5368 = ~n5160 & ~n5366;
  assign n5369 = ~n5367 & ~n5368;
  assign n5370 = ~n5362 & n5369;
  assign n5371 = n5362 & ~n5369;
  assign n5372 = ~n5370 & ~n5371;
  assign n5373 = pi70  & n4182;
  assign n5374 = pi68  & n4416;
  assign n5375 = pi69  & n4177;
  assign n5376 = ~n5374 & ~n5375;
  assign n5377 = ~n5373 & n5376;
  assign n5378 = n430 & n4185;
  assign n5379 = n5377 & ~n5378;
  assign n5380 = pi35  & ~n5379;
  assign n5381 = pi35  & ~n5380;
  assign n5382 = ~n5379 & ~n5380;
  assign n5383 = ~n5381 & ~n5382;
  assign n5384 = n5372 & ~n5383;
  assign n5385 = ~n5372 & n5383;
  assign n5386 = ~n5384 & ~n5385;
  assign n5387 = n5351 & ~n5386;
  assign n5388 = ~n5351 & n5386;
  assign n5389 = ~n5387 & ~n5388;
  assign n5390 = pi73  & n3550;
  assign n5391 = pi71  & n3735;
  assign n5392 = pi72  & n3545;
  assign n5393 = ~n5391 & ~n5392;
  assign n5394 = ~n5390 & n5393;
  assign n5395 = n639 & n3553;
  assign n5396 = n5394 & ~n5395;
  assign n5397 = pi32  & ~n5396;
  assign n5398 = pi32  & ~n5397;
  assign n5399 = ~n5396 & ~n5397;
  assign n5400 = ~n5398 & ~n5399;
  assign n5401 = n5389 & ~n5400;
  assign n5402 = ~n5389 & n5400;
  assign n5403 = ~n5401 & ~n5402;
  assign n5404 = n5350 & ~n5403;
  assign n5405 = ~n5350 & n5403;
  assign n5406 = ~n5404 & ~n5405;
  assign n5407 = pi76  & n2976;
  assign n5408 = pi74  & n3182;
  assign n5409 = pi75  & n2971;
  assign n5410 = ~n5408 & ~n5409;
  assign n5411 = ~n5407 & n5410;
  assign n5412 = n881 & n2979;
  assign n5413 = n5411 & ~n5412;
  assign n5414 = pi29  & ~n5413;
  assign n5415 = pi29  & ~n5414;
  assign n5416 = ~n5413 & ~n5414;
  assign n5417 = ~n5415 & ~n5416;
  assign n5418 = ~n5406 & n5417;
  assign n5419 = n5406 & ~n5417;
  assign n5420 = ~n5418 & ~n5419;
  assign n5421 = ~n5185 & ~n5188;
  assign n5422 = n5420 & ~n5421;
  assign n5423 = ~n5420 & n5421;
  assign n5424 = ~n5422 & ~n5423;
  assign n5425 = pi79  & n2486;
  assign n5426 = pi77  & n2644;
  assign n5427 = pi78  & n2481;
  assign n5428 = ~n5426 & ~n5427;
  assign n5429 = ~n5425 & n5428;
  assign n5430 = n1105 & n2489;
  assign n5431 = n5429 & ~n5430;
  assign n5432 = pi26  & ~n5431;
  assign n5433 = pi26  & ~n5432;
  assign n5434 = ~n5431 & ~n5432;
  assign n5435 = ~n5433 & ~n5434;
  assign n5436 = n5424 & ~n5435;
  assign n5437 = n5424 & ~n5436;
  assign n5438 = ~n5435 & ~n5436;
  assign n5439 = ~n5437 & ~n5438;
  assign n5440 = ~n5349 & ~n5439;
  assign n5441 = n5349 & n5439;
  assign n5442 = ~n5440 & ~n5441;
  assign n5443 = ~n5348 & n5442;
  assign n5444 = n5348 & ~n5442;
  assign n5445 = ~n5443 & ~n5444;
  assign n5446 = n5337 & ~n5445;
  assign n5447 = ~n5337 & n5445;
  assign n5448 = ~n5446 & ~n5447;
  assign n5449 = pi85  & n1582;
  assign n5450 = pi83  & n1713;
  assign n5451 = pi84  & n1577;
  assign n5452 = ~n5450 & ~n5451;
  assign n5453 = ~n5449 & n5452;
  assign n5454 = n1585 & n1943;
  assign n5455 = n5453 & ~n5454;
  assign n5456 = pi20  & ~n5455;
  assign n5457 = pi20  & ~n5456;
  assign n5458 = ~n5455 & ~n5456;
  assign n5459 = ~n5457 & ~n5458;
  assign n5460 = n5448 & ~n5459;
  assign n5461 = ~n5448 & n5459;
  assign n5462 = ~n5460 & ~n5461;
  assign n5463 = n5336 & ~n5462;
  assign n5464 = ~n5336 & n5462;
  assign n5465 = ~n5463 & ~n5464;
  assign n5466 = pi88  & n1269;
  assign n5467 = pi86  & n1340;
  assign n5468 = pi87  & n1264;
  assign n5469 = ~n5467 & ~n5468;
  assign n5470 = ~n5466 & n5469;
  assign n5471 = n1272 & n2277;
  assign n5472 = n5470 & ~n5471;
  assign n5473 = pi17  & ~n5472;
  assign n5474 = pi17  & ~n5473;
  assign n5475 = ~n5472 & ~n5473;
  assign n5476 = ~n5474 & ~n5475;
  assign n5477 = ~n5465 & n5476;
  assign n5478 = n5465 & ~n5476;
  assign n5479 = ~n5477 & ~n5478;
  assign n5480 = ~n5247 & n5479;
  assign n5481 = n5247 & ~n5479;
  assign n5482 = ~n5480 & ~n5481;
  assign n5483 = pi91  & n918;
  assign n5484 = pi89  & n1031;
  assign n5485 = pi90  & n913;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = ~n5483 & n5486;
  assign n5488 = n921 & n2926;
  assign n5489 = n5487 & ~n5488;
  assign n5490 = pi14  & ~n5489;
  assign n5491 = pi14  & ~n5490;
  assign n5492 = ~n5489 & ~n5490;
  assign n5493 = ~n5491 & ~n5492;
  assign n5494 = n5482 & ~n5493;
  assign n5495 = ~n5482 & n5493;
  assign n5496 = ~n5494 & ~n5495;
  assign n5497 = ~n5335 & n5496;
  assign n5498 = n5335 & ~n5496;
  assign n5499 = ~n5497 & ~n5498;
  assign n5500 = ~n5334 & n5499;
  assign n5501 = n5334 & ~n5499;
  assign n5502 = ~n5500 & ~n5501;
  assign n5503 = ~n5323 & n5502;
  assign n5504 = n5323 & ~n5502;
  assign n5505 = ~n5503 & ~n5504;
  assign n5506 = pi97  & n493;
  assign n5507 = pi95  & n533;
  assign n5508 = pi96  & n488;
  assign n5509 = ~n5507 & ~n5508;
  assign n5510 = ~n5506 & n5509;
  assign n5511 = n496 & n3946;
  assign n5512 = n5510 & ~n5511;
  assign n5513 = pi8  & ~n5512;
  assign n5514 = pi8  & ~n5513;
  assign n5515 = ~n5512 & ~n5513;
  assign n5516 = ~n5514 & ~n5515;
  assign n5517 = n5505 & ~n5516;
  assign n5518 = ~n5505 & n5516;
  assign n5519 = ~n5517 & ~n5518;
  assign n5520 = ~n5322 & n5519;
  assign n5521 = n5322 & ~n5519;
  assign n5522 = ~n5520 & ~n5521;
  assign n5523 = n5321 & ~n5522;
  assign n5524 = ~n5321 & n5522;
  assign n5525 = ~n5523 & ~n5524;
  assign n5526 = ~n5310 & n5525;
  assign n5527 = n5310 & ~n5525;
  assign n5528 = ~n5526 & ~n5527;
  assign n5529 = pi103  & n264;
  assign n5530 = pi101  & n281;
  assign n5531 = pi102  & n259;
  assign n5532 = ~n5530 & ~n5531;
  assign n5533 = ~n5529 & n5532;
  assign n5534 = ~n5292 & ~n5294;
  assign n5535 = ~pi102  & ~pi103 ;
  assign n5536 = pi102  & pi103 ;
  assign n5537 = ~n5535 & ~n5536;
  assign n5538 = ~n5534 & n5537;
  assign n5539 = n5534 & ~n5537;
  assign n5540 = ~n5538 & ~n5539;
  assign n5541 = n267 & n5540;
  assign n5542 = n5533 & ~n5541;
  assign n5543 = pi2  & ~n5542;
  assign n5544 = pi2  & ~n5543;
  assign n5545 = ~n5542 & ~n5543;
  assign n5546 = ~n5544 & ~n5545;
  assign n5547 = n5528 & ~n5546;
  assign n5548 = ~n5528 & n5546;
  assign n5549 = ~n5547 & ~n5548;
  assign n5550 = ~n5309 & n5549;
  assign n5551 = n5309 & ~n5549;
  assign po39  = ~n5550 & ~n5551;
  assign n5553 = ~n5547 & ~n5550;
  assign n5554 = pi104  & n264;
  assign n5555 = pi102  & n281;
  assign n5556 = pi103  & n259;
  assign n5557 = ~n5555 & ~n5556;
  assign n5558 = ~n5554 & n5557;
  assign n5559 = ~n5536 & ~n5538;
  assign n5560 = ~pi103  & ~pi104 ;
  assign n5561 = pi103  & pi104 ;
  assign n5562 = ~n5560 & ~n5561;
  assign n5563 = ~n5559 & n5562;
  assign n5564 = n5559 & ~n5562;
  assign n5565 = ~n5563 & ~n5564;
  assign n5566 = n267 & n5565;
  assign n5567 = n5558 & ~n5566;
  assign n5568 = pi2  & ~n5567;
  assign n5569 = pi2  & ~n5568;
  assign n5570 = ~n5567 & ~n5568;
  assign n5571 = ~n5569 & ~n5570;
  assign n5572 = ~n5524 & ~n5526;
  assign n5573 = ~n5517 & ~n5520;
  assign n5574 = pi98  & n493;
  assign n5575 = pi96  & n533;
  assign n5576 = pi97  & n488;
  assign n5577 = ~n5575 & ~n5576;
  assign n5578 = ~n5574 & n5577;
  assign n5579 = n496 & n4360;
  assign n5580 = n5578 & ~n5579;
  assign n5581 = pi8  & ~n5580;
  assign n5582 = pi8  & ~n5581;
  assign n5583 = ~n5580 & ~n5581;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = ~n5500 & ~n5503;
  assign n5586 = pi95  & n675;
  assign n5587 = pi93  & n769;
  assign n5588 = pi94  & n670;
  assign n5589 = ~n5587 & ~n5588;
  assign n5590 = ~n5586 & n5589;
  assign n5591 = n678 & n3710;
  assign n5592 = n5590 & ~n5591;
  assign n5593 = pi11  & ~n5592;
  assign n5594 = pi11  & ~n5593;
  assign n5595 = ~n5592 & ~n5593;
  assign n5596 = ~n5594 & ~n5595;
  assign n5597 = ~n5494 & ~n5497;
  assign n5598 = pi92  & n918;
  assign n5599 = pi90  & n1031;
  assign n5600 = pi91  & n913;
  assign n5601 = ~n5599 & ~n5600;
  assign n5602 = ~n5598 & n5601;
  assign n5603 = n921 & n3119;
  assign n5604 = n5602 & ~n5603;
  assign n5605 = pi14  & ~n5604;
  assign n5606 = pi14  & ~n5605;
  assign n5607 = ~n5604 & ~n5605;
  assign n5608 = ~n5606 & ~n5607;
  assign n5609 = ~n5478 & ~n5480;
  assign n5610 = ~n5460 & ~n5464;
  assign n5611 = ~n5436 & ~n5440;
  assign n5612 = ~n5419 & ~n5422;
  assign n5613 = ~n5401 & ~n5405;
  assign n5614 = ~n5384 & ~n5388;
  assign n5615 = ~n5367 & ~n5370;
  assign n5616 = pi68  & n4896;
  assign n5617 = pi66  & n5148;
  assign n5618 = pi67  & n4891;
  assign n5619 = ~n5617 & ~n5618;
  assign n5620 = ~n5616 & n5619;
  assign n5621 = n364 & n4899;
  assign n5622 = n5620 & ~n5621;
  assign n5623 = pi38  & ~n5622;
  assign n5624 = pi38  & ~n5623;
  assign n5625 = ~n5622 & ~n5623;
  assign n5626 = ~n5624 & ~n5625;
  assign n5627 = pi41  & ~n5366;
  assign n5628 = ~pi39  & pi40 ;
  assign n5629 = pi39  & ~pi40 ;
  assign n5630 = ~n5628 & ~n5629;
  assign n5631 = n5365 & ~n5630;
  assign n5632 = pi64  & n5631;
  assign n5633 = ~pi40  & pi41 ;
  assign n5634 = pi40  & ~pi41 ;
  assign n5635 = ~n5633 & ~n5634;
  assign n5636 = ~n5365 & n5635;
  assign n5637 = pi65  & n5636;
  assign n5638 = ~n5632 & ~n5637;
  assign n5639 = ~n5365 & ~n5635;
  assign n5640 = n270 & n5639;
  assign n5641 = n5638 & ~n5640;
  assign n5642 = pi41  & ~n5641;
  assign n5643 = pi41  & ~n5642;
  assign n5644 = ~n5641 & ~n5642;
  assign n5645 = ~n5643 & ~n5644;
  assign n5646 = n5627 & ~n5645;
  assign n5647 = ~n5627 & n5645;
  assign n5648 = ~n5646 & ~n5647;
  assign n5649 = n5626 & ~n5648;
  assign n5650 = ~n5626 & n5648;
  assign n5651 = ~n5649 & ~n5650;
  assign n5652 = ~n5615 & n5651;
  assign n5653 = n5615 & ~n5651;
  assign n5654 = ~n5652 & ~n5653;
  assign n5655 = pi71  & n4182;
  assign n5656 = pi69  & n4416;
  assign n5657 = pi70  & n4177;
  assign n5658 = ~n5656 & ~n5657;
  assign n5659 = ~n5655 & n5658;
  assign n5660 = n476 & n4185;
  assign n5661 = n5659 & ~n5660;
  assign n5662 = pi35  & ~n5661;
  assign n5663 = pi35  & ~n5662;
  assign n5664 = ~n5661 & ~n5662;
  assign n5665 = ~n5663 & ~n5664;
  assign n5666 = n5654 & ~n5665;
  assign n5667 = ~n5654 & n5665;
  assign n5668 = ~n5666 & ~n5667;
  assign n5669 = n5614 & ~n5668;
  assign n5670 = ~n5614 & n5668;
  assign n5671 = ~n5669 & ~n5670;
  assign n5672 = pi74  & n3550;
  assign n5673 = pi72  & n3735;
  assign n5674 = pi73  & n3545;
  assign n5675 = ~n5673 & ~n5674;
  assign n5676 = ~n5672 & n5675;
  assign n5677 = n722 & n3553;
  assign n5678 = n5676 & ~n5677;
  assign n5679 = pi32  & ~n5678;
  assign n5680 = pi32  & ~n5679;
  assign n5681 = ~n5678 & ~n5679;
  assign n5682 = ~n5680 & ~n5681;
  assign n5683 = n5671 & ~n5682;
  assign n5684 = ~n5671 & n5682;
  assign n5685 = ~n5613 & ~n5684;
  assign n5686 = ~n5683 & n5685;
  assign n5687 = ~n5613 & ~n5686;
  assign n5688 = ~n5683 & ~n5686;
  assign n5689 = ~n5684 & n5688;
  assign n5690 = ~n5687 & ~n5689;
  assign n5691 = pi77  & n2976;
  assign n5692 = pi75  & n3182;
  assign n5693 = pi76  & n2971;
  assign n5694 = ~n5692 & ~n5693;
  assign n5695 = ~n5691 & n5694;
  assign n5696 = n984 & n2979;
  assign n5697 = n5695 & ~n5696;
  assign n5698 = pi29  & ~n5697;
  assign n5699 = pi29  & ~n5698;
  assign n5700 = ~n5697 & ~n5698;
  assign n5701 = ~n5699 & ~n5700;
  assign n5702 = n5690 & n5701;
  assign n5703 = ~n5690 & ~n5701;
  assign n5704 = ~n5702 & ~n5703;
  assign n5705 = ~n5612 & n5704;
  assign n5706 = n5612 & ~n5704;
  assign n5707 = ~n5705 & ~n5706;
  assign n5708 = pi80  & n2486;
  assign n5709 = pi78  & n2644;
  assign n5710 = pi79  & n2481;
  assign n5711 = ~n5709 & ~n5710;
  assign n5712 = ~n5708 & n5711;
  assign n5713 = n1205 & n2489;
  assign n5714 = n5712 & ~n5713;
  assign n5715 = pi26  & ~n5714;
  assign n5716 = pi26  & ~n5715;
  assign n5717 = ~n5714 & ~n5715;
  assign n5718 = ~n5716 & ~n5717;
  assign n5719 = n5707 & ~n5718;
  assign n5720 = ~n5707 & n5718;
  assign n5721 = ~n5719 & ~n5720;
  assign n5722 = n5611 & ~n5721;
  assign n5723 = ~n5611 & n5721;
  assign n5724 = ~n5722 & ~n5723;
  assign n5725 = pi83  & n2004;
  assign n5726 = pi81  & n2141;
  assign n5727 = pi82  & n1999;
  assign n5728 = ~n5726 & ~n5727;
  assign n5729 = ~n5725 & n5728;
  assign n5730 = n1672 & n2007;
  assign n5731 = n5729 & ~n5730;
  assign n5732 = pi23  & ~n5731;
  assign n5733 = pi23  & ~n5732;
  assign n5734 = ~n5731 & ~n5732;
  assign n5735 = ~n5733 & ~n5734;
  assign n5736 = n5724 & ~n5735;
  assign n5737 = n5724 & ~n5736;
  assign n5738 = ~n5735 & ~n5736;
  assign n5739 = ~n5737 & ~n5738;
  assign n5740 = ~n5443 & ~n5447;
  assign n5741 = n5739 & n5740;
  assign n5742 = ~n5739 & ~n5740;
  assign n5743 = ~n5741 & ~n5742;
  assign n5744 = pi86  & n1582;
  assign n5745 = pi84  & n1713;
  assign n5746 = pi85  & n1577;
  assign n5747 = ~n5745 & ~n5746;
  assign n5748 = ~n5744 & n5747;
  assign n5749 = n1585 & n2099;
  assign n5750 = n5748 & ~n5749;
  assign n5751 = pi20  & ~n5750;
  assign n5752 = pi20  & ~n5751;
  assign n5753 = ~n5750 & ~n5751;
  assign n5754 = ~n5752 & ~n5753;
  assign n5755 = n5743 & ~n5754;
  assign n5756 = ~n5743 & n5754;
  assign n5757 = ~n5755 & ~n5756;
  assign n5758 = n5610 & ~n5757;
  assign n5759 = ~n5610 & n5757;
  assign n5760 = ~n5758 & ~n5759;
  assign n5761 = pi89  & n1269;
  assign n5762 = pi87  & n1340;
  assign n5763 = pi88  & n1264;
  assign n5764 = ~n5762 & ~n5763;
  assign n5765 = ~n5761 & n5764;
  assign n5766 = n1272 & n2432;
  assign n5767 = n5765 & ~n5766;
  assign n5768 = pi17  & ~n5767;
  assign n5769 = pi17  & ~n5768;
  assign n5770 = ~n5767 & ~n5768;
  assign n5771 = ~n5769 & ~n5770;
  assign n5772 = n5760 & ~n5771;
  assign n5773 = ~n5760 & n5771;
  assign n5774 = ~n5772 & ~n5773;
  assign n5775 = ~n5609 & n5774;
  assign n5776 = n5609 & ~n5774;
  assign n5777 = ~n5775 & ~n5776;
  assign n5778 = ~n5608 & n5777;
  assign n5779 = n5608 & ~n5777;
  assign n5780 = ~n5778 & ~n5779;
  assign n5781 = ~n5597 & n5780;
  assign n5782 = n5597 & ~n5780;
  assign n5783 = ~n5781 & ~n5782;
  assign n5784 = n5596 & ~n5783;
  assign n5785 = ~n5596 & n5783;
  assign n5786 = ~n5784 & ~n5785;
  assign n5787 = ~n5585 & n5786;
  assign n5788 = n5585 & ~n5786;
  assign n5789 = ~n5787 & ~n5788;
  assign n5790 = n5584 & ~n5789;
  assign n5791 = ~n5584 & n5789;
  assign n5792 = ~n5790 & ~n5791;
  assign n5793 = ~n5573 & n5792;
  assign n5794 = n5573 & ~n5792;
  assign n5795 = ~n5793 & ~n5794;
  assign n5796 = pi101  & n340;
  assign n5797 = pi99  & n380;
  assign n5798 = pi100  & n335;
  assign n5799 = ~n5797 & ~n5798;
  assign n5800 = ~n5796 & n5799;
  assign n5801 = n343 & n5056;
  assign n5802 = n5800 & ~n5801;
  assign n5803 = pi5  & ~n5802;
  assign n5804 = pi5  & ~n5803;
  assign n5805 = ~n5802 & ~n5803;
  assign n5806 = ~n5804 & ~n5805;
  assign n5807 = n5795 & ~n5806;
  assign n5808 = ~n5795 & n5806;
  assign n5809 = ~n5807 & ~n5808;
  assign n5810 = ~n5572 & n5809;
  assign n5811 = n5572 & ~n5809;
  assign n5812 = ~n5810 & ~n5811;
  assign n5813 = ~n5571 & n5812;
  assign n5814 = n5571 & ~n5812;
  assign n5815 = ~n5813 & ~n5814;
  assign n5816 = ~n5553 & n5815;
  assign n5817 = n5553 & ~n5815;
  assign po40  = ~n5816 & ~n5817;
  assign n5819 = ~n5813 & ~n5816;
  assign n5820 = ~n5807 & ~n5810;
  assign n5821 = pi102  & n340;
  assign n5822 = pi100  & n380;
  assign n5823 = pi101  & n335;
  assign n5824 = ~n5822 & ~n5823;
  assign n5825 = ~n5821 & n5824;
  assign n5826 = n343 & n5296;
  assign n5827 = n5825 & ~n5826;
  assign n5828 = pi5  & ~n5827;
  assign n5829 = pi5  & ~n5828;
  assign n5830 = ~n5827 & ~n5828;
  assign n5831 = ~n5829 & ~n5830;
  assign n5832 = ~n5791 & ~n5793;
  assign n5833 = ~n5785 & ~n5787;
  assign n5834 = pi96  & n675;
  assign n5835 = pi94  & n769;
  assign n5836 = pi95  & n670;
  assign n5837 = ~n5835 & ~n5836;
  assign n5838 = ~n5834 & n5837;
  assign n5839 = n678 & n3921;
  assign n5840 = n5838 & ~n5839;
  assign n5841 = pi11  & ~n5840;
  assign n5842 = pi11  & ~n5841;
  assign n5843 = ~n5840 & ~n5841;
  assign n5844 = ~n5842 & ~n5843;
  assign n5845 = ~n5778 & ~n5781;
  assign n5846 = pi93  & n918;
  assign n5847 = pi91  & n1031;
  assign n5848 = pi92  & n913;
  assign n5849 = ~n5847 & ~n5848;
  assign n5850 = ~n5846 & n5849;
  assign n5851 = n921 & n3144;
  assign n5852 = n5850 & ~n5851;
  assign n5853 = pi14  & ~n5852;
  assign n5854 = pi14  & ~n5853;
  assign n5855 = ~n5852 & ~n5853;
  assign n5856 = ~n5854 & ~n5855;
  assign n5857 = ~n5772 & ~n5775;
  assign n5858 = ~n5755 & ~n5759;
  assign n5859 = ~n5719 & ~n5723;
  assign n5860 = pi81  & n2486;
  assign n5861 = pi79  & n2644;
  assign n5862 = pi80  & n2481;
  assign n5863 = ~n5861 & ~n5862;
  assign n5864 = ~n5860 & n5863;
  assign n5865 = n1413 & n2489;
  assign n5866 = n5864 & ~n5865;
  assign n5867 = pi26  & ~n5866;
  assign n5868 = pi26  & ~n5867;
  assign n5869 = ~n5866 & ~n5867;
  assign n5870 = ~n5868 & ~n5869;
  assign n5871 = ~n5703 & ~n5705;
  assign n5872 = pi78  & n2976;
  assign n5873 = pi76  & n3182;
  assign n5874 = pi77  & n2971;
  assign n5875 = ~n5873 & ~n5874;
  assign n5876 = ~n5872 & n5875;
  assign n5877 = n1009 & n2979;
  assign n5878 = n5876 & ~n5877;
  assign n5879 = pi29  & ~n5878;
  assign n5880 = pi29  & ~n5879;
  assign n5881 = ~n5878 & ~n5879;
  assign n5882 = ~n5880 & ~n5881;
  assign n5883 = pi75  & n3550;
  assign n5884 = pi73  & n3735;
  assign n5885 = pi74  & n3545;
  assign n5886 = ~n5884 & ~n5885;
  assign n5887 = ~n5883 & n5886;
  assign n5888 = n747 & n3553;
  assign n5889 = n5887 & ~n5888;
  assign n5890 = pi32  & ~n5889;
  assign n5891 = pi32  & ~n5890;
  assign n5892 = ~n5889 & ~n5890;
  assign n5893 = ~n5891 & ~n5892;
  assign n5894 = ~n5666 & ~n5670;
  assign n5895 = pi72  & n4182;
  assign n5896 = pi70  & n4416;
  assign n5897 = pi71  & n4177;
  assign n5898 = ~n5896 & ~n5897;
  assign n5899 = ~n5895 & n5898;
  assign n5900 = n575 & n4185;
  assign n5901 = n5899 & ~n5900;
  assign n5902 = pi35  & ~n5901;
  assign n5903 = pi35  & ~n5902;
  assign n5904 = ~n5901 & ~n5902;
  assign n5905 = ~n5903 & ~n5904;
  assign n5906 = ~n5650 & ~n5652;
  assign n5907 = pi66  & n5636;
  assign n5908 = n5365 & ~n5635;
  assign n5909 = n5630 & n5908;
  assign n5910 = pi64  & n5909;
  assign n5911 = pi65  & n5631;
  assign n5912 = ~n5910 & ~n5911;
  assign n5913 = ~n5907 & n5912;
  assign n5914 = n291 & n5639;
  assign n5915 = n5913 & ~n5914;
  assign n5916 = pi41  & ~n5915;
  assign n5917 = pi41  & ~n5916;
  assign n5918 = ~n5915 & ~n5916;
  assign n5919 = ~n5917 & ~n5918;
  assign n5920 = ~n5646 & n5919;
  assign n5921 = n5646 & ~n5919;
  assign n5922 = ~n5920 & ~n5921;
  assign n5923 = pi69  & n4896;
  assign n5924 = pi67  & n5148;
  assign n5925 = pi68  & n4891;
  assign n5926 = ~n5924 & ~n5925;
  assign n5927 = ~n5923 & n5926;
  assign n5928 = n405 & n4899;
  assign n5929 = n5927 & ~n5928;
  assign n5930 = pi38  & ~n5929;
  assign n5931 = pi38  & ~n5930;
  assign n5932 = ~n5929 & ~n5930;
  assign n5933 = ~n5931 & ~n5932;
  assign n5934 = n5922 & ~n5933;
  assign n5935 = ~n5922 & n5933;
  assign n5936 = ~n5934 & ~n5935;
  assign n5937 = ~n5906 & n5936;
  assign n5938 = n5906 & ~n5936;
  assign n5939 = ~n5937 & ~n5938;
  assign n5940 = ~n5905 & n5939;
  assign n5941 = n5905 & ~n5939;
  assign n5942 = ~n5940 & ~n5941;
  assign n5943 = ~n5894 & n5942;
  assign n5944 = n5894 & ~n5942;
  assign n5945 = ~n5943 & ~n5944;
  assign n5946 = n5893 & ~n5945;
  assign n5947 = ~n5893 & n5945;
  assign n5948 = ~n5946 & ~n5947;
  assign n5949 = ~n5688 & n5948;
  assign n5950 = n5688 & ~n5948;
  assign n5951 = ~n5949 & ~n5950;
  assign n5952 = n5882 & ~n5951;
  assign n5953 = ~n5882 & n5951;
  assign n5954 = ~n5952 & ~n5953;
  assign n5955 = ~n5871 & n5954;
  assign n5956 = n5871 & ~n5954;
  assign n5957 = ~n5955 & ~n5956;
  assign n5958 = n5870 & ~n5957;
  assign n5959 = ~n5870 & n5957;
  assign n5960 = ~n5958 & ~n5959;
  assign n5961 = ~n5859 & n5960;
  assign n5962 = n5859 & ~n5960;
  assign n5963 = ~n5961 & ~n5962;
  assign n5964 = pi84  & n2004;
  assign n5965 = pi82  & n2141;
  assign n5966 = pi83  & n1999;
  assign n5967 = ~n5965 & ~n5966;
  assign n5968 = ~n5964 & n5967;
  assign n5969 = n1805 & n2007;
  assign n5970 = n5968 & ~n5969;
  assign n5971 = pi23  & ~n5970;
  assign n5972 = pi23  & ~n5971;
  assign n5973 = ~n5970 & ~n5971;
  assign n5974 = ~n5972 & ~n5973;
  assign n5975 = n5963 & ~n5974;
  assign n5976 = n5963 & ~n5975;
  assign n5977 = ~n5974 & ~n5975;
  assign n5978 = ~n5976 & ~n5977;
  assign n5979 = ~n5736 & ~n5742;
  assign n5980 = n5978 & n5979;
  assign n5981 = ~n5978 & ~n5979;
  assign n5982 = ~n5980 & ~n5981;
  assign n5983 = pi87  & n1582;
  assign n5984 = pi85  & n1713;
  assign n5985 = pi86  & n1577;
  assign n5986 = ~n5984 & ~n5985;
  assign n5987 = ~n5983 & n5986;
  assign n5988 = n1585 & n2252;
  assign n5989 = n5987 & ~n5988;
  assign n5990 = pi20  & ~n5989;
  assign n5991 = pi20  & ~n5990;
  assign n5992 = ~n5989 & ~n5990;
  assign n5993 = ~n5991 & ~n5992;
  assign n5994 = n5982 & ~n5993;
  assign n5995 = ~n5982 & n5993;
  assign n5996 = ~n5858 & ~n5995;
  assign n5997 = ~n5994 & n5996;
  assign n5998 = ~n5858 & ~n5997;
  assign n5999 = ~n5994 & ~n5997;
  assign n6000 = ~n5995 & n5999;
  assign n6001 = ~n5998 & ~n6000;
  assign n6002 = pi90  & n1269;
  assign n6003 = pi88  & n1340;
  assign n6004 = pi89  & n1264;
  assign n6005 = ~n6003 & ~n6004;
  assign n6006 = ~n6002 & n6005;
  assign n6007 = n1272 & n2606;
  assign n6008 = n6006 & ~n6007;
  assign n6009 = pi17  & ~n6008;
  assign n6010 = pi17  & ~n6009;
  assign n6011 = ~n6008 & ~n6009;
  assign n6012 = ~n6010 & ~n6011;
  assign n6013 = n6001 & n6012;
  assign n6014 = ~n6001 & ~n6012;
  assign n6015 = ~n6013 & ~n6014;
  assign n6016 = ~n5857 & n6015;
  assign n6017 = n5857 & ~n6015;
  assign n6018 = ~n6016 & ~n6017;
  assign n6019 = n5856 & ~n6018;
  assign n6020 = ~n5856 & n6018;
  assign n6021 = ~n6019 & ~n6020;
  assign n6022 = ~n5845 & n6021;
  assign n6023 = n5845 & ~n6021;
  assign n6024 = ~n6022 & ~n6023;
  assign n6025 = n5844 & ~n6024;
  assign n6026 = ~n5844 & n6024;
  assign n6027 = ~n6025 & ~n6026;
  assign n6028 = ~n5833 & n6027;
  assign n6029 = n5833 & ~n6027;
  assign n6030 = ~n6028 & ~n6029;
  assign n6031 = pi99  & n493;
  assign n6032 = pi97  & n533;
  assign n6033 = pi98  & n488;
  assign n6034 = ~n6032 & ~n6033;
  assign n6035 = ~n6031 & n6034;
  assign n6036 = n496 & n4584;
  assign n6037 = n6035 & ~n6036;
  assign n6038 = pi8  & ~n6037;
  assign n6039 = pi8  & ~n6038;
  assign n6040 = ~n6037 & ~n6038;
  assign n6041 = ~n6039 & ~n6040;
  assign n6042 = n6030 & ~n6041;
  assign n6043 = ~n6030 & n6041;
  assign n6044 = ~n6042 & ~n6043;
  assign n6045 = ~n5832 & n6044;
  assign n6046 = n5832 & ~n6044;
  assign n6047 = ~n6045 & ~n6046;
  assign n6048 = ~n5831 & n6047;
  assign n6049 = n5831 & ~n6047;
  assign n6050 = ~n6048 & ~n6049;
  assign n6051 = n5820 & ~n6050;
  assign n6052 = ~n5820 & n6050;
  assign n6053 = ~n6051 & ~n6052;
  assign n6054 = pi105  & n264;
  assign n6055 = pi103  & n281;
  assign n6056 = pi104  & n259;
  assign n6057 = ~n6055 & ~n6056;
  assign n6058 = ~n6054 & n6057;
  assign n6059 = ~n5561 & ~n5563;
  assign n6060 = ~pi104  & ~pi105 ;
  assign n6061 = pi104  & pi105 ;
  assign n6062 = ~n6060 & ~n6061;
  assign n6063 = ~n6059 & n6062;
  assign n6064 = n6059 & ~n6062;
  assign n6065 = ~n6063 & ~n6064;
  assign n6066 = n267 & n6065;
  assign n6067 = n6058 & ~n6066;
  assign n6068 = pi2  & ~n6067;
  assign n6069 = pi2  & ~n6068;
  assign n6070 = ~n6067 & ~n6068;
  assign n6071 = ~n6069 & ~n6070;
  assign n6072 = ~n6053 & n6071;
  assign n6073 = n6053 & ~n6071;
  assign n6074 = ~n6072 & ~n6073;
  assign n6075 = ~n5819 & n6074;
  assign n6076 = n5819 & ~n6074;
  assign po41  = ~n6075 & ~n6076;
  assign n6078 = ~n6073 & ~n6075;
  assign n6079 = pi106  & n264;
  assign n6080 = pi104  & n281;
  assign n6081 = pi105  & n259;
  assign n6082 = ~n6080 & ~n6081;
  assign n6083 = ~n6079 & n6082;
  assign n6084 = ~n6061 & ~n6063;
  assign n6085 = ~pi105  & ~pi106 ;
  assign n6086 = pi105  & pi106 ;
  assign n6087 = ~n6085 & ~n6086;
  assign n6088 = ~n6084 & n6087;
  assign n6089 = n6084 & ~n6087;
  assign n6090 = ~n6088 & ~n6089;
  assign n6091 = n267 & n6090;
  assign n6092 = n6083 & ~n6091;
  assign n6093 = pi2  & ~n6092;
  assign n6094 = pi2  & ~n6093;
  assign n6095 = ~n6092 & ~n6093;
  assign n6096 = ~n6094 & ~n6095;
  assign n6097 = ~n6048 & ~n6052;
  assign n6098 = pi103  & n340;
  assign n6099 = pi101  & n380;
  assign n6100 = pi102  & n335;
  assign n6101 = ~n6099 & ~n6100;
  assign n6102 = ~n6098 & n6101;
  assign n6103 = n343 & n5540;
  assign n6104 = n6102 & ~n6103;
  assign n6105 = pi5  & ~n6104;
  assign n6106 = pi5  & ~n6105;
  assign n6107 = ~n6104 & ~n6105;
  assign n6108 = ~n6106 & ~n6107;
  assign n6109 = ~n6042 & ~n6045;
  assign n6110 = pi100  & n493;
  assign n6111 = pi98  & n533;
  assign n6112 = pi99  & n488;
  assign n6113 = ~n6111 & ~n6112;
  assign n6114 = ~n6110 & n6113;
  assign n6115 = n496 & n4808;
  assign n6116 = n6114 & ~n6115;
  assign n6117 = pi8  & ~n6116;
  assign n6118 = pi8  & ~n6117;
  assign n6119 = ~n6116 & ~n6117;
  assign n6120 = ~n6118 & ~n6119;
  assign n6121 = ~n6026 & ~n6028;
  assign n6122 = ~n6020 & ~n6022;
  assign n6123 = pi94  & n918;
  assign n6124 = pi92  & n1031;
  assign n6125 = pi93  & n913;
  assign n6126 = ~n6124 & ~n6125;
  assign n6127 = ~n6123 & n6126;
  assign n6128 = n921 & n3499;
  assign n6129 = n6127 & ~n6128;
  assign n6130 = pi14  & ~n6129;
  assign n6131 = pi14  & ~n6130;
  assign n6132 = ~n6129 & ~n6130;
  assign n6133 = ~n6131 & ~n6132;
  assign n6134 = ~n6014 & ~n6016;
  assign n6135 = ~n5959 & ~n5961;
  assign n6136 = pi82  & n2486;
  assign n6137 = pi80  & n2644;
  assign n6138 = pi81  & n2481;
  assign n6139 = ~n6137 & ~n6138;
  assign n6140 = ~n6136 & n6139;
  assign n6141 = n1532 & n2489;
  assign n6142 = n6140 & ~n6141;
  assign n6143 = pi26  & ~n6142;
  assign n6144 = pi26  & ~n6143;
  assign n6145 = ~n6142 & ~n6143;
  assign n6146 = ~n6144 & ~n6145;
  assign n6147 = ~n5953 & ~n5955;
  assign n6148 = ~n5947 & ~n5949;
  assign n6149 = pi76  & n3550;
  assign n6150 = pi74  & n3735;
  assign n6151 = pi75  & n3545;
  assign n6152 = ~n6150 & ~n6151;
  assign n6153 = ~n6149 & n6152;
  assign n6154 = n881 & n3553;
  assign n6155 = n6153 & ~n6154;
  assign n6156 = pi32  & ~n6155;
  assign n6157 = pi32  & ~n6156;
  assign n6158 = ~n6155 & ~n6156;
  assign n6159 = ~n6157 & ~n6158;
  assign n6160 = ~n5940 & ~n5943;
  assign n6161 = ~n5934 & ~n5937;
  assign n6162 = pi67  & n5636;
  assign n6163 = pi65  & n5909;
  assign n6164 = pi66  & n5631;
  assign n6165 = ~n6163 & ~n6164;
  assign n6166 = ~n6162 & n6165;
  assign n6167 = n313 & n5639;
  assign n6168 = n6166 & ~n6167;
  assign n6169 = pi41  & ~n6168;
  assign n6170 = pi41  & ~n6169;
  assign n6171 = ~n6168 & ~n6169;
  assign n6172 = ~n6170 & ~n6171;
  assign n6173 = pi41  & ~pi42 ;
  assign n6174 = ~pi41  & pi42 ;
  assign n6175 = ~n6173 & ~n6174;
  assign n6176 = pi64  & ~n6175;
  assign n6177 = n5921 & n6176;
  assign n6178 = ~n5921 & ~n6176;
  assign n6179 = ~n6177 & ~n6178;
  assign n6180 = ~n6172 & n6179;
  assign n6181 = n6172 & ~n6179;
  assign n6182 = ~n6180 & ~n6181;
  assign n6183 = pi70  & n4896;
  assign n6184 = pi68  & n5148;
  assign n6185 = pi69  & n4891;
  assign n6186 = ~n6184 & ~n6185;
  assign n6187 = ~n6183 & n6186;
  assign n6188 = n430 & n4899;
  assign n6189 = n6187 & ~n6188;
  assign n6190 = pi38  & ~n6189;
  assign n6191 = pi38  & ~n6190;
  assign n6192 = ~n6189 & ~n6190;
  assign n6193 = ~n6191 & ~n6192;
  assign n6194 = n6182 & ~n6193;
  assign n6195 = ~n6182 & n6193;
  assign n6196 = ~n6194 & ~n6195;
  assign n6197 = n6161 & ~n6196;
  assign n6198 = ~n6161 & n6196;
  assign n6199 = ~n6197 & ~n6198;
  assign n6200 = pi73  & n4182;
  assign n6201 = pi71  & n4416;
  assign n6202 = pi72  & n4177;
  assign n6203 = ~n6201 & ~n6202;
  assign n6204 = ~n6200 & n6203;
  assign n6205 = n639 & n4185;
  assign n6206 = n6204 & ~n6205;
  assign n6207 = pi35  & ~n6206;
  assign n6208 = pi35  & ~n6207;
  assign n6209 = ~n6206 & ~n6207;
  assign n6210 = ~n6208 & ~n6209;
  assign n6211 = ~n6199 & n6210;
  assign n6212 = n6199 & ~n6210;
  assign n6213 = ~n6211 & ~n6212;
  assign n6214 = ~n6160 & n6213;
  assign n6215 = n6160 & ~n6213;
  assign n6216 = ~n6214 & ~n6215;
  assign n6217 = ~n6159 & n6216;
  assign n6218 = n6159 & ~n6216;
  assign n6219 = ~n6217 & ~n6218;
  assign n6220 = ~n6148 & n6219;
  assign n6221 = n6148 & ~n6219;
  assign n6222 = ~n6220 & ~n6221;
  assign n6223 = pi79  & n2976;
  assign n6224 = pi77  & n3182;
  assign n6225 = pi78  & n2971;
  assign n6226 = ~n6224 & ~n6225;
  assign n6227 = ~n6223 & n6226;
  assign n6228 = n1105 & n2979;
  assign n6229 = n6227 & ~n6228;
  assign n6230 = pi29  & ~n6229;
  assign n6231 = pi29  & ~n6230;
  assign n6232 = ~n6229 & ~n6230;
  assign n6233 = ~n6231 & ~n6232;
  assign n6234 = n6222 & ~n6233;
  assign n6235 = n6222 & ~n6234;
  assign n6236 = ~n6233 & ~n6234;
  assign n6237 = ~n6235 & ~n6236;
  assign n6238 = ~n6147 & ~n6237;
  assign n6239 = n6147 & n6237;
  assign n6240 = ~n6238 & ~n6239;
  assign n6241 = ~n6146 & n6240;
  assign n6242 = n6146 & ~n6240;
  assign n6243 = ~n6241 & ~n6242;
  assign n6244 = ~n6135 & n6243;
  assign n6245 = n6135 & ~n6243;
  assign n6246 = ~n6244 & ~n6245;
  assign n6247 = pi85  & n2004;
  assign n6248 = pi83  & n2141;
  assign n6249 = pi84  & n1999;
  assign n6250 = ~n6248 & ~n6249;
  assign n6251 = ~n6247 & n6250;
  assign n6252 = n1943 & n2007;
  assign n6253 = n6251 & ~n6252;
  assign n6254 = pi23  & ~n6253;
  assign n6255 = pi23  & ~n6254;
  assign n6256 = ~n6253 & ~n6254;
  assign n6257 = ~n6255 & ~n6256;
  assign n6258 = n6246 & ~n6257;
  assign n6259 = n6246 & ~n6258;
  assign n6260 = ~n6257 & ~n6258;
  assign n6261 = ~n6259 & ~n6260;
  assign n6262 = ~n5975 & ~n5981;
  assign n6263 = n6261 & n6262;
  assign n6264 = ~n6261 & ~n6262;
  assign n6265 = ~n6263 & ~n6264;
  assign n6266 = pi88  & n1582;
  assign n6267 = pi86  & n1713;
  assign n6268 = pi87  & n1577;
  assign n6269 = ~n6267 & ~n6268;
  assign n6270 = ~n6266 & n6269;
  assign n6271 = n1585 & n2277;
  assign n6272 = n6270 & ~n6271;
  assign n6273 = pi20  & ~n6272;
  assign n6274 = pi20  & ~n6273;
  assign n6275 = ~n6272 & ~n6273;
  assign n6276 = ~n6274 & ~n6275;
  assign n6277 = ~n6265 & n6276;
  assign n6278 = n6265 & ~n6276;
  assign n6279 = ~n6277 & ~n6278;
  assign n6280 = ~n5999 & n6279;
  assign n6281 = n5999 & ~n6279;
  assign n6282 = ~n6280 & ~n6281;
  assign n6283 = pi91  & n1269;
  assign n6284 = pi89  & n1340;
  assign n6285 = pi90  & n1264;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = ~n6283 & n6286;
  assign n6288 = n1272 & n2926;
  assign n6289 = n6287 & ~n6288;
  assign n6290 = pi17  & ~n6289;
  assign n6291 = pi17  & ~n6290;
  assign n6292 = ~n6289 & ~n6290;
  assign n6293 = ~n6291 & ~n6292;
  assign n6294 = n6282 & ~n6293;
  assign n6295 = ~n6282 & n6293;
  assign n6296 = ~n6294 & ~n6295;
  assign n6297 = ~n6134 & n6296;
  assign n6298 = n6134 & ~n6296;
  assign n6299 = ~n6297 & ~n6298;
  assign n6300 = ~n6133 & n6299;
  assign n6301 = n6133 & ~n6299;
  assign n6302 = ~n6300 & ~n6301;
  assign n6303 = ~n6122 & n6302;
  assign n6304 = n6122 & ~n6302;
  assign n6305 = ~n6303 & ~n6304;
  assign n6306 = pi97  & n675;
  assign n6307 = pi95  & n769;
  assign n6308 = pi96  & n670;
  assign n6309 = ~n6307 & ~n6308;
  assign n6310 = ~n6306 & n6309;
  assign n6311 = n678 & n3946;
  assign n6312 = n6310 & ~n6311;
  assign n6313 = pi11  & ~n6312;
  assign n6314 = pi11  & ~n6313;
  assign n6315 = ~n6312 & ~n6313;
  assign n6316 = ~n6314 & ~n6315;
  assign n6317 = n6305 & ~n6316;
  assign n6318 = ~n6305 & n6316;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = ~n6121 & n6319;
  assign n6321 = n6121 & ~n6319;
  assign n6322 = ~n6320 & ~n6321;
  assign n6323 = n6120 & ~n6322;
  assign n6324 = ~n6120 & n6322;
  assign n6325 = ~n6323 & ~n6324;
  assign n6326 = ~n6109 & n6325;
  assign n6327 = n6109 & ~n6325;
  assign n6328 = ~n6326 & ~n6327;
  assign n6329 = ~n6108 & n6328;
  assign n6330 = n6108 & ~n6328;
  assign n6331 = ~n6329 & ~n6330;
  assign n6332 = ~n6097 & n6331;
  assign n6333 = n6097 & ~n6331;
  assign n6334 = ~n6332 & ~n6333;
  assign n6335 = ~n6096 & n6334;
  assign n6336 = n6096 & ~n6334;
  assign n6337 = ~n6335 & ~n6336;
  assign n6338 = ~n6078 & n6337;
  assign n6339 = n6078 & ~n6337;
  assign po42  = ~n6338 & ~n6339;
  assign n6341 = ~n6335 & ~n6338;
  assign n6342 = ~n6329 & ~n6332;
  assign n6343 = ~n6324 & ~n6326;
  assign n6344 = ~n6317 & ~n6320;
  assign n6345 = ~n6300 & ~n6303;
  assign n6346 = pi95  & n918;
  assign n6347 = pi93  & n1031;
  assign n6348 = pi94  & n913;
  assign n6349 = ~n6347 & ~n6348;
  assign n6350 = ~n6346 & n6349;
  assign n6351 = n921 & n3710;
  assign n6352 = n6350 & ~n6351;
  assign n6353 = pi14  & ~n6352;
  assign n6354 = pi14  & ~n6353;
  assign n6355 = ~n6352 & ~n6353;
  assign n6356 = ~n6354 & ~n6355;
  assign n6357 = ~n6294 & ~n6297;
  assign n6358 = pi92  & n1269;
  assign n6359 = pi90  & n1340;
  assign n6360 = pi91  & n1264;
  assign n6361 = ~n6359 & ~n6360;
  assign n6362 = ~n6358 & n6361;
  assign n6363 = n1272 & n3119;
  assign n6364 = n6362 & ~n6363;
  assign n6365 = pi17  & ~n6364;
  assign n6366 = pi17  & ~n6365;
  assign n6367 = ~n6364 & ~n6365;
  assign n6368 = ~n6366 & ~n6367;
  assign n6369 = ~n6278 & ~n6280;
  assign n6370 = ~n6258 & ~n6264;
  assign n6371 = ~n6234 & ~n6238;
  assign n6372 = ~n6217 & ~n6220;
  assign n6373 = ~n6212 & ~n6214;
  assign n6374 = ~n6194 & ~n6198;
  assign n6375 = ~n6177 & ~n6180;
  assign n6376 = pi68  & n5636;
  assign n6377 = pi66  & n5909;
  assign n6378 = pi67  & n5631;
  assign n6379 = ~n6377 & ~n6378;
  assign n6380 = ~n6376 & n6379;
  assign n6381 = n364 & n5639;
  assign n6382 = n6380 & ~n6381;
  assign n6383 = pi41  & ~n6382;
  assign n6384 = pi41  & ~n6383;
  assign n6385 = ~n6382 & ~n6383;
  assign n6386 = ~n6384 & ~n6385;
  assign n6387 = pi44  & ~n6176;
  assign n6388 = ~pi42  & pi43 ;
  assign n6389 = pi42  & ~pi43 ;
  assign n6390 = ~n6388 & ~n6389;
  assign n6391 = n6175 & ~n6390;
  assign n6392 = pi64  & n6391;
  assign n6393 = ~pi43  & pi44 ;
  assign n6394 = pi43  & ~pi44 ;
  assign n6395 = ~n6393 & ~n6394;
  assign n6396 = ~n6175 & n6395;
  assign n6397 = pi65  & n6396;
  assign n6398 = ~n6392 & ~n6397;
  assign n6399 = ~n6175 & ~n6395;
  assign n6400 = n270 & n6399;
  assign n6401 = n6398 & ~n6400;
  assign n6402 = pi44  & ~n6401;
  assign n6403 = pi44  & ~n6402;
  assign n6404 = ~n6401 & ~n6402;
  assign n6405 = ~n6403 & ~n6404;
  assign n6406 = n6387 & ~n6405;
  assign n6407 = ~n6387 & n6405;
  assign n6408 = ~n6406 & ~n6407;
  assign n6409 = n6386 & ~n6408;
  assign n6410 = ~n6386 & n6408;
  assign n6411 = ~n6409 & ~n6410;
  assign n6412 = ~n6375 & n6411;
  assign n6413 = n6375 & ~n6411;
  assign n6414 = ~n6412 & ~n6413;
  assign n6415 = pi71  & n4896;
  assign n6416 = pi69  & n5148;
  assign n6417 = pi70  & n4891;
  assign n6418 = ~n6416 & ~n6417;
  assign n6419 = ~n6415 & n6418;
  assign n6420 = n476 & n4899;
  assign n6421 = n6419 & ~n6420;
  assign n6422 = pi38  & ~n6421;
  assign n6423 = pi38  & ~n6422;
  assign n6424 = ~n6421 & ~n6422;
  assign n6425 = ~n6423 & ~n6424;
  assign n6426 = n6414 & ~n6425;
  assign n6427 = ~n6414 & n6425;
  assign n6428 = ~n6426 & ~n6427;
  assign n6429 = n6374 & ~n6428;
  assign n6430 = ~n6374 & n6428;
  assign n6431 = ~n6429 & ~n6430;
  assign n6432 = pi74  & n4182;
  assign n6433 = pi72  & n4416;
  assign n6434 = pi73  & n4177;
  assign n6435 = ~n6433 & ~n6434;
  assign n6436 = ~n6432 & n6435;
  assign n6437 = n722 & n4185;
  assign n6438 = n6436 & ~n6437;
  assign n6439 = pi35  & ~n6438;
  assign n6440 = pi35  & ~n6439;
  assign n6441 = ~n6438 & ~n6439;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = n6431 & ~n6442;
  assign n6444 = ~n6431 & n6442;
  assign n6445 = ~n6373 & ~n6444;
  assign n6446 = ~n6443 & n6445;
  assign n6447 = ~n6373 & ~n6446;
  assign n6448 = ~n6443 & ~n6446;
  assign n6449 = ~n6444 & n6448;
  assign n6450 = ~n6447 & ~n6449;
  assign n6451 = pi77  & n3550;
  assign n6452 = pi75  & n3735;
  assign n6453 = pi76  & n3545;
  assign n6454 = ~n6452 & ~n6453;
  assign n6455 = ~n6451 & n6454;
  assign n6456 = n984 & n3553;
  assign n6457 = n6455 & ~n6456;
  assign n6458 = pi32  & ~n6457;
  assign n6459 = pi32  & ~n6458;
  assign n6460 = ~n6457 & ~n6458;
  assign n6461 = ~n6459 & ~n6460;
  assign n6462 = n6450 & n6461;
  assign n6463 = ~n6450 & ~n6461;
  assign n6464 = ~n6462 & ~n6463;
  assign n6465 = ~n6372 & n6464;
  assign n6466 = n6372 & ~n6464;
  assign n6467 = ~n6465 & ~n6466;
  assign n6468 = pi80  & n2976;
  assign n6469 = pi78  & n3182;
  assign n6470 = pi79  & n2971;
  assign n6471 = ~n6469 & ~n6470;
  assign n6472 = ~n6468 & n6471;
  assign n6473 = n1205 & n2979;
  assign n6474 = n6472 & ~n6473;
  assign n6475 = pi29  & ~n6474;
  assign n6476 = pi29  & ~n6475;
  assign n6477 = ~n6474 & ~n6475;
  assign n6478 = ~n6476 & ~n6477;
  assign n6479 = n6467 & ~n6478;
  assign n6480 = ~n6467 & n6478;
  assign n6481 = ~n6479 & ~n6480;
  assign n6482 = n6371 & ~n6481;
  assign n6483 = ~n6371 & n6481;
  assign n6484 = ~n6482 & ~n6483;
  assign n6485 = pi83  & n2486;
  assign n6486 = pi81  & n2644;
  assign n6487 = pi82  & n2481;
  assign n6488 = ~n6486 & ~n6487;
  assign n6489 = ~n6485 & n6488;
  assign n6490 = n1672 & n2489;
  assign n6491 = n6489 & ~n6490;
  assign n6492 = pi26  & ~n6491;
  assign n6493 = pi26  & ~n6492;
  assign n6494 = ~n6491 & ~n6492;
  assign n6495 = ~n6493 & ~n6494;
  assign n6496 = n6484 & ~n6495;
  assign n6497 = n6484 & ~n6496;
  assign n6498 = ~n6495 & ~n6496;
  assign n6499 = ~n6497 & ~n6498;
  assign n6500 = ~n6241 & ~n6244;
  assign n6501 = n6499 & n6500;
  assign n6502 = ~n6499 & ~n6500;
  assign n6503 = ~n6501 & ~n6502;
  assign n6504 = pi86  & n2004;
  assign n6505 = pi84  & n2141;
  assign n6506 = pi85  & n1999;
  assign n6507 = ~n6505 & ~n6506;
  assign n6508 = ~n6504 & n6507;
  assign n6509 = n2007 & n2099;
  assign n6510 = n6508 & ~n6509;
  assign n6511 = pi23  & ~n6510;
  assign n6512 = pi23  & ~n6511;
  assign n6513 = ~n6510 & ~n6511;
  assign n6514 = ~n6512 & ~n6513;
  assign n6515 = n6503 & ~n6514;
  assign n6516 = ~n6503 & n6514;
  assign n6517 = ~n6515 & ~n6516;
  assign n6518 = n6370 & ~n6517;
  assign n6519 = ~n6370 & n6517;
  assign n6520 = ~n6518 & ~n6519;
  assign n6521 = pi89  & n1582;
  assign n6522 = pi87  & n1713;
  assign n6523 = pi88  & n1577;
  assign n6524 = ~n6522 & ~n6523;
  assign n6525 = ~n6521 & n6524;
  assign n6526 = n1585 & n2432;
  assign n6527 = n6525 & ~n6526;
  assign n6528 = pi20  & ~n6527;
  assign n6529 = pi20  & ~n6528;
  assign n6530 = ~n6527 & ~n6528;
  assign n6531 = ~n6529 & ~n6530;
  assign n6532 = n6520 & ~n6531;
  assign n6533 = ~n6520 & n6531;
  assign n6534 = ~n6532 & ~n6533;
  assign n6535 = ~n6369 & n6534;
  assign n6536 = n6369 & ~n6534;
  assign n6537 = ~n6535 & ~n6536;
  assign n6538 = ~n6368 & n6537;
  assign n6539 = n6368 & ~n6537;
  assign n6540 = ~n6538 & ~n6539;
  assign n6541 = ~n6357 & n6540;
  assign n6542 = n6357 & ~n6540;
  assign n6543 = ~n6541 & ~n6542;
  assign n6544 = n6356 & ~n6543;
  assign n6545 = ~n6356 & n6543;
  assign n6546 = ~n6544 & ~n6545;
  assign n6547 = ~n6345 & n6546;
  assign n6548 = n6345 & ~n6546;
  assign n6549 = ~n6547 & ~n6548;
  assign n6550 = pi98  & n675;
  assign n6551 = pi96  & n769;
  assign n6552 = pi97  & n670;
  assign n6553 = ~n6551 & ~n6552;
  assign n6554 = ~n6550 & n6553;
  assign n6555 = n678 & n4360;
  assign n6556 = n6554 & ~n6555;
  assign n6557 = pi11  & ~n6556;
  assign n6558 = pi11  & ~n6557;
  assign n6559 = ~n6556 & ~n6557;
  assign n6560 = ~n6558 & ~n6559;
  assign n6561 = n6549 & ~n6560;
  assign n6562 = ~n6549 & n6560;
  assign n6563 = ~n6561 & ~n6562;
  assign n6564 = n6344 & ~n6563;
  assign n6565 = ~n6344 & n6563;
  assign n6566 = ~n6564 & ~n6565;
  assign n6567 = pi101  & n493;
  assign n6568 = pi99  & n533;
  assign n6569 = pi100  & n488;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = ~n6567 & n6570;
  assign n6572 = n496 & n5056;
  assign n6573 = n6571 & ~n6572;
  assign n6574 = pi8  & ~n6573;
  assign n6575 = pi8  & ~n6574;
  assign n6576 = ~n6573 & ~n6574;
  assign n6577 = ~n6575 & ~n6576;
  assign n6578 = n6566 & ~n6577;
  assign n6579 = ~n6566 & n6577;
  assign n6580 = ~n6343 & ~n6579;
  assign n6581 = ~n6578 & n6580;
  assign n6582 = ~n6343 & ~n6581;
  assign n6583 = ~n6578 & ~n6581;
  assign n6584 = ~n6579 & n6583;
  assign n6585 = ~n6582 & ~n6584;
  assign n6586 = pi104  & n340;
  assign n6587 = pi102  & n380;
  assign n6588 = pi103  & n335;
  assign n6589 = ~n6587 & ~n6588;
  assign n6590 = ~n6586 & n6589;
  assign n6591 = n343 & n5565;
  assign n6592 = n6590 & ~n6591;
  assign n6593 = pi5  & ~n6592;
  assign n6594 = pi5  & ~n6593;
  assign n6595 = ~n6592 & ~n6593;
  assign n6596 = ~n6594 & ~n6595;
  assign n6597 = n6585 & n6596;
  assign n6598 = ~n6585 & ~n6596;
  assign n6599 = ~n6597 & ~n6598;
  assign n6600 = ~n6342 & n6599;
  assign n6601 = n6342 & ~n6599;
  assign n6602 = ~n6600 & ~n6601;
  assign n6603 = pi107  & n264;
  assign n6604 = pi105  & n281;
  assign n6605 = pi106  & n259;
  assign n6606 = ~n6604 & ~n6605;
  assign n6607 = ~n6603 & n6606;
  assign n6608 = ~n6086 & ~n6088;
  assign n6609 = ~pi106  & ~pi107 ;
  assign n6610 = pi106  & pi107 ;
  assign n6611 = ~n6609 & ~n6610;
  assign n6612 = ~n6608 & n6611;
  assign n6613 = n6608 & ~n6611;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = n267 & n6614;
  assign n6616 = n6607 & ~n6615;
  assign n6617 = pi2  & ~n6616;
  assign n6618 = pi2  & ~n6617;
  assign n6619 = ~n6616 & ~n6617;
  assign n6620 = ~n6618 & ~n6619;
  assign n6621 = n6602 & ~n6620;
  assign n6622 = ~n6602 & n6620;
  assign n6623 = ~n6621 & ~n6622;
  assign n6624 = ~n6341 & n6623;
  assign n6625 = n6341 & ~n6623;
  assign po43  = ~n6624 & ~n6625;
  assign n6627 = ~n6621 & ~n6624;
  assign n6628 = pi108  & n264;
  assign n6629 = pi106  & n281;
  assign n6630 = pi107  & n259;
  assign n6631 = ~n6629 & ~n6630;
  assign n6632 = ~n6628 & n6631;
  assign n6633 = ~n6610 & ~n6612;
  assign n6634 = ~pi107  & ~pi108 ;
  assign n6635 = pi107  & pi108 ;
  assign n6636 = ~n6634 & ~n6635;
  assign n6637 = ~n6633 & n6636;
  assign n6638 = n6633 & ~n6636;
  assign n6639 = ~n6637 & ~n6638;
  assign n6640 = n267 & n6639;
  assign n6641 = n6632 & ~n6640;
  assign n6642 = pi2  & ~n6641;
  assign n6643 = pi2  & ~n6642;
  assign n6644 = ~n6641 & ~n6642;
  assign n6645 = ~n6643 & ~n6644;
  assign n6646 = ~n6598 & ~n6600;
  assign n6647 = pi105  & n340;
  assign n6648 = pi103  & n380;
  assign n6649 = pi104  & n335;
  assign n6650 = ~n6648 & ~n6649;
  assign n6651 = ~n6647 & n6650;
  assign n6652 = n343 & n6065;
  assign n6653 = n6651 & ~n6652;
  assign n6654 = pi5  & ~n6653;
  assign n6655 = pi5  & ~n6654;
  assign n6656 = ~n6653 & ~n6654;
  assign n6657 = ~n6655 & ~n6656;
  assign n6658 = ~n6561 & ~n6565;
  assign n6659 = ~n6545 & ~n6547;
  assign n6660 = pi96  & n918;
  assign n6661 = pi94  & n1031;
  assign n6662 = pi95  & n913;
  assign n6663 = ~n6661 & ~n6662;
  assign n6664 = ~n6660 & n6663;
  assign n6665 = n921 & n3921;
  assign n6666 = n6664 & ~n6665;
  assign n6667 = pi14  & ~n6666;
  assign n6668 = pi14  & ~n6667;
  assign n6669 = ~n6666 & ~n6667;
  assign n6670 = ~n6668 & ~n6669;
  assign n6671 = ~n6538 & ~n6541;
  assign n6672 = pi93  & n1269;
  assign n6673 = pi91  & n1340;
  assign n6674 = pi92  & n1264;
  assign n6675 = ~n6673 & ~n6674;
  assign n6676 = ~n6672 & n6675;
  assign n6677 = n1272 & n3144;
  assign n6678 = n6676 & ~n6677;
  assign n6679 = pi17  & ~n6678;
  assign n6680 = pi17  & ~n6679;
  assign n6681 = ~n6678 & ~n6679;
  assign n6682 = ~n6680 & ~n6681;
  assign n6683 = ~n6532 & ~n6535;
  assign n6684 = ~n6515 & ~n6519;
  assign n6685 = ~n6479 & ~n6483;
  assign n6686 = pi81  & n2976;
  assign n6687 = pi79  & n3182;
  assign n6688 = pi80  & n2971;
  assign n6689 = ~n6687 & ~n6688;
  assign n6690 = ~n6686 & n6689;
  assign n6691 = n1413 & n2979;
  assign n6692 = n6690 & ~n6691;
  assign n6693 = pi29  & ~n6692;
  assign n6694 = pi29  & ~n6693;
  assign n6695 = ~n6692 & ~n6693;
  assign n6696 = ~n6694 & ~n6695;
  assign n6697 = ~n6463 & ~n6465;
  assign n6698 = pi78  & n3550;
  assign n6699 = pi76  & n3735;
  assign n6700 = pi77  & n3545;
  assign n6701 = ~n6699 & ~n6700;
  assign n6702 = ~n6698 & n6701;
  assign n6703 = n1009 & n3553;
  assign n6704 = n6702 & ~n6703;
  assign n6705 = pi32  & ~n6704;
  assign n6706 = pi32  & ~n6705;
  assign n6707 = ~n6704 & ~n6705;
  assign n6708 = ~n6706 & ~n6707;
  assign n6709 = pi75  & n4182;
  assign n6710 = pi73  & n4416;
  assign n6711 = pi74  & n4177;
  assign n6712 = ~n6710 & ~n6711;
  assign n6713 = ~n6709 & n6712;
  assign n6714 = n747 & n4185;
  assign n6715 = n6713 & ~n6714;
  assign n6716 = pi35  & ~n6715;
  assign n6717 = pi35  & ~n6716;
  assign n6718 = ~n6715 & ~n6716;
  assign n6719 = ~n6717 & ~n6718;
  assign n6720 = ~n6426 & ~n6430;
  assign n6721 = pi72  & n4896;
  assign n6722 = pi70  & n5148;
  assign n6723 = pi71  & n4891;
  assign n6724 = ~n6722 & ~n6723;
  assign n6725 = ~n6721 & n6724;
  assign n6726 = n575 & n4899;
  assign n6727 = n6725 & ~n6726;
  assign n6728 = pi38  & ~n6727;
  assign n6729 = pi38  & ~n6728;
  assign n6730 = ~n6727 & ~n6728;
  assign n6731 = ~n6729 & ~n6730;
  assign n6732 = ~n6410 & ~n6412;
  assign n6733 = pi66  & n6396;
  assign n6734 = n6175 & ~n6395;
  assign n6735 = n6390 & n6734;
  assign n6736 = pi64  & n6735;
  assign n6737 = pi65  & n6391;
  assign n6738 = ~n6736 & ~n6737;
  assign n6739 = ~n6733 & n6738;
  assign n6740 = n291 & n6399;
  assign n6741 = n6739 & ~n6740;
  assign n6742 = pi44  & ~n6741;
  assign n6743 = pi44  & ~n6742;
  assign n6744 = ~n6741 & ~n6742;
  assign n6745 = ~n6743 & ~n6744;
  assign n6746 = ~n6406 & n6745;
  assign n6747 = n6406 & ~n6745;
  assign n6748 = ~n6746 & ~n6747;
  assign n6749 = pi69  & n5636;
  assign n6750 = pi67  & n5909;
  assign n6751 = pi68  & n5631;
  assign n6752 = ~n6750 & ~n6751;
  assign n6753 = ~n6749 & n6752;
  assign n6754 = n405 & n5639;
  assign n6755 = n6753 & ~n6754;
  assign n6756 = pi41  & ~n6755;
  assign n6757 = pi41  & ~n6756;
  assign n6758 = ~n6755 & ~n6756;
  assign n6759 = ~n6757 & ~n6758;
  assign n6760 = n6748 & ~n6759;
  assign n6761 = ~n6748 & n6759;
  assign n6762 = ~n6760 & ~n6761;
  assign n6763 = ~n6732 & n6762;
  assign n6764 = n6732 & ~n6762;
  assign n6765 = ~n6763 & ~n6764;
  assign n6766 = ~n6731 & n6765;
  assign n6767 = n6731 & ~n6765;
  assign n6768 = ~n6766 & ~n6767;
  assign n6769 = ~n6720 & n6768;
  assign n6770 = n6720 & ~n6768;
  assign n6771 = ~n6769 & ~n6770;
  assign n6772 = n6719 & ~n6771;
  assign n6773 = ~n6719 & n6771;
  assign n6774 = ~n6772 & ~n6773;
  assign n6775 = ~n6448 & n6774;
  assign n6776 = n6448 & ~n6774;
  assign n6777 = ~n6775 & ~n6776;
  assign n6778 = n6708 & ~n6777;
  assign n6779 = ~n6708 & n6777;
  assign n6780 = ~n6778 & ~n6779;
  assign n6781 = ~n6697 & n6780;
  assign n6782 = n6697 & ~n6780;
  assign n6783 = ~n6781 & ~n6782;
  assign n6784 = n6696 & ~n6783;
  assign n6785 = ~n6696 & n6783;
  assign n6786 = ~n6784 & ~n6785;
  assign n6787 = ~n6685 & n6786;
  assign n6788 = n6685 & ~n6786;
  assign n6789 = ~n6787 & ~n6788;
  assign n6790 = pi84  & n2486;
  assign n6791 = pi82  & n2644;
  assign n6792 = pi83  & n2481;
  assign n6793 = ~n6791 & ~n6792;
  assign n6794 = ~n6790 & n6793;
  assign n6795 = n1805 & n2489;
  assign n6796 = n6794 & ~n6795;
  assign n6797 = pi26  & ~n6796;
  assign n6798 = pi26  & ~n6797;
  assign n6799 = ~n6796 & ~n6797;
  assign n6800 = ~n6798 & ~n6799;
  assign n6801 = n6789 & ~n6800;
  assign n6802 = n6789 & ~n6801;
  assign n6803 = ~n6800 & ~n6801;
  assign n6804 = ~n6802 & ~n6803;
  assign n6805 = ~n6496 & ~n6502;
  assign n6806 = n6804 & n6805;
  assign n6807 = ~n6804 & ~n6805;
  assign n6808 = ~n6806 & ~n6807;
  assign n6809 = pi87  & n2004;
  assign n6810 = pi85  & n2141;
  assign n6811 = pi86  & n1999;
  assign n6812 = ~n6810 & ~n6811;
  assign n6813 = ~n6809 & n6812;
  assign n6814 = n2007 & n2252;
  assign n6815 = n6813 & ~n6814;
  assign n6816 = pi23  & ~n6815;
  assign n6817 = pi23  & ~n6816;
  assign n6818 = ~n6815 & ~n6816;
  assign n6819 = ~n6817 & ~n6818;
  assign n6820 = n6808 & ~n6819;
  assign n6821 = ~n6808 & n6819;
  assign n6822 = ~n6684 & ~n6821;
  assign n6823 = ~n6820 & n6822;
  assign n6824 = ~n6684 & ~n6823;
  assign n6825 = ~n6820 & ~n6823;
  assign n6826 = ~n6821 & n6825;
  assign n6827 = ~n6824 & ~n6826;
  assign n6828 = pi90  & n1582;
  assign n6829 = pi88  & n1713;
  assign n6830 = pi89  & n1577;
  assign n6831 = ~n6829 & ~n6830;
  assign n6832 = ~n6828 & n6831;
  assign n6833 = n1585 & n2606;
  assign n6834 = n6832 & ~n6833;
  assign n6835 = pi20  & ~n6834;
  assign n6836 = pi20  & ~n6835;
  assign n6837 = ~n6834 & ~n6835;
  assign n6838 = ~n6836 & ~n6837;
  assign n6839 = n6827 & n6838;
  assign n6840 = ~n6827 & ~n6838;
  assign n6841 = ~n6839 & ~n6840;
  assign n6842 = ~n6683 & n6841;
  assign n6843 = n6683 & ~n6841;
  assign n6844 = ~n6842 & ~n6843;
  assign n6845 = n6682 & ~n6844;
  assign n6846 = ~n6682 & n6844;
  assign n6847 = ~n6845 & ~n6846;
  assign n6848 = ~n6671 & n6847;
  assign n6849 = n6671 & ~n6847;
  assign n6850 = ~n6848 & ~n6849;
  assign n6851 = n6670 & ~n6850;
  assign n6852 = ~n6670 & n6850;
  assign n6853 = ~n6851 & ~n6852;
  assign n6854 = ~n6659 & n6853;
  assign n6855 = n6659 & ~n6853;
  assign n6856 = ~n6854 & ~n6855;
  assign n6857 = pi99  & n675;
  assign n6858 = pi97  & n769;
  assign n6859 = pi98  & n670;
  assign n6860 = ~n6858 & ~n6859;
  assign n6861 = ~n6857 & n6860;
  assign n6862 = n678 & n4584;
  assign n6863 = n6861 & ~n6862;
  assign n6864 = pi11  & ~n6863;
  assign n6865 = pi11  & ~n6864;
  assign n6866 = ~n6863 & ~n6864;
  assign n6867 = ~n6865 & ~n6866;
  assign n6868 = n6856 & ~n6867;
  assign n6869 = ~n6856 & n6867;
  assign n6870 = ~n6868 & ~n6869;
  assign n6871 = n6658 & ~n6870;
  assign n6872 = ~n6658 & n6870;
  assign n6873 = ~n6871 & ~n6872;
  assign n6874 = pi102  & n493;
  assign n6875 = pi100  & n533;
  assign n6876 = pi101  & n488;
  assign n6877 = ~n6875 & ~n6876;
  assign n6878 = ~n6874 & n6877;
  assign n6879 = n496 & n5296;
  assign n6880 = n6878 & ~n6879;
  assign n6881 = pi8  & ~n6880;
  assign n6882 = pi8  & ~n6881;
  assign n6883 = ~n6880 & ~n6881;
  assign n6884 = ~n6882 & ~n6883;
  assign n6885 = n6873 & ~n6884;
  assign n6886 = ~n6873 & n6884;
  assign n6887 = ~n6885 & ~n6886;
  assign n6888 = ~n6583 & n6887;
  assign n6889 = n6583 & ~n6887;
  assign n6890 = ~n6888 & ~n6889;
  assign n6891 = ~n6657 & n6890;
  assign n6892 = n6657 & ~n6890;
  assign n6893 = ~n6891 & ~n6892;
  assign n6894 = ~n6646 & n6893;
  assign n6895 = n6646 & ~n6893;
  assign n6896 = ~n6894 & ~n6895;
  assign n6897 = ~n6645 & n6896;
  assign n6898 = n6645 & ~n6896;
  assign n6899 = ~n6897 & ~n6898;
  assign n6900 = ~n6627 & n6899;
  assign n6901 = n6627 & ~n6899;
  assign po44  = ~n6900 & ~n6901;
  assign n6903 = ~n6897 & ~n6900;
  assign n6904 = ~n6891 & ~n6894;
  assign n6905 = ~n6885 & ~n6888;
  assign n6906 = ~n6868 & ~n6872;
  assign n6907 = pi100  & n675;
  assign n6908 = pi98  & n769;
  assign n6909 = pi99  & n670;
  assign n6910 = ~n6908 & ~n6909;
  assign n6911 = ~n6907 & n6910;
  assign n6912 = n678 & n4808;
  assign n6913 = n6911 & ~n6912;
  assign n6914 = pi11  & ~n6913;
  assign n6915 = pi11  & ~n6914;
  assign n6916 = ~n6913 & ~n6914;
  assign n6917 = ~n6915 & ~n6916;
  assign n6918 = ~n6852 & ~n6854;
  assign n6919 = ~n6846 & ~n6848;
  assign n6920 = pi94  & n1269;
  assign n6921 = pi92  & n1340;
  assign n6922 = pi93  & n1264;
  assign n6923 = ~n6921 & ~n6922;
  assign n6924 = ~n6920 & n6923;
  assign n6925 = n1272 & n3499;
  assign n6926 = n6924 & ~n6925;
  assign n6927 = pi17  & ~n6926;
  assign n6928 = pi17  & ~n6927;
  assign n6929 = ~n6926 & ~n6927;
  assign n6930 = ~n6928 & ~n6929;
  assign n6931 = ~n6840 & ~n6842;
  assign n6932 = ~n6785 & ~n6787;
  assign n6933 = pi82  & n2976;
  assign n6934 = pi80  & n3182;
  assign n6935 = pi81  & n2971;
  assign n6936 = ~n6934 & ~n6935;
  assign n6937 = ~n6933 & n6936;
  assign n6938 = n1532 & n2979;
  assign n6939 = n6937 & ~n6938;
  assign n6940 = pi29  & ~n6939;
  assign n6941 = pi29  & ~n6940;
  assign n6942 = ~n6939 & ~n6940;
  assign n6943 = ~n6941 & ~n6942;
  assign n6944 = ~n6779 & ~n6781;
  assign n6945 = ~n6773 & ~n6775;
  assign n6946 = pi76  & n4182;
  assign n6947 = pi74  & n4416;
  assign n6948 = pi75  & n4177;
  assign n6949 = ~n6947 & ~n6948;
  assign n6950 = ~n6946 & n6949;
  assign n6951 = n881 & n4185;
  assign n6952 = n6950 & ~n6951;
  assign n6953 = pi35  & ~n6952;
  assign n6954 = pi35  & ~n6953;
  assign n6955 = ~n6952 & ~n6953;
  assign n6956 = ~n6954 & ~n6955;
  assign n6957 = ~n6766 & ~n6769;
  assign n6958 = ~n6760 & ~n6763;
  assign n6959 = pi67  & n6396;
  assign n6960 = pi65  & n6735;
  assign n6961 = pi66  & n6391;
  assign n6962 = ~n6960 & ~n6961;
  assign n6963 = ~n6959 & n6962;
  assign n6964 = n313 & n6399;
  assign n6965 = n6963 & ~n6964;
  assign n6966 = pi44  & ~n6965;
  assign n6967 = pi44  & ~n6966;
  assign n6968 = ~n6965 & ~n6966;
  assign n6969 = ~n6967 & ~n6968;
  assign n6970 = pi44  & ~pi45 ;
  assign n6971 = ~pi44  & pi45 ;
  assign n6972 = ~n6970 & ~n6971;
  assign n6973 = pi64  & ~n6972;
  assign n6974 = n6747 & n6973;
  assign n6975 = ~n6747 & ~n6973;
  assign n6976 = ~n6974 & ~n6975;
  assign n6977 = ~n6969 & n6976;
  assign n6978 = n6969 & ~n6976;
  assign n6979 = ~n6977 & ~n6978;
  assign n6980 = pi70  & n5636;
  assign n6981 = pi68  & n5909;
  assign n6982 = pi69  & n5631;
  assign n6983 = ~n6981 & ~n6982;
  assign n6984 = ~n6980 & n6983;
  assign n6985 = n430 & n5639;
  assign n6986 = n6984 & ~n6985;
  assign n6987 = pi41  & ~n6986;
  assign n6988 = pi41  & ~n6987;
  assign n6989 = ~n6986 & ~n6987;
  assign n6990 = ~n6988 & ~n6989;
  assign n6991 = n6979 & ~n6990;
  assign n6992 = ~n6979 & n6990;
  assign n6993 = ~n6991 & ~n6992;
  assign n6994 = n6958 & ~n6993;
  assign n6995 = ~n6958 & n6993;
  assign n6996 = ~n6994 & ~n6995;
  assign n6997 = pi73  & n4896;
  assign n6998 = pi71  & n5148;
  assign n6999 = pi72  & n4891;
  assign n7000 = ~n6998 & ~n6999;
  assign n7001 = ~n6997 & n7000;
  assign n7002 = n639 & n4899;
  assign n7003 = n7001 & ~n7002;
  assign n7004 = pi38  & ~n7003;
  assign n7005 = pi38  & ~n7004;
  assign n7006 = ~n7003 & ~n7004;
  assign n7007 = ~n7005 & ~n7006;
  assign n7008 = ~n6996 & n7007;
  assign n7009 = n6996 & ~n7007;
  assign n7010 = ~n7008 & ~n7009;
  assign n7011 = ~n6957 & n7010;
  assign n7012 = n6957 & ~n7010;
  assign n7013 = ~n7011 & ~n7012;
  assign n7014 = ~n6956 & n7013;
  assign n7015 = n6956 & ~n7013;
  assign n7016 = ~n7014 & ~n7015;
  assign n7017 = ~n6945 & n7016;
  assign n7018 = n6945 & ~n7016;
  assign n7019 = ~n7017 & ~n7018;
  assign n7020 = pi79  & n3550;
  assign n7021 = pi77  & n3735;
  assign n7022 = pi78  & n3545;
  assign n7023 = ~n7021 & ~n7022;
  assign n7024 = ~n7020 & n7023;
  assign n7025 = n1105 & n3553;
  assign n7026 = n7024 & ~n7025;
  assign n7027 = pi32  & ~n7026;
  assign n7028 = pi32  & ~n7027;
  assign n7029 = ~n7026 & ~n7027;
  assign n7030 = ~n7028 & ~n7029;
  assign n7031 = n7019 & ~n7030;
  assign n7032 = ~n7019 & n7030;
  assign n7033 = ~n7031 & ~n7032;
  assign n7034 = ~n6944 & n7033;
  assign n7035 = n6944 & ~n7033;
  assign n7036 = ~n7034 & ~n7035;
  assign n7037 = ~n6943 & n7036;
  assign n7038 = n6943 & ~n7036;
  assign n7039 = ~n7037 & ~n7038;
  assign n7040 = ~n6932 & n7039;
  assign n7041 = n6932 & ~n7039;
  assign n7042 = ~n7040 & ~n7041;
  assign n7043 = pi85  & n2486;
  assign n7044 = pi83  & n2644;
  assign n7045 = pi84  & n2481;
  assign n7046 = ~n7044 & ~n7045;
  assign n7047 = ~n7043 & n7046;
  assign n7048 = n1943 & n2489;
  assign n7049 = n7047 & ~n7048;
  assign n7050 = pi26  & ~n7049;
  assign n7051 = pi26  & ~n7050;
  assign n7052 = ~n7049 & ~n7050;
  assign n7053 = ~n7051 & ~n7052;
  assign n7054 = n7042 & ~n7053;
  assign n7055 = n7042 & ~n7054;
  assign n7056 = ~n7053 & ~n7054;
  assign n7057 = ~n7055 & ~n7056;
  assign n7058 = ~n6801 & ~n6807;
  assign n7059 = n7057 & n7058;
  assign n7060 = ~n7057 & ~n7058;
  assign n7061 = ~n7059 & ~n7060;
  assign n7062 = pi88  & n2004;
  assign n7063 = pi86  & n2141;
  assign n7064 = pi87  & n1999;
  assign n7065 = ~n7063 & ~n7064;
  assign n7066 = ~n7062 & n7065;
  assign n7067 = n2007 & n2277;
  assign n7068 = n7066 & ~n7067;
  assign n7069 = pi23  & ~n7068;
  assign n7070 = pi23  & ~n7069;
  assign n7071 = ~n7068 & ~n7069;
  assign n7072 = ~n7070 & ~n7071;
  assign n7073 = ~n7061 & n7072;
  assign n7074 = n7061 & ~n7072;
  assign n7075 = ~n7073 & ~n7074;
  assign n7076 = ~n6825 & n7075;
  assign n7077 = n6825 & ~n7075;
  assign n7078 = ~n7076 & ~n7077;
  assign n7079 = pi91  & n1582;
  assign n7080 = pi89  & n1713;
  assign n7081 = pi90  & n1577;
  assign n7082 = ~n7080 & ~n7081;
  assign n7083 = ~n7079 & n7082;
  assign n7084 = n1585 & n2926;
  assign n7085 = n7083 & ~n7084;
  assign n7086 = pi20  & ~n7085;
  assign n7087 = pi20  & ~n7086;
  assign n7088 = ~n7085 & ~n7086;
  assign n7089 = ~n7087 & ~n7088;
  assign n7090 = n7078 & ~n7089;
  assign n7091 = ~n7078 & n7089;
  assign n7092 = ~n7090 & ~n7091;
  assign n7093 = ~n6931 & n7092;
  assign n7094 = n6931 & ~n7092;
  assign n7095 = ~n7093 & ~n7094;
  assign n7096 = ~n6930 & n7095;
  assign n7097 = n6930 & ~n7095;
  assign n7098 = ~n7096 & ~n7097;
  assign n7099 = ~n6919 & n7098;
  assign n7100 = n6919 & ~n7098;
  assign n7101 = ~n7099 & ~n7100;
  assign n7102 = pi97  & n918;
  assign n7103 = pi95  & n1031;
  assign n7104 = pi96  & n913;
  assign n7105 = ~n7103 & ~n7104;
  assign n7106 = ~n7102 & n7105;
  assign n7107 = n921 & n3946;
  assign n7108 = n7106 & ~n7107;
  assign n7109 = pi14  & ~n7108;
  assign n7110 = pi14  & ~n7109;
  assign n7111 = ~n7108 & ~n7109;
  assign n7112 = ~n7110 & ~n7111;
  assign n7113 = n7101 & ~n7112;
  assign n7114 = ~n7101 & n7112;
  assign n7115 = ~n7113 & ~n7114;
  assign n7116 = ~n6918 & n7115;
  assign n7117 = n6918 & ~n7115;
  assign n7118 = ~n7116 & ~n7117;
  assign n7119 = ~n6917 & n7118;
  assign n7120 = n6917 & ~n7118;
  assign n7121 = ~n7119 & ~n7120;
  assign n7122 = n6906 & ~n7121;
  assign n7123 = ~n6906 & n7121;
  assign n7124 = ~n7122 & ~n7123;
  assign n7125 = pi103  & n493;
  assign n7126 = pi101  & n533;
  assign n7127 = pi102  & n488;
  assign n7128 = ~n7126 & ~n7127;
  assign n7129 = ~n7125 & n7128;
  assign n7130 = n496 & n5540;
  assign n7131 = n7129 & ~n7130;
  assign n7132 = pi8  & ~n7131;
  assign n7133 = pi8  & ~n7132;
  assign n7134 = ~n7131 & ~n7132;
  assign n7135 = ~n7133 & ~n7134;
  assign n7136 = n7124 & ~n7135;
  assign n7137 = ~n7124 & n7135;
  assign n7138 = ~n7136 & ~n7137;
  assign n7139 = n6905 & ~n7138;
  assign n7140 = ~n6905 & n7138;
  assign n7141 = ~n7139 & ~n7140;
  assign n7142 = pi106  & n340;
  assign n7143 = pi104  & n380;
  assign n7144 = pi105  & n335;
  assign n7145 = ~n7143 & ~n7144;
  assign n7146 = ~n7142 & n7145;
  assign n7147 = n343 & n6090;
  assign n7148 = n7146 & ~n7147;
  assign n7149 = pi5  & ~n7148;
  assign n7150 = pi5  & ~n7149;
  assign n7151 = ~n7148 & ~n7149;
  assign n7152 = ~n7150 & ~n7151;
  assign n7153 = n7141 & ~n7152;
  assign n7154 = ~n7141 & n7152;
  assign n7155 = ~n7153 & ~n7154;
  assign n7156 = n6904 & ~n7155;
  assign n7157 = ~n6904 & n7155;
  assign n7158 = ~n7156 & ~n7157;
  assign n7159 = pi109  & n264;
  assign n7160 = pi107  & n281;
  assign n7161 = pi108  & n259;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = ~n7159 & n7162;
  assign n7164 = ~n6635 & ~n6637;
  assign n7165 = ~pi108  & ~pi109 ;
  assign n7166 = pi108  & pi109 ;
  assign n7167 = ~n7165 & ~n7166;
  assign n7168 = ~n7164 & n7167;
  assign n7169 = n7164 & ~n7167;
  assign n7170 = ~n7168 & ~n7169;
  assign n7171 = n267 & n7170;
  assign n7172 = n7163 & ~n7171;
  assign n7173 = pi2  & ~n7172;
  assign n7174 = pi2  & ~n7173;
  assign n7175 = ~n7172 & ~n7173;
  assign n7176 = ~n7174 & ~n7175;
  assign n7177 = ~n7158 & n7176;
  assign n7178 = n7158 & ~n7176;
  assign n7179 = ~n7177 & ~n7178;
  assign n7180 = ~n6903 & n7179;
  assign n7181 = n6903 & ~n7179;
  assign po45  = ~n7180 & ~n7181;
  assign n7183 = ~n7178 & ~n7180;
  assign n7184 = ~n7153 & ~n7157;
  assign n7185 = ~n7136 & ~n7140;
  assign n7186 = ~n7119 & ~n7123;
  assign n7187 = ~n7113 & ~n7116;
  assign n7188 = ~n7096 & ~n7099;
  assign n7189 = pi95  & n1269;
  assign n7190 = pi93  & n1340;
  assign n7191 = pi94  & n1264;
  assign n7192 = ~n7190 & ~n7191;
  assign n7193 = ~n7189 & n7192;
  assign n7194 = n1272 & n3710;
  assign n7195 = n7193 & ~n7194;
  assign n7196 = pi17  & ~n7195;
  assign n7197 = pi17  & ~n7196;
  assign n7198 = ~n7195 & ~n7196;
  assign n7199 = ~n7197 & ~n7198;
  assign n7200 = ~n7090 & ~n7093;
  assign n7201 = pi92  & n1582;
  assign n7202 = pi90  & n1713;
  assign n7203 = pi91  & n1577;
  assign n7204 = ~n7202 & ~n7203;
  assign n7205 = ~n7201 & n7204;
  assign n7206 = n1585 & n3119;
  assign n7207 = n7205 & ~n7206;
  assign n7208 = pi20  & ~n7207;
  assign n7209 = pi20  & ~n7208;
  assign n7210 = ~n7207 & ~n7208;
  assign n7211 = ~n7209 & ~n7210;
  assign n7212 = ~n7074 & ~n7076;
  assign n7213 = ~n7037 & ~n7040;
  assign n7214 = ~n7031 & ~n7034;
  assign n7215 = ~n7014 & ~n7017;
  assign n7216 = ~n7009 & ~n7011;
  assign n7217 = ~n6991 & ~n6995;
  assign n7218 = ~n6974 & ~n6977;
  assign n7219 = pi68  & n6396;
  assign n7220 = pi66  & n6735;
  assign n7221 = pi67  & n6391;
  assign n7222 = ~n7220 & ~n7221;
  assign n7223 = ~n7219 & n7222;
  assign n7224 = n364 & n6399;
  assign n7225 = n7223 & ~n7224;
  assign n7226 = pi44  & ~n7225;
  assign n7227 = pi44  & ~n7226;
  assign n7228 = ~n7225 & ~n7226;
  assign n7229 = ~n7227 & ~n7228;
  assign n7230 = pi47  & ~n6973;
  assign n7231 = ~pi45  & pi46 ;
  assign n7232 = pi45  & ~pi46 ;
  assign n7233 = ~n7231 & ~n7232;
  assign n7234 = n6972 & ~n7233;
  assign n7235 = pi64  & n7234;
  assign n7236 = ~pi46  & pi47 ;
  assign n7237 = pi46  & ~pi47 ;
  assign n7238 = ~n7236 & ~n7237;
  assign n7239 = ~n6972 & n7238;
  assign n7240 = pi65  & n7239;
  assign n7241 = ~n7235 & ~n7240;
  assign n7242 = ~n6972 & ~n7238;
  assign n7243 = n270 & n7242;
  assign n7244 = n7241 & ~n7243;
  assign n7245 = pi47  & ~n7244;
  assign n7246 = pi47  & ~n7245;
  assign n7247 = ~n7244 & ~n7245;
  assign n7248 = ~n7246 & ~n7247;
  assign n7249 = n7230 & ~n7248;
  assign n7250 = ~n7230 & n7248;
  assign n7251 = ~n7249 & ~n7250;
  assign n7252 = n7229 & ~n7251;
  assign n7253 = ~n7229 & n7251;
  assign n7254 = ~n7252 & ~n7253;
  assign n7255 = ~n7218 & n7254;
  assign n7256 = n7218 & ~n7254;
  assign n7257 = ~n7255 & ~n7256;
  assign n7258 = pi71  & n5636;
  assign n7259 = pi69  & n5909;
  assign n7260 = pi70  & n5631;
  assign n7261 = ~n7259 & ~n7260;
  assign n7262 = ~n7258 & n7261;
  assign n7263 = n476 & n5639;
  assign n7264 = n7262 & ~n7263;
  assign n7265 = pi41  & ~n7264;
  assign n7266 = pi41  & ~n7265;
  assign n7267 = ~n7264 & ~n7265;
  assign n7268 = ~n7266 & ~n7267;
  assign n7269 = n7257 & ~n7268;
  assign n7270 = ~n7257 & n7268;
  assign n7271 = ~n7269 & ~n7270;
  assign n7272 = n7217 & ~n7271;
  assign n7273 = ~n7217 & n7271;
  assign n7274 = ~n7272 & ~n7273;
  assign n7275 = pi74  & n4896;
  assign n7276 = pi72  & n5148;
  assign n7277 = pi73  & n4891;
  assign n7278 = ~n7276 & ~n7277;
  assign n7279 = ~n7275 & n7278;
  assign n7280 = n722 & n4899;
  assign n7281 = n7279 & ~n7280;
  assign n7282 = pi38  & ~n7281;
  assign n7283 = pi38  & ~n7282;
  assign n7284 = ~n7281 & ~n7282;
  assign n7285 = ~n7283 & ~n7284;
  assign n7286 = n7274 & ~n7285;
  assign n7287 = ~n7274 & n7285;
  assign n7288 = ~n7216 & ~n7287;
  assign n7289 = ~n7286 & n7288;
  assign n7290 = ~n7216 & ~n7289;
  assign n7291 = ~n7286 & ~n7289;
  assign n7292 = ~n7287 & n7291;
  assign n7293 = ~n7290 & ~n7292;
  assign n7294 = pi77  & n4182;
  assign n7295 = pi75  & n4416;
  assign n7296 = pi76  & n4177;
  assign n7297 = ~n7295 & ~n7296;
  assign n7298 = ~n7294 & n7297;
  assign n7299 = n984 & n4185;
  assign n7300 = n7298 & ~n7299;
  assign n7301 = pi35  & ~n7300;
  assign n7302 = pi35  & ~n7301;
  assign n7303 = ~n7300 & ~n7301;
  assign n7304 = ~n7302 & ~n7303;
  assign n7305 = n7293 & n7304;
  assign n7306 = ~n7293 & ~n7304;
  assign n7307 = ~n7305 & ~n7306;
  assign n7308 = ~n7215 & n7307;
  assign n7309 = n7215 & ~n7307;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = pi80  & n3550;
  assign n7312 = pi78  & n3735;
  assign n7313 = pi79  & n3545;
  assign n7314 = ~n7312 & ~n7313;
  assign n7315 = ~n7311 & n7314;
  assign n7316 = n1205 & n3553;
  assign n7317 = n7315 & ~n7316;
  assign n7318 = pi32  & ~n7317;
  assign n7319 = pi32  & ~n7318;
  assign n7320 = ~n7317 & ~n7318;
  assign n7321 = ~n7319 & ~n7320;
  assign n7322 = n7310 & ~n7321;
  assign n7323 = ~n7310 & n7321;
  assign n7324 = ~n7322 & ~n7323;
  assign n7325 = n7214 & ~n7324;
  assign n7326 = ~n7214 & n7324;
  assign n7327 = ~n7325 & ~n7326;
  assign n7328 = pi83  & n2976;
  assign n7329 = pi81  & n3182;
  assign n7330 = pi82  & n2971;
  assign n7331 = ~n7329 & ~n7330;
  assign n7332 = ~n7328 & n7331;
  assign n7333 = n1672 & n2979;
  assign n7334 = n7332 & ~n7333;
  assign n7335 = pi29  & ~n7334;
  assign n7336 = pi29  & ~n7335;
  assign n7337 = ~n7334 & ~n7335;
  assign n7338 = ~n7336 & ~n7337;
  assign n7339 = n7327 & ~n7338;
  assign n7340 = ~n7327 & n7338;
  assign n7341 = ~n7339 & ~n7340;
  assign n7342 = n7213 & ~n7341;
  assign n7343 = ~n7213 & n7341;
  assign n7344 = ~n7342 & ~n7343;
  assign n7345 = pi86  & n2486;
  assign n7346 = pi84  & n2644;
  assign n7347 = pi85  & n2481;
  assign n7348 = ~n7346 & ~n7347;
  assign n7349 = ~n7345 & n7348;
  assign n7350 = n2099 & n2489;
  assign n7351 = n7349 & ~n7350;
  assign n7352 = pi26  & ~n7351;
  assign n7353 = pi26  & ~n7352;
  assign n7354 = ~n7351 & ~n7352;
  assign n7355 = ~n7353 & ~n7354;
  assign n7356 = n7344 & ~n7355;
  assign n7357 = n7344 & ~n7356;
  assign n7358 = ~n7355 & ~n7356;
  assign n7359 = ~n7357 & ~n7358;
  assign n7360 = ~n7054 & ~n7060;
  assign n7361 = n7359 & n7360;
  assign n7362 = ~n7359 & ~n7360;
  assign n7363 = ~n7361 & ~n7362;
  assign n7364 = pi89  & n2004;
  assign n7365 = pi87  & n2141;
  assign n7366 = pi88  & n1999;
  assign n7367 = ~n7365 & ~n7366;
  assign n7368 = ~n7364 & n7367;
  assign n7369 = n2007 & n2432;
  assign n7370 = n7368 & ~n7369;
  assign n7371 = pi23  & ~n7370;
  assign n7372 = pi23  & ~n7371;
  assign n7373 = ~n7370 & ~n7371;
  assign n7374 = ~n7372 & ~n7373;
  assign n7375 = n7363 & ~n7374;
  assign n7376 = ~n7363 & n7374;
  assign n7377 = ~n7375 & ~n7376;
  assign n7378 = ~n7212 & n7377;
  assign n7379 = n7212 & ~n7377;
  assign n7380 = ~n7378 & ~n7379;
  assign n7381 = ~n7211 & n7380;
  assign n7382 = n7211 & ~n7380;
  assign n7383 = ~n7381 & ~n7382;
  assign n7384 = ~n7200 & n7383;
  assign n7385 = n7200 & ~n7383;
  assign n7386 = ~n7384 & ~n7385;
  assign n7387 = n7199 & ~n7386;
  assign n7388 = ~n7199 & n7386;
  assign n7389 = ~n7387 & ~n7388;
  assign n7390 = ~n7188 & n7389;
  assign n7391 = n7188 & ~n7389;
  assign n7392 = ~n7390 & ~n7391;
  assign n7393 = pi98  & n918;
  assign n7394 = pi96  & n1031;
  assign n7395 = pi97  & n913;
  assign n7396 = ~n7394 & ~n7395;
  assign n7397 = ~n7393 & n7396;
  assign n7398 = n921 & n4360;
  assign n7399 = n7397 & ~n7398;
  assign n7400 = pi14  & ~n7399;
  assign n7401 = pi14  & ~n7400;
  assign n7402 = ~n7399 & ~n7400;
  assign n7403 = ~n7401 & ~n7402;
  assign n7404 = n7392 & ~n7403;
  assign n7405 = ~n7392 & n7403;
  assign n7406 = ~n7404 & ~n7405;
  assign n7407 = n7187 & ~n7406;
  assign n7408 = ~n7187 & n7406;
  assign n7409 = ~n7407 & ~n7408;
  assign n7410 = pi101  & n675;
  assign n7411 = pi99  & n769;
  assign n7412 = pi100  & n670;
  assign n7413 = ~n7411 & ~n7412;
  assign n7414 = ~n7410 & n7413;
  assign n7415 = n678 & n5056;
  assign n7416 = n7414 & ~n7415;
  assign n7417 = pi11  & ~n7416;
  assign n7418 = pi11  & ~n7417;
  assign n7419 = ~n7416 & ~n7417;
  assign n7420 = ~n7418 & ~n7419;
  assign n7421 = n7409 & ~n7420;
  assign n7422 = ~n7409 & n7420;
  assign n7423 = ~n7421 & ~n7422;
  assign n7424 = n7186 & ~n7423;
  assign n7425 = ~n7186 & n7423;
  assign n7426 = ~n7424 & ~n7425;
  assign n7427 = pi104  & n493;
  assign n7428 = pi102  & n533;
  assign n7429 = pi103  & n488;
  assign n7430 = ~n7428 & ~n7429;
  assign n7431 = ~n7427 & n7430;
  assign n7432 = n496 & n5565;
  assign n7433 = n7431 & ~n7432;
  assign n7434 = pi8  & ~n7433;
  assign n7435 = pi8  & ~n7434;
  assign n7436 = ~n7433 & ~n7434;
  assign n7437 = ~n7435 & ~n7436;
  assign n7438 = n7426 & ~n7437;
  assign n7439 = ~n7426 & n7437;
  assign n7440 = ~n7185 & ~n7439;
  assign n7441 = ~n7438 & n7440;
  assign n7442 = ~n7185 & ~n7441;
  assign n7443 = ~n7438 & ~n7441;
  assign n7444 = ~n7439 & n7443;
  assign n7445 = ~n7442 & ~n7444;
  assign n7446 = pi107  & n340;
  assign n7447 = pi105  & n380;
  assign n7448 = pi106  & n335;
  assign n7449 = ~n7447 & ~n7448;
  assign n7450 = ~n7446 & n7449;
  assign n7451 = n343 & n6614;
  assign n7452 = n7450 & ~n7451;
  assign n7453 = pi5  & ~n7452;
  assign n7454 = pi5  & ~n7453;
  assign n7455 = ~n7452 & ~n7453;
  assign n7456 = ~n7454 & ~n7455;
  assign n7457 = ~n7445 & ~n7456;
  assign n7458 = n7445 & n7456;
  assign n7459 = ~n7457 & ~n7458;
  assign n7460 = n7184 & ~n7459;
  assign n7461 = ~n7184 & n7459;
  assign n7462 = ~n7460 & ~n7461;
  assign n7463 = pi110  & n264;
  assign n7464 = pi108  & n281;
  assign n7465 = pi109  & n259;
  assign n7466 = ~n7464 & ~n7465;
  assign n7467 = ~n7463 & n7466;
  assign n7468 = ~n7166 & ~n7168;
  assign n7469 = ~pi109  & ~pi110 ;
  assign n7470 = pi109  & pi110 ;
  assign n7471 = ~n7469 & ~n7470;
  assign n7472 = ~n7468 & n7471;
  assign n7473 = n7468 & ~n7471;
  assign n7474 = ~n7472 & ~n7473;
  assign n7475 = n267 & n7474;
  assign n7476 = n7467 & ~n7475;
  assign n7477 = pi2  & ~n7476;
  assign n7478 = pi2  & ~n7477;
  assign n7479 = ~n7476 & ~n7477;
  assign n7480 = ~n7478 & ~n7479;
  assign n7481 = n7462 & ~n7480;
  assign n7482 = ~n7462 & n7480;
  assign n7483 = ~n7481 & ~n7482;
  assign n7484 = ~n7183 & n7483;
  assign n7485 = n7183 & ~n7483;
  assign po46  = ~n7484 & ~n7485;
  assign n7487 = ~n7481 & ~n7484;
  assign n7488 = ~n7457 & ~n7461;
  assign n7489 = ~n7421 & ~n7425;
  assign n7490 = ~n7404 & ~n7408;
  assign n7491 = ~n7388 & ~n7390;
  assign n7492 = pi96  & n1269;
  assign n7493 = pi94  & n1340;
  assign n7494 = pi95  & n1264;
  assign n7495 = ~n7493 & ~n7494;
  assign n7496 = ~n7492 & n7495;
  assign n7497 = n1272 & n3921;
  assign n7498 = n7496 & ~n7497;
  assign n7499 = pi17  & ~n7498;
  assign n7500 = pi17  & ~n7499;
  assign n7501 = ~n7498 & ~n7499;
  assign n7502 = ~n7500 & ~n7501;
  assign n7503 = ~n7381 & ~n7384;
  assign n7504 = pi93  & n1582;
  assign n7505 = pi91  & n1713;
  assign n7506 = pi92  & n1577;
  assign n7507 = ~n7505 & ~n7506;
  assign n7508 = ~n7504 & n7507;
  assign n7509 = n1585 & n3144;
  assign n7510 = n7508 & ~n7509;
  assign n7511 = pi20  & ~n7510;
  assign n7512 = pi20  & ~n7511;
  assign n7513 = ~n7510 & ~n7511;
  assign n7514 = ~n7512 & ~n7513;
  assign n7515 = ~n7375 & ~n7378;
  assign n7516 = ~n7356 & ~n7362;
  assign n7517 = ~n7322 & ~n7326;
  assign n7518 = pi81  & n3550;
  assign n7519 = pi79  & n3735;
  assign n7520 = pi80  & n3545;
  assign n7521 = ~n7519 & ~n7520;
  assign n7522 = ~n7518 & n7521;
  assign n7523 = n1413 & n3553;
  assign n7524 = n7522 & ~n7523;
  assign n7525 = pi32  & ~n7524;
  assign n7526 = pi32  & ~n7525;
  assign n7527 = ~n7524 & ~n7525;
  assign n7528 = ~n7526 & ~n7527;
  assign n7529 = ~n7306 & ~n7308;
  assign n7530 = pi75  & n4896;
  assign n7531 = pi73  & n5148;
  assign n7532 = pi74  & n4891;
  assign n7533 = ~n7531 & ~n7532;
  assign n7534 = ~n7530 & n7533;
  assign n7535 = n747 & n4899;
  assign n7536 = n7534 & ~n7535;
  assign n7537 = pi38  & ~n7536;
  assign n7538 = pi38  & ~n7537;
  assign n7539 = ~n7536 & ~n7537;
  assign n7540 = ~n7538 & ~n7539;
  assign n7541 = ~n7269 & ~n7273;
  assign n7542 = pi72  & n5636;
  assign n7543 = pi70  & n5909;
  assign n7544 = pi71  & n5631;
  assign n7545 = ~n7543 & ~n7544;
  assign n7546 = ~n7542 & n7545;
  assign n7547 = n575 & n5639;
  assign n7548 = n7546 & ~n7547;
  assign n7549 = pi41  & ~n7548;
  assign n7550 = pi41  & ~n7549;
  assign n7551 = ~n7548 & ~n7549;
  assign n7552 = ~n7550 & ~n7551;
  assign n7553 = ~n7253 & ~n7255;
  assign n7554 = pi66  & n7239;
  assign n7555 = n6972 & ~n7238;
  assign n7556 = n7233 & n7555;
  assign n7557 = pi64  & n7556;
  assign n7558 = pi65  & n7234;
  assign n7559 = ~n7557 & ~n7558;
  assign n7560 = ~n7554 & n7559;
  assign n7561 = n291 & n7242;
  assign n7562 = n7560 & ~n7561;
  assign n7563 = pi47  & ~n7562;
  assign n7564 = pi47  & ~n7563;
  assign n7565 = ~n7562 & ~n7563;
  assign n7566 = ~n7564 & ~n7565;
  assign n7567 = ~n7249 & n7566;
  assign n7568 = n7249 & ~n7566;
  assign n7569 = ~n7567 & ~n7568;
  assign n7570 = pi69  & n6396;
  assign n7571 = pi67  & n6735;
  assign n7572 = pi68  & n6391;
  assign n7573 = ~n7571 & ~n7572;
  assign n7574 = ~n7570 & n7573;
  assign n7575 = n405 & n6399;
  assign n7576 = n7574 & ~n7575;
  assign n7577 = pi44  & ~n7576;
  assign n7578 = pi44  & ~n7577;
  assign n7579 = ~n7576 & ~n7577;
  assign n7580 = ~n7578 & ~n7579;
  assign n7581 = n7569 & ~n7580;
  assign n7582 = ~n7569 & n7580;
  assign n7583 = ~n7581 & ~n7582;
  assign n7584 = ~n7553 & n7583;
  assign n7585 = n7553 & ~n7583;
  assign n7586 = ~n7584 & ~n7585;
  assign n7587 = ~n7552 & n7586;
  assign n7588 = n7552 & ~n7586;
  assign n7589 = ~n7587 & ~n7588;
  assign n7590 = ~n7541 & n7589;
  assign n7591 = n7541 & ~n7589;
  assign n7592 = ~n7590 & ~n7591;
  assign n7593 = n7540 & ~n7592;
  assign n7594 = ~n7540 & n7592;
  assign n7595 = ~n7593 & ~n7594;
  assign n7596 = ~n7291 & n7595;
  assign n7597 = n7291 & ~n7595;
  assign n7598 = ~n7596 & ~n7597;
  assign n7599 = pi78  & n4182;
  assign n7600 = pi76  & n4416;
  assign n7601 = pi77  & n4177;
  assign n7602 = ~n7600 & ~n7601;
  assign n7603 = ~n7599 & n7602;
  assign n7604 = n1009 & n4185;
  assign n7605 = n7603 & ~n7604;
  assign n7606 = pi35  & ~n7605;
  assign n7607 = pi35  & ~n7606;
  assign n7608 = ~n7605 & ~n7606;
  assign n7609 = ~n7607 & ~n7608;
  assign n7610 = n7598 & ~n7609;
  assign n7611 = ~n7598 & n7609;
  assign n7612 = ~n7610 & ~n7611;
  assign n7613 = ~n7529 & n7612;
  assign n7614 = n7529 & ~n7612;
  assign n7615 = ~n7613 & ~n7614;
  assign n7616 = ~n7528 & n7615;
  assign n7617 = n7528 & ~n7615;
  assign n7618 = ~n7616 & ~n7617;
  assign n7619 = ~n7517 & n7618;
  assign n7620 = n7517 & ~n7618;
  assign n7621 = ~n7619 & ~n7620;
  assign n7622 = pi84  & n2976;
  assign n7623 = pi82  & n3182;
  assign n7624 = pi83  & n2971;
  assign n7625 = ~n7623 & ~n7624;
  assign n7626 = ~n7622 & n7625;
  assign n7627 = n1805 & n2979;
  assign n7628 = n7626 & ~n7627;
  assign n7629 = pi29  & ~n7628;
  assign n7630 = pi29  & ~n7629;
  assign n7631 = ~n7628 & ~n7629;
  assign n7632 = ~n7630 & ~n7631;
  assign n7633 = n7621 & ~n7632;
  assign n7634 = n7621 & ~n7633;
  assign n7635 = ~n7632 & ~n7633;
  assign n7636 = ~n7634 & ~n7635;
  assign n7637 = ~n7339 & ~n7343;
  assign n7638 = n7636 & n7637;
  assign n7639 = ~n7636 & ~n7637;
  assign n7640 = ~n7638 & ~n7639;
  assign n7641 = pi87  & n2486;
  assign n7642 = pi85  & n2644;
  assign n7643 = pi86  & n2481;
  assign n7644 = ~n7642 & ~n7643;
  assign n7645 = ~n7641 & n7644;
  assign n7646 = n2252 & n2489;
  assign n7647 = n7645 & ~n7646;
  assign n7648 = pi26  & ~n7647;
  assign n7649 = pi26  & ~n7648;
  assign n7650 = ~n7647 & ~n7648;
  assign n7651 = ~n7649 & ~n7650;
  assign n7652 = n7640 & ~n7651;
  assign n7653 = ~n7640 & n7651;
  assign n7654 = ~n7516 & ~n7653;
  assign n7655 = ~n7652 & n7654;
  assign n7656 = ~n7516 & ~n7655;
  assign n7657 = ~n7652 & ~n7655;
  assign n7658 = ~n7653 & n7657;
  assign n7659 = ~n7656 & ~n7658;
  assign n7660 = pi90  & n2004;
  assign n7661 = pi88  & n2141;
  assign n7662 = pi89  & n1999;
  assign n7663 = ~n7661 & ~n7662;
  assign n7664 = ~n7660 & n7663;
  assign n7665 = n2007 & n2606;
  assign n7666 = n7664 & ~n7665;
  assign n7667 = pi23  & ~n7666;
  assign n7668 = pi23  & ~n7667;
  assign n7669 = ~n7666 & ~n7667;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = n7659 & n7670;
  assign n7672 = ~n7659 & ~n7670;
  assign n7673 = ~n7671 & ~n7672;
  assign n7674 = ~n7515 & n7673;
  assign n7675 = n7515 & ~n7673;
  assign n7676 = ~n7674 & ~n7675;
  assign n7677 = n7514 & ~n7676;
  assign n7678 = ~n7514 & n7676;
  assign n7679 = ~n7677 & ~n7678;
  assign n7680 = ~n7503 & n7679;
  assign n7681 = n7503 & ~n7679;
  assign n7682 = ~n7680 & ~n7681;
  assign n7683 = n7502 & ~n7682;
  assign n7684 = ~n7502 & n7682;
  assign n7685 = ~n7683 & ~n7684;
  assign n7686 = ~n7491 & n7685;
  assign n7687 = n7491 & ~n7685;
  assign n7688 = ~n7686 & ~n7687;
  assign n7689 = pi99  & n918;
  assign n7690 = pi97  & n1031;
  assign n7691 = pi98  & n913;
  assign n7692 = ~n7690 & ~n7691;
  assign n7693 = ~n7689 & n7692;
  assign n7694 = n921 & n4584;
  assign n7695 = n7693 & ~n7694;
  assign n7696 = pi14  & ~n7695;
  assign n7697 = pi14  & ~n7696;
  assign n7698 = ~n7695 & ~n7696;
  assign n7699 = ~n7697 & ~n7698;
  assign n7700 = n7688 & ~n7699;
  assign n7701 = ~n7688 & n7699;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = n7490 & ~n7702;
  assign n7704 = ~n7490 & n7702;
  assign n7705 = ~n7703 & ~n7704;
  assign n7706 = pi102  & n675;
  assign n7707 = pi100  & n769;
  assign n7708 = pi101  & n670;
  assign n7709 = ~n7707 & ~n7708;
  assign n7710 = ~n7706 & n7709;
  assign n7711 = n678 & n5296;
  assign n7712 = n7710 & ~n7711;
  assign n7713 = pi11  & ~n7712;
  assign n7714 = pi11  & ~n7713;
  assign n7715 = ~n7712 & ~n7713;
  assign n7716 = ~n7714 & ~n7715;
  assign n7717 = n7705 & ~n7716;
  assign n7718 = ~n7705 & n7716;
  assign n7719 = ~n7717 & ~n7718;
  assign n7720 = n7489 & ~n7719;
  assign n7721 = ~n7489 & n7719;
  assign n7722 = ~n7720 & ~n7721;
  assign n7723 = pi105  & n493;
  assign n7724 = pi103  & n533;
  assign n7725 = pi104  & n488;
  assign n7726 = ~n7724 & ~n7725;
  assign n7727 = ~n7723 & n7726;
  assign n7728 = n496 & n6065;
  assign n7729 = n7727 & ~n7728;
  assign n7730 = pi8  & ~n7729;
  assign n7731 = pi8  & ~n7730;
  assign n7732 = ~n7729 & ~n7730;
  assign n7733 = ~n7731 & ~n7732;
  assign n7734 = n7722 & ~n7733;
  assign n7735 = ~n7722 & n7733;
  assign n7736 = ~n7443 & ~n7735;
  assign n7737 = ~n7734 & n7736;
  assign n7738 = ~n7443 & ~n7737;
  assign n7739 = ~n7734 & ~n7737;
  assign n7740 = ~n7735 & n7739;
  assign n7741 = ~n7738 & ~n7740;
  assign n7742 = pi108  & n340;
  assign n7743 = pi106  & n380;
  assign n7744 = pi107  & n335;
  assign n7745 = ~n7743 & ~n7744;
  assign n7746 = ~n7742 & n7745;
  assign n7747 = n343 & n6639;
  assign n7748 = n7746 & ~n7747;
  assign n7749 = pi5  & ~n7748;
  assign n7750 = pi5  & ~n7749;
  assign n7751 = ~n7748 & ~n7749;
  assign n7752 = ~n7750 & ~n7751;
  assign n7753 = n7741 & n7752;
  assign n7754 = ~n7741 & ~n7752;
  assign n7755 = ~n7753 & ~n7754;
  assign n7756 = ~n7488 & n7755;
  assign n7757 = n7488 & ~n7755;
  assign n7758 = ~n7756 & ~n7757;
  assign n7759 = pi111  & n264;
  assign n7760 = pi109  & n281;
  assign n7761 = pi110  & n259;
  assign n7762 = ~n7760 & ~n7761;
  assign n7763 = ~n7759 & n7762;
  assign n7764 = ~n7470 & ~n7472;
  assign n7765 = ~pi110  & ~pi111 ;
  assign n7766 = pi110  & pi111 ;
  assign n7767 = ~n7765 & ~n7766;
  assign n7768 = ~n7764 & n7767;
  assign n7769 = n7764 & ~n7767;
  assign n7770 = ~n7768 & ~n7769;
  assign n7771 = n267 & n7770;
  assign n7772 = n7763 & ~n7771;
  assign n7773 = pi2  & ~n7772;
  assign n7774 = pi2  & ~n7773;
  assign n7775 = ~n7772 & ~n7773;
  assign n7776 = ~n7774 & ~n7775;
  assign n7777 = n7758 & ~n7776;
  assign n7778 = ~n7758 & n7776;
  assign n7779 = ~n7777 & ~n7778;
  assign n7780 = ~n7487 & n7779;
  assign n7781 = n7487 & ~n7779;
  assign po47  = ~n7780 & ~n7781;
  assign n7783 = ~n7777 & ~n7780;
  assign n7784 = pi112  & n264;
  assign n7785 = pi110  & n281;
  assign n7786 = pi111  & n259;
  assign n7787 = ~n7785 & ~n7786;
  assign n7788 = ~n7784 & n7787;
  assign n7789 = ~n7766 & ~n7768;
  assign n7790 = ~pi111  & ~pi112 ;
  assign n7791 = pi111  & pi112 ;
  assign n7792 = ~n7790 & ~n7791;
  assign n7793 = ~n7789 & n7792;
  assign n7794 = n7789 & ~n7792;
  assign n7795 = ~n7793 & ~n7794;
  assign n7796 = n267 & n7795;
  assign n7797 = n7788 & ~n7796;
  assign n7798 = pi2  & ~n7797;
  assign n7799 = pi2  & ~n7798;
  assign n7800 = ~n7797 & ~n7798;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = ~n7754 & ~n7756;
  assign n7803 = pi109  & n340;
  assign n7804 = pi107  & n380;
  assign n7805 = pi108  & n335;
  assign n7806 = ~n7804 & ~n7805;
  assign n7807 = ~n7803 & n7806;
  assign n7808 = n343 & n7170;
  assign n7809 = n7807 & ~n7808;
  assign n7810 = pi5  & ~n7809;
  assign n7811 = pi5  & ~n7810;
  assign n7812 = ~n7809 & ~n7810;
  assign n7813 = ~n7811 & ~n7812;
  assign n7814 = ~n7717 & ~n7721;
  assign n7815 = ~n7700 & ~n7704;
  assign n7816 = pi100  & n918;
  assign n7817 = pi98  & n1031;
  assign n7818 = pi99  & n913;
  assign n7819 = ~n7817 & ~n7818;
  assign n7820 = ~n7816 & n7819;
  assign n7821 = n921 & n4808;
  assign n7822 = n7820 & ~n7821;
  assign n7823 = pi14  & ~n7822;
  assign n7824 = pi14  & ~n7823;
  assign n7825 = ~n7822 & ~n7823;
  assign n7826 = ~n7824 & ~n7825;
  assign n7827 = ~n7684 & ~n7686;
  assign n7828 = ~n7678 & ~n7680;
  assign n7829 = pi94  & n1582;
  assign n7830 = pi92  & n1713;
  assign n7831 = pi93  & n1577;
  assign n7832 = ~n7830 & ~n7831;
  assign n7833 = ~n7829 & n7832;
  assign n7834 = n1585 & n3499;
  assign n7835 = n7833 & ~n7834;
  assign n7836 = pi20  & ~n7835;
  assign n7837 = pi20  & ~n7836;
  assign n7838 = ~n7835 & ~n7836;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = ~n7672 & ~n7674;
  assign n7841 = ~n7633 & ~n7639;
  assign n7842 = ~n7610 & ~n7613;
  assign n7843 = pi79  & n4182;
  assign n7844 = pi77  & n4416;
  assign n7845 = pi78  & n4177;
  assign n7846 = ~n7844 & ~n7845;
  assign n7847 = ~n7843 & n7846;
  assign n7848 = n1105 & n4185;
  assign n7849 = n7847 & ~n7848;
  assign n7850 = pi35  & ~n7849;
  assign n7851 = pi35  & ~n7850;
  assign n7852 = ~n7849 & ~n7850;
  assign n7853 = ~n7851 & ~n7852;
  assign n7854 = ~n7594 & ~n7596;
  assign n7855 = pi76  & n4896;
  assign n7856 = pi74  & n5148;
  assign n7857 = pi75  & n4891;
  assign n7858 = ~n7856 & ~n7857;
  assign n7859 = ~n7855 & n7858;
  assign n7860 = n881 & n4899;
  assign n7861 = n7859 & ~n7860;
  assign n7862 = pi38  & ~n7861;
  assign n7863 = pi38  & ~n7862;
  assign n7864 = ~n7861 & ~n7862;
  assign n7865 = ~n7863 & ~n7864;
  assign n7866 = ~n7587 & ~n7590;
  assign n7867 = ~n7581 & ~n7584;
  assign n7868 = pi67  & n7239;
  assign n7869 = pi65  & n7556;
  assign n7870 = pi66  & n7234;
  assign n7871 = ~n7869 & ~n7870;
  assign n7872 = ~n7868 & n7871;
  assign n7873 = n313 & n7242;
  assign n7874 = n7872 & ~n7873;
  assign n7875 = pi47  & ~n7874;
  assign n7876 = pi47  & ~n7875;
  assign n7877 = ~n7874 & ~n7875;
  assign n7878 = ~n7876 & ~n7877;
  assign n7879 = pi47  & ~pi48 ;
  assign n7880 = ~pi47  & pi48 ;
  assign n7881 = ~n7879 & ~n7880;
  assign n7882 = pi64  & ~n7881;
  assign n7883 = n7568 & n7882;
  assign n7884 = ~n7568 & ~n7882;
  assign n7885 = ~n7883 & ~n7884;
  assign n7886 = ~n7878 & n7885;
  assign n7887 = n7878 & ~n7885;
  assign n7888 = ~n7886 & ~n7887;
  assign n7889 = pi70  & n6396;
  assign n7890 = pi68  & n6735;
  assign n7891 = pi69  & n6391;
  assign n7892 = ~n7890 & ~n7891;
  assign n7893 = ~n7889 & n7892;
  assign n7894 = n430 & n6399;
  assign n7895 = n7893 & ~n7894;
  assign n7896 = pi44  & ~n7895;
  assign n7897 = pi44  & ~n7896;
  assign n7898 = ~n7895 & ~n7896;
  assign n7899 = ~n7897 & ~n7898;
  assign n7900 = n7888 & ~n7899;
  assign n7901 = ~n7888 & n7899;
  assign n7902 = ~n7900 & ~n7901;
  assign n7903 = n7867 & ~n7902;
  assign n7904 = ~n7867 & n7902;
  assign n7905 = ~n7903 & ~n7904;
  assign n7906 = pi73  & n5636;
  assign n7907 = pi71  & n5909;
  assign n7908 = pi72  & n5631;
  assign n7909 = ~n7907 & ~n7908;
  assign n7910 = ~n7906 & n7909;
  assign n7911 = n639 & n5639;
  assign n7912 = n7910 & ~n7911;
  assign n7913 = pi41  & ~n7912;
  assign n7914 = pi41  & ~n7913;
  assign n7915 = ~n7912 & ~n7913;
  assign n7916 = ~n7914 & ~n7915;
  assign n7917 = ~n7905 & n7916;
  assign n7918 = n7905 & ~n7916;
  assign n7919 = ~n7917 & ~n7918;
  assign n7920 = ~n7866 & n7919;
  assign n7921 = n7866 & ~n7919;
  assign n7922 = ~n7920 & ~n7921;
  assign n7923 = ~n7865 & n7922;
  assign n7924 = n7865 & ~n7922;
  assign n7925 = ~n7923 & ~n7924;
  assign n7926 = ~n7854 & n7925;
  assign n7927 = n7854 & ~n7925;
  assign n7928 = ~n7926 & ~n7927;
  assign n7929 = ~n7853 & n7928;
  assign n7930 = n7853 & ~n7928;
  assign n7931 = ~n7929 & ~n7930;
  assign n7932 = ~n7842 & n7931;
  assign n7933 = n7842 & ~n7931;
  assign n7934 = ~n7932 & ~n7933;
  assign n7935 = pi82  & n3550;
  assign n7936 = pi80  & n3735;
  assign n7937 = pi81  & n3545;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = ~n7935 & n7938;
  assign n7940 = n1532 & n3553;
  assign n7941 = n7939 & ~n7940;
  assign n7942 = pi32  & ~n7941;
  assign n7943 = pi32  & ~n7942;
  assign n7944 = ~n7941 & ~n7942;
  assign n7945 = ~n7943 & ~n7944;
  assign n7946 = n7934 & ~n7945;
  assign n7947 = n7934 & ~n7946;
  assign n7948 = ~n7945 & ~n7946;
  assign n7949 = ~n7947 & ~n7948;
  assign n7950 = ~n7616 & ~n7619;
  assign n7951 = n7949 & n7950;
  assign n7952 = ~n7949 & ~n7950;
  assign n7953 = ~n7951 & ~n7952;
  assign n7954 = pi85  & n2976;
  assign n7955 = pi83  & n3182;
  assign n7956 = pi84  & n2971;
  assign n7957 = ~n7955 & ~n7956;
  assign n7958 = ~n7954 & n7957;
  assign n7959 = n1943 & n2979;
  assign n7960 = n7958 & ~n7959;
  assign n7961 = pi29  & ~n7960;
  assign n7962 = pi29  & ~n7961;
  assign n7963 = ~n7960 & ~n7961;
  assign n7964 = ~n7962 & ~n7963;
  assign n7965 = n7953 & ~n7964;
  assign n7966 = ~n7953 & n7964;
  assign n7967 = ~n7965 & ~n7966;
  assign n7968 = n7841 & ~n7967;
  assign n7969 = ~n7841 & n7967;
  assign n7970 = ~n7968 & ~n7969;
  assign n7971 = pi88  & n2486;
  assign n7972 = pi86  & n2644;
  assign n7973 = pi87  & n2481;
  assign n7974 = ~n7972 & ~n7973;
  assign n7975 = ~n7971 & n7974;
  assign n7976 = n2277 & n2489;
  assign n7977 = n7975 & ~n7976;
  assign n7978 = pi26  & ~n7977;
  assign n7979 = pi26  & ~n7978;
  assign n7980 = ~n7977 & ~n7978;
  assign n7981 = ~n7979 & ~n7980;
  assign n7982 = ~n7970 & n7981;
  assign n7983 = n7970 & ~n7981;
  assign n7984 = ~n7982 & ~n7983;
  assign n7985 = ~n7657 & n7984;
  assign n7986 = n7657 & ~n7984;
  assign n7987 = ~n7985 & ~n7986;
  assign n7988 = pi91  & n2004;
  assign n7989 = pi89  & n2141;
  assign n7990 = pi90  & n1999;
  assign n7991 = ~n7989 & ~n7990;
  assign n7992 = ~n7988 & n7991;
  assign n7993 = n2007 & n2926;
  assign n7994 = n7992 & ~n7993;
  assign n7995 = pi23  & ~n7994;
  assign n7996 = pi23  & ~n7995;
  assign n7997 = ~n7994 & ~n7995;
  assign n7998 = ~n7996 & ~n7997;
  assign n7999 = n7987 & ~n7998;
  assign n8000 = ~n7987 & n7998;
  assign n8001 = ~n7999 & ~n8000;
  assign n8002 = ~n7840 & n8001;
  assign n8003 = n7840 & ~n8001;
  assign n8004 = ~n8002 & ~n8003;
  assign n8005 = ~n7839 & n8004;
  assign n8006 = n7839 & ~n8004;
  assign n8007 = ~n8005 & ~n8006;
  assign n8008 = ~n7828 & n8007;
  assign n8009 = n7828 & ~n8007;
  assign n8010 = ~n8008 & ~n8009;
  assign n8011 = pi97  & n1269;
  assign n8012 = pi95  & n1340;
  assign n8013 = pi96  & n1264;
  assign n8014 = ~n8012 & ~n8013;
  assign n8015 = ~n8011 & n8014;
  assign n8016 = n1272 & n3946;
  assign n8017 = n8015 & ~n8016;
  assign n8018 = pi17  & ~n8017;
  assign n8019 = pi17  & ~n8018;
  assign n8020 = ~n8017 & ~n8018;
  assign n8021 = ~n8019 & ~n8020;
  assign n8022 = n8010 & ~n8021;
  assign n8023 = ~n8010 & n8021;
  assign n8024 = ~n8022 & ~n8023;
  assign n8025 = ~n7827 & n8024;
  assign n8026 = n7827 & ~n8024;
  assign n8027 = ~n8025 & ~n8026;
  assign n8028 = ~n7826 & n8027;
  assign n8029 = n7826 & ~n8027;
  assign n8030 = ~n8028 & ~n8029;
  assign n8031 = n7815 & ~n8030;
  assign n8032 = ~n7815 & n8030;
  assign n8033 = ~n8031 & ~n8032;
  assign n8034 = pi103  & n675;
  assign n8035 = pi101  & n769;
  assign n8036 = pi102  & n670;
  assign n8037 = ~n8035 & ~n8036;
  assign n8038 = ~n8034 & n8037;
  assign n8039 = n678 & n5540;
  assign n8040 = n8038 & ~n8039;
  assign n8041 = pi11  & ~n8040;
  assign n8042 = pi11  & ~n8041;
  assign n8043 = ~n8040 & ~n8041;
  assign n8044 = ~n8042 & ~n8043;
  assign n8045 = n8033 & ~n8044;
  assign n8046 = ~n8033 & n8044;
  assign n8047 = ~n8045 & ~n8046;
  assign n8048 = n7814 & ~n8047;
  assign n8049 = ~n7814 & n8047;
  assign n8050 = ~n8048 & ~n8049;
  assign n8051 = pi106  & n493;
  assign n8052 = pi104  & n533;
  assign n8053 = pi105  & n488;
  assign n8054 = ~n8052 & ~n8053;
  assign n8055 = ~n8051 & n8054;
  assign n8056 = n496 & n6090;
  assign n8057 = n8055 & ~n8056;
  assign n8058 = pi8  & ~n8057;
  assign n8059 = pi8  & ~n8058;
  assign n8060 = ~n8057 & ~n8058;
  assign n8061 = ~n8059 & ~n8060;
  assign n8062 = n8050 & ~n8061;
  assign n8063 = ~n8050 & n8061;
  assign n8064 = ~n8062 & ~n8063;
  assign n8065 = ~n7739 & n8064;
  assign n8066 = n7739 & ~n8064;
  assign n8067 = ~n8065 & ~n8066;
  assign n8068 = ~n7813 & n8067;
  assign n8069 = n7813 & ~n8067;
  assign n8070 = ~n8068 & ~n8069;
  assign n8071 = ~n7802 & n8070;
  assign n8072 = n7802 & ~n8070;
  assign n8073 = ~n8071 & ~n8072;
  assign n8074 = n7801 & ~n8073;
  assign n8075 = ~n7801 & n8073;
  assign n8076 = ~n8074 & ~n8075;
  assign n8077 = ~n7783 & n8076;
  assign n8078 = n7783 & ~n8076;
  assign po48  = ~n8077 & ~n8078;
  assign n8080 = ~n8075 & ~n8077;
  assign n8081 = ~n8068 & ~n8071;
  assign n8082 = ~n8062 & ~n8065;
  assign n8083 = ~n8045 & ~n8049;
  assign n8084 = ~n8028 & ~n8032;
  assign n8085 = ~n8022 & ~n8025;
  assign n8086 = ~n8005 & ~n8008;
  assign n8087 = pi95  & n1582;
  assign n8088 = pi93  & n1713;
  assign n8089 = pi94  & n1577;
  assign n8090 = ~n8088 & ~n8089;
  assign n8091 = ~n8087 & n8090;
  assign n8092 = n1585 & n3710;
  assign n8093 = n8091 & ~n8092;
  assign n8094 = pi20  & ~n8093;
  assign n8095 = pi20  & ~n8094;
  assign n8096 = ~n8093 & ~n8094;
  assign n8097 = ~n8095 & ~n8096;
  assign n8098 = ~n7999 & ~n8002;
  assign n8099 = pi92  & n2004;
  assign n8100 = pi90  & n2141;
  assign n8101 = pi91  & n1999;
  assign n8102 = ~n8100 & ~n8101;
  assign n8103 = ~n8099 & n8102;
  assign n8104 = n2007 & n3119;
  assign n8105 = n8103 & ~n8104;
  assign n8106 = pi23  & ~n8105;
  assign n8107 = pi23  & ~n8106;
  assign n8108 = ~n8105 & ~n8106;
  assign n8109 = ~n8107 & ~n8108;
  assign n8110 = ~n7983 & ~n7985;
  assign n8111 = ~n7946 & ~n7952;
  assign n8112 = ~n7929 & ~n7932;
  assign n8113 = ~n7923 & ~n7926;
  assign n8114 = ~n7918 & ~n7920;
  assign n8115 = ~n7900 & ~n7904;
  assign n8116 = ~n7883 & ~n7886;
  assign n8117 = pi68  & n7239;
  assign n8118 = pi66  & n7556;
  assign n8119 = pi67  & n7234;
  assign n8120 = ~n8118 & ~n8119;
  assign n8121 = ~n8117 & n8120;
  assign n8122 = n364 & n7242;
  assign n8123 = n8121 & ~n8122;
  assign n8124 = pi47  & ~n8123;
  assign n8125 = pi47  & ~n8124;
  assign n8126 = ~n8123 & ~n8124;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = pi50  & ~n7882;
  assign n8129 = ~pi48  & pi49 ;
  assign n8130 = pi48  & ~pi49 ;
  assign n8131 = ~n8129 & ~n8130;
  assign n8132 = n7881 & ~n8131;
  assign n8133 = pi64  & n8132;
  assign n8134 = ~pi49  & pi50 ;
  assign n8135 = pi49  & ~pi50 ;
  assign n8136 = ~n8134 & ~n8135;
  assign n8137 = ~n7881 & n8136;
  assign n8138 = pi65  & n8137;
  assign n8139 = ~n8133 & ~n8138;
  assign n8140 = ~n7881 & ~n8136;
  assign n8141 = n270 & n8140;
  assign n8142 = n8139 & ~n8141;
  assign n8143 = pi50  & ~n8142;
  assign n8144 = pi50  & ~n8143;
  assign n8145 = ~n8142 & ~n8143;
  assign n8146 = ~n8144 & ~n8145;
  assign n8147 = n8128 & ~n8146;
  assign n8148 = ~n8128 & n8146;
  assign n8149 = ~n8147 & ~n8148;
  assign n8150 = n8127 & ~n8149;
  assign n8151 = ~n8127 & n8149;
  assign n8152 = ~n8150 & ~n8151;
  assign n8153 = ~n8116 & n8152;
  assign n8154 = n8116 & ~n8152;
  assign n8155 = ~n8153 & ~n8154;
  assign n8156 = pi71  & n6396;
  assign n8157 = pi69  & n6735;
  assign n8158 = pi70  & n6391;
  assign n8159 = ~n8157 & ~n8158;
  assign n8160 = ~n8156 & n8159;
  assign n8161 = n476 & n6399;
  assign n8162 = n8160 & ~n8161;
  assign n8163 = pi44  & ~n8162;
  assign n8164 = pi44  & ~n8163;
  assign n8165 = ~n8162 & ~n8163;
  assign n8166 = ~n8164 & ~n8165;
  assign n8167 = n8155 & ~n8166;
  assign n8168 = ~n8155 & n8166;
  assign n8169 = ~n8167 & ~n8168;
  assign n8170 = n8115 & ~n8169;
  assign n8171 = ~n8115 & n8169;
  assign n8172 = ~n8170 & ~n8171;
  assign n8173 = pi74  & n5636;
  assign n8174 = pi72  & n5909;
  assign n8175 = pi73  & n5631;
  assign n8176 = ~n8174 & ~n8175;
  assign n8177 = ~n8173 & n8176;
  assign n8178 = n722 & n5639;
  assign n8179 = n8177 & ~n8178;
  assign n8180 = pi41  & ~n8179;
  assign n8181 = pi41  & ~n8180;
  assign n8182 = ~n8179 & ~n8180;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = n8172 & ~n8183;
  assign n8185 = ~n8172 & n8183;
  assign n8186 = ~n8114 & ~n8185;
  assign n8187 = ~n8184 & n8186;
  assign n8188 = ~n8114 & ~n8187;
  assign n8189 = ~n8184 & ~n8187;
  assign n8190 = ~n8185 & n8189;
  assign n8191 = ~n8188 & ~n8190;
  assign n8192 = pi77  & n4896;
  assign n8193 = pi75  & n5148;
  assign n8194 = pi76  & n4891;
  assign n8195 = ~n8193 & ~n8194;
  assign n8196 = ~n8192 & n8195;
  assign n8197 = n984 & n4899;
  assign n8198 = n8196 & ~n8197;
  assign n8199 = pi38  & ~n8198;
  assign n8200 = pi38  & ~n8199;
  assign n8201 = ~n8198 & ~n8199;
  assign n8202 = ~n8200 & ~n8201;
  assign n8203 = n8191 & n8202;
  assign n8204 = ~n8191 & ~n8202;
  assign n8205 = ~n8203 & ~n8204;
  assign n8206 = ~n8113 & n8205;
  assign n8207 = n8113 & ~n8205;
  assign n8208 = ~n8206 & ~n8207;
  assign n8209 = pi80  & n4182;
  assign n8210 = pi78  & n4416;
  assign n8211 = pi79  & n4177;
  assign n8212 = ~n8210 & ~n8211;
  assign n8213 = ~n8209 & n8212;
  assign n8214 = n1205 & n4185;
  assign n8215 = n8213 & ~n8214;
  assign n8216 = pi35  & ~n8215;
  assign n8217 = pi35  & ~n8216;
  assign n8218 = ~n8215 & ~n8216;
  assign n8219 = ~n8217 & ~n8218;
  assign n8220 = n8208 & ~n8219;
  assign n8221 = ~n8208 & n8219;
  assign n8222 = ~n8220 & ~n8221;
  assign n8223 = n8112 & ~n8222;
  assign n8224 = ~n8112 & n8222;
  assign n8225 = ~n8223 & ~n8224;
  assign n8226 = pi83  & n3550;
  assign n8227 = pi81  & n3735;
  assign n8228 = pi82  & n3545;
  assign n8229 = ~n8227 & ~n8228;
  assign n8230 = ~n8226 & n8229;
  assign n8231 = n1672 & n3553;
  assign n8232 = n8230 & ~n8231;
  assign n8233 = pi32  & ~n8232;
  assign n8234 = pi32  & ~n8233;
  assign n8235 = ~n8232 & ~n8233;
  assign n8236 = ~n8234 & ~n8235;
  assign n8237 = n8225 & ~n8236;
  assign n8238 = ~n8225 & n8236;
  assign n8239 = ~n8237 & ~n8238;
  assign n8240 = n8111 & ~n8239;
  assign n8241 = ~n8111 & n8239;
  assign n8242 = ~n8240 & ~n8241;
  assign n8243 = pi86  & n2976;
  assign n8244 = pi84  & n3182;
  assign n8245 = pi85  & n2971;
  assign n8246 = ~n8244 & ~n8245;
  assign n8247 = ~n8243 & n8246;
  assign n8248 = n2099 & n2979;
  assign n8249 = n8247 & ~n8248;
  assign n8250 = pi29  & ~n8249;
  assign n8251 = pi29  & ~n8250;
  assign n8252 = ~n8249 & ~n8250;
  assign n8253 = ~n8251 & ~n8252;
  assign n8254 = n8242 & ~n8253;
  assign n8255 = n8242 & ~n8254;
  assign n8256 = ~n8253 & ~n8254;
  assign n8257 = ~n8255 & ~n8256;
  assign n8258 = ~n7965 & ~n7969;
  assign n8259 = n8257 & n8258;
  assign n8260 = ~n8257 & ~n8258;
  assign n8261 = ~n8259 & ~n8260;
  assign n8262 = pi89  & n2486;
  assign n8263 = pi87  & n2644;
  assign n8264 = pi88  & n2481;
  assign n8265 = ~n8263 & ~n8264;
  assign n8266 = ~n8262 & n8265;
  assign n8267 = n2432 & n2489;
  assign n8268 = n8266 & ~n8267;
  assign n8269 = pi26  & ~n8268;
  assign n8270 = pi26  & ~n8269;
  assign n8271 = ~n8268 & ~n8269;
  assign n8272 = ~n8270 & ~n8271;
  assign n8273 = n8261 & ~n8272;
  assign n8274 = ~n8261 & n8272;
  assign n8275 = ~n8273 & ~n8274;
  assign n8276 = ~n8110 & n8275;
  assign n8277 = n8110 & ~n8275;
  assign n8278 = ~n8276 & ~n8277;
  assign n8279 = ~n8109 & n8278;
  assign n8280 = n8109 & ~n8278;
  assign n8281 = ~n8279 & ~n8280;
  assign n8282 = ~n8098 & n8281;
  assign n8283 = n8098 & ~n8281;
  assign n8284 = ~n8282 & ~n8283;
  assign n8285 = ~n8097 & n8284;
  assign n8286 = n8097 & ~n8284;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = n8086 & ~n8287;
  assign n8289 = ~n8086 & n8287;
  assign n8290 = ~n8288 & ~n8289;
  assign n8291 = pi98  & n1269;
  assign n8292 = pi96  & n1340;
  assign n8293 = pi97  & n1264;
  assign n8294 = ~n8292 & ~n8293;
  assign n8295 = ~n8291 & n8294;
  assign n8296 = n1272 & n4360;
  assign n8297 = n8295 & ~n8296;
  assign n8298 = pi17  & ~n8297;
  assign n8299 = pi17  & ~n8298;
  assign n8300 = ~n8297 & ~n8298;
  assign n8301 = ~n8299 & ~n8300;
  assign n8302 = n8290 & ~n8301;
  assign n8303 = ~n8290 & n8301;
  assign n8304 = ~n8302 & ~n8303;
  assign n8305 = n8085 & ~n8304;
  assign n8306 = ~n8085 & n8304;
  assign n8307 = ~n8305 & ~n8306;
  assign n8308 = pi101  & n918;
  assign n8309 = pi99  & n1031;
  assign n8310 = pi100  & n913;
  assign n8311 = ~n8309 & ~n8310;
  assign n8312 = ~n8308 & n8311;
  assign n8313 = n921 & n5056;
  assign n8314 = n8312 & ~n8313;
  assign n8315 = pi14  & ~n8314;
  assign n8316 = pi14  & ~n8315;
  assign n8317 = ~n8314 & ~n8315;
  assign n8318 = ~n8316 & ~n8317;
  assign n8319 = n8307 & ~n8318;
  assign n8320 = ~n8307 & n8318;
  assign n8321 = ~n8319 & ~n8320;
  assign n8322 = n8084 & ~n8321;
  assign n8323 = ~n8084 & n8321;
  assign n8324 = ~n8322 & ~n8323;
  assign n8325 = pi104  & n675;
  assign n8326 = pi102  & n769;
  assign n8327 = pi103  & n670;
  assign n8328 = ~n8326 & ~n8327;
  assign n8329 = ~n8325 & n8328;
  assign n8330 = n678 & n5565;
  assign n8331 = n8329 & ~n8330;
  assign n8332 = pi11  & ~n8331;
  assign n8333 = pi11  & ~n8332;
  assign n8334 = ~n8331 & ~n8332;
  assign n8335 = ~n8333 & ~n8334;
  assign n8336 = n8324 & ~n8335;
  assign n8337 = ~n8324 & n8335;
  assign n8338 = ~n8336 & ~n8337;
  assign n8339 = n8083 & ~n8338;
  assign n8340 = ~n8083 & n8338;
  assign n8341 = ~n8339 & ~n8340;
  assign n8342 = pi107  & n493;
  assign n8343 = pi105  & n533;
  assign n8344 = pi106  & n488;
  assign n8345 = ~n8343 & ~n8344;
  assign n8346 = ~n8342 & n8345;
  assign n8347 = n496 & n6614;
  assign n8348 = n8346 & ~n8347;
  assign n8349 = pi8  & ~n8348;
  assign n8350 = pi8  & ~n8349;
  assign n8351 = ~n8348 & ~n8349;
  assign n8352 = ~n8350 & ~n8351;
  assign n8353 = n8341 & ~n8352;
  assign n8354 = ~n8341 & n8352;
  assign n8355 = ~n8353 & ~n8354;
  assign n8356 = n8082 & ~n8355;
  assign n8357 = ~n8082 & n8355;
  assign n8358 = ~n8356 & ~n8357;
  assign n8359 = pi110  & n340;
  assign n8360 = pi108  & n380;
  assign n8361 = pi109  & n335;
  assign n8362 = ~n8360 & ~n8361;
  assign n8363 = ~n8359 & n8362;
  assign n8364 = n343 & n7474;
  assign n8365 = n8363 & ~n8364;
  assign n8366 = pi5  & ~n8365;
  assign n8367 = pi5  & ~n8366;
  assign n8368 = ~n8365 & ~n8366;
  assign n8369 = ~n8367 & ~n8368;
  assign n8370 = n8358 & ~n8369;
  assign n8371 = ~n8358 & n8369;
  assign n8372 = ~n8370 & ~n8371;
  assign n8373 = n8081 & ~n8372;
  assign n8374 = ~n8081 & n8372;
  assign n8375 = ~n8373 & ~n8374;
  assign n8376 = pi113  & n264;
  assign n8377 = pi111  & n281;
  assign n8378 = pi112  & n259;
  assign n8379 = ~n8377 & ~n8378;
  assign n8380 = ~n8376 & n8379;
  assign n8381 = ~n7791 & ~n7793;
  assign n8382 = ~pi112  & ~pi113 ;
  assign n8383 = pi112  & pi113 ;
  assign n8384 = ~n8382 & ~n8383;
  assign n8385 = ~n8381 & n8384;
  assign n8386 = n8381 & ~n8384;
  assign n8387 = ~n8385 & ~n8386;
  assign n8388 = n267 & n8387;
  assign n8389 = n8380 & ~n8388;
  assign n8390 = pi2  & ~n8389;
  assign n8391 = pi2  & ~n8390;
  assign n8392 = ~n8389 & ~n8390;
  assign n8393 = ~n8391 & ~n8392;
  assign n8394 = ~n8375 & n8393;
  assign n8395 = n8375 & ~n8393;
  assign n8396 = ~n8394 & ~n8395;
  assign n8397 = ~n8080 & n8396;
  assign n8398 = n8080 & ~n8396;
  assign po49  = ~n8397 & ~n8398;
  assign n8400 = ~n8395 & ~n8397;
  assign n8401 = ~n8370 & ~n8374;
  assign n8402 = ~n8353 & ~n8357;
  assign n8403 = ~n8336 & ~n8340;
  assign n8404 = ~n8319 & ~n8323;
  assign n8405 = ~n8302 & ~n8306;
  assign n8406 = ~n8285 & ~n8289;
  assign n8407 = pi96  & n1582;
  assign n8408 = pi94  & n1713;
  assign n8409 = pi95  & n1577;
  assign n8410 = ~n8408 & ~n8409;
  assign n8411 = ~n8407 & n8410;
  assign n8412 = n1585 & n3921;
  assign n8413 = n8411 & ~n8412;
  assign n8414 = pi20  & ~n8413;
  assign n8415 = pi20  & ~n8414;
  assign n8416 = ~n8413 & ~n8414;
  assign n8417 = ~n8415 & ~n8416;
  assign n8418 = ~n8279 & ~n8282;
  assign n8419 = pi93  & n2004;
  assign n8420 = pi91  & n2141;
  assign n8421 = pi92  & n1999;
  assign n8422 = ~n8420 & ~n8421;
  assign n8423 = ~n8419 & n8422;
  assign n8424 = n2007 & n3144;
  assign n8425 = n8423 & ~n8424;
  assign n8426 = pi23  & ~n8425;
  assign n8427 = pi23  & ~n8426;
  assign n8428 = ~n8425 & ~n8426;
  assign n8429 = ~n8427 & ~n8428;
  assign n8430 = ~n8273 & ~n8276;
  assign n8431 = ~n8254 & ~n8260;
  assign n8432 = ~n8220 & ~n8224;
  assign n8433 = pi81  & n4182;
  assign n8434 = pi79  & n4416;
  assign n8435 = pi80  & n4177;
  assign n8436 = ~n8434 & ~n8435;
  assign n8437 = ~n8433 & n8436;
  assign n8438 = n1413 & n4185;
  assign n8439 = n8437 & ~n8438;
  assign n8440 = pi35  & ~n8439;
  assign n8441 = pi35  & ~n8440;
  assign n8442 = ~n8439 & ~n8440;
  assign n8443 = ~n8441 & ~n8442;
  assign n8444 = ~n8204 & ~n8206;
  assign n8445 = pi75  & n5636;
  assign n8446 = pi73  & n5909;
  assign n8447 = pi74  & n5631;
  assign n8448 = ~n8446 & ~n8447;
  assign n8449 = ~n8445 & n8448;
  assign n8450 = n747 & n5639;
  assign n8451 = n8449 & ~n8450;
  assign n8452 = pi41  & ~n8451;
  assign n8453 = pi41  & ~n8452;
  assign n8454 = ~n8451 & ~n8452;
  assign n8455 = ~n8453 & ~n8454;
  assign n8456 = ~n8167 & ~n8171;
  assign n8457 = pi72  & n6396;
  assign n8458 = pi70  & n6735;
  assign n8459 = pi71  & n6391;
  assign n8460 = ~n8458 & ~n8459;
  assign n8461 = ~n8457 & n8460;
  assign n8462 = n575 & n6399;
  assign n8463 = n8461 & ~n8462;
  assign n8464 = pi44  & ~n8463;
  assign n8465 = pi44  & ~n8464;
  assign n8466 = ~n8463 & ~n8464;
  assign n8467 = ~n8465 & ~n8466;
  assign n8468 = ~n8151 & ~n8153;
  assign n8469 = pi66  & n8137;
  assign n8470 = n7881 & ~n8136;
  assign n8471 = n8131 & n8470;
  assign n8472 = pi64  & n8471;
  assign n8473 = pi65  & n8132;
  assign n8474 = ~n8472 & ~n8473;
  assign n8475 = ~n8469 & n8474;
  assign n8476 = n291 & n8140;
  assign n8477 = n8475 & ~n8476;
  assign n8478 = pi50  & ~n8477;
  assign n8479 = pi50  & ~n8478;
  assign n8480 = ~n8477 & ~n8478;
  assign n8481 = ~n8479 & ~n8480;
  assign n8482 = ~n8147 & n8481;
  assign n8483 = n8147 & ~n8481;
  assign n8484 = ~n8482 & ~n8483;
  assign n8485 = pi69  & n7239;
  assign n8486 = pi67  & n7556;
  assign n8487 = pi68  & n7234;
  assign n8488 = ~n8486 & ~n8487;
  assign n8489 = ~n8485 & n8488;
  assign n8490 = n405 & n7242;
  assign n8491 = n8489 & ~n8490;
  assign n8492 = pi47  & ~n8491;
  assign n8493 = pi47  & ~n8492;
  assign n8494 = ~n8491 & ~n8492;
  assign n8495 = ~n8493 & ~n8494;
  assign n8496 = n8484 & ~n8495;
  assign n8497 = ~n8484 & n8495;
  assign n8498 = ~n8496 & ~n8497;
  assign n8499 = ~n8468 & n8498;
  assign n8500 = n8468 & ~n8498;
  assign n8501 = ~n8499 & ~n8500;
  assign n8502 = ~n8467 & n8501;
  assign n8503 = n8467 & ~n8501;
  assign n8504 = ~n8502 & ~n8503;
  assign n8505 = ~n8456 & n8504;
  assign n8506 = n8456 & ~n8504;
  assign n8507 = ~n8505 & ~n8506;
  assign n8508 = n8455 & ~n8507;
  assign n8509 = ~n8455 & n8507;
  assign n8510 = ~n8508 & ~n8509;
  assign n8511 = ~n8189 & n8510;
  assign n8512 = n8189 & ~n8510;
  assign n8513 = ~n8511 & ~n8512;
  assign n8514 = pi78  & n4896;
  assign n8515 = pi76  & n5148;
  assign n8516 = pi77  & n4891;
  assign n8517 = ~n8515 & ~n8516;
  assign n8518 = ~n8514 & n8517;
  assign n8519 = n1009 & n4899;
  assign n8520 = n8518 & ~n8519;
  assign n8521 = pi38  & ~n8520;
  assign n8522 = pi38  & ~n8521;
  assign n8523 = ~n8520 & ~n8521;
  assign n8524 = ~n8522 & ~n8523;
  assign n8525 = n8513 & ~n8524;
  assign n8526 = ~n8513 & n8524;
  assign n8527 = ~n8525 & ~n8526;
  assign n8528 = ~n8444 & n8527;
  assign n8529 = n8444 & ~n8527;
  assign n8530 = ~n8528 & ~n8529;
  assign n8531 = ~n8443 & n8530;
  assign n8532 = n8443 & ~n8530;
  assign n8533 = ~n8531 & ~n8532;
  assign n8534 = ~n8432 & n8533;
  assign n8535 = n8432 & ~n8533;
  assign n8536 = ~n8534 & ~n8535;
  assign n8537 = pi84  & n3550;
  assign n8538 = pi82  & n3735;
  assign n8539 = pi83  & n3545;
  assign n8540 = ~n8538 & ~n8539;
  assign n8541 = ~n8537 & n8540;
  assign n8542 = n1805 & n3553;
  assign n8543 = n8541 & ~n8542;
  assign n8544 = pi32  & ~n8543;
  assign n8545 = pi32  & ~n8544;
  assign n8546 = ~n8543 & ~n8544;
  assign n8547 = ~n8545 & ~n8546;
  assign n8548 = n8536 & ~n8547;
  assign n8549 = n8536 & ~n8548;
  assign n8550 = ~n8547 & ~n8548;
  assign n8551 = ~n8549 & ~n8550;
  assign n8552 = ~n8237 & ~n8241;
  assign n8553 = n8551 & n8552;
  assign n8554 = ~n8551 & ~n8552;
  assign n8555 = ~n8553 & ~n8554;
  assign n8556 = pi87  & n2976;
  assign n8557 = pi85  & n3182;
  assign n8558 = pi86  & n2971;
  assign n8559 = ~n8557 & ~n8558;
  assign n8560 = ~n8556 & n8559;
  assign n8561 = n2252 & n2979;
  assign n8562 = n8560 & ~n8561;
  assign n8563 = pi29  & ~n8562;
  assign n8564 = pi29  & ~n8563;
  assign n8565 = ~n8562 & ~n8563;
  assign n8566 = ~n8564 & ~n8565;
  assign n8567 = n8555 & ~n8566;
  assign n8568 = ~n8555 & n8566;
  assign n8569 = ~n8431 & ~n8568;
  assign n8570 = ~n8567 & n8569;
  assign n8571 = ~n8431 & ~n8570;
  assign n8572 = ~n8567 & ~n8570;
  assign n8573 = ~n8568 & n8572;
  assign n8574 = ~n8571 & ~n8573;
  assign n8575 = pi90  & n2486;
  assign n8576 = pi88  & n2644;
  assign n8577 = pi89  & n2481;
  assign n8578 = ~n8576 & ~n8577;
  assign n8579 = ~n8575 & n8578;
  assign n8580 = n2489 & n2606;
  assign n8581 = n8579 & ~n8580;
  assign n8582 = pi26  & ~n8581;
  assign n8583 = pi26  & ~n8582;
  assign n8584 = ~n8581 & ~n8582;
  assign n8585 = ~n8583 & ~n8584;
  assign n8586 = n8574 & n8585;
  assign n8587 = ~n8574 & ~n8585;
  assign n8588 = ~n8586 & ~n8587;
  assign n8589 = ~n8430 & n8588;
  assign n8590 = n8430 & ~n8588;
  assign n8591 = ~n8589 & ~n8590;
  assign n8592 = n8429 & ~n8591;
  assign n8593 = ~n8429 & n8591;
  assign n8594 = ~n8592 & ~n8593;
  assign n8595 = ~n8418 & n8594;
  assign n8596 = n8418 & ~n8594;
  assign n8597 = ~n8595 & ~n8596;
  assign n8598 = n8417 & ~n8597;
  assign n8599 = ~n8417 & n8597;
  assign n8600 = ~n8598 & ~n8599;
  assign n8601 = ~n8406 & n8600;
  assign n8602 = n8406 & ~n8600;
  assign n8603 = ~n8601 & ~n8602;
  assign n8604 = pi99  & n1269;
  assign n8605 = pi97  & n1340;
  assign n8606 = pi98  & n1264;
  assign n8607 = ~n8605 & ~n8606;
  assign n8608 = ~n8604 & n8607;
  assign n8609 = n1272 & n4584;
  assign n8610 = n8608 & ~n8609;
  assign n8611 = pi17  & ~n8610;
  assign n8612 = pi17  & ~n8611;
  assign n8613 = ~n8610 & ~n8611;
  assign n8614 = ~n8612 & ~n8613;
  assign n8615 = n8603 & ~n8614;
  assign n8616 = ~n8603 & n8614;
  assign n8617 = ~n8615 & ~n8616;
  assign n8618 = n8405 & ~n8617;
  assign n8619 = ~n8405 & n8617;
  assign n8620 = ~n8618 & ~n8619;
  assign n8621 = pi102  & n918;
  assign n8622 = pi100  & n1031;
  assign n8623 = pi101  & n913;
  assign n8624 = ~n8622 & ~n8623;
  assign n8625 = ~n8621 & n8624;
  assign n8626 = n921 & n5296;
  assign n8627 = n8625 & ~n8626;
  assign n8628 = pi14  & ~n8627;
  assign n8629 = pi14  & ~n8628;
  assign n8630 = ~n8627 & ~n8628;
  assign n8631 = ~n8629 & ~n8630;
  assign n8632 = n8620 & ~n8631;
  assign n8633 = ~n8620 & n8631;
  assign n8634 = ~n8632 & ~n8633;
  assign n8635 = n8404 & ~n8634;
  assign n8636 = ~n8404 & n8634;
  assign n8637 = ~n8635 & ~n8636;
  assign n8638 = pi105  & n675;
  assign n8639 = pi103  & n769;
  assign n8640 = pi104  & n670;
  assign n8641 = ~n8639 & ~n8640;
  assign n8642 = ~n8638 & n8641;
  assign n8643 = n678 & n6065;
  assign n8644 = n8642 & ~n8643;
  assign n8645 = pi11  & ~n8644;
  assign n8646 = pi11  & ~n8645;
  assign n8647 = ~n8644 & ~n8645;
  assign n8648 = ~n8646 & ~n8647;
  assign n8649 = n8637 & ~n8648;
  assign n8650 = ~n8637 & n8648;
  assign n8651 = ~n8649 & ~n8650;
  assign n8652 = n8403 & ~n8651;
  assign n8653 = ~n8403 & n8651;
  assign n8654 = ~n8652 & ~n8653;
  assign n8655 = pi108  & n493;
  assign n8656 = pi106  & n533;
  assign n8657 = pi107  & n488;
  assign n8658 = ~n8656 & ~n8657;
  assign n8659 = ~n8655 & n8658;
  assign n8660 = n496 & n6639;
  assign n8661 = n8659 & ~n8660;
  assign n8662 = pi8  & ~n8661;
  assign n8663 = pi8  & ~n8662;
  assign n8664 = ~n8661 & ~n8662;
  assign n8665 = ~n8663 & ~n8664;
  assign n8666 = n8654 & ~n8665;
  assign n8667 = ~n8654 & n8665;
  assign n8668 = ~n8402 & ~n8667;
  assign n8669 = ~n8666 & n8668;
  assign n8670 = ~n8402 & ~n8669;
  assign n8671 = ~n8666 & ~n8669;
  assign n8672 = ~n8667 & n8671;
  assign n8673 = ~n8670 & ~n8672;
  assign n8674 = pi111  & n340;
  assign n8675 = pi109  & n380;
  assign n8676 = pi110  & n335;
  assign n8677 = ~n8675 & ~n8676;
  assign n8678 = ~n8674 & n8677;
  assign n8679 = n343 & n7770;
  assign n8680 = n8678 & ~n8679;
  assign n8681 = pi5  & ~n8680;
  assign n8682 = pi5  & ~n8681;
  assign n8683 = ~n8680 & ~n8681;
  assign n8684 = ~n8682 & ~n8683;
  assign n8685 = ~n8673 & ~n8684;
  assign n8686 = n8673 & n8684;
  assign n8687 = ~n8685 & ~n8686;
  assign n8688 = n8401 & ~n8687;
  assign n8689 = ~n8401 & n8687;
  assign n8690 = ~n8688 & ~n8689;
  assign n8691 = pi114  & n264;
  assign n8692 = pi112  & n281;
  assign n8693 = pi113  & n259;
  assign n8694 = ~n8692 & ~n8693;
  assign n8695 = ~n8691 & n8694;
  assign n8696 = ~n8383 & ~n8385;
  assign n8697 = ~pi113  & ~pi114 ;
  assign n8698 = pi113  & pi114 ;
  assign n8699 = ~n8697 & ~n8698;
  assign n8700 = ~n8696 & n8699;
  assign n8701 = n8696 & ~n8699;
  assign n8702 = ~n8700 & ~n8701;
  assign n8703 = n267 & n8702;
  assign n8704 = n8695 & ~n8703;
  assign n8705 = pi2  & ~n8704;
  assign n8706 = pi2  & ~n8705;
  assign n8707 = ~n8704 & ~n8705;
  assign n8708 = ~n8706 & ~n8707;
  assign n8709 = n8690 & ~n8708;
  assign n8710 = ~n8690 & n8708;
  assign n8711 = ~n8709 & ~n8710;
  assign n8712 = ~n8400 & n8711;
  assign n8713 = n8400 & ~n8711;
  assign po50  = ~n8712 & ~n8713;
  assign n8715 = ~n8709 & ~n8712;
  assign n8716 = pi115  & n264;
  assign n8717 = pi113  & n281;
  assign n8718 = pi114  & n259;
  assign n8719 = ~n8717 & ~n8718;
  assign n8720 = ~n8716 & n8719;
  assign n8721 = ~n8698 & ~n8700;
  assign n8722 = ~pi114  & ~pi115 ;
  assign n8723 = pi114  & pi115 ;
  assign n8724 = ~n8722 & ~n8723;
  assign n8725 = ~n8721 & n8724;
  assign n8726 = n8721 & ~n8724;
  assign n8727 = ~n8725 & ~n8726;
  assign n8728 = n267 & n8727;
  assign n8729 = n8720 & ~n8728;
  assign n8730 = pi2  & ~n8729;
  assign n8731 = pi2  & ~n8730;
  assign n8732 = ~n8729 & ~n8730;
  assign n8733 = ~n8731 & ~n8732;
  assign n8734 = ~n8685 & ~n8689;
  assign n8735 = pi112  & n340;
  assign n8736 = pi110  & n380;
  assign n8737 = pi111  & n335;
  assign n8738 = ~n8736 & ~n8737;
  assign n8739 = ~n8735 & n8738;
  assign n8740 = n343 & n7795;
  assign n8741 = n8739 & ~n8740;
  assign n8742 = pi5  & ~n8741;
  assign n8743 = pi5  & ~n8742;
  assign n8744 = ~n8741 & ~n8742;
  assign n8745 = ~n8743 & ~n8744;
  assign n8746 = ~n8632 & ~n8636;
  assign n8747 = ~n8615 & ~n8619;
  assign n8748 = pi100  & n1269;
  assign n8749 = pi98  & n1340;
  assign n8750 = pi99  & n1264;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = ~n8748 & n8751;
  assign n8753 = n1272 & n4808;
  assign n8754 = n8752 & ~n8753;
  assign n8755 = pi17  & ~n8754;
  assign n8756 = pi17  & ~n8755;
  assign n8757 = ~n8754 & ~n8755;
  assign n8758 = ~n8756 & ~n8757;
  assign n8759 = ~n8599 & ~n8601;
  assign n8760 = ~n8593 & ~n8595;
  assign n8761 = pi94  & n2004;
  assign n8762 = pi92  & n2141;
  assign n8763 = pi93  & n1999;
  assign n8764 = ~n8762 & ~n8763;
  assign n8765 = ~n8761 & n8764;
  assign n8766 = n2007 & n3499;
  assign n8767 = n8765 & ~n8766;
  assign n8768 = pi23  & ~n8767;
  assign n8769 = pi23  & ~n8768;
  assign n8770 = ~n8767 & ~n8768;
  assign n8771 = ~n8769 & ~n8770;
  assign n8772 = ~n8587 & ~n8589;
  assign n8773 = ~n8531 & ~n8534;
  assign n8774 = pi82  & n4182;
  assign n8775 = pi80  & n4416;
  assign n8776 = pi81  & n4177;
  assign n8777 = ~n8775 & ~n8776;
  assign n8778 = ~n8774 & n8777;
  assign n8779 = n1532 & n4185;
  assign n8780 = n8778 & ~n8779;
  assign n8781 = pi35  & ~n8780;
  assign n8782 = pi35  & ~n8781;
  assign n8783 = ~n8780 & ~n8781;
  assign n8784 = ~n8782 & ~n8783;
  assign n8785 = ~n8525 & ~n8528;
  assign n8786 = pi79  & n4896;
  assign n8787 = pi77  & n5148;
  assign n8788 = pi78  & n4891;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = ~n8786 & n8789;
  assign n8791 = n1105 & n4899;
  assign n8792 = n8790 & ~n8791;
  assign n8793 = pi38  & ~n8792;
  assign n8794 = pi38  & ~n8793;
  assign n8795 = ~n8792 & ~n8793;
  assign n8796 = ~n8794 & ~n8795;
  assign n8797 = ~n8509 & ~n8511;
  assign n8798 = pi76  & n5636;
  assign n8799 = pi74  & n5909;
  assign n8800 = pi75  & n5631;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = ~n8798 & n8801;
  assign n8803 = n881 & n5639;
  assign n8804 = n8802 & ~n8803;
  assign n8805 = pi41  & ~n8804;
  assign n8806 = pi41  & ~n8805;
  assign n8807 = ~n8804 & ~n8805;
  assign n8808 = ~n8806 & ~n8807;
  assign n8809 = ~n8502 & ~n8505;
  assign n8810 = ~n8496 & ~n8499;
  assign n8811 = pi67  & n8137;
  assign n8812 = pi65  & n8471;
  assign n8813 = pi66  & n8132;
  assign n8814 = ~n8812 & ~n8813;
  assign n8815 = ~n8811 & n8814;
  assign n8816 = n313 & n8140;
  assign n8817 = n8815 & ~n8816;
  assign n8818 = pi50  & ~n8817;
  assign n8819 = pi50  & ~n8818;
  assign n8820 = ~n8817 & ~n8818;
  assign n8821 = ~n8819 & ~n8820;
  assign n8822 = pi50  & ~pi51 ;
  assign n8823 = ~pi50  & pi51 ;
  assign n8824 = ~n8822 & ~n8823;
  assign n8825 = pi64  & ~n8824;
  assign n8826 = n8483 & n8825;
  assign n8827 = ~n8483 & ~n8825;
  assign n8828 = ~n8826 & ~n8827;
  assign n8829 = ~n8821 & n8828;
  assign n8830 = n8821 & ~n8828;
  assign n8831 = ~n8829 & ~n8830;
  assign n8832 = pi70  & n7239;
  assign n8833 = pi68  & n7556;
  assign n8834 = pi69  & n7234;
  assign n8835 = ~n8833 & ~n8834;
  assign n8836 = ~n8832 & n8835;
  assign n8837 = n430 & n7242;
  assign n8838 = n8836 & ~n8837;
  assign n8839 = pi47  & ~n8838;
  assign n8840 = pi47  & ~n8839;
  assign n8841 = ~n8838 & ~n8839;
  assign n8842 = ~n8840 & ~n8841;
  assign n8843 = n8831 & ~n8842;
  assign n8844 = ~n8831 & n8842;
  assign n8845 = ~n8843 & ~n8844;
  assign n8846 = n8810 & ~n8845;
  assign n8847 = ~n8810 & n8845;
  assign n8848 = ~n8846 & ~n8847;
  assign n8849 = pi73  & n6396;
  assign n8850 = pi71  & n6735;
  assign n8851 = pi72  & n6391;
  assign n8852 = ~n8850 & ~n8851;
  assign n8853 = ~n8849 & n8852;
  assign n8854 = n639 & n6399;
  assign n8855 = n8853 & ~n8854;
  assign n8856 = pi44  & ~n8855;
  assign n8857 = pi44  & ~n8856;
  assign n8858 = ~n8855 & ~n8856;
  assign n8859 = ~n8857 & ~n8858;
  assign n8860 = ~n8848 & n8859;
  assign n8861 = n8848 & ~n8859;
  assign n8862 = ~n8860 & ~n8861;
  assign n8863 = ~n8809 & n8862;
  assign n8864 = n8809 & ~n8862;
  assign n8865 = ~n8863 & ~n8864;
  assign n8866 = ~n8808 & n8865;
  assign n8867 = n8808 & ~n8865;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = ~n8797 & n8868;
  assign n8870 = n8797 & ~n8868;
  assign n8871 = ~n8869 & ~n8870;
  assign n8872 = ~n8796 & n8871;
  assign n8873 = n8796 & ~n8871;
  assign n8874 = ~n8872 & ~n8873;
  assign n8875 = ~n8785 & n8874;
  assign n8876 = n8785 & ~n8874;
  assign n8877 = ~n8875 & ~n8876;
  assign n8878 = ~n8784 & n8877;
  assign n8879 = n8784 & ~n8877;
  assign n8880 = ~n8878 & ~n8879;
  assign n8881 = ~n8773 & n8880;
  assign n8882 = n8773 & ~n8880;
  assign n8883 = ~n8881 & ~n8882;
  assign n8884 = pi85  & n3550;
  assign n8885 = pi83  & n3735;
  assign n8886 = pi84  & n3545;
  assign n8887 = ~n8885 & ~n8886;
  assign n8888 = ~n8884 & n8887;
  assign n8889 = n1943 & n3553;
  assign n8890 = n8888 & ~n8889;
  assign n8891 = pi32  & ~n8890;
  assign n8892 = pi32  & ~n8891;
  assign n8893 = ~n8890 & ~n8891;
  assign n8894 = ~n8892 & ~n8893;
  assign n8895 = n8883 & ~n8894;
  assign n8896 = n8883 & ~n8895;
  assign n8897 = ~n8894 & ~n8895;
  assign n8898 = ~n8896 & ~n8897;
  assign n8899 = ~n8548 & ~n8554;
  assign n8900 = n8898 & n8899;
  assign n8901 = ~n8898 & ~n8899;
  assign n8902 = ~n8900 & ~n8901;
  assign n8903 = pi88  & n2976;
  assign n8904 = pi86  & n3182;
  assign n8905 = pi87  & n2971;
  assign n8906 = ~n8904 & ~n8905;
  assign n8907 = ~n8903 & n8906;
  assign n8908 = n2277 & n2979;
  assign n8909 = n8907 & ~n8908;
  assign n8910 = pi29  & ~n8909;
  assign n8911 = pi29  & ~n8910;
  assign n8912 = ~n8909 & ~n8910;
  assign n8913 = ~n8911 & ~n8912;
  assign n8914 = ~n8902 & n8913;
  assign n8915 = n8902 & ~n8913;
  assign n8916 = ~n8914 & ~n8915;
  assign n8917 = ~n8572 & n8916;
  assign n8918 = n8572 & ~n8916;
  assign n8919 = ~n8917 & ~n8918;
  assign n8920 = pi91  & n2486;
  assign n8921 = pi89  & n2644;
  assign n8922 = pi90  & n2481;
  assign n8923 = ~n8921 & ~n8922;
  assign n8924 = ~n8920 & n8923;
  assign n8925 = n2489 & n2926;
  assign n8926 = n8924 & ~n8925;
  assign n8927 = pi26  & ~n8926;
  assign n8928 = pi26  & ~n8927;
  assign n8929 = ~n8926 & ~n8927;
  assign n8930 = ~n8928 & ~n8929;
  assign n8931 = n8919 & ~n8930;
  assign n8932 = ~n8919 & n8930;
  assign n8933 = ~n8931 & ~n8932;
  assign n8934 = ~n8772 & n8933;
  assign n8935 = n8772 & ~n8933;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = ~n8771 & n8936;
  assign n8938 = n8771 & ~n8936;
  assign n8939 = ~n8937 & ~n8938;
  assign n8940 = ~n8760 & n8939;
  assign n8941 = n8760 & ~n8939;
  assign n8942 = ~n8940 & ~n8941;
  assign n8943 = pi97  & n1582;
  assign n8944 = pi95  & n1713;
  assign n8945 = pi96  & n1577;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = ~n8943 & n8946;
  assign n8948 = n1585 & n3946;
  assign n8949 = n8947 & ~n8948;
  assign n8950 = pi20  & ~n8949;
  assign n8951 = pi20  & ~n8950;
  assign n8952 = ~n8949 & ~n8950;
  assign n8953 = ~n8951 & ~n8952;
  assign n8954 = n8942 & ~n8953;
  assign n8955 = ~n8942 & n8953;
  assign n8956 = ~n8954 & ~n8955;
  assign n8957 = ~n8759 & n8956;
  assign n8958 = n8759 & ~n8956;
  assign n8959 = ~n8957 & ~n8958;
  assign n8960 = ~n8758 & n8959;
  assign n8961 = n8758 & ~n8959;
  assign n8962 = ~n8960 & ~n8961;
  assign n8963 = n8747 & ~n8962;
  assign n8964 = ~n8747 & n8962;
  assign n8965 = ~n8963 & ~n8964;
  assign n8966 = pi103  & n918;
  assign n8967 = pi101  & n1031;
  assign n8968 = pi102  & n913;
  assign n8969 = ~n8967 & ~n8968;
  assign n8970 = ~n8966 & n8969;
  assign n8971 = n921 & n5540;
  assign n8972 = n8970 & ~n8971;
  assign n8973 = pi14  & ~n8972;
  assign n8974 = pi14  & ~n8973;
  assign n8975 = ~n8972 & ~n8973;
  assign n8976 = ~n8974 & ~n8975;
  assign n8977 = n8965 & ~n8976;
  assign n8978 = ~n8965 & n8976;
  assign n8979 = ~n8977 & ~n8978;
  assign n8980 = n8746 & ~n8979;
  assign n8981 = ~n8746 & n8979;
  assign n8982 = ~n8980 & ~n8981;
  assign n8983 = pi106  & n675;
  assign n8984 = pi104  & n769;
  assign n8985 = pi105  & n670;
  assign n8986 = ~n8984 & ~n8985;
  assign n8987 = ~n8983 & n8986;
  assign n8988 = n678 & n6090;
  assign n8989 = n8987 & ~n8988;
  assign n8990 = pi11  & ~n8989;
  assign n8991 = pi11  & ~n8990;
  assign n8992 = ~n8989 & ~n8990;
  assign n8993 = ~n8991 & ~n8992;
  assign n8994 = ~n8982 & n8993;
  assign n8995 = n8982 & ~n8993;
  assign n8996 = ~n8994 & ~n8995;
  assign n8997 = ~n8649 & ~n8653;
  assign n8998 = n8996 & ~n8997;
  assign n8999 = ~n8996 & n8997;
  assign n9000 = ~n8998 & ~n8999;
  assign n9001 = pi109  & n493;
  assign n9002 = pi107  & n533;
  assign n9003 = pi108  & n488;
  assign n9004 = ~n9002 & ~n9003;
  assign n9005 = ~n9001 & n9004;
  assign n9006 = n496 & n7170;
  assign n9007 = n9005 & ~n9006;
  assign n9008 = pi8  & ~n9007;
  assign n9009 = pi8  & ~n9008;
  assign n9010 = ~n9007 & ~n9008;
  assign n9011 = ~n9009 & ~n9010;
  assign n9012 = n9000 & ~n9011;
  assign n9013 = ~n9000 & n9011;
  assign n9014 = ~n9012 & ~n9013;
  assign n9015 = ~n8671 & n9014;
  assign n9016 = n8671 & ~n9014;
  assign n9017 = ~n9015 & ~n9016;
  assign n9018 = n8745 & ~n9017;
  assign n9019 = ~n8745 & n9017;
  assign n9020 = ~n9018 & ~n9019;
  assign n9021 = ~n8734 & n9020;
  assign n9022 = n8734 & ~n9020;
  assign n9023 = ~n9021 & ~n9022;
  assign n9024 = ~n8733 & n9023;
  assign n9025 = n8733 & ~n9023;
  assign n9026 = ~n9024 & ~n9025;
  assign n9027 = ~n8715 & n9026;
  assign n9028 = n8715 & ~n9026;
  assign po51  = ~n9027 & ~n9028;
  assign n9030 = ~n9024 & ~n9027;
  assign n9031 = pi116  & n264;
  assign n9032 = pi114  & n281;
  assign n9033 = pi115  & n259;
  assign n9034 = ~n9032 & ~n9033;
  assign n9035 = ~n9031 & n9034;
  assign n9036 = ~n8723 & ~n8725;
  assign n9037 = ~pi115  & ~pi116 ;
  assign n9038 = pi115  & pi116 ;
  assign n9039 = ~n9037 & ~n9038;
  assign n9040 = ~n9036 & n9039;
  assign n9041 = n9036 & ~n9039;
  assign n9042 = ~n9040 & ~n9041;
  assign n9043 = n267 & n9042;
  assign n9044 = n9035 & ~n9043;
  assign n9045 = pi2  & ~n9044;
  assign n9046 = pi2  & ~n9045;
  assign n9047 = ~n9044 & ~n9045;
  assign n9048 = ~n9046 & ~n9047;
  assign n9049 = ~n9019 & ~n9021;
  assign n9050 = ~n9012 & ~n9015;
  assign n9051 = ~n8995 & ~n8998;
  assign n9052 = ~n8977 & ~n8981;
  assign n9053 = ~n8960 & ~n8964;
  assign n9054 = ~n8954 & ~n8957;
  assign n9055 = ~n8937 & ~n8940;
  assign n9056 = ~n8931 & ~n8934;
  assign n9057 = pi92  & n2486;
  assign n9058 = pi90  & n2644;
  assign n9059 = pi91  & n2481;
  assign n9060 = ~n9058 & ~n9059;
  assign n9061 = ~n9057 & n9060;
  assign n9062 = n2489 & n3119;
  assign n9063 = n9061 & ~n9062;
  assign n9064 = pi26  & ~n9063;
  assign n9065 = pi26  & ~n9064;
  assign n9066 = ~n9063 & ~n9064;
  assign n9067 = ~n9065 & ~n9066;
  assign n9068 = ~n8915 & ~n8917;
  assign n9069 = ~n8895 & ~n8901;
  assign n9070 = ~n8878 & ~n8881;
  assign n9071 = ~n8872 & ~n8875;
  assign n9072 = ~n8866 & ~n8869;
  assign n9073 = ~n8861 & ~n8863;
  assign n9074 = ~n8843 & ~n8847;
  assign n9075 = ~n8826 & ~n8829;
  assign n9076 = pi68  & n8137;
  assign n9077 = pi66  & n8471;
  assign n9078 = pi67  & n8132;
  assign n9079 = ~n9077 & ~n9078;
  assign n9080 = ~n9076 & n9079;
  assign n9081 = n364 & n8140;
  assign n9082 = n9080 & ~n9081;
  assign n9083 = pi50  & ~n9082;
  assign n9084 = pi50  & ~n9083;
  assign n9085 = ~n9082 & ~n9083;
  assign n9086 = ~n9084 & ~n9085;
  assign n9087 = pi53  & ~n8825;
  assign n9088 = ~pi51  & pi52 ;
  assign n9089 = pi51  & ~pi52 ;
  assign n9090 = ~n9088 & ~n9089;
  assign n9091 = n8824 & ~n9090;
  assign n9092 = pi64  & n9091;
  assign n9093 = ~pi52  & pi53 ;
  assign n9094 = pi52  & ~pi53 ;
  assign n9095 = ~n9093 & ~n9094;
  assign n9096 = ~n8824 & n9095;
  assign n9097 = pi65  & n9096;
  assign n9098 = ~n9092 & ~n9097;
  assign n9099 = ~n8824 & ~n9095;
  assign n9100 = n270 & n9099;
  assign n9101 = n9098 & ~n9100;
  assign n9102 = pi53  & ~n9101;
  assign n9103 = pi53  & ~n9102;
  assign n9104 = ~n9101 & ~n9102;
  assign n9105 = ~n9103 & ~n9104;
  assign n9106 = n9087 & ~n9105;
  assign n9107 = ~n9087 & n9105;
  assign n9108 = ~n9106 & ~n9107;
  assign n9109 = n9086 & ~n9108;
  assign n9110 = ~n9086 & n9108;
  assign n9111 = ~n9109 & ~n9110;
  assign n9112 = ~n9075 & n9111;
  assign n9113 = n9075 & ~n9111;
  assign n9114 = ~n9112 & ~n9113;
  assign n9115 = pi71  & n7239;
  assign n9116 = pi69  & n7556;
  assign n9117 = pi70  & n7234;
  assign n9118 = ~n9116 & ~n9117;
  assign n9119 = ~n9115 & n9118;
  assign n9120 = n476 & n7242;
  assign n9121 = n9119 & ~n9120;
  assign n9122 = pi47  & ~n9121;
  assign n9123 = pi47  & ~n9122;
  assign n9124 = ~n9121 & ~n9122;
  assign n9125 = ~n9123 & ~n9124;
  assign n9126 = n9114 & ~n9125;
  assign n9127 = ~n9114 & n9125;
  assign n9128 = ~n9126 & ~n9127;
  assign n9129 = n9074 & ~n9128;
  assign n9130 = ~n9074 & n9128;
  assign n9131 = ~n9129 & ~n9130;
  assign n9132 = pi74  & n6396;
  assign n9133 = pi72  & n6735;
  assign n9134 = pi73  & n6391;
  assign n9135 = ~n9133 & ~n9134;
  assign n9136 = ~n9132 & n9135;
  assign n9137 = n722 & n6399;
  assign n9138 = n9136 & ~n9137;
  assign n9139 = pi44  & ~n9138;
  assign n9140 = pi44  & ~n9139;
  assign n9141 = ~n9138 & ~n9139;
  assign n9142 = ~n9140 & ~n9141;
  assign n9143 = n9131 & ~n9142;
  assign n9144 = ~n9131 & n9142;
  assign n9145 = ~n9073 & ~n9144;
  assign n9146 = ~n9143 & n9145;
  assign n9147 = ~n9073 & ~n9146;
  assign n9148 = ~n9143 & ~n9146;
  assign n9149 = ~n9144 & n9148;
  assign n9150 = ~n9147 & ~n9149;
  assign n9151 = pi77  & n5636;
  assign n9152 = pi75  & n5909;
  assign n9153 = pi76  & n5631;
  assign n9154 = ~n9152 & ~n9153;
  assign n9155 = ~n9151 & n9154;
  assign n9156 = n984 & n5639;
  assign n9157 = n9155 & ~n9156;
  assign n9158 = pi41  & ~n9157;
  assign n9159 = pi41  & ~n9158;
  assign n9160 = ~n9157 & ~n9158;
  assign n9161 = ~n9159 & ~n9160;
  assign n9162 = n9150 & n9161;
  assign n9163 = ~n9150 & ~n9161;
  assign n9164 = ~n9162 & ~n9163;
  assign n9165 = ~n9072 & n9164;
  assign n9166 = n9072 & ~n9164;
  assign n9167 = ~n9165 & ~n9166;
  assign n9168 = pi80  & n4896;
  assign n9169 = pi78  & n5148;
  assign n9170 = pi79  & n4891;
  assign n9171 = ~n9169 & ~n9170;
  assign n9172 = ~n9168 & n9171;
  assign n9173 = n1205 & n4899;
  assign n9174 = n9172 & ~n9173;
  assign n9175 = pi38  & ~n9174;
  assign n9176 = pi38  & ~n9175;
  assign n9177 = ~n9174 & ~n9175;
  assign n9178 = ~n9176 & ~n9177;
  assign n9179 = n9167 & ~n9178;
  assign n9180 = ~n9167 & n9178;
  assign n9181 = ~n9179 & ~n9180;
  assign n9182 = n9071 & ~n9181;
  assign n9183 = ~n9071 & n9181;
  assign n9184 = ~n9182 & ~n9183;
  assign n9185 = pi83  & n4182;
  assign n9186 = pi81  & n4416;
  assign n9187 = pi82  & n4177;
  assign n9188 = ~n9186 & ~n9187;
  assign n9189 = ~n9185 & n9188;
  assign n9190 = n1672 & n4185;
  assign n9191 = n9189 & ~n9190;
  assign n9192 = pi35  & ~n9191;
  assign n9193 = pi35  & ~n9192;
  assign n9194 = ~n9191 & ~n9192;
  assign n9195 = ~n9193 & ~n9194;
  assign n9196 = n9184 & ~n9195;
  assign n9197 = ~n9184 & n9195;
  assign n9198 = ~n9070 & ~n9197;
  assign n9199 = ~n9196 & n9198;
  assign n9200 = ~n9070 & ~n9199;
  assign n9201 = ~n9196 & ~n9199;
  assign n9202 = ~n9197 & n9201;
  assign n9203 = ~n9200 & ~n9202;
  assign n9204 = pi86  & n3550;
  assign n9205 = pi84  & n3735;
  assign n9206 = pi85  & n3545;
  assign n9207 = ~n9205 & ~n9206;
  assign n9208 = ~n9204 & n9207;
  assign n9209 = n2099 & n3553;
  assign n9210 = n9208 & ~n9209;
  assign n9211 = pi32  & ~n9210;
  assign n9212 = pi32  & ~n9211;
  assign n9213 = ~n9210 & ~n9211;
  assign n9214 = ~n9212 & ~n9213;
  assign n9215 = ~n9203 & ~n9214;
  assign n9216 = n9203 & n9214;
  assign n9217 = ~n9215 & ~n9216;
  assign n9218 = n9069 & ~n9217;
  assign n9219 = ~n9069 & n9217;
  assign n9220 = ~n9218 & ~n9219;
  assign n9221 = pi89  & n2976;
  assign n9222 = pi87  & n3182;
  assign n9223 = pi88  & n2971;
  assign n9224 = ~n9222 & ~n9223;
  assign n9225 = ~n9221 & n9224;
  assign n9226 = n2432 & n2979;
  assign n9227 = n9225 & ~n9226;
  assign n9228 = pi29  & ~n9227;
  assign n9229 = pi29  & ~n9228;
  assign n9230 = ~n9227 & ~n9228;
  assign n9231 = ~n9229 & ~n9230;
  assign n9232 = n9220 & ~n9231;
  assign n9233 = ~n9220 & n9231;
  assign n9234 = ~n9232 & ~n9233;
  assign n9235 = ~n9068 & n9234;
  assign n9236 = n9068 & ~n9234;
  assign n9237 = ~n9235 & ~n9236;
  assign n9238 = ~n9067 & n9237;
  assign n9239 = n9067 & ~n9237;
  assign n9240 = ~n9238 & ~n9239;
  assign n9241 = n9056 & ~n9240;
  assign n9242 = ~n9056 & n9240;
  assign n9243 = ~n9241 & ~n9242;
  assign n9244 = pi95  & n2004;
  assign n9245 = pi93  & n2141;
  assign n9246 = pi94  & n1999;
  assign n9247 = ~n9245 & ~n9246;
  assign n9248 = ~n9244 & n9247;
  assign n9249 = n2007 & n3710;
  assign n9250 = n9248 & ~n9249;
  assign n9251 = pi23  & ~n9250;
  assign n9252 = pi23  & ~n9251;
  assign n9253 = ~n9250 & ~n9251;
  assign n9254 = ~n9252 & ~n9253;
  assign n9255 = n9243 & ~n9254;
  assign n9256 = ~n9243 & n9254;
  assign n9257 = ~n9255 & ~n9256;
  assign n9258 = n9055 & ~n9257;
  assign n9259 = ~n9055 & n9257;
  assign n9260 = ~n9258 & ~n9259;
  assign n9261 = pi98  & n1582;
  assign n9262 = pi96  & n1713;
  assign n9263 = pi97  & n1577;
  assign n9264 = ~n9262 & ~n9263;
  assign n9265 = ~n9261 & n9264;
  assign n9266 = n1585 & n4360;
  assign n9267 = n9265 & ~n9266;
  assign n9268 = pi20  & ~n9267;
  assign n9269 = pi20  & ~n9268;
  assign n9270 = ~n9267 & ~n9268;
  assign n9271 = ~n9269 & ~n9270;
  assign n9272 = n9260 & ~n9271;
  assign n9273 = ~n9260 & n9271;
  assign n9274 = ~n9272 & ~n9273;
  assign n9275 = n9054 & ~n9274;
  assign n9276 = ~n9054 & n9274;
  assign n9277 = ~n9275 & ~n9276;
  assign n9278 = pi101  & n1269;
  assign n9279 = pi99  & n1340;
  assign n9280 = pi100  & n1264;
  assign n9281 = ~n9279 & ~n9280;
  assign n9282 = ~n9278 & n9281;
  assign n9283 = n1272 & n5056;
  assign n9284 = n9282 & ~n9283;
  assign n9285 = pi17  & ~n9284;
  assign n9286 = pi17  & ~n9285;
  assign n9287 = ~n9284 & ~n9285;
  assign n9288 = ~n9286 & ~n9287;
  assign n9289 = n9277 & ~n9288;
  assign n9290 = ~n9277 & n9288;
  assign n9291 = ~n9289 & ~n9290;
  assign n9292 = n9053 & ~n9291;
  assign n9293 = ~n9053 & n9291;
  assign n9294 = ~n9292 & ~n9293;
  assign n9295 = pi104  & n918;
  assign n9296 = pi102  & n1031;
  assign n9297 = pi103  & n913;
  assign n9298 = ~n9296 & ~n9297;
  assign n9299 = ~n9295 & n9298;
  assign n9300 = n921 & n5565;
  assign n9301 = n9299 & ~n9300;
  assign n9302 = pi14  & ~n9301;
  assign n9303 = pi14  & ~n9302;
  assign n9304 = ~n9301 & ~n9302;
  assign n9305 = ~n9303 & ~n9304;
  assign n9306 = n9294 & ~n9305;
  assign n9307 = ~n9294 & n9305;
  assign n9308 = ~n9306 & ~n9307;
  assign n9309 = n9052 & ~n9308;
  assign n9310 = ~n9052 & n9308;
  assign n9311 = ~n9309 & ~n9310;
  assign n9312 = pi107  & n675;
  assign n9313 = pi105  & n769;
  assign n9314 = pi106  & n670;
  assign n9315 = ~n9313 & ~n9314;
  assign n9316 = ~n9312 & n9315;
  assign n9317 = n678 & n6614;
  assign n9318 = n9316 & ~n9317;
  assign n9319 = pi11  & ~n9318;
  assign n9320 = pi11  & ~n9319;
  assign n9321 = ~n9318 & ~n9319;
  assign n9322 = ~n9320 & ~n9321;
  assign n9323 = n9311 & ~n9322;
  assign n9324 = ~n9311 & n9322;
  assign n9325 = ~n9051 & ~n9324;
  assign n9326 = ~n9323 & n9325;
  assign n9327 = ~n9051 & ~n9326;
  assign n9328 = ~n9323 & ~n9326;
  assign n9329 = ~n9324 & n9328;
  assign n9330 = ~n9327 & ~n9329;
  assign n9331 = pi110  & n493;
  assign n9332 = pi108  & n533;
  assign n9333 = pi109  & n488;
  assign n9334 = ~n9332 & ~n9333;
  assign n9335 = ~n9331 & n9334;
  assign n9336 = n496 & n7474;
  assign n9337 = n9335 & ~n9336;
  assign n9338 = pi8  & ~n9337;
  assign n9339 = pi8  & ~n9338;
  assign n9340 = ~n9337 & ~n9338;
  assign n9341 = ~n9339 & ~n9340;
  assign n9342 = ~n9330 & ~n9341;
  assign n9343 = n9330 & n9341;
  assign n9344 = ~n9342 & ~n9343;
  assign n9345 = n9050 & ~n9344;
  assign n9346 = ~n9050 & n9344;
  assign n9347 = ~n9345 & ~n9346;
  assign n9348 = pi113  & n340;
  assign n9349 = pi111  & n380;
  assign n9350 = pi112  & n335;
  assign n9351 = ~n9349 & ~n9350;
  assign n9352 = ~n9348 & n9351;
  assign n9353 = n343 & n8387;
  assign n9354 = n9352 & ~n9353;
  assign n9355 = pi5  & ~n9354;
  assign n9356 = pi5  & ~n9355;
  assign n9357 = ~n9354 & ~n9355;
  assign n9358 = ~n9356 & ~n9357;
  assign n9359 = n9347 & ~n9358;
  assign n9360 = ~n9347 & n9358;
  assign n9361 = ~n9359 & ~n9360;
  assign n9362 = ~n9049 & n9361;
  assign n9363 = n9049 & ~n9361;
  assign n9364 = ~n9362 & ~n9363;
  assign n9365 = ~n9048 & n9364;
  assign n9366 = n9048 & ~n9364;
  assign n9367 = ~n9365 & ~n9366;
  assign n9368 = ~n9030 & n9367;
  assign n9369 = n9030 & ~n9367;
  assign po52  = ~n9368 & ~n9369;
  assign n9371 = ~n9365 & ~n9368;
  assign n9372 = ~n9359 & ~n9362;
  assign n9373 = ~n9342 & ~n9346;
  assign n9374 = ~n9306 & ~n9310;
  assign n9375 = ~n9289 & ~n9293;
  assign n9376 = ~n9272 & ~n9276;
  assign n9377 = ~n9255 & ~n9259;
  assign n9378 = pi96  & n2004;
  assign n9379 = pi94  & n2141;
  assign n9380 = pi95  & n1999;
  assign n9381 = ~n9379 & ~n9380;
  assign n9382 = ~n9378 & n9381;
  assign n9383 = n2007 & n3921;
  assign n9384 = n9382 & ~n9383;
  assign n9385 = pi23  & ~n9384;
  assign n9386 = pi23  & ~n9385;
  assign n9387 = ~n9384 & ~n9385;
  assign n9388 = ~n9386 & ~n9387;
  assign n9389 = ~n9238 & ~n9242;
  assign n9390 = pi93  & n2486;
  assign n9391 = pi91  & n2644;
  assign n9392 = pi92  & n2481;
  assign n9393 = ~n9391 & ~n9392;
  assign n9394 = ~n9390 & n9393;
  assign n9395 = n2489 & n3144;
  assign n9396 = n9394 & ~n9395;
  assign n9397 = pi26  & ~n9396;
  assign n9398 = pi26  & ~n9397;
  assign n9399 = ~n9396 & ~n9397;
  assign n9400 = ~n9398 & ~n9399;
  assign n9401 = ~n9232 & ~n9235;
  assign n9402 = pi90  & n2976;
  assign n9403 = pi88  & n3182;
  assign n9404 = pi89  & n2971;
  assign n9405 = ~n9403 & ~n9404;
  assign n9406 = ~n9402 & n9405;
  assign n9407 = n2606 & n2979;
  assign n9408 = n9406 & ~n9407;
  assign n9409 = pi29  & ~n9408;
  assign n9410 = pi29  & ~n9409;
  assign n9411 = ~n9408 & ~n9409;
  assign n9412 = ~n9410 & ~n9411;
  assign n9413 = ~n9215 & ~n9219;
  assign n9414 = pi87  & n3550;
  assign n9415 = pi85  & n3735;
  assign n9416 = pi86  & n3545;
  assign n9417 = ~n9415 & ~n9416;
  assign n9418 = ~n9414 & n9417;
  assign n9419 = n2252 & n3553;
  assign n9420 = n9418 & ~n9419;
  assign n9421 = pi32  & ~n9420;
  assign n9422 = pi32  & ~n9421;
  assign n9423 = ~n9420 & ~n9421;
  assign n9424 = ~n9422 & ~n9423;
  assign n9425 = ~n9179 & ~n9183;
  assign n9426 = pi81  & n4896;
  assign n9427 = pi79  & n5148;
  assign n9428 = pi80  & n4891;
  assign n9429 = ~n9427 & ~n9428;
  assign n9430 = ~n9426 & n9429;
  assign n9431 = n1413 & n4899;
  assign n9432 = n9430 & ~n9431;
  assign n9433 = pi38  & ~n9432;
  assign n9434 = pi38  & ~n9433;
  assign n9435 = ~n9432 & ~n9433;
  assign n9436 = ~n9434 & ~n9435;
  assign n9437 = ~n9163 & ~n9165;
  assign n9438 = pi75  & n6396;
  assign n9439 = pi73  & n6735;
  assign n9440 = pi74  & n6391;
  assign n9441 = ~n9439 & ~n9440;
  assign n9442 = ~n9438 & n9441;
  assign n9443 = n747 & n6399;
  assign n9444 = n9442 & ~n9443;
  assign n9445 = pi44  & ~n9444;
  assign n9446 = pi44  & ~n9445;
  assign n9447 = ~n9444 & ~n9445;
  assign n9448 = ~n9446 & ~n9447;
  assign n9449 = ~n9126 & ~n9130;
  assign n9450 = ~n9110 & ~n9112;
  assign n9451 = pi66  & n9096;
  assign n9452 = n8824 & ~n9095;
  assign n9453 = n9090 & n9452;
  assign n9454 = pi64  & n9453;
  assign n9455 = pi65  & n9091;
  assign n9456 = ~n9454 & ~n9455;
  assign n9457 = ~n9451 & n9456;
  assign n9458 = n291 & n9099;
  assign n9459 = n9457 & ~n9458;
  assign n9460 = pi53  & ~n9459;
  assign n9461 = pi53  & ~n9460;
  assign n9462 = ~n9459 & ~n9460;
  assign n9463 = ~n9461 & ~n9462;
  assign n9464 = ~n9106 & n9463;
  assign n9465 = n9106 & ~n9463;
  assign n9466 = ~n9464 & ~n9465;
  assign n9467 = pi69  & n8137;
  assign n9468 = pi67  & n8471;
  assign n9469 = pi68  & n8132;
  assign n9470 = ~n9468 & ~n9469;
  assign n9471 = ~n9467 & n9470;
  assign n9472 = n405 & n8140;
  assign n9473 = n9471 & ~n9472;
  assign n9474 = pi50  & ~n9473;
  assign n9475 = pi50  & ~n9474;
  assign n9476 = ~n9473 & ~n9474;
  assign n9477 = ~n9475 & ~n9476;
  assign n9478 = n9466 & ~n9477;
  assign n9479 = ~n9466 & n9477;
  assign n9480 = ~n9450 & ~n9479;
  assign n9481 = ~n9478 & n9480;
  assign n9482 = ~n9450 & ~n9481;
  assign n9483 = ~n9478 & ~n9481;
  assign n9484 = ~n9479 & n9483;
  assign n9485 = ~n9482 & ~n9484;
  assign n9486 = pi72  & n7239;
  assign n9487 = pi70  & n7556;
  assign n9488 = pi71  & n7234;
  assign n9489 = ~n9487 & ~n9488;
  assign n9490 = ~n9486 & n9489;
  assign n9491 = n575 & n7242;
  assign n9492 = n9490 & ~n9491;
  assign n9493 = pi47  & ~n9492;
  assign n9494 = pi47  & ~n9493;
  assign n9495 = ~n9492 & ~n9493;
  assign n9496 = ~n9494 & ~n9495;
  assign n9497 = n9485 & n9496;
  assign n9498 = ~n9485 & ~n9496;
  assign n9499 = ~n9497 & ~n9498;
  assign n9500 = ~n9449 & n9499;
  assign n9501 = n9449 & ~n9499;
  assign n9502 = ~n9500 & ~n9501;
  assign n9503 = n9448 & ~n9502;
  assign n9504 = ~n9448 & n9502;
  assign n9505 = ~n9503 & ~n9504;
  assign n9506 = ~n9148 & n9505;
  assign n9507 = n9148 & ~n9505;
  assign n9508 = ~n9506 & ~n9507;
  assign n9509 = pi78  & n5636;
  assign n9510 = pi76  & n5909;
  assign n9511 = pi77  & n5631;
  assign n9512 = ~n9510 & ~n9511;
  assign n9513 = ~n9509 & n9512;
  assign n9514 = n1009 & n5639;
  assign n9515 = n9513 & ~n9514;
  assign n9516 = pi41  & ~n9515;
  assign n9517 = pi41  & ~n9516;
  assign n9518 = ~n9515 & ~n9516;
  assign n9519 = ~n9517 & ~n9518;
  assign n9520 = n9508 & ~n9519;
  assign n9521 = ~n9508 & n9519;
  assign n9522 = ~n9520 & ~n9521;
  assign n9523 = ~n9437 & n9522;
  assign n9524 = n9437 & ~n9522;
  assign n9525 = ~n9523 & ~n9524;
  assign n9526 = ~n9436 & n9525;
  assign n9527 = n9436 & ~n9525;
  assign n9528 = ~n9526 & ~n9527;
  assign n9529 = ~n9425 & n9528;
  assign n9530 = n9425 & ~n9528;
  assign n9531 = ~n9529 & ~n9530;
  assign n9532 = pi84  & n4182;
  assign n9533 = pi82  & n4416;
  assign n9534 = pi83  & n4177;
  assign n9535 = ~n9533 & ~n9534;
  assign n9536 = ~n9532 & n9535;
  assign n9537 = n1805 & n4185;
  assign n9538 = n9536 & ~n9537;
  assign n9539 = pi35  & ~n9538;
  assign n9540 = pi35  & ~n9539;
  assign n9541 = ~n9538 & ~n9539;
  assign n9542 = ~n9540 & ~n9541;
  assign n9543 = n9531 & ~n9542;
  assign n9544 = n9531 & ~n9543;
  assign n9545 = ~n9542 & ~n9543;
  assign n9546 = ~n9544 & ~n9545;
  assign n9547 = ~n9201 & ~n9546;
  assign n9548 = n9201 & n9546;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = ~n9424 & n9549;
  assign n9551 = n9424 & ~n9549;
  assign n9552 = ~n9550 & ~n9551;
  assign n9553 = ~n9413 & n9552;
  assign n9554 = n9413 & ~n9552;
  assign n9555 = ~n9553 & ~n9554;
  assign n9556 = n9412 & ~n9555;
  assign n9557 = ~n9412 & n9555;
  assign n9558 = ~n9556 & ~n9557;
  assign n9559 = ~n9401 & n9558;
  assign n9560 = n9401 & ~n9558;
  assign n9561 = ~n9559 & ~n9560;
  assign n9562 = n9400 & ~n9561;
  assign n9563 = ~n9400 & n9561;
  assign n9564 = ~n9562 & ~n9563;
  assign n9565 = ~n9389 & n9564;
  assign n9566 = n9389 & ~n9564;
  assign n9567 = ~n9565 & ~n9566;
  assign n9568 = n9388 & ~n9567;
  assign n9569 = ~n9388 & n9567;
  assign n9570 = ~n9568 & ~n9569;
  assign n9571 = ~n9377 & n9570;
  assign n9572 = n9377 & ~n9570;
  assign n9573 = ~n9571 & ~n9572;
  assign n9574 = pi99  & n1582;
  assign n9575 = pi97  & n1713;
  assign n9576 = pi98  & n1577;
  assign n9577 = ~n9575 & ~n9576;
  assign n9578 = ~n9574 & n9577;
  assign n9579 = n1585 & n4584;
  assign n9580 = n9578 & ~n9579;
  assign n9581 = pi20  & ~n9580;
  assign n9582 = pi20  & ~n9581;
  assign n9583 = ~n9580 & ~n9581;
  assign n9584 = ~n9582 & ~n9583;
  assign n9585 = n9573 & ~n9584;
  assign n9586 = ~n9573 & n9584;
  assign n9587 = ~n9585 & ~n9586;
  assign n9588 = n9376 & ~n9587;
  assign n9589 = ~n9376 & n9587;
  assign n9590 = ~n9588 & ~n9589;
  assign n9591 = pi102  & n1269;
  assign n9592 = pi100  & n1340;
  assign n9593 = pi101  & n1264;
  assign n9594 = ~n9592 & ~n9593;
  assign n9595 = ~n9591 & n9594;
  assign n9596 = n1272 & n5296;
  assign n9597 = n9595 & ~n9596;
  assign n9598 = pi17  & ~n9597;
  assign n9599 = pi17  & ~n9598;
  assign n9600 = ~n9597 & ~n9598;
  assign n9601 = ~n9599 & ~n9600;
  assign n9602 = n9590 & ~n9601;
  assign n9603 = ~n9590 & n9601;
  assign n9604 = ~n9602 & ~n9603;
  assign n9605 = n9375 & ~n9604;
  assign n9606 = ~n9375 & n9604;
  assign n9607 = ~n9605 & ~n9606;
  assign n9608 = pi105  & n918;
  assign n9609 = pi103  & n1031;
  assign n9610 = pi104  & n913;
  assign n9611 = ~n9609 & ~n9610;
  assign n9612 = ~n9608 & n9611;
  assign n9613 = n921 & n6065;
  assign n9614 = n9612 & ~n9613;
  assign n9615 = pi14  & ~n9614;
  assign n9616 = pi14  & ~n9615;
  assign n9617 = ~n9614 & ~n9615;
  assign n9618 = ~n9616 & ~n9617;
  assign n9619 = n9607 & ~n9618;
  assign n9620 = ~n9607 & n9618;
  assign n9621 = ~n9619 & ~n9620;
  assign n9622 = n9374 & ~n9621;
  assign n9623 = ~n9374 & n9621;
  assign n9624 = ~n9622 & ~n9623;
  assign n9625 = pi108  & n675;
  assign n9626 = pi106  & n769;
  assign n9627 = pi107  & n670;
  assign n9628 = ~n9626 & ~n9627;
  assign n9629 = ~n9625 & n9628;
  assign n9630 = n678 & n6639;
  assign n9631 = n9629 & ~n9630;
  assign n9632 = pi11  & ~n9631;
  assign n9633 = pi11  & ~n9632;
  assign n9634 = ~n9631 & ~n9632;
  assign n9635 = ~n9633 & ~n9634;
  assign n9636 = n9624 & ~n9635;
  assign n9637 = ~n9624 & n9635;
  assign n9638 = ~n9328 & ~n9637;
  assign n9639 = ~n9636 & n9638;
  assign n9640 = ~n9328 & ~n9639;
  assign n9641 = ~n9636 & ~n9639;
  assign n9642 = ~n9637 & n9641;
  assign n9643 = ~n9640 & ~n9642;
  assign n9644 = pi111  & n493;
  assign n9645 = pi109  & n533;
  assign n9646 = pi110  & n488;
  assign n9647 = ~n9645 & ~n9646;
  assign n9648 = ~n9644 & n9647;
  assign n9649 = n496 & n7770;
  assign n9650 = n9648 & ~n9649;
  assign n9651 = pi8  & ~n9650;
  assign n9652 = pi8  & ~n9651;
  assign n9653 = ~n9650 & ~n9651;
  assign n9654 = ~n9652 & ~n9653;
  assign n9655 = ~n9643 & ~n9654;
  assign n9656 = n9643 & n9654;
  assign n9657 = ~n9655 & ~n9656;
  assign n9658 = n9373 & ~n9657;
  assign n9659 = ~n9373 & n9657;
  assign n9660 = ~n9658 & ~n9659;
  assign n9661 = pi114  & n340;
  assign n9662 = pi112  & n380;
  assign n9663 = pi113  & n335;
  assign n9664 = ~n9662 & ~n9663;
  assign n9665 = ~n9661 & n9664;
  assign n9666 = n343 & n8702;
  assign n9667 = n9665 & ~n9666;
  assign n9668 = pi5  & ~n9667;
  assign n9669 = pi5  & ~n9668;
  assign n9670 = ~n9667 & ~n9668;
  assign n9671 = ~n9669 & ~n9670;
  assign n9672 = n9660 & ~n9671;
  assign n9673 = ~n9660 & n9671;
  assign n9674 = ~n9372 & ~n9673;
  assign n9675 = ~n9672 & n9674;
  assign n9676 = ~n9372 & ~n9675;
  assign n9677 = ~n9672 & ~n9675;
  assign n9678 = ~n9673 & n9677;
  assign n9679 = ~n9676 & ~n9678;
  assign n9680 = pi117  & n264;
  assign n9681 = pi115  & n281;
  assign n9682 = pi116  & n259;
  assign n9683 = ~n9681 & ~n9682;
  assign n9684 = ~n9680 & n9683;
  assign n9685 = ~n9038 & ~n9040;
  assign n9686 = ~pi116  & ~pi117 ;
  assign n9687 = pi116  & pi117 ;
  assign n9688 = ~n9686 & ~n9687;
  assign n9689 = ~n9685 & n9688;
  assign n9690 = n9685 & ~n9688;
  assign n9691 = ~n9689 & ~n9690;
  assign n9692 = n267 & n9691;
  assign n9693 = n9684 & ~n9692;
  assign n9694 = pi2  & ~n9693;
  assign n9695 = pi2  & ~n9694;
  assign n9696 = ~n9693 & ~n9694;
  assign n9697 = ~n9695 & ~n9696;
  assign n9698 = ~n9679 & ~n9697;
  assign n9699 = n9679 & n9697;
  assign n9700 = ~n9698 & ~n9699;
  assign n9701 = ~n9371 & n9700;
  assign n9702 = n9371 & ~n9700;
  assign po53  = ~n9701 & ~n9702;
  assign n9704 = ~n9698 & ~n9701;
  assign n9705 = pi118  & n264;
  assign n9706 = pi116  & n281;
  assign n9707 = pi117  & n259;
  assign n9708 = ~n9706 & ~n9707;
  assign n9709 = ~n9705 & n9708;
  assign n9710 = ~n9687 & ~n9689;
  assign n9711 = ~pi117  & ~pi118 ;
  assign n9712 = pi117  & pi118 ;
  assign n9713 = ~n9711 & ~n9712;
  assign n9714 = ~n9710 & n9713;
  assign n9715 = n9710 & ~n9713;
  assign n9716 = ~n9714 & ~n9715;
  assign n9717 = n267 & n9716;
  assign n9718 = n9709 & ~n9717;
  assign n9719 = pi2  & ~n9718;
  assign n9720 = pi2  & ~n9719;
  assign n9721 = ~n9718 & ~n9719;
  assign n9722 = ~n9720 & ~n9721;
  assign n9723 = ~n9655 & ~n9659;
  assign n9724 = pi112  & n493;
  assign n9725 = pi110  & n533;
  assign n9726 = pi111  & n488;
  assign n9727 = ~n9725 & ~n9726;
  assign n9728 = ~n9724 & n9727;
  assign n9729 = n496 & n7795;
  assign n9730 = n9728 & ~n9729;
  assign n9731 = pi8  & ~n9730;
  assign n9732 = pi8  & ~n9731;
  assign n9733 = ~n9730 & ~n9731;
  assign n9734 = ~n9732 & ~n9733;
  assign n9735 = pi109  & n675;
  assign n9736 = pi107  & n769;
  assign n9737 = pi108  & n670;
  assign n9738 = ~n9736 & ~n9737;
  assign n9739 = ~n9735 & n9738;
  assign n9740 = n678 & n7170;
  assign n9741 = n9739 & ~n9740;
  assign n9742 = pi11  & ~n9741;
  assign n9743 = pi11  & ~n9742;
  assign n9744 = ~n9741 & ~n9742;
  assign n9745 = ~n9743 & ~n9744;
  assign n9746 = ~n9619 & ~n9623;
  assign n9747 = ~n9602 & ~n9606;
  assign n9748 = ~n9585 & ~n9589;
  assign n9749 = pi100  & n1582;
  assign n9750 = pi98  & n1713;
  assign n9751 = pi99  & n1577;
  assign n9752 = ~n9750 & ~n9751;
  assign n9753 = ~n9749 & n9752;
  assign n9754 = n1585 & n4808;
  assign n9755 = n9753 & ~n9754;
  assign n9756 = pi20  & ~n9755;
  assign n9757 = pi20  & ~n9756;
  assign n9758 = ~n9755 & ~n9756;
  assign n9759 = ~n9757 & ~n9758;
  assign n9760 = ~n9569 & ~n9571;
  assign n9761 = ~n9563 & ~n9565;
  assign n9762 = pi94  & n2486;
  assign n9763 = pi92  & n2644;
  assign n9764 = pi93  & n2481;
  assign n9765 = ~n9763 & ~n9764;
  assign n9766 = ~n9762 & n9765;
  assign n9767 = n2489 & n3499;
  assign n9768 = n9766 & ~n9767;
  assign n9769 = pi26  & ~n9768;
  assign n9770 = pi26  & ~n9769;
  assign n9771 = ~n9768 & ~n9769;
  assign n9772 = ~n9770 & ~n9771;
  assign n9773 = ~n9557 & ~n9559;
  assign n9774 = pi91  & n2976;
  assign n9775 = pi89  & n3182;
  assign n9776 = pi90  & n2971;
  assign n9777 = ~n9775 & ~n9776;
  assign n9778 = ~n9774 & n9777;
  assign n9779 = n2926 & n2979;
  assign n9780 = n9778 & ~n9779;
  assign n9781 = pi29  & ~n9780;
  assign n9782 = pi29  & ~n9781;
  assign n9783 = ~n9780 & ~n9781;
  assign n9784 = ~n9782 & ~n9783;
  assign n9785 = ~n9550 & ~n9553;
  assign n9786 = pi88  & n3550;
  assign n9787 = pi86  & n3735;
  assign n9788 = pi87  & n3545;
  assign n9789 = ~n9787 & ~n9788;
  assign n9790 = ~n9786 & n9789;
  assign n9791 = n2277 & n3553;
  assign n9792 = n9790 & ~n9791;
  assign n9793 = pi32  & ~n9792;
  assign n9794 = pi32  & ~n9793;
  assign n9795 = ~n9792 & ~n9793;
  assign n9796 = ~n9794 & ~n9795;
  assign n9797 = ~n9543 & ~n9547;
  assign n9798 = pi85  & n4182;
  assign n9799 = pi83  & n4416;
  assign n9800 = pi84  & n4177;
  assign n9801 = ~n9799 & ~n9800;
  assign n9802 = ~n9798 & n9801;
  assign n9803 = n1943 & n4185;
  assign n9804 = n9802 & ~n9803;
  assign n9805 = pi35  & ~n9804;
  assign n9806 = pi35  & ~n9805;
  assign n9807 = ~n9804 & ~n9805;
  assign n9808 = ~n9806 & ~n9807;
  assign n9809 = ~n9526 & ~n9529;
  assign n9810 = pi82  & n4896;
  assign n9811 = pi80  & n5148;
  assign n9812 = pi81  & n4891;
  assign n9813 = ~n9811 & ~n9812;
  assign n9814 = ~n9810 & n9813;
  assign n9815 = n1532 & n4899;
  assign n9816 = n9814 & ~n9815;
  assign n9817 = pi38  & ~n9816;
  assign n9818 = pi38  & ~n9817;
  assign n9819 = ~n9816 & ~n9817;
  assign n9820 = ~n9818 & ~n9819;
  assign n9821 = ~n9520 & ~n9523;
  assign n9822 = pi79  & n5636;
  assign n9823 = pi77  & n5909;
  assign n9824 = pi78  & n5631;
  assign n9825 = ~n9823 & ~n9824;
  assign n9826 = ~n9822 & n9825;
  assign n9827 = n1105 & n5639;
  assign n9828 = n9826 & ~n9827;
  assign n9829 = pi41  & ~n9828;
  assign n9830 = pi41  & ~n9829;
  assign n9831 = ~n9828 & ~n9829;
  assign n9832 = ~n9830 & ~n9831;
  assign n9833 = ~n9504 & ~n9506;
  assign n9834 = pi76  & n6396;
  assign n9835 = pi74  & n6735;
  assign n9836 = pi75  & n6391;
  assign n9837 = ~n9835 & ~n9836;
  assign n9838 = ~n9834 & n9837;
  assign n9839 = n881 & n6399;
  assign n9840 = n9838 & ~n9839;
  assign n9841 = pi44  & ~n9840;
  assign n9842 = pi44  & ~n9841;
  assign n9843 = ~n9840 & ~n9841;
  assign n9844 = ~n9842 & ~n9843;
  assign n9845 = ~n9498 & ~n9500;
  assign n9846 = pi73  & n7239;
  assign n9847 = pi71  & n7556;
  assign n9848 = pi72  & n7234;
  assign n9849 = ~n9847 & ~n9848;
  assign n9850 = ~n9846 & n9849;
  assign n9851 = n639 & n7242;
  assign n9852 = n9850 & ~n9851;
  assign n9853 = pi47  & ~n9852;
  assign n9854 = pi47  & ~n9853;
  assign n9855 = ~n9852 & ~n9853;
  assign n9856 = ~n9854 & ~n9855;
  assign n9857 = pi67  & n9096;
  assign n9858 = pi65  & n9453;
  assign n9859 = pi66  & n9091;
  assign n9860 = ~n9858 & ~n9859;
  assign n9861 = ~n9857 & n9860;
  assign n9862 = n313 & n9099;
  assign n9863 = n9861 & ~n9862;
  assign n9864 = pi53  & ~n9863;
  assign n9865 = pi53  & ~n9864;
  assign n9866 = ~n9863 & ~n9864;
  assign n9867 = ~n9865 & ~n9866;
  assign n9868 = pi53  & ~pi54 ;
  assign n9869 = ~pi53  & pi54 ;
  assign n9870 = ~n9868 & ~n9869;
  assign n9871 = pi64  & ~n9870;
  assign n9872 = n9465 & n9871;
  assign n9873 = ~n9465 & ~n9871;
  assign n9874 = ~n9872 & ~n9873;
  assign n9875 = ~n9867 & n9874;
  assign n9876 = n9867 & ~n9874;
  assign n9877 = ~n9875 & ~n9876;
  assign n9878 = pi70  & n8137;
  assign n9879 = pi68  & n8471;
  assign n9880 = pi69  & n8132;
  assign n9881 = ~n9879 & ~n9880;
  assign n9882 = ~n9878 & n9881;
  assign n9883 = n430 & n8140;
  assign n9884 = n9882 & ~n9883;
  assign n9885 = pi50  & ~n9884;
  assign n9886 = pi50  & ~n9885;
  assign n9887 = ~n9884 & ~n9885;
  assign n9888 = ~n9886 & ~n9887;
  assign n9889 = n9877 & ~n9888;
  assign n9890 = ~n9877 & n9888;
  assign n9891 = ~n9889 & ~n9890;
  assign n9892 = ~n9483 & n9891;
  assign n9893 = n9483 & ~n9891;
  assign n9894 = ~n9892 & ~n9893;
  assign n9895 = ~n9856 & n9894;
  assign n9896 = n9856 & ~n9894;
  assign n9897 = ~n9895 & ~n9896;
  assign n9898 = ~n9845 & n9897;
  assign n9899 = n9845 & ~n9897;
  assign n9900 = ~n9898 & ~n9899;
  assign n9901 = ~n9844 & n9900;
  assign n9902 = n9844 & ~n9900;
  assign n9903 = ~n9901 & ~n9902;
  assign n9904 = ~n9833 & n9903;
  assign n9905 = n9833 & ~n9903;
  assign n9906 = ~n9904 & ~n9905;
  assign n9907 = ~n9832 & n9906;
  assign n9908 = n9832 & ~n9906;
  assign n9909 = ~n9907 & ~n9908;
  assign n9910 = ~n9821 & n9909;
  assign n9911 = n9821 & ~n9909;
  assign n9912 = ~n9910 & ~n9911;
  assign n9913 = ~n9820 & n9912;
  assign n9914 = ~n9820 & ~n9913;
  assign n9915 = n9912 & ~n9913;
  assign n9916 = ~n9914 & ~n9915;
  assign n9917 = ~n9809 & ~n9916;
  assign n9918 = n9809 & n9916;
  assign n9919 = ~n9917 & ~n9918;
  assign n9920 = ~n9808 & n9919;
  assign n9921 = n9808 & ~n9919;
  assign n9922 = ~n9920 & ~n9921;
  assign n9923 = ~n9797 & n9922;
  assign n9924 = n9797 & ~n9922;
  assign n9925 = ~n9923 & ~n9924;
  assign n9926 = ~n9796 & n9925;
  assign n9927 = n9796 & ~n9925;
  assign n9928 = ~n9926 & ~n9927;
  assign n9929 = ~n9785 & n9928;
  assign n9930 = n9785 & ~n9928;
  assign n9931 = ~n9929 & ~n9930;
  assign n9932 = ~n9784 & n9931;
  assign n9933 = n9784 & ~n9931;
  assign n9934 = ~n9932 & ~n9933;
  assign n9935 = ~n9773 & n9934;
  assign n9936 = n9773 & ~n9934;
  assign n9937 = ~n9935 & ~n9936;
  assign n9938 = ~n9772 & n9937;
  assign n9939 = n9772 & ~n9937;
  assign n9940 = ~n9938 & ~n9939;
  assign n9941 = ~n9761 & n9940;
  assign n9942 = n9761 & ~n9940;
  assign n9943 = ~n9941 & ~n9942;
  assign n9944 = pi97  & n2004;
  assign n9945 = pi95  & n2141;
  assign n9946 = pi96  & n1999;
  assign n9947 = ~n9945 & ~n9946;
  assign n9948 = ~n9944 & n9947;
  assign n9949 = n2007 & n3946;
  assign n9950 = n9948 & ~n9949;
  assign n9951 = pi23  & ~n9950;
  assign n9952 = pi23  & ~n9951;
  assign n9953 = ~n9950 & ~n9951;
  assign n9954 = ~n9952 & ~n9953;
  assign n9955 = n9943 & ~n9954;
  assign n9956 = ~n9943 & n9954;
  assign n9957 = ~n9955 & ~n9956;
  assign n9958 = ~n9760 & n9957;
  assign n9959 = n9760 & ~n9957;
  assign n9960 = ~n9958 & ~n9959;
  assign n9961 = ~n9759 & n9960;
  assign n9962 = n9759 & ~n9960;
  assign n9963 = ~n9961 & ~n9962;
  assign n9964 = n9748 & ~n9963;
  assign n9965 = ~n9748 & n9963;
  assign n9966 = ~n9964 & ~n9965;
  assign n9967 = pi103  & n1269;
  assign n9968 = pi101  & n1340;
  assign n9969 = pi102  & n1264;
  assign n9970 = ~n9968 & ~n9969;
  assign n9971 = ~n9967 & n9970;
  assign n9972 = n1272 & n5540;
  assign n9973 = n9971 & ~n9972;
  assign n9974 = pi17  & ~n9973;
  assign n9975 = pi17  & ~n9974;
  assign n9976 = ~n9973 & ~n9974;
  assign n9977 = ~n9975 & ~n9976;
  assign n9978 = n9966 & ~n9977;
  assign n9979 = ~n9966 & n9977;
  assign n9980 = ~n9978 & ~n9979;
  assign n9981 = n9747 & ~n9980;
  assign n9982 = ~n9747 & n9980;
  assign n9983 = ~n9981 & ~n9982;
  assign n9984 = pi106  & n918;
  assign n9985 = pi104  & n1031;
  assign n9986 = pi105  & n913;
  assign n9987 = ~n9985 & ~n9986;
  assign n9988 = ~n9984 & n9987;
  assign n9989 = n921 & n6090;
  assign n9990 = n9988 & ~n9989;
  assign n9991 = pi14  & ~n9990;
  assign n9992 = pi14  & ~n9991;
  assign n9993 = ~n9990 & ~n9991;
  assign n9994 = ~n9992 & ~n9993;
  assign n9995 = ~n9983 & n9994;
  assign n9996 = n9983 & ~n9994;
  assign n9997 = ~n9995 & ~n9996;
  assign n9998 = ~n9746 & n9997;
  assign n9999 = n9746 & ~n9997;
  assign n10000 = ~n9998 & ~n9999;
  assign n10001 = ~n9745 & n10000;
  assign n10002 = n9745 & ~n10000;
  assign n10003 = ~n10001 & ~n10002;
  assign n10004 = ~n9641 & n10003;
  assign n10005 = n9641 & ~n10003;
  assign n10006 = ~n10004 & ~n10005;
  assign n10007 = ~n9734 & n10006;
  assign n10008 = n9734 & ~n10006;
  assign n10009 = ~n10007 & ~n10008;
  assign n10010 = n9723 & ~n10009;
  assign n10011 = ~n9723 & n10009;
  assign n10012 = ~n10010 & ~n10011;
  assign n10013 = pi115  & n340;
  assign n10014 = pi113  & n380;
  assign n10015 = pi114  & n335;
  assign n10016 = ~n10014 & ~n10015;
  assign n10017 = ~n10013 & n10016;
  assign n10018 = n343 & n8727;
  assign n10019 = n10017 & ~n10018;
  assign n10020 = pi5  & ~n10019;
  assign n10021 = pi5  & ~n10020;
  assign n10022 = ~n10019 & ~n10020;
  assign n10023 = ~n10021 & ~n10022;
  assign n10024 = ~n10012 & n10023;
  assign n10025 = n10012 & ~n10023;
  assign n10026 = ~n10024 & ~n10025;
  assign n10027 = ~n9677 & n10026;
  assign n10028 = n9677 & ~n10026;
  assign n10029 = ~n10027 & ~n10028;
  assign n10030 = ~n9722 & n10029;
  assign n10031 = n9722 & ~n10029;
  assign n10032 = ~n10030 & ~n10031;
  assign n10033 = ~n9704 & n10032;
  assign n10034 = n9704 & ~n10032;
  assign po54  = ~n10033 & ~n10034;
  assign n10036 = ~n10030 & ~n10033;
  assign n10037 = pi119  & n264;
  assign n10038 = pi117  & n281;
  assign n10039 = pi118  & n259;
  assign n10040 = ~n10038 & ~n10039;
  assign n10041 = ~n10037 & n10040;
  assign n10042 = ~n9712 & ~n9714;
  assign n10043 = ~pi118  & ~pi119 ;
  assign n10044 = pi118  & pi119 ;
  assign n10045 = ~n10043 & ~n10044;
  assign n10046 = ~n10042 & n10045;
  assign n10047 = n10042 & ~n10045;
  assign n10048 = ~n10046 & ~n10047;
  assign n10049 = n267 & n10048;
  assign n10050 = n10041 & ~n10049;
  assign n10051 = pi2  & ~n10050;
  assign n10052 = pi2  & ~n10051;
  assign n10053 = ~n10050 & ~n10051;
  assign n10054 = ~n10052 & ~n10053;
  assign n10055 = ~n10025 & ~n10027;
  assign n10056 = ~n10007 & ~n10011;
  assign n10057 = pi113  & n493;
  assign n10058 = pi111  & n533;
  assign n10059 = pi112  & n488;
  assign n10060 = ~n10058 & ~n10059;
  assign n10061 = ~n10057 & n10060;
  assign n10062 = n496 & n8387;
  assign n10063 = n10061 & ~n10062;
  assign n10064 = pi8  & ~n10063;
  assign n10065 = pi8  & ~n10064;
  assign n10066 = ~n10063 & ~n10064;
  assign n10067 = ~n10065 & ~n10066;
  assign n10068 = ~n10001 & ~n10004;
  assign n10069 = ~n9996 & ~n9998;
  assign n10070 = ~n9978 & ~n9982;
  assign n10071 = ~n9961 & ~n9965;
  assign n10072 = ~n9955 & ~n9958;
  assign n10073 = ~n9938 & ~n9941;
  assign n10074 = ~n9932 & ~n9935;
  assign n10075 = ~n9926 & ~n9929;
  assign n10076 = ~n9920 & ~n9923;
  assign n10077 = ~n9913 & ~n9917;
  assign n10078 = ~n9901 & ~n9904;
  assign n10079 = pi77  & n6396;
  assign n10080 = pi75  & n6735;
  assign n10081 = pi76  & n6391;
  assign n10082 = ~n10080 & ~n10081;
  assign n10083 = ~n10079 & n10082;
  assign n10084 = n984 & n6399;
  assign n10085 = n10083 & ~n10084;
  assign n10086 = pi44  & ~n10085;
  assign n10087 = pi44  & ~n10086;
  assign n10088 = ~n10085 & ~n10086;
  assign n10089 = ~n10087 & ~n10088;
  assign n10090 = ~n9895 & ~n9898;
  assign n10091 = pi74  & n7239;
  assign n10092 = pi72  & n7556;
  assign n10093 = pi73  & n7234;
  assign n10094 = ~n10092 & ~n10093;
  assign n10095 = ~n10091 & n10094;
  assign n10096 = n722 & n7242;
  assign n10097 = n10095 & ~n10096;
  assign n10098 = pi47  & ~n10097;
  assign n10099 = pi47  & ~n10098;
  assign n10100 = ~n10097 & ~n10098;
  assign n10101 = ~n10099 & ~n10100;
  assign n10102 = ~n9889 & ~n9892;
  assign n10103 = pi71  & n8137;
  assign n10104 = pi69  & n8471;
  assign n10105 = pi70  & n8132;
  assign n10106 = ~n10104 & ~n10105;
  assign n10107 = ~n10103 & n10106;
  assign n10108 = n476 & n8140;
  assign n10109 = n10107 & ~n10108;
  assign n10110 = pi50  & ~n10109;
  assign n10111 = pi50  & ~n10110;
  assign n10112 = ~n10109 & ~n10110;
  assign n10113 = ~n10111 & ~n10112;
  assign n10114 = ~n9872 & ~n9875;
  assign n10115 = pi68  & n9096;
  assign n10116 = pi66  & n9453;
  assign n10117 = pi67  & n9091;
  assign n10118 = ~n10116 & ~n10117;
  assign n10119 = ~n10115 & n10118;
  assign n10120 = n364 & n9099;
  assign n10121 = n10119 & ~n10120;
  assign n10122 = pi53  & ~n10121;
  assign n10123 = pi53  & ~n10122;
  assign n10124 = ~n10121 & ~n10122;
  assign n10125 = ~n10123 & ~n10124;
  assign n10126 = pi56  & ~n9871;
  assign n10127 = ~pi54  & pi55 ;
  assign n10128 = pi54  & ~pi55 ;
  assign n10129 = ~n10127 & ~n10128;
  assign n10130 = n9870 & ~n10129;
  assign n10131 = pi64  & n10130;
  assign n10132 = ~pi55  & pi56 ;
  assign n10133 = pi55  & ~pi56 ;
  assign n10134 = ~n10132 & ~n10133;
  assign n10135 = ~n9870 & n10134;
  assign n10136 = pi65  & n10135;
  assign n10137 = ~n10131 & ~n10136;
  assign n10138 = ~n9870 & ~n10134;
  assign n10139 = n270 & n10138;
  assign n10140 = n10137 & ~n10139;
  assign n10141 = pi56  & ~n10140;
  assign n10142 = pi56  & ~n10141;
  assign n10143 = ~n10140 & ~n10141;
  assign n10144 = ~n10142 & ~n10143;
  assign n10145 = n10126 & ~n10144;
  assign n10146 = ~n10126 & n10144;
  assign n10147 = ~n10145 & ~n10146;
  assign n10148 = n10125 & ~n10147;
  assign n10149 = ~n10125 & n10147;
  assign n10150 = ~n10148 & ~n10149;
  assign n10151 = ~n10114 & n10150;
  assign n10152 = n10114 & ~n10150;
  assign n10153 = ~n10151 & ~n10152;
  assign n10154 = n10113 & ~n10153;
  assign n10155 = ~n10113 & n10153;
  assign n10156 = ~n10154 & ~n10155;
  assign n10157 = ~n10102 & n10156;
  assign n10158 = n10102 & ~n10156;
  assign n10159 = ~n10157 & ~n10158;
  assign n10160 = n10101 & ~n10159;
  assign n10161 = ~n10101 & n10159;
  assign n10162 = ~n10160 & ~n10161;
  assign n10163 = ~n10090 & n10162;
  assign n10164 = n10090 & ~n10162;
  assign n10165 = ~n10163 & ~n10164;
  assign n10166 = n10089 & ~n10165;
  assign n10167 = ~n10089 & n10165;
  assign n10168 = ~n10166 & ~n10167;
  assign n10169 = ~n10078 & n10168;
  assign n10170 = n10078 & ~n10168;
  assign n10171 = ~n10169 & ~n10170;
  assign n10172 = pi80  & n5636;
  assign n10173 = pi78  & n5909;
  assign n10174 = pi79  & n5631;
  assign n10175 = ~n10173 & ~n10174;
  assign n10176 = ~n10172 & n10175;
  assign n10177 = n1205 & n5639;
  assign n10178 = n10176 & ~n10177;
  assign n10179 = pi41  & ~n10178;
  assign n10180 = pi41  & ~n10179;
  assign n10181 = ~n10178 & ~n10179;
  assign n10182 = ~n10180 & ~n10181;
  assign n10183 = n10171 & ~n10182;
  assign n10184 = n10171 & ~n10183;
  assign n10185 = ~n10182 & ~n10183;
  assign n10186 = ~n10184 & ~n10185;
  assign n10187 = ~n9907 & ~n9910;
  assign n10188 = n10186 & n10187;
  assign n10189 = ~n10186 & ~n10187;
  assign n10190 = ~n10188 & ~n10189;
  assign n10191 = pi83  & n4896;
  assign n10192 = pi81  & n5148;
  assign n10193 = pi82  & n4891;
  assign n10194 = ~n10192 & ~n10193;
  assign n10195 = ~n10191 & n10194;
  assign n10196 = n1672 & n4899;
  assign n10197 = n10195 & ~n10196;
  assign n10198 = pi38  & ~n10197;
  assign n10199 = pi38  & ~n10198;
  assign n10200 = ~n10197 & ~n10198;
  assign n10201 = ~n10199 & ~n10200;
  assign n10202 = n10190 & ~n10201;
  assign n10203 = ~n10190 & n10201;
  assign n10204 = ~n10077 & ~n10203;
  assign n10205 = ~n10202 & n10204;
  assign n10206 = ~n10077 & ~n10205;
  assign n10207 = ~n10202 & ~n10205;
  assign n10208 = ~n10203 & n10207;
  assign n10209 = ~n10206 & ~n10208;
  assign n10210 = pi86  & n4182;
  assign n10211 = pi84  & n4416;
  assign n10212 = pi85  & n4177;
  assign n10213 = ~n10211 & ~n10212;
  assign n10214 = ~n10210 & n10213;
  assign n10215 = n2099 & n4185;
  assign n10216 = n10214 & ~n10215;
  assign n10217 = pi35  & ~n10216;
  assign n10218 = pi35  & ~n10217;
  assign n10219 = ~n10216 & ~n10217;
  assign n10220 = ~n10218 & ~n10219;
  assign n10221 = ~n10209 & ~n10220;
  assign n10222 = n10209 & n10220;
  assign n10223 = ~n10221 & ~n10222;
  assign n10224 = n10076 & ~n10223;
  assign n10225 = ~n10076 & n10223;
  assign n10226 = ~n10224 & ~n10225;
  assign n10227 = pi89  & n3550;
  assign n10228 = pi87  & n3735;
  assign n10229 = pi88  & n3545;
  assign n10230 = ~n10228 & ~n10229;
  assign n10231 = ~n10227 & n10230;
  assign n10232 = n2432 & n3553;
  assign n10233 = n10231 & ~n10232;
  assign n10234 = pi32  & ~n10233;
  assign n10235 = pi32  & ~n10234;
  assign n10236 = ~n10233 & ~n10234;
  assign n10237 = ~n10235 & ~n10236;
  assign n10238 = n10226 & ~n10237;
  assign n10239 = ~n10226 & n10237;
  assign n10240 = ~n10238 & ~n10239;
  assign n10241 = n10075 & ~n10240;
  assign n10242 = ~n10075 & n10240;
  assign n10243 = ~n10241 & ~n10242;
  assign n10244 = pi92  & n2976;
  assign n10245 = pi90  & n3182;
  assign n10246 = pi91  & n2971;
  assign n10247 = ~n10245 & ~n10246;
  assign n10248 = ~n10244 & n10247;
  assign n10249 = n2979 & n3119;
  assign n10250 = n10248 & ~n10249;
  assign n10251 = pi29  & ~n10250;
  assign n10252 = pi29  & ~n10251;
  assign n10253 = ~n10250 & ~n10251;
  assign n10254 = ~n10252 & ~n10253;
  assign n10255 = n10243 & ~n10254;
  assign n10256 = ~n10243 & n10254;
  assign n10257 = ~n10255 & ~n10256;
  assign n10258 = n10074 & ~n10257;
  assign n10259 = ~n10074 & n10257;
  assign n10260 = ~n10258 & ~n10259;
  assign n10261 = pi95  & n2486;
  assign n10262 = pi93  & n2644;
  assign n10263 = pi94  & n2481;
  assign n10264 = ~n10262 & ~n10263;
  assign n10265 = ~n10261 & n10264;
  assign n10266 = n2489 & n3710;
  assign n10267 = n10265 & ~n10266;
  assign n10268 = pi26  & ~n10267;
  assign n10269 = pi26  & ~n10268;
  assign n10270 = ~n10267 & ~n10268;
  assign n10271 = ~n10269 & ~n10270;
  assign n10272 = n10260 & ~n10271;
  assign n10273 = ~n10260 & n10271;
  assign n10274 = ~n10272 & ~n10273;
  assign n10275 = n10073 & ~n10274;
  assign n10276 = ~n10073 & n10274;
  assign n10277 = ~n10275 & ~n10276;
  assign n10278 = pi98  & n2004;
  assign n10279 = pi96  & n2141;
  assign n10280 = pi97  & n1999;
  assign n10281 = ~n10279 & ~n10280;
  assign n10282 = ~n10278 & n10281;
  assign n10283 = n2007 & n4360;
  assign n10284 = n10282 & ~n10283;
  assign n10285 = pi23  & ~n10284;
  assign n10286 = pi23  & ~n10285;
  assign n10287 = ~n10284 & ~n10285;
  assign n10288 = ~n10286 & ~n10287;
  assign n10289 = n10277 & ~n10288;
  assign n10290 = ~n10277 & n10288;
  assign n10291 = ~n10289 & ~n10290;
  assign n10292 = n10072 & ~n10291;
  assign n10293 = ~n10072 & n10291;
  assign n10294 = ~n10292 & ~n10293;
  assign n10295 = pi101  & n1582;
  assign n10296 = pi99  & n1713;
  assign n10297 = pi100  & n1577;
  assign n10298 = ~n10296 & ~n10297;
  assign n10299 = ~n10295 & n10298;
  assign n10300 = n1585 & n5056;
  assign n10301 = n10299 & ~n10300;
  assign n10302 = pi20  & ~n10301;
  assign n10303 = pi20  & ~n10302;
  assign n10304 = ~n10301 & ~n10302;
  assign n10305 = ~n10303 & ~n10304;
  assign n10306 = n10294 & ~n10305;
  assign n10307 = ~n10294 & n10305;
  assign n10308 = ~n10306 & ~n10307;
  assign n10309 = n10071 & ~n10308;
  assign n10310 = ~n10071 & n10308;
  assign n10311 = ~n10309 & ~n10310;
  assign n10312 = pi104  & n1269;
  assign n10313 = pi102  & n1340;
  assign n10314 = pi103  & n1264;
  assign n10315 = ~n10313 & ~n10314;
  assign n10316 = ~n10312 & n10315;
  assign n10317 = n1272 & n5565;
  assign n10318 = n10316 & ~n10317;
  assign n10319 = pi17  & ~n10318;
  assign n10320 = pi17  & ~n10319;
  assign n10321 = ~n10318 & ~n10319;
  assign n10322 = ~n10320 & ~n10321;
  assign n10323 = n10311 & ~n10322;
  assign n10324 = ~n10311 & n10322;
  assign n10325 = ~n10323 & ~n10324;
  assign n10326 = n10070 & ~n10325;
  assign n10327 = ~n10070 & n10325;
  assign n10328 = ~n10326 & ~n10327;
  assign n10329 = pi107  & n918;
  assign n10330 = pi105  & n1031;
  assign n10331 = pi106  & n913;
  assign n10332 = ~n10330 & ~n10331;
  assign n10333 = ~n10329 & n10332;
  assign n10334 = n921 & n6614;
  assign n10335 = n10333 & ~n10334;
  assign n10336 = pi14  & ~n10335;
  assign n10337 = pi14  & ~n10336;
  assign n10338 = ~n10335 & ~n10336;
  assign n10339 = ~n10337 & ~n10338;
  assign n10340 = n10328 & ~n10339;
  assign n10341 = ~n10328 & n10339;
  assign n10342 = ~n10069 & ~n10341;
  assign n10343 = ~n10340 & n10342;
  assign n10344 = ~n10069 & ~n10343;
  assign n10345 = ~n10340 & ~n10343;
  assign n10346 = ~n10341 & n10345;
  assign n10347 = ~n10344 & ~n10346;
  assign n10348 = pi110  & n675;
  assign n10349 = pi108  & n769;
  assign n10350 = pi109  & n670;
  assign n10351 = ~n10349 & ~n10350;
  assign n10352 = ~n10348 & n10351;
  assign n10353 = n678 & n7474;
  assign n10354 = n10352 & ~n10353;
  assign n10355 = pi11  & ~n10354;
  assign n10356 = pi11  & ~n10355;
  assign n10357 = ~n10354 & ~n10355;
  assign n10358 = ~n10356 & ~n10357;
  assign n10359 = n10347 & n10358;
  assign n10360 = ~n10347 & ~n10358;
  assign n10361 = ~n10359 & ~n10360;
  assign n10362 = ~n10068 & n10361;
  assign n10363 = n10068 & ~n10361;
  assign n10364 = ~n10362 & ~n10363;
  assign n10365 = n10067 & ~n10364;
  assign n10366 = ~n10067 & n10364;
  assign n10367 = ~n10365 & ~n10366;
  assign n10368 = ~n10056 & n10367;
  assign n10369 = n10056 & ~n10367;
  assign n10370 = ~n10368 & ~n10369;
  assign n10371 = pi116  & n340;
  assign n10372 = pi114  & n380;
  assign n10373 = pi115  & n335;
  assign n10374 = ~n10372 & ~n10373;
  assign n10375 = ~n10371 & n10374;
  assign n10376 = n343 & n9042;
  assign n10377 = n10375 & ~n10376;
  assign n10378 = pi5  & ~n10377;
  assign n10379 = pi5  & ~n10378;
  assign n10380 = ~n10377 & ~n10378;
  assign n10381 = ~n10379 & ~n10380;
  assign n10382 = n10370 & ~n10381;
  assign n10383 = ~n10370 & n10381;
  assign n10384 = ~n10382 & ~n10383;
  assign n10385 = ~n10055 & n10384;
  assign n10386 = n10055 & ~n10384;
  assign n10387 = ~n10385 & ~n10386;
  assign n10388 = ~n10054 & n10387;
  assign n10389 = n10054 & ~n10387;
  assign n10390 = ~n10388 & ~n10389;
  assign n10391 = ~n10036 & n10390;
  assign n10392 = n10036 & ~n10390;
  assign po55  = ~n10391 & ~n10392;
  assign n10394 = ~n10388 & ~n10391;
  assign n10395 = ~n10382 & ~n10385;
  assign n10396 = pi117  & n340;
  assign n10397 = pi115  & n380;
  assign n10398 = pi116  & n335;
  assign n10399 = ~n10397 & ~n10398;
  assign n10400 = ~n10396 & n10399;
  assign n10401 = n343 & n9691;
  assign n10402 = n10400 & ~n10401;
  assign n10403 = pi5  & ~n10402;
  assign n10404 = pi5  & ~n10403;
  assign n10405 = ~n10402 & ~n10403;
  assign n10406 = ~n10404 & ~n10405;
  assign n10407 = ~n10366 & ~n10368;
  assign n10408 = pi114  & n493;
  assign n10409 = pi112  & n533;
  assign n10410 = pi113  & n488;
  assign n10411 = ~n10409 & ~n10410;
  assign n10412 = ~n10408 & n10411;
  assign n10413 = n496 & n8702;
  assign n10414 = n10412 & ~n10413;
  assign n10415 = pi8  & ~n10414;
  assign n10416 = pi8  & ~n10415;
  assign n10417 = ~n10414 & ~n10415;
  assign n10418 = ~n10416 & ~n10417;
  assign n10419 = ~n10360 & ~n10362;
  assign n10420 = ~n10323 & ~n10327;
  assign n10421 = ~n10306 & ~n10310;
  assign n10422 = ~n10289 & ~n10293;
  assign n10423 = ~n10272 & ~n10276;
  assign n10424 = pi96  & n2486;
  assign n10425 = pi94  & n2644;
  assign n10426 = pi95  & n2481;
  assign n10427 = ~n10425 & ~n10426;
  assign n10428 = ~n10424 & n10427;
  assign n10429 = n2489 & n3921;
  assign n10430 = n10428 & ~n10429;
  assign n10431 = pi26  & ~n10430;
  assign n10432 = pi26  & ~n10431;
  assign n10433 = ~n10430 & ~n10431;
  assign n10434 = ~n10432 & ~n10433;
  assign n10435 = ~n10255 & ~n10259;
  assign n10436 = ~n10238 & ~n10242;
  assign n10437 = ~n10221 & ~n10225;
  assign n10438 = pi87  & n4182;
  assign n10439 = pi85  & n4416;
  assign n10440 = pi86  & n4177;
  assign n10441 = ~n10439 & ~n10440;
  assign n10442 = ~n10438 & n10441;
  assign n10443 = n2252 & n4185;
  assign n10444 = n10442 & ~n10443;
  assign n10445 = pi35  & ~n10444;
  assign n10446 = pi35  & ~n10445;
  assign n10447 = ~n10444 & ~n10445;
  assign n10448 = ~n10446 & ~n10447;
  assign n10449 = ~n10183 & ~n10189;
  assign n10450 = pi81  & n5636;
  assign n10451 = pi79  & n5909;
  assign n10452 = pi80  & n5631;
  assign n10453 = ~n10451 & ~n10452;
  assign n10454 = ~n10450 & n10453;
  assign n10455 = n1413 & n5639;
  assign n10456 = n10454 & ~n10455;
  assign n10457 = pi41  & ~n10456;
  assign n10458 = pi41  & ~n10457;
  assign n10459 = ~n10456 & ~n10457;
  assign n10460 = ~n10458 & ~n10459;
  assign n10461 = ~n10167 & ~n10169;
  assign n10462 = ~n10161 & ~n10163;
  assign n10463 = pi75  & n7239;
  assign n10464 = pi73  & n7556;
  assign n10465 = pi74  & n7234;
  assign n10466 = ~n10464 & ~n10465;
  assign n10467 = ~n10463 & n10466;
  assign n10468 = n747 & n7242;
  assign n10469 = n10467 & ~n10468;
  assign n10470 = pi47  & ~n10469;
  assign n10471 = pi47  & ~n10470;
  assign n10472 = ~n10469 & ~n10470;
  assign n10473 = ~n10471 & ~n10472;
  assign n10474 = ~n10155 & ~n10157;
  assign n10475 = ~n10149 & ~n10151;
  assign n10476 = pi66  & n10135;
  assign n10477 = n9870 & ~n10134;
  assign n10478 = n10129 & n10477;
  assign n10479 = pi64  & n10478;
  assign n10480 = pi65  & n10130;
  assign n10481 = ~n10479 & ~n10480;
  assign n10482 = ~n10476 & n10481;
  assign n10483 = n291 & n10138;
  assign n10484 = n10482 & ~n10483;
  assign n10485 = pi56  & ~n10484;
  assign n10486 = pi56  & ~n10485;
  assign n10487 = ~n10484 & ~n10485;
  assign n10488 = ~n10486 & ~n10487;
  assign n10489 = ~n10145 & n10488;
  assign n10490 = n10145 & ~n10488;
  assign n10491 = ~n10489 & ~n10490;
  assign n10492 = pi69  & n9096;
  assign n10493 = pi67  & n9453;
  assign n10494 = pi68  & n9091;
  assign n10495 = ~n10493 & ~n10494;
  assign n10496 = ~n10492 & n10495;
  assign n10497 = n405 & n9099;
  assign n10498 = n10496 & ~n10497;
  assign n10499 = pi53  & ~n10498;
  assign n10500 = pi53  & ~n10499;
  assign n10501 = ~n10498 & ~n10499;
  assign n10502 = ~n10500 & ~n10501;
  assign n10503 = n10491 & ~n10502;
  assign n10504 = ~n10491 & n10502;
  assign n10505 = ~n10475 & ~n10504;
  assign n10506 = ~n10503 & n10505;
  assign n10507 = ~n10475 & ~n10506;
  assign n10508 = ~n10503 & ~n10506;
  assign n10509 = ~n10504 & n10508;
  assign n10510 = ~n10507 & ~n10509;
  assign n10511 = pi72  & n8137;
  assign n10512 = pi70  & n8471;
  assign n10513 = pi71  & n8132;
  assign n10514 = ~n10512 & ~n10513;
  assign n10515 = ~n10511 & n10514;
  assign n10516 = n575 & n8140;
  assign n10517 = n10515 & ~n10516;
  assign n10518 = pi50  & ~n10517;
  assign n10519 = pi50  & ~n10518;
  assign n10520 = ~n10517 & ~n10518;
  assign n10521 = ~n10519 & ~n10520;
  assign n10522 = n10510 & n10521;
  assign n10523 = ~n10510 & ~n10521;
  assign n10524 = ~n10522 & ~n10523;
  assign n10525 = ~n10474 & n10524;
  assign n10526 = n10474 & ~n10524;
  assign n10527 = ~n10525 & ~n10526;
  assign n10528 = n10473 & ~n10527;
  assign n10529 = ~n10473 & n10527;
  assign n10530 = ~n10528 & ~n10529;
  assign n10531 = ~n10462 & n10530;
  assign n10532 = n10462 & ~n10530;
  assign n10533 = ~n10531 & ~n10532;
  assign n10534 = pi78  & n6396;
  assign n10535 = pi76  & n6735;
  assign n10536 = pi77  & n6391;
  assign n10537 = ~n10535 & ~n10536;
  assign n10538 = ~n10534 & n10537;
  assign n10539 = n1009 & n6399;
  assign n10540 = n10538 & ~n10539;
  assign n10541 = pi44  & ~n10540;
  assign n10542 = pi44  & ~n10541;
  assign n10543 = ~n10540 & ~n10541;
  assign n10544 = ~n10542 & ~n10543;
  assign n10545 = n10533 & ~n10544;
  assign n10546 = n10533 & ~n10545;
  assign n10547 = ~n10544 & ~n10545;
  assign n10548 = ~n10546 & ~n10547;
  assign n10549 = ~n10461 & ~n10548;
  assign n10550 = n10461 & n10548;
  assign n10551 = ~n10549 & ~n10550;
  assign n10552 = ~n10460 & n10551;
  assign n10553 = n10460 & ~n10551;
  assign n10554 = ~n10552 & ~n10553;
  assign n10555 = ~n10449 & n10554;
  assign n10556 = n10449 & ~n10554;
  assign n10557 = ~n10555 & ~n10556;
  assign n10558 = pi84  & n4896;
  assign n10559 = pi82  & n5148;
  assign n10560 = pi83  & n4891;
  assign n10561 = ~n10559 & ~n10560;
  assign n10562 = ~n10558 & n10561;
  assign n10563 = n1805 & n4899;
  assign n10564 = n10562 & ~n10563;
  assign n10565 = pi38  & ~n10564;
  assign n10566 = pi38  & ~n10565;
  assign n10567 = ~n10564 & ~n10565;
  assign n10568 = ~n10566 & ~n10567;
  assign n10569 = n10557 & ~n10568;
  assign n10570 = n10557 & ~n10569;
  assign n10571 = ~n10568 & ~n10569;
  assign n10572 = ~n10570 & ~n10571;
  assign n10573 = ~n10207 & ~n10572;
  assign n10574 = n10207 & n10572;
  assign n10575 = ~n10573 & ~n10574;
  assign n10576 = ~n10448 & n10575;
  assign n10577 = n10448 & ~n10575;
  assign n10578 = ~n10576 & ~n10577;
  assign n10579 = n10437 & ~n10578;
  assign n10580 = ~n10437 & n10578;
  assign n10581 = ~n10579 & ~n10580;
  assign n10582 = pi90  & n3550;
  assign n10583 = pi88  & n3735;
  assign n10584 = pi89  & n3545;
  assign n10585 = ~n10583 & ~n10584;
  assign n10586 = ~n10582 & n10585;
  assign n10587 = n2606 & n3553;
  assign n10588 = n10586 & ~n10587;
  assign n10589 = pi32  & ~n10588;
  assign n10590 = pi32  & ~n10589;
  assign n10591 = ~n10588 & ~n10589;
  assign n10592 = ~n10590 & ~n10591;
  assign n10593 = n10581 & ~n10592;
  assign n10594 = ~n10581 & n10592;
  assign n10595 = ~n10436 & ~n10594;
  assign n10596 = ~n10593 & n10595;
  assign n10597 = ~n10436 & ~n10596;
  assign n10598 = ~n10593 & ~n10596;
  assign n10599 = ~n10594 & n10598;
  assign n10600 = ~n10597 & ~n10599;
  assign n10601 = pi93  & n2976;
  assign n10602 = pi91  & n3182;
  assign n10603 = pi92  & n2971;
  assign n10604 = ~n10602 & ~n10603;
  assign n10605 = ~n10601 & n10604;
  assign n10606 = n2979 & n3144;
  assign n10607 = n10605 & ~n10606;
  assign n10608 = pi29  & ~n10607;
  assign n10609 = pi29  & ~n10608;
  assign n10610 = ~n10607 & ~n10608;
  assign n10611 = ~n10609 & ~n10610;
  assign n10612 = n10600 & n10611;
  assign n10613 = ~n10600 & ~n10611;
  assign n10614 = ~n10612 & ~n10613;
  assign n10615 = ~n10435 & n10614;
  assign n10616 = n10435 & ~n10614;
  assign n10617 = ~n10615 & ~n10616;
  assign n10618 = n10434 & ~n10617;
  assign n10619 = ~n10434 & n10617;
  assign n10620 = ~n10618 & ~n10619;
  assign n10621 = ~n10423 & n10620;
  assign n10622 = n10423 & ~n10620;
  assign n10623 = ~n10621 & ~n10622;
  assign n10624 = pi99  & n2004;
  assign n10625 = pi97  & n2141;
  assign n10626 = pi98  & n1999;
  assign n10627 = ~n10625 & ~n10626;
  assign n10628 = ~n10624 & n10627;
  assign n10629 = n2007 & n4584;
  assign n10630 = n10628 & ~n10629;
  assign n10631 = pi23  & ~n10630;
  assign n10632 = pi23  & ~n10631;
  assign n10633 = ~n10630 & ~n10631;
  assign n10634 = ~n10632 & ~n10633;
  assign n10635 = n10623 & ~n10634;
  assign n10636 = ~n10623 & n10634;
  assign n10637 = ~n10635 & ~n10636;
  assign n10638 = n10422 & ~n10637;
  assign n10639 = ~n10422 & n10637;
  assign n10640 = ~n10638 & ~n10639;
  assign n10641 = pi102  & n1582;
  assign n10642 = pi100  & n1713;
  assign n10643 = pi101  & n1577;
  assign n10644 = ~n10642 & ~n10643;
  assign n10645 = ~n10641 & n10644;
  assign n10646 = n1585 & n5296;
  assign n10647 = n10645 & ~n10646;
  assign n10648 = pi20  & ~n10647;
  assign n10649 = pi20  & ~n10648;
  assign n10650 = ~n10647 & ~n10648;
  assign n10651 = ~n10649 & ~n10650;
  assign n10652 = n10640 & ~n10651;
  assign n10653 = ~n10640 & n10651;
  assign n10654 = ~n10652 & ~n10653;
  assign n10655 = n10421 & ~n10654;
  assign n10656 = ~n10421 & n10654;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = pi105  & n1269;
  assign n10659 = pi103  & n1340;
  assign n10660 = pi104  & n1264;
  assign n10661 = ~n10659 & ~n10660;
  assign n10662 = ~n10658 & n10661;
  assign n10663 = n1272 & n6065;
  assign n10664 = n10662 & ~n10663;
  assign n10665 = pi17  & ~n10664;
  assign n10666 = pi17  & ~n10665;
  assign n10667 = ~n10664 & ~n10665;
  assign n10668 = ~n10666 & ~n10667;
  assign n10669 = n10657 & ~n10668;
  assign n10670 = ~n10657 & n10668;
  assign n10671 = ~n10669 & ~n10670;
  assign n10672 = n10420 & ~n10671;
  assign n10673 = ~n10420 & n10671;
  assign n10674 = ~n10672 & ~n10673;
  assign n10675 = pi108  & n918;
  assign n10676 = pi106  & n1031;
  assign n10677 = pi107  & n913;
  assign n10678 = ~n10676 & ~n10677;
  assign n10679 = ~n10675 & n10678;
  assign n10680 = n921 & n6639;
  assign n10681 = n10679 & ~n10680;
  assign n10682 = pi14  & ~n10681;
  assign n10683 = pi14  & ~n10682;
  assign n10684 = ~n10681 & ~n10682;
  assign n10685 = ~n10683 & ~n10684;
  assign n10686 = n10674 & ~n10685;
  assign n10687 = ~n10674 & n10685;
  assign n10688 = ~n10345 & ~n10687;
  assign n10689 = ~n10686 & n10688;
  assign n10690 = ~n10345 & ~n10689;
  assign n10691 = ~n10686 & ~n10689;
  assign n10692 = ~n10687 & n10691;
  assign n10693 = ~n10690 & ~n10692;
  assign n10694 = pi111  & n675;
  assign n10695 = pi109  & n769;
  assign n10696 = pi110  & n670;
  assign n10697 = ~n10695 & ~n10696;
  assign n10698 = ~n10694 & n10697;
  assign n10699 = n678 & n7770;
  assign n10700 = n10698 & ~n10699;
  assign n10701 = pi11  & ~n10700;
  assign n10702 = pi11  & ~n10701;
  assign n10703 = ~n10700 & ~n10701;
  assign n10704 = ~n10702 & ~n10703;
  assign n10705 = ~n10693 & ~n10704;
  assign n10706 = n10693 & n10704;
  assign n10707 = ~n10705 & ~n10706;
  assign n10708 = ~n10419 & n10707;
  assign n10709 = n10419 & ~n10707;
  assign n10710 = ~n10708 & ~n10709;
  assign n10711 = ~n10418 & n10710;
  assign n10712 = n10418 & ~n10710;
  assign n10713 = ~n10711 & ~n10712;
  assign n10714 = ~n10407 & n10713;
  assign n10715 = n10407 & ~n10713;
  assign n10716 = ~n10714 & ~n10715;
  assign n10717 = n10406 & ~n10716;
  assign n10718 = ~n10406 & n10716;
  assign n10719 = ~n10717 & ~n10718;
  assign n10720 = ~n10395 & n10719;
  assign n10721 = n10395 & ~n10719;
  assign n10722 = ~n10720 & ~n10721;
  assign n10723 = pi120  & n264;
  assign n10724 = pi118  & n281;
  assign n10725 = pi119  & n259;
  assign n10726 = ~n10724 & ~n10725;
  assign n10727 = ~n10723 & n10726;
  assign n10728 = ~n10044 & ~n10046;
  assign n10729 = ~pi119  & ~pi120 ;
  assign n10730 = pi119  & pi120 ;
  assign n10731 = ~n10729 & ~n10730;
  assign n10732 = ~n10728 & n10731;
  assign n10733 = n10728 & ~n10731;
  assign n10734 = ~n10732 & ~n10733;
  assign n10735 = n267 & n10734;
  assign n10736 = n10727 & ~n10735;
  assign n10737 = pi2  & ~n10736;
  assign n10738 = pi2  & ~n10737;
  assign n10739 = ~n10736 & ~n10737;
  assign n10740 = ~n10738 & ~n10739;
  assign n10741 = n10722 & ~n10740;
  assign n10742 = ~n10722 & n10740;
  assign n10743 = ~n10741 & ~n10742;
  assign n10744 = ~n10394 & n10743;
  assign n10745 = n10394 & ~n10743;
  assign po56  = ~n10744 & ~n10745;
  assign n10747 = ~n10741 & ~n10744;
  assign n10748 = ~n10718 & ~n10720;
  assign n10749 = pi118  & n340;
  assign n10750 = pi116  & n380;
  assign n10751 = pi117  & n335;
  assign n10752 = ~n10750 & ~n10751;
  assign n10753 = ~n10749 & n10752;
  assign n10754 = n343 & n9716;
  assign n10755 = n10753 & ~n10754;
  assign n10756 = pi5  & ~n10755;
  assign n10757 = pi5  & ~n10756;
  assign n10758 = ~n10755 & ~n10756;
  assign n10759 = ~n10757 & ~n10758;
  assign n10760 = ~n10711 & ~n10714;
  assign n10761 = pi115  & n493;
  assign n10762 = pi113  & n533;
  assign n10763 = pi114  & n488;
  assign n10764 = ~n10762 & ~n10763;
  assign n10765 = ~n10761 & n10764;
  assign n10766 = n496 & n8727;
  assign n10767 = n10765 & ~n10766;
  assign n10768 = pi8  & ~n10767;
  assign n10769 = pi8  & ~n10768;
  assign n10770 = ~n10767 & ~n10768;
  assign n10771 = ~n10769 & ~n10770;
  assign n10772 = ~n10705 & ~n10708;
  assign n10773 = pi112  & n675;
  assign n10774 = pi110  & n769;
  assign n10775 = pi111  & n670;
  assign n10776 = ~n10774 & ~n10775;
  assign n10777 = ~n10773 & n10776;
  assign n10778 = n678 & n7795;
  assign n10779 = n10777 & ~n10778;
  assign n10780 = pi11  & ~n10779;
  assign n10781 = pi11  & ~n10780;
  assign n10782 = ~n10779 & ~n10780;
  assign n10783 = ~n10781 & ~n10782;
  assign n10784 = pi109  & n918;
  assign n10785 = pi107  & n1031;
  assign n10786 = pi108  & n913;
  assign n10787 = ~n10785 & ~n10786;
  assign n10788 = ~n10784 & n10787;
  assign n10789 = n921 & n7170;
  assign n10790 = n10788 & ~n10789;
  assign n10791 = pi14  & ~n10790;
  assign n10792 = pi14  & ~n10791;
  assign n10793 = ~n10790 & ~n10791;
  assign n10794 = ~n10792 & ~n10793;
  assign n10795 = ~n10669 & ~n10673;
  assign n10796 = ~n10652 & ~n10656;
  assign n10797 = ~n10635 & ~n10639;
  assign n10798 = pi100  & n2004;
  assign n10799 = pi98  & n2141;
  assign n10800 = pi99  & n1999;
  assign n10801 = ~n10799 & ~n10800;
  assign n10802 = ~n10798 & n10801;
  assign n10803 = n2007 & n4808;
  assign n10804 = n10802 & ~n10803;
  assign n10805 = pi23  & ~n10804;
  assign n10806 = pi23  & ~n10805;
  assign n10807 = ~n10804 & ~n10805;
  assign n10808 = ~n10806 & ~n10807;
  assign n10809 = ~n10619 & ~n10621;
  assign n10810 = ~n10613 & ~n10615;
  assign n10811 = pi94  & n2976;
  assign n10812 = pi92  & n3182;
  assign n10813 = pi93  & n2971;
  assign n10814 = ~n10812 & ~n10813;
  assign n10815 = ~n10811 & n10814;
  assign n10816 = n2979 & n3499;
  assign n10817 = n10815 & ~n10816;
  assign n10818 = pi29  & ~n10817;
  assign n10819 = pi29  & ~n10818;
  assign n10820 = ~n10817 & ~n10818;
  assign n10821 = ~n10819 & ~n10820;
  assign n10822 = ~n10569 & ~n10573;
  assign n10823 = pi85  & n4896;
  assign n10824 = pi83  & n5148;
  assign n10825 = pi84  & n4891;
  assign n10826 = ~n10824 & ~n10825;
  assign n10827 = ~n10823 & n10826;
  assign n10828 = n1943 & n4899;
  assign n10829 = n10827 & ~n10828;
  assign n10830 = pi38  & ~n10829;
  assign n10831 = pi38  & ~n10830;
  assign n10832 = ~n10829 & ~n10830;
  assign n10833 = ~n10831 & ~n10832;
  assign n10834 = ~n10552 & ~n10555;
  assign n10835 = pi82  & n5636;
  assign n10836 = pi80  & n5909;
  assign n10837 = pi81  & n5631;
  assign n10838 = ~n10836 & ~n10837;
  assign n10839 = ~n10835 & n10838;
  assign n10840 = n1532 & n5639;
  assign n10841 = n10839 & ~n10840;
  assign n10842 = pi41  & ~n10841;
  assign n10843 = pi41  & ~n10842;
  assign n10844 = ~n10841 & ~n10842;
  assign n10845 = ~n10843 & ~n10844;
  assign n10846 = ~n10545 & ~n10549;
  assign n10847 = pi79  & n6396;
  assign n10848 = pi77  & n6735;
  assign n10849 = pi78  & n6391;
  assign n10850 = ~n10848 & ~n10849;
  assign n10851 = ~n10847 & n10850;
  assign n10852 = n1105 & n6399;
  assign n10853 = n10851 & ~n10852;
  assign n10854 = pi44  & ~n10853;
  assign n10855 = pi44  & ~n10854;
  assign n10856 = ~n10853 & ~n10854;
  assign n10857 = ~n10855 & ~n10856;
  assign n10858 = ~n10529 & ~n10531;
  assign n10859 = pi76  & n7239;
  assign n10860 = pi74  & n7556;
  assign n10861 = pi75  & n7234;
  assign n10862 = ~n10860 & ~n10861;
  assign n10863 = ~n10859 & n10862;
  assign n10864 = n881 & n7242;
  assign n10865 = n10863 & ~n10864;
  assign n10866 = pi47  & ~n10865;
  assign n10867 = pi47  & ~n10866;
  assign n10868 = ~n10865 & ~n10866;
  assign n10869 = ~n10867 & ~n10868;
  assign n10870 = ~n10523 & ~n10525;
  assign n10871 = pi73  & n8137;
  assign n10872 = pi71  & n8471;
  assign n10873 = pi72  & n8132;
  assign n10874 = ~n10872 & ~n10873;
  assign n10875 = ~n10871 & n10874;
  assign n10876 = n639 & n8140;
  assign n10877 = n10875 & ~n10876;
  assign n10878 = pi50  & ~n10877;
  assign n10879 = pi50  & ~n10878;
  assign n10880 = ~n10877 & ~n10878;
  assign n10881 = ~n10879 & ~n10880;
  assign n10882 = pi67  & n10135;
  assign n10883 = pi65  & n10478;
  assign n10884 = pi66  & n10130;
  assign n10885 = ~n10883 & ~n10884;
  assign n10886 = ~n10882 & n10885;
  assign n10887 = n313 & n10138;
  assign n10888 = n10886 & ~n10887;
  assign n10889 = pi56  & ~n10888;
  assign n10890 = pi56  & ~n10889;
  assign n10891 = ~n10888 & ~n10889;
  assign n10892 = ~n10890 & ~n10891;
  assign n10893 = pi56  & ~pi57 ;
  assign n10894 = ~pi56  & pi57 ;
  assign n10895 = ~n10893 & ~n10894;
  assign n10896 = pi64  & ~n10895;
  assign n10897 = n10490 & n10896;
  assign n10898 = ~n10490 & ~n10896;
  assign n10899 = ~n10897 & ~n10898;
  assign n10900 = ~n10892 & n10899;
  assign n10901 = n10892 & ~n10899;
  assign n10902 = ~n10900 & ~n10901;
  assign n10903 = pi70  & n9096;
  assign n10904 = pi68  & n9453;
  assign n10905 = pi69  & n9091;
  assign n10906 = ~n10904 & ~n10905;
  assign n10907 = ~n10903 & n10906;
  assign n10908 = n430 & n9099;
  assign n10909 = n10907 & ~n10908;
  assign n10910 = pi53  & ~n10909;
  assign n10911 = pi53  & ~n10910;
  assign n10912 = ~n10909 & ~n10910;
  assign n10913 = ~n10911 & ~n10912;
  assign n10914 = n10902 & ~n10913;
  assign n10915 = ~n10902 & n10913;
  assign n10916 = ~n10914 & ~n10915;
  assign n10917 = ~n10508 & n10916;
  assign n10918 = n10508 & ~n10916;
  assign n10919 = ~n10917 & ~n10918;
  assign n10920 = ~n10881 & n10919;
  assign n10921 = n10881 & ~n10919;
  assign n10922 = ~n10920 & ~n10921;
  assign n10923 = ~n10870 & n10922;
  assign n10924 = n10870 & ~n10922;
  assign n10925 = ~n10923 & ~n10924;
  assign n10926 = n10869 & ~n10925;
  assign n10927 = ~n10869 & n10925;
  assign n10928 = ~n10926 & ~n10927;
  assign n10929 = ~n10858 & n10928;
  assign n10930 = n10858 & ~n10928;
  assign n10931 = ~n10929 & ~n10930;
  assign n10932 = ~n10857 & n10931;
  assign n10933 = n10857 & ~n10931;
  assign n10934 = ~n10932 & ~n10933;
  assign n10935 = ~n10846 & n10934;
  assign n10936 = n10846 & ~n10934;
  assign n10937 = ~n10935 & ~n10936;
  assign n10938 = ~n10845 & n10937;
  assign n10939 = ~n10845 & ~n10938;
  assign n10940 = n10937 & ~n10938;
  assign n10941 = ~n10939 & ~n10940;
  assign n10942 = ~n10834 & ~n10941;
  assign n10943 = n10834 & n10941;
  assign n10944 = ~n10942 & ~n10943;
  assign n10945 = ~n10833 & n10944;
  assign n10946 = n10833 & ~n10944;
  assign n10947 = ~n10945 & ~n10946;
  assign n10948 = ~n10822 & n10947;
  assign n10949 = n10822 & ~n10947;
  assign n10950 = ~n10948 & ~n10949;
  assign n10951 = pi88  & n4182;
  assign n10952 = pi86  & n4416;
  assign n10953 = pi87  & n4177;
  assign n10954 = ~n10952 & ~n10953;
  assign n10955 = ~n10951 & n10954;
  assign n10956 = n2277 & n4185;
  assign n10957 = n10955 & ~n10956;
  assign n10958 = pi35  & ~n10957;
  assign n10959 = pi35  & ~n10958;
  assign n10960 = ~n10957 & ~n10958;
  assign n10961 = ~n10959 & ~n10960;
  assign n10962 = n10950 & ~n10961;
  assign n10963 = n10950 & ~n10962;
  assign n10964 = ~n10961 & ~n10962;
  assign n10965 = ~n10963 & ~n10964;
  assign n10966 = ~n10576 & ~n10580;
  assign n10967 = n10965 & n10966;
  assign n10968 = ~n10965 & ~n10966;
  assign n10969 = ~n10967 & ~n10968;
  assign n10970 = pi91  & n3550;
  assign n10971 = pi89  & n3735;
  assign n10972 = pi90  & n3545;
  assign n10973 = ~n10971 & ~n10972;
  assign n10974 = ~n10970 & n10973;
  assign n10975 = n2926 & n3553;
  assign n10976 = n10974 & ~n10975;
  assign n10977 = pi32  & ~n10976;
  assign n10978 = pi32  & ~n10977;
  assign n10979 = ~n10976 & ~n10977;
  assign n10980 = ~n10978 & ~n10979;
  assign n10981 = ~n10969 & n10980;
  assign n10982 = n10969 & ~n10980;
  assign n10983 = ~n10981 & ~n10982;
  assign n10984 = ~n10598 & n10983;
  assign n10985 = n10598 & ~n10983;
  assign n10986 = ~n10984 & ~n10985;
  assign n10987 = ~n10821 & n10986;
  assign n10988 = n10821 & ~n10986;
  assign n10989 = ~n10987 & ~n10988;
  assign n10990 = ~n10810 & n10989;
  assign n10991 = n10810 & ~n10989;
  assign n10992 = ~n10990 & ~n10991;
  assign n10993 = pi97  & n2486;
  assign n10994 = pi95  & n2644;
  assign n10995 = pi96  & n2481;
  assign n10996 = ~n10994 & ~n10995;
  assign n10997 = ~n10993 & n10996;
  assign n10998 = n2489 & n3946;
  assign n10999 = n10997 & ~n10998;
  assign n11000 = pi26  & ~n10999;
  assign n11001 = pi26  & ~n11000;
  assign n11002 = ~n10999 & ~n11000;
  assign n11003 = ~n11001 & ~n11002;
  assign n11004 = n10992 & ~n11003;
  assign n11005 = ~n10992 & n11003;
  assign n11006 = ~n11004 & ~n11005;
  assign n11007 = ~n10809 & n11006;
  assign n11008 = n10809 & ~n11006;
  assign n11009 = ~n11007 & ~n11008;
  assign n11010 = ~n10808 & n11009;
  assign n11011 = n10808 & ~n11009;
  assign n11012 = ~n11010 & ~n11011;
  assign n11013 = n10797 & ~n11012;
  assign n11014 = ~n10797 & n11012;
  assign n11015 = ~n11013 & ~n11014;
  assign n11016 = pi103  & n1582;
  assign n11017 = pi101  & n1713;
  assign n11018 = pi102  & n1577;
  assign n11019 = ~n11017 & ~n11018;
  assign n11020 = ~n11016 & n11019;
  assign n11021 = n1585 & n5540;
  assign n11022 = n11020 & ~n11021;
  assign n11023 = pi20  & ~n11022;
  assign n11024 = pi20  & ~n11023;
  assign n11025 = ~n11022 & ~n11023;
  assign n11026 = ~n11024 & ~n11025;
  assign n11027 = n11015 & ~n11026;
  assign n11028 = ~n11015 & n11026;
  assign n11029 = ~n11027 & ~n11028;
  assign n11030 = n10796 & ~n11029;
  assign n11031 = ~n10796 & n11029;
  assign n11032 = ~n11030 & ~n11031;
  assign n11033 = pi106  & n1269;
  assign n11034 = pi104  & n1340;
  assign n11035 = pi105  & n1264;
  assign n11036 = ~n11034 & ~n11035;
  assign n11037 = ~n11033 & n11036;
  assign n11038 = n1272 & n6090;
  assign n11039 = n11037 & ~n11038;
  assign n11040 = pi17  & ~n11039;
  assign n11041 = pi17  & ~n11040;
  assign n11042 = ~n11039 & ~n11040;
  assign n11043 = ~n11041 & ~n11042;
  assign n11044 = ~n11032 & n11043;
  assign n11045 = n11032 & ~n11043;
  assign n11046 = ~n11044 & ~n11045;
  assign n11047 = ~n10795 & n11046;
  assign n11048 = n10795 & ~n11046;
  assign n11049 = ~n11047 & ~n11048;
  assign n11050 = ~n10794 & n11049;
  assign n11051 = n10794 & ~n11049;
  assign n11052 = ~n11050 & ~n11051;
  assign n11053 = ~n10691 & n11052;
  assign n11054 = n10691 & ~n11052;
  assign n11055 = ~n11053 & ~n11054;
  assign n11056 = ~n10783 & n11055;
  assign n11057 = n10783 & ~n11055;
  assign n11058 = ~n11056 & ~n11057;
  assign n11059 = ~n10772 & n11058;
  assign n11060 = n10772 & ~n11058;
  assign n11061 = ~n11059 & ~n11060;
  assign n11062 = ~n10771 & n11061;
  assign n11063 = n10771 & ~n11061;
  assign n11064 = ~n11062 & ~n11063;
  assign n11065 = ~n10760 & n11064;
  assign n11066 = n10760 & ~n11064;
  assign n11067 = ~n11065 & ~n11066;
  assign n11068 = ~n10759 & n11067;
  assign n11069 = ~n10759 & ~n11068;
  assign n11070 = n11067 & ~n11068;
  assign n11071 = ~n11069 & ~n11070;
  assign n11072 = ~n10748 & ~n11071;
  assign n11073 = n10748 & n11071;
  assign n11074 = ~n11072 & ~n11073;
  assign n11075 = pi121  & n264;
  assign n11076 = pi119  & n281;
  assign n11077 = pi120  & n259;
  assign n11078 = ~n11076 & ~n11077;
  assign n11079 = ~n11075 & n11078;
  assign n11080 = ~n10730 & ~n10732;
  assign n11081 = ~pi120  & ~pi121 ;
  assign n11082 = pi120  & pi121 ;
  assign n11083 = ~n11081 & ~n11082;
  assign n11084 = ~n11080 & n11083;
  assign n11085 = n11080 & ~n11083;
  assign n11086 = ~n11084 & ~n11085;
  assign n11087 = n267 & n11086;
  assign n11088 = n11079 & ~n11087;
  assign n11089 = pi2  & ~n11088;
  assign n11090 = pi2  & ~n11089;
  assign n11091 = ~n11088 & ~n11089;
  assign n11092 = ~n11090 & ~n11091;
  assign n11093 = n11074 & ~n11092;
  assign n11094 = ~n11074 & n11092;
  assign n11095 = ~n11093 & ~n11094;
  assign n11096 = ~n10747 & n11095;
  assign n11097 = n10747 & ~n11095;
  assign po57  = ~n11096 & ~n11097;
  assign n11099 = ~n11093 & ~n11096;
  assign n11100 = ~n11068 & ~n11072;
  assign n11101 = pi119  & n340;
  assign n11102 = pi117  & n380;
  assign n11103 = pi118  & n335;
  assign n11104 = ~n11102 & ~n11103;
  assign n11105 = ~n11101 & n11104;
  assign n11106 = n343 & n10048;
  assign n11107 = n11105 & ~n11106;
  assign n11108 = pi5  & ~n11107;
  assign n11109 = pi5  & ~n11108;
  assign n11110 = ~n11107 & ~n11108;
  assign n11111 = ~n11109 & ~n11110;
  assign n11112 = ~n11062 & ~n11065;
  assign n11113 = pi116  & n493;
  assign n11114 = pi114  & n533;
  assign n11115 = pi115  & n488;
  assign n11116 = ~n11114 & ~n11115;
  assign n11117 = ~n11113 & n11116;
  assign n11118 = n496 & n9042;
  assign n11119 = n11117 & ~n11118;
  assign n11120 = pi8  & ~n11119;
  assign n11121 = pi8  & ~n11120;
  assign n11122 = ~n11119 & ~n11120;
  assign n11123 = ~n11121 & ~n11122;
  assign n11124 = ~n11056 & ~n11059;
  assign n11125 = pi113  & n675;
  assign n11126 = pi111  & n769;
  assign n11127 = pi112  & n670;
  assign n11128 = ~n11126 & ~n11127;
  assign n11129 = ~n11125 & n11128;
  assign n11130 = n678 & n8387;
  assign n11131 = n11129 & ~n11130;
  assign n11132 = pi11  & ~n11131;
  assign n11133 = pi11  & ~n11132;
  assign n11134 = ~n11131 & ~n11132;
  assign n11135 = ~n11133 & ~n11134;
  assign n11136 = ~n11050 & ~n11053;
  assign n11137 = ~n11045 & ~n11047;
  assign n11138 = ~n11027 & ~n11031;
  assign n11139 = ~n11010 & ~n11014;
  assign n11140 = ~n11004 & ~n11007;
  assign n11141 = ~n10987 & ~n10990;
  assign n11142 = pi95  & n2976;
  assign n11143 = pi93  & n3182;
  assign n11144 = pi94  & n2971;
  assign n11145 = ~n11143 & ~n11144;
  assign n11146 = ~n11142 & n11145;
  assign n11147 = n2979 & n3710;
  assign n11148 = n11146 & ~n11147;
  assign n11149 = pi29  & ~n11148;
  assign n11150 = pi29  & ~n11149;
  assign n11151 = ~n11148 & ~n11149;
  assign n11152 = ~n11150 & ~n11151;
  assign n11153 = ~n10982 & ~n10984;
  assign n11154 = ~n10962 & ~n10968;
  assign n11155 = ~n10945 & ~n10948;
  assign n11156 = ~n10938 & ~n10942;
  assign n11157 = ~n10932 & ~n10935;
  assign n11158 = ~n10927 & ~n10929;
  assign n11159 = ~n10920 & ~n10923;
  assign n11160 = ~n10914 & ~n10917;
  assign n11161 = pi71  & n9096;
  assign n11162 = pi69  & n9453;
  assign n11163 = pi70  & n9091;
  assign n11164 = ~n11162 & ~n11163;
  assign n11165 = ~n11161 & n11164;
  assign n11166 = n476 & n9099;
  assign n11167 = n11165 & ~n11166;
  assign n11168 = pi53  & ~n11167;
  assign n11169 = pi53  & ~n11168;
  assign n11170 = ~n11167 & ~n11168;
  assign n11171 = ~n11169 & ~n11170;
  assign n11172 = ~n10897 & ~n10900;
  assign n11173 = pi68  & n10135;
  assign n11174 = pi66  & n10478;
  assign n11175 = pi67  & n10130;
  assign n11176 = ~n11174 & ~n11175;
  assign n11177 = ~n11173 & n11176;
  assign n11178 = n364 & n10138;
  assign n11179 = n11177 & ~n11178;
  assign n11180 = pi56  & ~n11179;
  assign n11181 = pi56  & ~n11180;
  assign n11182 = ~n11179 & ~n11180;
  assign n11183 = ~n11181 & ~n11182;
  assign n11184 = pi59  & ~n10896;
  assign n11185 = ~pi57  & pi58 ;
  assign n11186 = pi57  & ~pi58 ;
  assign n11187 = ~n11185 & ~n11186;
  assign n11188 = n10895 & ~n11187;
  assign n11189 = pi64  & n11188;
  assign n11190 = ~pi58  & pi59 ;
  assign n11191 = pi58  & ~pi59 ;
  assign n11192 = ~n11190 & ~n11191;
  assign n11193 = ~n10895 & n11192;
  assign n11194 = pi65  & n11193;
  assign n11195 = ~n11189 & ~n11194;
  assign n11196 = ~n10895 & ~n11192;
  assign n11197 = n270 & n11196;
  assign n11198 = n11195 & ~n11197;
  assign n11199 = pi59  & ~n11198;
  assign n11200 = pi59  & ~n11199;
  assign n11201 = ~n11198 & ~n11199;
  assign n11202 = ~n11200 & ~n11201;
  assign n11203 = n11184 & ~n11202;
  assign n11204 = ~n11184 & n11202;
  assign n11205 = ~n11203 & ~n11204;
  assign n11206 = n11183 & ~n11205;
  assign n11207 = ~n11183 & n11205;
  assign n11208 = ~n11206 & ~n11207;
  assign n11209 = ~n11172 & n11208;
  assign n11210 = n11172 & ~n11208;
  assign n11211 = ~n11209 & ~n11210;
  assign n11212 = n11171 & ~n11211;
  assign n11213 = ~n11171 & n11211;
  assign n11214 = ~n11212 & ~n11213;
  assign n11215 = ~n11160 & n11214;
  assign n11216 = n11160 & ~n11214;
  assign n11217 = ~n11215 & ~n11216;
  assign n11218 = pi74  & n8137;
  assign n11219 = pi72  & n8471;
  assign n11220 = pi73  & n8132;
  assign n11221 = ~n11219 & ~n11220;
  assign n11222 = ~n11218 & n11221;
  assign n11223 = n722 & n8140;
  assign n11224 = n11222 & ~n11223;
  assign n11225 = pi50  & ~n11224;
  assign n11226 = pi50  & ~n11225;
  assign n11227 = ~n11224 & ~n11225;
  assign n11228 = ~n11226 & ~n11227;
  assign n11229 = n11217 & ~n11228;
  assign n11230 = ~n11217 & n11228;
  assign n11231 = ~n11229 & ~n11230;
  assign n11232 = n11159 & ~n11231;
  assign n11233 = ~n11159 & n11231;
  assign n11234 = ~n11232 & ~n11233;
  assign n11235 = pi77  & n7239;
  assign n11236 = pi75  & n7556;
  assign n11237 = pi76  & n7234;
  assign n11238 = ~n11236 & ~n11237;
  assign n11239 = ~n11235 & n11238;
  assign n11240 = n984 & n7242;
  assign n11241 = n11239 & ~n11240;
  assign n11242 = pi47  & ~n11241;
  assign n11243 = pi47  & ~n11242;
  assign n11244 = ~n11241 & ~n11242;
  assign n11245 = ~n11243 & ~n11244;
  assign n11246 = n11234 & ~n11245;
  assign n11247 = ~n11234 & n11245;
  assign n11248 = ~n11158 & ~n11247;
  assign n11249 = ~n11246 & n11248;
  assign n11250 = ~n11158 & ~n11249;
  assign n11251 = ~n11246 & ~n11249;
  assign n11252 = ~n11247 & n11251;
  assign n11253 = ~n11250 & ~n11252;
  assign n11254 = pi80  & n6396;
  assign n11255 = pi78  & n6735;
  assign n11256 = pi79  & n6391;
  assign n11257 = ~n11255 & ~n11256;
  assign n11258 = ~n11254 & n11257;
  assign n11259 = n1205 & n6399;
  assign n11260 = n11258 & ~n11259;
  assign n11261 = pi44  & ~n11260;
  assign n11262 = pi44  & ~n11261;
  assign n11263 = ~n11260 & ~n11261;
  assign n11264 = ~n11262 & ~n11263;
  assign n11265 = ~n11253 & ~n11264;
  assign n11266 = n11253 & n11264;
  assign n11267 = ~n11265 & ~n11266;
  assign n11268 = n11157 & ~n11267;
  assign n11269 = ~n11157 & n11267;
  assign n11270 = ~n11268 & ~n11269;
  assign n11271 = pi83  & n5636;
  assign n11272 = pi81  & n5909;
  assign n11273 = pi82  & n5631;
  assign n11274 = ~n11272 & ~n11273;
  assign n11275 = ~n11271 & n11274;
  assign n11276 = n1672 & n5639;
  assign n11277 = n11275 & ~n11276;
  assign n11278 = pi41  & ~n11277;
  assign n11279 = pi41  & ~n11278;
  assign n11280 = ~n11277 & ~n11278;
  assign n11281 = ~n11279 & ~n11280;
  assign n11282 = n11270 & ~n11281;
  assign n11283 = ~n11270 & n11281;
  assign n11284 = ~n11156 & ~n11283;
  assign n11285 = ~n11282 & n11284;
  assign n11286 = ~n11156 & ~n11285;
  assign n11287 = ~n11282 & ~n11285;
  assign n11288 = ~n11283 & n11287;
  assign n11289 = ~n11286 & ~n11288;
  assign n11290 = pi86  & n4896;
  assign n11291 = pi84  & n5148;
  assign n11292 = pi85  & n4891;
  assign n11293 = ~n11291 & ~n11292;
  assign n11294 = ~n11290 & n11293;
  assign n11295 = n2099 & n4899;
  assign n11296 = n11294 & ~n11295;
  assign n11297 = pi38  & ~n11296;
  assign n11298 = pi38  & ~n11297;
  assign n11299 = ~n11296 & ~n11297;
  assign n11300 = ~n11298 & ~n11299;
  assign n11301 = ~n11289 & ~n11300;
  assign n11302 = n11289 & n11300;
  assign n11303 = ~n11301 & ~n11302;
  assign n11304 = n11155 & ~n11303;
  assign n11305 = ~n11155 & n11303;
  assign n11306 = ~n11304 & ~n11305;
  assign n11307 = pi89  & n4182;
  assign n11308 = pi87  & n4416;
  assign n11309 = pi88  & n4177;
  assign n11310 = ~n11308 & ~n11309;
  assign n11311 = ~n11307 & n11310;
  assign n11312 = n2432 & n4185;
  assign n11313 = n11311 & ~n11312;
  assign n11314 = pi35  & ~n11313;
  assign n11315 = pi35  & ~n11314;
  assign n11316 = ~n11313 & ~n11314;
  assign n11317 = ~n11315 & ~n11316;
  assign n11318 = n11306 & ~n11317;
  assign n11319 = ~n11306 & n11317;
  assign n11320 = ~n11318 & ~n11319;
  assign n11321 = n11154 & ~n11320;
  assign n11322 = ~n11154 & n11320;
  assign n11323 = ~n11321 & ~n11322;
  assign n11324 = pi92  & n3550;
  assign n11325 = pi90  & n3735;
  assign n11326 = pi91  & n3545;
  assign n11327 = ~n11325 & ~n11326;
  assign n11328 = ~n11324 & n11327;
  assign n11329 = n3119 & n3553;
  assign n11330 = n11328 & ~n11329;
  assign n11331 = pi32  & ~n11330;
  assign n11332 = pi32  & ~n11331;
  assign n11333 = ~n11330 & ~n11331;
  assign n11334 = ~n11332 & ~n11333;
  assign n11335 = n11323 & ~n11334;
  assign n11336 = ~n11323 & n11334;
  assign n11337 = ~n11335 & ~n11336;
  assign n11338 = ~n11153 & n11337;
  assign n11339 = n11153 & ~n11337;
  assign n11340 = ~n11338 & ~n11339;
  assign n11341 = ~n11152 & n11340;
  assign n11342 = n11152 & ~n11340;
  assign n11343 = ~n11341 & ~n11342;
  assign n11344 = n11141 & ~n11343;
  assign n11345 = ~n11141 & n11343;
  assign n11346 = ~n11344 & ~n11345;
  assign n11347 = pi98  & n2486;
  assign n11348 = pi96  & n2644;
  assign n11349 = pi97  & n2481;
  assign n11350 = ~n11348 & ~n11349;
  assign n11351 = ~n11347 & n11350;
  assign n11352 = n2489 & n4360;
  assign n11353 = n11351 & ~n11352;
  assign n11354 = pi26  & ~n11353;
  assign n11355 = pi26  & ~n11354;
  assign n11356 = ~n11353 & ~n11354;
  assign n11357 = ~n11355 & ~n11356;
  assign n11358 = n11346 & ~n11357;
  assign n11359 = ~n11346 & n11357;
  assign n11360 = ~n11358 & ~n11359;
  assign n11361 = n11140 & ~n11360;
  assign n11362 = ~n11140 & n11360;
  assign n11363 = ~n11361 & ~n11362;
  assign n11364 = pi101  & n2004;
  assign n11365 = pi99  & n2141;
  assign n11366 = pi100  & n1999;
  assign n11367 = ~n11365 & ~n11366;
  assign n11368 = ~n11364 & n11367;
  assign n11369 = n2007 & n5056;
  assign n11370 = n11368 & ~n11369;
  assign n11371 = pi23  & ~n11370;
  assign n11372 = pi23  & ~n11371;
  assign n11373 = ~n11370 & ~n11371;
  assign n11374 = ~n11372 & ~n11373;
  assign n11375 = n11363 & ~n11374;
  assign n11376 = ~n11363 & n11374;
  assign n11377 = ~n11375 & ~n11376;
  assign n11378 = n11139 & ~n11377;
  assign n11379 = ~n11139 & n11377;
  assign n11380 = ~n11378 & ~n11379;
  assign n11381 = pi104  & n1582;
  assign n11382 = pi102  & n1713;
  assign n11383 = pi103  & n1577;
  assign n11384 = ~n11382 & ~n11383;
  assign n11385 = ~n11381 & n11384;
  assign n11386 = n1585 & n5565;
  assign n11387 = n11385 & ~n11386;
  assign n11388 = pi20  & ~n11387;
  assign n11389 = pi20  & ~n11388;
  assign n11390 = ~n11387 & ~n11388;
  assign n11391 = ~n11389 & ~n11390;
  assign n11392 = n11380 & ~n11391;
  assign n11393 = ~n11380 & n11391;
  assign n11394 = ~n11392 & ~n11393;
  assign n11395 = n11138 & ~n11394;
  assign n11396 = ~n11138 & n11394;
  assign n11397 = ~n11395 & ~n11396;
  assign n11398 = pi107  & n1269;
  assign n11399 = pi105  & n1340;
  assign n11400 = pi106  & n1264;
  assign n11401 = ~n11399 & ~n11400;
  assign n11402 = ~n11398 & n11401;
  assign n11403 = n1272 & n6614;
  assign n11404 = n11402 & ~n11403;
  assign n11405 = pi17  & ~n11404;
  assign n11406 = pi17  & ~n11405;
  assign n11407 = ~n11404 & ~n11405;
  assign n11408 = ~n11406 & ~n11407;
  assign n11409 = n11397 & ~n11408;
  assign n11410 = ~n11397 & n11408;
  assign n11411 = ~n11137 & ~n11410;
  assign n11412 = ~n11409 & n11411;
  assign n11413 = ~n11137 & ~n11412;
  assign n11414 = ~n11409 & ~n11412;
  assign n11415 = ~n11410 & n11414;
  assign n11416 = ~n11413 & ~n11415;
  assign n11417 = pi110  & n918;
  assign n11418 = pi108  & n1031;
  assign n11419 = pi109  & n913;
  assign n11420 = ~n11418 & ~n11419;
  assign n11421 = ~n11417 & n11420;
  assign n11422 = n921 & n7474;
  assign n11423 = n11421 & ~n11422;
  assign n11424 = pi14  & ~n11423;
  assign n11425 = pi14  & ~n11424;
  assign n11426 = ~n11423 & ~n11424;
  assign n11427 = ~n11425 & ~n11426;
  assign n11428 = n11416 & n11427;
  assign n11429 = ~n11416 & ~n11427;
  assign n11430 = ~n11428 & ~n11429;
  assign n11431 = ~n11136 & n11430;
  assign n11432 = n11136 & ~n11430;
  assign n11433 = ~n11431 & ~n11432;
  assign n11434 = n11135 & ~n11433;
  assign n11435 = ~n11135 & n11433;
  assign n11436 = ~n11434 & ~n11435;
  assign n11437 = ~n11124 & n11436;
  assign n11438 = n11124 & ~n11436;
  assign n11439 = ~n11437 & ~n11438;
  assign n11440 = n11123 & ~n11439;
  assign n11441 = ~n11123 & n11439;
  assign n11442 = ~n11440 & ~n11441;
  assign n11443 = ~n11112 & n11442;
  assign n11444 = n11112 & ~n11442;
  assign n11445 = ~n11443 & ~n11444;
  assign n11446 = n11111 & ~n11445;
  assign n11447 = ~n11111 & n11445;
  assign n11448 = ~n11446 & ~n11447;
  assign n11449 = ~n11100 & n11448;
  assign n11450 = n11100 & ~n11448;
  assign n11451 = ~n11449 & ~n11450;
  assign n11452 = pi122  & n264;
  assign n11453 = pi120  & n281;
  assign n11454 = pi121  & n259;
  assign n11455 = ~n11453 & ~n11454;
  assign n11456 = ~n11452 & n11455;
  assign n11457 = ~n11082 & ~n11084;
  assign n11458 = ~pi121  & ~pi122 ;
  assign n11459 = pi121  & pi122 ;
  assign n11460 = ~n11458 & ~n11459;
  assign n11461 = ~n11457 & n11460;
  assign n11462 = n11457 & ~n11460;
  assign n11463 = ~n11461 & ~n11462;
  assign n11464 = n267 & n11463;
  assign n11465 = n11456 & ~n11464;
  assign n11466 = pi2  & ~n11465;
  assign n11467 = pi2  & ~n11466;
  assign n11468 = ~n11465 & ~n11466;
  assign n11469 = ~n11467 & ~n11468;
  assign n11470 = n11451 & ~n11469;
  assign n11471 = ~n11451 & n11469;
  assign n11472 = ~n11470 & ~n11471;
  assign n11473 = ~n11099 & n11472;
  assign n11474 = n11099 & ~n11472;
  assign po58  = ~n11473 & ~n11474;
  assign n11476 = ~n11470 & ~n11473;
  assign n11477 = ~n11447 & ~n11449;
  assign n11478 = pi123  & n264;
  assign n11479 = pi121  & n281;
  assign n11480 = pi122  & n259;
  assign n11481 = ~n11479 & ~n11480;
  assign n11482 = ~n11478 & n11481;
  assign n11483 = ~n11459 & ~n11461;
  assign n11484 = ~pi122  & ~pi123 ;
  assign n11485 = pi122  & pi123 ;
  assign n11486 = ~n11484 & ~n11485;
  assign n11487 = ~n11483 & n11486;
  assign n11488 = n11483 & ~n11486;
  assign n11489 = ~n11487 & ~n11488;
  assign n11490 = n267 & n11489;
  assign n11491 = n11482 & ~n11490;
  assign n11492 = pi2  & ~n11491;
  assign n11493 = pi2  & ~n11492;
  assign n11494 = ~n11491 & ~n11492;
  assign n11495 = ~n11493 & ~n11494;
  assign n11496 = pi120  & n340;
  assign n11497 = pi118  & n380;
  assign n11498 = pi119  & n335;
  assign n11499 = ~n11497 & ~n11498;
  assign n11500 = ~n11496 & n11499;
  assign n11501 = n343 & n10734;
  assign n11502 = n11500 & ~n11501;
  assign n11503 = pi5  & ~n11502;
  assign n11504 = pi5  & ~n11503;
  assign n11505 = ~n11502 & ~n11503;
  assign n11506 = ~n11504 & ~n11505;
  assign n11507 = ~n11441 & ~n11443;
  assign n11508 = pi117  & n493;
  assign n11509 = pi115  & n533;
  assign n11510 = pi116  & n488;
  assign n11511 = ~n11509 & ~n11510;
  assign n11512 = ~n11508 & n11511;
  assign n11513 = n496 & n9691;
  assign n11514 = n11512 & ~n11513;
  assign n11515 = pi8  & ~n11514;
  assign n11516 = pi8  & ~n11515;
  assign n11517 = ~n11514 & ~n11515;
  assign n11518 = ~n11516 & ~n11517;
  assign n11519 = ~n11435 & ~n11437;
  assign n11520 = ~n11429 & ~n11431;
  assign n11521 = ~n11392 & ~n11396;
  assign n11522 = ~n11375 & ~n11379;
  assign n11523 = ~n11358 & ~n11362;
  assign n11524 = ~n11341 & ~n11345;
  assign n11525 = ~n11335 & ~n11338;
  assign n11526 = ~n11318 & ~n11322;
  assign n11527 = ~n11301 & ~n11305;
  assign n11528 = pi84  & n5636;
  assign n11529 = pi82  & n5909;
  assign n11530 = pi83  & n5631;
  assign n11531 = ~n11529 & ~n11530;
  assign n11532 = ~n11528 & n11531;
  assign n11533 = n1805 & n5639;
  assign n11534 = n11532 & ~n11533;
  assign n11535 = pi41  & ~n11534;
  assign n11536 = pi41  & ~n11535;
  assign n11537 = ~n11534 & ~n11535;
  assign n11538 = ~n11536 & ~n11537;
  assign n11539 = ~n11265 & ~n11269;
  assign n11540 = pi81  & n6396;
  assign n11541 = pi79  & n6735;
  assign n11542 = pi80  & n6391;
  assign n11543 = ~n11541 & ~n11542;
  assign n11544 = ~n11540 & n11543;
  assign n11545 = n1413 & n6399;
  assign n11546 = n11544 & ~n11545;
  assign n11547 = pi44  & ~n11546;
  assign n11548 = pi44  & ~n11547;
  assign n11549 = ~n11546 & ~n11547;
  assign n11550 = ~n11548 & ~n11549;
  assign n11551 = ~n11229 & ~n11233;
  assign n11552 = pi75  & n8137;
  assign n11553 = pi73  & n8471;
  assign n11554 = pi74  & n8132;
  assign n11555 = ~n11553 & ~n11554;
  assign n11556 = ~n11552 & n11555;
  assign n11557 = n747 & n8140;
  assign n11558 = n11556 & ~n11557;
  assign n11559 = pi50  & ~n11558;
  assign n11560 = pi50  & ~n11559;
  assign n11561 = ~n11558 & ~n11559;
  assign n11562 = ~n11560 & ~n11561;
  assign n11563 = ~n11213 & ~n11215;
  assign n11564 = ~n11207 & ~n11209;
  assign n11565 = pi66  & n11193;
  assign n11566 = n10895 & ~n11192;
  assign n11567 = n11187 & n11566;
  assign n11568 = pi64  & n11567;
  assign n11569 = pi65  & n11188;
  assign n11570 = ~n11568 & ~n11569;
  assign n11571 = ~n11565 & n11570;
  assign n11572 = n291 & n11196;
  assign n11573 = n11571 & ~n11572;
  assign n11574 = pi59  & ~n11573;
  assign n11575 = pi59  & ~n11574;
  assign n11576 = ~n11573 & ~n11574;
  assign n11577 = ~n11575 & ~n11576;
  assign n11578 = ~n11203 & n11577;
  assign n11579 = n11203 & ~n11577;
  assign n11580 = ~n11578 & ~n11579;
  assign n11581 = pi69  & n10135;
  assign n11582 = pi67  & n10478;
  assign n11583 = pi68  & n10130;
  assign n11584 = ~n11582 & ~n11583;
  assign n11585 = ~n11581 & n11584;
  assign n11586 = n405 & n10138;
  assign n11587 = n11585 & ~n11586;
  assign n11588 = pi56  & ~n11587;
  assign n11589 = pi56  & ~n11588;
  assign n11590 = ~n11587 & ~n11588;
  assign n11591 = ~n11589 & ~n11590;
  assign n11592 = n11580 & ~n11591;
  assign n11593 = ~n11580 & n11591;
  assign n11594 = ~n11564 & ~n11593;
  assign n11595 = ~n11592 & n11594;
  assign n11596 = ~n11564 & ~n11595;
  assign n11597 = ~n11592 & ~n11595;
  assign n11598 = ~n11593 & n11597;
  assign n11599 = ~n11596 & ~n11598;
  assign n11600 = pi72  & n9096;
  assign n11601 = pi70  & n9453;
  assign n11602 = pi71  & n9091;
  assign n11603 = ~n11601 & ~n11602;
  assign n11604 = ~n11600 & n11603;
  assign n11605 = n575 & n9099;
  assign n11606 = n11604 & ~n11605;
  assign n11607 = pi53  & ~n11606;
  assign n11608 = pi53  & ~n11607;
  assign n11609 = ~n11606 & ~n11607;
  assign n11610 = ~n11608 & ~n11609;
  assign n11611 = n11599 & n11610;
  assign n11612 = ~n11599 & ~n11610;
  assign n11613 = ~n11611 & ~n11612;
  assign n11614 = ~n11563 & n11613;
  assign n11615 = n11563 & ~n11613;
  assign n11616 = ~n11614 & ~n11615;
  assign n11617 = n11562 & ~n11616;
  assign n11618 = ~n11562 & n11616;
  assign n11619 = ~n11617 & ~n11618;
  assign n11620 = ~n11551 & n11619;
  assign n11621 = n11551 & ~n11619;
  assign n11622 = ~n11620 & ~n11621;
  assign n11623 = pi78  & n7239;
  assign n11624 = pi76  & n7556;
  assign n11625 = pi77  & n7234;
  assign n11626 = ~n11624 & ~n11625;
  assign n11627 = ~n11623 & n11626;
  assign n11628 = n1009 & n7242;
  assign n11629 = n11627 & ~n11628;
  assign n11630 = pi47  & ~n11629;
  assign n11631 = pi47  & ~n11630;
  assign n11632 = ~n11629 & ~n11630;
  assign n11633 = ~n11631 & ~n11632;
  assign n11634 = n11622 & ~n11633;
  assign n11635 = n11622 & ~n11634;
  assign n11636 = ~n11633 & ~n11634;
  assign n11637 = ~n11635 & ~n11636;
  assign n11638 = ~n11251 & ~n11637;
  assign n11639 = n11251 & n11637;
  assign n11640 = ~n11638 & ~n11639;
  assign n11641 = ~n11550 & n11640;
  assign n11642 = n11550 & ~n11640;
  assign n11643 = ~n11641 & ~n11642;
  assign n11644 = ~n11539 & n11643;
  assign n11645 = n11539 & ~n11643;
  assign n11646 = ~n11644 & ~n11645;
  assign n11647 = ~n11538 & n11646;
  assign n11648 = n11538 & ~n11646;
  assign n11649 = ~n11647 & ~n11648;
  assign n11650 = ~n11287 & ~n11649;
  assign n11651 = n11287 & n11649;
  assign n11652 = ~n11650 & ~n11651;
  assign n11653 = pi87  & n4896;
  assign n11654 = pi85  & n5148;
  assign n11655 = pi86  & n4891;
  assign n11656 = ~n11654 & ~n11655;
  assign n11657 = ~n11653 & n11656;
  assign n11658 = n2252 & n4899;
  assign n11659 = n11657 & ~n11658;
  assign n11660 = pi38  & ~n11659;
  assign n11661 = pi38  & ~n11660;
  assign n11662 = ~n11659 & ~n11660;
  assign n11663 = ~n11661 & ~n11662;
  assign n11664 = ~n11652 & ~n11663;
  assign n11665 = n11652 & n11663;
  assign n11666 = ~n11664 & ~n11665;
  assign n11667 = n11527 & ~n11666;
  assign n11668 = ~n11527 & n11666;
  assign n11669 = ~n11667 & ~n11668;
  assign n11670 = pi90  & n4182;
  assign n11671 = pi88  & n4416;
  assign n11672 = pi89  & n4177;
  assign n11673 = ~n11671 & ~n11672;
  assign n11674 = ~n11670 & n11673;
  assign n11675 = n2606 & n4185;
  assign n11676 = n11674 & ~n11675;
  assign n11677 = pi35  & ~n11676;
  assign n11678 = pi35  & ~n11677;
  assign n11679 = ~n11676 & ~n11677;
  assign n11680 = ~n11678 & ~n11679;
  assign n11681 = n11669 & ~n11680;
  assign n11682 = ~n11669 & n11680;
  assign n11683 = ~n11681 & ~n11682;
  assign n11684 = n11526 & ~n11683;
  assign n11685 = ~n11526 & n11683;
  assign n11686 = ~n11684 & ~n11685;
  assign n11687 = pi93  & n3550;
  assign n11688 = pi91  & n3735;
  assign n11689 = pi92  & n3545;
  assign n11690 = ~n11688 & ~n11689;
  assign n11691 = ~n11687 & n11690;
  assign n11692 = n3144 & n3553;
  assign n11693 = n11691 & ~n11692;
  assign n11694 = pi32  & ~n11693;
  assign n11695 = pi32  & ~n11694;
  assign n11696 = ~n11693 & ~n11694;
  assign n11697 = ~n11695 & ~n11696;
  assign n11698 = n11686 & ~n11697;
  assign n11699 = ~n11686 & n11697;
  assign n11700 = ~n11525 & ~n11699;
  assign n11701 = ~n11698 & n11700;
  assign n11702 = ~n11525 & ~n11701;
  assign n11703 = ~n11698 & ~n11701;
  assign n11704 = ~n11699 & n11703;
  assign n11705 = ~n11702 & ~n11704;
  assign n11706 = pi96  & n2976;
  assign n11707 = pi94  & n3182;
  assign n11708 = pi95  & n2971;
  assign n11709 = ~n11707 & ~n11708;
  assign n11710 = ~n11706 & n11709;
  assign n11711 = n2979 & n3921;
  assign n11712 = n11710 & ~n11711;
  assign n11713 = pi29  & ~n11712;
  assign n11714 = pi29  & ~n11713;
  assign n11715 = ~n11712 & ~n11713;
  assign n11716 = ~n11714 & ~n11715;
  assign n11717 = n11705 & n11716;
  assign n11718 = ~n11705 & ~n11716;
  assign n11719 = ~n11717 & ~n11718;
  assign n11720 = ~n11524 & n11719;
  assign n11721 = n11524 & ~n11719;
  assign n11722 = ~n11720 & ~n11721;
  assign n11723 = pi99  & n2486;
  assign n11724 = pi97  & n2644;
  assign n11725 = pi98  & n2481;
  assign n11726 = ~n11724 & ~n11725;
  assign n11727 = ~n11723 & n11726;
  assign n11728 = n2489 & n4584;
  assign n11729 = n11727 & ~n11728;
  assign n11730 = pi26  & ~n11729;
  assign n11731 = pi26  & ~n11730;
  assign n11732 = ~n11729 & ~n11730;
  assign n11733 = ~n11731 & ~n11732;
  assign n11734 = n11722 & ~n11733;
  assign n11735 = ~n11722 & n11733;
  assign n11736 = ~n11734 & ~n11735;
  assign n11737 = n11523 & ~n11736;
  assign n11738 = ~n11523 & n11736;
  assign n11739 = ~n11737 & ~n11738;
  assign n11740 = pi102  & n2004;
  assign n11741 = pi100  & n2141;
  assign n11742 = pi101  & n1999;
  assign n11743 = ~n11741 & ~n11742;
  assign n11744 = ~n11740 & n11743;
  assign n11745 = n2007 & n5296;
  assign n11746 = n11744 & ~n11745;
  assign n11747 = pi23  & ~n11746;
  assign n11748 = pi23  & ~n11747;
  assign n11749 = ~n11746 & ~n11747;
  assign n11750 = ~n11748 & ~n11749;
  assign n11751 = n11739 & ~n11750;
  assign n11752 = ~n11739 & n11750;
  assign n11753 = ~n11751 & ~n11752;
  assign n11754 = n11522 & ~n11753;
  assign n11755 = ~n11522 & n11753;
  assign n11756 = ~n11754 & ~n11755;
  assign n11757 = pi105  & n1582;
  assign n11758 = pi103  & n1713;
  assign n11759 = pi104  & n1577;
  assign n11760 = ~n11758 & ~n11759;
  assign n11761 = ~n11757 & n11760;
  assign n11762 = n1585 & n6065;
  assign n11763 = n11761 & ~n11762;
  assign n11764 = pi20  & ~n11763;
  assign n11765 = pi20  & ~n11764;
  assign n11766 = ~n11763 & ~n11764;
  assign n11767 = ~n11765 & ~n11766;
  assign n11768 = n11756 & ~n11767;
  assign n11769 = ~n11756 & n11767;
  assign n11770 = ~n11521 & ~n11769;
  assign n11771 = ~n11768 & n11770;
  assign n11772 = ~n11521 & ~n11771;
  assign n11773 = ~n11768 & ~n11771;
  assign n11774 = ~n11769 & n11773;
  assign n11775 = ~n11772 & ~n11774;
  assign n11776 = pi108  & n1269;
  assign n11777 = pi106  & n1340;
  assign n11778 = pi107  & n1264;
  assign n11779 = ~n11777 & ~n11778;
  assign n11780 = ~n11776 & n11779;
  assign n11781 = n1272 & n6639;
  assign n11782 = n11780 & ~n11781;
  assign n11783 = pi17  & ~n11782;
  assign n11784 = pi17  & ~n11783;
  assign n11785 = ~n11782 & ~n11783;
  assign n11786 = ~n11784 & ~n11785;
  assign n11787 = ~n11775 & ~n11786;
  assign n11788 = n11775 & n11786;
  assign n11789 = ~n11787 & ~n11788;
  assign n11790 = ~n11414 & ~n11789;
  assign n11791 = n11414 & n11789;
  assign n11792 = ~n11790 & ~n11791;
  assign n11793 = pi111  & n918;
  assign n11794 = pi109  & n1031;
  assign n11795 = pi110  & n913;
  assign n11796 = ~n11794 & ~n11795;
  assign n11797 = ~n11793 & n11796;
  assign n11798 = n921 & n7770;
  assign n11799 = n11797 & ~n11798;
  assign n11800 = pi14  & ~n11799;
  assign n11801 = pi14  & ~n11800;
  assign n11802 = ~n11799 & ~n11800;
  assign n11803 = ~n11801 & ~n11802;
  assign n11804 = ~n11792 & ~n11803;
  assign n11805 = n11792 & n11803;
  assign n11806 = ~n11804 & ~n11805;
  assign n11807 = ~n11520 & n11806;
  assign n11808 = n11520 & ~n11806;
  assign n11809 = ~n11807 & ~n11808;
  assign n11810 = pi114  & n675;
  assign n11811 = pi112  & n769;
  assign n11812 = pi113  & n670;
  assign n11813 = ~n11811 & ~n11812;
  assign n11814 = ~n11810 & n11813;
  assign n11815 = n678 & n8702;
  assign n11816 = n11814 & ~n11815;
  assign n11817 = pi11  & ~n11816;
  assign n11818 = pi11  & ~n11817;
  assign n11819 = ~n11816 & ~n11817;
  assign n11820 = ~n11818 & ~n11819;
  assign n11821 = n11809 & ~n11820;
  assign n11822 = ~n11809 & n11820;
  assign n11823 = ~n11821 & ~n11822;
  assign n11824 = ~n11519 & n11823;
  assign n11825 = n11519 & ~n11823;
  assign n11826 = ~n11824 & ~n11825;
  assign n11827 = ~n11518 & n11826;
  assign n11828 = n11518 & ~n11826;
  assign n11829 = ~n11827 & ~n11828;
  assign n11830 = ~n11507 & n11829;
  assign n11831 = n11507 & ~n11829;
  assign n11832 = ~n11830 & ~n11831;
  assign n11833 = ~n11506 & n11832;
  assign n11834 = n11506 & ~n11832;
  assign n11835 = ~n11833 & ~n11834;
  assign n11836 = ~n11495 & n11835;
  assign n11837 = n11495 & ~n11835;
  assign n11838 = ~n11836 & ~n11837;
  assign n11839 = ~n11477 & n11838;
  assign n11840 = n11477 & ~n11838;
  assign n11841 = ~n11839 & ~n11840;
  assign n11842 = ~n11476 & n11841;
  assign n11843 = n11476 & ~n11841;
  assign po59  = ~n11842 & ~n11843;
  assign n11845 = ~n11839 & ~n11842;
  assign n11846 = ~n11833 & ~n11836;
  assign n11847 = pi124  & n264;
  assign n11848 = pi122  & n281;
  assign n11849 = pi123  & n259;
  assign n11850 = ~n11848 & ~n11849;
  assign n11851 = ~n11847 & n11850;
  assign n11852 = ~n11485 & ~n11487;
  assign n11853 = ~pi123  & ~pi124 ;
  assign n11854 = pi123  & pi124 ;
  assign n11855 = ~n11853 & ~n11854;
  assign n11856 = ~n11852 & n11855;
  assign n11857 = n11852 & ~n11855;
  assign n11858 = ~n11856 & ~n11857;
  assign n11859 = n267 & n11858;
  assign n11860 = n11851 & ~n11859;
  assign n11861 = pi2  & ~n11860;
  assign n11862 = pi2  & ~n11861;
  assign n11863 = ~n11860 & ~n11861;
  assign n11864 = ~n11862 & ~n11863;
  assign n11865 = pi121  & n340;
  assign n11866 = pi119  & n380;
  assign n11867 = pi120  & n335;
  assign n11868 = ~n11866 & ~n11867;
  assign n11869 = ~n11865 & n11868;
  assign n11870 = n343 & n11086;
  assign n11871 = n11869 & ~n11870;
  assign n11872 = pi5  & ~n11871;
  assign n11873 = pi5  & ~n11872;
  assign n11874 = ~n11871 & ~n11872;
  assign n11875 = ~n11873 & ~n11874;
  assign n11876 = ~n11827 & ~n11830;
  assign n11877 = pi118  & n493;
  assign n11878 = pi116  & n533;
  assign n11879 = pi117  & n488;
  assign n11880 = ~n11878 & ~n11879;
  assign n11881 = ~n11877 & n11880;
  assign n11882 = n496 & n9716;
  assign n11883 = n11881 & ~n11882;
  assign n11884 = pi8  & ~n11883;
  assign n11885 = pi8  & ~n11884;
  assign n11886 = ~n11883 & ~n11884;
  assign n11887 = ~n11885 & ~n11886;
  assign n11888 = ~n11821 & ~n11824;
  assign n11889 = pi115  & n675;
  assign n11890 = pi113  & n769;
  assign n11891 = pi114  & n670;
  assign n11892 = ~n11890 & ~n11891;
  assign n11893 = ~n11889 & n11892;
  assign n11894 = n678 & n8727;
  assign n11895 = n11893 & ~n11894;
  assign n11896 = pi11  & ~n11895;
  assign n11897 = pi11  & ~n11896;
  assign n11898 = ~n11895 & ~n11896;
  assign n11899 = ~n11897 & ~n11898;
  assign n11900 = ~n11804 & ~n11807;
  assign n11901 = pi112  & n918;
  assign n11902 = pi110  & n1031;
  assign n11903 = pi111  & n913;
  assign n11904 = ~n11902 & ~n11903;
  assign n11905 = ~n11901 & n11904;
  assign n11906 = n921 & n7795;
  assign n11907 = n11905 & ~n11906;
  assign n11908 = pi14  & ~n11907;
  assign n11909 = pi14  & ~n11908;
  assign n11910 = ~n11907 & ~n11908;
  assign n11911 = ~n11909 & ~n11910;
  assign n11912 = ~n11788 & ~n11791;
  assign n11913 = pi109  & n1269;
  assign n11914 = pi107  & n1340;
  assign n11915 = pi108  & n1264;
  assign n11916 = ~n11914 & ~n11915;
  assign n11917 = ~n11913 & n11916;
  assign n11918 = n1272 & n7170;
  assign n11919 = n11917 & ~n11918;
  assign n11920 = pi17  & ~n11919;
  assign n11921 = pi17  & ~n11920;
  assign n11922 = ~n11919 & ~n11920;
  assign n11923 = ~n11921 & ~n11922;
  assign n11924 = ~n11751 & ~n11755;
  assign n11925 = ~n11734 & ~n11738;
  assign n11926 = ~n11718 & ~n11720;
  assign n11927 = ~n11681 & ~n11685;
  assign n11928 = ~n11664 & ~n11668;
  assign n11929 = pi85  & n5636;
  assign n11930 = pi83  & n5909;
  assign n11931 = pi84  & n5631;
  assign n11932 = ~n11930 & ~n11931;
  assign n11933 = ~n11929 & n11932;
  assign n11934 = n1943 & n5639;
  assign n11935 = n11933 & ~n11934;
  assign n11936 = pi41  & ~n11935;
  assign n11937 = pi41  & ~n11936;
  assign n11938 = ~n11935 & ~n11936;
  assign n11939 = ~n11937 & ~n11938;
  assign n11940 = ~n11641 & ~n11644;
  assign n11941 = pi82  & n6396;
  assign n11942 = pi80  & n6735;
  assign n11943 = pi81  & n6391;
  assign n11944 = ~n11942 & ~n11943;
  assign n11945 = ~n11941 & n11944;
  assign n11946 = n1532 & n6399;
  assign n11947 = n11945 & ~n11946;
  assign n11948 = pi44  & ~n11947;
  assign n11949 = pi44  & ~n11948;
  assign n11950 = ~n11947 & ~n11948;
  assign n11951 = ~n11949 & ~n11950;
  assign n11952 = ~n11634 & ~n11638;
  assign n11953 = pi79  & n7239;
  assign n11954 = pi77  & n7556;
  assign n11955 = pi78  & n7234;
  assign n11956 = ~n11954 & ~n11955;
  assign n11957 = ~n11953 & n11956;
  assign n11958 = n1105 & n7242;
  assign n11959 = n11957 & ~n11958;
  assign n11960 = pi47  & ~n11959;
  assign n11961 = pi47  & ~n11960;
  assign n11962 = ~n11959 & ~n11960;
  assign n11963 = ~n11961 & ~n11962;
  assign n11964 = ~n11618 & ~n11620;
  assign n11965 = pi76  & n8137;
  assign n11966 = pi74  & n8471;
  assign n11967 = pi75  & n8132;
  assign n11968 = ~n11966 & ~n11967;
  assign n11969 = ~n11965 & n11968;
  assign n11970 = n881 & n8140;
  assign n11971 = n11969 & ~n11970;
  assign n11972 = pi50  & ~n11971;
  assign n11973 = pi50  & ~n11972;
  assign n11974 = ~n11971 & ~n11972;
  assign n11975 = ~n11973 & ~n11974;
  assign n11976 = ~n11612 & ~n11614;
  assign n11977 = pi73  & n9096;
  assign n11978 = pi71  & n9453;
  assign n11979 = pi72  & n9091;
  assign n11980 = ~n11978 & ~n11979;
  assign n11981 = ~n11977 & n11980;
  assign n11982 = n639 & n9099;
  assign n11983 = n11981 & ~n11982;
  assign n11984 = pi53  & ~n11983;
  assign n11985 = pi53  & ~n11984;
  assign n11986 = ~n11983 & ~n11984;
  assign n11987 = ~n11985 & ~n11986;
  assign n11988 = pi67  & n11193;
  assign n11989 = pi65  & n11567;
  assign n11990 = pi66  & n11188;
  assign n11991 = ~n11989 & ~n11990;
  assign n11992 = ~n11988 & n11991;
  assign n11993 = n313 & n11196;
  assign n11994 = n11992 & ~n11993;
  assign n11995 = pi59  & ~n11994;
  assign n11996 = pi59  & ~n11995;
  assign n11997 = ~n11994 & ~n11995;
  assign n11998 = ~n11996 & ~n11997;
  assign n11999 = pi59  & ~pi60 ;
  assign n12000 = ~pi59  & pi60 ;
  assign n12001 = ~n11999 & ~n12000;
  assign n12002 = pi64  & ~n12001;
  assign n12003 = n11579 & n12002;
  assign n12004 = ~n11579 & ~n12002;
  assign n12005 = ~n12003 & ~n12004;
  assign n12006 = ~n11998 & n12005;
  assign n12007 = n11998 & ~n12005;
  assign n12008 = ~n12006 & ~n12007;
  assign n12009 = pi70  & n10135;
  assign n12010 = pi68  & n10478;
  assign n12011 = pi69  & n10130;
  assign n12012 = ~n12010 & ~n12011;
  assign n12013 = ~n12009 & n12012;
  assign n12014 = n430 & n10138;
  assign n12015 = n12013 & ~n12014;
  assign n12016 = pi56  & ~n12015;
  assign n12017 = pi56  & ~n12016;
  assign n12018 = ~n12015 & ~n12016;
  assign n12019 = ~n12017 & ~n12018;
  assign n12020 = n12008 & ~n12019;
  assign n12021 = ~n12008 & n12019;
  assign n12022 = ~n12020 & ~n12021;
  assign n12023 = ~n11597 & n12022;
  assign n12024 = n11597 & ~n12022;
  assign n12025 = ~n12023 & ~n12024;
  assign n12026 = ~n11987 & n12025;
  assign n12027 = n11987 & ~n12025;
  assign n12028 = ~n12026 & ~n12027;
  assign n12029 = ~n11976 & n12028;
  assign n12030 = n11976 & ~n12028;
  assign n12031 = ~n12029 & ~n12030;
  assign n12032 = n11975 & ~n12031;
  assign n12033 = ~n11975 & n12031;
  assign n12034 = ~n12032 & ~n12033;
  assign n12035 = ~n11964 & n12034;
  assign n12036 = n11964 & ~n12034;
  assign n12037 = ~n12035 & ~n12036;
  assign n12038 = ~n11963 & n12037;
  assign n12039 = n11963 & ~n12037;
  assign n12040 = ~n12038 & ~n12039;
  assign n12041 = ~n11952 & n12040;
  assign n12042 = n11952 & ~n12040;
  assign n12043 = ~n12041 & ~n12042;
  assign n12044 = ~n11951 & n12043;
  assign n12045 = ~n11951 & ~n12044;
  assign n12046 = n12043 & ~n12044;
  assign n12047 = ~n12045 & ~n12046;
  assign n12048 = ~n11940 & ~n12047;
  assign n12049 = n11940 & n12047;
  assign n12050 = ~n12048 & ~n12049;
  assign n12051 = ~n11939 & n12050;
  assign n12052 = n11939 & ~n12050;
  assign n12053 = ~n12051 & ~n12052;
  assign n12054 = ~n11648 & ~n11651;
  assign n12055 = n12053 & n12054;
  assign n12056 = ~n12053 & ~n12054;
  assign n12057 = ~n12055 & ~n12056;
  assign n12058 = pi88  & n4896;
  assign n12059 = pi86  & n5148;
  assign n12060 = pi87  & n4891;
  assign n12061 = ~n12059 & ~n12060;
  assign n12062 = ~n12058 & n12061;
  assign n12063 = n2277 & n4899;
  assign n12064 = n12062 & ~n12063;
  assign n12065 = pi38  & ~n12064;
  assign n12066 = pi38  & ~n12065;
  assign n12067 = ~n12064 & ~n12065;
  assign n12068 = ~n12066 & ~n12067;
  assign n12069 = n12057 & ~n12068;
  assign n12070 = ~n12057 & n12068;
  assign n12071 = ~n12069 & ~n12070;
  assign n12072 = n11928 & ~n12071;
  assign n12073 = ~n11928 & n12071;
  assign n12074 = ~n12072 & ~n12073;
  assign n12075 = pi91  & n4182;
  assign n12076 = pi89  & n4416;
  assign n12077 = pi90  & n4177;
  assign n12078 = ~n12076 & ~n12077;
  assign n12079 = ~n12075 & n12078;
  assign n12080 = n2926 & n4185;
  assign n12081 = n12079 & ~n12080;
  assign n12082 = pi35  & ~n12081;
  assign n12083 = pi35  & ~n12082;
  assign n12084 = ~n12081 & ~n12082;
  assign n12085 = ~n12083 & ~n12084;
  assign n12086 = n12074 & ~n12085;
  assign n12087 = ~n12074 & n12085;
  assign n12088 = ~n12086 & ~n12087;
  assign n12089 = n11927 & ~n12088;
  assign n12090 = ~n11927 & n12088;
  assign n12091 = ~n12089 & ~n12090;
  assign n12092 = pi94  & n3550;
  assign n12093 = pi92  & n3735;
  assign n12094 = pi93  & n3545;
  assign n12095 = ~n12093 & ~n12094;
  assign n12096 = ~n12092 & n12095;
  assign n12097 = n3499 & n3553;
  assign n12098 = n12096 & ~n12097;
  assign n12099 = pi32  & ~n12098;
  assign n12100 = pi32  & ~n12099;
  assign n12101 = ~n12098 & ~n12099;
  assign n12102 = ~n12100 & ~n12101;
  assign n12103 = ~n12091 & n12102;
  assign n12104 = n12091 & ~n12102;
  assign n12105 = ~n12103 & ~n12104;
  assign n12106 = ~n11703 & n12105;
  assign n12107 = n11703 & ~n12105;
  assign n12108 = ~n12106 & ~n12107;
  assign n12109 = pi97  & n2976;
  assign n12110 = pi95  & n3182;
  assign n12111 = pi96  & n2971;
  assign n12112 = ~n12110 & ~n12111;
  assign n12113 = ~n12109 & n12112;
  assign n12114 = n2979 & n3946;
  assign n12115 = n12113 & ~n12114;
  assign n12116 = pi29  & ~n12115;
  assign n12117 = pi29  & ~n12116;
  assign n12118 = ~n12115 & ~n12116;
  assign n12119 = ~n12117 & ~n12118;
  assign n12120 = n12108 & ~n12119;
  assign n12121 = ~n12108 & n12119;
  assign n12122 = ~n12120 & ~n12121;
  assign n12123 = ~n11926 & ~n12122;
  assign n12124 = n11926 & n12122;
  assign n12125 = ~n12123 & ~n12124;
  assign n12126 = pi100  & n2486;
  assign n12127 = pi98  & n2644;
  assign n12128 = pi99  & n2481;
  assign n12129 = ~n12127 & ~n12128;
  assign n12130 = ~n12126 & n12129;
  assign n12131 = n2489 & n4808;
  assign n12132 = n12130 & ~n12131;
  assign n12133 = pi26  & ~n12132;
  assign n12134 = pi26  & ~n12133;
  assign n12135 = ~n12132 & ~n12133;
  assign n12136 = ~n12134 & ~n12135;
  assign n12137 = ~n12125 & ~n12136;
  assign n12138 = n12125 & n12136;
  assign n12139 = ~n12137 & ~n12138;
  assign n12140 = n11925 & ~n12139;
  assign n12141 = ~n11925 & n12139;
  assign n12142 = ~n12140 & ~n12141;
  assign n12143 = pi103  & n2004;
  assign n12144 = pi101  & n2141;
  assign n12145 = pi102  & n1999;
  assign n12146 = ~n12144 & ~n12145;
  assign n12147 = ~n12143 & n12146;
  assign n12148 = n2007 & n5540;
  assign n12149 = n12147 & ~n12148;
  assign n12150 = pi23  & ~n12149;
  assign n12151 = pi23  & ~n12150;
  assign n12152 = ~n12149 & ~n12150;
  assign n12153 = ~n12151 & ~n12152;
  assign n12154 = n12142 & ~n12153;
  assign n12155 = ~n12142 & n12153;
  assign n12156 = ~n12154 & ~n12155;
  assign n12157 = n11924 & ~n12156;
  assign n12158 = ~n11924 & n12156;
  assign n12159 = ~n12157 & ~n12158;
  assign n12160 = pi106  & n1582;
  assign n12161 = pi104  & n1713;
  assign n12162 = pi105  & n1577;
  assign n12163 = ~n12161 & ~n12162;
  assign n12164 = ~n12160 & n12163;
  assign n12165 = n1585 & n6090;
  assign n12166 = n12164 & ~n12165;
  assign n12167 = pi20  & ~n12166;
  assign n12168 = pi20  & ~n12167;
  assign n12169 = ~n12166 & ~n12167;
  assign n12170 = ~n12168 & ~n12169;
  assign n12171 = ~n12159 & n12170;
  assign n12172 = n12159 & ~n12170;
  assign n12173 = ~n12171 & ~n12172;
  assign n12174 = ~n11773 & n12173;
  assign n12175 = n11773 & ~n12173;
  assign n12176 = ~n12174 & ~n12175;
  assign n12177 = ~n11923 & n12176;
  assign n12178 = n11923 & ~n12176;
  assign n12179 = ~n12177 & ~n12178;
  assign n12180 = n11912 & n12179;
  assign n12181 = ~n11912 & ~n12179;
  assign n12182 = ~n12180 & ~n12181;
  assign n12183 = ~n11911 & n12182;
  assign n12184 = n11911 & ~n12182;
  assign n12185 = ~n12183 & ~n12184;
  assign n12186 = ~n11900 & n12185;
  assign n12187 = n11900 & ~n12185;
  assign n12188 = ~n12186 & ~n12187;
  assign n12189 = ~n11899 & n12188;
  assign n12190 = n11899 & ~n12188;
  assign n12191 = ~n12189 & ~n12190;
  assign n12192 = ~n11888 & n12191;
  assign n12193 = n11888 & ~n12191;
  assign n12194 = ~n12192 & ~n12193;
  assign n12195 = ~n11887 & n12194;
  assign n12196 = n11887 & ~n12194;
  assign n12197 = ~n12195 & ~n12196;
  assign n12198 = ~n11876 & n12197;
  assign n12199 = n11876 & ~n12197;
  assign n12200 = ~n12198 & ~n12199;
  assign n12201 = ~n11875 & n12200;
  assign n12202 = n11875 & ~n12200;
  assign n12203 = ~n12201 & ~n12202;
  assign n12204 = ~n11864 & n12203;
  assign n12205 = n11864 & ~n12203;
  assign n12206 = ~n12204 & ~n12205;
  assign n12207 = ~n11846 & n12206;
  assign n12208 = n11846 & ~n12206;
  assign n12209 = ~n12207 & ~n12208;
  assign n12210 = ~n11845 & n12209;
  assign n12211 = n11845 & ~n12209;
  assign po60  = ~n12210 & ~n12211;
  assign n12213 = ~n12201 & ~n12204;
  assign n12214 = ~n12195 & ~n12198;
  assign n12215 = ~n12189 & ~n12192;
  assign n12216 = pi116  & n675;
  assign n12217 = pi114  & n769;
  assign n12218 = pi115  & n670;
  assign n12219 = ~n12217 & ~n12218;
  assign n12220 = ~n12216 & n12219;
  assign n12221 = n678 & n9042;
  assign n12222 = n12220 & ~n12221;
  assign n12223 = pi11  & ~n12222;
  assign n12224 = pi11  & ~n12223;
  assign n12225 = ~n12222 & ~n12223;
  assign n12226 = ~n12224 & ~n12225;
  assign n12227 = ~n12183 & ~n12186;
  assign n12228 = pi113  & n918;
  assign n12229 = pi111  & n1031;
  assign n12230 = pi112  & n913;
  assign n12231 = ~n12229 & ~n12230;
  assign n12232 = ~n12228 & n12231;
  assign n12233 = n921 & n8387;
  assign n12234 = n12232 & ~n12233;
  assign n12235 = pi14  & ~n12234;
  assign n12236 = pi14  & ~n12235;
  assign n12237 = ~n12234 & ~n12235;
  assign n12238 = ~n12236 & ~n12237;
  assign n12239 = ~n12177 & ~n12180;
  assign n12240 = ~n12172 & ~n12174;
  assign n12241 = ~n12154 & ~n12158;
  assign n12242 = ~n12137 & ~n12141;
  assign n12243 = pi98  & n2976;
  assign n12244 = pi96  & n3182;
  assign n12245 = pi97  & n2971;
  assign n12246 = ~n12244 & ~n12245;
  assign n12247 = ~n12243 & n12246;
  assign n12248 = n2979 & n4360;
  assign n12249 = n12247 & ~n12248;
  assign n12250 = pi29  & ~n12249;
  assign n12251 = pi29  & ~n12250;
  assign n12252 = ~n12249 & ~n12250;
  assign n12253 = ~n12251 & ~n12252;
  assign n12254 = ~n12104 & ~n12106;
  assign n12255 = ~n12086 & ~n12090;
  assign n12256 = ~n12069 & ~n12073;
  assign n12257 = ~n12051 & ~n12055;
  assign n12258 = ~n12044 & ~n12048;
  assign n12259 = ~n12038 & ~n12041;
  assign n12260 = ~n12033 & ~n12035;
  assign n12261 = ~n12026 & ~n12029;
  assign n12262 = ~n12020 & ~n12023;
  assign n12263 = pi71  & n10135;
  assign n12264 = pi69  & n10478;
  assign n12265 = pi70  & n10130;
  assign n12266 = ~n12264 & ~n12265;
  assign n12267 = ~n12263 & n12266;
  assign n12268 = n476 & n10138;
  assign n12269 = n12267 & ~n12268;
  assign n12270 = pi56  & ~n12269;
  assign n12271 = pi56  & ~n12270;
  assign n12272 = ~n12269 & ~n12270;
  assign n12273 = ~n12271 & ~n12272;
  assign n12274 = ~n12003 & ~n12006;
  assign n12275 = pi68  & n11193;
  assign n12276 = pi66  & n11567;
  assign n12277 = pi67  & n11188;
  assign n12278 = ~n12276 & ~n12277;
  assign n12279 = ~n12275 & n12278;
  assign n12280 = n364 & n11196;
  assign n12281 = n12279 & ~n12280;
  assign n12282 = pi59  & ~n12281;
  assign n12283 = pi59  & ~n12282;
  assign n12284 = ~n12281 & ~n12282;
  assign n12285 = ~n12283 & ~n12284;
  assign n12286 = pi62  & ~n12002;
  assign n12287 = ~pi60  & pi61 ;
  assign n12288 = pi60  & ~pi61 ;
  assign n12289 = ~n12287 & ~n12288;
  assign n12290 = n12001 & ~n12289;
  assign n12291 = pi64  & n12290;
  assign n12292 = ~pi61  & pi62 ;
  assign n12293 = pi61  & ~pi62 ;
  assign n12294 = ~n12292 & ~n12293;
  assign n12295 = ~n12001 & n12294;
  assign n12296 = pi65  & n12295;
  assign n12297 = ~n12291 & ~n12296;
  assign n12298 = ~n12001 & ~n12294;
  assign n12299 = n270 & n12298;
  assign n12300 = n12297 & ~n12299;
  assign n12301 = pi62  & ~n12300;
  assign n12302 = pi62  & ~n12301;
  assign n12303 = ~n12300 & ~n12301;
  assign n12304 = ~n12302 & ~n12303;
  assign n12305 = n12286 & ~n12304;
  assign n12306 = ~n12286 & n12304;
  assign n12307 = ~n12305 & ~n12306;
  assign n12308 = n12285 & ~n12307;
  assign n12309 = ~n12285 & n12307;
  assign n12310 = ~n12308 & ~n12309;
  assign n12311 = ~n12274 & n12310;
  assign n12312 = n12274 & ~n12310;
  assign n12313 = ~n12311 & ~n12312;
  assign n12314 = n12273 & ~n12313;
  assign n12315 = ~n12273 & n12313;
  assign n12316 = ~n12314 & ~n12315;
  assign n12317 = ~n12262 & n12316;
  assign n12318 = n12262 & ~n12316;
  assign n12319 = ~n12317 & ~n12318;
  assign n12320 = pi74  & n9096;
  assign n12321 = pi72  & n9453;
  assign n12322 = pi73  & n9091;
  assign n12323 = ~n12321 & ~n12322;
  assign n12324 = ~n12320 & n12323;
  assign n12325 = n722 & n9099;
  assign n12326 = n12324 & ~n12325;
  assign n12327 = pi53  & ~n12326;
  assign n12328 = pi53  & ~n12327;
  assign n12329 = ~n12326 & ~n12327;
  assign n12330 = ~n12328 & ~n12329;
  assign n12331 = n12319 & ~n12330;
  assign n12332 = ~n12319 & n12330;
  assign n12333 = ~n12331 & ~n12332;
  assign n12334 = n12261 & ~n12333;
  assign n12335 = ~n12261 & n12333;
  assign n12336 = ~n12334 & ~n12335;
  assign n12337 = pi77  & n8137;
  assign n12338 = pi75  & n8471;
  assign n12339 = pi76  & n8132;
  assign n12340 = ~n12338 & ~n12339;
  assign n12341 = ~n12337 & n12340;
  assign n12342 = n984 & n8140;
  assign n12343 = n12341 & ~n12342;
  assign n12344 = pi50  & ~n12343;
  assign n12345 = pi50  & ~n12344;
  assign n12346 = ~n12343 & ~n12344;
  assign n12347 = ~n12345 & ~n12346;
  assign n12348 = n12336 & ~n12347;
  assign n12349 = ~n12336 & n12347;
  assign n12350 = ~n12260 & ~n12349;
  assign n12351 = ~n12348 & n12350;
  assign n12352 = ~n12260 & ~n12351;
  assign n12353 = ~n12348 & ~n12351;
  assign n12354 = ~n12349 & n12353;
  assign n12355 = ~n12352 & ~n12354;
  assign n12356 = pi80  & n7239;
  assign n12357 = pi78  & n7556;
  assign n12358 = pi79  & n7234;
  assign n12359 = ~n12357 & ~n12358;
  assign n12360 = ~n12356 & n12359;
  assign n12361 = n1205 & n7242;
  assign n12362 = n12360 & ~n12361;
  assign n12363 = pi47  & ~n12362;
  assign n12364 = pi47  & ~n12363;
  assign n12365 = ~n12362 & ~n12363;
  assign n12366 = ~n12364 & ~n12365;
  assign n12367 = ~n12355 & ~n12366;
  assign n12368 = n12355 & n12366;
  assign n12369 = ~n12367 & ~n12368;
  assign n12370 = n12259 & ~n12369;
  assign n12371 = ~n12259 & n12369;
  assign n12372 = ~n12370 & ~n12371;
  assign n12373 = pi83  & n6396;
  assign n12374 = pi81  & n6735;
  assign n12375 = pi82  & n6391;
  assign n12376 = ~n12374 & ~n12375;
  assign n12377 = ~n12373 & n12376;
  assign n12378 = n1672 & n6399;
  assign n12379 = n12377 & ~n12378;
  assign n12380 = pi44  & ~n12379;
  assign n12381 = pi44  & ~n12380;
  assign n12382 = ~n12379 & ~n12380;
  assign n12383 = ~n12381 & ~n12382;
  assign n12384 = n12372 & ~n12383;
  assign n12385 = ~n12372 & n12383;
  assign n12386 = ~n12258 & ~n12385;
  assign n12387 = ~n12384 & n12386;
  assign n12388 = ~n12258 & ~n12387;
  assign n12389 = ~n12384 & ~n12387;
  assign n12390 = ~n12385 & n12389;
  assign n12391 = ~n12388 & ~n12390;
  assign n12392 = pi86  & n5636;
  assign n12393 = pi84  & n5909;
  assign n12394 = pi85  & n5631;
  assign n12395 = ~n12393 & ~n12394;
  assign n12396 = ~n12392 & n12395;
  assign n12397 = n2099 & n5639;
  assign n12398 = n12396 & ~n12397;
  assign n12399 = pi41  & ~n12398;
  assign n12400 = pi41  & ~n12399;
  assign n12401 = ~n12398 & ~n12399;
  assign n12402 = ~n12400 & ~n12401;
  assign n12403 = ~n12391 & ~n12402;
  assign n12404 = n12391 & n12402;
  assign n12405 = ~n12403 & ~n12404;
  assign n12406 = n12257 & ~n12405;
  assign n12407 = ~n12257 & n12405;
  assign n12408 = ~n12406 & ~n12407;
  assign n12409 = pi89  & n4896;
  assign n12410 = pi87  & n5148;
  assign n12411 = pi88  & n4891;
  assign n12412 = ~n12410 & ~n12411;
  assign n12413 = ~n12409 & n12412;
  assign n12414 = n2432 & n4899;
  assign n12415 = n12413 & ~n12414;
  assign n12416 = pi38  & ~n12415;
  assign n12417 = pi38  & ~n12416;
  assign n12418 = ~n12415 & ~n12416;
  assign n12419 = ~n12417 & ~n12418;
  assign n12420 = n12408 & ~n12419;
  assign n12421 = ~n12408 & n12419;
  assign n12422 = ~n12420 & ~n12421;
  assign n12423 = n12256 & ~n12422;
  assign n12424 = ~n12256 & n12422;
  assign n12425 = ~n12423 & ~n12424;
  assign n12426 = pi92  & n4182;
  assign n12427 = pi90  & n4416;
  assign n12428 = pi91  & n4177;
  assign n12429 = ~n12427 & ~n12428;
  assign n12430 = ~n12426 & n12429;
  assign n12431 = n3119 & n4185;
  assign n12432 = n12430 & ~n12431;
  assign n12433 = pi35  & ~n12432;
  assign n12434 = pi35  & ~n12433;
  assign n12435 = ~n12432 & ~n12433;
  assign n12436 = ~n12434 & ~n12435;
  assign n12437 = n12425 & ~n12436;
  assign n12438 = ~n12425 & n12436;
  assign n12439 = ~n12437 & ~n12438;
  assign n12440 = n12255 & ~n12439;
  assign n12441 = ~n12255 & n12439;
  assign n12442 = ~n12440 & ~n12441;
  assign n12443 = pi95  & n3550;
  assign n12444 = pi93  & n3735;
  assign n12445 = pi94  & n3545;
  assign n12446 = ~n12444 & ~n12445;
  assign n12447 = ~n12443 & n12446;
  assign n12448 = n3553 & n3710;
  assign n12449 = n12447 & ~n12448;
  assign n12450 = pi32  & ~n12449;
  assign n12451 = pi32  & ~n12450;
  assign n12452 = ~n12449 & ~n12450;
  assign n12453 = ~n12451 & ~n12452;
  assign n12454 = n12442 & ~n12453;
  assign n12455 = ~n12442 & n12453;
  assign n12456 = ~n12454 & ~n12455;
  assign n12457 = ~n12254 & n12456;
  assign n12458 = n12254 & ~n12456;
  assign n12459 = ~n12457 & ~n12458;
  assign n12460 = ~n12253 & n12459;
  assign n12461 = n12253 & ~n12459;
  assign n12462 = ~n12460 & ~n12461;
  assign n12463 = ~n12121 & ~n12124;
  assign n12464 = ~n12462 & ~n12463;
  assign n12465 = n12462 & n12463;
  assign n12466 = ~n12464 & ~n12465;
  assign n12467 = pi101  & n2486;
  assign n12468 = pi99  & n2644;
  assign n12469 = pi100  & n2481;
  assign n12470 = ~n12468 & ~n12469;
  assign n12471 = ~n12467 & n12470;
  assign n12472 = n2489 & n5056;
  assign n12473 = n12471 & ~n12472;
  assign n12474 = pi26  & ~n12473;
  assign n12475 = pi26  & ~n12474;
  assign n12476 = ~n12473 & ~n12474;
  assign n12477 = ~n12475 & ~n12476;
  assign n12478 = n12466 & ~n12477;
  assign n12479 = ~n12466 & n12477;
  assign n12480 = ~n12478 & ~n12479;
  assign n12481 = n12242 & ~n12480;
  assign n12482 = ~n12242 & n12480;
  assign n12483 = ~n12481 & ~n12482;
  assign n12484 = pi104  & n2004;
  assign n12485 = pi102  & n2141;
  assign n12486 = pi103  & n1999;
  assign n12487 = ~n12485 & ~n12486;
  assign n12488 = ~n12484 & n12487;
  assign n12489 = n2007 & n5565;
  assign n12490 = n12488 & ~n12489;
  assign n12491 = pi23  & ~n12490;
  assign n12492 = pi23  & ~n12491;
  assign n12493 = ~n12490 & ~n12491;
  assign n12494 = ~n12492 & ~n12493;
  assign n12495 = n12483 & ~n12494;
  assign n12496 = ~n12483 & n12494;
  assign n12497 = ~n12495 & ~n12496;
  assign n12498 = n12241 & ~n12497;
  assign n12499 = ~n12241 & n12497;
  assign n12500 = ~n12498 & ~n12499;
  assign n12501 = pi107  & n1582;
  assign n12502 = pi105  & n1713;
  assign n12503 = pi106  & n1577;
  assign n12504 = ~n12502 & ~n12503;
  assign n12505 = ~n12501 & n12504;
  assign n12506 = n1585 & n6614;
  assign n12507 = n12505 & ~n12506;
  assign n12508 = pi20  & ~n12507;
  assign n12509 = pi20  & ~n12508;
  assign n12510 = ~n12507 & ~n12508;
  assign n12511 = ~n12509 & ~n12510;
  assign n12512 = n12500 & ~n12511;
  assign n12513 = ~n12500 & n12511;
  assign n12514 = ~n12240 & ~n12513;
  assign n12515 = ~n12512 & n12514;
  assign n12516 = ~n12240 & ~n12515;
  assign n12517 = ~n12512 & ~n12515;
  assign n12518 = ~n12513 & n12517;
  assign n12519 = ~n12516 & ~n12518;
  assign n12520 = pi110  & n1269;
  assign n12521 = pi108  & n1340;
  assign n12522 = pi109  & n1264;
  assign n12523 = ~n12521 & ~n12522;
  assign n12524 = ~n12520 & n12523;
  assign n12525 = n1272 & n7474;
  assign n12526 = n12524 & ~n12525;
  assign n12527 = pi17  & ~n12526;
  assign n12528 = pi17  & ~n12527;
  assign n12529 = ~n12526 & ~n12527;
  assign n12530 = ~n12528 & ~n12529;
  assign n12531 = n12519 & n12530;
  assign n12532 = ~n12519 & ~n12530;
  assign n12533 = ~n12531 & ~n12532;
  assign n12534 = ~n12239 & n12533;
  assign n12535 = n12239 & ~n12533;
  assign n12536 = ~n12534 & ~n12535;
  assign n12537 = n12238 & ~n12536;
  assign n12538 = ~n12238 & n12536;
  assign n12539 = ~n12537 & ~n12538;
  assign n12540 = ~n12227 & n12539;
  assign n12541 = n12227 & ~n12539;
  assign n12542 = ~n12540 & ~n12541;
  assign n12543 = n12226 & ~n12542;
  assign n12544 = ~n12226 & n12542;
  assign n12545 = ~n12543 & ~n12544;
  assign n12546 = ~n12215 & n12545;
  assign n12547 = n12215 & ~n12545;
  assign n12548 = ~n12546 & ~n12547;
  assign n12549 = pi119  & n493;
  assign n12550 = pi117  & n533;
  assign n12551 = pi118  & n488;
  assign n12552 = ~n12550 & ~n12551;
  assign n12553 = ~n12549 & n12552;
  assign n12554 = n496 & n10048;
  assign n12555 = n12553 & ~n12554;
  assign n12556 = pi8  & ~n12555;
  assign n12557 = pi8  & ~n12556;
  assign n12558 = ~n12555 & ~n12556;
  assign n12559 = ~n12557 & ~n12558;
  assign n12560 = n12548 & ~n12559;
  assign n12561 = ~n12548 & n12559;
  assign n12562 = ~n12560 & ~n12561;
  assign n12563 = n12214 & ~n12562;
  assign n12564 = ~n12214 & n12562;
  assign n12565 = ~n12563 & ~n12564;
  assign n12566 = pi122  & n340;
  assign n12567 = pi120  & n380;
  assign n12568 = pi121  & n335;
  assign n12569 = ~n12567 & ~n12568;
  assign n12570 = ~n12566 & n12569;
  assign n12571 = n343 & n11463;
  assign n12572 = n12570 & ~n12571;
  assign n12573 = pi5  & ~n12572;
  assign n12574 = pi5  & ~n12573;
  assign n12575 = ~n12572 & ~n12573;
  assign n12576 = ~n12574 & ~n12575;
  assign n12577 = ~n12565 & n12576;
  assign n12578 = n12565 & ~n12576;
  assign n12579 = ~n12577 & ~n12578;
  assign n12580 = pi125  & n264;
  assign n12581 = pi123  & n281;
  assign n12582 = pi124  & n259;
  assign n12583 = ~n12581 & ~n12582;
  assign n12584 = ~n12580 & n12583;
  assign n12585 = ~n11854 & ~n11856;
  assign n12586 = ~pi124  & ~pi125 ;
  assign n12587 = pi124  & pi125 ;
  assign n12588 = ~n12586 & ~n12587;
  assign n12589 = ~n12585 & n12588;
  assign n12590 = n12585 & ~n12588;
  assign n12591 = ~n12589 & ~n12590;
  assign n12592 = n267 & n12591;
  assign n12593 = n12584 & ~n12592;
  assign n12594 = pi2  & ~n12593;
  assign n12595 = pi2  & ~n12594;
  assign n12596 = ~n12593 & ~n12594;
  assign n12597 = ~n12595 & ~n12596;
  assign n12598 = n12579 & ~n12597;
  assign n12599 = ~n12579 & n12597;
  assign n12600 = ~n12598 & ~n12599;
  assign n12601 = n12213 & ~n12600;
  assign n12602 = ~n12213 & n12600;
  assign n12603 = ~n12601 & ~n12602;
  assign n12604 = ~n12207 & ~n12210;
  assign n12605 = n12603 & ~n12604;
  assign n12606 = ~n12603 & n12604;
  assign po61  = ~n12605 & ~n12606;
  assign n12608 = ~n12602 & ~n12605;
  assign n12609 = ~n12578 & ~n12598;
  assign n12610 = ~n12560 & ~n12564;
  assign n12611 = ~n12544 & ~n12546;
  assign n12612 = pi117  & n675;
  assign n12613 = pi115  & n769;
  assign n12614 = pi116  & n670;
  assign n12615 = ~n12613 & ~n12614;
  assign n12616 = ~n12612 & n12615;
  assign n12617 = n678 & n9691;
  assign n12618 = n12616 & ~n12617;
  assign n12619 = pi11  & ~n12618;
  assign n12620 = pi11  & ~n12619;
  assign n12621 = ~n12618 & ~n12619;
  assign n12622 = ~n12620 & ~n12621;
  assign n12623 = ~n12538 & ~n12540;
  assign n12624 = ~n12532 & ~n12534;
  assign n12625 = pi111  & n1269;
  assign n12626 = pi109  & n1340;
  assign n12627 = pi110  & n1264;
  assign n12628 = ~n12626 & ~n12627;
  assign n12629 = ~n12625 & n12628;
  assign n12630 = n1272 & n7770;
  assign n12631 = n12629 & ~n12630;
  assign n12632 = pi17  & ~n12631;
  assign n12633 = pi17  & ~n12632;
  assign n12634 = ~n12631 & ~n12632;
  assign n12635 = ~n12633 & ~n12634;
  assign n12636 = ~n12495 & ~n12499;
  assign n12637 = ~n12478 & ~n12482;
  assign n12638 = ~n12460 & ~n12465;
  assign n12639 = ~n12454 & ~n12457;
  assign n12640 = ~n12437 & ~n12441;
  assign n12641 = ~n12420 & ~n12424;
  assign n12642 = ~n12403 & ~n12407;
  assign n12643 = pi87  & n5636;
  assign n12644 = pi85  & n5909;
  assign n12645 = pi86  & n5631;
  assign n12646 = ~n12644 & ~n12645;
  assign n12647 = ~n12643 & n12646;
  assign n12648 = n2252 & n5639;
  assign n12649 = n12647 & ~n12648;
  assign n12650 = pi41  & ~n12649;
  assign n12651 = pi41  & ~n12650;
  assign n12652 = ~n12649 & ~n12650;
  assign n12653 = ~n12651 & ~n12652;
  assign n12654 = pi84  & n6396;
  assign n12655 = pi82  & n6735;
  assign n12656 = pi83  & n6391;
  assign n12657 = ~n12655 & ~n12656;
  assign n12658 = ~n12654 & n12657;
  assign n12659 = n1805 & n6399;
  assign n12660 = n12658 & ~n12659;
  assign n12661 = pi44  & ~n12660;
  assign n12662 = pi44  & ~n12661;
  assign n12663 = ~n12660 & ~n12661;
  assign n12664 = ~n12662 & ~n12663;
  assign n12665 = ~n12367 & ~n12371;
  assign n12666 = pi81  & n7239;
  assign n12667 = pi79  & n7556;
  assign n12668 = pi80  & n7234;
  assign n12669 = ~n12667 & ~n12668;
  assign n12670 = ~n12666 & n12669;
  assign n12671 = n1413 & n7242;
  assign n12672 = n12670 & ~n12671;
  assign n12673 = pi47  & ~n12672;
  assign n12674 = pi47  & ~n12673;
  assign n12675 = ~n12672 & ~n12673;
  assign n12676 = ~n12674 & ~n12675;
  assign n12677 = ~n12331 & ~n12335;
  assign n12678 = pi75  & n9096;
  assign n12679 = pi73  & n9453;
  assign n12680 = pi74  & n9091;
  assign n12681 = ~n12679 & ~n12680;
  assign n12682 = ~n12678 & n12681;
  assign n12683 = n747 & n9099;
  assign n12684 = n12682 & ~n12683;
  assign n12685 = pi53  & ~n12684;
  assign n12686 = pi53  & ~n12685;
  assign n12687 = ~n12684 & ~n12685;
  assign n12688 = ~n12686 & ~n12687;
  assign n12689 = ~n12315 & ~n12317;
  assign n12690 = ~n12309 & ~n12311;
  assign n12691 = pi66  & n12295;
  assign n12692 = n12001 & ~n12294;
  assign n12693 = n12289 & n12692;
  assign n12694 = pi64  & n12693;
  assign n12695 = pi65  & n12290;
  assign n12696 = ~n12694 & ~n12695;
  assign n12697 = ~n12691 & n12696;
  assign n12698 = n291 & n12298;
  assign n12699 = n12697 & ~n12698;
  assign n12700 = pi62  & ~n12699;
  assign n12701 = pi62  & ~n12700;
  assign n12702 = ~n12699 & ~n12700;
  assign n12703 = ~n12701 & ~n12702;
  assign n12704 = ~n12305 & n12703;
  assign n12705 = n12305 & ~n12703;
  assign n12706 = ~n12704 & ~n12705;
  assign n12707 = pi69  & n11193;
  assign n12708 = pi67  & n11567;
  assign n12709 = pi68  & n11188;
  assign n12710 = ~n12708 & ~n12709;
  assign n12711 = ~n12707 & n12710;
  assign n12712 = n405 & n11196;
  assign n12713 = n12711 & ~n12712;
  assign n12714 = pi59  & ~n12713;
  assign n12715 = pi59  & ~n12714;
  assign n12716 = ~n12713 & ~n12714;
  assign n12717 = ~n12715 & ~n12716;
  assign n12718 = n12706 & ~n12717;
  assign n12719 = ~n12706 & n12717;
  assign n12720 = ~n12690 & ~n12719;
  assign n12721 = ~n12718 & n12720;
  assign n12722 = ~n12690 & ~n12721;
  assign n12723 = ~n12718 & ~n12721;
  assign n12724 = ~n12719 & n12723;
  assign n12725 = ~n12722 & ~n12724;
  assign n12726 = pi72  & n10135;
  assign n12727 = pi70  & n10478;
  assign n12728 = pi71  & n10130;
  assign n12729 = ~n12727 & ~n12728;
  assign n12730 = ~n12726 & n12729;
  assign n12731 = n575 & n10138;
  assign n12732 = n12730 & ~n12731;
  assign n12733 = pi56  & ~n12732;
  assign n12734 = pi56  & ~n12733;
  assign n12735 = ~n12732 & ~n12733;
  assign n12736 = ~n12734 & ~n12735;
  assign n12737 = n12725 & n12736;
  assign n12738 = ~n12725 & ~n12736;
  assign n12739 = ~n12737 & ~n12738;
  assign n12740 = ~n12689 & n12739;
  assign n12741 = n12689 & ~n12739;
  assign n12742 = ~n12740 & ~n12741;
  assign n12743 = n12688 & ~n12742;
  assign n12744 = ~n12688 & n12742;
  assign n12745 = ~n12743 & ~n12744;
  assign n12746 = ~n12677 & n12745;
  assign n12747 = n12677 & ~n12745;
  assign n12748 = ~n12746 & ~n12747;
  assign n12749 = pi78  & n8137;
  assign n12750 = pi76  & n8471;
  assign n12751 = pi77  & n8132;
  assign n12752 = ~n12750 & ~n12751;
  assign n12753 = ~n12749 & n12752;
  assign n12754 = n1009 & n8140;
  assign n12755 = n12753 & ~n12754;
  assign n12756 = pi50  & ~n12755;
  assign n12757 = pi50  & ~n12756;
  assign n12758 = ~n12755 & ~n12756;
  assign n12759 = ~n12757 & ~n12758;
  assign n12760 = n12748 & ~n12759;
  assign n12761 = n12748 & ~n12760;
  assign n12762 = ~n12759 & ~n12760;
  assign n12763 = ~n12761 & ~n12762;
  assign n12764 = ~n12353 & ~n12763;
  assign n12765 = n12353 & n12763;
  assign n12766 = ~n12764 & ~n12765;
  assign n12767 = ~n12676 & n12766;
  assign n12768 = n12676 & ~n12766;
  assign n12769 = ~n12767 & ~n12768;
  assign n12770 = ~n12665 & n12769;
  assign n12771 = n12665 & ~n12769;
  assign n12772 = ~n12770 & ~n12771;
  assign n12773 = ~n12664 & n12772;
  assign n12774 = n12664 & ~n12772;
  assign n12775 = ~n12773 & ~n12774;
  assign n12776 = ~n12389 & n12775;
  assign n12777 = n12389 & ~n12775;
  assign n12778 = ~n12776 & ~n12777;
  assign n12779 = ~n12653 & n12778;
  assign n12780 = n12653 & ~n12778;
  assign n12781 = ~n12779 & ~n12780;
  assign n12782 = n12642 & ~n12781;
  assign n12783 = ~n12642 & n12781;
  assign n12784 = ~n12782 & ~n12783;
  assign n12785 = pi90  & n4896;
  assign n12786 = pi88  & n5148;
  assign n12787 = pi89  & n4891;
  assign n12788 = ~n12786 & ~n12787;
  assign n12789 = ~n12785 & n12788;
  assign n12790 = n2606 & n4899;
  assign n12791 = n12789 & ~n12790;
  assign n12792 = pi38  & ~n12791;
  assign n12793 = pi38  & ~n12792;
  assign n12794 = ~n12791 & ~n12792;
  assign n12795 = ~n12793 & ~n12794;
  assign n12796 = n12784 & ~n12795;
  assign n12797 = ~n12784 & n12795;
  assign n12798 = ~n12796 & ~n12797;
  assign n12799 = n12641 & ~n12798;
  assign n12800 = ~n12641 & n12798;
  assign n12801 = ~n12799 & ~n12800;
  assign n12802 = pi93  & n4182;
  assign n12803 = pi91  & n4416;
  assign n12804 = pi92  & n4177;
  assign n12805 = ~n12803 & ~n12804;
  assign n12806 = ~n12802 & n12805;
  assign n12807 = n3144 & n4185;
  assign n12808 = n12806 & ~n12807;
  assign n12809 = pi35  & ~n12808;
  assign n12810 = pi35  & ~n12809;
  assign n12811 = ~n12808 & ~n12809;
  assign n12812 = ~n12810 & ~n12811;
  assign n12813 = n12801 & ~n12812;
  assign n12814 = ~n12801 & n12812;
  assign n12815 = ~n12813 & ~n12814;
  assign n12816 = n12640 & ~n12815;
  assign n12817 = ~n12640 & n12815;
  assign n12818 = ~n12816 & ~n12817;
  assign n12819 = pi96  & n3550;
  assign n12820 = pi94  & n3735;
  assign n12821 = pi95  & n3545;
  assign n12822 = ~n12820 & ~n12821;
  assign n12823 = ~n12819 & n12822;
  assign n12824 = n3553 & n3921;
  assign n12825 = n12823 & ~n12824;
  assign n12826 = pi32  & ~n12825;
  assign n12827 = pi32  & ~n12826;
  assign n12828 = ~n12825 & ~n12826;
  assign n12829 = ~n12827 & ~n12828;
  assign n12830 = n12818 & ~n12829;
  assign n12831 = ~n12818 & n12829;
  assign n12832 = ~n12639 & ~n12831;
  assign n12833 = ~n12830 & n12832;
  assign n12834 = ~n12639 & ~n12833;
  assign n12835 = ~n12830 & ~n12833;
  assign n12836 = ~n12831 & n12835;
  assign n12837 = ~n12834 & ~n12836;
  assign n12838 = pi99  & n2976;
  assign n12839 = pi97  & n3182;
  assign n12840 = pi98  & n2971;
  assign n12841 = ~n12839 & ~n12840;
  assign n12842 = ~n12838 & n12841;
  assign n12843 = n2979 & n4584;
  assign n12844 = n12842 & ~n12843;
  assign n12845 = pi29  & ~n12844;
  assign n12846 = pi29  & ~n12845;
  assign n12847 = ~n12844 & ~n12845;
  assign n12848 = ~n12846 & ~n12847;
  assign n12849 = ~n12837 & ~n12848;
  assign n12850 = n12837 & n12848;
  assign n12851 = ~n12849 & ~n12850;
  assign n12852 = n12638 & ~n12851;
  assign n12853 = ~n12638 & n12851;
  assign n12854 = ~n12852 & ~n12853;
  assign n12855 = pi102  & n2486;
  assign n12856 = pi100  & n2644;
  assign n12857 = pi101  & n2481;
  assign n12858 = ~n12856 & ~n12857;
  assign n12859 = ~n12855 & n12858;
  assign n12860 = n2489 & n5296;
  assign n12861 = n12859 & ~n12860;
  assign n12862 = pi26  & ~n12861;
  assign n12863 = pi26  & ~n12862;
  assign n12864 = ~n12861 & ~n12862;
  assign n12865 = ~n12863 & ~n12864;
  assign n12866 = n12854 & ~n12865;
  assign n12867 = ~n12854 & n12865;
  assign n12868 = ~n12866 & ~n12867;
  assign n12869 = n12637 & ~n12868;
  assign n12870 = ~n12637 & n12868;
  assign n12871 = ~n12869 & ~n12870;
  assign n12872 = pi105  & n2004;
  assign n12873 = pi103  & n2141;
  assign n12874 = pi104  & n1999;
  assign n12875 = ~n12873 & ~n12874;
  assign n12876 = ~n12872 & n12875;
  assign n12877 = n2007 & n6065;
  assign n12878 = n12876 & ~n12877;
  assign n12879 = pi23  & ~n12878;
  assign n12880 = pi23  & ~n12879;
  assign n12881 = ~n12878 & ~n12879;
  assign n12882 = ~n12880 & ~n12881;
  assign n12883 = n12871 & ~n12882;
  assign n12884 = ~n12871 & n12882;
  assign n12885 = ~n12636 & ~n12884;
  assign n12886 = ~n12883 & n12885;
  assign n12887 = ~n12636 & ~n12886;
  assign n12888 = ~n12883 & ~n12886;
  assign n12889 = ~n12884 & n12888;
  assign n12890 = ~n12887 & ~n12889;
  assign n12891 = pi108  & n1582;
  assign n12892 = pi106  & n1713;
  assign n12893 = pi107  & n1577;
  assign n12894 = ~n12892 & ~n12893;
  assign n12895 = ~n12891 & n12894;
  assign n12896 = n1585 & n6639;
  assign n12897 = n12895 & ~n12896;
  assign n12898 = pi20  & ~n12897;
  assign n12899 = pi20  & ~n12898;
  assign n12900 = ~n12897 & ~n12898;
  assign n12901 = ~n12899 & ~n12900;
  assign n12902 = ~n12890 & ~n12901;
  assign n12903 = n12890 & n12901;
  assign n12904 = ~n12902 & ~n12903;
  assign n12905 = ~n12517 & n12904;
  assign n12906 = n12517 & ~n12904;
  assign n12907 = ~n12905 & ~n12906;
  assign n12908 = ~n12635 & n12907;
  assign n12909 = n12635 & ~n12907;
  assign n12910 = ~n12908 & ~n12909;
  assign n12911 = ~n12624 & n12910;
  assign n12912 = n12624 & ~n12910;
  assign n12913 = ~n12911 & ~n12912;
  assign n12914 = pi114  & n918;
  assign n12915 = pi112  & n1031;
  assign n12916 = pi113  & n913;
  assign n12917 = ~n12915 & ~n12916;
  assign n12918 = ~n12914 & n12917;
  assign n12919 = n921 & n8702;
  assign n12920 = n12918 & ~n12919;
  assign n12921 = pi14  & ~n12920;
  assign n12922 = pi14  & ~n12921;
  assign n12923 = ~n12920 & ~n12921;
  assign n12924 = ~n12922 & ~n12923;
  assign n12925 = n12913 & ~n12924;
  assign n12926 = ~n12913 & n12924;
  assign n12927 = ~n12925 & ~n12926;
  assign n12928 = ~n12623 & n12927;
  assign n12929 = n12623 & ~n12927;
  assign n12930 = ~n12928 & ~n12929;
  assign n12931 = ~n12622 & n12930;
  assign n12932 = n12622 & ~n12930;
  assign n12933 = ~n12931 & ~n12932;
  assign n12934 = ~n12611 & n12933;
  assign n12935 = n12611 & ~n12933;
  assign n12936 = ~n12934 & ~n12935;
  assign n12937 = pi120  & n493;
  assign n12938 = pi118  & n533;
  assign n12939 = pi119  & n488;
  assign n12940 = ~n12938 & ~n12939;
  assign n12941 = ~n12937 & n12940;
  assign n12942 = n496 & n10734;
  assign n12943 = n12941 & ~n12942;
  assign n12944 = pi8  & ~n12943;
  assign n12945 = pi8  & ~n12944;
  assign n12946 = ~n12943 & ~n12944;
  assign n12947 = ~n12945 & ~n12946;
  assign n12948 = ~n12936 & n12947;
  assign n12949 = n12936 & ~n12947;
  assign n12950 = ~n12948 & ~n12949;
  assign n12951 = pi123  & n340;
  assign n12952 = pi121  & n380;
  assign n12953 = pi122  & n335;
  assign n12954 = ~n12952 & ~n12953;
  assign n12955 = ~n12951 & n12954;
  assign n12956 = n343 & n11489;
  assign n12957 = n12955 & ~n12956;
  assign n12958 = pi5  & ~n12957;
  assign n12959 = pi5  & ~n12958;
  assign n12960 = ~n12957 & ~n12958;
  assign n12961 = ~n12959 & ~n12960;
  assign n12962 = n12950 & ~n12961;
  assign n12963 = ~n12950 & n12961;
  assign n12964 = ~n12962 & ~n12963;
  assign n12965 = n12610 & ~n12964;
  assign n12966 = ~n12610 & n12964;
  assign n12967 = ~n12965 & ~n12966;
  assign n12968 = pi126  & n264;
  assign n12969 = pi124  & n281;
  assign n12970 = pi125  & n259;
  assign n12971 = ~n12969 & ~n12970;
  assign n12972 = ~n12968 & n12971;
  assign n12973 = ~n12587 & ~n12589;
  assign n12974 = ~pi125  & ~pi126 ;
  assign n12975 = pi125  & pi126 ;
  assign n12976 = ~n12974 & ~n12975;
  assign n12977 = ~n12973 & n12976;
  assign n12978 = n12973 & ~n12976;
  assign n12979 = ~n12977 & ~n12978;
  assign n12980 = n267 & n12979;
  assign n12981 = n12972 & ~n12980;
  assign n12982 = pi2  & ~n12981;
  assign n12983 = pi2  & ~n12982;
  assign n12984 = ~n12981 & ~n12982;
  assign n12985 = ~n12983 & ~n12984;
  assign n12986 = ~n12967 & n12985;
  assign n12987 = n12967 & ~n12985;
  assign n12988 = ~n12986 & ~n12987;
  assign n12989 = ~n12609 & n12988;
  assign n12990 = n12609 & ~n12988;
  assign n12991 = ~n12989 & ~n12990;
  assign n12992 = ~n12608 & n12991;
  assign n12993 = n12608 & ~n12991;
  assign po62  = ~n12992 & ~n12993;
  assign n12995 = ~n12989 & ~n12992;
  assign n12996 = ~n12966 & ~n12987;
  assign n12997 = ~n12949 & ~n12962;
  assign n12998 = pi124  & n340;
  assign n12999 = pi122  & n380;
  assign n13000 = pi123  & n335;
  assign n13001 = ~n12999 & ~n13000;
  assign n13002 = ~n12998 & n13001;
  assign n13003 = n343 & n11858;
  assign n13004 = n13002 & ~n13003;
  assign n13005 = pi5  & ~n13004;
  assign n13006 = pi5  & ~n13005;
  assign n13007 = ~n13004 & ~n13005;
  assign n13008 = ~n13006 & ~n13007;
  assign n13009 = ~n12931 & ~n12934;
  assign n13010 = ~n12925 & ~n12928;
  assign n13011 = pi115  & n918;
  assign n13012 = pi113  & n1031;
  assign n13013 = pi114  & n913;
  assign n13014 = ~n13012 & ~n13013;
  assign n13015 = ~n13011 & n13014;
  assign n13016 = n921 & n8727;
  assign n13017 = n13015 & ~n13016;
  assign n13018 = pi14  & ~n13017;
  assign n13019 = pi14  & ~n13018;
  assign n13020 = ~n13017 & ~n13018;
  assign n13021 = ~n13019 & ~n13020;
  assign n13022 = ~n12908 & ~n12911;
  assign n13023 = pi112  & n1269;
  assign n13024 = pi110  & n1340;
  assign n13025 = pi111  & n1264;
  assign n13026 = ~n13024 & ~n13025;
  assign n13027 = ~n13023 & n13026;
  assign n13028 = n1272 & n7795;
  assign n13029 = n13027 & ~n13028;
  assign n13030 = pi17  & ~n13029;
  assign n13031 = pi17  & ~n13030;
  assign n13032 = ~n13029 & ~n13030;
  assign n13033 = ~n13031 & ~n13032;
  assign n13034 = ~n12902 & ~n12905;
  assign n13035 = pi109  & n1582;
  assign n13036 = pi107  & n1713;
  assign n13037 = pi108  & n1577;
  assign n13038 = ~n13036 & ~n13037;
  assign n13039 = ~n13035 & n13038;
  assign n13040 = n1585 & n7170;
  assign n13041 = n13039 & ~n13040;
  assign n13042 = pi20  & ~n13041;
  assign n13043 = pi20  & ~n13042;
  assign n13044 = ~n13041 & ~n13042;
  assign n13045 = ~n13043 & ~n13044;
  assign n13046 = pi106  & n2004;
  assign n13047 = pi104  & n2141;
  assign n13048 = pi105  & n1999;
  assign n13049 = ~n13047 & ~n13048;
  assign n13050 = ~n13046 & n13049;
  assign n13051 = n2007 & n6090;
  assign n13052 = n13050 & ~n13051;
  assign n13053 = pi23  & ~n13052;
  assign n13054 = pi23  & ~n13053;
  assign n13055 = ~n13052 & ~n13053;
  assign n13056 = ~n13054 & ~n13055;
  assign n13057 = ~n12866 & ~n12870;
  assign n13058 = ~n12849 & ~n12853;
  assign n13059 = pi100  & n2976;
  assign n13060 = pi98  & n3182;
  assign n13061 = pi99  & n2971;
  assign n13062 = ~n13060 & ~n13061;
  assign n13063 = ~n13059 & n13062;
  assign n13064 = n2979 & n4808;
  assign n13065 = n13063 & ~n13064;
  assign n13066 = pi29  & ~n13065;
  assign n13067 = pi29  & ~n13066;
  assign n13068 = ~n13065 & ~n13066;
  assign n13069 = ~n13067 & ~n13068;
  assign n13070 = ~n12796 & ~n12800;
  assign n13071 = ~n12779 & ~n12783;
  assign n13072 = ~n12773 & ~n12776;
  assign n13073 = pi85  & n6396;
  assign n13074 = pi83  & n6735;
  assign n13075 = pi84  & n6391;
  assign n13076 = ~n13074 & ~n13075;
  assign n13077 = ~n13073 & n13076;
  assign n13078 = n1943 & n6399;
  assign n13079 = n13077 & ~n13078;
  assign n13080 = pi44  & ~n13079;
  assign n13081 = pi44  & ~n13080;
  assign n13082 = ~n13079 & ~n13080;
  assign n13083 = ~n13081 & ~n13082;
  assign n13084 = ~n12767 & ~n12770;
  assign n13085 = ~n12744 & ~n12746;
  assign n13086 = pi76  & n9096;
  assign n13087 = pi74  & n9453;
  assign n13088 = pi75  & n9091;
  assign n13089 = ~n13087 & ~n13088;
  assign n13090 = ~n13086 & n13089;
  assign n13091 = n881 & n9099;
  assign n13092 = n13090 & ~n13091;
  assign n13093 = pi53  & ~n13092;
  assign n13094 = pi53  & ~n13093;
  assign n13095 = ~n13092 & ~n13093;
  assign n13096 = ~n13094 & ~n13095;
  assign n13097 = ~n12738 & ~n12740;
  assign n13098 = pi70  & n11193;
  assign n13099 = pi68  & n11567;
  assign n13100 = pi69  & n11188;
  assign n13101 = ~n13099 & ~n13100;
  assign n13102 = ~n13098 & n13101;
  assign n13103 = n430 & n11196;
  assign n13104 = n13102 & ~n13103;
  assign n13105 = pi59  & ~n13104;
  assign n13106 = pi59  & ~n13105;
  assign n13107 = ~n13104 & ~n13105;
  assign n13108 = ~n13106 & ~n13107;
  assign n13109 = pi67  & n12295;
  assign n13110 = pi65  & n12693;
  assign n13111 = pi66  & n12290;
  assign n13112 = ~n13110 & ~n13111;
  assign n13113 = ~n13109 & n13112;
  assign n13114 = n313 & n12298;
  assign n13115 = n13113 & ~n13114;
  assign n13116 = pi62  & ~n13115;
  assign n13117 = pi62  & ~n13116;
  assign n13118 = ~n13115 & ~n13116;
  assign n13119 = ~n13117 & ~n13118;
  assign n13120 = pi62  & ~pi63 ;
  assign n13121 = ~pi62  & pi63 ;
  assign n13122 = ~n13120 & ~n13121;
  assign n13123 = pi64  & ~n13122;
  assign n13124 = n12705 & n13123;
  assign n13125 = ~n12705 & ~n13123;
  assign n13126 = ~n13124 & ~n13125;
  assign n13127 = ~n13119 & n13126;
  assign n13128 = n13119 & ~n13126;
  assign n13129 = ~n13127 & ~n13128;
  assign n13130 = n13108 & ~n13129;
  assign n13131 = ~n13108 & n13129;
  assign n13132 = ~n13130 & ~n13131;
  assign n13133 = ~n12723 & n13132;
  assign n13134 = n12723 & ~n13132;
  assign n13135 = ~n13133 & ~n13134;
  assign n13136 = pi73  & n10135;
  assign n13137 = pi71  & n10478;
  assign n13138 = pi72  & n10130;
  assign n13139 = ~n13137 & ~n13138;
  assign n13140 = ~n13136 & n13139;
  assign n13141 = n639 & n10138;
  assign n13142 = n13140 & ~n13141;
  assign n13143 = pi56  & ~n13142;
  assign n13144 = pi56  & ~n13143;
  assign n13145 = ~n13142 & ~n13143;
  assign n13146 = ~n13144 & ~n13145;
  assign n13147 = n13135 & ~n13146;
  assign n13148 = ~n13135 & n13146;
  assign n13149 = ~n13147 & ~n13148;
  assign n13150 = ~n13097 & n13149;
  assign n13151 = n13097 & ~n13149;
  assign n13152 = ~n13150 & ~n13151;
  assign n13153 = n13096 & ~n13152;
  assign n13154 = ~n13096 & n13152;
  assign n13155 = ~n13153 & ~n13154;
  assign n13156 = ~n13085 & n13155;
  assign n13157 = n13085 & ~n13155;
  assign n13158 = ~n13156 & ~n13157;
  assign n13159 = pi79  & n8137;
  assign n13160 = pi77  & n8471;
  assign n13161 = pi78  & n8132;
  assign n13162 = ~n13160 & ~n13161;
  assign n13163 = ~n13159 & n13162;
  assign n13164 = n1105 & n8140;
  assign n13165 = n13163 & ~n13164;
  assign n13166 = pi50  & ~n13165;
  assign n13167 = pi50  & ~n13166;
  assign n13168 = ~n13165 & ~n13166;
  assign n13169 = ~n13167 & ~n13168;
  assign n13170 = n13158 & ~n13169;
  assign n13171 = n13158 & ~n13170;
  assign n13172 = ~n13169 & ~n13170;
  assign n13173 = ~n13171 & ~n13172;
  assign n13174 = ~n12760 & ~n12764;
  assign n13175 = n13173 & n13174;
  assign n13176 = ~n13173 & ~n13174;
  assign n13177 = ~n13175 & ~n13176;
  assign n13178 = pi82  & n7239;
  assign n13179 = pi80  & n7556;
  assign n13180 = pi81  & n7234;
  assign n13181 = ~n13179 & ~n13180;
  assign n13182 = ~n13178 & n13181;
  assign n13183 = n1532 & n7242;
  assign n13184 = n13182 & ~n13183;
  assign n13185 = pi47  & ~n13184;
  assign n13186 = pi47  & ~n13185;
  assign n13187 = ~n13184 & ~n13185;
  assign n13188 = ~n13186 & ~n13187;
  assign n13189 = ~n13177 & n13188;
  assign n13190 = n13177 & ~n13188;
  assign n13191 = ~n13189 & ~n13190;
  assign n13192 = ~n13084 & n13191;
  assign n13193 = n13084 & ~n13191;
  assign n13194 = ~n13192 & ~n13193;
  assign n13195 = ~n13083 & n13194;
  assign n13196 = n13083 & ~n13194;
  assign n13197 = ~n13195 & ~n13196;
  assign n13198 = ~n13072 & n13197;
  assign n13199 = n13072 & ~n13197;
  assign n13200 = ~n13198 & ~n13199;
  assign n13201 = pi88  & n5636;
  assign n13202 = pi86  & n5909;
  assign n13203 = pi87  & n5631;
  assign n13204 = ~n13202 & ~n13203;
  assign n13205 = ~n13201 & n13204;
  assign n13206 = n2277 & n5639;
  assign n13207 = n13205 & ~n13206;
  assign n13208 = pi41  & ~n13207;
  assign n13209 = pi41  & ~n13208;
  assign n13210 = ~n13207 & ~n13208;
  assign n13211 = ~n13209 & ~n13210;
  assign n13212 = n13200 & ~n13211;
  assign n13213 = ~n13200 & n13211;
  assign n13214 = ~n13212 & ~n13213;
  assign n13215 = n13071 & ~n13214;
  assign n13216 = ~n13071 & n13214;
  assign n13217 = ~n13215 & ~n13216;
  assign n13218 = pi91  & n4896;
  assign n13219 = pi89  & n5148;
  assign n13220 = pi90  & n4891;
  assign n13221 = ~n13219 & ~n13220;
  assign n13222 = ~n13218 & n13221;
  assign n13223 = n2926 & n4899;
  assign n13224 = n13222 & ~n13223;
  assign n13225 = pi38  & ~n13224;
  assign n13226 = pi38  & ~n13225;
  assign n13227 = ~n13224 & ~n13225;
  assign n13228 = ~n13226 & ~n13227;
  assign n13229 = n13217 & ~n13228;
  assign n13230 = ~n13217 & n13228;
  assign n13231 = ~n13229 & ~n13230;
  assign n13232 = n13070 & ~n13231;
  assign n13233 = ~n13070 & n13231;
  assign n13234 = ~n13232 & ~n13233;
  assign n13235 = pi94  & n4182;
  assign n13236 = pi92  & n4416;
  assign n13237 = pi93  & n4177;
  assign n13238 = ~n13236 & ~n13237;
  assign n13239 = ~n13235 & n13238;
  assign n13240 = n3499 & n4185;
  assign n13241 = n13239 & ~n13240;
  assign n13242 = pi35  & ~n13241;
  assign n13243 = pi35  & ~n13242;
  assign n13244 = ~n13241 & ~n13242;
  assign n13245 = ~n13243 & ~n13244;
  assign n13246 = ~n13234 & n13245;
  assign n13247 = n13234 & ~n13245;
  assign n13248 = ~n13246 & ~n13247;
  assign n13249 = ~n12813 & ~n12817;
  assign n13250 = n13248 & ~n13249;
  assign n13251 = ~n13248 & n13249;
  assign n13252 = ~n13250 & ~n13251;
  assign n13253 = pi97  & n3550;
  assign n13254 = pi95  & n3735;
  assign n13255 = pi96  & n3545;
  assign n13256 = ~n13254 & ~n13255;
  assign n13257 = ~n13253 & n13256;
  assign n13258 = n3553 & n3946;
  assign n13259 = n13257 & ~n13258;
  assign n13260 = pi32  & ~n13259;
  assign n13261 = pi32  & ~n13260;
  assign n13262 = ~n13259 & ~n13260;
  assign n13263 = ~n13261 & ~n13262;
  assign n13264 = n13252 & ~n13263;
  assign n13265 = ~n13252 & n13263;
  assign n13266 = ~n13264 & ~n13265;
  assign n13267 = ~n12835 & n13266;
  assign n13268 = n12835 & ~n13266;
  assign n13269 = ~n13267 & ~n13268;
  assign n13270 = ~n13069 & n13269;
  assign n13271 = n13069 & ~n13269;
  assign n13272 = ~n13270 & ~n13271;
  assign n13273 = n13058 & ~n13272;
  assign n13274 = ~n13058 & n13272;
  assign n13275 = ~n13273 & ~n13274;
  assign n13276 = pi103  & n2486;
  assign n13277 = pi101  & n2644;
  assign n13278 = pi102  & n2481;
  assign n13279 = ~n13277 & ~n13278;
  assign n13280 = ~n13276 & n13279;
  assign n13281 = n2489 & n5540;
  assign n13282 = n13280 & ~n13281;
  assign n13283 = pi26  & ~n13282;
  assign n13284 = pi26  & ~n13283;
  assign n13285 = ~n13282 & ~n13283;
  assign n13286 = ~n13284 & ~n13285;
  assign n13287 = ~n13275 & n13286;
  assign n13288 = n13275 & ~n13286;
  assign n13289 = ~n13287 & ~n13288;
  assign n13290 = ~n13057 & n13289;
  assign n13291 = n13057 & ~n13289;
  assign n13292 = ~n13290 & ~n13291;
  assign n13293 = ~n13056 & n13292;
  assign n13294 = n13056 & ~n13292;
  assign n13295 = ~n13293 & ~n13294;
  assign n13296 = ~n12888 & n13295;
  assign n13297 = n12888 & ~n13295;
  assign n13298 = ~n13296 & ~n13297;
  assign n13299 = ~n13045 & n13298;
  assign n13300 = n13045 & ~n13298;
  assign n13301 = ~n13299 & ~n13300;
  assign n13302 = ~n13034 & n13301;
  assign n13303 = n13034 & ~n13301;
  assign n13304 = ~n13302 & ~n13303;
  assign n13305 = ~n13033 & n13304;
  assign n13306 = n13033 & ~n13304;
  assign n13307 = ~n13305 & ~n13306;
  assign n13308 = ~n13022 & n13307;
  assign n13309 = n13022 & ~n13307;
  assign n13310 = ~n13308 & ~n13309;
  assign n13311 = ~n13021 & n13310;
  assign n13312 = n13021 & ~n13310;
  assign n13313 = ~n13311 & ~n13312;
  assign n13314 = ~n13010 & n13313;
  assign n13315 = n13010 & ~n13313;
  assign n13316 = ~n13314 & ~n13315;
  assign n13317 = pi118  & n675;
  assign n13318 = pi116  & n769;
  assign n13319 = pi117  & n670;
  assign n13320 = ~n13318 & ~n13319;
  assign n13321 = ~n13317 & n13320;
  assign n13322 = n678 & n9716;
  assign n13323 = n13321 & ~n13322;
  assign n13324 = pi11  & ~n13323;
  assign n13325 = pi11  & ~n13324;
  assign n13326 = ~n13323 & ~n13324;
  assign n13327 = ~n13325 & ~n13326;
  assign n13328 = n13316 & ~n13327;
  assign n13329 = ~n13316 & n13327;
  assign n13330 = ~n13328 & ~n13329;
  assign n13331 = n13009 & ~n13330;
  assign n13332 = ~n13009 & n13330;
  assign n13333 = ~n13331 & ~n13332;
  assign n13334 = pi121  & n493;
  assign n13335 = pi119  & n533;
  assign n13336 = pi120  & n488;
  assign n13337 = ~n13335 & ~n13336;
  assign n13338 = ~n13334 & n13337;
  assign n13339 = n496 & n11086;
  assign n13340 = n13338 & ~n13339;
  assign n13341 = pi8  & ~n13340;
  assign n13342 = pi8  & ~n13341;
  assign n13343 = ~n13340 & ~n13341;
  assign n13344 = ~n13342 & ~n13343;
  assign n13345 = n13333 & ~n13344;
  assign n13346 = ~n13333 & n13344;
  assign n13347 = ~n13345 & ~n13346;
  assign n13348 = ~n13008 & n13347;
  assign n13349 = n13008 & ~n13347;
  assign n13350 = ~n13348 & ~n13349;
  assign n13351 = n12997 & ~n13350;
  assign n13352 = ~n12997 & n13350;
  assign n13353 = ~n13351 & ~n13352;
  assign n13354 = pi127  & n264;
  assign n13355 = pi125  & n281;
  assign n13356 = pi126  & n259;
  assign n13357 = ~n13355 & ~n13356;
  assign n13358 = ~n13354 & n13357;
  assign n13359 = ~n12975 & ~n12977;
  assign n13360 = pi126  & ~pi127 ;
  assign n13361 = ~pi126  & pi127 ;
  assign n13362 = ~n13360 & ~n13361;
  assign n13363 = ~n13359 & ~n13362;
  assign n13364 = n13359 & n13362;
  assign n13365 = ~n13363 & ~n13364;
  assign n13366 = n267 & n13365;
  assign n13367 = n13358 & ~n13366;
  assign n13368 = pi2  & ~n13367;
  assign n13369 = pi2  & ~n13368;
  assign n13370 = ~n13367 & ~n13368;
  assign n13371 = ~n13369 & ~n13370;
  assign n13372 = n13353 & ~n13371;
  assign n13373 = ~n13353 & n13371;
  assign n13374 = ~n13372 & ~n13373;
  assign n13375 = ~n12996 & n13374;
  assign n13376 = n12996 & ~n13374;
  assign n13377 = ~n13375 & ~n13376;
  assign n13378 = ~n12995 & n13377;
  assign n13379 = n12995 & ~n13377;
  assign po63  = ~n13378 & ~n13379;
  assign n13381 = ~n13375 & ~n13378;
  assign n13382 = ~n13352 & ~n13372;
  assign n13383 = pi126  & n281;
  assign n13384 = pi127  & n259;
  assign n13385 = ~n13383 & ~n13384;
  assign n13386 = ~pi126  & ~n13363;
  assign n13387 = pi127  & ~n13386;
  assign n13388 = ~pi127  & ~n13363;
  assign n13389 = ~n13387 & ~n13388;
  assign n13390 = n267 & n13389;
  assign n13391 = n13385 & ~n13390;
  assign n13392 = pi2  & ~n13391;
  assign n13393 = pi2  & ~n13392;
  assign n13394 = ~n13391 & ~n13392;
  assign n13395 = ~n13393 & ~n13394;
  assign n13396 = ~n13345 & ~n13348;
  assign n13397 = pi125  & n340;
  assign n13398 = pi123  & n380;
  assign n13399 = pi124  & n335;
  assign n13400 = ~n13398 & ~n13399;
  assign n13401 = ~n13397 & n13400;
  assign n13402 = n343 & n12591;
  assign n13403 = n13401 & ~n13402;
  assign n13404 = pi5  & ~n13403;
  assign n13405 = pi5  & ~n13404;
  assign n13406 = ~n13403 & ~n13404;
  assign n13407 = ~n13405 & ~n13406;
  assign n13408 = ~n13328 & ~n13332;
  assign n13409 = pi119  & n675;
  assign n13410 = pi117  & n769;
  assign n13411 = pi118  & n670;
  assign n13412 = ~n13410 & ~n13411;
  assign n13413 = ~n13409 & n13412;
  assign n13414 = n678 & n10048;
  assign n13415 = n13413 & ~n13414;
  assign n13416 = pi11  & ~n13415;
  assign n13417 = pi11  & ~n13416;
  assign n13418 = ~n13415 & ~n13416;
  assign n13419 = ~n13417 & ~n13418;
  assign n13420 = ~n13311 & ~n13314;
  assign n13421 = pi116  & n918;
  assign n13422 = pi114  & n1031;
  assign n13423 = pi115  & n913;
  assign n13424 = ~n13422 & ~n13423;
  assign n13425 = ~n13421 & n13424;
  assign n13426 = n921 & n9042;
  assign n13427 = n13425 & ~n13426;
  assign n13428 = pi14  & ~n13427;
  assign n13429 = pi14  & ~n13428;
  assign n13430 = ~n13427 & ~n13428;
  assign n13431 = ~n13429 & ~n13430;
  assign n13432 = ~n13305 & ~n13308;
  assign n13433 = pi113  & n1269;
  assign n13434 = pi111  & n1340;
  assign n13435 = pi112  & n1264;
  assign n13436 = ~n13434 & ~n13435;
  assign n13437 = ~n13433 & n13436;
  assign n13438 = n1272 & n8387;
  assign n13439 = n13437 & ~n13438;
  assign n13440 = pi17  & ~n13439;
  assign n13441 = pi17  & ~n13440;
  assign n13442 = ~n13439 & ~n13440;
  assign n13443 = ~n13441 & ~n13442;
  assign n13444 = ~n13299 & ~n13302;
  assign n13445 = pi110  & n1582;
  assign n13446 = pi108  & n1713;
  assign n13447 = pi109  & n1577;
  assign n13448 = ~n13446 & ~n13447;
  assign n13449 = ~n13445 & n13448;
  assign n13450 = n1585 & n7474;
  assign n13451 = n13449 & ~n13450;
  assign n13452 = pi20  & ~n13451;
  assign n13453 = pi20  & ~n13452;
  assign n13454 = ~n13451 & ~n13452;
  assign n13455 = ~n13453 & ~n13454;
  assign n13456 = ~n13293 & ~n13296;
  assign n13457 = pi107  & n2004;
  assign n13458 = pi105  & n2141;
  assign n13459 = pi106  & n1999;
  assign n13460 = ~n13458 & ~n13459;
  assign n13461 = ~n13457 & n13460;
  assign n13462 = n2007 & n6614;
  assign n13463 = n13461 & ~n13462;
  assign n13464 = pi23  & ~n13463;
  assign n13465 = pi23  & ~n13464;
  assign n13466 = ~n13463 & ~n13464;
  assign n13467 = ~n13465 & ~n13466;
  assign n13468 = ~n13288 & ~n13290;
  assign n13469 = ~n13270 & ~n13274;
  assign n13470 = ~n13264 & ~n13267;
  assign n13471 = ~n13229 & ~n13233;
  assign n13472 = ~n13212 & ~n13216;
  assign n13473 = ~n13195 & ~n13198;
  assign n13474 = ~n13147 & ~n13150;
  assign n13475 = ~n13131 & ~n13133;
  assign n13476 = ~n13124 & ~n13127;
  assign n13477 = pi63  & n13122;
  assign n13478 = pi64  & n13477;
  assign n13479 = pi65  & ~n13122;
  assign n13480 = ~n13478 & ~n13479;
  assign n13481 = pi68  & n12295;
  assign n13482 = pi66  & n12693;
  assign n13483 = pi67  & n12290;
  assign n13484 = ~n13482 & ~n13483;
  assign n13485 = ~n13481 & n13484;
  assign n13486 = n364 & n12298;
  assign n13487 = n13485 & ~n13486;
  assign n13488 = pi62  & ~n13487;
  assign n13489 = pi62  & ~n13488;
  assign n13490 = ~n13487 & ~n13488;
  assign n13491 = ~n13489 & ~n13490;
  assign n13492 = ~n13480 & ~n13491;
  assign n13493 = n13480 & n13491;
  assign n13494 = ~n13492 & ~n13493;
  assign n13495 = n13476 & ~n13494;
  assign n13496 = ~n13476 & n13494;
  assign n13497 = ~n13495 & ~n13496;
  assign n13498 = pi71  & n11193;
  assign n13499 = pi69  & n11567;
  assign n13500 = pi70  & n11188;
  assign n13501 = ~n13499 & ~n13500;
  assign n13502 = ~n13498 & n13501;
  assign n13503 = n476 & n11196;
  assign n13504 = n13502 & ~n13503;
  assign n13505 = pi59  & ~n13504;
  assign n13506 = pi59  & ~n13505;
  assign n13507 = ~n13504 & ~n13505;
  assign n13508 = ~n13506 & ~n13507;
  assign n13509 = ~n13497 & n13508;
  assign n13510 = n13497 & ~n13508;
  assign n13511 = ~n13509 & ~n13510;
  assign n13512 = ~n13475 & n13511;
  assign n13513 = n13475 & ~n13511;
  assign n13514 = ~n13512 & ~n13513;
  assign n13515 = pi74  & n10135;
  assign n13516 = pi72  & n10478;
  assign n13517 = pi73  & n10130;
  assign n13518 = ~n13516 & ~n13517;
  assign n13519 = ~n13515 & n13518;
  assign n13520 = n722 & n10138;
  assign n13521 = n13519 & ~n13520;
  assign n13522 = pi56  & ~n13521;
  assign n13523 = pi56  & ~n13522;
  assign n13524 = ~n13521 & ~n13522;
  assign n13525 = ~n13523 & ~n13524;
  assign n13526 = n13514 & ~n13525;
  assign n13527 = ~n13514 & n13525;
  assign n13528 = ~n13526 & ~n13527;
  assign n13529 = n13474 & ~n13528;
  assign n13530 = ~n13474 & n13528;
  assign n13531 = ~n13529 & ~n13530;
  assign n13532 = pi77  & n9096;
  assign n13533 = pi75  & n9453;
  assign n13534 = pi76  & n9091;
  assign n13535 = ~n13533 & ~n13534;
  assign n13536 = ~n13532 & n13535;
  assign n13537 = n984 & n9099;
  assign n13538 = n13536 & ~n13537;
  assign n13539 = pi53  & ~n13538;
  assign n13540 = pi53  & ~n13539;
  assign n13541 = ~n13538 & ~n13539;
  assign n13542 = ~n13540 & ~n13541;
  assign n13543 = ~n13531 & n13542;
  assign n13544 = n13531 & ~n13542;
  assign n13545 = ~n13543 & ~n13544;
  assign n13546 = ~n13154 & ~n13156;
  assign n13547 = n13545 & ~n13546;
  assign n13548 = ~n13545 & n13546;
  assign n13549 = ~n13547 & ~n13548;
  assign n13550 = pi80  & n8137;
  assign n13551 = pi78  & n8471;
  assign n13552 = pi79  & n8132;
  assign n13553 = ~n13551 & ~n13552;
  assign n13554 = ~n13550 & n13553;
  assign n13555 = n1205 & n8140;
  assign n13556 = n13554 & ~n13555;
  assign n13557 = pi50  & ~n13556;
  assign n13558 = pi50  & ~n13557;
  assign n13559 = ~n13556 & ~n13557;
  assign n13560 = ~n13558 & ~n13559;
  assign n13561 = n13549 & ~n13560;
  assign n13562 = n13549 & ~n13561;
  assign n13563 = ~n13560 & ~n13561;
  assign n13564 = ~n13562 & ~n13563;
  assign n13565 = ~n13170 & ~n13176;
  assign n13566 = n13564 & n13565;
  assign n13567 = ~n13564 & ~n13565;
  assign n13568 = ~n13566 & ~n13567;
  assign n13569 = pi83  & n7239;
  assign n13570 = pi81  & n7556;
  assign n13571 = pi82  & n7234;
  assign n13572 = ~n13570 & ~n13571;
  assign n13573 = ~n13569 & n13572;
  assign n13574 = n1672 & n7242;
  assign n13575 = n13573 & ~n13574;
  assign n13576 = pi47  & ~n13575;
  assign n13577 = pi47  & ~n13576;
  assign n13578 = ~n13575 & ~n13576;
  assign n13579 = ~n13577 & ~n13578;
  assign n13580 = ~n13568 & n13579;
  assign n13581 = n13568 & ~n13579;
  assign n13582 = ~n13580 & ~n13581;
  assign n13583 = ~n13190 & ~n13192;
  assign n13584 = n13582 & ~n13583;
  assign n13585 = ~n13582 & n13583;
  assign n13586 = ~n13584 & ~n13585;
  assign n13587 = pi86  & n6396;
  assign n13588 = pi84  & n6735;
  assign n13589 = pi85  & n6391;
  assign n13590 = ~n13588 & ~n13589;
  assign n13591 = ~n13587 & n13590;
  assign n13592 = n2099 & n6399;
  assign n13593 = n13591 & ~n13592;
  assign n13594 = pi44  & ~n13593;
  assign n13595 = pi44  & ~n13594;
  assign n13596 = ~n13593 & ~n13594;
  assign n13597 = ~n13595 & ~n13596;
  assign n13598 = n13586 & ~n13597;
  assign n13599 = ~n13586 & n13597;
  assign n13600 = ~n13598 & ~n13599;
  assign n13601 = n13473 & ~n13600;
  assign n13602 = ~n13473 & n13600;
  assign n13603 = ~n13601 & ~n13602;
  assign n13604 = pi89  & n5636;
  assign n13605 = pi87  & n5909;
  assign n13606 = pi88  & n5631;
  assign n13607 = ~n13605 & ~n13606;
  assign n13608 = ~n13604 & n13607;
  assign n13609 = n2432 & n5639;
  assign n13610 = n13608 & ~n13609;
  assign n13611 = pi41  & ~n13610;
  assign n13612 = pi41  & ~n13611;
  assign n13613 = ~n13610 & ~n13611;
  assign n13614 = ~n13612 & ~n13613;
  assign n13615 = n13603 & ~n13614;
  assign n13616 = ~n13603 & n13614;
  assign n13617 = ~n13615 & ~n13616;
  assign n13618 = n13472 & ~n13617;
  assign n13619 = ~n13472 & n13617;
  assign n13620 = ~n13618 & ~n13619;
  assign n13621 = pi92  & n4896;
  assign n13622 = pi90  & n5148;
  assign n13623 = pi91  & n4891;
  assign n13624 = ~n13622 & ~n13623;
  assign n13625 = ~n13621 & n13624;
  assign n13626 = n3119 & n4899;
  assign n13627 = n13625 & ~n13626;
  assign n13628 = pi38  & ~n13627;
  assign n13629 = pi38  & ~n13628;
  assign n13630 = ~n13627 & ~n13628;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = n13620 & ~n13631;
  assign n13633 = ~n13620 & n13631;
  assign n13634 = ~n13632 & ~n13633;
  assign n13635 = n13471 & ~n13634;
  assign n13636 = ~n13471 & n13634;
  assign n13637 = ~n13635 & ~n13636;
  assign n13638 = pi95  & n4182;
  assign n13639 = pi93  & n4416;
  assign n13640 = pi94  & n4177;
  assign n13641 = ~n13639 & ~n13640;
  assign n13642 = ~n13638 & n13641;
  assign n13643 = n3710 & n4185;
  assign n13644 = n13642 & ~n13643;
  assign n13645 = pi35  & ~n13644;
  assign n13646 = pi35  & ~n13645;
  assign n13647 = ~n13644 & ~n13645;
  assign n13648 = ~n13646 & ~n13647;
  assign n13649 = ~n13637 & n13648;
  assign n13650 = n13637 & ~n13648;
  assign n13651 = ~n13649 & ~n13650;
  assign n13652 = ~n13247 & ~n13250;
  assign n13653 = n13651 & ~n13652;
  assign n13654 = ~n13651 & n13652;
  assign n13655 = ~n13653 & ~n13654;
  assign n13656 = pi98  & n3550;
  assign n13657 = pi96  & n3735;
  assign n13658 = pi97  & n3545;
  assign n13659 = ~n13657 & ~n13658;
  assign n13660 = ~n13656 & n13659;
  assign n13661 = n3553 & n4360;
  assign n13662 = n13660 & ~n13661;
  assign n13663 = pi32  & ~n13662;
  assign n13664 = pi32  & ~n13663;
  assign n13665 = ~n13662 & ~n13663;
  assign n13666 = ~n13664 & ~n13665;
  assign n13667 = n13655 & ~n13666;
  assign n13668 = ~n13655 & n13666;
  assign n13669 = ~n13667 & ~n13668;
  assign n13670 = n13470 & ~n13669;
  assign n13671 = ~n13470 & n13669;
  assign n13672 = ~n13670 & ~n13671;
  assign n13673 = pi101  & n2976;
  assign n13674 = pi99  & n3182;
  assign n13675 = pi100  & n2971;
  assign n13676 = ~n13674 & ~n13675;
  assign n13677 = ~n13673 & n13676;
  assign n13678 = n2979 & n5056;
  assign n13679 = n13677 & ~n13678;
  assign n13680 = pi29  & ~n13679;
  assign n13681 = pi29  & ~n13680;
  assign n13682 = ~n13679 & ~n13680;
  assign n13683 = ~n13681 & ~n13682;
  assign n13684 = n13672 & ~n13683;
  assign n13685 = ~n13672 & n13683;
  assign n13686 = ~n13684 & ~n13685;
  assign n13687 = n13469 & ~n13686;
  assign n13688 = ~n13469 & n13686;
  assign n13689 = ~n13687 & ~n13688;
  assign n13690 = pi104  & n2486;
  assign n13691 = pi102  & n2644;
  assign n13692 = pi103  & n2481;
  assign n13693 = ~n13691 & ~n13692;
  assign n13694 = ~n13690 & n13693;
  assign n13695 = n2489 & n5565;
  assign n13696 = n13694 & ~n13695;
  assign n13697 = pi26  & ~n13696;
  assign n13698 = pi26  & ~n13697;
  assign n13699 = ~n13696 & ~n13697;
  assign n13700 = ~n13698 & ~n13699;
  assign n13701 = n13689 & ~n13700;
  assign n13702 = ~n13689 & n13700;
  assign n13703 = ~n13701 & ~n13702;
  assign n13704 = ~n13468 & n13703;
  assign n13705 = n13468 & ~n13703;
  assign n13706 = ~n13704 & ~n13705;
  assign n13707 = ~n13467 & n13706;
  assign n13708 = n13467 & ~n13706;
  assign n13709 = ~n13707 & ~n13708;
  assign n13710 = ~n13456 & n13709;
  assign n13711 = n13456 & ~n13709;
  assign n13712 = ~n13710 & ~n13711;
  assign n13713 = ~n13455 & n13712;
  assign n13714 = n13455 & ~n13712;
  assign n13715 = ~n13713 & ~n13714;
  assign n13716 = ~n13444 & n13715;
  assign n13717 = n13444 & ~n13715;
  assign n13718 = ~n13716 & ~n13717;
  assign n13719 = ~n13443 & n13718;
  assign n13720 = n13443 & ~n13718;
  assign n13721 = ~n13719 & ~n13720;
  assign n13722 = ~n13432 & n13721;
  assign n13723 = n13432 & ~n13721;
  assign n13724 = ~n13722 & ~n13723;
  assign n13725 = ~n13431 & n13724;
  assign n13726 = n13431 & ~n13724;
  assign n13727 = ~n13725 & ~n13726;
  assign n13728 = ~n13420 & n13727;
  assign n13729 = n13420 & ~n13727;
  assign n13730 = ~n13728 & ~n13729;
  assign n13731 = ~n13419 & n13730;
  assign n13732 = n13419 & ~n13730;
  assign n13733 = ~n13731 & ~n13732;
  assign n13734 = ~n13408 & n13733;
  assign n13735 = n13408 & ~n13733;
  assign n13736 = ~n13734 & ~n13735;
  assign n13737 = pi122  & n493;
  assign n13738 = pi120  & n533;
  assign n13739 = pi121  & n488;
  assign n13740 = ~n13738 & ~n13739;
  assign n13741 = ~n13737 & n13740;
  assign n13742 = n496 & n11463;
  assign n13743 = n13741 & ~n13742;
  assign n13744 = pi8  & ~n13743;
  assign n13745 = pi8  & ~n13744;
  assign n13746 = ~n13743 & ~n13744;
  assign n13747 = ~n13745 & ~n13746;
  assign n13748 = n13736 & ~n13747;
  assign n13749 = ~n13736 & n13747;
  assign n13750 = ~n13748 & ~n13749;
  assign n13751 = ~n13407 & n13750;
  assign n13752 = n13407 & ~n13750;
  assign n13753 = ~n13751 & ~n13752;
  assign n13754 = ~n13396 & n13753;
  assign n13755 = n13396 & ~n13753;
  assign n13756 = ~n13754 & ~n13755;
  assign n13757 = ~n13395 & n13756;
  assign n13758 = n13395 & ~n13756;
  assign n13759 = ~n13757 & ~n13758;
  assign n13760 = ~n13382 & n13759;
  assign n13761 = n13382 & ~n13759;
  assign n13762 = ~n13760 & ~n13761;
  assign n13763 = ~n13381 & n13762;
  assign n13764 = n13381 & ~n13762;
  assign po64  = ~n13763 & ~n13764;
  assign n13766 = ~n13754 & ~n13757;
  assign n13767 = ~n13748 & ~n13751;
  assign n13768 = n267 & n13387;
  assign n13769 = ~pi2  & ~n13768;
  assign n13770 = pi127  & n281;
  assign n13771 = ~n13768 & ~n13770;
  assign n13772 = pi2  & ~n13771;
  assign n13773 = ~n13769 & ~n13772;
  assign n13774 = ~n13767 & n13773;
  assign n13775 = n13767 & ~n13773;
  assign n13776 = ~n13774 & ~n13775;
  assign n13777 = ~n13731 & ~n13734;
  assign n13778 = ~n13725 & ~n13728;
  assign n13779 = ~n13719 & ~n13722;
  assign n13780 = pi114  & n1269;
  assign n13781 = pi112  & n1340;
  assign n13782 = pi113  & n1264;
  assign n13783 = ~n13781 & ~n13782;
  assign n13784 = ~n13780 & n13783;
  assign n13785 = n1272 & n8702;
  assign n13786 = n13784 & ~n13785;
  assign n13787 = pi17  & ~n13786;
  assign n13788 = pi17  & ~n13787;
  assign n13789 = ~n13786 & ~n13787;
  assign n13790 = ~n13788 & ~n13789;
  assign n13791 = ~n13713 & ~n13716;
  assign n13792 = pi111  & n1582;
  assign n13793 = pi109  & n1713;
  assign n13794 = pi110  & n1577;
  assign n13795 = ~n13793 & ~n13794;
  assign n13796 = ~n13792 & n13795;
  assign n13797 = n1585 & n7770;
  assign n13798 = n13796 & ~n13797;
  assign n13799 = pi20  & ~n13798;
  assign n13800 = pi20  & ~n13799;
  assign n13801 = ~n13798 & ~n13799;
  assign n13802 = ~n13800 & ~n13801;
  assign n13803 = ~n13707 & ~n13710;
  assign n13804 = ~n13701 & ~n13704;
  assign n13805 = ~n13684 & ~n13688;
  assign n13806 = ~n13667 & ~n13671;
  assign n13807 = ~n13650 & ~n13653;
  assign n13808 = ~n13632 & ~n13636;
  assign n13809 = ~n13615 & ~n13619;
  assign n13810 = ~n13598 & ~n13602;
  assign n13811 = pi87  & n6396;
  assign n13812 = pi85  & n6735;
  assign n13813 = pi86  & n6391;
  assign n13814 = ~n13812 & ~n13813;
  assign n13815 = ~n13811 & n13814;
  assign n13816 = n2252 & n6399;
  assign n13817 = n13815 & ~n13816;
  assign n13818 = pi44  & ~n13817;
  assign n13819 = pi44  & ~n13818;
  assign n13820 = ~n13817 & ~n13818;
  assign n13821 = ~n13819 & ~n13820;
  assign n13822 = ~n13581 & ~n13584;
  assign n13823 = ~n13561 & ~n13567;
  assign n13824 = pi81  & n8137;
  assign n13825 = pi79  & n8471;
  assign n13826 = pi80  & n8132;
  assign n13827 = ~n13825 & ~n13826;
  assign n13828 = ~n13824 & n13827;
  assign n13829 = n1413 & n8140;
  assign n13830 = n13828 & ~n13829;
  assign n13831 = pi50  & ~n13830;
  assign n13832 = pi50  & ~n13831;
  assign n13833 = ~n13830 & ~n13831;
  assign n13834 = ~n13832 & ~n13833;
  assign n13835 = ~n13544 & ~n13547;
  assign n13836 = ~n13526 & ~n13530;
  assign n13837 = ~n13510 & ~n13512;
  assign n13838 = ~n13492 & ~n13496;
  assign n13839 = pi65  & n13477;
  assign n13840 = pi66  & ~n13122;
  assign n13841 = ~n13839 & ~n13840;
  assign n13842 = pi69  & n12295;
  assign n13843 = pi67  & n12693;
  assign n13844 = pi68  & n12290;
  assign n13845 = ~n13843 & ~n13844;
  assign n13846 = ~n13842 & n13845;
  assign n13847 = n405 & n12298;
  assign n13848 = n13846 & ~n13847;
  assign n13849 = pi62  & ~n13848;
  assign n13850 = pi62  & ~n13849;
  assign n13851 = ~n13848 & ~n13849;
  assign n13852 = ~n13850 & ~n13851;
  assign n13853 = ~n13841 & ~n13852;
  assign n13854 = n13841 & n13852;
  assign n13855 = ~n13853 & ~n13854;
  assign n13856 = n13838 & ~n13855;
  assign n13857 = ~n13838 & n13855;
  assign n13858 = ~n13856 & ~n13857;
  assign n13859 = pi72  & n11193;
  assign n13860 = pi70  & n11567;
  assign n13861 = pi71  & n11188;
  assign n13862 = ~n13860 & ~n13861;
  assign n13863 = ~n13859 & n13862;
  assign n13864 = n575 & n11196;
  assign n13865 = n13863 & ~n13864;
  assign n13866 = pi59  & ~n13865;
  assign n13867 = pi59  & ~n13866;
  assign n13868 = ~n13865 & ~n13866;
  assign n13869 = ~n13867 & ~n13868;
  assign n13870 = n13858 & ~n13869;
  assign n13871 = ~n13858 & n13869;
  assign n13872 = ~n13837 & ~n13871;
  assign n13873 = ~n13870 & n13872;
  assign n13874 = ~n13837 & ~n13873;
  assign n13875 = ~n13870 & ~n13873;
  assign n13876 = ~n13871 & n13875;
  assign n13877 = ~n13874 & ~n13876;
  assign n13878 = pi75  & n10135;
  assign n13879 = pi73  & n10478;
  assign n13880 = pi74  & n10130;
  assign n13881 = ~n13879 & ~n13880;
  assign n13882 = ~n13878 & n13881;
  assign n13883 = n747 & n10138;
  assign n13884 = n13882 & ~n13883;
  assign n13885 = pi56  & ~n13884;
  assign n13886 = pi56  & ~n13885;
  assign n13887 = ~n13884 & ~n13885;
  assign n13888 = ~n13886 & ~n13887;
  assign n13889 = n13877 & n13888;
  assign n13890 = ~n13877 & ~n13888;
  assign n13891 = ~n13889 & ~n13890;
  assign n13892 = ~n13836 & n13891;
  assign n13893 = n13836 & ~n13891;
  assign n13894 = ~n13892 & ~n13893;
  assign n13895 = pi78  & n9096;
  assign n13896 = pi76  & n9453;
  assign n13897 = pi77  & n9091;
  assign n13898 = ~n13896 & ~n13897;
  assign n13899 = ~n13895 & n13898;
  assign n13900 = n1009 & n9099;
  assign n13901 = n13899 & ~n13900;
  assign n13902 = pi53  & ~n13901;
  assign n13903 = pi53  & ~n13902;
  assign n13904 = ~n13901 & ~n13902;
  assign n13905 = ~n13903 & ~n13904;
  assign n13906 = n13894 & ~n13905;
  assign n13907 = ~n13894 & n13905;
  assign n13908 = ~n13906 & ~n13907;
  assign n13909 = ~n13835 & n13908;
  assign n13910 = n13835 & ~n13908;
  assign n13911 = ~n13909 & ~n13910;
  assign n13912 = ~n13834 & n13911;
  assign n13913 = n13834 & ~n13911;
  assign n13914 = ~n13912 & ~n13913;
  assign n13915 = n13823 & ~n13914;
  assign n13916 = ~n13823 & n13914;
  assign n13917 = ~n13915 & ~n13916;
  assign n13918 = pi84  & n7239;
  assign n13919 = pi82  & n7556;
  assign n13920 = pi83  & n7234;
  assign n13921 = ~n13919 & ~n13920;
  assign n13922 = ~n13918 & n13921;
  assign n13923 = n1805 & n7242;
  assign n13924 = n13922 & ~n13923;
  assign n13925 = pi47  & ~n13924;
  assign n13926 = pi47  & ~n13925;
  assign n13927 = ~n13924 & ~n13925;
  assign n13928 = ~n13926 & ~n13927;
  assign n13929 = n13917 & ~n13928;
  assign n13930 = n13917 & ~n13929;
  assign n13931 = ~n13928 & ~n13929;
  assign n13932 = ~n13930 & ~n13931;
  assign n13933 = ~n13822 & ~n13932;
  assign n13934 = n13822 & n13932;
  assign n13935 = ~n13933 & ~n13934;
  assign n13936 = ~n13821 & n13935;
  assign n13937 = n13821 & ~n13935;
  assign n13938 = ~n13936 & ~n13937;
  assign n13939 = n13810 & ~n13938;
  assign n13940 = ~n13810 & n13938;
  assign n13941 = ~n13939 & ~n13940;
  assign n13942 = pi90  & n5636;
  assign n13943 = pi88  & n5909;
  assign n13944 = pi89  & n5631;
  assign n13945 = ~n13943 & ~n13944;
  assign n13946 = ~n13942 & n13945;
  assign n13947 = n2606 & n5639;
  assign n13948 = n13946 & ~n13947;
  assign n13949 = pi41  & ~n13948;
  assign n13950 = pi41  & ~n13949;
  assign n13951 = ~n13948 & ~n13949;
  assign n13952 = ~n13950 & ~n13951;
  assign n13953 = n13941 & ~n13952;
  assign n13954 = ~n13941 & n13952;
  assign n13955 = ~n13953 & ~n13954;
  assign n13956 = n13809 & ~n13955;
  assign n13957 = ~n13809 & n13955;
  assign n13958 = ~n13956 & ~n13957;
  assign n13959 = pi93  & n4896;
  assign n13960 = pi91  & n5148;
  assign n13961 = pi92  & n4891;
  assign n13962 = ~n13960 & ~n13961;
  assign n13963 = ~n13959 & n13962;
  assign n13964 = n3144 & n4899;
  assign n13965 = n13963 & ~n13964;
  assign n13966 = pi38  & ~n13965;
  assign n13967 = pi38  & ~n13966;
  assign n13968 = ~n13965 & ~n13966;
  assign n13969 = ~n13967 & ~n13968;
  assign n13970 = n13958 & ~n13969;
  assign n13971 = ~n13958 & n13969;
  assign n13972 = ~n13970 & ~n13971;
  assign n13973 = n13808 & ~n13972;
  assign n13974 = ~n13808 & n13972;
  assign n13975 = ~n13973 & ~n13974;
  assign n13976 = pi96  & n4182;
  assign n13977 = pi94  & n4416;
  assign n13978 = pi95  & n4177;
  assign n13979 = ~n13977 & ~n13978;
  assign n13980 = ~n13976 & n13979;
  assign n13981 = n3921 & n4185;
  assign n13982 = n13980 & ~n13981;
  assign n13983 = pi35  & ~n13982;
  assign n13984 = pi35  & ~n13983;
  assign n13985 = ~n13982 & ~n13983;
  assign n13986 = ~n13984 & ~n13985;
  assign n13987 = n13975 & ~n13986;
  assign n13988 = ~n13975 & n13986;
  assign n13989 = ~n13807 & ~n13988;
  assign n13990 = ~n13987 & n13989;
  assign n13991 = ~n13807 & ~n13990;
  assign n13992 = ~n13987 & ~n13990;
  assign n13993 = ~n13988 & n13992;
  assign n13994 = ~n13991 & ~n13993;
  assign n13995 = pi99  & n3550;
  assign n13996 = pi97  & n3735;
  assign n13997 = pi98  & n3545;
  assign n13998 = ~n13996 & ~n13997;
  assign n13999 = ~n13995 & n13998;
  assign n14000 = n3553 & n4584;
  assign n14001 = n13999 & ~n14000;
  assign n14002 = pi32  & ~n14001;
  assign n14003 = pi32  & ~n14002;
  assign n14004 = ~n14001 & ~n14002;
  assign n14005 = ~n14003 & ~n14004;
  assign n14006 = ~n13994 & ~n14005;
  assign n14007 = n13994 & n14005;
  assign n14008 = ~n14006 & ~n14007;
  assign n14009 = n13806 & ~n14008;
  assign n14010 = ~n13806 & n14008;
  assign n14011 = ~n14009 & ~n14010;
  assign n14012 = pi102  & n2976;
  assign n14013 = pi100  & n3182;
  assign n14014 = pi101  & n2971;
  assign n14015 = ~n14013 & ~n14014;
  assign n14016 = ~n14012 & n14015;
  assign n14017 = n2979 & n5296;
  assign n14018 = n14016 & ~n14017;
  assign n14019 = pi29  & ~n14018;
  assign n14020 = pi29  & ~n14019;
  assign n14021 = ~n14018 & ~n14019;
  assign n14022 = ~n14020 & ~n14021;
  assign n14023 = n14011 & ~n14022;
  assign n14024 = ~n14011 & n14022;
  assign n14025 = ~n14023 & ~n14024;
  assign n14026 = n13805 & ~n14025;
  assign n14027 = ~n13805 & n14025;
  assign n14028 = ~n14026 & ~n14027;
  assign n14029 = pi105  & n2486;
  assign n14030 = pi103  & n2644;
  assign n14031 = pi104  & n2481;
  assign n14032 = ~n14030 & ~n14031;
  assign n14033 = ~n14029 & n14032;
  assign n14034 = n2489 & n6065;
  assign n14035 = n14033 & ~n14034;
  assign n14036 = pi26  & ~n14035;
  assign n14037 = pi26  & ~n14036;
  assign n14038 = ~n14035 & ~n14036;
  assign n14039 = ~n14037 & ~n14038;
  assign n14040 = n14028 & ~n14039;
  assign n14041 = ~n14028 & n14039;
  assign n14042 = ~n13804 & ~n14041;
  assign n14043 = ~n14040 & n14042;
  assign n14044 = ~n13804 & ~n14043;
  assign n14045 = ~n14040 & ~n14043;
  assign n14046 = ~n14041 & n14045;
  assign n14047 = ~n14044 & ~n14046;
  assign n14048 = pi108  & n2004;
  assign n14049 = pi106  & n2141;
  assign n14050 = pi107  & n1999;
  assign n14051 = ~n14049 & ~n14050;
  assign n14052 = ~n14048 & n14051;
  assign n14053 = n2007 & n6639;
  assign n14054 = n14052 & ~n14053;
  assign n14055 = pi23  & ~n14054;
  assign n14056 = pi23  & ~n14055;
  assign n14057 = ~n14054 & ~n14055;
  assign n14058 = ~n14056 & ~n14057;
  assign n14059 = ~n14047 & ~n14058;
  assign n14060 = n14047 & n14058;
  assign n14061 = ~n14059 & ~n14060;
  assign n14062 = ~n13803 & n14061;
  assign n14063 = n13803 & ~n14061;
  assign n14064 = ~n14062 & ~n14063;
  assign n14065 = ~n13802 & n14064;
  assign n14066 = n13802 & ~n14064;
  assign n14067 = ~n14065 & ~n14066;
  assign n14068 = ~n13791 & n14067;
  assign n14069 = n13791 & ~n14067;
  assign n14070 = ~n14068 & ~n14069;
  assign n14071 = n13790 & ~n14070;
  assign n14072 = ~n13790 & n14070;
  assign n14073 = ~n14071 & ~n14072;
  assign n14074 = ~n13779 & n14073;
  assign n14075 = n13779 & ~n14073;
  assign n14076 = ~n14074 & ~n14075;
  assign n14077 = pi117  & n918;
  assign n14078 = pi115  & n1031;
  assign n14079 = pi116  & n913;
  assign n14080 = ~n14078 & ~n14079;
  assign n14081 = ~n14077 & n14080;
  assign n14082 = n921 & n9691;
  assign n14083 = n14081 & ~n14082;
  assign n14084 = pi14  & ~n14083;
  assign n14085 = pi14  & ~n14084;
  assign n14086 = ~n14083 & ~n14084;
  assign n14087 = ~n14085 & ~n14086;
  assign n14088 = n14076 & ~n14087;
  assign n14089 = ~n14076 & n14087;
  assign n14090 = ~n14088 & ~n14089;
  assign n14091 = n13778 & ~n14090;
  assign n14092 = ~n13778 & n14090;
  assign n14093 = ~n14091 & ~n14092;
  assign n14094 = pi120  & n675;
  assign n14095 = pi118  & n769;
  assign n14096 = pi119  & n670;
  assign n14097 = ~n14095 & ~n14096;
  assign n14098 = ~n14094 & n14097;
  assign n14099 = n678 & n10734;
  assign n14100 = n14098 & ~n14099;
  assign n14101 = pi11  & ~n14100;
  assign n14102 = pi11  & ~n14101;
  assign n14103 = ~n14100 & ~n14101;
  assign n14104 = ~n14102 & ~n14103;
  assign n14105 = ~n14093 & n14104;
  assign n14106 = n14093 & ~n14104;
  assign n14107 = ~n14105 & ~n14106;
  assign n14108 = pi123  & n493;
  assign n14109 = pi121  & n533;
  assign n14110 = pi122  & n488;
  assign n14111 = ~n14109 & ~n14110;
  assign n14112 = ~n14108 & n14111;
  assign n14113 = n496 & n11489;
  assign n14114 = n14112 & ~n14113;
  assign n14115 = pi8  & ~n14114;
  assign n14116 = pi8  & ~n14115;
  assign n14117 = ~n14114 & ~n14115;
  assign n14118 = ~n14116 & ~n14117;
  assign n14119 = n14107 & ~n14118;
  assign n14120 = ~n14107 & n14118;
  assign n14121 = ~n14119 & ~n14120;
  assign n14122 = n13777 & ~n14121;
  assign n14123 = ~n13777 & n14121;
  assign n14124 = ~n14122 & ~n14123;
  assign n14125 = pi126  & n340;
  assign n14126 = pi124  & n380;
  assign n14127 = pi125  & n335;
  assign n14128 = ~n14126 & ~n14127;
  assign n14129 = ~n14125 & n14128;
  assign n14130 = n343 & n12979;
  assign n14131 = n14129 & ~n14130;
  assign n14132 = pi5  & ~n14131;
  assign n14133 = pi5  & ~n14132;
  assign n14134 = ~n14131 & ~n14132;
  assign n14135 = ~n14133 & ~n14134;
  assign n14136 = n14124 & ~n14135;
  assign n14137 = ~n14124 & n14135;
  assign n14138 = ~n14136 & ~n14137;
  assign n14139 = n13776 & n14138;
  assign n14140 = ~n13776 & ~n14138;
  assign n14141 = ~n14139 & ~n14140;
  assign n14142 = n13766 & ~n14141;
  assign n14143 = ~n13766 & n14141;
  assign n14144 = ~n14142 & ~n14143;
  assign n14145 = ~n13760 & ~n13763;
  assign n14146 = n14144 & ~n14145;
  assign n14147 = ~n14144 & n14145;
  assign po65  = ~n14146 & ~n14147;
  assign n14149 = ~n13774 & ~n14139;
  assign n14150 = pi124  & n493;
  assign n14151 = pi122  & n533;
  assign n14152 = pi123  & n488;
  assign n14153 = ~n14151 & ~n14152;
  assign n14154 = ~n14150 & n14153;
  assign n14155 = n496 & n11858;
  assign n14156 = n14154 & ~n14155;
  assign n14157 = pi8  & ~n14156;
  assign n14158 = pi8  & ~n14157;
  assign n14159 = ~n14156 & ~n14157;
  assign n14160 = ~n14158 & ~n14159;
  assign n14161 = ~n14106 & ~n14119;
  assign n14162 = ~n14160 & ~n14161;
  assign n14163 = ~n14160 & ~n14162;
  assign n14164 = ~n14161 & ~n14162;
  assign n14165 = ~n14163 & ~n14164;
  assign n14166 = pi121  & n675;
  assign n14167 = pi119  & n769;
  assign n14168 = pi120  & n670;
  assign n14169 = ~n14167 & ~n14168;
  assign n14170 = ~n14166 & n14169;
  assign n14171 = n678 & n11086;
  assign n14172 = n14170 & ~n14171;
  assign n14173 = pi11  & ~n14172;
  assign n14174 = pi11  & ~n14173;
  assign n14175 = ~n14172 & ~n14173;
  assign n14176 = ~n14174 & ~n14175;
  assign n14177 = ~n14088 & ~n14092;
  assign n14178 = n14176 & n14177;
  assign n14179 = ~n14176 & ~n14177;
  assign n14180 = ~n14178 & ~n14179;
  assign n14181 = pi115  & n1269;
  assign n14182 = pi113  & n1340;
  assign n14183 = pi114  & n1264;
  assign n14184 = ~n14182 & ~n14183;
  assign n14185 = ~n14181 & n14184;
  assign n14186 = n1272 & n8727;
  assign n14187 = n14185 & ~n14186;
  assign n14188 = pi17  & ~n14187;
  assign n14189 = pi17  & ~n14188;
  assign n14190 = ~n14187 & ~n14188;
  assign n14191 = ~n14189 & ~n14190;
  assign n14192 = ~n14065 & ~n14068;
  assign n14193 = n14191 & n14192;
  assign n14194 = ~n14191 & ~n14192;
  assign n14195 = ~n14193 & ~n14194;
  assign n14196 = pi112  & n1582;
  assign n14197 = pi110  & n1713;
  assign n14198 = pi111  & n1577;
  assign n14199 = ~n14197 & ~n14198;
  assign n14200 = ~n14196 & n14199;
  assign n14201 = n1585 & n7795;
  assign n14202 = n14200 & ~n14201;
  assign n14203 = pi20  & ~n14202;
  assign n14204 = pi20  & ~n14203;
  assign n14205 = ~n14202 & ~n14203;
  assign n14206 = ~n14204 & ~n14205;
  assign n14207 = ~n14059 & ~n14062;
  assign n14208 = n14206 & n14207;
  assign n14209 = ~n14206 & ~n14207;
  assign n14210 = ~n14208 & ~n14209;
  assign n14211 = pi109  & n2004;
  assign n14212 = pi107  & n2141;
  assign n14213 = pi108  & n1999;
  assign n14214 = ~n14212 & ~n14213;
  assign n14215 = ~n14211 & n14214;
  assign n14216 = n2007 & n7170;
  assign n14217 = n14215 & ~n14216;
  assign n14218 = pi23  & ~n14217;
  assign n14219 = pi23  & ~n14218;
  assign n14220 = ~n14217 & ~n14218;
  assign n14221 = ~n14219 & ~n14220;
  assign n14222 = ~n14045 & n14221;
  assign n14223 = n14045 & ~n14221;
  assign n14224 = ~n14222 & ~n14223;
  assign n14225 = pi106  & n2486;
  assign n14226 = pi104  & n2644;
  assign n14227 = pi105  & n2481;
  assign n14228 = ~n14226 & ~n14227;
  assign n14229 = ~n14225 & n14228;
  assign n14230 = n2489 & n6090;
  assign n14231 = n14229 & ~n14230;
  assign n14232 = pi26  & ~n14231;
  assign n14233 = pi26  & ~n14232;
  assign n14234 = ~n14231 & ~n14232;
  assign n14235 = ~n14233 & ~n14234;
  assign n14236 = ~n14023 & ~n14027;
  assign n14237 = n14235 & n14236;
  assign n14238 = ~n14235 & ~n14236;
  assign n14239 = ~n14237 & ~n14238;
  assign n14240 = ~n14006 & ~n14010;
  assign n14241 = pi103  & n2976;
  assign n14242 = pi101  & n3182;
  assign n14243 = pi102  & n2971;
  assign n14244 = ~n14242 & ~n14243;
  assign n14245 = ~n14241 & n14244;
  assign n14246 = ~n2979 & n14245;
  assign n14247 = ~n5540 & n14245;
  assign n14248 = ~n14246 & ~n14247;
  assign n14249 = pi29  & ~n14248;
  assign n14250 = ~pi29  & n14248;
  assign n14251 = ~n14249 & ~n14250;
  assign n14252 = ~n14240 & ~n14251;
  assign n14253 = n14240 & n14251;
  assign n14254 = ~n14252 & ~n14253;
  assign n14255 = ~n13953 & ~n13957;
  assign n14256 = ~n13936 & ~n13940;
  assign n14257 = ~n13912 & ~n13916;
  assign n14258 = ~n13906 & ~n13909;
  assign n14259 = ~n13890 & ~n13892;
  assign n14260 = pi76  & n10135;
  assign n14261 = pi74  & n10478;
  assign n14262 = pi75  & n10130;
  assign n14263 = ~n14261 & ~n14262;
  assign n14264 = ~n14260 & n14263;
  assign n14265 = n881 & n10138;
  assign n14266 = n14264 & ~n14265;
  assign n14267 = pi56  & ~n14266;
  assign n14268 = pi56  & ~n14267;
  assign n14269 = ~n14266 & ~n14267;
  assign n14270 = ~n14268 & ~n14269;
  assign n14271 = ~n13853 & ~n13857;
  assign n14272 = pi66  & n13477;
  assign n14273 = pi67  & ~n13122;
  assign n14274 = ~n14272 & ~n14273;
  assign n14275 = pi2  & ~n14274;
  assign n14276 = ~pi2  & n14274;
  assign n14277 = ~n14275 & ~n14276;
  assign n14278 = pi70  & n12295;
  assign n14279 = pi68  & n12693;
  assign n14280 = pi69  & n12290;
  assign n14281 = ~n14279 & ~n14280;
  assign n14282 = ~n14278 & n14281;
  assign n14283 = ~n12298 & n14282;
  assign n14284 = ~n430 & n14282;
  assign n14285 = ~n14283 & ~n14284;
  assign n14286 = pi62  & ~n14285;
  assign n14287 = ~pi62  & n14285;
  assign n14288 = ~n14286 & ~n14287;
  assign n14289 = n14277 & ~n14288;
  assign n14290 = ~n14277 & n14288;
  assign n14291 = ~n14289 & ~n14290;
  assign n14292 = ~n14271 & n14291;
  assign n14293 = n14271 & ~n14291;
  assign n14294 = ~n14292 & ~n14293;
  assign n14295 = pi73  & n11193;
  assign n14296 = pi71  & n11567;
  assign n14297 = pi72  & n11188;
  assign n14298 = ~n14296 & ~n14297;
  assign n14299 = ~n14295 & n14298;
  assign n14300 = n639 & n11196;
  assign n14301 = n14299 & ~n14300;
  assign n14302 = pi59  & ~n14301;
  assign n14303 = pi59  & ~n14302;
  assign n14304 = ~n14301 & ~n14302;
  assign n14305 = ~n14303 & ~n14304;
  assign n14306 = n14294 & ~n14305;
  assign n14307 = ~n14294 & n14305;
  assign n14308 = ~n14306 & ~n14307;
  assign n14309 = ~n13875 & n14308;
  assign n14310 = n13875 & ~n14308;
  assign n14311 = ~n14309 & ~n14310;
  assign n14312 = n14270 & ~n14311;
  assign n14313 = ~n14270 & n14311;
  assign n14314 = ~n14312 & ~n14313;
  assign n14315 = ~n14259 & n14314;
  assign n14316 = n14259 & ~n14314;
  assign n14317 = ~n14315 & ~n14316;
  assign n14318 = pi79  & n9096;
  assign n14319 = pi77  & n9453;
  assign n14320 = pi78  & n9091;
  assign n14321 = ~n14319 & ~n14320;
  assign n14322 = ~n14318 & n14321;
  assign n14323 = n1105 & n9099;
  assign n14324 = n14322 & ~n14323;
  assign n14325 = pi53  & ~n14324;
  assign n14326 = pi53  & ~n14325;
  assign n14327 = ~n14324 & ~n14325;
  assign n14328 = ~n14326 & ~n14327;
  assign n14329 = n14317 & ~n14328;
  assign n14330 = ~n14317 & n14328;
  assign n14331 = ~n14329 & ~n14330;
  assign n14332 = n14258 & ~n14331;
  assign n14333 = ~n14258 & n14331;
  assign n14334 = ~n14332 & ~n14333;
  assign n14335 = pi82  & n8137;
  assign n14336 = pi80  & n8471;
  assign n14337 = pi81  & n8132;
  assign n14338 = ~n14336 & ~n14337;
  assign n14339 = ~n14335 & n14338;
  assign n14340 = n1532 & n8140;
  assign n14341 = n14339 & ~n14340;
  assign n14342 = pi50  & ~n14341;
  assign n14343 = pi50  & ~n14342;
  assign n14344 = ~n14341 & ~n14342;
  assign n14345 = ~n14343 & ~n14344;
  assign n14346 = n14334 & ~n14345;
  assign n14347 = ~n14334 & n14345;
  assign n14348 = ~n14346 & ~n14347;
  assign n14349 = n14257 & ~n14348;
  assign n14350 = ~n14257 & n14348;
  assign n14351 = ~n14349 & ~n14350;
  assign n14352 = pi85  & n7239;
  assign n14353 = pi83  & n7556;
  assign n14354 = pi84  & n7234;
  assign n14355 = ~n14353 & ~n14354;
  assign n14356 = ~n14352 & n14355;
  assign n14357 = n1943 & n7242;
  assign n14358 = n14356 & ~n14357;
  assign n14359 = pi47  & ~n14358;
  assign n14360 = pi47  & ~n14359;
  assign n14361 = ~n14358 & ~n14359;
  assign n14362 = ~n14360 & ~n14361;
  assign n14363 = ~n14351 & n14362;
  assign n14364 = n14351 & ~n14362;
  assign n14365 = ~n14363 & ~n14364;
  assign n14366 = ~n13929 & ~n13933;
  assign n14367 = n14365 & ~n14366;
  assign n14368 = ~n14365 & n14366;
  assign n14369 = ~n14367 & ~n14368;
  assign n14370 = pi88  & n6396;
  assign n14371 = pi86  & n6735;
  assign n14372 = pi87  & n6391;
  assign n14373 = ~n14371 & ~n14372;
  assign n14374 = ~n14370 & n14373;
  assign n14375 = n2277 & n6399;
  assign n14376 = n14374 & ~n14375;
  assign n14377 = pi44  & ~n14376;
  assign n14378 = pi44  & ~n14377;
  assign n14379 = ~n14376 & ~n14377;
  assign n14380 = ~n14378 & ~n14379;
  assign n14381 = n14369 & ~n14380;
  assign n14382 = ~n14369 & n14380;
  assign n14383 = ~n14381 & ~n14382;
  assign n14384 = n14256 & ~n14383;
  assign n14385 = ~n14256 & n14383;
  assign n14386 = ~n14384 & ~n14385;
  assign n14387 = pi91  & n5636;
  assign n14388 = pi89  & n5909;
  assign n14389 = pi90  & n5631;
  assign n14390 = ~n14388 & ~n14389;
  assign n14391 = ~n14387 & n14390;
  assign n14392 = n2926 & n5639;
  assign n14393 = n14391 & ~n14392;
  assign n14394 = pi41  & ~n14393;
  assign n14395 = pi41  & ~n14394;
  assign n14396 = ~n14393 & ~n14394;
  assign n14397 = ~n14395 & ~n14396;
  assign n14398 = n14386 & ~n14397;
  assign n14399 = ~n14386 & n14397;
  assign n14400 = ~n14398 & ~n14399;
  assign n14401 = n14255 & ~n14400;
  assign n14402 = ~n14255 & n14400;
  assign n14403 = ~n14401 & ~n14402;
  assign n14404 = pi94  & n4896;
  assign n14405 = pi92  & n5148;
  assign n14406 = pi93  & n4891;
  assign n14407 = ~n14405 & ~n14406;
  assign n14408 = ~n14404 & n14407;
  assign n14409 = n3499 & n4899;
  assign n14410 = n14408 & ~n14409;
  assign n14411 = pi38  & ~n14410;
  assign n14412 = pi38  & ~n14411;
  assign n14413 = ~n14410 & ~n14411;
  assign n14414 = ~n14412 & ~n14413;
  assign n14415 = ~n14403 & n14414;
  assign n14416 = n14403 & ~n14414;
  assign n14417 = ~n14415 & ~n14416;
  assign n14418 = ~n13970 & ~n13974;
  assign n14419 = n14417 & ~n14418;
  assign n14420 = ~n14417 & n14418;
  assign n14421 = ~n14419 & ~n14420;
  assign n14422 = pi97  & n4182;
  assign n14423 = pi95  & n4416;
  assign n14424 = pi96  & n4177;
  assign n14425 = ~n14423 & ~n14424;
  assign n14426 = ~n14422 & n14425;
  assign n14427 = n3946 & n4185;
  assign n14428 = n14426 & ~n14427;
  assign n14429 = pi35  & ~n14428;
  assign n14430 = pi35  & ~n14429;
  assign n14431 = ~n14428 & ~n14429;
  assign n14432 = ~n14430 & ~n14431;
  assign n14433 = n14421 & ~n14432;
  assign n14434 = ~n14421 & n14432;
  assign n14435 = ~n14433 & ~n14434;
  assign n14436 = pi100  & n3550;
  assign n14437 = pi98  & n3735;
  assign n14438 = pi99  & n3545;
  assign n14439 = ~n14437 & ~n14438;
  assign n14440 = ~n14436 & n14439;
  assign n14441 = ~n3553 & n14440;
  assign n14442 = ~n4808 & n14440;
  assign n14443 = ~n14441 & ~n14442;
  assign n14444 = pi32  & ~n14443;
  assign n14445 = ~pi32  & n14443;
  assign n14446 = ~n14444 & ~n14445;
  assign n14447 = ~n13992 & ~n14446;
  assign n14448 = n13992 & n14446;
  assign n14449 = ~n14447 & ~n14448;
  assign n14450 = n14435 & n14449;
  assign n14451 = ~n14435 & ~n14449;
  assign n14452 = ~n14450 & ~n14451;
  assign n14453 = n14254 & n14452;
  assign n14454 = ~n14254 & ~n14452;
  assign n14455 = ~n14453 & ~n14454;
  assign n14456 = n14239 & n14455;
  assign n14457 = ~n14239 & ~n14455;
  assign n14458 = ~n14224 & ~n14457;
  assign n14459 = ~n14456 & n14458;
  assign n14460 = ~n14224 & ~n14459;
  assign n14461 = ~n14457 & ~n14459;
  assign n14462 = ~n14456 & n14461;
  assign n14463 = ~n14460 & ~n14462;
  assign n14464 = n14210 & ~n14463;
  assign n14465 = ~n14210 & n14463;
  assign n14466 = n14195 & ~n14465;
  assign n14467 = ~n14464 & n14466;
  assign n14468 = n14195 & ~n14467;
  assign n14469 = ~n14465 & ~n14467;
  assign n14470 = ~n14464 & n14469;
  assign n14471 = ~n14468 & ~n14470;
  assign n14472 = ~n14072 & ~n14074;
  assign n14473 = pi118  & n918;
  assign n14474 = pi116  & n1031;
  assign n14475 = pi117  & n913;
  assign n14476 = ~n14474 & ~n14475;
  assign n14477 = ~n14473 & n14476;
  assign n14478 = ~n921 & n14477;
  assign n14479 = ~n9716 & n14477;
  assign n14480 = ~n14478 & ~n14479;
  assign n14481 = pi14  & ~n14480;
  assign n14482 = ~pi14  & n14480;
  assign n14483 = ~n14481 & ~n14482;
  assign n14484 = ~n14472 & ~n14483;
  assign n14485 = n14472 & n14483;
  assign n14486 = ~n14484 & ~n14485;
  assign n14487 = ~n14471 & n14486;
  assign n14488 = n14471 & ~n14486;
  assign n14489 = ~n14487 & ~n14488;
  assign n14490 = n14180 & n14489;
  assign n14491 = ~n14180 & ~n14489;
  assign n14492 = ~n14490 & ~n14491;
  assign n14493 = ~n14165 & n14492;
  assign n14494 = n14165 & ~n14492;
  assign n14495 = ~n14493 & ~n14494;
  assign n14496 = ~n14123 & ~n14136;
  assign n14497 = pi127  & n340;
  assign n14498 = pi125  & n380;
  assign n14499 = pi126  & n335;
  assign n14500 = ~n14498 & ~n14499;
  assign n14501 = ~n14497 & n14500;
  assign n14502 = n343 & n13365;
  assign n14503 = n14501 & ~n14502;
  assign n14504 = pi5  & ~n14503;
  assign n14505 = pi5  & ~n14504;
  assign n14506 = ~n14503 & ~n14504;
  assign n14507 = ~n14505 & ~n14506;
  assign n14508 = ~n14496 & ~n14507;
  assign n14509 = n14496 & n14507;
  assign n14510 = ~n14508 & ~n14509;
  assign n14511 = n14495 & n14510;
  assign n14512 = ~n14495 & ~n14510;
  assign n14513 = ~n14511 & ~n14512;
  assign n14514 = n14149 & ~n14513;
  assign n14515 = ~n14149 & n14513;
  assign n14516 = ~n14514 & ~n14515;
  assign n14517 = ~n14143 & ~n14146;
  assign n14518 = n14516 & ~n14517;
  assign n14519 = ~n14516 & n14517;
  assign po66  = ~n14518 & ~n14519;
  assign n14521 = ~n14515 & ~n14518;
  assign n14522 = ~n14508 & ~n14511;
  assign n14523 = ~n14484 & ~n14487;
  assign n14524 = pi122  & n675;
  assign n14525 = pi120  & n769;
  assign n14526 = pi121  & n670;
  assign n14527 = ~n14525 & ~n14526;
  assign n14528 = ~n14524 & n14527;
  assign n14529 = ~n678 & n14528;
  assign n14530 = ~n11463 & n14528;
  assign n14531 = ~n14529 & ~n14530;
  assign n14532 = pi11  & ~n14531;
  assign n14533 = ~pi11  & n14531;
  assign n14534 = ~n14532 & ~n14533;
  assign n14535 = ~n14523 & ~n14534;
  assign n14536 = n14523 & n14534;
  assign n14537 = ~n14535 & ~n14536;
  assign n14538 = pi119  & n918;
  assign n14539 = pi117  & n1031;
  assign n14540 = pi118  & n913;
  assign n14541 = ~n14539 & ~n14540;
  assign n14542 = ~n14538 & n14541;
  assign n14543 = n921 & n10048;
  assign n14544 = n14542 & ~n14543;
  assign n14545 = pi14  & ~n14544;
  assign n14546 = pi14  & ~n14545;
  assign n14547 = ~n14544 & ~n14545;
  assign n14548 = ~n14546 & ~n14547;
  assign n14549 = ~n14194 & ~n14467;
  assign n14550 = n14548 & n14549;
  assign n14551 = ~n14548 & ~n14549;
  assign n14552 = ~n14550 & ~n14551;
  assign n14553 = pi113  & n1582;
  assign n14554 = pi111  & n1713;
  assign n14555 = pi112  & n1577;
  assign n14556 = ~n14554 & ~n14555;
  assign n14557 = ~n14553 & n14556;
  assign n14558 = n1585 & n8387;
  assign n14559 = n14557 & ~n14558;
  assign n14560 = pi20  & ~n14559;
  assign n14561 = pi20  & ~n14560;
  assign n14562 = ~n14559 & ~n14560;
  assign n14563 = ~n14561 & ~n14562;
  assign n14564 = ~n14045 & ~n14221;
  assign n14565 = ~n14459 & ~n14564;
  assign n14566 = n14563 & n14565;
  assign n14567 = ~n14563 & ~n14565;
  assign n14568 = ~n14566 & ~n14567;
  assign n14569 = pi107  & n2486;
  assign n14570 = pi105  & n2644;
  assign n14571 = pi106  & n2481;
  assign n14572 = ~n14570 & ~n14571;
  assign n14573 = ~n14569 & n14572;
  assign n14574 = n2489 & n6614;
  assign n14575 = n14573 & ~n14574;
  assign n14576 = pi26  & ~n14575;
  assign n14577 = pi26  & ~n14576;
  assign n14578 = ~n14575 & ~n14576;
  assign n14579 = ~n14577 & ~n14578;
  assign n14580 = ~n14252 & ~n14453;
  assign n14581 = n14579 & n14580;
  assign n14582 = ~n14579 & ~n14580;
  assign n14583 = ~n14581 & ~n14582;
  assign n14584 = ~n14419 & ~n14433;
  assign n14585 = pi101  & n3550;
  assign n14586 = pi99  & n3735;
  assign n14587 = pi100  & n3545;
  assign n14588 = ~n14586 & ~n14587;
  assign n14589 = ~n14585 & n14588;
  assign n14590 = ~n3553 & n14589;
  assign n14591 = ~n5056 & n14589;
  assign n14592 = ~n14590 & ~n14591;
  assign n14593 = pi32  & ~n14592;
  assign n14594 = ~pi32  & n14592;
  assign n14595 = ~n14593 & ~n14594;
  assign n14596 = ~n14584 & ~n14595;
  assign n14597 = n14584 & n14595;
  assign n14598 = ~n14596 & ~n14597;
  assign n14599 = pi98  & n4182;
  assign n14600 = pi96  & n4416;
  assign n14601 = pi97  & n4177;
  assign n14602 = ~n14600 & ~n14601;
  assign n14603 = ~n14599 & n14602;
  assign n14604 = n4185 & n4360;
  assign n14605 = n14603 & ~n14604;
  assign n14606 = pi35  & ~n14605;
  assign n14607 = pi35  & ~n14606;
  assign n14608 = ~n14605 & ~n14606;
  assign n14609 = ~n14607 & ~n14608;
  assign n14610 = ~n14402 & ~n14416;
  assign n14611 = ~n14385 & ~n14398;
  assign n14612 = ~n14367 & ~n14381;
  assign n14613 = pi89  & n6396;
  assign n14614 = pi87  & n6735;
  assign n14615 = pi88  & n6391;
  assign n14616 = ~n14614 & ~n14615;
  assign n14617 = ~n14613 & n14616;
  assign n14618 = n2432 & n6399;
  assign n14619 = n14617 & ~n14618;
  assign n14620 = pi44  & ~n14619;
  assign n14621 = pi44  & ~n14620;
  assign n14622 = ~n14619 & ~n14620;
  assign n14623 = ~n14621 & ~n14622;
  assign n14624 = ~n14350 & ~n14364;
  assign n14625 = ~n14333 & ~n14346;
  assign n14626 = ~n14292 & ~n14306;
  assign n14627 = ~n14275 & ~n14289;
  assign n14628 = pi71  & n12295;
  assign n14629 = pi69  & n12693;
  assign n14630 = pi70  & n12290;
  assign n14631 = ~n14629 & ~n14630;
  assign n14632 = ~n14628 & n14631;
  assign n14633 = n476 & n12298;
  assign n14634 = n14632 & ~n14633;
  assign n14635 = pi62  & ~n14634;
  assign n14636 = pi62  & ~n14635;
  assign n14637 = ~n14634 & ~n14635;
  assign n14638 = ~n14636 & ~n14637;
  assign n14639 = pi67  & n13477;
  assign n14640 = pi68  & ~n13122;
  assign n14641 = ~n14639 & ~n14640;
  assign n14642 = pi2  & ~n14641;
  assign n14643 = ~pi2  & n14641;
  assign n14644 = ~n14642 & ~n14643;
  assign n14645 = ~n14638 & n14644;
  assign n14646 = n14638 & ~n14644;
  assign n14647 = ~n14645 & ~n14646;
  assign n14648 = n14627 & ~n14647;
  assign n14649 = ~n14627 & n14647;
  assign n14650 = ~n14648 & ~n14649;
  assign n14651 = pi74  & n11193;
  assign n14652 = pi72  & n11567;
  assign n14653 = pi73  & n11188;
  assign n14654 = ~n14652 & ~n14653;
  assign n14655 = ~n14651 & n14654;
  assign n14656 = n722 & n11196;
  assign n14657 = n14655 & ~n14656;
  assign n14658 = pi59  & ~n14657;
  assign n14659 = pi59  & ~n14658;
  assign n14660 = ~n14657 & ~n14658;
  assign n14661 = ~n14659 & ~n14660;
  assign n14662 = n14650 & ~n14661;
  assign n14663 = ~n14650 & n14661;
  assign n14664 = ~n14662 & ~n14663;
  assign n14665 = n14626 & ~n14664;
  assign n14666 = ~n14626 & n14664;
  assign n14667 = ~n14665 & ~n14666;
  assign n14668 = pi77  & n10135;
  assign n14669 = pi75  & n10478;
  assign n14670 = pi76  & n10130;
  assign n14671 = ~n14669 & ~n14670;
  assign n14672 = ~n14668 & n14671;
  assign n14673 = n984 & n10138;
  assign n14674 = n14672 & ~n14673;
  assign n14675 = pi56  & ~n14674;
  assign n14676 = pi56  & ~n14675;
  assign n14677 = ~n14674 & ~n14675;
  assign n14678 = ~n14676 & ~n14677;
  assign n14679 = ~n14667 & n14678;
  assign n14680 = n14667 & ~n14678;
  assign n14681 = ~n14679 & ~n14680;
  assign n14682 = ~n14309 & ~n14313;
  assign n14683 = n14681 & ~n14682;
  assign n14684 = ~n14681 & n14682;
  assign n14685 = ~n14683 & ~n14684;
  assign n14686 = pi80  & n9096;
  assign n14687 = pi78  & n9453;
  assign n14688 = pi79  & n9091;
  assign n14689 = ~n14687 & ~n14688;
  assign n14690 = ~n14686 & n14689;
  assign n14691 = n1205 & n9099;
  assign n14692 = n14690 & ~n14691;
  assign n14693 = pi53  & ~n14692;
  assign n14694 = pi53  & ~n14693;
  assign n14695 = ~n14692 & ~n14693;
  assign n14696 = ~n14694 & ~n14695;
  assign n14697 = n14685 & ~n14696;
  assign n14698 = n14685 & ~n14697;
  assign n14699 = ~n14696 & ~n14697;
  assign n14700 = ~n14698 & ~n14699;
  assign n14701 = ~n14315 & ~n14329;
  assign n14702 = n14700 & n14701;
  assign n14703 = ~n14700 & ~n14701;
  assign n14704 = ~n14702 & ~n14703;
  assign n14705 = pi83  & n8137;
  assign n14706 = pi81  & n8471;
  assign n14707 = pi82  & n8132;
  assign n14708 = ~n14706 & ~n14707;
  assign n14709 = ~n14705 & n14708;
  assign n14710 = n1672 & n8140;
  assign n14711 = n14709 & ~n14710;
  assign n14712 = pi50  & ~n14711;
  assign n14713 = pi50  & ~n14712;
  assign n14714 = ~n14711 & ~n14712;
  assign n14715 = ~n14713 & ~n14714;
  assign n14716 = n14704 & ~n14715;
  assign n14717 = ~n14704 & n14715;
  assign n14718 = ~n14716 & ~n14717;
  assign n14719 = n14625 & ~n14718;
  assign n14720 = ~n14625 & n14718;
  assign n14721 = ~n14719 & ~n14720;
  assign n14722 = pi86  & n7239;
  assign n14723 = pi84  & n7556;
  assign n14724 = pi85  & n7234;
  assign n14725 = ~n14723 & ~n14724;
  assign n14726 = ~n14722 & n14725;
  assign n14727 = n2099 & n7242;
  assign n14728 = n14726 & ~n14727;
  assign n14729 = pi47  & ~n14728;
  assign n14730 = pi47  & ~n14729;
  assign n14731 = ~n14728 & ~n14729;
  assign n14732 = ~n14730 & ~n14731;
  assign n14733 = n14721 & ~n14732;
  assign n14734 = ~n14721 & n14732;
  assign n14735 = ~n14733 & ~n14734;
  assign n14736 = ~n14624 & n14735;
  assign n14737 = n14624 & ~n14735;
  assign n14738 = ~n14736 & ~n14737;
  assign n14739 = ~n14623 & n14738;
  assign n14740 = n14623 & ~n14738;
  assign n14741 = ~n14739 & ~n14740;
  assign n14742 = n14612 & ~n14741;
  assign n14743 = ~n14612 & n14741;
  assign n14744 = ~n14742 & ~n14743;
  assign n14745 = pi92  & n5636;
  assign n14746 = pi90  & n5909;
  assign n14747 = pi91  & n5631;
  assign n14748 = ~n14746 & ~n14747;
  assign n14749 = ~n14745 & n14748;
  assign n14750 = n3119 & n5639;
  assign n14751 = n14749 & ~n14750;
  assign n14752 = pi41  & ~n14751;
  assign n14753 = pi41  & ~n14752;
  assign n14754 = ~n14751 & ~n14752;
  assign n14755 = ~n14753 & ~n14754;
  assign n14756 = n14744 & ~n14755;
  assign n14757 = ~n14744 & n14755;
  assign n14758 = ~n14756 & ~n14757;
  assign n14759 = n14611 & ~n14758;
  assign n14760 = ~n14611 & n14758;
  assign n14761 = ~n14759 & ~n14760;
  assign n14762 = pi95  & n4896;
  assign n14763 = pi93  & n5148;
  assign n14764 = pi94  & n4891;
  assign n14765 = ~n14763 & ~n14764;
  assign n14766 = ~n14762 & n14765;
  assign n14767 = n3710 & n4899;
  assign n14768 = n14766 & ~n14767;
  assign n14769 = pi38  & ~n14768;
  assign n14770 = pi38  & ~n14769;
  assign n14771 = ~n14768 & ~n14769;
  assign n14772 = ~n14770 & ~n14771;
  assign n14773 = ~n14761 & n14772;
  assign n14774 = n14761 & ~n14772;
  assign n14775 = ~n14773 & ~n14774;
  assign n14776 = ~n14610 & n14775;
  assign n14777 = n14610 & ~n14775;
  assign n14778 = ~n14776 & ~n14777;
  assign n14779 = ~n14609 & n14778;
  assign n14780 = n14609 & ~n14778;
  assign n14781 = ~n14779 & ~n14780;
  assign n14782 = ~n14598 & ~n14781;
  assign n14783 = n14598 & n14781;
  assign n14784 = ~n14782 & ~n14783;
  assign n14785 = ~n14447 & ~n14450;
  assign n14786 = pi104  & n2976;
  assign n14787 = pi102  & n3182;
  assign n14788 = pi103  & n2971;
  assign n14789 = ~n14787 & ~n14788;
  assign n14790 = ~n14786 & n14789;
  assign n14791 = ~n2979 & n14790;
  assign n14792 = ~n5565 & n14790;
  assign n14793 = ~n14791 & ~n14792;
  assign n14794 = pi29  & ~n14793;
  assign n14795 = ~pi29  & n14793;
  assign n14796 = ~n14794 & ~n14795;
  assign n14797 = ~n14785 & ~n14796;
  assign n14798 = n14785 & n14796;
  assign n14799 = ~n14797 & ~n14798;
  assign n14800 = n14784 & n14799;
  assign n14801 = ~n14784 & ~n14799;
  assign n14802 = ~n14800 & ~n14801;
  assign n14803 = n14583 & n14802;
  assign n14804 = ~n14583 & ~n14802;
  assign n14805 = ~n14803 & ~n14804;
  assign n14806 = pi110  & n2004;
  assign n14807 = pi108  & n2141;
  assign n14808 = pi109  & n1999;
  assign n14809 = ~n14807 & ~n14808;
  assign n14810 = ~n14806 & n14809;
  assign n14811 = n2007 & n7474;
  assign n14812 = n14810 & ~n14811;
  assign n14813 = pi23  & ~n14812;
  assign n14814 = pi23  & ~n14813;
  assign n14815 = ~n14812 & ~n14813;
  assign n14816 = ~n14814 & ~n14815;
  assign n14817 = ~n14238 & ~n14456;
  assign n14818 = ~n14816 & ~n14817;
  assign n14819 = n14816 & n14817;
  assign n14820 = ~n14818 & ~n14819;
  assign n14821 = n14805 & n14820;
  assign n14822 = ~n14805 & ~n14820;
  assign n14823 = ~n14821 & ~n14822;
  assign n14824 = n14568 & n14823;
  assign n14825 = ~n14568 & ~n14823;
  assign n14826 = ~n14824 & ~n14825;
  assign n14827 = pi116  & n1269;
  assign n14828 = pi114  & n1340;
  assign n14829 = pi115  & n1264;
  assign n14830 = ~n14828 & ~n14829;
  assign n14831 = ~n14827 & n14830;
  assign n14832 = n1272 & n9042;
  assign n14833 = n14831 & ~n14832;
  assign n14834 = pi17  & ~n14833;
  assign n14835 = pi17  & ~n14834;
  assign n14836 = ~n14833 & ~n14834;
  assign n14837 = ~n14835 & ~n14836;
  assign n14838 = ~n14209 & ~n14464;
  assign n14839 = ~n14837 & ~n14838;
  assign n14840 = n14837 & n14838;
  assign n14841 = ~n14839 & ~n14840;
  assign n14842 = n14826 & n14841;
  assign n14843 = ~n14826 & ~n14841;
  assign n14844 = ~n14842 & ~n14843;
  assign n14845 = n14552 & n14844;
  assign n14846 = ~n14552 & ~n14844;
  assign n14847 = ~n14845 & ~n14846;
  assign n14848 = n14537 & n14847;
  assign n14849 = ~n14537 & ~n14847;
  assign n14850 = ~n14848 & ~n14849;
  assign n14851 = ~n14179 & ~n14490;
  assign n14852 = pi125  & n493;
  assign n14853 = pi123  & n533;
  assign n14854 = pi124  & n488;
  assign n14855 = ~n14853 & ~n14854;
  assign n14856 = ~n14852 & n14855;
  assign n14857 = ~n496 & n14856;
  assign n14858 = ~n12591 & n14856;
  assign n14859 = ~n14857 & ~n14858;
  assign n14860 = pi8  & ~n14859;
  assign n14861 = ~pi8  & n14859;
  assign n14862 = ~n14860 & ~n14861;
  assign n14863 = ~n14851 & ~n14862;
  assign n14864 = n14851 & n14862;
  assign n14865 = ~n14863 & ~n14864;
  assign n14866 = n14850 & n14865;
  assign n14867 = ~n14850 & ~n14865;
  assign n14868 = ~n14866 & ~n14867;
  assign n14869 = ~n14162 & ~n14493;
  assign n14870 = pi126  & n380;
  assign n14871 = pi127  & n335;
  assign n14872 = ~n14870 & ~n14871;
  assign n14873 = ~n343 & n14872;
  assign n14874 = ~n13389 & n14872;
  assign n14875 = ~n14873 & ~n14874;
  assign n14876 = pi5  & ~n14875;
  assign n14877 = ~pi5  & n14875;
  assign n14878 = ~n14876 & ~n14877;
  assign n14879 = ~n14869 & ~n14878;
  assign n14880 = n14869 & n14878;
  assign n14881 = ~n14879 & ~n14880;
  assign n14882 = n14868 & n14881;
  assign n14883 = ~n14868 & ~n14881;
  assign n14884 = ~n14882 & ~n14883;
  assign n14885 = ~n14522 & n14884;
  assign n14886 = n14522 & ~n14884;
  assign n14887 = ~n14885 & ~n14886;
  assign n14888 = ~n14521 & n14887;
  assign n14889 = n14521 & ~n14887;
  assign po67  = ~n14888 & ~n14889;
  assign n14891 = ~n14885 & ~n14888;
  assign n14892 = ~n14879 & ~n14882;
  assign n14893 = pi123  & n675;
  assign n14894 = pi121  & n769;
  assign n14895 = pi122  & n670;
  assign n14896 = ~n14894 & ~n14895;
  assign n14897 = ~n14893 & n14896;
  assign n14898 = n678 & n11489;
  assign n14899 = n14897 & ~n14898;
  assign n14900 = pi11  & ~n14899;
  assign n14901 = pi11  & ~n14900;
  assign n14902 = ~n14899 & ~n14900;
  assign n14903 = ~n14901 & ~n14902;
  assign n14904 = ~n14551 & ~n14845;
  assign n14905 = n14903 & n14904;
  assign n14906 = ~n14903 & ~n14904;
  assign n14907 = ~n14905 & ~n14906;
  assign n14908 = ~n14567 & ~n14824;
  assign n14909 = pi117  & n1269;
  assign n14910 = pi115  & n1340;
  assign n14911 = pi116  & n1264;
  assign n14912 = ~n14910 & ~n14911;
  assign n14913 = ~n14909 & n14912;
  assign n14914 = ~n1272 & n14913;
  assign n14915 = ~n9691 & n14913;
  assign n14916 = ~n14914 & ~n14915;
  assign n14917 = pi17  & ~n14916;
  assign n14918 = ~pi17  & n14916;
  assign n14919 = ~n14917 & ~n14918;
  assign n14920 = ~n14908 & ~n14919;
  assign n14921 = n14908 & n14919;
  assign n14922 = ~n14920 & ~n14921;
  assign n14923 = pi114  & n1582;
  assign n14924 = pi112  & n1713;
  assign n14925 = pi113  & n1577;
  assign n14926 = ~n14924 & ~n14925;
  assign n14927 = ~n14923 & n14926;
  assign n14928 = n1585 & n8702;
  assign n14929 = n14927 & ~n14928;
  assign n14930 = pi20  & ~n14929;
  assign n14931 = pi20  & ~n14930;
  assign n14932 = ~n14929 & ~n14930;
  assign n14933 = ~n14931 & ~n14932;
  assign n14934 = ~n14818 & ~n14821;
  assign n14935 = ~n14933 & ~n14934;
  assign n14936 = n14933 & n14934;
  assign n14937 = ~n14935 & ~n14936;
  assign n14938 = pi111  & n2004;
  assign n14939 = pi109  & n2141;
  assign n14940 = pi110  & n1999;
  assign n14941 = ~n14939 & ~n14940;
  assign n14942 = ~n14938 & n14941;
  assign n14943 = n2007 & n7770;
  assign n14944 = n14942 & ~n14943;
  assign n14945 = pi23  & ~n14944;
  assign n14946 = pi23  & ~n14945;
  assign n14947 = ~n14944 & ~n14945;
  assign n14948 = ~n14946 & ~n14947;
  assign n14949 = ~n14582 & ~n14803;
  assign n14950 = n14948 & n14949;
  assign n14951 = ~n14948 & ~n14949;
  assign n14952 = ~n14950 & ~n14951;
  assign n14953 = pi105  & n2976;
  assign n14954 = pi103  & n3182;
  assign n14955 = pi104  & n2971;
  assign n14956 = ~n14954 & ~n14955;
  assign n14957 = ~n14953 & n14956;
  assign n14958 = n2979 & n6065;
  assign n14959 = n14957 & ~n14958;
  assign n14960 = pi29  & ~n14959;
  assign n14961 = pi29  & ~n14960;
  assign n14962 = ~n14959 & ~n14960;
  assign n14963 = ~n14961 & ~n14962;
  assign n14964 = ~n14596 & ~n14783;
  assign n14965 = n14963 & n14964;
  assign n14966 = ~n14963 & ~n14964;
  assign n14967 = ~n14965 & ~n14966;
  assign n14968 = ~n14776 & ~n14779;
  assign n14969 = pi102  & n3550;
  assign n14970 = pi100  & n3735;
  assign n14971 = pi101  & n3545;
  assign n14972 = ~n14970 & ~n14971;
  assign n14973 = ~n14969 & n14972;
  assign n14974 = ~n3553 & n14973;
  assign n14975 = ~n5296 & n14973;
  assign n14976 = ~n14974 & ~n14975;
  assign n14977 = pi32  & ~n14976;
  assign n14978 = ~pi32  & n14976;
  assign n14979 = ~n14977 & ~n14978;
  assign n14980 = ~n14968 & ~n14979;
  assign n14981 = n14968 & n14979;
  assign n14982 = ~n14980 & ~n14981;
  assign n14983 = ~n14743 & ~n14756;
  assign n14984 = ~n14736 & ~n14739;
  assign n14985 = ~n14720 & ~n14733;
  assign n14986 = ~n14683 & ~n14697;
  assign n14987 = ~n14642 & ~n14645;
  assign n14988 = pi72  & n12295;
  assign n14989 = pi70  & n12693;
  assign n14990 = pi71  & n12290;
  assign n14991 = ~n14989 & ~n14990;
  assign n14992 = ~n14988 & n14991;
  assign n14993 = n575 & n12298;
  assign n14994 = n14992 & ~n14993;
  assign n14995 = pi62  & ~n14994;
  assign n14996 = pi62  & ~n14995;
  assign n14997 = ~n14994 & ~n14995;
  assign n14998 = ~n14996 & ~n14997;
  assign n14999 = pi68  & n13477;
  assign n15000 = pi69  & ~n13122;
  assign n15001 = ~n14999 & ~n15000;
  assign n15002 = pi2  & ~n15001;
  assign n15003 = ~pi2  & n15001;
  assign n15004 = ~n15002 & ~n15003;
  assign n15005 = ~n14998 & n15004;
  assign n15006 = n14998 & ~n15004;
  assign n15007 = ~n15005 & ~n15006;
  assign n15008 = n14987 & ~n15007;
  assign n15009 = ~n14987 & n15007;
  assign n15010 = ~n15008 & ~n15009;
  assign n15011 = pi75  & n11193;
  assign n15012 = pi73  & n11567;
  assign n15013 = pi74  & n11188;
  assign n15014 = ~n15012 & ~n15013;
  assign n15015 = ~n15011 & n15014;
  assign n15016 = n747 & n11196;
  assign n15017 = n15015 & ~n15016;
  assign n15018 = pi59  & ~n15017;
  assign n15019 = pi59  & ~n15018;
  assign n15020 = ~n15017 & ~n15018;
  assign n15021 = ~n15019 & ~n15020;
  assign n15022 = ~n15010 & n15021;
  assign n15023 = n15010 & ~n15021;
  assign n15024 = ~n15022 & ~n15023;
  assign n15025 = ~n14649 & ~n14662;
  assign n15026 = n15024 & ~n15025;
  assign n15027 = ~n15024 & n15025;
  assign n15028 = ~n15026 & ~n15027;
  assign n15029 = pi78  & n10135;
  assign n15030 = pi76  & n10478;
  assign n15031 = pi77  & n10130;
  assign n15032 = ~n15030 & ~n15031;
  assign n15033 = ~n15029 & n15032;
  assign n15034 = n1009 & n10138;
  assign n15035 = n15033 & ~n15034;
  assign n15036 = pi56  & ~n15035;
  assign n15037 = pi56  & ~n15036;
  assign n15038 = ~n15035 & ~n15036;
  assign n15039 = ~n15037 & ~n15038;
  assign n15040 = n15028 & ~n15039;
  assign n15041 = n15028 & ~n15040;
  assign n15042 = ~n15039 & ~n15040;
  assign n15043 = ~n15041 & ~n15042;
  assign n15044 = ~n14666 & ~n14680;
  assign n15045 = ~n15043 & ~n15044;
  assign n15046 = n15043 & n15044;
  assign n15047 = ~n15045 & ~n15046;
  assign n15048 = pi81  & n9096;
  assign n15049 = pi79  & n9453;
  assign n15050 = pi80  & n9091;
  assign n15051 = ~n15049 & ~n15050;
  assign n15052 = ~n15048 & n15051;
  assign n15053 = n1413 & n9099;
  assign n15054 = n15052 & ~n15053;
  assign n15055 = pi53  & ~n15054;
  assign n15056 = pi53  & ~n15055;
  assign n15057 = ~n15054 & ~n15055;
  assign n15058 = ~n15056 & ~n15057;
  assign n15059 = n15047 & ~n15058;
  assign n15060 = ~n15047 & n15058;
  assign n15061 = ~n15059 & ~n15060;
  assign n15062 = n14986 & ~n15061;
  assign n15063 = ~n14986 & n15061;
  assign n15064 = ~n15062 & ~n15063;
  assign n15065 = pi84  & n8137;
  assign n15066 = pi82  & n8471;
  assign n15067 = pi83  & n8132;
  assign n15068 = ~n15066 & ~n15067;
  assign n15069 = ~n15065 & n15068;
  assign n15070 = n1805 & n8140;
  assign n15071 = n15069 & ~n15070;
  assign n15072 = pi50  & ~n15071;
  assign n15073 = pi50  & ~n15072;
  assign n15074 = ~n15071 & ~n15072;
  assign n15075 = ~n15073 & ~n15074;
  assign n15076 = ~n15064 & n15075;
  assign n15077 = n15064 & ~n15075;
  assign n15078 = ~n15076 & ~n15077;
  assign n15079 = ~n14703 & ~n14716;
  assign n15080 = n15078 & ~n15079;
  assign n15081 = ~n15078 & n15079;
  assign n15082 = ~n15080 & ~n15081;
  assign n15083 = pi87  & n7239;
  assign n15084 = pi85  & n7556;
  assign n15085 = pi86  & n7234;
  assign n15086 = ~n15084 & ~n15085;
  assign n15087 = ~n15083 & n15086;
  assign n15088 = n2252 & n7242;
  assign n15089 = n15087 & ~n15088;
  assign n15090 = pi47  & ~n15089;
  assign n15091 = pi47  & ~n15090;
  assign n15092 = ~n15089 & ~n15090;
  assign n15093 = ~n15091 & ~n15092;
  assign n15094 = n15082 & ~n15093;
  assign n15095 = ~n15082 & n15093;
  assign n15096 = ~n15094 & ~n15095;
  assign n15097 = n14985 & ~n15096;
  assign n15098 = ~n14985 & n15096;
  assign n15099 = ~n15097 & ~n15098;
  assign n15100 = pi90  & n6396;
  assign n15101 = pi88  & n6735;
  assign n15102 = pi89  & n6391;
  assign n15103 = ~n15101 & ~n15102;
  assign n15104 = ~n15100 & n15103;
  assign n15105 = n2606 & n6399;
  assign n15106 = n15104 & ~n15105;
  assign n15107 = pi44  & ~n15106;
  assign n15108 = pi44  & ~n15107;
  assign n15109 = ~n15106 & ~n15107;
  assign n15110 = ~n15108 & ~n15109;
  assign n15111 = n15099 & ~n15110;
  assign n15112 = ~n15099 & n15110;
  assign n15113 = ~n15111 & ~n15112;
  assign n15114 = n14984 & ~n15113;
  assign n15115 = ~n14984 & n15113;
  assign n15116 = ~n15114 & ~n15115;
  assign n15117 = pi93  & n5636;
  assign n15118 = pi91  & n5909;
  assign n15119 = pi92  & n5631;
  assign n15120 = ~n15118 & ~n15119;
  assign n15121 = ~n15117 & n15120;
  assign n15122 = n3144 & n5639;
  assign n15123 = n15121 & ~n15122;
  assign n15124 = pi41  & ~n15123;
  assign n15125 = pi41  & ~n15124;
  assign n15126 = ~n15123 & ~n15124;
  assign n15127 = ~n15125 & ~n15126;
  assign n15128 = n15116 & ~n15127;
  assign n15129 = ~n15116 & n15127;
  assign n15130 = ~n15128 & ~n15129;
  assign n15131 = n14983 & ~n15130;
  assign n15132 = ~n14983 & n15130;
  assign n15133 = ~n15131 & ~n15132;
  assign n15134 = pi96  & n4896;
  assign n15135 = pi94  & n5148;
  assign n15136 = pi95  & n4891;
  assign n15137 = ~n15135 & ~n15136;
  assign n15138 = ~n15134 & n15137;
  assign n15139 = n3921 & n4899;
  assign n15140 = n15138 & ~n15139;
  assign n15141 = pi38  & ~n15140;
  assign n15142 = pi38  & ~n15141;
  assign n15143 = ~n15140 & ~n15141;
  assign n15144 = ~n15142 & ~n15143;
  assign n15145 = ~n15133 & n15144;
  assign n15146 = n15133 & ~n15144;
  assign n15147 = ~n15145 & ~n15146;
  assign n15148 = ~n14760 & ~n14774;
  assign n15149 = n15147 & ~n15148;
  assign n15150 = ~n15147 & n15148;
  assign n15151 = ~n15149 & ~n15150;
  assign n15152 = pi99  & n4182;
  assign n15153 = pi97  & n4416;
  assign n15154 = pi98  & n4177;
  assign n15155 = ~n15153 & ~n15154;
  assign n15156 = ~n15152 & n15155;
  assign n15157 = n4185 & n4584;
  assign n15158 = n15156 & ~n15157;
  assign n15159 = pi35  & ~n15158;
  assign n15160 = pi35  & ~n15159;
  assign n15161 = ~n15158 & ~n15159;
  assign n15162 = ~n15160 & ~n15161;
  assign n15163 = n15151 & ~n15162;
  assign n15164 = ~n15151 & n15162;
  assign n15165 = ~n15163 & ~n15164;
  assign n15166 = n14982 & n15165;
  assign n15167 = ~n14982 & ~n15165;
  assign n15168 = ~n15166 & ~n15167;
  assign n15169 = n14967 & n15168;
  assign n15170 = ~n14967 & ~n15168;
  assign n15171 = ~n15169 & ~n15170;
  assign n15172 = ~n14797 & ~n14800;
  assign n15173 = pi108  & n2486;
  assign n15174 = pi106  & n2644;
  assign n15175 = pi107  & n2481;
  assign n15176 = ~n15174 & ~n15175;
  assign n15177 = ~n15173 & n15176;
  assign n15178 = ~n2489 & n15177;
  assign n15179 = ~n6639 & n15177;
  assign n15180 = ~n15178 & ~n15179;
  assign n15181 = pi26  & ~n15180;
  assign n15182 = ~pi26  & n15180;
  assign n15183 = ~n15181 & ~n15182;
  assign n15184 = ~n15172 & ~n15183;
  assign n15185 = n15172 & n15183;
  assign n15186 = ~n15184 & ~n15185;
  assign n15187 = n15171 & n15186;
  assign n15188 = ~n15171 & ~n15186;
  assign n15189 = ~n15187 & ~n15188;
  assign n15190 = n14952 & n15189;
  assign n15191 = ~n14952 & ~n15189;
  assign n15192 = ~n15190 & ~n15191;
  assign n15193 = n14937 & ~n15192;
  assign n15194 = ~n14937 & n15192;
  assign n15195 = ~n15193 & ~n15194;
  assign n15196 = n14922 & ~n15195;
  assign n15197 = ~n14922 & n15195;
  assign n15198 = ~n15196 & ~n15197;
  assign n15199 = pi120  & n918;
  assign n15200 = pi118  & n1031;
  assign n15201 = pi119  & n913;
  assign n15202 = ~n15200 & ~n15201;
  assign n15203 = ~n15199 & n15202;
  assign n15204 = n921 & n10734;
  assign n15205 = n15203 & ~n15204;
  assign n15206 = pi14  & ~n15205;
  assign n15207 = pi14  & ~n15206;
  assign n15208 = ~n15205 & ~n15206;
  assign n15209 = ~n15207 & ~n15208;
  assign n15210 = ~n14839 & ~n14842;
  assign n15211 = ~n15209 & ~n15210;
  assign n15212 = n15209 & n15210;
  assign n15213 = ~n15211 & ~n15212;
  assign n15214 = n15198 & n15213;
  assign n15215 = ~n15198 & ~n15213;
  assign n15216 = ~n15214 & ~n15215;
  assign n15217 = n14907 & n15216;
  assign n15218 = ~n14907 & ~n15216;
  assign n15219 = ~n15217 & ~n15218;
  assign n15220 = ~n14535 & ~n14848;
  assign n15221 = pi126  & n493;
  assign n15222 = pi124  & n533;
  assign n15223 = pi125  & n488;
  assign n15224 = ~n15222 & ~n15223;
  assign n15225 = ~n15221 & n15224;
  assign n15226 = ~n496 & n15225;
  assign n15227 = ~n12979 & n15225;
  assign n15228 = ~n15226 & ~n15227;
  assign n15229 = pi8  & ~n15228;
  assign n15230 = ~pi8  & n15228;
  assign n15231 = ~n15229 & ~n15230;
  assign n15232 = ~n15220 & ~n15231;
  assign n15233 = n15220 & n15231;
  assign n15234 = ~n15232 & ~n15233;
  assign n15235 = n15219 & n15234;
  assign n15236 = ~n15219 & ~n15234;
  assign n15237 = ~n15235 & ~n15236;
  assign n15238 = ~n14863 & ~n14866;
  assign n15239 = pi127  & n380;
  assign n15240 = n343 & n13387;
  assign n15241 = ~n15239 & ~n15240;
  assign n15242 = pi5  & ~n15241;
  assign n15243 = pi5  & ~n15242;
  assign n15244 = ~n15241 & ~n15242;
  assign n15245 = ~n15243 & ~n15244;
  assign n15246 = ~n15238 & ~n15245;
  assign n15247 = n15238 & n15245;
  assign n15248 = ~n15246 & ~n15247;
  assign n15249 = n15237 & n15248;
  assign n15250 = ~n15237 & ~n15248;
  assign n15251 = ~n15249 & ~n15250;
  assign n15252 = ~n14892 & n15251;
  assign n15253 = n14892 & ~n15251;
  assign n15254 = ~n15252 & ~n15253;
  assign n15255 = ~n14891 & n15254;
  assign n15256 = n14891 & ~n15254;
  assign po68  = ~n15255 & ~n15256;
  assign n15258 = ~n15252 & ~n15255;
  assign n15259 = ~n15246 & ~n15249;
  assign n15260 = ~n15232 & ~n15235;
  assign n15261 = pi127  & n493;
  assign n15262 = pi125  & n533;
  assign n15263 = pi126  & n488;
  assign n15264 = ~n15262 & ~n15263;
  assign n15265 = ~n15261 & n15264;
  assign n15266 = n496 & n13365;
  assign n15267 = n15265 & ~n15266;
  assign n15268 = pi8  & ~n15267;
  assign n15269 = pi8  & ~n15268;
  assign n15270 = ~n15267 & ~n15268;
  assign n15271 = ~n15269 & ~n15270;
  assign n15272 = ~n15260 & ~n15271;
  assign n15273 = n15260 & n15271;
  assign n15274 = ~n15272 & ~n15273;
  assign n15275 = pi124  & n675;
  assign n15276 = pi122  & n769;
  assign n15277 = pi123  & n670;
  assign n15278 = ~n15276 & ~n15277;
  assign n15279 = ~n15275 & n15278;
  assign n15280 = n678 & n11858;
  assign n15281 = n15279 & ~n15280;
  assign n15282 = pi11  & ~n15281;
  assign n15283 = pi11  & ~n15282;
  assign n15284 = ~n15281 & ~n15282;
  assign n15285 = ~n15283 & ~n15284;
  assign n15286 = ~n14906 & ~n15217;
  assign n15287 = n15285 & n15286;
  assign n15288 = ~n15285 & ~n15286;
  assign n15289 = ~n15287 & ~n15288;
  assign n15290 = pi121  & n918;
  assign n15291 = pi119  & n1031;
  assign n15292 = pi120  & n913;
  assign n15293 = ~n15291 & ~n15292;
  assign n15294 = ~n15290 & n15293;
  assign n15295 = n921 & n11086;
  assign n15296 = n15294 & ~n15295;
  assign n15297 = pi14  & ~n15296;
  assign n15298 = pi14  & ~n15297;
  assign n15299 = ~n15296 & ~n15297;
  assign n15300 = ~n15298 & ~n15299;
  assign n15301 = ~n15211 & ~n15214;
  assign n15302 = ~n15300 & ~n15301;
  assign n15303 = n15300 & n15301;
  assign n15304 = ~n15302 & ~n15303;
  assign n15305 = ~n14920 & ~n15196;
  assign n15306 = pi118  & n1269;
  assign n15307 = pi116  & n1340;
  assign n15308 = pi117  & n1264;
  assign n15309 = ~n15307 & ~n15308;
  assign n15310 = ~n15306 & n15309;
  assign n15311 = n1272 & n9716;
  assign n15312 = n15310 & ~n15311;
  assign n15313 = pi17  & ~n15312;
  assign n15314 = pi17  & ~n15313;
  assign n15315 = ~n15312 & ~n15313;
  assign n15316 = ~n15314 & ~n15315;
  assign n15317 = ~n15305 & ~n15316;
  assign n15318 = ~n15305 & ~n15317;
  assign n15319 = ~n15316 & ~n15317;
  assign n15320 = ~n15318 & ~n15319;
  assign n15321 = pi115  & n1582;
  assign n15322 = pi113  & n1713;
  assign n15323 = pi114  & n1577;
  assign n15324 = ~n15322 & ~n15323;
  assign n15325 = ~n15321 & n15324;
  assign n15326 = n1585 & n8727;
  assign n15327 = n15325 & ~n15326;
  assign n15328 = pi20  & ~n15327;
  assign n15329 = pi20  & ~n15328;
  assign n15330 = ~n15327 & ~n15328;
  assign n15331 = ~n15329 & ~n15330;
  assign n15332 = ~n14936 & ~n15193;
  assign n15333 = ~n15331 & n15332;
  assign n15334 = n15331 & ~n15332;
  assign n15335 = ~n15333 & ~n15334;
  assign n15336 = pi112  & n2004;
  assign n15337 = pi110  & n2141;
  assign n15338 = pi111  & n1999;
  assign n15339 = ~n15337 & ~n15338;
  assign n15340 = ~n15336 & n15339;
  assign n15341 = n2007 & n7795;
  assign n15342 = n15340 & ~n15341;
  assign n15343 = pi23  & ~n15342;
  assign n15344 = pi23  & ~n15343;
  assign n15345 = ~n15342 & ~n15343;
  assign n15346 = ~n15344 & ~n15345;
  assign n15347 = ~n14951 & ~n15190;
  assign n15348 = n15346 & n15347;
  assign n15349 = ~n15346 & ~n15347;
  assign n15350 = ~n15348 & ~n15349;
  assign n15351 = ~n15184 & ~n15187;
  assign n15352 = pi109  & n2486;
  assign n15353 = pi107  & n2644;
  assign n15354 = pi108  & n2481;
  assign n15355 = ~n15353 & ~n15354;
  assign n15356 = ~n15352 & n15355;
  assign n15357 = n2489 & n7170;
  assign n15358 = n15356 & ~n15357;
  assign n15359 = pi26  & ~n15358;
  assign n15360 = pi26  & ~n15359;
  assign n15361 = ~n15358 & ~n15359;
  assign n15362 = ~n15360 & ~n15361;
  assign n15363 = ~n15351 & ~n15362;
  assign n15364 = ~n15351 & ~n15363;
  assign n15365 = ~n15362 & ~n15363;
  assign n15366 = ~n15364 & ~n15365;
  assign n15367 = pi106  & n2976;
  assign n15368 = pi104  & n3182;
  assign n15369 = pi105  & n2971;
  assign n15370 = ~n15368 & ~n15369;
  assign n15371 = ~n15367 & n15370;
  assign n15372 = n2979 & n6090;
  assign n15373 = n15371 & ~n15372;
  assign n15374 = pi29  & ~n15373;
  assign n15375 = pi29  & ~n15374;
  assign n15376 = ~n15373 & ~n15374;
  assign n15377 = ~n15375 & ~n15376;
  assign n15378 = ~n14966 & ~n15169;
  assign n15379 = n15377 & n15378;
  assign n15380 = ~n15377 & ~n15378;
  assign n15381 = ~n15379 & ~n15380;
  assign n15382 = ~n15149 & ~n15163;
  assign n15383 = pi100  & n4182;
  assign n15384 = pi98  & n4416;
  assign n15385 = pi99  & n4177;
  assign n15386 = ~n15384 & ~n15385;
  assign n15387 = ~n15383 & n15386;
  assign n15388 = n4185 & n4808;
  assign n15389 = n15387 & ~n15388;
  assign n15390 = pi35  & ~n15389;
  assign n15391 = pi35  & ~n15390;
  assign n15392 = ~n15389 & ~n15390;
  assign n15393 = ~n15391 & ~n15392;
  assign n15394 = ~n15132 & ~n15146;
  assign n15395 = ~n15115 & ~n15128;
  assign n15396 = ~n15098 & ~n15111;
  assign n15397 = ~n15080 & ~n15094;
  assign n15398 = pi88  & n7239;
  assign n15399 = pi86  & n7556;
  assign n15400 = pi87  & n7234;
  assign n15401 = ~n15399 & ~n15400;
  assign n15402 = ~n15398 & n15401;
  assign n15403 = n2277 & n7242;
  assign n15404 = n15402 & ~n15403;
  assign n15405 = pi47  & ~n15404;
  assign n15406 = pi47  & ~n15405;
  assign n15407 = ~n15404 & ~n15405;
  assign n15408 = ~n15406 & ~n15407;
  assign n15409 = ~n15063 & ~n15077;
  assign n15410 = ~n15045 & ~n15059;
  assign n15411 = ~n15026 & ~n15040;
  assign n15412 = ~n15009 & ~n15023;
  assign n15413 = pi76  & n11193;
  assign n15414 = pi74  & n11567;
  assign n15415 = pi75  & n11188;
  assign n15416 = ~n15414 & ~n15415;
  assign n15417 = ~n15413 & n15416;
  assign n15418 = n881 & n11196;
  assign n15419 = n15417 & ~n15418;
  assign n15420 = pi59  & ~n15419;
  assign n15421 = pi59  & ~n15420;
  assign n15422 = ~n15419 & ~n15420;
  assign n15423 = ~n15421 & ~n15422;
  assign n15424 = ~n15002 & ~n15005;
  assign n15425 = pi69  & n13477;
  assign n15426 = pi70  & ~n13122;
  assign n15427 = ~n15425 & ~n15426;
  assign n15428 = pi2  & ~pi5 ;
  assign n15429 = ~pi2  & pi5 ;
  assign n15430 = ~n15428 & ~n15429;
  assign n15431 = ~n15427 & ~n15430;
  assign n15432 = n15427 & n15430;
  assign n15433 = ~n15431 & ~n15432;
  assign n15434 = n15424 & ~n15433;
  assign n15435 = ~n15424 & n15433;
  assign n15436 = ~n15434 & ~n15435;
  assign n15437 = pi73  & n12295;
  assign n15438 = pi71  & n12693;
  assign n15439 = pi72  & n12290;
  assign n15440 = ~n15438 & ~n15439;
  assign n15441 = ~n15437 & n15440;
  assign n15442 = n639 & n12298;
  assign n15443 = n15441 & ~n15442;
  assign n15444 = pi62  & ~n15443;
  assign n15445 = pi62  & ~n15444;
  assign n15446 = ~n15443 & ~n15444;
  assign n15447 = ~n15445 & ~n15446;
  assign n15448 = ~n15436 & n15447;
  assign n15449 = n15436 & ~n15447;
  assign n15450 = ~n15448 & ~n15449;
  assign n15451 = ~n15423 & n15450;
  assign n15452 = n15423 & ~n15450;
  assign n15453 = ~n15451 & ~n15452;
  assign n15454 = ~n15412 & n15453;
  assign n15455 = n15412 & ~n15453;
  assign n15456 = ~n15454 & ~n15455;
  assign n15457 = pi79  & n10135;
  assign n15458 = pi77  & n10478;
  assign n15459 = pi78  & n10130;
  assign n15460 = ~n15458 & ~n15459;
  assign n15461 = ~n15457 & n15460;
  assign n15462 = n1105 & n10138;
  assign n15463 = n15461 & ~n15462;
  assign n15464 = pi56  & ~n15463;
  assign n15465 = pi56  & ~n15464;
  assign n15466 = ~n15463 & ~n15464;
  assign n15467 = ~n15465 & ~n15466;
  assign n15468 = n15456 & ~n15467;
  assign n15469 = ~n15456 & n15467;
  assign n15470 = ~n15468 & ~n15469;
  assign n15471 = n15411 & ~n15470;
  assign n15472 = ~n15411 & n15470;
  assign n15473 = ~n15471 & ~n15472;
  assign n15474 = pi82  & n9096;
  assign n15475 = pi80  & n9453;
  assign n15476 = pi81  & n9091;
  assign n15477 = ~n15475 & ~n15476;
  assign n15478 = ~n15474 & n15477;
  assign n15479 = n1532 & n9099;
  assign n15480 = n15478 & ~n15479;
  assign n15481 = pi53  & ~n15480;
  assign n15482 = pi53  & ~n15481;
  assign n15483 = ~n15480 & ~n15481;
  assign n15484 = ~n15482 & ~n15483;
  assign n15485 = n15473 & ~n15484;
  assign n15486 = ~n15473 & n15484;
  assign n15487 = ~n15485 & ~n15486;
  assign n15488 = n15410 & ~n15487;
  assign n15489 = ~n15410 & n15487;
  assign n15490 = ~n15488 & ~n15489;
  assign n15491 = pi85  & n8137;
  assign n15492 = pi83  & n8471;
  assign n15493 = pi84  & n8132;
  assign n15494 = ~n15492 & ~n15493;
  assign n15495 = ~n15491 & n15494;
  assign n15496 = n1943 & n8140;
  assign n15497 = n15495 & ~n15496;
  assign n15498 = pi50  & ~n15497;
  assign n15499 = pi50  & ~n15498;
  assign n15500 = ~n15497 & ~n15498;
  assign n15501 = ~n15499 & ~n15500;
  assign n15502 = n15490 & ~n15501;
  assign n15503 = ~n15490 & n15501;
  assign n15504 = ~n15502 & ~n15503;
  assign n15505 = ~n15409 & n15504;
  assign n15506 = n15409 & ~n15504;
  assign n15507 = ~n15505 & ~n15506;
  assign n15508 = ~n15408 & n15507;
  assign n15509 = n15408 & ~n15507;
  assign n15510 = ~n15508 & ~n15509;
  assign n15511 = n15397 & ~n15510;
  assign n15512 = ~n15397 & n15510;
  assign n15513 = ~n15511 & ~n15512;
  assign n15514 = pi91  & n6396;
  assign n15515 = pi89  & n6735;
  assign n15516 = pi90  & n6391;
  assign n15517 = ~n15515 & ~n15516;
  assign n15518 = ~n15514 & n15517;
  assign n15519 = n2926 & n6399;
  assign n15520 = n15518 & ~n15519;
  assign n15521 = pi44  & ~n15520;
  assign n15522 = pi44  & ~n15521;
  assign n15523 = ~n15520 & ~n15521;
  assign n15524 = ~n15522 & ~n15523;
  assign n15525 = n15513 & ~n15524;
  assign n15526 = ~n15513 & n15524;
  assign n15527 = ~n15525 & ~n15526;
  assign n15528 = n15396 & ~n15527;
  assign n15529 = ~n15396 & n15527;
  assign n15530 = ~n15528 & ~n15529;
  assign n15531 = pi94  & n5636;
  assign n15532 = pi92  & n5909;
  assign n15533 = pi93  & n5631;
  assign n15534 = ~n15532 & ~n15533;
  assign n15535 = ~n15531 & n15534;
  assign n15536 = n3499 & n5639;
  assign n15537 = n15535 & ~n15536;
  assign n15538 = pi41  & ~n15537;
  assign n15539 = pi41  & ~n15538;
  assign n15540 = ~n15537 & ~n15538;
  assign n15541 = ~n15539 & ~n15540;
  assign n15542 = n15530 & ~n15541;
  assign n15543 = ~n15530 & n15541;
  assign n15544 = ~n15395 & ~n15543;
  assign n15545 = ~n15542 & n15544;
  assign n15546 = ~n15395 & ~n15545;
  assign n15547 = ~n15542 & ~n15545;
  assign n15548 = ~n15543 & n15547;
  assign n15549 = ~n15546 & ~n15548;
  assign n15550 = pi97  & n4896;
  assign n15551 = pi95  & n5148;
  assign n15552 = pi96  & n4891;
  assign n15553 = ~n15551 & ~n15552;
  assign n15554 = ~n15550 & n15553;
  assign n15555 = n3946 & n4899;
  assign n15556 = n15554 & ~n15555;
  assign n15557 = pi38  & ~n15556;
  assign n15558 = pi38  & ~n15557;
  assign n15559 = ~n15556 & ~n15557;
  assign n15560 = ~n15558 & ~n15559;
  assign n15561 = ~n15549 & ~n15560;
  assign n15562 = n15549 & n15560;
  assign n15563 = ~n15561 & ~n15562;
  assign n15564 = ~n15394 & n15563;
  assign n15565 = n15394 & ~n15563;
  assign n15566 = ~n15564 & ~n15565;
  assign n15567 = ~n15393 & n15566;
  assign n15568 = n15393 & ~n15566;
  assign n15569 = ~n15567 & ~n15568;
  assign n15570 = n15382 & ~n15569;
  assign n15571 = ~n15382 & n15569;
  assign n15572 = ~n15570 & ~n15571;
  assign n15573 = pi103  & n3550;
  assign n15574 = pi101  & n3735;
  assign n15575 = pi102  & n3545;
  assign n15576 = ~n15574 & ~n15575;
  assign n15577 = ~n15573 & n15576;
  assign n15578 = n3553 & n5540;
  assign n15579 = n15577 & ~n15578;
  assign n15580 = pi32  & ~n15579;
  assign n15581 = pi32  & ~n15580;
  assign n15582 = ~n15579 & ~n15580;
  assign n15583 = ~n15581 & ~n15582;
  assign n15584 = ~n14980 & ~n15166;
  assign n15585 = n15583 & n15584;
  assign n15586 = ~n15583 & ~n15584;
  assign n15587 = ~n15585 & ~n15586;
  assign n15588 = n15572 & n15587;
  assign n15589 = ~n15572 & ~n15587;
  assign n15590 = ~n15588 & ~n15589;
  assign n15591 = n15381 & n15590;
  assign n15592 = ~n15381 & ~n15590;
  assign n15593 = ~n15591 & ~n15592;
  assign n15594 = ~n15366 & n15593;
  assign n15595 = n15366 & ~n15593;
  assign n15596 = ~n15594 & ~n15595;
  assign n15597 = n15350 & n15596;
  assign n15598 = ~n15350 & ~n15596;
  assign n15599 = ~n15597 & ~n15598;
  assign n15600 = n15335 & n15599;
  assign n15601 = ~n15335 & ~n15599;
  assign n15602 = ~n15600 & ~n15601;
  assign n15603 = ~n15320 & n15602;
  assign n15604 = n15320 & ~n15602;
  assign n15605 = ~n15603 & ~n15604;
  assign n15606 = n15304 & n15605;
  assign n15607 = ~n15304 & ~n15605;
  assign n15608 = ~n15606 & ~n15607;
  assign n15609 = n15289 & n15608;
  assign n15610 = ~n15289 & ~n15608;
  assign n15611 = ~n15609 & ~n15610;
  assign n15612 = n15274 & n15611;
  assign n15613 = ~n15274 & ~n15611;
  assign n15614 = ~n15612 & ~n15613;
  assign n15615 = ~n15259 & n15614;
  assign n15616 = n15259 & ~n15614;
  assign n15617 = ~n15615 & ~n15616;
  assign n15618 = ~n15258 & n15617;
  assign n15619 = n15258 & ~n15617;
  assign po69  = ~n15618 & ~n15619;
  assign n15621 = ~n15615 & ~n15618;
  assign n15622 = ~n15288 & ~n15609;
  assign n15623 = pi126  & n533;
  assign n15624 = pi127  & n488;
  assign n15625 = ~n15623 & ~n15624;
  assign n15626 = ~n496 & n15625;
  assign n15627 = ~n13389 & n15625;
  assign n15628 = ~n15626 & ~n15627;
  assign n15629 = pi8  & ~n15628;
  assign n15630 = ~pi8  & n15628;
  assign n15631 = ~n15629 & ~n15630;
  assign n15632 = ~n15622 & ~n15631;
  assign n15633 = n15622 & n15631;
  assign n15634 = ~n15632 & ~n15633;
  assign n15635 = pi125  & n675;
  assign n15636 = pi123  & n769;
  assign n15637 = pi124  & n670;
  assign n15638 = ~n15636 & ~n15637;
  assign n15639 = ~n15635 & n15638;
  assign n15640 = n678 & n12591;
  assign n15641 = n15639 & ~n15640;
  assign n15642 = pi11  & ~n15641;
  assign n15643 = pi11  & ~n15642;
  assign n15644 = ~n15641 & ~n15642;
  assign n15645 = ~n15643 & ~n15644;
  assign n15646 = ~n15302 & ~n15606;
  assign n15647 = n15645 & n15646;
  assign n15648 = ~n15645 & ~n15646;
  assign n15649 = ~n15647 & ~n15648;
  assign n15650 = ~n15317 & ~n15603;
  assign n15651 = pi122  & n918;
  assign n15652 = pi120  & n1031;
  assign n15653 = pi121  & n913;
  assign n15654 = ~n15652 & ~n15653;
  assign n15655 = ~n15651 & n15654;
  assign n15656 = ~n921 & n15655;
  assign n15657 = ~n11463 & n15655;
  assign n15658 = ~n15656 & ~n15657;
  assign n15659 = pi14  & ~n15658;
  assign n15660 = ~pi14  & n15658;
  assign n15661 = ~n15659 & ~n15660;
  assign n15662 = ~n15650 & ~n15661;
  assign n15663 = n15650 & n15661;
  assign n15664 = ~n15662 & ~n15663;
  assign n15665 = pi119  & n1269;
  assign n15666 = pi117  & n1340;
  assign n15667 = pi118  & n1264;
  assign n15668 = ~n15666 & ~n15667;
  assign n15669 = ~n15665 & n15668;
  assign n15670 = n1272 & n10048;
  assign n15671 = n15669 & ~n15670;
  assign n15672 = pi17  & ~n15671;
  assign n15673 = pi17  & ~n15672;
  assign n15674 = ~n15671 & ~n15672;
  assign n15675 = ~n15673 & ~n15674;
  assign n15676 = ~n15333 & ~n15600;
  assign n15677 = n15675 & n15676;
  assign n15678 = ~n15675 & ~n15676;
  assign n15679 = ~n15677 & ~n15678;
  assign n15680 = pi116  & n1582;
  assign n15681 = pi114  & n1713;
  assign n15682 = pi115  & n1577;
  assign n15683 = ~n15681 & ~n15682;
  assign n15684 = ~n15680 & n15683;
  assign n15685 = n1585 & n9042;
  assign n15686 = n15684 & ~n15685;
  assign n15687 = pi20  & ~n15686;
  assign n15688 = pi20  & ~n15687;
  assign n15689 = ~n15686 & ~n15687;
  assign n15690 = ~n15688 & ~n15689;
  assign n15691 = ~n15349 & ~n15597;
  assign n15692 = n15690 & n15691;
  assign n15693 = ~n15690 & ~n15691;
  assign n15694 = ~n15692 & ~n15693;
  assign n15695 = pi113  & n2004;
  assign n15696 = pi111  & n2141;
  assign n15697 = pi112  & n1999;
  assign n15698 = ~n15696 & ~n15697;
  assign n15699 = ~n15695 & n15698;
  assign n15700 = n2007 & n8387;
  assign n15701 = n15699 & ~n15700;
  assign n15702 = pi23  & ~n15701;
  assign n15703 = pi23  & ~n15702;
  assign n15704 = ~n15701 & ~n15702;
  assign n15705 = ~n15703 & ~n15704;
  assign n15706 = ~n15363 & ~n15594;
  assign n15707 = ~n15705 & ~n15706;
  assign n15708 = n15705 & n15706;
  assign n15709 = ~n15707 & ~n15708;
  assign n15710 = ~n15380 & ~n15591;
  assign n15711 = pi110  & n2486;
  assign n15712 = pi108  & n2644;
  assign n15713 = pi109  & n2481;
  assign n15714 = ~n15712 & ~n15713;
  assign n15715 = ~n15711 & n15714;
  assign n15716 = ~n2489 & n15715;
  assign n15717 = ~n7474 & n15715;
  assign n15718 = ~n15716 & ~n15717;
  assign n15719 = pi26  & ~n15718;
  assign n15720 = ~pi26  & n15718;
  assign n15721 = ~n15719 & ~n15720;
  assign n15722 = ~n15710 & ~n15721;
  assign n15723 = n15710 & n15721;
  assign n15724 = ~n15722 & ~n15723;
  assign n15725 = pi107  & n2976;
  assign n15726 = pi105  & n3182;
  assign n15727 = pi106  & n2971;
  assign n15728 = ~n15726 & ~n15727;
  assign n15729 = ~n15725 & n15728;
  assign n15730 = n2979 & n6614;
  assign n15731 = n15729 & ~n15730;
  assign n15732 = pi29  & ~n15731;
  assign n15733 = pi29  & ~n15732;
  assign n15734 = ~n15731 & ~n15732;
  assign n15735 = ~n15733 & ~n15734;
  assign n15736 = ~n15586 & ~n15588;
  assign n15737 = ~n15735 & ~n15736;
  assign n15738 = n15735 & n15736;
  assign n15739 = ~n15737 & ~n15738;
  assign n15740 = pi104  & n3550;
  assign n15741 = pi102  & n3735;
  assign n15742 = pi103  & n3545;
  assign n15743 = ~n15741 & ~n15742;
  assign n15744 = ~n15740 & n15743;
  assign n15745 = n3553 & n5565;
  assign n15746 = n15744 & ~n15745;
  assign n15747 = pi32  & ~n15746;
  assign n15748 = pi32  & ~n15747;
  assign n15749 = ~n15746 & ~n15747;
  assign n15750 = ~n15748 & ~n15749;
  assign n15751 = ~n15567 & ~n15571;
  assign n15752 = n15750 & n15751;
  assign n15753 = ~n15750 & ~n15751;
  assign n15754 = ~n15752 & ~n15753;
  assign n15755 = pi101  & n4182;
  assign n15756 = pi99  & n4416;
  assign n15757 = pi100  & n4177;
  assign n15758 = ~n15756 & ~n15757;
  assign n15759 = ~n15755 & n15758;
  assign n15760 = n4185 & n5056;
  assign n15761 = n15759 & ~n15760;
  assign n15762 = pi35  & ~n15761;
  assign n15763 = pi35  & ~n15762;
  assign n15764 = ~n15761 & ~n15762;
  assign n15765 = ~n15763 & ~n15764;
  assign n15766 = ~n15561 & ~n15564;
  assign n15767 = pi98  & n4896;
  assign n15768 = pi96  & n5148;
  assign n15769 = pi97  & n4891;
  assign n15770 = ~n15768 & ~n15769;
  assign n15771 = ~n15767 & n15770;
  assign n15772 = n4360 & n4899;
  assign n15773 = n15771 & ~n15772;
  assign n15774 = pi38  & ~n15773;
  assign n15775 = pi38  & ~n15774;
  assign n15776 = ~n15773 & ~n15774;
  assign n15777 = ~n15775 & ~n15776;
  assign n15778 = ~n15525 & ~n15529;
  assign n15779 = ~n15508 & ~n15512;
  assign n15780 = ~n15502 & ~n15505;
  assign n15781 = ~n15485 & ~n15489;
  assign n15782 = ~n15468 & ~n15472;
  assign n15783 = ~n15435 & ~n15449;
  assign n15784 = ~pi2  & ~pi5 ;
  assign n15785 = ~n15431 & ~n15784;
  assign n15786 = pi70  & n13477;
  assign n15787 = pi71  & ~n13122;
  assign n15788 = ~n15786 & ~n15787;
  assign n15789 = ~n15785 & n15788;
  assign n15790 = n15785 & ~n15788;
  assign n15791 = ~n15789 & ~n15790;
  assign n15792 = pi74  & n12295;
  assign n15793 = pi72  & n12693;
  assign n15794 = pi73  & n12290;
  assign n15795 = ~n15793 & ~n15794;
  assign n15796 = ~n15792 & n15795;
  assign n15797 = ~n12298 & n15796;
  assign n15798 = ~n722 & n15796;
  assign n15799 = ~n15797 & ~n15798;
  assign n15800 = pi62  & ~n15799;
  assign n15801 = ~pi62  & n15799;
  assign n15802 = ~n15800 & ~n15801;
  assign n15803 = n15791 & ~n15802;
  assign n15804 = ~n15791 & n15802;
  assign n15805 = ~n15803 & ~n15804;
  assign n15806 = ~n15783 & n15805;
  assign n15807 = n15783 & ~n15805;
  assign n15808 = ~n15806 & ~n15807;
  assign n15809 = pi77  & n11193;
  assign n15810 = pi75  & n11567;
  assign n15811 = pi76  & n11188;
  assign n15812 = ~n15810 & ~n15811;
  assign n15813 = ~n15809 & n15812;
  assign n15814 = n984 & n11196;
  assign n15815 = n15813 & ~n15814;
  assign n15816 = pi59  & ~n15815;
  assign n15817 = pi59  & ~n15816;
  assign n15818 = ~n15815 & ~n15816;
  assign n15819 = ~n15817 & ~n15818;
  assign n15820 = n15808 & ~n15819;
  assign n15821 = n15808 & ~n15820;
  assign n15822 = ~n15819 & ~n15820;
  assign n15823 = ~n15821 & ~n15822;
  assign n15824 = ~n15451 & ~n15454;
  assign n15825 = n15823 & n15824;
  assign n15826 = ~n15823 & ~n15824;
  assign n15827 = ~n15825 & ~n15826;
  assign n15828 = pi80  & n10135;
  assign n15829 = pi78  & n10478;
  assign n15830 = pi79  & n10130;
  assign n15831 = ~n15829 & ~n15830;
  assign n15832 = ~n15828 & n15831;
  assign n15833 = n1205 & n10138;
  assign n15834 = n15832 & ~n15833;
  assign n15835 = pi56  & ~n15834;
  assign n15836 = pi56  & ~n15835;
  assign n15837 = ~n15834 & ~n15835;
  assign n15838 = ~n15836 & ~n15837;
  assign n15839 = n15827 & ~n15838;
  assign n15840 = ~n15827 & n15838;
  assign n15841 = ~n15839 & ~n15840;
  assign n15842 = n15782 & ~n15841;
  assign n15843 = ~n15782 & n15841;
  assign n15844 = ~n15842 & ~n15843;
  assign n15845 = pi83  & n9096;
  assign n15846 = pi81  & n9453;
  assign n15847 = pi82  & n9091;
  assign n15848 = ~n15846 & ~n15847;
  assign n15849 = ~n15845 & n15848;
  assign n15850 = n1672 & n9099;
  assign n15851 = n15849 & ~n15850;
  assign n15852 = pi53  & ~n15851;
  assign n15853 = pi53  & ~n15852;
  assign n15854 = ~n15851 & ~n15852;
  assign n15855 = ~n15853 & ~n15854;
  assign n15856 = n15844 & ~n15855;
  assign n15857 = ~n15844 & n15855;
  assign n15858 = ~n15856 & ~n15857;
  assign n15859 = n15781 & ~n15858;
  assign n15860 = ~n15781 & n15858;
  assign n15861 = ~n15859 & ~n15860;
  assign n15862 = pi86  & n8137;
  assign n15863 = pi84  & n8471;
  assign n15864 = pi85  & n8132;
  assign n15865 = ~n15863 & ~n15864;
  assign n15866 = ~n15862 & n15865;
  assign n15867 = n2099 & n8140;
  assign n15868 = n15866 & ~n15867;
  assign n15869 = pi50  & ~n15868;
  assign n15870 = pi50  & ~n15869;
  assign n15871 = ~n15868 & ~n15869;
  assign n15872 = ~n15870 & ~n15871;
  assign n15873 = n15861 & ~n15872;
  assign n15874 = ~n15861 & n15872;
  assign n15875 = ~n15873 & ~n15874;
  assign n15876 = n15780 & ~n15875;
  assign n15877 = ~n15780 & n15875;
  assign n15878 = ~n15876 & ~n15877;
  assign n15879 = pi89  & n7239;
  assign n15880 = pi87  & n7556;
  assign n15881 = pi88  & n7234;
  assign n15882 = ~n15880 & ~n15881;
  assign n15883 = ~n15879 & n15882;
  assign n15884 = n2432 & n7242;
  assign n15885 = n15883 & ~n15884;
  assign n15886 = pi47  & ~n15885;
  assign n15887 = pi47  & ~n15886;
  assign n15888 = ~n15885 & ~n15886;
  assign n15889 = ~n15887 & ~n15888;
  assign n15890 = n15878 & ~n15889;
  assign n15891 = ~n15878 & n15889;
  assign n15892 = ~n15890 & ~n15891;
  assign n15893 = n15779 & ~n15892;
  assign n15894 = ~n15779 & n15892;
  assign n15895 = ~n15893 & ~n15894;
  assign n15896 = pi92  & n6396;
  assign n15897 = pi90  & n6735;
  assign n15898 = pi91  & n6391;
  assign n15899 = ~n15897 & ~n15898;
  assign n15900 = ~n15896 & n15899;
  assign n15901 = n3119 & n6399;
  assign n15902 = n15900 & ~n15901;
  assign n15903 = pi44  & ~n15902;
  assign n15904 = pi44  & ~n15903;
  assign n15905 = ~n15902 & ~n15903;
  assign n15906 = ~n15904 & ~n15905;
  assign n15907 = n15895 & ~n15906;
  assign n15908 = ~n15895 & n15906;
  assign n15909 = ~n15907 & ~n15908;
  assign n15910 = n15778 & ~n15909;
  assign n15911 = ~n15778 & n15909;
  assign n15912 = ~n15910 & ~n15911;
  assign n15913 = pi95  & n5636;
  assign n15914 = pi93  & n5909;
  assign n15915 = pi94  & n5631;
  assign n15916 = ~n15914 & ~n15915;
  assign n15917 = ~n15913 & n15916;
  assign n15918 = n3710 & n5639;
  assign n15919 = n15917 & ~n15918;
  assign n15920 = pi41  & ~n15919;
  assign n15921 = pi41  & ~n15920;
  assign n15922 = ~n15919 & ~n15920;
  assign n15923 = ~n15921 & ~n15922;
  assign n15924 = ~n15912 & n15923;
  assign n15925 = n15912 & ~n15923;
  assign n15926 = ~n15924 & ~n15925;
  assign n15927 = ~n15547 & n15926;
  assign n15928 = n15547 & ~n15926;
  assign n15929 = ~n15927 & ~n15928;
  assign n15930 = ~n15777 & n15929;
  assign n15931 = n15777 & ~n15929;
  assign n15932 = ~n15930 & ~n15931;
  assign n15933 = ~n15766 & n15932;
  assign n15934 = n15766 & ~n15932;
  assign n15935 = ~n15933 & ~n15934;
  assign n15936 = ~n15765 & n15935;
  assign n15937 = n15765 & ~n15935;
  assign n15938 = ~n15936 & ~n15937;
  assign n15939 = n15754 & n15938;
  assign n15940 = ~n15754 & ~n15938;
  assign n15941 = ~n15939 & ~n15940;
  assign n15942 = n15739 & ~n15941;
  assign n15943 = ~n15739 & n15941;
  assign n15944 = ~n15942 & ~n15943;
  assign n15945 = n15724 & ~n15944;
  assign n15946 = ~n15724 & n15944;
  assign n15947 = ~n15945 & ~n15946;
  assign n15948 = n15709 & n15947;
  assign n15949 = ~n15709 & ~n15947;
  assign n15950 = ~n15948 & ~n15949;
  assign n15951 = n15694 & n15950;
  assign n15952 = ~n15694 & ~n15950;
  assign n15953 = ~n15951 & ~n15952;
  assign n15954 = n15679 & n15953;
  assign n15955 = ~n15679 & ~n15953;
  assign n15956 = n15664 & ~n15955;
  assign n15957 = ~n15954 & n15956;
  assign n15958 = n15664 & ~n15957;
  assign n15959 = ~n15955 & ~n15957;
  assign n15960 = ~n15954 & n15959;
  assign n15961 = ~n15958 & ~n15960;
  assign n15962 = n15649 & ~n15961;
  assign n15963 = ~n15649 & n15961;
  assign n15964 = n15634 & ~n15963;
  assign n15965 = ~n15962 & n15964;
  assign n15966 = n15634 & ~n15965;
  assign n15967 = ~n15963 & ~n15965;
  assign n15968 = ~n15962 & n15967;
  assign n15969 = ~n15966 & ~n15968;
  assign n15970 = ~n15272 & ~n15612;
  assign n15971 = ~n15969 & ~n15970;
  assign n15972 = n15969 & n15970;
  assign n15973 = ~n15971 & ~n15972;
  assign n15974 = ~n15621 & n15973;
  assign n15975 = n15621 & ~n15973;
  assign po70  = ~n15974 & ~n15975;
  assign n15977 = ~n15971 & ~n15974;
  assign n15978 = ~n15632 & ~n15965;
  assign n15979 = ~n15662 & ~n15957;
  assign n15980 = pi126  & n675;
  assign n15981 = pi124  & n769;
  assign n15982 = pi125  & n670;
  assign n15983 = ~n15981 & ~n15982;
  assign n15984 = ~n15980 & n15983;
  assign n15985 = ~n678 & n15984;
  assign n15986 = ~n12979 & n15984;
  assign n15987 = ~n15985 & ~n15986;
  assign n15988 = pi11  & ~n15987;
  assign n15989 = ~pi11  & n15987;
  assign n15990 = ~n15988 & ~n15989;
  assign n15991 = ~n15979 & ~n15990;
  assign n15992 = ~n15979 & ~n15991;
  assign n15993 = ~n15990 & ~n15991;
  assign n15994 = ~n15992 & ~n15993;
  assign n15995 = pi120  & n1269;
  assign n15996 = pi118  & n1340;
  assign n15997 = pi119  & n1264;
  assign n15998 = ~n15996 & ~n15997;
  assign n15999 = ~n15995 & n15998;
  assign n16000 = n1272 & n10734;
  assign n16001 = n15999 & ~n16000;
  assign n16002 = pi17  & ~n16001;
  assign n16003 = pi17  & ~n16002;
  assign n16004 = ~n16001 & ~n16002;
  assign n16005 = ~n16003 & ~n16004;
  assign n16006 = ~n15693 & ~n15951;
  assign n16007 = n16005 & n16006;
  assign n16008 = ~n16005 & ~n16006;
  assign n16009 = ~n16007 & ~n16008;
  assign n16010 = pi114  & n2004;
  assign n16011 = pi112  & n2141;
  assign n16012 = pi113  & n1999;
  assign n16013 = ~n16011 & ~n16012;
  assign n16014 = ~n16010 & n16013;
  assign n16015 = n2007 & n8702;
  assign n16016 = n16014 & ~n16015;
  assign n16017 = pi23  & ~n16016;
  assign n16018 = pi23  & ~n16017;
  assign n16019 = ~n16016 & ~n16017;
  assign n16020 = ~n16018 & ~n16019;
  assign n16021 = ~n15722 & ~n15945;
  assign n16022 = n16020 & n16021;
  assign n16023 = ~n16020 & ~n16021;
  assign n16024 = ~n16022 & ~n16023;
  assign n16025 = pi111  & n2486;
  assign n16026 = pi109  & n2644;
  assign n16027 = pi110  & n2481;
  assign n16028 = ~n16026 & ~n16027;
  assign n16029 = ~n16025 & n16028;
  assign n16030 = n2489 & n7770;
  assign n16031 = n16029 & ~n16030;
  assign n16032 = pi26  & ~n16031;
  assign n16033 = pi26  & ~n16032;
  assign n16034 = ~n16031 & ~n16032;
  assign n16035 = ~n16033 & ~n16034;
  assign n16036 = ~n15738 & ~n15942;
  assign n16037 = ~n16035 & n16036;
  assign n16038 = ~n16035 & ~n16037;
  assign n16039 = n16036 & ~n16037;
  assign n16040 = ~n16038 & ~n16039;
  assign n16041 = pi105  & n3550;
  assign n16042 = pi103  & n3735;
  assign n16043 = pi104  & n3545;
  assign n16044 = ~n16042 & ~n16043;
  assign n16045 = ~n16041 & n16044;
  assign n16046 = n3553 & n6065;
  assign n16047 = n16045 & ~n16046;
  assign n16048 = pi32  & ~n16047;
  assign n16049 = pi32  & ~n16048;
  assign n16050 = ~n16047 & ~n16048;
  assign n16051 = ~n16049 & ~n16050;
  assign n16052 = ~n15933 & ~n15936;
  assign n16053 = n16051 & n16052;
  assign n16054 = ~n16051 & ~n16052;
  assign n16055 = ~n16053 & ~n16054;
  assign n16056 = ~n15894 & ~n15907;
  assign n16057 = ~n15877 & ~n15890;
  assign n16058 = ~n15860 & ~n15873;
  assign n16059 = pi87  & n8137;
  assign n16060 = pi85  & n8471;
  assign n16061 = pi86  & n8132;
  assign n16062 = ~n16060 & ~n16061;
  assign n16063 = ~n16059 & n16062;
  assign n16064 = n2252 & n8140;
  assign n16065 = n16063 & ~n16064;
  assign n16066 = pi50  & ~n16065;
  assign n16067 = pi50  & ~n16066;
  assign n16068 = ~n16065 & ~n16066;
  assign n16069 = ~n16067 & ~n16068;
  assign n16070 = ~n15843 & ~n15856;
  assign n16071 = ~n15826 & ~n15839;
  assign n16072 = ~n15806 & ~n15820;
  assign n16073 = pi78  & n11193;
  assign n16074 = pi76  & n11567;
  assign n16075 = pi77  & n11188;
  assign n16076 = ~n16074 & ~n16075;
  assign n16077 = ~n16073 & n16076;
  assign n16078 = n1009 & n11196;
  assign n16079 = n16077 & ~n16078;
  assign n16080 = pi59  & ~n16079;
  assign n16081 = pi59  & ~n16080;
  assign n16082 = ~n16079 & ~n16080;
  assign n16083 = ~n16081 & ~n16082;
  assign n16084 = ~n15789 & ~n15803;
  assign n16085 = pi71  & n13477;
  assign n16086 = pi72  & ~n13122;
  assign n16087 = ~n16085 & ~n16086;
  assign n16088 = n15788 & ~n16087;
  assign n16089 = ~n15788 & n16087;
  assign n16090 = ~n16084 & ~n16089;
  assign n16091 = ~n16088 & n16090;
  assign n16092 = ~n16084 & ~n16091;
  assign n16093 = ~n16089 & ~n16091;
  assign n16094 = ~n16088 & n16093;
  assign n16095 = ~n16092 & ~n16094;
  assign n16096 = pi75  & n12295;
  assign n16097 = pi73  & n12693;
  assign n16098 = pi74  & n12290;
  assign n16099 = ~n16097 & ~n16098;
  assign n16100 = ~n16096 & n16099;
  assign n16101 = n747 & n12298;
  assign n16102 = n16100 & ~n16101;
  assign n16103 = pi62  & ~n16102;
  assign n16104 = pi62  & ~n16103;
  assign n16105 = ~n16102 & ~n16103;
  assign n16106 = ~n16104 & ~n16105;
  assign n16107 = ~n16095 & ~n16106;
  assign n16108 = n16095 & n16106;
  assign n16109 = ~n16107 & ~n16108;
  assign n16110 = ~n16083 & n16109;
  assign n16111 = n16083 & ~n16109;
  assign n16112 = ~n16110 & ~n16111;
  assign n16113 = n16072 & ~n16112;
  assign n16114 = ~n16072 & n16112;
  assign n16115 = ~n16113 & ~n16114;
  assign n16116 = pi81  & n10135;
  assign n16117 = pi79  & n10478;
  assign n16118 = pi80  & n10130;
  assign n16119 = ~n16117 & ~n16118;
  assign n16120 = ~n16116 & n16119;
  assign n16121 = n1413 & n10138;
  assign n16122 = n16120 & ~n16121;
  assign n16123 = pi56  & ~n16122;
  assign n16124 = pi56  & ~n16123;
  assign n16125 = ~n16122 & ~n16123;
  assign n16126 = ~n16124 & ~n16125;
  assign n16127 = n16115 & ~n16126;
  assign n16128 = ~n16115 & n16126;
  assign n16129 = ~n16127 & ~n16128;
  assign n16130 = n16071 & ~n16129;
  assign n16131 = ~n16071 & n16129;
  assign n16132 = ~n16130 & ~n16131;
  assign n16133 = pi84  & n9096;
  assign n16134 = pi82  & n9453;
  assign n16135 = pi83  & n9091;
  assign n16136 = ~n16134 & ~n16135;
  assign n16137 = ~n16133 & n16136;
  assign n16138 = n1805 & n9099;
  assign n16139 = n16137 & ~n16138;
  assign n16140 = pi53  & ~n16139;
  assign n16141 = pi53  & ~n16140;
  assign n16142 = ~n16139 & ~n16140;
  assign n16143 = ~n16141 & ~n16142;
  assign n16144 = ~n16132 & n16143;
  assign n16145 = n16132 & ~n16143;
  assign n16146 = ~n16144 & ~n16145;
  assign n16147 = ~n16070 & n16146;
  assign n16148 = n16070 & ~n16146;
  assign n16149 = ~n16147 & ~n16148;
  assign n16150 = ~n16069 & n16149;
  assign n16151 = n16069 & ~n16149;
  assign n16152 = ~n16150 & ~n16151;
  assign n16153 = ~n16058 & n16152;
  assign n16154 = n16058 & ~n16152;
  assign n16155 = ~n16153 & ~n16154;
  assign n16156 = pi90  & n7239;
  assign n16157 = pi88  & n7556;
  assign n16158 = pi89  & n7234;
  assign n16159 = ~n16157 & ~n16158;
  assign n16160 = ~n16156 & n16159;
  assign n16161 = n2606 & n7242;
  assign n16162 = n16160 & ~n16161;
  assign n16163 = pi47  & ~n16162;
  assign n16164 = pi47  & ~n16163;
  assign n16165 = ~n16162 & ~n16163;
  assign n16166 = ~n16164 & ~n16165;
  assign n16167 = n16155 & ~n16166;
  assign n16168 = ~n16155 & n16166;
  assign n16169 = ~n16167 & ~n16168;
  assign n16170 = n16057 & ~n16169;
  assign n16171 = ~n16057 & n16169;
  assign n16172 = ~n16170 & ~n16171;
  assign n16173 = pi93  & n6396;
  assign n16174 = pi91  & n6735;
  assign n16175 = pi92  & n6391;
  assign n16176 = ~n16174 & ~n16175;
  assign n16177 = ~n16173 & n16176;
  assign n16178 = n3144 & n6399;
  assign n16179 = n16177 & ~n16178;
  assign n16180 = pi44  & ~n16179;
  assign n16181 = pi44  & ~n16180;
  assign n16182 = ~n16179 & ~n16180;
  assign n16183 = ~n16181 & ~n16182;
  assign n16184 = n16172 & ~n16183;
  assign n16185 = ~n16172 & n16183;
  assign n16186 = ~n16184 & ~n16185;
  assign n16187 = n16056 & ~n16186;
  assign n16188 = ~n16056 & n16186;
  assign n16189 = ~n16187 & ~n16188;
  assign n16190 = pi96  & n5636;
  assign n16191 = pi94  & n5909;
  assign n16192 = pi95  & n5631;
  assign n16193 = ~n16191 & ~n16192;
  assign n16194 = ~n16190 & n16193;
  assign n16195 = n3921 & n5639;
  assign n16196 = n16194 & ~n16195;
  assign n16197 = pi41  & ~n16196;
  assign n16198 = pi41  & ~n16197;
  assign n16199 = ~n16196 & ~n16197;
  assign n16200 = ~n16198 & ~n16199;
  assign n16201 = ~n16189 & n16200;
  assign n16202 = n16189 & ~n16200;
  assign n16203 = ~n16201 & ~n16202;
  assign n16204 = ~n15911 & ~n15925;
  assign n16205 = n16203 & ~n16204;
  assign n16206 = ~n16203 & n16204;
  assign n16207 = ~n16205 & ~n16206;
  assign n16208 = pi99  & n4896;
  assign n16209 = pi97  & n5148;
  assign n16210 = pi98  & n4891;
  assign n16211 = ~n16209 & ~n16210;
  assign n16212 = ~n16208 & n16211;
  assign n16213 = n4584 & n4899;
  assign n16214 = n16212 & ~n16213;
  assign n16215 = pi38  & ~n16214;
  assign n16216 = pi38  & ~n16215;
  assign n16217 = ~n16214 & ~n16215;
  assign n16218 = ~n16216 & ~n16217;
  assign n16219 = n16207 & ~n16218;
  assign n16220 = n16207 & ~n16219;
  assign n16221 = ~n16218 & ~n16219;
  assign n16222 = ~n16220 & ~n16221;
  assign n16223 = ~n15927 & ~n15930;
  assign n16224 = n16222 & n16223;
  assign n16225 = ~n16222 & ~n16223;
  assign n16226 = ~n16224 & ~n16225;
  assign n16227 = pi102  & n4182;
  assign n16228 = pi100  & n4416;
  assign n16229 = pi101  & n4177;
  assign n16230 = ~n16228 & ~n16229;
  assign n16231 = ~n16227 & n16230;
  assign n16232 = n4185 & n5296;
  assign n16233 = n16231 & ~n16232;
  assign n16234 = pi35  & ~n16233;
  assign n16235 = pi35  & ~n16234;
  assign n16236 = ~n16233 & ~n16234;
  assign n16237 = ~n16235 & ~n16236;
  assign n16238 = n16226 & ~n16237;
  assign n16239 = ~n16226 & n16237;
  assign n16240 = n16055 & ~n16239;
  assign n16241 = ~n16238 & n16240;
  assign n16242 = n16055 & ~n16241;
  assign n16243 = ~n16239 & ~n16241;
  assign n16244 = ~n16238 & n16243;
  assign n16245 = ~n16242 & ~n16244;
  assign n16246 = ~n15753 & ~n15939;
  assign n16247 = pi108  & n2976;
  assign n16248 = pi106  & n3182;
  assign n16249 = pi107  & n2971;
  assign n16250 = ~n16248 & ~n16249;
  assign n16251 = ~n16247 & n16250;
  assign n16252 = ~n2979 & n16251;
  assign n16253 = ~n6639 & n16251;
  assign n16254 = ~n16252 & ~n16253;
  assign n16255 = pi29  & ~n16254;
  assign n16256 = ~pi29  & n16254;
  assign n16257 = ~n16255 & ~n16256;
  assign n16258 = ~n16246 & ~n16257;
  assign n16259 = n16246 & n16257;
  assign n16260 = ~n16258 & ~n16259;
  assign n16261 = ~n16245 & n16260;
  assign n16262 = n16245 & ~n16260;
  assign n16263 = ~n16261 & ~n16262;
  assign n16264 = ~n16040 & n16263;
  assign n16265 = ~n16040 & ~n16264;
  assign n16266 = n16263 & ~n16264;
  assign n16267 = ~n16265 & ~n16266;
  assign n16268 = ~n16024 & n16267;
  assign n16269 = n16024 & ~n16267;
  assign n16270 = ~n16268 & ~n16269;
  assign n16271 = ~n15707 & ~n15948;
  assign n16272 = pi117  & n1582;
  assign n16273 = pi115  & n1713;
  assign n16274 = pi116  & n1577;
  assign n16275 = ~n16273 & ~n16274;
  assign n16276 = ~n16272 & n16275;
  assign n16277 = ~n1585 & n16276;
  assign n16278 = ~n9691 & n16276;
  assign n16279 = ~n16277 & ~n16278;
  assign n16280 = pi20  & ~n16279;
  assign n16281 = ~pi20  & n16279;
  assign n16282 = ~n16280 & ~n16281;
  assign n16283 = ~n16271 & ~n16282;
  assign n16284 = n16271 & n16282;
  assign n16285 = ~n16283 & ~n16284;
  assign n16286 = n16270 & n16285;
  assign n16287 = ~n16270 & ~n16285;
  assign n16288 = ~n16286 & ~n16287;
  assign n16289 = n16009 & n16288;
  assign n16290 = ~n16009 & ~n16288;
  assign n16291 = ~n16289 & ~n16290;
  assign n16292 = pi123  & n918;
  assign n16293 = pi121  & n1031;
  assign n16294 = pi122  & n913;
  assign n16295 = ~n16293 & ~n16294;
  assign n16296 = ~n16292 & n16295;
  assign n16297 = n921 & n11489;
  assign n16298 = n16296 & ~n16297;
  assign n16299 = pi14  & ~n16298;
  assign n16300 = pi14  & ~n16299;
  assign n16301 = ~n16298 & ~n16299;
  assign n16302 = ~n16300 & ~n16301;
  assign n16303 = ~n15678 & ~n15954;
  assign n16304 = ~n16302 & ~n16303;
  assign n16305 = n16302 & n16303;
  assign n16306 = ~n16304 & ~n16305;
  assign n16307 = n16291 & n16306;
  assign n16308 = ~n16291 & ~n16306;
  assign n16309 = ~n16307 & ~n16308;
  assign n16310 = ~n15994 & n16309;
  assign n16311 = n15994 & ~n16309;
  assign n16312 = ~n16310 & ~n16311;
  assign n16313 = ~n15648 & ~n15962;
  assign n16314 = pi127  & n533;
  assign n16315 = n496 & n13387;
  assign n16316 = ~n16314 & ~n16315;
  assign n16317 = pi8  & ~n16316;
  assign n16318 = pi8  & ~n16317;
  assign n16319 = ~n16316 & ~n16317;
  assign n16320 = ~n16318 & ~n16319;
  assign n16321 = ~n16313 & ~n16320;
  assign n16322 = n16313 & n16320;
  assign n16323 = ~n16321 & ~n16322;
  assign n16324 = n16312 & n16323;
  assign n16325 = ~n16312 & ~n16323;
  assign n16326 = ~n16324 & ~n16325;
  assign n16327 = ~n15978 & n16326;
  assign n16328 = n15978 & ~n16326;
  assign n16329 = ~n16327 & ~n16328;
  assign n16330 = ~n15977 & n16329;
  assign n16331 = n15977 & ~n16329;
  assign po71  = ~n16330 & ~n16331;
  assign n16333 = ~n16327 & ~n16330;
  assign n16334 = ~n16321 & ~n16324;
  assign n16335 = ~n16304 & ~n16307;
  assign n16336 = pi124  & n918;
  assign n16337 = pi122  & n1031;
  assign n16338 = pi123  & n913;
  assign n16339 = ~n16337 & ~n16338;
  assign n16340 = ~n16336 & n16339;
  assign n16341 = n921 & n11858;
  assign n16342 = n16340 & ~n16341;
  assign n16343 = pi14  & ~n16342;
  assign n16344 = pi14  & ~n16343;
  assign n16345 = ~n16342 & ~n16343;
  assign n16346 = ~n16344 & ~n16345;
  assign n16347 = ~n16335 & n16346;
  assign n16348 = n16335 & ~n16346;
  assign n16349 = ~n16347 & ~n16348;
  assign n16350 = pi121  & n1269;
  assign n16351 = pi119  & n1340;
  assign n16352 = pi120  & n1264;
  assign n16353 = ~n16351 & ~n16352;
  assign n16354 = ~n16350 & n16353;
  assign n16355 = n1272 & n11086;
  assign n16356 = n16354 & ~n16355;
  assign n16357 = pi17  & ~n16356;
  assign n16358 = pi17  & ~n16357;
  assign n16359 = ~n16356 & ~n16357;
  assign n16360 = ~n16358 & ~n16359;
  assign n16361 = ~n16008 & ~n16289;
  assign n16362 = n16360 & n16361;
  assign n16363 = ~n16360 & ~n16361;
  assign n16364 = ~n16362 & ~n16363;
  assign n16365 = pi115  & n2004;
  assign n16366 = pi113  & n2141;
  assign n16367 = pi114  & n1999;
  assign n16368 = ~n16366 & ~n16367;
  assign n16369 = ~n16365 & n16368;
  assign n16370 = n2007 & n8727;
  assign n16371 = n16369 & ~n16370;
  assign n16372 = pi23  & ~n16371;
  assign n16373 = pi23  & ~n16372;
  assign n16374 = ~n16371 & ~n16372;
  assign n16375 = ~n16373 & ~n16374;
  assign n16376 = ~n16023 & ~n16269;
  assign n16377 = ~n16375 & ~n16376;
  assign n16378 = n16375 & n16376;
  assign n16379 = ~n16377 & ~n16378;
  assign n16380 = pi112  & n2486;
  assign n16381 = pi110  & n2644;
  assign n16382 = pi111  & n2481;
  assign n16383 = ~n16381 & ~n16382;
  assign n16384 = ~n16380 & n16383;
  assign n16385 = n2489 & n7795;
  assign n16386 = n16384 & ~n16385;
  assign n16387 = pi26  & ~n16386;
  assign n16388 = pi26  & ~n16387;
  assign n16389 = ~n16386 & ~n16387;
  assign n16390 = ~n16388 & ~n16389;
  assign n16391 = ~n16037 & ~n16264;
  assign n16392 = n16390 & n16391;
  assign n16393 = ~n16390 & ~n16391;
  assign n16394 = ~n16392 & ~n16393;
  assign n16395 = ~n16258 & ~n16261;
  assign n16396 = pi109  & n2976;
  assign n16397 = pi107  & n3182;
  assign n16398 = pi108  & n2971;
  assign n16399 = ~n16397 & ~n16398;
  assign n16400 = ~n16396 & n16399;
  assign n16401 = n2979 & n7170;
  assign n16402 = n16400 & ~n16401;
  assign n16403 = pi29  & ~n16402;
  assign n16404 = pi29  & ~n16403;
  assign n16405 = ~n16402 & ~n16403;
  assign n16406 = ~n16404 & ~n16405;
  assign n16407 = ~n16395 & ~n16406;
  assign n16408 = n16395 & n16406;
  assign n16409 = ~n16407 & ~n16408;
  assign n16410 = ~n16054 & ~n16241;
  assign n16411 = pi106  & n3550;
  assign n16412 = pi104  & n3735;
  assign n16413 = pi105  & n3545;
  assign n16414 = ~n16412 & ~n16413;
  assign n16415 = ~n16411 & n16414;
  assign n16416 = n3553 & n6090;
  assign n16417 = n16415 & ~n16416;
  assign n16418 = pi32  & ~n16417;
  assign n16419 = pi32  & ~n16418;
  assign n16420 = ~n16417 & ~n16418;
  assign n16421 = ~n16419 & ~n16420;
  assign n16422 = ~n16410 & ~n16421;
  assign n16423 = n16410 & n16421;
  assign n16424 = ~n16422 & ~n16423;
  assign n16425 = ~n16205 & ~n16219;
  assign n16426 = pi100  & n4896;
  assign n16427 = pi98  & n5148;
  assign n16428 = pi99  & n4891;
  assign n16429 = ~n16427 & ~n16428;
  assign n16430 = ~n16426 & n16429;
  assign n16431 = n4808 & n4899;
  assign n16432 = n16430 & ~n16431;
  assign n16433 = pi38  & ~n16432;
  assign n16434 = pi38  & ~n16433;
  assign n16435 = ~n16432 & ~n16433;
  assign n16436 = ~n16434 & ~n16435;
  assign n16437 = ~n16188 & ~n16202;
  assign n16438 = ~n16171 & ~n16184;
  assign n16439 = ~n16153 & ~n16167;
  assign n16440 = ~n16147 & ~n16150;
  assign n16441 = pi88  & n8137;
  assign n16442 = pi86  & n8471;
  assign n16443 = pi87  & n8132;
  assign n16444 = ~n16442 & ~n16443;
  assign n16445 = ~n16441 & n16444;
  assign n16446 = n2277 & n8140;
  assign n16447 = n16445 & ~n16446;
  assign n16448 = pi50  & ~n16447;
  assign n16449 = pi50  & ~n16448;
  assign n16450 = ~n16447 & ~n16448;
  assign n16451 = ~n16449 & ~n16450;
  assign n16452 = ~n16114 & ~n16127;
  assign n16453 = ~n16107 & ~n16110;
  assign n16454 = pi76  & n12295;
  assign n16455 = pi74  & n12693;
  assign n16456 = pi75  & n12290;
  assign n16457 = ~n16455 & ~n16456;
  assign n16458 = ~n16454 & n16457;
  assign n16459 = n881 & n12298;
  assign n16460 = n16458 & ~n16459;
  assign n16461 = pi62  & ~n16460;
  assign n16462 = pi62  & ~n16461;
  assign n16463 = ~n16460 & ~n16461;
  assign n16464 = ~n16462 & ~n16463;
  assign n16465 = pi72  & n13477;
  assign n16466 = pi73  & ~n13122;
  assign n16467 = ~n16465 & ~n16466;
  assign n16468 = ~pi8  & ~n16087;
  assign n16469 = pi8  & n16087;
  assign n16470 = ~n16468 & ~n16469;
  assign n16471 = ~n16467 & n16470;
  assign n16472 = n16467 & ~n16470;
  assign n16473 = ~n16471 & ~n16472;
  assign n16474 = ~n16093 & n16473;
  assign n16475 = n16093 & ~n16473;
  assign n16476 = ~n16474 & ~n16475;
  assign n16477 = n16464 & n16476;
  assign n16478 = ~n16464 & ~n16476;
  assign n16479 = ~n16477 & ~n16478;
  assign n16480 = pi79  & n11193;
  assign n16481 = pi77  & n11567;
  assign n16482 = pi78  & n11188;
  assign n16483 = ~n16481 & ~n16482;
  assign n16484 = ~n16480 & n16483;
  assign n16485 = n1105 & n11196;
  assign n16486 = n16484 & ~n16485;
  assign n16487 = pi59  & ~n16486;
  assign n16488 = pi59  & ~n16487;
  assign n16489 = ~n16486 & ~n16487;
  assign n16490 = ~n16488 & ~n16489;
  assign n16491 = ~n16479 & ~n16490;
  assign n16492 = n16479 & n16490;
  assign n16493 = ~n16491 & ~n16492;
  assign n16494 = ~n16453 & n16493;
  assign n16495 = n16453 & ~n16493;
  assign n16496 = ~n16494 & ~n16495;
  assign n16497 = pi82  & n10135;
  assign n16498 = pi80  & n10478;
  assign n16499 = pi81  & n10130;
  assign n16500 = ~n16498 & ~n16499;
  assign n16501 = ~n16497 & n16500;
  assign n16502 = n1532 & n10138;
  assign n16503 = n16501 & ~n16502;
  assign n16504 = pi56  & ~n16503;
  assign n16505 = pi56  & ~n16504;
  assign n16506 = ~n16503 & ~n16504;
  assign n16507 = ~n16505 & ~n16506;
  assign n16508 = n16496 & ~n16507;
  assign n16509 = ~n16496 & n16507;
  assign n16510 = ~n16508 & ~n16509;
  assign n16511 = n16452 & ~n16510;
  assign n16512 = ~n16452 & n16510;
  assign n16513 = ~n16511 & ~n16512;
  assign n16514 = pi85  & n9096;
  assign n16515 = pi83  & n9453;
  assign n16516 = pi84  & n9091;
  assign n16517 = ~n16515 & ~n16516;
  assign n16518 = ~n16514 & n16517;
  assign n16519 = n1943 & n9099;
  assign n16520 = n16518 & ~n16519;
  assign n16521 = pi53  & ~n16520;
  assign n16522 = pi53  & ~n16521;
  assign n16523 = ~n16520 & ~n16521;
  assign n16524 = ~n16522 & ~n16523;
  assign n16525 = n16513 & ~n16524;
  assign n16526 = n16513 & ~n16525;
  assign n16527 = ~n16524 & ~n16525;
  assign n16528 = ~n16526 & ~n16527;
  assign n16529 = ~n16131 & ~n16145;
  assign n16530 = ~n16528 & ~n16529;
  assign n16531 = n16528 & n16529;
  assign n16532 = ~n16530 & ~n16531;
  assign n16533 = ~n16451 & n16532;
  assign n16534 = n16451 & ~n16532;
  assign n16535 = ~n16533 & ~n16534;
  assign n16536 = ~n16440 & n16535;
  assign n16537 = n16440 & ~n16535;
  assign n16538 = ~n16536 & ~n16537;
  assign n16539 = pi91  & n7239;
  assign n16540 = pi89  & n7556;
  assign n16541 = pi90  & n7234;
  assign n16542 = ~n16540 & ~n16541;
  assign n16543 = ~n16539 & n16542;
  assign n16544 = n2926 & n7242;
  assign n16545 = n16543 & ~n16544;
  assign n16546 = pi47  & ~n16545;
  assign n16547 = pi47  & ~n16546;
  assign n16548 = ~n16545 & ~n16546;
  assign n16549 = ~n16547 & ~n16548;
  assign n16550 = n16538 & ~n16549;
  assign n16551 = ~n16538 & n16549;
  assign n16552 = ~n16550 & ~n16551;
  assign n16553 = n16439 & ~n16552;
  assign n16554 = ~n16439 & n16552;
  assign n16555 = ~n16553 & ~n16554;
  assign n16556 = pi94  & n6396;
  assign n16557 = pi92  & n6735;
  assign n16558 = pi93  & n6391;
  assign n16559 = ~n16557 & ~n16558;
  assign n16560 = ~n16556 & n16559;
  assign n16561 = n3499 & n6399;
  assign n16562 = n16560 & ~n16561;
  assign n16563 = pi44  & ~n16562;
  assign n16564 = pi44  & ~n16563;
  assign n16565 = ~n16562 & ~n16563;
  assign n16566 = ~n16564 & ~n16565;
  assign n16567 = n16555 & ~n16566;
  assign n16568 = ~n16555 & n16566;
  assign n16569 = ~n16438 & ~n16568;
  assign n16570 = ~n16567 & n16569;
  assign n16571 = ~n16438 & ~n16570;
  assign n16572 = ~n16567 & ~n16570;
  assign n16573 = ~n16568 & n16572;
  assign n16574 = ~n16571 & ~n16573;
  assign n16575 = pi97  & n5636;
  assign n16576 = pi95  & n5909;
  assign n16577 = pi96  & n5631;
  assign n16578 = ~n16576 & ~n16577;
  assign n16579 = ~n16575 & n16578;
  assign n16580 = n3946 & n5639;
  assign n16581 = n16579 & ~n16580;
  assign n16582 = pi41  & ~n16581;
  assign n16583 = pi41  & ~n16582;
  assign n16584 = ~n16581 & ~n16582;
  assign n16585 = ~n16583 & ~n16584;
  assign n16586 = ~n16574 & ~n16585;
  assign n16587 = n16574 & n16585;
  assign n16588 = ~n16586 & ~n16587;
  assign n16589 = ~n16437 & n16588;
  assign n16590 = n16437 & ~n16588;
  assign n16591 = ~n16589 & ~n16590;
  assign n16592 = ~n16436 & n16591;
  assign n16593 = n16436 & ~n16591;
  assign n16594 = ~n16592 & ~n16593;
  assign n16595 = n16425 & ~n16594;
  assign n16596 = ~n16425 & n16594;
  assign n16597 = ~n16595 & ~n16596;
  assign n16598 = pi103  & n4182;
  assign n16599 = pi101  & n4416;
  assign n16600 = pi102  & n4177;
  assign n16601 = ~n16599 & ~n16600;
  assign n16602 = ~n16598 & n16601;
  assign n16603 = n4185 & n5540;
  assign n16604 = n16602 & ~n16603;
  assign n16605 = pi35  & ~n16604;
  assign n16606 = pi35  & ~n16605;
  assign n16607 = ~n16604 & ~n16605;
  assign n16608 = ~n16606 & ~n16607;
  assign n16609 = n16597 & ~n16608;
  assign n16610 = n16597 & ~n16609;
  assign n16611 = ~n16608 & ~n16609;
  assign n16612 = ~n16610 & ~n16611;
  assign n16613 = ~n16225 & ~n16238;
  assign n16614 = ~n16612 & ~n16613;
  assign n16615 = n16612 & n16613;
  assign n16616 = ~n16614 & ~n16615;
  assign n16617 = n16424 & n16616;
  assign n16618 = ~n16424 & ~n16616;
  assign n16619 = ~n16617 & ~n16618;
  assign n16620 = n16409 & n16619;
  assign n16621 = ~n16409 & ~n16619;
  assign n16622 = ~n16620 & ~n16621;
  assign n16623 = n16394 & n16622;
  assign n16624 = ~n16394 & ~n16622;
  assign n16625 = ~n16623 & ~n16624;
  assign n16626 = n16379 & n16625;
  assign n16627 = ~n16379 & ~n16625;
  assign n16628 = ~n16626 & ~n16627;
  assign n16629 = ~n16283 & ~n16286;
  assign n16630 = pi118  & n1582;
  assign n16631 = pi116  & n1713;
  assign n16632 = pi117  & n1577;
  assign n16633 = ~n16631 & ~n16632;
  assign n16634 = ~n16630 & n16633;
  assign n16635 = n1585 & n9716;
  assign n16636 = n16634 & ~n16635;
  assign n16637 = pi20  & ~n16636;
  assign n16638 = pi20  & ~n16637;
  assign n16639 = ~n16636 & ~n16637;
  assign n16640 = ~n16638 & ~n16639;
  assign n16641 = ~n16629 & ~n16640;
  assign n16642 = n16629 & n16640;
  assign n16643 = ~n16641 & ~n16642;
  assign n16644 = n16628 & n16643;
  assign n16645 = ~n16628 & ~n16643;
  assign n16646 = ~n16644 & ~n16645;
  assign n16647 = n16364 & n16646;
  assign n16648 = ~n16364 & ~n16646;
  assign n16649 = ~n16349 & ~n16648;
  assign n16650 = ~n16647 & n16649;
  assign n16651 = ~n16349 & ~n16650;
  assign n16652 = ~n16648 & ~n16650;
  assign n16653 = ~n16647 & n16652;
  assign n16654 = ~n16651 & ~n16653;
  assign n16655 = ~n15991 & ~n16310;
  assign n16656 = pi127  & n675;
  assign n16657 = pi125  & n769;
  assign n16658 = pi126  & n670;
  assign n16659 = ~n16657 & ~n16658;
  assign n16660 = ~n16656 & n16659;
  assign n16661 = n678 & n13365;
  assign n16662 = n16660 & ~n16661;
  assign n16663 = pi11  & ~n16662;
  assign n16664 = pi11  & ~n16663;
  assign n16665 = ~n16662 & ~n16663;
  assign n16666 = ~n16664 & ~n16665;
  assign n16667 = ~n16655 & ~n16666;
  assign n16668 = n16655 & n16666;
  assign n16669 = ~n16667 & ~n16668;
  assign n16670 = ~n16654 & n16669;
  assign n16671 = n16654 & ~n16669;
  assign n16672 = ~n16670 & ~n16671;
  assign n16673 = ~n16334 & n16672;
  assign n16674 = n16334 & ~n16672;
  assign n16675 = ~n16673 & ~n16674;
  assign n16676 = ~n16333 & n16675;
  assign n16677 = n16333 & ~n16675;
  assign po72  = ~n16676 & ~n16677;
  assign n16679 = ~n16673 & ~n16676;
  assign n16680 = ~n16667 & ~n16670;
  assign n16681 = pi119  & n1582;
  assign n16682 = pi117  & n1713;
  assign n16683 = pi118  & n1577;
  assign n16684 = ~n16682 & ~n16683;
  assign n16685 = ~n16681 & n16684;
  assign n16686 = n1585 & n10048;
  assign n16687 = n16685 & ~n16686;
  assign n16688 = pi20  & ~n16687;
  assign n16689 = pi20  & ~n16688;
  assign n16690 = ~n16687 & ~n16688;
  assign n16691 = ~n16689 & ~n16690;
  assign n16692 = ~n16377 & ~n16626;
  assign n16693 = n16691 & n16692;
  assign n16694 = ~n16691 & ~n16692;
  assign n16695 = ~n16693 & ~n16694;
  assign n16696 = pi116  & n2004;
  assign n16697 = pi114  & n2141;
  assign n16698 = pi115  & n1999;
  assign n16699 = ~n16697 & ~n16698;
  assign n16700 = ~n16696 & n16699;
  assign n16701 = n2007 & n9042;
  assign n16702 = n16700 & ~n16701;
  assign n16703 = pi23  & ~n16702;
  assign n16704 = pi23  & ~n16703;
  assign n16705 = ~n16702 & ~n16703;
  assign n16706 = ~n16704 & ~n16705;
  assign n16707 = ~n16393 & ~n16623;
  assign n16708 = n16706 & n16707;
  assign n16709 = ~n16706 & ~n16707;
  assign n16710 = ~n16708 & ~n16709;
  assign n16711 = pi113  & n2486;
  assign n16712 = pi111  & n2644;
  assign n16713 = pi112  & n2481;
  assign n16714 = ~n16712 & ~n16713;
  assign n16715 = ~n16711 & n16714;
  assign n16716 = n2489 & n8387;
  assign n16717 = n16715 & ~n16716;
  assign n16718 = pi26  & ~n16717;
  assign n16719 = pi26  & ~n16718;
  assign n16720 = ~n16717 & ~n16718;
  assign n16721 = ~n16719 & ~n16720;
  assign n16722 = ~n16407 & ~n16620;
  assign n16723 = ~n16721 & ~n16722;
  assign n16724 = n16721 & n16722;
  assign n16725 = ~n16723 & ~n16724;
  assign n16726 = pi107  & n3550;
  assign n16727 = pi105  & n3735;
  assign n16728 = pi106  & n3545;
  assign n16729 = ~n16727 & ~n16728;
  assign n16730 = ~n16726 & n16729;
  assign n16731 = n3553 & n6614;
  assign n16732 = n16730 & ~n16731;
  assign n16733 = pi32  & ~n16732;
  assign n16734 = pi32  & ~n16733;
  assign n16735 = ~n16732 & ~n16733;
  assign n16736 = ~n16734 & ~n16735;
  assign n16737 = ~n16609 & ~n16614;
  assign n16738 = n16736 & n16737;
  assign n16739 = ~n16736 & ~n16737;
  assign n16740 = ~n16738 & ~n16739;
  assign n16741 = pi104  & n4182;
  assign n16742 = pi102  & n4416;
  assign n16743 = pi103  & n4177;
  assign n16744 = ~n16742 & ~n16743;
  assign n16745 = ~n16741 & n16744;
  assign n16746 = n4185 & n5565;
  assign n16747 = n16745 & ~n16746;
  assign n16748 = pi35  & ~n16747;
  assign n16749 = pi35  & ~n16748;
  assign n16750 = ~n16747 & ~n16748;
  assign n16751 = ~n16749 & ~n16750;
  assign n16752 = ~n16592 & ~n16596;
  assign n16753 = pi101  & n4896;
  assign n16754 = pi99  & n5148;
  assign n16755 = pi100  & n4891;
  assign n16756 = ~n16754 & ~n16755;
  assign n16757 = ~n16753 & n16756;
  assign n16758 = n4899 & n5056;
  assign n16759 = n16757 & ~n16758;
  assign n16760 = pi38  & ~n16759;
  assign n16761 = pi38  & ~n16760;
  assign n16762 = ~n16759 & ~n16760;
  assign n16763 = ~n16761 & ~n16762;
  assign n16764 = ~n16586 & ~n16589;
  assign n16765 = pi98  & n5636;
  assign n16766 = pi96  & n5909;
  assign n16767 = pi97  & n5631;
  assign n16768 = ~n16766 & ~n16767;
  assign n16769 = ~n16765 & n16768;
  assign n16770 = n4360 & n5639;
  assign n16771 = n16769 & ~n16770;
  assign n16772 = pi41  & ~n16771;
  assign n16773 = pi41  & ~n16772;
  assign n16774 = ~n16771 & ~n16772;
  assign n16775 = ~n16773 & ~n16774;
  assign n16776 = ~n16550 & ~n16554;
  assign n16777 = ~n16533 & ~n16536;
  assign n16778 = ~n16525 & ~n16530;
  assign n16779 = ~n16508 & ~n16512;
  assign n16780 = ~n16491 & ~n16494;
  assign n16781 = pi80  & n11193;
  assign n16782 = pi78  & n11567;
  assign n16783 = pi79  & n11188;
  assign n16784 = ~n16782 & ~n16783;
  assign n16785 = ~n16781 & n16784;
  assign n16786 = n1205 & n11196;
  assign n16787 = n16785 & ~n16786;
  assign n16788 = pi59  & ~n16787;
  assign n16789 = pi59  & ~n16788;
  assign n16790 = ~n16787 & ~n16788;
  assign n16791 = ~n16789 & ~n16790;
  assign n16792 = ~n16475 & ~n16477;
  assign n16793 = pi77  & n12295;
  assign n16794 = pi75  & n12693;
  assign n16795 = pi76  & n12290;
  assign n16796 = ~n16794 & ~n16795;
  assign n16797 = ~n16793 & n16796;
  assign n16798 = n984 & n12298;
  assign n16799 = n16797 & ~n16798;
  assign n16800 = pi62  & ~n16799;
  assign n16801 = pi62  & ~n16800;
  assign n16802 = ~n16799 & ~n16800;
  assign n16803 = ~n16801 & ~n16802;
  assign n16804 = pi73  & n13477;
  assign n16805 = pi74  & ~n13122;
  assign n16806 = ~n16804 & ~n16805;
  assign n16807 = ~n16468 & ~n16471;
  assign n16808 = n16806 & ~n16807;
  assign n16809 = ~n16806 & n16807;
  assign n16810 = ~n16808 & ~n16809;
  assign n16811 = ~n16803 & n16810;
  assign n16812 = n16803 & ~n16810;
  assign n16813 = ~n16811 & ~n16812;
  assign n16814 = n16792 & n16813;
  assign n16815 = ~n16792 & ~n16813;
  assign n16816 = ~n16814 & ~n16815;
  assign n16817 = ~n16791 & n16816;
  assign n16818 = n16791 & ~n16816;
  assign n16819 = ~n16817 & ~n16818;
  assign n16820 = n16780 & ~n16819;
  assign n16821 = ~n16780 & n16819;
  assign n16822 = ~n16820 & ~n16821;
  assign n16823 = pi83  & n10135;
  assign n16824 = pi81  & n10478;
  assign n16825 = pi82  & n10130;
  assign n16826 = ~n16824 & ~n16825;
  assign n16827 = ~n16823 & n16826;
  assign n16828 = n1672 & n10138;
  assign n16829 = n16827 & ~n16828;
  assign n16830 = pi56  & ~n16829;
  assign n16831 = pi56  & ~n16830;
  assign n16832 = ~n16829 & ~n16830;
  assign n16833 = ~n16831 & ~n16832;
  assign n16834 = n16822 & ~n16833;
  assign n16835 = ~n16822 & n16833;
  assign n16836 = ~n16834 & ~n16835;
  assign n16837 = n16779 & ~n16836;
  assign n16838 = ~n16779 & n16836;
  assign n16839 = ~n16837 & ~n16838;
  assign n16840 = pi86  & n9096;
  assign n16841 = pi84  & n9453;
  assign n16842 = pi85  & n9091;
  assign n16843 = ~n16841 & ~n16842;
  assign n16844 = ~n16840 & n16843;
  assign n16845 = n2099 & n9099;
  assign n16846 = n16844 & ~n16845;
  assign n16847 = pi53  & ~n16846;
  assign n16848 = pi53  & ~n16847;
  assign n16849 = ~n16846 & ~n16847;
  assign n16850 = ~n16848 & ~n16849;
  assign n16851 = n16839 & ~n16850;
  assign n16852 = ~n16839 & n16850;
  assign n16853 = ~n16851 & ~n16852;
  assign n16854 = n16778 & ~n16853;
  assign n16855 = ~n16778 & n16853;
  assign n16856 = ~n16854 & ~n16855;
  assign n16857 = pi89  & n8137;
  assign n16858 = pi87  & n8471;
  assign n16859 = pi88  & n8132;
  assign n16860 = ~n16858 & ~n16859;
  assign n16861 = ~n16857 & n16860;
  assign n16862 = n2432 & n8140;
  assign n16863 = n16861 & ~n16862;
  assign n16864 = pi50  & ~n16863;
  assign n16865 = pi50  & ~n16864;
  assign n16866 = ~n16863 & ~n16864;
  assign n16867 = ~n16865 & ~n16866;
  assign n16868 = n16856 & ~n16867;
  assign n16869 = ~n16856 & n16867;
  assign n16870 = ~n16868 & ~n16869;
  assign n16871 = n16777 & ~n16870;
  assign n16872 = ~n16777 & n16870;
  assign n16873 = ~n16871 & ~n16872;
  assign n16874 = pi92  & n7239;
  assign n16875 = pi90  & n7556;
  assign n16876 = pi91  & n7234;
  assign n16877 = ~n16875 & ~n16876;
  assign n16878 = ~n16874 & n16877;
  assign n16879 = n3119 & n7242;
  assign n16880 = n16878 & ~n16879;
  assign n16881 = pi47  & ~n16880;
  assign n16882 = pi47  & ~n16881;
  assign n16883 = ~n16880 & ~n16881;
  assign n16884 = ~n16882 & ~n16883;
  assign n16885 = n16873 & ~n16884;
  assign n16886 = ~n16873 & n16884;
  assign n16887 = ~n16885 & ~n16886;
  assign n16888 = n16776 & ~n16887;
  assign n16889 = ~n16776 & n16887;
  assign n16890 = ~n16888 & ~n16889;
  assign n16891 = pi95  & n6396;
  assign n16892 = pi93  & n6735;
  assign n16893 = pi94  & n6391;
  assign n16894 = ~n16892 & ~n16893;
  assign n16895 = ~n16891 & n16894;
  assign n16896 = n3710 & n6399;
  assign n16897 = n16895 & ~n16896;
  assign n16898 = pi44  & ~n16897;
  assign n16899 = pi44  & ~n16898;
  assign n16900 = ~n16897 & ~n16898;
  assign n16901 = ~n16899 & ~n16900;
  assign n16902 = ~n16890 & n16901;
  assign n16903 = n16890 & ~n16901;
  assign n16904 = ~n16902 & ~n16903;
  assign n16905 = ~n16572 & n16904;
  assign n16906 = n16572 & ~n16904;
  assign n16907 = ~n16905 & ~n16906;
  assign n16908 = ~n16775 & n16907;
  assign n16909 = n16775 & ~n16907;
  assign n16910 = ~n16908 & ~n16909;
  assign n16911 = ~n16764 & n16910;
  assign n16912 = n16764 & ~n16910;
  assign n16913 = ~n16911 & ~n16912;
  assign n16914 = ~n16763 & n16913;
  assign n16915 = n16763 & ~n16913;
  assign n16916 = ~n16914 & ~n16915;
  assign n16917 = ~n16752 & n16916;
  assign n16918 = n16752 & ~n16916;
  assign n16919 = ~n16917 & ~n16918;
  assign n16920 = ~n16751 & n16919;
  assign n16921 = n16751 & ~n16919;
  assign n16922 = ~n16920 & ~n16921;
  assign n16923 = n16740 & n16922;
  assign n16924 = ~n16740 & ~n16922;
  assign n16925 = ~n16923 & ~n16924;
  assign n16926 = ~n16422 & ~n16617;
  assign n16927 = pi110  & n2976;
  assign n16928 = pi108  & n3182;
  assign n16929 = pi109  & n2971;
  assign n16930 = ~n16928 & ~n16929;
  assign n16931 = ~n16927 & n16930;
  assign n16932 = ~n2979 & n16931;
  assign n16933 = ~n7474 & n16931;
  assign n16934 = ~n16932 & ~n16933;
  assign n16935 = pi29  & ~n16934;
  assign n16936 = ~pi29  & n16934;
  assign n16937 = ~n16935 & ~n16936;
  assign n16938 = ~n16926 & ~n16937;
  assign n16939 = n16926 & n16937;
  assign n16940 = ~n16938 & ~n16939;
  assign n16941 = n16925 & n16940;
  assign n16942 = ~n16925 & ~n16940;
  assign n16943 = ~n16941 & ~n16942;
  assign n16944 = n16725 & n16943;
  assign n16945 = ~n16725 & ~n16943;
  assign n16946 = ~n16944 & ~n16945;
  assign n16947 = n16710 & n16946;
  assign n16948 = ~n16710 & ~n16946;
  assign n16949 = n16695 & ~n16948;
  assign n16950 = ~n16947 & n16949;
  assign n16951 = n16695 & ~n16950;
  assign n16952 = ~n16948 & ~n16950;
  assign n16953 = ~n16947 & n16952;
  assign n16954 = ~n16951 & ~n16953;
  assign n16955 = ~n16641 & ~n16644;
  assign n16956 = pi122  & n1269;
  assign n16957 = pi120  & n1340;
  assign n16958 = pi121  & n1264;
  assign n16959 = ~n16957 & ~n16958;
  assign n16960 = ~n16956 & n16959;
  assign n16961 = ~n1272 & n16960;
  assign n16962 = ~n11463 & n16960;
  assign n16963 = ~n16961 & ~n16962;
  assign n16964 = pi17  & ~n16963;
  assign n16965 = ~pi17  & n16963;
  assign n16966 = ~n16964 & ~n16965;
  assign n16967 = ~n16955 & ~n16966;
  assign n16968 = n16955 & n16966;
  assign n16969 = ~n16967 & ~n16968;
  assign n16970 = ~n16954 & n16969;
  assign n16971 = ~n16954 & ~n16970;
  assign n16972 = n16969 & ~n16970;
  assign n16973 = ~n16971 & ~n16972;
  assign n16974 = pi125  & n918;
  assign n16975 = pi123  & n1031;
  assign n16976 = pi124  & n913;
  assign n16977 = ~n16975 & ~n16976;
  assign n16978 = ~n16974 & n16977;
  assign n16979 = n921 & n12591;
  assign n16980 = n16978 & ~n16979;
  assign n16981 = pi14  & ~n16980;
  assign n16982 = pi14  & ~n16981;
  assign n16983 = ~n16980 & ~n16981;
  assign n16984 = ~n16982 & ~n16983;
  assign n16985 = ~n16363 & ~n16647;
  assign n16986 = ~n16984 & ~n16985;
  assign n16987 = n16984 & n16985;
  assign n16988 = ~n16986 & ~n16987;
  assign n16989 = ~n16973 & n16988;
  assign n16990 = n16973 & ~n16988;
  assign n16991 = ~n16989 & ~n16990;
  assign n16992 = ~n16335 & ~n16346;
  assign n16993 = ~n16650 & ~n16992;
  assign n16994 = pi126  & n769;
  assign n16995 = pi127  & n670;
  assign n16996 = ~n16994 & ~n16995;
  assign n16997 = ~n678 & n16996;
  assign n16998 = ~n13389 & n16996;
  assign n16999 = ~n16997 & ~n16998;
  assign n17000 = pi11  & ~n16999;
  assign n17001 = ~pi11  & n16999;
  assign n17002 = ~n17000 & ~n17001;
  assign n17003 = ~n16993 & ~n17002;
  assign n17004 = n16993 & n17002;
  assign n17005 = ~n17003 & ~n17004;
  assign n17006 = n16991 & n17005;
  assign n17007 = ~n16991 & ~n17005;
  assign n17008 = ~n17006 & ~n17007;
  assign n17009 = ~n16680 & n17008;
  assign n17010 = n16680 & ~n17008;
  assign n17011 = ~n17009 & ~n17010;
  assign n17012 = ~n16679 & n17011;
  assign n17013 = n16679 & ~n17011;
  assign po73  = ~n17012 & ~n17013;
  assign n17015 = ~n17009 & ~n17012;
  assign n17016 = ~n17003 & ~n17006;
  assign n17017 = ~n16967 & ~n16970;
  assign n17018 = pi126  & n918;
  assign n17019 = pi124  & n1031;
  assign n17020 = pi125  & n913;
  assign n17021 = ~n17019 & ~n17020;
  assign n17022 = ~n17018 & n17021;
  assign n17023 = ~n921 & n17022;
  assign n17024 = ~n12979 & n17022;
  assign n17025 = ~n17023 & ~n17024;
  assign n17026 = pi14  & ~n17025;
  assign n17027 = ~pi14  & n17025;
  assign n17028 = ~n17026 & ~n17027;
  assign n17029 = ~n17017 & ~n17028;
  assign n17030 = n17017 & n17028;
  assign n17031 = ~n17029 & ~n17030;
  assign n17032 = pi123  & n1269;
  assign n17033 = pi121  & n1340;
  assign n17034 = pi122  & n1264;
  assign n17035 = ~n17033 & ~n17034;
  assign n17036 = ~n17032 & n17035;
  assign n17037 = n1272 & n11489;
  assign n17038 = n17036 & ~n17037;
  assign n17039 = pi17  & ~n17038;
  assign n17040 = pi17  & ~n17039;
  assign n17041 = ~n17038 & ~n17039;
  assign n17042 = ~n17040 & ~n17041;
  assign n17043 = ~n16694 & ~n16950;
  assign n17044 = n17042 & n17043;
  assign n17045 = ~n17042 & ~n17043;
  assign n17046 = ~n17044 & ~n17045;
  assign n17047 = pi120  & n1582;
  assign n17048 = pi118  & n1713;
  assign n17049 = pi119  & n1577;
  assign n17050 = ~n17048 & ~n17049;
  assign n17051 = ~n17047 & n17050;
  assign n17052 = n1585 & n10734;
  assign n17053 = n17051 & ~n17052;
  assign n17054 = pi20  & ~n17053;
  assign n17055 = pi20  & ~n17054;
  assign n17056 = ~n17053 & ~n17054;
  assign n17057 = ~n17055 & ~n17056;
  assign n17058 = ~n16709 & ~n16947;
  assign n17059 = ~n17057 & ~n17058;
  assign n17060 = n17057 & n17058;
  assign n17061 = ~n17059 & ~n17060;
  assign n17062 = ~n16938 & ~n16941;
  assign n17063 = pi114  & n2486;
  assign n17064 = pi112  & n2644;
  assign n17065 = pi113  & n2481;
  assign n17066 = ~n17064 & ~n17065;
  assign n17067 = ~n17063 & n17066;
  assign n17068 = ~n2489 & n17067;
  assign n17069 = ~n8702 & n17067;
  assign n17070 = ~n17068 & ~n17069;
  assign n17071 = pi26  & ~n17070;
  assign n17072 = ~pi26  & n17070;
  assign n17073 = ~n17071 & ~n17072;
  assign n17074 = ~n17062 & ~n17073;
  assign n17075 = n17062 & n17073;
  assign n17076 = ~n17074 & ~n17075;
  assign n17077 = pi111  & n2976;
  assign n17078 = pi109  & n3182;
  assign n17079 = pi110  & n2971;
  assign n17080 = ~n17078 & ~n17079;
  assign n17081 = ~n17077 & n17080;
  assign n17082 = n2979 & n7770;
  assign n17083 = n17081 & ~n17082;
  assign n17084 = pi29  & ~n17083;
  assign n17085 = pi29  & ~n17084;
  assign n17086 = ~n17083 & ~n17084;
  assign n17087 = ~n17085 & ~n17086;
  assign n17088 = ~n16739 & ~n16923;
  assign n17089 = n17087 & n17088;
  assign n17090 = ~n17087 & ~n17088;
  assign n17091 = ~n17089 & ~n17090;
  assign n17092 = ~n16917 & ~n16920;
  assign n17093 = pi108  & n3550;
  assign n17094 = pi106  & n3735;
  assign n17095 = pi107  & n3545;
  assign n17096 = ~n17094 & ~n17095;
  assign n17097 = ~n17093 & n17096;
  assign n17098 = ~n3553 & n17097;
  assign n17099 = ~n6639 & n17097;
  assign n17100 = ~n17098 & ~n17099;
  assign n17101 = pi32  & ~n17100;
  assign n17102 = ~pi32  & n17100;
  assign n17103 = ~n17101 & ~n17102;
  assign n17104 = ~n17092 & ~n17103;
  assign n17105 = n17092 & n17103;
  assign n17106 = ~n17104 & ~n17105;
  assign n17107 = pi105  & n4182;
  assign n17108 = pi103  & n4416;
  assign n17109 = pi104  & n4177;
  assign n17110 = ~n17108 & ~n17109;
  assign n17111 = ~n17107 & n17110;
  assign n17112 = n4185 & n6065;
  assign n17113 = n17111 & ~n17112;
  assign n17114 = pi35  & ~n17113;
  assign n17115 = pi35  & ~n17114;
  assign n17116 = ~n17113 & ~n17114;
  assign n17117 = ~n17115 & ~n17116;
  assign n17118 = ~n16911 & ~n16914;
  assign n17119 = ~n16905 & ~n16908;
  assign n17120 = ~n16855 & ~n16868;
  assign n17121 = pi90  & n8137;
  assign n17122 = pi88  & n8471;
  assign n17123 = pi89  & n8132;
  assign n17124 = ~n17122 & ~n17123;
  assign n17125 = ~n17121 & n17124;
  assign n17126 = n2606 & n8140;
  assign n17127 = n17125 & ~n17126;
  assign n17128 = pi50  & ~n17127;
  assign n17129 = pi50  & ~n17128;
  assign n17130 = ~n17127 & ~n17128;
  assign n17131 = ~n17129 & ~n17130;
  assign n17132 = ~n16838 & ~n16851;
  assign n17133 = pi87  & n9096;
  assign n17134 = pi85  & n9453;
  assign n17135 = pi86  & n9091;
  assign n17136 = ~n17134 & ~n17135;
  assign n17137 = ~n17133 & n17136;
  assign n17138 = n2252 & n9099;
  assign n17139 = n17137 & ~n17138;
  assign n17140 = pi53  & ~n17139;
  assign n17141 = pi53  & ~n17140;
  assign n17142 = ~n17139 & ~n17140;
  assign n17143 = ~n17141 & ~n17142;
  assign n17144 = ~n16821 & ~n16834;
  assign n17145 = ~n16814 & ~n16817;
  assign n17146 = ~n16808 & ~n16811;
  assign n17147 = pi74  & n13477;
  assign n17148 = pi75  & ~n13122;
  assign n17149 = ~n17147 & ~n17148;
  assign n17150 = n16806 & ~n17149;
  assign n17151 = ~n16806 & n17149;
  assign n17152 = ~n17150 & ~n17151;
  assign n17153 = ~n17146 & n17152;
  assign n17154 = n17146 & ~n17152;
  assign n17155 = ~n17153 & ~n17154;
  assign n17156 = pi78  & n12295;
  assign n17157 = pi76  & n12693;
  assign n17158 = pi77  & n12290;
  assign n17159 = ~n17157 & ~n17158;
  assign n17160 = ~n17156 & n17159;
  assign n17161 = n1009 & n12298;
  assign n17162 = n17160 & ~n17161;
  assign n17163 = pi62  & ~n17162;
  assign n17164 = pi62  & ~n17163;
  assign n17165 = ~n17162 & ~n17163;
  assign n17166 = ~n17164 & ~n17165;
  assign n17167 = n17155 & ~n17166;
  assign n17168 = n17155 & ~n17167;
  assign n17169 = ~n17166 & ~n17167;
  assign n17170 = ~n17168 & ~n17169;
  assign n17171 = pi81  & n11193;
  assign n17172 = pi79  & n11567;
  assign n17173 = pi80  & n11188;
  assign n17174 = ~n17172 & ~n17173;
  assign n17175 = ~n17171 & n17174;
  assign n17176 = n1413 & n11196;
  assign n17177 = n17175 & ~n17176;
  assign n17178 = pi59  & ~n17177;
  assign n17179 = pi59  & ~n17178;
  assign n17180 = ~n17177 & ~n17178;
  assign n17181 = ~n17179 & ~n17180;
  assign n17182 = ~n17170 & ~n17181;
  assign n17183 = n17170 & n17181;
  assign n17184 = ~n17182 & ~n17183;
  assign n17185 = n17145 & ~n17184;
  assign n17186 = ~n17145 & n17184;
  assign n17187 = ~n17185 & ~n17186;
  assign n17188 = pi84  & n10135;
  assign n17189 = pi82  & n10478;
  assign n17190 = pi83  & n10130;
  assign n17191 = ~n17189 & ~n17190;
  assign n17192 = ~n17188 & n17191;
  assign n17193 = n1805 & n10138;
  assign n17194 = n17192 & ~n17193;
  assign n17195 = pi56  & ~n17194;
  assign n17196 = pi56  & ~n17195;
  assign n17197 = ~n17194 & ~n17195;
  assign n17198 = ~n17196 & ~n17197;
  assign n17199 = ~n17187 & n17198;
  assign n17200 = n17187 & ~n17198;
  assign n17201 = ~n17199 & ~n17200;
  assign n17202 = ~n17144 & n17201;
  assign n17203 = n17144 & ~n17201;
  assign n17204 = ~n17202 & ~n17203;
  assign n17205 = ~n17143 & n17204;
  assign n17206 = n17143 & ~n17204;
  assign n17207 = ~n17205 & ~n17206;
  assign n17208 = ~n17132 & n17207;
  assign n17209 = n17132 & ~n17207;
  assign n17210 = ~n17208 & ~n17209;
  assign n17211 = ~n17131 & n17210;
  assign n17212 = n17131 & ~n17210;
  assign n17213 = ~n17211 & ~n17212;
  assign n17214 = ~n17120 & n17213;
  assign n17215 = n17120 & ~n17213;
  assign n17216 = ~n17214 & ~n17215;
  assign n17217 = pi93  & n7239;
  assign n17218 = pi91  & n7556;
  assign n17219 = pi92  & n7234;
  assign n17220 = ~n17218 & ~n17219;
  assign n17221 = ~n17217 & n17220;
  assign n17222 = n3144 & n7242;
  assign n17223 = n17221 & ~n17222;
  assign n17224 = pi47  & ~n17223;
  assign n17225 = pi47  & ~n17224;
  assign n17226 = ~n17223 & ~n17224;
  assign n17227 = ~n17225 & ~n17226;
  assign n17228 = n17216 & ~n17227;
  assign n17229 = n17216 & ~n17228;
  assign n17230 = ~n17227 & ~n17228;
  assign n17231 = ~n17229 & ~n17230;
  assign n17232 = ~n16872 & ~n16885;
  assign n17233 = n17231 & n17232;
  assign n17234 = ~n17231 & ~n17232;
  assign n17235 = ~n17233 & ~n17234;
  assign n17236 = pi96  & n6396;
  assign n17237 = pi94  & n6735;
  assign n17238 = pi95  & n6391;
  assign n17239 = ~n17237 & ~n17238;
  assign n17240 = ~n17236 & n17239;
  assign n17241 = n3921 & n6399;
  assign n17242 = n17240 & ~n17241;
  assign n17243 = pi44  & ~n17242;
  assign n17244 = pi44  & ~n17243;
  assign n17245 = ~n17242 & ~n17243;
  assign n17246 = ~n17244 & ~n17245;
  assign n17247 = ~n17235 & n17246;
  assign n17248 = n17235 & ~n17246;
  assign n17249 = ~n17247 & ~n17248;
  assign n17250 = ~n16889 & ~n16903;
  assign n17251 = n17249 & ~n17250;
  assign n17252 = ~n17249 & n17250;
  assign n17253 = ~n17251 & ~n17252;
  assign n17254 = pi99  & n5636;
  assign n17255 = pi97  & n5909;
  assign n17256 = pi98  & n5631;
  assign n17257 = ~n17255 & ~n17256;
  assign n17258 = ~n17254 & n17257;
  assign n17259 = n4584 & n5639;
  assign n17260 = n17258 & ~n17259;
  assign n17261 = pi41  & ~n17260;
  assign n17262 = pi41  & ~n17261;
  assign n17263 = ~n17260 & ~n17261;
  assign n17264 = ~n17262 & ~n17263;
  assign n17265 = n17253 & ~n17264;
  assign n17266 = ~n17253 & n17264;
  assign n17267 = ~n17265 & ~n17266;
  assign n17268 = n17119 & ~n17267;
  assign n17269 = ~n17119 & n17267;
  assign n17270 = ~n17268 & ~n17269;
  assign n17271 = pi102  & n4896;
  assign n17272 = pi100  & n5148;
  assign n17273 = pi101  & n4891;
  assign n17274 = ~n17272 & ~n17273;
  assign n17275 = ~n17271 & n17274;
  assign n17276 = n4899 & n5296;
  assign n17277 = n17275 & ~n17276;
  assign n17278 = pi38  & ~n17277;
  assign n17279 = pi38  & ~n17278;
  assign n17280 = ~n17277 & ~n17278;
  assign n17281 = ~n17279 & ~n17280;
  assign n17282 = ~n17270 & n17281;
  assign n17283 = n17270 & ~n17281;
  assign n17284 = ~n17282 & ~n17283;
  assign n17285 = ~n17118 & n17284;
  assign n17286 = n17118 & ~n17284;
  assign n17287 = ~n17285 & ~n17286;
  assign n17288 = ~n17117 & n17287;
  assign n17289 = n17117 & ~n17287;
  assign n17290 = ~n17288 & ~n17289;
  assign n17291 = n17106 & n17290;
  assign n17292 = ~n17106 & ~n17290;
  assign n17293 = ~n17291 & ~n17292;
  assign n17294 = n17091 & n17293;
  assign n17295 = ~n17091 & ~n17293;
  assign n17296 = n17076 & ~n17295;
  assign n17297 = ~n17294 & n17296;
  assign n17298 = n17076 & ~n17297;
  assign n17299 = ~n17295 & ~n17297;
  assign n17300 = ~n17294 & n17299;
  assign n17301 = ~n17298 & ~n17300;
  assign n17302 = ~n16723 & ~n16944;
  assign n17303 = pi117  & n2004;
  assign n17304 = pi115  & n2141;
  assign n17305 = pi116  & n1999;
  assign n17306 = ~n17304 & ~n17305;
  assign n17307 = ~n17303 & n17306;
  assign n17308 = ~n2007 & n17307;
  assign n17309 = ~n9691 & n17307;
  assign n17310 = ~n17308 & ~n17309;
  assign n17311 = pi23  & ~n17310;
  assign n17312 = ~pi23  & n17310;
  assign n17313 = ~n17311 & ~n17312;
  assign n17314 = ~n17302 & ~n17313;
  assign n17315 = n17302 & n17313;
  assign n17316 = ~n17314 & ~n17315;
  assign n17317 = ~n17301 & n17316;
  assign n17318 = n17301 & ~n17316;
  assign n17319 = ~n17317 & ~n17318;
  assign n17320 = n17061 & n17319;
  assign n17321 = ~n17061 & ~n17319;
  assign n17322 = ~n17320 & ~n17321;
  assign n17323 = n17046 & n17322;
  assign n17324 = ~n17046 & ~n17322;
  assign n17325 = n17031 & ~n17324;
  assign n17326 = ~n17323 & n17325;
  assign n17327 = n17031 & ~n17326;
  assign n17328 = ~n17324 & ~n17326;
  assign n17329 = ~n17323 & n17328;
  assign n17330 = ~n17327 & ~n17329;
  assign n17331 = ~n16986 & ~n16989;
  assign n17332 = pi127  & n769;
  assign n17333 = n678 & n13387;
  assign n17334 = ~n17332 & ~n17333;
  assign n17335 = pi11  & ~n17334;
  assign n17336 = pi11  & ~n17335;
  assign n17337 = ~n17334 & ~n17335;
  assign n17338 = ~n17336 & ~n17337;
  assign n17339 = ~n17331 & ~n17338;
  assign n17340 = n17331 & n17338;
  assign n17341 = ~n17339 & ~n17340;
  assign n17342 = n17330 & n17341;
  assign n17343 = ~n17330 & ~n17341;
  assign n17344 = ~n17342 & ~n17343;
  assign n17345 = ~n17016 & ~n17344;
  assign n17346 = n17016 & n17344;
  assign n17347 = ~n17345 & ~n17346;
  assign n17348 = ~n17015 & n17347;
  assign n17349 = n17015 & ~n17347;
  assign po74  = ~n17348 & ~n17349;
  assign n17351 = ~n17345 & ~n17348;
  assign n17352 = ~n17340 & ~n17342;
  assign n17353 = pi121  & n1582;
  assign n17354 = pi119  & n1713;
  assign n17355 = pi120  & n1577;
  assign n17356 = ~n17354 & ~n17355;
  assign n17357 = ~n17353 & n17356;
  assign n17358 = n1585 & n11086;
  assign n17359 = n17357 & ~n17358;
  assign n17360 = pi20  & ~n17359;
  assign n17361 = pi20  & ~n17360;
  assign n17362 = ~n17359 & ~n17360;
  assign n17363 = ~n17361 & ~n17362;
  assign n17364 = ~n17059 & ~n17320;
  assign n17365 = n17363 & n17364;
  assign n17366 = ~n17363 & ~n17364;
  assign n17367 = ~n17365 & ~n17366;
  assign n17368 = ~n17314 & ~n17317;
  assign n17369 = pi118  & n2004;
  assign n17370 = pi116  & n2141;
  assign n17371 = pi117  & n1999;
  assign n17372 = ~n17370 & ~n17371;
  assign n17373 = ~n17369 & n17372;
  assign n17374 = n2007 & n9716;
  assign n17375 = n17373 & ~n17374;
  assign n17376 = pi23  & ~n17375;
  assign n17377 = pi23  & ~n17376;
  assign n17378 = ~n17375 & ~n17376;
  assign n17379 = ~n17377 & ~n17378;
  assign n17380 = ~n17368 & ~n17379;
  assign n17381 = ~n17368 & ~n17380;
  assign n17382 = ~n17379 & ~n17380;
  assign n17383 = ~n17381 & ~n17382;
  assign n17384 = pi115  & n2486;
  assign n17385 = pi113  & n2644;
  assign n17386 = pi114  & n2481;
  assign n17387 = ~n17385 & ~n17386;
  assign n17388 = ~n17384 & n17387;
  assign n17389 = n2489 & n8727;
  assign n17390 = n17388 & ~n17389;
  assign n17391 = pi26  & ~n17390;
  assign n17392 = pi26  & ~n17391;
  assign n17393 = ~n17390 & ~n17391;
  assign n17394 = ~n17392 & ~n17393;
  assign n17395 = ~n17074 & ~n17297;
  assign n17396 = n17394 & n17395;
  assign n17397 = ~n17394 & ~n17395;
  assign n17398 = ~n17396 & ~n17397;
  assign n17399 = ~n17285 & ~n17288;
  assign n17400 = pi106  & n4182;
  assign n17401 = pi104  & n4416;
  assign n17402 = pi105  & n4177;
  assign n17403 = ~n17401 & ~n17402;
  assign n17404 = ~n17400 & n17403;
  assign n17405 = n4185 & n6090;
  assign n17406 = n17404 & ~n17405;
  assign n17407 = pi35  & ~n17406;
  assign n17408 = pi35  & ~n17407;
  assign n17409 = ~n17406 & ~n17407;
  assign n17410 = ~n17408 & ~n17409;
  assign n17411 = ~n17269 & ~n17283;
  assign n17412 = ~n17251 & ~n17265;
  assign n17413 = pi100  & n5636;
  assign n17414 = pi98  & n5909;
  assign n17415 = pi99  & n5631;
  assign n17416 = ~n17414 & ~n17415;
  assign n17417 = ~n17413 & n17416;
  assign n17418 = n4808 & n5639;
  assign n17419 = n17417 & ~n17418;
  assign n17420 = pi41  & ~n17419;
  assign n17421 = pi41  & ~n17420;
  assign n17422 = ~n17419 & ~n17420;
  assign n17423 = ~n17421 & ~n17422;
  assign n17424 = ~n17234 & ~n17248;
  assign n17425 = ~n17214 & ~n17228;
  assign n17426 = ~n17208 & ~n17211;
  assign n17427 = ~n17202 & ~n17205;
  assign n17428 = pi88  & n9096;
  assign n17429 = pi86  & n9453;
  assign n17430 = pi87  & n9091;
  assign n17431 = ~n17429 & ~n17430;
  assign n17432 = ~n17428 & n17431;
  assign n17433 = n2277 & n9099;
  assign n17434 = n17432 & ~n17433;
  assign n17435 = pi53  & ~n17434;
  assign n17436 = pi53  & ~n17435;
  assign n17437 = ~n17434 & ~n17435;
  assign n17438 = ~n17436 & ~n17437;
  assign n17439 = ~n17186 & ~n17200;
  assign n17440 = ~n17150 & ~n17153;
  assign n17441 = pi79  & n12295;
  assign n17442 = pi77  & n12693;
  assign n17443 = pi78  & n12290;
  assign n17444 = ~n17442 & ~n17443;
  assign n17445 = ~n17441 & n17444;
  assign n17446 = n1105 & n12298;
  assign n17447 = n17445 & ~n17446;
  assign n17448 = pi62  & ~n17447;
  assign n17449 = pi62  & ~n17448;
  assign n17450 = ~n17447 & ~n17448;
  assign n17451 = ~n17449 & ~n17450;
  assign n17452 = pi75  & n13477;
  assign n17453 = pi76  & ~n13122;
  assign n17454 = ~n17452 & ~n17453;
  assign n17455 = ~pi11  & ~n16806;
  assign n17456 = pi11  & n16806;
  assign n17457 = ~n17455 & ~n17456;
  assign n17458 = ~n17454 & n17457;
  assign n17459 = n17454 & ~n17457;
  assign n17460 = ~n17458 & ~n17459;
  assign n17461 = ~n17451 & n17460;
  assign n17462 = n17451 & ~n17460;
  assign n17463 = ~n17461 & ~n17462;
  assign n17464 = ~n17440 & n17463;
  assign n17465 = n17440 & ~n17463;
  assign n17466 = ~n17464 & ~n17465;
  assign n17467 = pi82  & n11193;
  assign n17468 = pi80  & n11567;
  assign n17469 = pi81  & n11188;
  assign n17470 = ~n17468 & ~n17469;
  assign n17471 = ~n17467 & n17470;
  assign n17472 = n1532 & n11196;
  assign n17473 = n17471 & ~n17472;
  assign n17474 = pi59  & ~n17473;
  assign n17475 = pi59  & ~n17474;
  assign n17476 = ~n17473 & ~n17474;
  assign n17477 = ~n17475 & ~n17476;
  assign n17478 = n17466 & ~n17477;
  assign n17479 = n17466 & ~n17478;
  assign n17480 = ~n17477 & ~n17478;
  assign n17481 = ~n17479 & ~n17480;
  assign n17482 = ~n17167 & ~n17182;
  assign n17483 = n17481 & n17482;
  assign n17484 = ~n17481 & ~n17482;
  assign n17485 = ~n17483 & ~n17484;
  assign n17486 = pi85  & n10135;
  assign n17487 = pi83  & n10478;
  assign n17488 = pi84  & n10130;
  assign n17489 = ~n17487 & ~n17488;
  assign n17490 = ~n17486 & n17489;
  assign n17491 = n1943 & n10138;
  assign n17492 = n17490 & ~n17491;
  assign n17493 = pi56  & ~n17492;
  assign n17494 = pi56  & ~n17493;
  assign n17495 = ~n17492 & ~n17493;
  assign n17496 = ~n17494 & ~n17495;
  assign n17497 = n17485 & ~n17496;
  assign n17498 = ~n17485 & n17496;
  assign n17499 = ~n17497 & ~n17498;
  assign n17500 = ~n17439 & n17499;
  assign n17501 = n17439 & ~n17499;
  assign n17502 = ~n17500 & ~n17501;
  assign n17503 = ~n17438 & n17502;
  assign n17504 = n17438 & ~n17502;
  assign n17505 = ~n17503 & ~n17504;
  assign n17506 = ~n17427 & n17505;
  assign n17507 = n17427 & ~n17505;
  assign n17508 = ~n17506 & ~n17507;
  assign n17509 = pi91  & n8137;
  assign n17510 = pi89  & n8471;
  assign n17511 = pi90  & n8132;
  assign n17512 = ~n17510 & ~n17511;
  assign n17513 = ~n17509 & n17512;
  assign n17514 = n2926 & n8140;
  assign n17515 = n17513 & ~n17514;
  assign n17516 = pi50  & ~n17515;
  assign n17517 = pi50  & ~n17516;
  assign n17518 = ~n17515 & ~n17516;
  assign n17519 = ~n17517 & ~n17518;
  assign n17520 = n17508 & ~n17519;
  assign n17521 = ~n17508 & n17519;
  assign n17522 = ~n17520 & ~n17521;
  assign n17523 = n17426 & ~n17522;
  assign n17524 = ~n17426 & n17522;
  assign n17525 = ~n17523 & ~n17524;
  assign n17526 = pi94  & n7239;
  assign n17527 = pi92  & n7556;
  assign n17528 = pi93  & n7234;
  assign n17529 = ~n17527 & ~n17528;
  assign n17530 = ~n17526 & n17529;
  assign n17531 = n3499 & n7242;
  assign n17532 = n17530 & ~n17531;
  assign n17533 = pi47  & ~n17532;
  assign n17534 = pi47  & ~n17533;
  assign n17535 = ~n17532 & ~n17533;
  assign n17536 = ~n17534 & ~n17535;
  assign n17537 = n17525 & ~n17536;
  assign n17538 = ~n17525 & n17536;
  assign n17539 = ~n17425 & ~n17538;
  assign n17540 = ~n17537 & n17539;
  assign n17541 = ~n17425 & ~n17540;
  assign n17542 = ~n17537 & ~n17540;
  assign n17543 = ~n17538 & n17542;
  assign n17544 = ~n17541 & ~n17543;
  assign n17545 = pi97  & n6396;
  assign n17546 = pi95  & n6735;
  assign n17547 = pi96  & n6391;
  assign n17548 = ~n17546 & ~n17547;
  assign n17549 = ~n17545 & n17548;
  assign n17550 = n3946 & n6399;
  assign n17551 = n17549 & ~n17550;
  assign n17552 = pi44  & ~n17551;
  assign n17553 = pi44  & ~n17552;
  assign n17554 = ~n17551 & ~n17552;
  assign n17555 = ~n17553 & ~n17554;
  assign n17556 = ~n17544 & ~n17555;
  assign n17557 = n17544 & n17555;
  assign n17558 = ~n17556 & ~n17557;
  assign n17559 = ~n17424 & n17558;
  assign n17560 = n17424 & ~n17558;
  assign n17561 = ~n17559 & ~n17560;
  assign n17562 = ~n17423 & n17561;
  assign n17563 = n17423 & ~n17561;
  assign n17564 = ~n17562 & ~n17563;
  assign n17565 = n17412 & ~n17564;
  assign n17566 = ~n17412 & n17564;
  assign n17567 = ~n17565 & ~n17566;
  assign n17568 = pi103  & n4896;
  assign n17569 = pi101  & n5148;
  assign n17570 = pi102  & n4891;
  assign n17571 = ~n17569 & ~n17570;
  assign n17572 = ~n17568 & n17571;
  assign n17573 = n4899 & n5540;
  assign n17574 = n17572 & ~n17573;
  assign n17575 = pi38  & ~n17574;
  assign n17576 = pi38  & ~n17575;
  assign n17577 = ~n17574 & ~n17575;
  assign n17578 = ~n17576 & ~n17577;
  assign n17579 = n17567 & ~n17578;
  assign n17580 = n17567 & ~n17579;
  assign n17581 = ~n17578 & ~n17579;
  assign n17582 = ~n17580 & ~n17581;
  assign n17583 = ~n17411 & ~n17582;
  assign n17584 = n17411 & n17582;
  assign n17585 = ~n17583 & ~n17584;
  assign n17586 = ~n17410 & n17585;
  assign n17587 = n17410 & ~n17585;
  assign n17588 = ~n17586 & ~n17587;
  assign n17589 = n17399 & ~n17588;
  assign n17590 = ~n17399 & n17588;
  assign n17591 = ~n17589 & ~n17590;
  assign n17592 = ~n17104 & ~n17291;
  assign n17593 = pi109  & n3550;
  assign n17594 = pi107  & n3735;
  assign n17595 = pi108  & n3545;
  assign n17596 = ~n17594 & ~n17595;
  assign n17597 = ~n17593 & n17596;
  assign n17598 = n3553 & n7170;
  assign n17599 = n17597 & ~n17598;
  assign n17600 = pi32  & ~n17599;
  assign n17601 = pi32  & ~n17600;
  assign n17602 = ~n17599 & ~n17600;
  assign n17603 = ~n17601 & ~n17602;
  assign n17604 = ~n17592 & ~n17603;
  assign n17605 = ~n17592 & ~n17604;
  assign n17606 = ~n17603 & ~n17604;
  assign n17607 = ~n17605 & ~n17606;
  assign n17608 = n17591 & ~n17607;
  assign n17609 = ~n17591 & n17607;
  assign n17610 = ~n17090 & ~n17294;
  assign n17611 = pi112  & n2976;
  assign n17612 = pi110  & n3182;
  assign n17613 = pi111  & n2971;
  assign n17614 = ~n17612 & ~n17613;
  assign n17615 = ~n17611 & n17614;
  assign n17616 = n2979 & n7795;
  assign n17617 = n17615 & ~n17616;
  assign n17618 = pi29  & ~n17617;
  assign n17619 = pi29  & ~n17618;
  assign n17620 = ~n17617 & ~n17618;
  assign n17621 = ~n17619 & ~n17620;
  assign n17622 = ~n17610 & ~n17621;
  assign n17623 = n17610 & n17621;
  assign n17624 = ~n17622 & ~n17623;
  assign n17625 = ~n17609 & n17624;
  assign n17626 = ~n17608 & n17625;
  assign n17627 = n17624 & ~n17626;
  assign n17628 = ~n17609 & ~n17626;
  assign n17629 = ~n17608 & n17628;
  assign n17630 = ~n17627 & ~n17629;
  assign n17631 = n17398 & ~n17630;
  assign n17632 = ~n17398 & n17630;
  assign n17633 = ~n17383 & ~n17632;
  assign n17634 = ~n17631 & n17633;
  assign n17635 = ~n17383 & ~n17634;
  assign n17636 = ~n17632 & ~n17634;
  assign n17637 = ~n17631 & n17636;
  assign n17638 = ~n17635 & ~n17637;
  assign n17639 = n17367 & ~n17638;
  assign n17640 = ~n17367 & n17638;
  assign n17641 = ~n17045 & ~n17323;
  assign n17642 = pi124  & n1269;
  assign n17643 = pi122  & n1340;
  assign n17644 = pi123  & n1264;
  assign n17645 = ~n17643 & ~n17644;
  assign n17646 = ~n17642 & n17645;
  assign n17647 = n1272 & n11858;
  assign n17648 = n17646 & ~n17647;
  assign n17649 = pi17  & ~n17648;
  assign n17650 = pi17  & ~n17649;
  assign n17651 = ~n17648 & ~n17649;
  assign n17652 = ~n17650 & ~n17651;
  assign n17653 = ~n17641 & ~n17652;
  assign n17654 = n17641 & n17652;
  assign n17655 = ~n17653 & ~n17654;
  assign n17656 = ~n17640 & n17655;
  assign n17657 = ~n17639 & n17656;
  assign n17658 = n17655 & ~n17657;
  assign n17659 = ~n17640 & ~n17657;
  assign n17660 = ~n17639 & n17659;
  assign n17661 = ~n17658 & ~n17660;
  assign n17662 = ~n17029 & ~n17326;
  assign n17663 = pi127  & n918;
  assign n17664 = pi125  & n1031;
  assign n17665 = pi126  & n913;
  assign n17666 = ~n17664 & ~n17665;
  assign n17667 = ~n17663 & n17666;
  assign n17668 = n921 & n13365;
  assign n17669 = n17667 & ~n17668;
  assign n17670 = pi14  & ~n17669;
  assign n17671 = pi14  & ~n17670;
  assign n17672 = ~n17669 & ~n17670;
  assign n17673 = ~n17671 & ~n17672;
  assign n17674 = ~n17662 & ~n17673;
  assign n17675 = n17662 & n17673;
  assign n17676 = ~n17674 & ~n17675;
  assign n17677 = ~n17661 & n17676;
  assign n17678 = n17661 & ~n17676;
  assign n17679 = ~n17677 & ~n17678;
  assign n17680 = n17352 & n17679;
  assign n17681 = ~n17352 & ~n17679;
  assign n17682 = ~n17680 & ~n17681;
  assign n17683 = ~n17351 & n17682;
  assign n17684 = n17351 & ~n17682;
  assign po75  = ~n17683 & ~n17684;
  assign n17686 = ~n17680 & ~n17683;
  assign n17687 = ~n17674 & ~n17677;
  assign n17688 = ~n17380 & ~n17634;
  assign n17689 = pi122  & n1582;
  assign n17690 = pi120  & n1713;
  assign n17691 = pi121  & n1577;
  assign n17692 = ~n17690 & ~n17691;
  assign n17693 = ~n17689 & n17692;
  assign n17694 = ~n1585 & n17693;
  assign n17695 = ~n11463 & n17693;
  assign n17696 = ~n17694 & ~n17695;
  assign n17697 = pi20  & ~n17696;
  assign n17698 = ~pi20  & n17696;
  assign n17699 = ~n17697 & ~n17698;
  assign n17700 = ~n17688 & ~n17699;
  assign n17701 = n17688 & n17699;
  assign n17702 = ~n17700 & ~n17701;
  assign n17703 = pi119  & n2004;
  assign n17704 = pi117  & n2141;
  assign n17705 = pi118  & n1999;
  assign n17706 = ~n17704 & ~n17705;
  assign n17707 = ~n17703 & n17706;
  assign n17708 = n2007 & n10048;
  assign n17709 = n17707 & ~n17708;
  assign n17710 = pi23  & ~n17709;
  assign n17711 = pi23  & ~n17710;
  assign n17712 = ~n17709 & ~n17710;
  assign n17713 = ~n17711 & ~n17712;
  assign n17714 = ~n17397 & ~n17631;
  assign n17715 = ~n17713 & ~n17714;
  assign n17716 = ~n17713 & ~n17715;
  assign n17717 = ~n17714 & ~n17715;
  assign n17718 = ~n17716 & ~n17717;
  assign n17719 = ~n17622 & ~n17626;
  assign n17720 = pi116  & n2486;
  assign n17721 = pi114  & n2644;
  assign n17722 = pi115  & n2481;
  assign n17723 = ~n17721 & ~n17722;
  assign n17724 = ~n17720 & n17723;
  assign n17725 = ~n2489 & n17724;
  assign n17726 = ~n9042 & n17724;
  assign n17727 = ~n17725 & ~n17726;
  assign n17728 = pi26  & ~n17727;
  assign n17729 = ~pi26  & n17727;
  assign n17730 = ~n17728 & ~n17729;
  assign n17731 = ~n17719 & ~n17730;
  assign n17732 = n17719 & n17730;
  assign n17733 = ~n17731 & ~n17732;
  assign n17734 = pi113  & n2976;
  assign n17735 = pi111  & n3182;
  assign n17736 = pi112  & n2971;
  assign n17737 = ~n17735 & ~n17736;
  assign n17738 = ~n17734 & n17737;
  assign n17739 = n2979 & n8387;
  assign n17740 = n17738 & ~n17739;
  assign n17741 = pi29  & ~n17740;
  assign n17742 = pi29  & ~n17741;
  assign n17743 = ~n17740 & ~n17741;
  assign n17744 = ~n17742 & ~n17743;
  assign n17745 = ~n17604 & ~n17608;
  assign n17746 = ~n17744 & ~n17745;
  assign n17747 = n17744 & n17745;
  assign n17748 = ~n17746 & ~n17747;
  assign n17749 = ~n17579 & ~n17583;
  assign n17750 = pi104  & n4896;
  assign n17751 = pi102  & n5148;
  assign n17752 = pi103  & n4891;
  assign n17753 = ~n17751 & ~n17752;
  assign n17754 = ~n17750 & n17753;
  assign n17755 = n4899 & n5565;
  assign n17756 = n17754 & ~n17755;
  assign n17757 = pi38  & ~n17756;
  assign n17758 = pi38  & ~n17757;
  assign n17759 = ~n17756 & ~n17757;
  assign n17760 = ~n17758 & ~n17759;
  assign n17761 = ~n17562 & ~n17566;
  assign n17762 = pi101  & n5636;
  assign n17763 = pi99  & n5909;
  assign n17764 = pi100  & n5631;
  assign n17765 = ~n17763 & ~n17764;
  assign n17766 = ~n17762 & n17765;
  assign n17767 = n5056 & n5639;
  assign n17768 = n17766 & ~n17767;
  assign n17769 = pi41  & ~n17768;
  assign n17770 = pi41  & ~n17769;
  assign n17771 = ~n17768 & ~n17769;
  assign n17772 = ~n17770 & ~n17771;
  assign n17773 = ~n17556 & ~n17559;
  assign n17774 = pi98  & n6396;
  assign n17775 = pi96  & n6735;
  assign n17776 = pi97  & n6391;
  assign n17777 = ~n17775 & ~n17776;
  assign n17778 = ~n17774 & n17777;
  assign n17779 = n4360 & n6399;
  assign n17780 = n17778 & ~n17779;
  assign n17781 = pi44  & ~n17780;
  assign n17782 = pi44  & ~n17781;
  assign n17783 = ~n17780 & ~n17781;
  assign n17784 = ~n17782 & ~n17783;
  assign n17785 = pi95  & n7239;
  assign n17786 = pi93  & n7556;
  assign n17787 = pi94  & n7234;
  assign n17788 = ~n17786 & ~n17787;
  assign n17789 = ~n17785 & n17788;
  assign n17790 = n3710 & n7242;
  assign n17791 = n17789 & ~n17790;
  assign n17792 = pi47  & ~n17791;
  assign n17793 = pi47  & ~n17792;
  assign n17794 = ~n17791 & ~n17792;
  assign n17795 = ~n17793 & ~n17794;
  assign n17796 = ~n17520 & ~n17524;
  assign n17797 = ~n17503 & ~n17506;
  assign n17798 = ~n17497 & ~n17500;
  assign n17799 = ~n17461 & ~n17464;
  assign n17800 = pi80  & n12295;
  assign n17801 = pi78  & n12693;
  assign n17802 = pi79  & n12290;
  assign n17803 = ~n17801 & ~n17802;
  assign n17804 = ~n17800 & n17803;
  assign n17805 = n1205 & n12298;
  assign n17806 = n17804 & ~n17805;
  assign n17807 = pi62  & ~n17806;
  assign n17808 = pi62  & ~n17807;
  assign n17809 = ~n17806 & ~n17807;
  assign n17810 = ~n17808 & ~n17809;
  assign n17811 = pi76  & n13477;
  assign n17812 = pi77  & ~n13122;
  assign n17813 = ~n17811 & ~n17812;
  assign n17814 = ~n17455 & ~n17458;
  assign n17815 = n17813 & ~n17814;
  assign n17816 = ~n17813 & n17814;
  assign n17817 = ~n17815 & ~n17816;
  assign n17818 = ~n17810 & n17817;
  assign n17819 = n17810 & ~n17817;
  assign n17820 = ~n17818 & ~n17819;
  assign n17821 = n17799 & ~n17820;
  assign n17822 = ~n17799 & n17820;
  assign n17823 = ~n17821 & ~n17822;
  assign n17824 = pi83  & n11193;
  assign n17825 = pi81  & n11567;
  assign n17826 = pi82  & n11188;
  assign n17827 = ~n17825 & ~n17826;
  assign n17828 = ~n17824 & n17827;
  assign n17829 = n1672 & n11196;
  assign n17830 = n17828 & ~n17829;
  assign n17831 = pi59  & ~n17830;
  assign n17832 = pi59  & ~n17831;
  assign n17833 = ~n17830 & ~n17831;
  assign n17834 = ~n17832 & ~n17833;
  assign n17835 = n17823 & ~n17834;
  assign n17836 = n17823 & ~n17835;
  assign n17837 = ~n17834 & ~n17835;
  assign n17838 = ~n17836 & ~n17837;
  assign n17839 = ~n17478 & ~n17484;
  assign n17840 = n17838 & n17839;
  assign n17841 = ~n17838 & ~n17839;
  assign n17842 = ~n17840 & ~n17841;
  assign n17843 = pi86  & n10135;
  assign n17844 = pi84  & n10478;
  assign n17845 = pi85  & n10130;
  assign n17846 = ~n17844 & ~n17845;
  assign n17847 = ~n17843 & n17846;
  assign n17848 = n2099 & n10138;
  assign n17849 = n17847 & ~n17848;
  assign n17850 = pi56  & ~n17849;
  assign n17851 = pi56  & ~n17850;
  assign n17852 = ~n17849 & ~n17850;
  assign n17853 = ~n17851 & ~n17852;
  assign n17854 = n17842 & ~n17853;
  assign n17855 = ~n17842 & n17853;
  assign n17856 = ~n17854 & ~n17855;
  assign n17857 = n17798 & ~n17856;
  assign n17858 = ~n17798 & n17856;
  assign n17859 = ~n17857 & ~n17858;
  assign n17860 = pi89  & n9096;
  assign n17861 = pi87  & n9453;
  assign n17862 = pi88  & n9091;
  assign n17863 = ~n17861 & ~n17862;
  assign n17864 = ~n17860 & n17863;
  assign n17865 = n2432 & n9099;
  assign n17866 = n17864 & ~n17865;
  assign n17867 = pi53  & ~n17866;
  assign n17868 = pi53  & ~n17867;
  assign n17869 = ~n17866 & ~n17867;
  assign n17870 = ~n17868 & ~n17869;
  assign n17871 = n17859 & ~n17870;
  assign n17872 = ~n17859 & n17870;
  assign n17873 = ~n17871 & ~n17872;
  assign n17874 = n17797 & ~n17873;
  assign n17875 = ~n17797 & n17873;
  assign n17876 = ~n17874 & ~n17875;
  assign n17877 = pi92  & n8137;
  assign n17878 = pi90  & n8471;
  assign n17879 = pi91  & n8132;
  assign n17880 = ~n17878 & ~n17879;
  assign n17881 = ~n17877 & n17880;
  assign n17882 = n3119 & n8140;
  assign n17883 = n17881 & ~n17882;
  assign n17884 = pi50  & ~n17883;
  assign n17885 = pi50  & ~n17884;
  assign n17886 = ~n17883 & ~n17884;
  assign n17887 = ~n17885 & ~n17886;
  assign n17888 = ~n17876 & n17887;
  assign n17889 = n17876 & ~n17887;
  assign n17890 = ~n17888 & ~n17889;
  assign n17891 = ~n17796 & n17890;
  assign n17892 = n17796 & ~n17890;
  assign n17893 = ~n17891 & ~n17892;
  assign n17894 = ~n17795 & n17893;
  assign n17895 = n17795 & ~n17893;
  assign n17896 = ~n17894 & ~n17895;
  assign n17897 = ~n17542 & n17896;
  assign n17898 = n17542 & ~n17896;
  assign n17899 = ~n17897 & ~n17898;
  assign n17900 = ~n17784 & n17899;
  assign n17901 = n17784 & ~n17899;
  assign n17902 = ~n17900 & ~n17901;
  assign n17903 = ~n17773 & n17902;
  assign n17904 = n17773 & ~n17902;
  assign n17905 = ~n17903 & ~n17904;
  assign n17906 = ~n17772 & n17905;
  assign n17907 = n17772 & ~n17905;
  assign n17908 = ~n17906 & ~n17907;
  assign n17909 = ~n17761 & n17908;
  assign n17910 = n17761 & ~n17908;
  assign n17911 = ~n17909 & ~n17910;
  assign n17912 = ~n17760 & n17911;
  assign n17913 = n17760 & ~n17911;
  assign n17914 = ~n17912 & ~n17913;
  assign n17915 = ~n17749 & n17914;
  assign n17916 = n17749 & ~n17914;
  assign n17917 = ~n17915 & ~n17916;
  assign n17918 = pi107  & n4182;
  assign n17919 = pi105  & n4416;
  assign n17920 = pi106  & n4177;
  assign n17921 = ~n17919 & ~n17920;
  assign n17922 = ~n17918 & n17921;
  assign n17923 = n4185 & n6614;
  assign n17924 = n17922 & ~n17923;
  assign n17925 = pi35  & ~n17924;
  assign n17926 = pi35  & ~n17925;
  assign n17927 = ~n17924 & ~n17925;
  assign n17928 = ~n17926 & ~n17927;
  assign n17929 = n17917 & ~n17928;
  assign n17930 = ~n17917 & n17928;
  assign n17931 = ~n17929 & ~n17930;
  assign n17932 = ~n17586 & ~n17590;
  assign n17933 = pi110  & n3550;
  assign n17934 = pi108  & n3735;
  assign n17935 = pi109  & n3545;
  assign n17936 = ~n17934 & ~n17935;
  assign n17937 = ~n17933 & n17936;
  assign n17938 = ~n3553 & n17937;
  assign n17939 = ~n7474 & n17937;
  assign n17940 = ~n17938 & ~n17939;
  assign n17941 = pi32  & ~n17940;
  assign n17942 = ~pi32  & n17940;
  assign n17943 = ~n17941 & ~n17942;
  assign n17944 = ~n17932 & ~n17943;
  assign n17945 = n17932 & n17943;
  assign n17946 = ~n17944 & ~n17945;
  assign n17947 = n17931 & n17946;
  assign n17948 = ~n17931 & ~n17946;
  assign n17949 = ~n17947 & ~n17948;
  assign n17950 = n17748 & n17949;
  assign n17951 = ~n17748 & ~n17949;
  assign n17952 = ~n17950 & ~n17951;
  assign n17953 = n17733 & n17952;
  assign n17954 = ~n17733 & ~n17952;
  assign n17955 = ~n17953 & ~n17954;
  assign n17956 = ~n17718 & n17955;
  assign n17957 = n17718 & ~n17955;
  assign n17958 = ~n17956 & ~n17957;
  assign n17959 = n17702 & n17958;
  assign n17960 = ~n17702 & ~n17958;
  assign n17961 = ~n17959 & ~n17960;
  assign n17962 = pi125  & n1269;
  assign n17963 = pi123  & n1340;
  assign n17964 = pi124  & n1264;
  assign n17965 = ~n17963 & ~n17964;
  assign n17966 = ~n17962 & n17965;
  assign n17967 = n1272 & n12591;
  assign n17968 = n17966 & ~n17967;
  assign n17969 = pi17  & ~n17968;
  assign n17970 = pi17  & ~n17969;
  assign n17971 = ~n17968 & ~n17969;
  assign n17972 = ~n17970 & ~n17971;
  assign n17973 = ~n17366 & ~n17639;
  assign n17974 = ~n17972 & ~n17973;
  assign n17975 = n17972 & n17973;
  assign n17976 = ~n17974 & ~n17975;
  assign n17977 = n17961 & n17976;
  assign n17978 = ~n17961 & ~n17976;
  assign n17979 = ~n17977 & ~n17978;
  assign n17980 = ~n17653 & ~n17657;
  assign n17981 = pi126  & n1031;
  assign n17982 = pi127  & n913;
  assign n17983 = ~n17981 & ~n17982;
  assign n17984 = ~n921 & n17983;
  assign n17985 = ~n13389 & n17983;
  assign n17986 = ~n17984 & ~n17985;
  assign n17987 = pi14  & ~n17986;
  assign n17988 = ~pi14  & n17986;
  assign n17989 = ~n17987 & ~n17988;
  assign n17990 = ~n17980 & ~n17989;
  assign n17991 = n17980 & n17989;
  assign n17992 = ~n17990 & ~n17991;
  assign n17993 = n17979 & n17992;
  assign n17994 = ~n17979 & ~n17992;
  assign n17995 = ~n17993 & ~n17994;
  assign n17996 = ~n17687 & n17995;
  assign n17997 = n17687 & ~n17995;
  assign n17998 = ~n17996 & ~n17997;
  assign n17999 = ~n17686 & n17998;
  assign n18000 = n17686 & ~n17998;
  assign po76  = ~n17999 & ~n18000;
  assign n18002 = ~n17996 & ~n17999;
  assign n18003 = ~n17990 & ~n17993;
  assign n18004 = pi123  & n1582;
  assign n18005 = pi121  & n1713;
  assign n18006 = pi122  & n1577;
  assign n18007 = ~n18005 & ~n18006;
  assign n18008 = ~n18004 & n18007;
  assign n18009 = n1585 & n11489;
  assign n18010 = n18008 & ~n18009;
  assign n18011 = pi20  & ~n18010;
  assign n18012 = pi20  & ~n18011;
  assign n18013 = ~n18010 & ~n18011;
  assign n18014 = ~n18012 & ~n18013;
  assign n18015 = ~n17715 & ~n17956;
  assign n18016 = n18014 & n18015;
  assign n18017 = ~n18014 & ~n18015;
  assign n18018 = ~n18016 & ~n18017;
  assign n18019 = pi120  & n2004;
  assign n18020 = pi118  & n2141;
  assign n18021 = pi119  & n1999;
  assign n18022 = ~n18020 & ~n18021;
  assign n18023 = ~n18019 & n18022;
  assign n18024 = n2007 & n10734;
  assign n18025 = n18023 & ~n18024;
  assign n18026 = pi23  & ~n18025;
  assign n18027 = pi23  & ~n18026;
  assign n18028 = ~n18025 & ~n18026;
  assign n18029 = ~n18027 & ~n18028;
  assign n18030 = ~n17731 & ~n17953;
  assign n18031 = n18029 & n18030;
  assign n18032 = ~n18029 & ~n18030;
  assign n18033 = ~n18031 & ~n18032;
  assign n18034 = pi117  & n2486;
  assign n18035 = pi115  & n2644;
  assign n18036 = pi116  & n2481;
  assign n18037 = ~n18035 & ~n18036;
  assign n18038 = ~n18034 & n18037;
  assign n18039 = n2489 & n9691;
  assign n18040 = n18038 & ~n18039;
  assign n18041 = pi26  & ~n18040;
  assign n18042 = pi26  & ~n18041;
  assign n18043 = ~n18040 & ~n18041;
  assign n18044 = ~n18042 & ~n18043;
  assign n18045 = ~n17746 & ~n17950;
  assign n18046 = n18044 & n18045;
  assign n18047 = ~n18044 & ~n18045;
  assign n18048 = ~n18046 & ~n18047;
  assign n18049 = ~n17944 & ~n17947;
  assign n18050 = pi114  & n2976;
  assign n18051 = pi112  & n3182;
  assign n18052 = pi113  & n2971;
  assign n18053 = ~n18051 & ~n18052;
  assign n18054 = ~n18050 & n18053;
  assign n18055 = ~n2979 & n18054;
  assign n18056 = ~n8702 & n18054;
  assign n18057 = ~n18055 & ~n18056;
  assign n18058 = pi29  & ~n18057;
  assign n18059 = ~pi29  & n18057;
  assign n18060 = ~n18058 & ~n18059;
  assign n18061 = ~n18049 & ~n18060;
  assign n18062 = n18049 & n18060;
  assign n18063 = ~n18061 & ~n18062;
  assign n18064 = ~n17915 & ~n17929;
  assign n18065 = pi111  & n3550;
  assign n18066 = pi109  & n3735;
  assign n18067 = pi110  & n3545;
  assign n18068 = ~n18066 & ~n18067;
  assign n18069 = ~n18065 & n18068;
  assign n18070 = ~n3553 & n18069;
  assign n18071 = ~n7770 & n18069;
  assign n18072 = ~n18070 & ~n18071;
  assign n18073 = pi32  & ~n18072;
  assign n18074 = ~pi32  & n18072;
  assign n18075 = ~n18073 & ~n18074;
  assign n18076 = ~n18064 & ~n18075;
  assign n18077 = n18064 & n18075;
  assign n18078 = ~n18076 & ~n18077;
  assign n18079 = pi108  & n4182;
  assign n18080 = pi106  & n4416;
  assign n18081 = pi107  & n4177;
  assign n18082 = ~n18080 & ~n18081;
  assign n18083 = ~n18079 & n18082;
  assign n18084 = n4185 & n6639;
  assign n18085 = n18083 & ~n18084;
  assign n18086 = pi35  & ~n18085;
  assign n18087 = pi35  & ~n18086;
  assign n18088 = ~n18085 & ~n18086;
  assign n18089 = ~n18087 & ~n18088;
  assign n18090 = ~n17909 & ~n17912;
  assign n18091 = pi105  & n4896;
  assign n18092 = pi103  & n5148;
  assign n18093 = pi104  & n4891;
  assign n18094 = ~n18092 & ~n18093;
  assign n18095 = ~n18091 & n18094;
  assign n18096 = n4899 & n6065;
  assign n18097 = n18095 & ~n18096;
  assign n18098 = pi38  & ~n18097;
  assign n18099 = pi38  & ~n18098;
  assign n18100 = ~n18097 & ~n18098;
  assign n18101 = ~n18099 & ~n18100;
  assign n18102 = ~n17903 & ~n17906;
  assign n18103 = ~n17897 & ~n17900;
  assign n18104 = ~n17891 & ~n17894;
  assign n18105 = pi96  & n7239;
  assign n18106 = pi94  & n7556;
  assign n18107 = pi95  & n7234;
  assign n18108 = ~n18106 & ~n18107;
  assign n18109 = ~n18105 & n18108;
  assign n18110 = n3921 & n7242;
  assign n18111 = n18109 & ~n18110;
  assign n18112 = pi47  & ~n18111;
  assign n18113 = pi47  & ~n18112;
  assign n18114 = ~n18111 & ~n18112;
  assign n18115 = ~n18113 & ~n18114;
  assign n18116 = ~n17858 & ~n17871;
  assign n18117 = pi90  & n9096;
  assign n18118 = pi88  & n9453;
  assign n18119 = pi89  & n9091;
  assign n18120 = ~n18118 & ~n18119;
  assign n18121 = ~n18117 & n18120;
  assign n18122 = n2606 & n9099;
  assign n18123 = n18121 & ~n18122;
  assign n18124 = pi53  & ~n18123;
  assign n18125 = pi53  & ~n18124;
  assign n18126 = ~n18123 & ~n18124;
  assign n18127 = ~n18125 & ~n18126;
  assign n18128 = ~n17841 & ~n17854;
  assign n18129 = ~n17815 & ~n17818;
  assign n18130 = pi77  & n13477;
  assign n18131 = pi78  & ~n13122;
  assign n18132 = ~n18130 & ~n18131;
  assign n18133 = n17813 & ~n18132;
  assign n18134 = ~n17813 & n18132;
  assign n18135 = ~n18133 & ~n18134;
  assign n18136 = pi81  & n12295;
  assign n18137 = pi79  & n12693;
  assign n18138 = pi80  & n12290;
  assign n18139 = ~n18137 & ~n18138;
  assign n18140 = ~n18136 & n18139;
  assign n18141 = ~n12298 & n18140;
  assign n18142 = ~n1413 & n18140;
  assign n18143 = ~n18141 & ~n18142;
  assign n18144 = pi62  & ~n18143;
  assign n18145 = ~pi62  & n18143;
  assign n18146 = ~n18144 & ~n18145;
  assign n18147 = n18135 & ~n18146;
  assign n18148 = ~n18135 & n18146;
  assign n18149 = ~n18147 & ~n18148;
  assign n18150 = ~n18129 & n18149;
  assign n18151 = n18129 & ~n18149;
  assign n18152 = ~n18150 & ~n18151;
  assign n18153 = pi84  & n11193;
  assign n18154 = pi82  & n11567;
  assign n18155 = pi83  & n11188;
  assign n18156 = ~n18154 & ~n18155;
  assign n18157 = ~n18153 & n18156;
  assign n18158 = n1805 & n11196;
  assign n18159 = n18157 & ~n18158;
  assign n18160 = pi59  & ~n18159;
  assign n18161 = pi59  & ~n18160;
  assign n18162 = ~n18159 & ~n18160;
  assign n18163 = ~n18161 & ~n18162;
  assign n18164 = n18152 & ~n18163;
  assign n18165 = n18152 & ~n18164;
  assign n18166 = ~n18163 & ~n18164;
  assign n18167 = ~n18165 & ~n18166;
  assign n18168 = ~n17822 & ~n17835;
  assign n18169 = n18167 & n18168;
  assign n18170 = ~n18167 & ~n18168;
  assign n18171 = ~n18169 & ~n18170;
  assign n18172 = pi87  & n10135;
  assign n18173 = pi85  & n10478;
  assign n18174 = pi86  & n10130;
  assign n18175 = ~n18173 & ~n18174;
  assign n18176 = ~n18172 & n18175;
  assign n18177 = n2252 & n10138;
  assign n18178 = n18176 & ~n18177;
  assign n18179 = pi56  & ~n18178;
  assign n18180 = pi56  & ~n18179;
  assign n18181 = ~n18178 & ~n18179;
  assign n18182 = ~n18180 & ~n18181;
  assign n18183 = ~n18171 & n18182;
  assign n18184 = n18171 & ~n18182;
  assign n18185 = ~n18183 & ~n18184;
  assign n18186 = ~n18128 & n18185;
  assign n18187 = n18128 & ~n18185;
  assign n18188 = ~n18186 & ~n18187;
  assign n18189 = ~n18127 & n18188;
  assign n18190 = n18127 & ~n18188;
  assign n18191 = ~n18189 & ~n18190;
  assign n18192 = ~n18116 & n18191;
  assign n18193 = n18116 & ~n18191;
  assign n18194 = ~n18192 & ~n18193;
  assign n18195 = pi93  & n8137;
  assign n18196 = pi91  & n8471;
  assign n18197 = pi92  & n8132;
  assign n18198 = ~n18196 & ~n18197;
  assign n18199 = ~n18195 & n18198;
  assign n18200 = n3144 & n8140;
  assign n18201 = n18199 & ~n18200;
  assign n18202 = pi50  & ~n18201;
  assign n18203 = pi50  & ~n18202;
  assign n18204 = ~n18201 & ~n18202;
  assign n18205 = ~n18203 & ~n18204;
  assign n18206 = n18194 & ~n18205;
  assign n18207 = n18194 & ~n18206;
  assign n18208 = ~n18205 & ~n18206;
  assign n18209 = ~n18207 & ~n18208;
  assign n18210 = ~n17875 & ~n17889;
  assign n18211 = ~n18209 & ~n18210;
  assign n18212 = n18209 & n18210;
  assign n18213 = ~n18211 & ~n18212;
  assign n18214 = n18115 & n18213;
  assign n18215 = ~n18115 & ~n18213;
  assign n18216 = ~n18214 & ~n18215;
  assign n18217 = n18104 & n18216;
  assign n18218 = ~n18104 & ~n18216;
  assign n18219 = ~n18217 & ~n18218;
  assign n18220 = pi99  & n6396;
  assign n18221 = pi97  & n6735;
  assign n18222 = pi98  & n6391;
  assign n18223 = ~n18221 & ~n18222;
  assign n18224 = ~n18220 & n18223;
  assign n18225 = n4584 & n6399;
  assign n18226 = n18224 & ~n18225;
  assign n18227 = pi44  & ~n18226;
  assign n18228 = pi44  & ~n18227;
  assign n18229 = ~n18226 & ~n18227;
  assign n18230 = ~n18228 & ~n18229;
  assign n18231 = n18219 & ~n18230;
  assign n18232 = ~n18219 & n18230;
  assign n18233 = ~n18231 & ~n18232;
  assign n18234 = n18103 & ~n18233;
  assign n18235 = ~n18103 & n18233;
  assign n18236 = ~n18234 & ~n18235;
  assign n18237 = pi102  & n5636;
  assign n18238 = pi100  & n5909;
  assign n18239 = pi101  & n5631;
  assign n18240 = ~n18238 & ~n18239;
  assign n18241 = ~n18237 & n18240;
  assign n18242 = n5296 & n5639;
  assign n18243 = n18241 & ~n18242;
  assign n18244 = pi41  & ~n18243;
  assign n18245 = pi41  & ~n18244;
  assign n18246 = ~n18243 & ~n18244;
  assign n18247 = ~n18245 & ~n18246;
  assign n18248 = ~n18236 & n18247;
  assign n18249 = n18236 & ~n18247;
  assign n18250 = ~n18248 & ~n18249;
  assign n18251 = ~n18102 & n18250;
  assign n18252 = n18102 & ~n18250;
  assign n18253 = ~n18251 & ~n18252;
  assign n18254 = ~n18101 & n18253;
  assign n18255 = n18101 & ~n18253;
  assign n18256 = ~n18254 & ~n18255;
  assign n18257 = ~n18090 & n18256;
  assign n18258 = n18090 & ~n18256;
  assign n18259 = ~n18257 & ~n18258;
  assign n18260 = ~n18089 & n18259;
  assign n18261 = ~n18089 & ~n18260;
  assign n18262 = n18259 & ~n18260;
  assign n18263 = ~n18261 & ~n18262;
  assign n18264 = n18078 & ~n18263;
  assign n18265 = ~n18078 & n18263;
  assign n18266 = ~n18264 & ~n18265;
  assign n18267 = n18063 & n18266;
  assign n18268 = ~n18063 & ~n18266;
  assign n18269 = ~n18267 & ~n18268;
  assign n18270 = n18048 & n18269;
  assign n18271 = ~n18048 & ~n18269;
  assign n18272 = ~n18270 & ~n18271;
  assign n18273 = n18033 & n18272;
  assign n18274 = ~n18033 & ~n18272;
  assign n18275 = n18018 & ~n18274;
  assign n18276 = ~n18273 & n18275;
  assign n18277 = n18018 & ~n18276;
  assign n18278 = ~n18274 & ~n18276;
  assign n18279 = ~n18273 & n18278;
  assign n18280 = ~n18277 & ~n18279;
  assign n18281 = ~n17700 & ~n17959;
  assign n18282 = pi126  & n1269;
  assign n18283 = pi124  & n1340;
  assign n18284 = pi125  & n1264;
  assign n18285 = ~n18283 & ~n18284;
  assign n18286 = ~n18282 & n18285;
  assign n18287 = ~n1272 & n18286;
  assign n18288 = ~n12979 & n18286;
  assign n18289 = ~n18287 & ~n18288;
  assign n18290 = pi17  & ~n18289;
  assign n18291 = ~pi17  & n18289;
  assign n18292 = ~n18290 & ~n18291;
  assign n18293 = ~n18281 & ~n18292;
  assign n18294 = ~n18281 & ~n18293;
  assign n18295 = ~n18292 & ~n18293;
  assign n18296 = ~n18294 & ~n18295;
  assign n18297 = ~n18280 & ~n18296;
  assign n18298 = n18280 & n18296;
  assign n18299 = ~n18297 & ~n18298;
  assign n18300 = ~n17974 & ~n17977;
  assign n18301 = pi127  & n1031;
  assign n18302 = n921 & n13387;
  assign n18303 = ~n18301 & ~n18302;
  assign n18304 = pi14  & ~n18303;
  assign n18305 = pi14  & ~n18304;
  assign n18306 = ~n18303 & ~n18304;
  assign n18307 = ~n18305 & ~n18306;
  assign n18308 = ~n18300 & ~n18307;
  assign n18309 = n18300 & n18307;
  assign n18310 = ~n18308 & ~n18309;
  assign n18311 = n18299 & n18310;
  assign n18312 = ~n18299 & ~n18310;
  assign n18313 = ~n18311 & ~n18312;
  assign n18314 = ~n18003 & n18313;
  assign n18315 = n18003 & ~n18313;
  assign n18316 = ~n18314 & ~n18315;
  assign n18317 = ~n18002 & n18316;
  assign n18318 = n18002 & ~n18316;
  assign po77  = ~n18317 & ~n18318;
  assign n18320 = ~n18293 & ~n18297;
  assign n18321 = pi127  & n1269;
  assign n18322 = pi125  & n1340;
  assign n18323 = pi126  & n1264;
  assign n18324 = ~n18322 & ~n18323;
  assign n18325 = ~n18321 & n18324;
  assign n18326 = n1272 & n13365;
  assign n18327 = n18325 & ~n18326;
  assign n18328 = pi17  & ~n18327;
  assign n18329 = pi17  & ~n18328;
  assign n18330 = ~n18327 & ~n18328;
  assign n18331 = ~n18329 & ~n18330;
  assign n18332 = ~n18320 & ~n18331;
  assign n18333 = n18320 & n18331;
  assign n18334 = ~n18332 & ~n18333;
  assign n18335 = pi124  & n1582;
  assign n18336 = pi122  & n1713;
  assign n18337 = pi123  & n1577;
  assign n18338 = ~n18336 & ~n18337;
  assign n18339 = ~n18335 & n18338;
  assign n18340 = n1585 & n11858;
  assign n18341 = n18339 & ~n18340;
  assign n18342 = pi20  & ~n18341;
  assign n18343 = pi20  & ~n18342;
  assign n18344 = ~n18341 & ~n18342;
  assign n18345 = ~n18343 & ~n18344;
  assign n18346 = ~n18017 & ~n18276;
  assign n18347 = n18345 & n18346;
  assign n18348 = ~n18345 & ~n18346;
  assign n18349 = ~n18347 & ~n18348;
  assign n18350 = ~n18032 & ~n18273;
  assign n18351 = pi121  & n2004;
  assign n18352 = pi119  & n2141;
  assign n18353 = pi120  & n1999;
  assign n18354 = ~n18352 & ~n18353;
  assign n18355 = ~n18351 & n18354;
  assign n18356 = n2007 & n11086;
  assign n18357 = n18355 & ~n18356;
  assign n18358 = pi23  & ~n18357;
  assign n18359 = pi23  & ~n18358;
  assign n18360 = ~n18357 & ~n18358;
  assign n18361 = ~n18359 & ~n18360;
  assign n18362 = ~n18350 & n18361;
  assign n18363 = n18350 & ~n18361;
  assign n18364 = ~n18362 & ~n18363;
  assign n18365 = pi118  & n2486;
  assign n18366 = pi116  & n2644;
  assign n18367 = pi117  & n2481;
  assign n18368 = ~n18366 & ~n18367;
  assign n18369 = ~n18365 & n18368;
  assign n18370 = n2489 & n9716;
  assign n18371 = n18369 & ~n18370;
  assign n18372 = pi26  & ~n18371;
  assign n18373 = pi26  & ~n18372;
  assign n18374 = ~n18371 & ~n18372;
  assign n18375 = ~n18373 & ~n18374;
  assign n18376 = ~n18047 & ~n18270;
  assign n18377 = n18375 & n18376;
  assign n18378 = ~n18375 & ~n18376;
  assign n18379 = ~n18377 & ~n18378;
  assign n18380 = pi115  & n2976;
  assign n18381 = pi113  & n3182;
  assign n18382 = pi114  & n2971;
  assign n18383 = ~n18381 & ~n18382;
  assign n18384 = ~n18380 & n18383;
  assign n18385 = n2979 & n8727;
  assign n18386 = n18384 & ~n18385;
  assign n18387 = pi29  & ~n18386;
  assign n18388 = pi29  & ~n18387;
  assign n18389 = ~n18386 & ~n18387;
  assign n18390 = ~n18388 & ~n18389;
  assign n18391 = ~n18061 & ~n18267;
  assign n18392 = n18390 & n18391;
  assign n18393 = ~n18390 & ~n18391;
  assign n18394 = ~n18392 & ~n18393;
  assign n18395 = ~n18251 & ~n18254;
  assign n18396 = pi106  & n4896;
  assign n18397 = pi104  & n5148;
  assign n18398 = pi105  & n4891;
  assign n18399 = ~n18397 & ~n18398;
  assign n18400 = ~n18396 & n18399;
  assign n18401 = n4899 & n6090;
  assign n18402 = n18400 & ~n18401;
  assign n18403 = pi38  & ~n18402;
  assign n18404 = pi38  & ~n18403;
  assign n18405 = ~n18402 & ~n18403;
  assign n18406 = ~n18404 & ~n18405;
  assign n18407 = ~n18235 & ~n18249;
  assign n18408 = ~n18218 & ~n18231;
  assign n18409 = ~n18212 & ~n18214;
  assign n18410 = ~n18192 & ~n18206;
  assign n18411 = ~n18186 & ~n18189;
  assign n18412 = ~n18170 & ~n18184;
  assign n18413 = ~n18150 & ~n18164;
  assign n18414 = ~n18133 & ~n18147;
  assign n18415 = pi82  & n12295;
  assign n18416 = pi80  & n12693;
  assign n18417 = pi81  & n12290;
  assign n18418 = ~n18416 & ~n18417;
  assign n18419 = ~n18415 & n18418;
  assign n18420 = n1532 & n12298;
  assign n18421 = n18419 & ~n18420;
  assign n18422 = pi62  & ~n18421;
  assign n18423 = pi62  & ~n18422;
  assign n18424 = ~n18421 & ~n18422;
  assign n18425 = ~n18423 & ~n18424;
  assign n18426 = pi78  & n13477;
  assign n18427 = pi79  & ~n13122;
  assign n18428 = ~n18426 & ~n18427;
  assign n18429 = ~pi14  & ~n18428;
  assign n18430 = pi14  & n18428;
  assign n18431 = ~n18429 & ~n18430;
  assign n18432 = ~n17813 & n18431;
  assign n18433 = n17813 & ~n18431;
  assign n18434 = ~n18432 & ~n18433;
  assign n18435 = ~n18425 & n18434;
  assign n18436 = n18425 & ~n18434;
  assign n18437 = ~n18435 & ~n18436;
  assign n18438 = n18414 & ~n18437;
  assign n18439 = ~n18414 & n18437;
  assign n18440 = ~n18438 & ~n18439;
  assign n18441 = pi85  & n11193;
  assign n18442 = pi83  & n11567;
  assign n18443 = pi84  & n11188;
  assign n18444 = ~n18442 & ~n18443;
  assign n18445 = ~n18441 & n18444;
  assign n18446 = n1943 & n11196;
  assign n18447 = n18445 & ~n18446;
  assign n18448 = pi59  & ~n18447;
  assign n18449 = pi59  & ~n18448;
  assign n18450 = ~n18447 & ~n18448;
  assign n18451 = ~n18449 & ~n18450;
  assign n18452 = n18440 & ~n18451;
  assign n18453 = ~n18440 & n18451;
  assign n18454 = ~n18452 & ~n18453;
  assign n18455 = n18413 & ~n18454;
  assign n18456 = ~n18413 & n18454;
  assign n18457 = ~n18455 & ~n18456;
  assign n18458 = pi88  & n10135;
  assign n18459 = pi86  & n10478;
  assign n18460 = pi87  & n10130;
  assign n18461 = ~n18459 & ~n18460;
  assign n18462 = ~n18458 & n18461;
  assign n18463 = n2277 & n10138;
  assign n18464 = n18462 & ~n18463;
  assign n18465 = pi56  & ~n18464;
  assign n18466 = pi56  & ~n18465;
  assign n18467 = ~n18464 & ~n18465;
  assign n18468 = ~n18466 & ~n18467;
  assign n18469 = n18457 & ~n18468;
  assign n18470 = ~n18457 & n18468;
  assign n18471 = ~n18412 & ~n18470;
  assign n18472 = ~n18469 & n18471;
  assign n18473 = ~n18412 & ~n18472;
  assign n18474 = ~n18469 & ~n18472;
  assign n18475 = ~n18470 & n18474;
  assign n18476 = ~n18473 & ~n18475;
  assign n18477 = pi91  & n9096;
  assign n18478 = pi89  & n9453;
  assign n18479 = pi90  & n9091;
  assign n18480 = ~n18478 & ~n18479;
  assign n18481 = ~n18477 & n18480;
  assign n18482 = n2926 & n9099;
  assign n18483 = n18481 & ~n18482;
  assign n18484 = pi53  & ~n18483;
  assign n18485 = pi53  & ~n18484;
  assign n18486 = ~n18483 & ~n18484;
  assign n18487 = ~n18485 & ~n18486;
  assign n18488 = ~n18476 & ~n18487;
  assign n18489 = n18476 & n18487;
  assign n18490 = ~n18488 & ~n18489;
  assign n18491 = n18411 & ~n18490;
  assign n18492 = ~n18411 & n18490;
  assign n18493 = ~n18491 & ~n18492;
  assign n18494 = pi94  & n8137;
  assign n18495 = pi92  & n8471;
  assign n18496 = pi93  & n8132;
  assign n18497 = ~n18495 & ~n18496;
  assign n18498 = ~n18494 & n18497;
  assign n18499 = n3499 & n8140;
  assign n18500 = n18498 & ~n18499;
  assign n18501 = pi50  & ~n18500;
  assign n18502 = pi50  & ~n18501;
  assign n18503 = ~n18500 & ~n18501;
  assign n18504 = ~n18502 & ~n18503;
  assign n18505 = n18493 & ~n18504;
  assign n18506 = ~n18493 & n18504;
  assign n18507 = ~n18505 & ~n18506;
  assign n18508 = n18410 & ~n18507;
  assign n18509 = ~n18410 & n18507;
  assign n18510 = ~n18508 & ~n18509;
  assign n18511 = pi97  & n7239;
  assign n18512 = pi95  & n7556;
  assign n18513 = pi96  & n7234;
  assign n18514 = ~n18512 & ~n18513;
  assign n18515 = ~n18511 & n18514;
  assign n18516 = n3946 & n7242;
  assign n18517 = n18515 & ~n18516;
  assign n18518 = pi47  & ~n18517;
  assign n18519 = pi47  & ~n18518;
  assign n18520 = ~n18517 & ~n18518;
  assign n18521 = ~n18519 & ~n18520;
  assign n18522 = n18510 & ~n18521;
  assign n18523 = ~n18510 & n18521;
  assign n18524 = ~n18522 & ~n18523;
  assign n18525 = n18409 & ~n18524;
  assign n18526 = ~n18409 & n18524;
  assign n18527 = ~n18525 & ~n18526;
  assign n18528 = pi100  & n6396;
  assign n18529 = pi98  & n6735;
  assign n18530 = pi99  & n6391;
  assign n18531 = ~n18529 & ~n18530;
  assign n18532 = ~n18528 & n18531;
  assign n18533 = n4808 & n6399;
  assign n18534 = n18532 & ~n18533;
  assign n18535 = pi44  & ~n18534;
  assign n18536 = pi44  & ~n18535;
  assign n18537 = ~n18534 & ~n18535;
  assign n18538 = ~n18536 & ~n18537;
  assign n18539 = ~n18527 & ~n18538;
  assign n18540 = n18527 & n18538;
  assign n18541 = ~n18539 & ~n18540;
  assign n18542 = n18408 & ~n18541;
  assign n18543 = ~n18408 & n18541;
  assign n18544 = ~n18542 & ~n18543;
  assign n18545 = pi103  & n5636;
  assign n18546 = pi101  & n5909;
  assign n18547 = pi102  & n5631;
  assign n18548 = ~n18546 & ~n18547;
  assign n18549 = ~n18545 & n18548;
  assign n18550 = n5540 & n5639;
  assign n18551 = n18549 & ~n18550;
  assign n18552 = pi41  & ~n18551;
  assign n18553 = pi41  & ~n18552;
  assign n18554 = ~n18551 & ~n18552;
  assign n18555 = ~n18553 & ~n18554;
  assign n18556 = n18544 & ~n18555;
  assign n18557 = ~n18544 & n18555;
  assign n18558 = ~n18556 & ~n18557;
  assign n18559 = ~n18407 & n18558;
  assign n18560 = n18407 & ~n18558;
  assign n18561 = ~n18559 & ~n18560;
  assign n18562 = ~n18406 & n18561;
  assign n18563 = n18406 & ~n18561;
  assign n18564 = ~n18562 & ~n18563;
  assign n18565 = n18395 & ~n18564;
  assign n18566 = ~n18395 & n18564;
  assign n18567 = ~n18565 & ~n18566;
  assign n18568 = pi109  & n4182;
  assign n18569 = pi107  & n4416;
  assign n18570 = pi108  & n4177;
  assign n18571 = ~n18569 & ~n18570;
  assign n18572 = ~n18568 & n18571;
  assign n18573 = n4185 & n7170;
  assign n18574 = n18572 & ~n18573;
  assign n18575 = pi35  & ~n18574;
  assign n18576 = pi35  & ~n18575;
  assign n18577 = ~n18574 & ~n18575;
  assign n18578 = ~n18576 & ~n18577;
  assign n18579 = n18567 & ~n18578;
  assign n18580 = n18567 & ~n18579;
  assign n18581 = ~n18578 & ~n18579;
  assign n18582 = ~n18580 & ~n18581;
  assign n18583 = ~n18257 & ~n18260;
  assign n18584 = n18582 & n18583;
  assign n18585 = ~n18582 & ~n18583;
  assign n18586 = ~n18584 & ~n18585;
  assign n18587 = ~n18076 & ~n18264;
  assign n18588 = pi112  & n3550;
  assign n18589 = pi110  & n3735;
  assign n18590 = pi111  & n3545;
  assign n18591 = ~n18589 & ~n18590;
  assign n18592 = ~n18588 & n18591;
  assign n18593 = n3553 & n7795;
  assign n18594 = n18592 & ~n18593;
  assign n18595 = pi32  & ~n18594;
  assign n18596 = pi32  & ~n18595;
  assign n18597 = ~n18594 & ~n18595;
  assign n18598 = ~n18596 & ~n18597;
  assign n18599 = ~n18587 & ~n18598;
  assign n18600 = ~n18587 & ~n18599;
  assign n18601 = ~n18598 & ~n18599;
  assign n18602 = ~n18600 & ~n18601;
  assign n18603 = n18586 & ~n18602;
  assign n18604 = ~n18586 & n18602;
  assign n18605 = n18394 & ~n18604;
  assign n18606 = ~n18603 & n18605;
  assign n18607 = n18394 & ~n18606;
  assign n18608 = ~n18604 & ~n18606;
  assign n18609 = ~n18603 & n18608;
  assign n18610 = ~n18607 & ~n18609;
  assign n18611 = n18379 & ~n18610;
  assign n18612 = ~n18379 & n18610;
  assign n18613 = ~n18364 & ~n18612;
  assign n18614 = ~n18611 & n18613;
  assign n18615 = ~n18364 & ~n18614;
  assign n18616 = ~n18612 & ~n18614;
  assign n18617 = ~n18611 & n18616;
  assign n18618 = ~n18615 & ~n18617;
  assign n18619 = n18349 & ~n18618;
  assign n18620 = ~n18349 & n18618;
  assign n18621 = n18334 & ~n18620;
  assign n18622 = ~n18619 & n18621;
  assign n18623 = n18334 & ~n18622;
  assign n18624 = ~n18620 & ~n18622;
  assign n18625 = ~n18619 & n18624;
  assign n18626 = ~n18623 & ~n18625;
  assign n18627 = ~n18308 & ~n18311;
  assign n18628 = n18626 & n18627;
  assign n18629 = ~n18626 & ~n18627;
  assign n18630 = ~n18628 & ~n18629;
  assign n18631 = ~n18314 & ~n18317;
  assign n18632 = n18630 & ~n18631;
  assign n18633 = ~n18630 & n18631;
  assign po78  = ~n18632 & ~n18633;
  assign n18635 = ~n18348 & ~n18619;
  assign n18636 = pi126  & n1340;
  assign n18637 = pi127  & n1264;
  assign n18638 = ~n18636 & ~n18637;
  assign n18639 = ~n1272 & n18638;
  assign n18640 = ~n13389 & n18638;
  assign n18641 = ~n18639 & ~n18640;
  assign n18642 = pi17  & ~n18641;
  assign n18643 = ~pi17  & n18641;
  assign n18644 = ~n18642 & ~n18643;
  assign n18645 = ~n18635 & ~n18644;
  assign n18646 = n18635 & n18644;
  assign n18647 = ~n18645 & ~n18646;
  assign n18648 = pi125  & n1582;
  assign n18649 = pi123  & n1713;
  assign n18650 = pi124  & n1577;
  assign n18651 = ~n18649 & ~n18650;
  assign n18652 = ~n18648 & n18651;
  assign n18653 = n1585 & n12591;
  assign n18654 = n18652 & ~n18653;
  assign n18655 = pi20  & ~n18654;
  assign n18656 = pi20  & ~n18655;
  assign n18657 = ~n18654 & ~n18655;
  assign n18658 = ~n18656 & ~n18657;
  assign n18659 = ~n18350 & ~n18361;
  assign n18660 = ~n18614 & ~n18659;
  assign n18661 = n18658 & n18660;
  assign n18662 = ~n18658 & ~n18660;
  assign n18663 = ~n18661 & ~n18662;
  assign n18664 = ~n18378 & ~n18611;
  assign n18665 = pi122  & n2004;
  assign n18666 = pi120  & n2141;
  assign n18667 = pi121  & n1999;
  assign n18668 = ~n18666 & ~n18667;
  assign n18669 = ~n18665 & n18668;
  assign n18670 = ~n2007 & n18669;
  assign n18671 = ~n11463 & n18669;
  assign n18672 = ~n18670 & ~n18671;
  assign n18673 = pi23  & ~n18672;
  assign n18674 = ~pi23  & n18672;
  assign n18675 = ~n18673 & ~n18674;
  assign n18676 = ~n18664 & ~n18675;
  assign n18677 = n18664 & n18675;
  assign n18678 = ~n18676 & ~n18677;
  assign n18679 = pi119  & n2486;
  assign n18680 = pi117  & n2644;
  assign n18681 = pi118  & n2481;
  assign n18682 = ~n18680 & ~n18681;
  assign n18683 = ~n18679 & n18682;
  assign n18684 = n2489 & n10048;
  assign n18685 = n18683 & ~n18684;
  assign n18686 = pi26  & ~n18685;
  assign n18687 = pi26  & ~n18686;
  assign n18688 = ~n18685 & ~n18686;
  assign n18689 = ~n18687 & ~n18688;
  assign n18690 = ~n18393 & ~n18606;
  assign n18691 = n18689 & n18690;
  assign n18692 = ~n18689 & ~n18690;
  assign n18693 = ~n18691 & ~n18692;
  assign n18694 = pi116  & n2976;
  assign n18695 = pi114  & n3182;
  assign n18696 = pi115  & n2971;
  assign n18697 = ~n18695 & ~n18696;
  assign n18698 = ~n18694 & n18697;
  assign n18699 = n2979 & n9042;
  assign n18700 = n18698 & ~n18699;
  assign n18701 = pi29  & ~n18700;
  assign n18702 = pi29  & ~n18701;
  assign n18703 = ~n18700 & ~n18701;
  assign n18704 = ~n18702 & ~n18703;
  assign n18705 = ~n18599 & ~n18603;
  assign n18706 = ~n18704 & ~n18705;
  assign n18707 = n18704 & n18705;
  assign n18708 = ~n18706 & ~n18707;
  assign n18709 = pi113  & n3550;
  assign n18710 = pi111  & n3735;
  assign n18711 = pi112  & n3545;
  assign n18712 = ~n18710 & ~n18711;
  assign n18713 = ~n18709 & n18712;
  assign n18714 = n3553 & n8387;
  assign n18715 = n18713 & ~n18714;
  assign n18716 = pi32  & ~n18715;
  assign n18717 = pi32  & ~n18716;
  assign n18718 = ~n18715 & ~n18716;
  assign n18719 = ~n18717 & ~n18718;
  assign n18720 = ~n18579 & ~n18585;
  assign n18721 = n18719 & n18720;
  assign n18722 = ~n18719 & ~n18720;
  assign n18723 = ~n18721 & ~n18722;
  assign n18724 = ~n18562 & ~n18566;
  assign n18725 = ~n18556 & ~n18559;
  assign n18726 = pi104  & n5636;
  assign n18727 = pi102  & n5909;
  assign n18728 = pi103  & n5631;
  assign n18729 = ~n18727 & ~n18728;
  assign n18730 = ~n18726 & n18729;
  assign n18731 = n5565 & n5639;
  assign n18732 = n18730 & ~n18731;
  assign n18733 = pi41  & ~n18732;
  assign n18734 = pi41  & ~n18733;
  assign n18735 = ~n18732 & ~n18733;
  assign n18736 = ~n18734 & ~n18735;
  assign n18737 = ~n18539 & ~n18543;
  assign n18738 = pi101  & n6396;
  assign n18739 = pi99  & n6735;
  assign n18740 = pi100  & n6391;
  assign n18741 = ~n18739 & ~n18740;
  assign n18742 = ~n18738 & n18741;
  assign n18743 = n5056 & n6399;
  assign n18744 = n18742 & ~n18743;
  assign n18745 = pi44  & ~n18744;
  assign n18746 = pi44  & ~n18745;
  assign n18747 = ~n18744 & ~n18745;
  assign n18748 = ~n18746 & ~n18747;
  assign n18749 = ~n18505 & ~n18509;
  assign n18750 = pi92  & n9096;
  assign n18751 = pi90  & n9453;
  assign n18752 = pi91  & n9091;
  assign n18753 = ~n18751 & ~n18752;
  assign n18754 = ~n18750 & n18753;
  assign n18755 = n3119 & n9099;
  assign n18756 = n18754 & ~n18755;
  assign n18757 = pi53  & ~n18756;
  assign n18758 = pi53  & ~n18757;
  assign n18759 = ~n18756 & ~n18757;
  assign n18760 = ~n18758 & ~n18759;
  assign n18761 = ~n18452 & ~n18456;
  assign n18762 = ~n18435 & ~n18439;
  assign n18763 = pi79  & n13477;
  assign n18764 = pi80  & ~n13122;
  assign n18765 = ~n18763 & ~n18764;
  assign n18766 = ~n18429 & ~n18432;
  assign n18767 = ~n18765 & n18766;
  assign n18768 = n18765 & ~n18766;
  assign n18769 = ~n18767 & ~n18768;
  assign n18770 = pi83  & n12295;
  assign n18771 = pi81  & n12693;
  assign n18772 = pi82  & n12290;
  assign n18773 = ~n18771 & ~n18772;
  assign n18774 = ~n18770 & n18773;
  assign n18775 = ~n12298 & n18774;
  assign n18776 = ~n1672 & n18774;
  assign n18777 = ~n18775 & ~n18776;
  assign n18778 = pi62  & ~n18777;
  assign n18779 = ~pi62  & n18777;
  assign n18780 = ~n18778 & ~n18779;
  assign n18781 = n18769 & ~n18780;
  assign n18782 = ~n18769 & n18780;
  assign n18783 = ~n18781 & ~n18782;
  assign n18784 = ~n18762 & n18783;
  assign n18785 = n18762 & ~n18783;
  assign n18786 = ~n18784 & ~n18785;
  assign n18787 = pi86  & n11193;
  assign n18788 = pi84  & n11567;
  assign n18789 = pi85  & n11188;
  assign n18790 = ~n18788 & ~n18789;
  assign n18791 = ~n18787 & n18790;
  assign n18792 = n2099 & n11196;
  assign n18793 = n18791 & ~n18792;
  assign n18794 = pi59  & ~n18793;
  assign n18795 = pi59  & ~n18794;
  assign n18796 = ~n18793 & ~n18794;
  assign n18797 = ~n18795 & ~n18796;
  assign n18798 = n18786 & ~n18797;
  assign n18799 = ~n18786 & n18797;
  assign n18800 = ~n18798 & ~n18799;
  assign n18801 = n18761 & ~n18800;
  assign n18802 = ~n18761 & n18800;
  assign n18803 = ~n18801 & ~n18802;
  assign n18804 = pi89  & n10135;
  assign n18805 = pi87  & n10478;
  assign n18806 = pi88  & n10130;
  assign n18807 = ~n18805 & ~n18806;
  assign n18808 = ~n18804 & n18807;
  assign n18809 = n2432 & n10138;
  assign n18810 = n18808 & ~n18809;
  assign n18811 = pi56  & ~n18810;
  assign n18812 = pi56  & ~n18811;
  assign n18813 = ~n18810 & ~n18811;
  assign n18814 = ~n18812 & ~n18813;
  assign n18815 = n18803 & ~n18814;
  assign n18816 = ~n18803 & n18814;
  assign n18817 = ~n18815 & ~n18816;
  assign n18818 = ~n18474 & n18817;
  assign n18819 = n18474 & ~n18817;
  assign n18820 = ~n18818 & ~n18819;
  assign n18821 = n18760 & ~n18820;
  assign n18822 = ~n18760 & n18820;
  assign n18823 = ~n18821 & ~n18822;
  assign n18824 = ~n18488 & ~n18492;
  assign n18825 = n18823 & ~n18824;
  assign n18826 = ~n18823 & n18824;
  assign n18827 = ~n18825 & ~n18826;
  assign n18828 = pi95  & n8137;
  assign n18829 = pi93  & n8471;
  assign n18830 = pi94  & n8132;
  assign n18831 = ~n18829 & ~n18830;
  assign n18832 = ~n18828 & n18831;
  assign n18833 = n3710 & n8140;
  assign n18834 = n18832 & ~n18833;
  assign n18835 = pi50  & ~n18834;
  assign n18836 = pi50  & ~n18835;
  assign n18837 = ~n18834 & ~n18835;
  assign n18838 = ~n18836 & ~n18837;
  assign n18839 = n18827 & ~n18838;
  assign n18840 = ~n18827 & n18838;
  assign n18841 = ~n18839 & ~n18840;
  assign n18842 = n18749 & ~n18841;
  assign n18843 = ~n18749 & n18841;
  assign n18844 = ~n18842 & ~n18843;
  assign n18845 = pi98  & n7239;
  assign n18846 = pi96  & n7556;
  assign n18847 = pi97  & n7234;
  assign n18848 = ~n18846 & ~n18847;
  assign n18849 = ~n18845 & n18848;
  assign n18850 = n4360 & n7242;
  assign n18851 = n18849 & ~n18850;
  assign n18852 = pi47  & ~n18851;
  assign n18853 = pi47  & ~n18852;
  assign n18854 = ~n18851 & ~n18852;
  assign n18855 = ~n18853 & ~n18854;
  assign n18856 = ~n18844 & n18855;
  assign n18857 = n18844 & ~n18855;
  assign n18858 = ~n18856 & ~n18857;
  assign n18859 = ~n18523 & ~n18526;
  assign n18860 = n18858 & n18859;
  assign n18861 = ~n18858 & ~n18859;
  assign n18862 = ~n18860 & ~n18861;
  assign n18863 = ~n18748 & n18862;
  assign n18864 = n18748 & ~n18862;
  assign n18865 = ~n18863 & ~n18864;
  assign n18866 = ~n18737 & n18865;
  assign n18867 = n18737 & ~n18865;
  assign n18868 = ~n18866 & ~n18867;
  assign n18869 = ~n18736 & n18868;
  assign n18870 = n18736 & ~n18868;
  assign n18871 = ~n18869 & ~n18870;
  assign n18872 = ~n18725 & n18871;
  assign n18873 = n18725 & ~n18871;
  assign n18874 = ~n18872 & ~n18873;
  assign n18875 = pi107  & n4896;
  assign n18876 = pi105  & n5148;
  assign n18877 = pi106  & n4891;
  assign n18878 = ~n18876 & ~n18877;
  assign n18879 = ~n18875 & n18878;
  assign n18880 = n4899 & n6614;
  assign n18881 = n18879 & ~n18880;
  assign n18882 = pi38  & ~n18881;
  assign n18883 = pi38  & ~n18882;
  assign n18884 = ~n18881 & ~n18882;
  assign n18885 = ~n18883 & ~n18884;
  assign n18886 = n18874 & ~n18885;
  assign n18887 = ~n18874 & n18885;
  assign n18888 = ~n18886 & ~n18887;
  assign n18889 = n18724 & ~n18888;
  assign n18890 = ~n18724 & n18888;
  assign n18891 = ~n18889 & ~n18890;
  assign n18892 = pi110  & n4182;
  assign n18893 = pi108  & n4416;
  assign n18894 = pi109  & n4177;
  assign n18895 = ~n18893 & ~n18894;
  assign n18896 = ~n18892 & n18895;
  assign n18897 = n4185 & n7474;
  assign n18898 = n18896 & ~n18897;
  assign n18899 = pi35  & ~n18898;
  assign n18900 = pi35  & ~n18899;
  assign n18901 = ~n18898 & ~n18899;
  assign n18902 = ~n18900 & ~n18901;
  assign n18903 = n18891 & ~n18902;
  assign n18904 = ~n18891 & n18902;
  assign n18905 = ~n18903 & ~n18904;
  assign n18906 = n18723 & n18905;
  assign n18907 = ~n18723 & ~n18905;
  assign n18908 = n18708 & ~n18907;
  assign n18909 = ~n18906 & n18908;
  assign n18910 = n18708 & ~n18909;
  assign n18911 = ~n18907 & ~n18909;
  assign n18912 = ~n18906 & n18911;
  assign n18913 = ~n18910 & ~n18912;
  assign n18914 = n18693 & ~n18913;
  assign n18915 = ~n18693 & n18913;
  assign n18916 = n18678 & ~n18915;
  assign n18917 = ~n18914 & n18916;
  assign n18918 = n18678 & ~n18917;
  assign n18919 = ~n18915 & ~n18917;
  assign n18920 = ~n18914 & n18919;
  assign n18921 = ~n18918 & ~n18920;
  assign n18922 = n18663 & ~n18921;
  assign n18923 = ~n18663 & n18921;
  assign n18924 = n18647 & ~n18923;
  assign n18925 = ~n18922 & n18924;
  assign n18926 = n18647 & ~n18925;
  assign n18927 = ~n18923 & ~n18925;
  assign n18928 = ~n18922 & n18927;
  assign n18929 = ~n18926 & ~n18928;
  assign n18930 = ~n18332 & ~n18622;
  assign n18931 = n18929 & n18930;
  assign n18932 = ~n18929 & ~n18930;
  assign n18933 = ~n18931 & ~n18932;
  assign n18934 = ~n18629 & ~n18632;
  assign n18935 = n18933 & ~n18934;
  assign n18936 = ~n18933 & n18934;
  assign po79  = ~n18935 & ~n18936;
  assign n18938 = ~n18932 & ~n18935;
  assign n18939 = ~n18645 & ~n18925;
  assign n18940 = pi126  & n1582;
  assign n18941 = pi124  & n1713;
  assign n18942 = pi125  & n1577;
  assign n18943 = ~n18941 & ~n18942;
  assign n18944 = ~n18940 & n18943;
  assign n18945 = n1585 & n12979;
  assign n18946 = n18944 & ~n18945;
  assign n18947 = pi20  & ~n18946;
  assign n18948 = pi20  & ~n18947;
  assign n18949 = ~n18946 & ~n18947;
  assign n18950 = ~n18948 & ~n18949;
  assign n18951 = ~n18676 & ~n18917;
  assign n18952 = n18950 & n18951;
  assign n18953 = ~n18950 & ~n18951;
  assign n18954 = ~n18952 & ~n18953;
  assign n18955 = pi123  & n2004;
  assign n18956 = pi121  & n2141;
  assign n18957 = pi122  & n1999;
  assign n18958 = ~n18956 & ~n18957;
  assign n18959 = ~n18955 & n18958;
  assign n18960 = n2007 & n11489;
  assign n18961 = n18959 & ~n18960;
  assign n18962 = pi23  & ~n18961;
  assign n18963 = pi23  & ~n18962;
  assign n18964 = ~n18961 & ~n18962;
  assign n18965 = ~n18963 & ~n18964;
  assign n18966 = ~n18692 & ~n18914;
  assign n18967 = ~n18965 & ~n18966;
  assign n18968 = n18965 & n18966;
  assign n18969 = ~n18967 & ~n18968;
  assign n18970 = pi120  & n2486;
  assign n18971 = pi118  & n2644;
  assign n18972 = pi119  & n2481;
  assign n18973 = ~n18971 & ~n18972;
  assign n18974 = ~n18970 & n18973;
  assign n18975 = n2489 & n10734;
  assign n18976 = n18974 & ~n18975;
  assign n18977 = pi26  & ~n18976;
  assign n18978 = pi26  & ~n18977;
  assign n18979 = ~n18976 & ~n18977;
  assign n18980 = ~n18978 & ~n18979;
  assign n18981 = ~n18706 & ~n18909;
  assign n18982 = n18980 & n18981;
  assign n18983 = ~n18980 & ~n18981;
  assign n18984 = ~n18982 & ~n18983;
  assign n18985 = pi117  & n2976;
  assign n18986 = pi115  & n3182;
  assign n18987 = pi116  & n2971;
  assign n18988 = ~n18986 & ~n18987;
  assign n18989 = ~n18985 & n18988;
  assign n18990 = n2979 & n9691;
  assign n18991 = n18989 & ~n18990;
  assign n18992 = pi29  & ~n18991;
  assign n18993 = pi29  & ~n18992;
  assign n18994 = ~n18991 & ~n18992;
  assign n18995 = ~n18993 & ~n18994;
  assign n18996 = ~n18722 & ~n18906;
  assign n18997 = ~n18995 & ~n18996;
  assign n18998 = n18995 & n18996;
  assign n18999 = ~n18997 & ~n18998;
  assign n19000 = pi114  & n3550;
  assign n19001 = pi112  & n3735;
  assign n19002 = pi113  & n3545;
  assign n19003 = ~n19001 & ~n19002;
  assign n19004 = ~n19000 & n19003;
  assign n19005 = n3553 & n8702;
  assign n19006 = n19004 & ~n19005;
  assign n19007 = pi32  & ~n19006;
  assign n19008 = pi32  & ~n19007;
  assign n19009 = ~n19006 & ~n19007;
  assign n19010 = ~n19008 & ~n19009;
  assign n19011 = ~n18890 & ~n18903;
  assign n19012 = n19010 & n19011;
  assign n19013 = ~n19010 & ~n19011;
  assign n19014 = ~n19012 & ~n19013;
  assign n19015 = ~n18872 & ~n18886;
  assign n19016 = pi108  & n4896;
  assign n19017 = pi106  & n5148;
  assign n19018 = pi107  & n4891;
  assign n19019 = ~n19017 & ~n19018;
  assign n19020 = ~n19016 & n19019;
  assign n19021 = n4899 & n6639;
  assign n19022 = n19020 & ~n19021;
  assign n19023 = pi38  & ~n19022;
  assign n19024 = pi38  & ~n19023;
  assign n19025 = ~n19022 & ~n19023;
  assign n19026 = ~n19024 & ~n19025;
  assign n19027 = ~n18866 & ~n18869;
  assign n19028 = pi105  & n5636;
  assign n19029 = pi103  & n5909;
  assign n19030 = pi104  & n5631;
  assign n19031 = ~n19029 & ~n19030;
  assign n19032 = ~n19028 & n19031;
  assign n19033 = n5639 & n6065;
  assign n19034 = n19032 & ~n19033;
  assign n19035 = pi41  & ~n19034;
  assign n19036 = pi41  & ~n19035;
  assign n19037 = ~n19034 & ~n19035;
  assign n19038 = ~n19036 & ~n19037;
  assign n19039 = ~n18860 & ~n18863;
  assign n19040 = pi102  & n6396;
  assign n19041 = pi100  & n6735;
  assign n19042 = pi101  & n6391;
  assign n19043 = ~n19041 & ~n19042;
  assign n19044 = ~n19040 & n19043;
  assign n19045 = n5296 & n6399;
  assign n19046 = n19044 & ~n19045;
  assign n19047 = pi44  & ~n19046;
  assign n19048 = pi44  & ~n19047;
  assign n19049 = ~n19046 & ~n19047;
  assign n19050 = ~n19048 & ~n19049;
  assign n19051 = ~n18843 & ~n18857;
  assign n19052 = pi96  & n8137;
  assign n19053 = pi94  & n8471;
  assign n19054 = pi95  & n8132;
  assign n19055 = ~n19053 & ~n19054;
  assign n19056 = ~n19052 & n19055;
  assign n19057 = n3921 & n8140;
  assign n19058 = n19056 & ~n19057;
  assign n19059 = pi50  & ~n19058;
  assign n19060 = pi50  & ~n19059;
  assign n19061 = ~n19058 & ~n19059;
  assign n19062 = ~n19060 & ~n19061;
  assign n19063 = ~n18818 & ~n18822;
  assign n19064 = ~n18802 & ~n18815;
  assign n19065 = pi90  & n10135;
  assign n19066 = pi88  & n10478;
  assign n19067 = pi89  & n10130;
  assign n19068 = ~n19066 & ~n19067;
  assign n19069 = ~n19065 & n19068;
  assign n19070 = n2606 & n10138;
  assign n19071 = n19069 & ~n19070;
  assign n19072 = pi56  & ~n19071;
  assign n19073 = pi56  & ~n19072;
  assign n19074 = ~n19071 & ~n19072;
  assign n19075 = ~n19073 & ~n19074;
  assign n19076 = ~n18784 & ~n18798;
  assign n19077 = pi84  & n12295;
  assign n19078 = pi82  & n12693;
  assign n19079 = pi83  & n12290;
  assign n19080 = ~n19078 & ~n19079;
  assign n19081 = ~n19077 & n19080;
  assign n19082 = n1805 & n12298;
  assign n19083 = n19081 & ~n19082;
  assign n19084 = pi62  & ~n19083;
  assign n19085 = pi62  & ~n19084;
  assign n19086 = ~n19083 & ~n19084;
  assign n19087 = ~n19085 & ~n19086;
  assign n19088 = pi80  & n13477;
  assign n19089 = pi81  & ~n13122;
  assign n19090 = ~n19088 & ~n19089;
  assign n19091 = n18765 & ~n19090;
  assign n19092 = ~n18765 & n19090;
  assign n19093 = ~n19087 & ~n19092;
  assign n19094 = ~n19091 & n19093;
  assign n19095 = ~n19087 & ~n19094;
  assign n19096 = ~n19092 & ~n19094;
  assign n19097 = ~n19091 & n19096;
  assign n19098 = ~n19095 & ~n19097;
  assign n19099 = ~n18768 & ~n18781;
  assign n19100 = n19098 & n19099;
  assign n19101 = ~n19098 & ~n19099;
  assign n19102 = ~n19100 & ~n19101;
  assign n19103 = pi87  & n11193;
  assign n19104 = pi85  & n11567;
  assign n19105 = pi86  & n11188;
  assign n19106 = ~n19104 & ~n19105;
  assign n19107 = ~n19103 & n19106;
  assign n19108 = n2252 & n11196;
  assign n19109 = n19107 & ~n19108;
  assign n19110 = pi59  & ~n19109;
  assign n19111 = pi59  & ~n19110;
  assign n19112 = ~n19109 & ~n19110;
  assign n19113 = ~n19111 & ~n19112;
  assign n19114 = ~n19102 & n19113;
  assign n19115 = n19102 & ~n19113;
  assign n19116 = ~n19114 & ~n19115;
  assign n19117 = ~n19076 & n19116;
  assign n19118 = n19076 & ~n19116;
  assign n19119 = ~n19117 & ~n19118;
  assign n19120 = ~n19075 & n19119;
  assign n19121 = n19075 & ~n19119;
  assign n19122 = ~n19120 & ~n19121;
  assign n19123 = ~n19064 & n19122;
  assign n19124 = n19064 & ~n19122;
  assign n19125 = ~n19123 & ~n19124;
  assign n19126 = pi93  & n9096;
  assign n19127 = pi91  & n9453;
  assign n19128 = pi92  & n9091;
  assign n19129 = ~n19127 & ~n19128;
  assign n19130 = ~n19126 & n19129;
  assign n19131 = n3144 & n9099;
  assign n19132 = n19130 & ~n19131;
  assign n19133 = pi53  & ~n19132;
  assign n19134 = pi53  & ~n19133;
  assign n19135 = ~n19132 & ~n19133;
  assign n19136 = ~n19134 & ~n19135;
  assign n19137 = n19125 & ~n19136;
  assign n19138 = ~n19125 & n19136;
  assign n19139 = ~n19137 & ~n19138;
  assign n19140 = ~n19063 & n19139;
  assign n19141 = n19063 & ~n19139;
  assign n19142 = ~n19140 & ~n19141;
  assign n19143 = n19062 & n19142;
  assign n19144 = ~n19062 & ~n19142;
  assign n19145 = ~n19143 & ~n19144;
  assign n19146 = ~n18825 & ~n18839;
  assign n19147 = n19145 & n19146;
  assign n19148 = ~n19145 & ~n19146;
  assign n19149 = ~n19147 & ~n19148;
  assign n19150 = pi99  & n7239;
  assign n19151 = pi97  & n7556;
  assign n19152 = pi98  & n7234;
  assign n19153 = ~n19151 & ~n19152;
  assign n19154 = ~n19150 & n19153;
  assign n19155 = n4584 & n7242;
  assign n19156 = n19154 & ~n19155;
  assign n19157 = pi47  & ~n19156;
  assign n19158 = pi47  & ~n19157;
  assign n19159 = ~n19156 & ~n19157;
  assign n19160 = ~n19158 & ~n19159;
  assign n19161 = n19149 & ~n19160;
  assign n19162 = ~n19149 & n19160;
  assign n19163 = ~n19161 & ~n19162;
  assign n19164 = ~n19051 & n19163;
  assign n19165 = n19051 & ~n19163;
  assign n19166 = ~n19164 & ~n19165;
  assign n19167 = n19050 & n19166;
  assign n19168 = ~n19050 & ~n19166;
  assign n19169 = ~n19167 & ~n19168;
  assign n19170 = ~n19039 & ~n19169;
  assign n19171 = n19039 & n19169;
  assign n19172 = ~n19170 & ~n19171;
  assign n19173 = ~n19038 & n19172;
  assign n19174 = n19038 & ~n19172;
  assign n19175 = ~n19173 & ~n19174;
  assign n19176 = ~n19027 & n19175;
  assign n19177 = n19027 & ~n19175;
  assign n19178 = ~n19176 & ~n19177;
  assign n19179 = ~n19026 & n19178;
  assign n19180 = n19026 & ~n19178;
  assign n19181 = ~n19179 & ~n19180;
  assign n19182 = ~n19015 & n19181;
  assign n19183 = n19015 & ~n19181;
  assign n19184 = ~n19182 & ~n19183;
  assign n19185 = pi111  & n4182;
  assign n19186 = pi109  & n4416;
  assign n19187 = pi110  & n4177;
  assign n19188 = ~n19186 & ~n19187;
  assign n19189 = ~n19185 & n19188;
  assign n19190 = n4185 & n7770;
  assign n19191 = n19189 & ~n19190;
  assign n19192 = pi35  & ~n19191;
  assign n19193 = pi35  & ~n19192;
  assign n19194 = ~n19191 & ~n19192;
  assign n19195 = ~n19193 & ~n19194;
  assign n19196 = n19184 & ~n19195;
  assign n19197 = n19184 & ~n19196;
  assign n19198 = ~n19195 & ~n19196;
  assign n19199 = ~n19197 & ~n19198;
  assign n19200 = n19014 & ~n19199;
  assign n19201 = ~n19014 & n19199;
  assign n19202 = n18999 & ~n19201;
  assign n19203 = ~n19200 & n19202;
  assign n19204 = n18999 & ~n19203;
  assign n19205 = ~n19201 & ~n19203;
  assign n19206 = ~n19200 & n19205;
  assign n19207 = ~n19204 & ~n19206;
  assign n19208 = n18984 & ~n19207;
  assign n19209 = ~n18984 & n19207;
  assign n19210 = n18969 & ~n19209;
  assign n19211 = ~n19208 & n19210;
  assign n19212 = n18969 & ~n19211;
  assign n19213 = ~n19209 & ~n19211;
  assign n19214 = ~n19208 & n19213;
  assign n19215 = ~n19212 & ~n19214;
  assign n19216 = ~n18954 & n19215;
  assign n19217 = n18954 & ~n19215;
  assign n19218 = ~n19216 & ~n19217;
  assign n19219 = ~n18662 & ~n18922;
  assign n19220 = pi127  & n1340;
  assign n19221 = n1272 & n13387;
  assign n19222 = ~n19220 & ~n19221;
  assign n19223 = pi17  & ~n19222;
  assign n19224 = pi17  & ~n19223;
  assign n19225 = ~n19222 & ~n19223;
  assign n19226 = ~n19224 & ~n19225;
  assign n19227 = ~n19219 & ~n19226;
  assign n19228 = n19219 & n19226;
  assign n19229 = ~n19227 & ~n19228;
  assign n19230 = n19218 & n19229;
  assign n19231 = ~n19218 & ~n19229;
  assign n19232 = ~n19230 & ~n19231;
  assign n19233 = ~n18939 & n19232;
  assign n19234 = n18939 & ~n19232;
  assign n19235 = ~n19233 & ~n19234;
  assign n19236 = ~n18938 & n19235;
  assign n19237 = n18938 & ~n19235;
  assign po80  = ~n19236 & ~n19237;
  assign n19239 = ~n19233 & ~n19236;
  assign n19240 = ~n19227 & ~n19230;
  assign n19241 = ~n18953 & ~n19217;
  assign n19242 = pi127  & n1582;
  assign n19243 = pi125  & n1713;
  assign n19244 = pi126  & n1577;
  assign n19245 = ~n19243 & ~n19244;
  assign n19246 = ~n19242 & n19245;
  assign n19247 = n1585 & n13365;
  assign n19248 = n19246 & ~n19247;
  assign n19249 = pi20  & ~n19248;
  assign n19250 = pi20  & ~n19249;
  assign n19251 = ~n19248 & ~n19249;
  assign n19252 = ~n19250 & ~n19251;
  assign n19253 = ~n19241 & ~n19252;
  assign n19254 = n19241 & n19252;
  assign n19255 = ~n19253 & ~n19254;
  assign n19256 = pi124  & n2004;
  assign n19257 = pi122  & n2141;
  assign n19258 = pi123  & n1999;
  assign n19259 = ~n19257 & ~n19258;
  assign n19260 = ~n19256 & n19259;
  assign n19261 = n2007 & n11858;
  assign n19262 = n19260 & ~n19261;
  assign n19263 = pi23  & ~n19262;
  assign n19264 = pi23  & ~n19263;
  assign n19265 = ~n19262 & ~n19263;
  assign n19266 = ~n19264 & ~n19265;
  assign n19267 = ~n18967 & ~n19211;
  assign n19268 = n19266 & n19267;
  assign n19269 = ~n19266 & ~n19267;
  assign n19270 = ~n19268 & ~n19269;
  assign n19271 = pi121  & n2486;
  assign n19272 = pi119  & n2644;
  assign n19273 = pi120  & n2481;
  assign n19274 = ~n19272 & ~n19273;
  assign n19275 = ~n19271 & n19274;
  assign n19276 = n2489 & n11086;
  assign n19277 = n19275 & ~n19276;
  assign n19278 = pi26  & ~n19277;
  assign n19279 = pi26  & ~n19278;
  assign n19280 = ~n19277 & ~n19278;
  assign n19281 = ~n19279 & ~n19280;
  assign n19282 = ~n18983 & ~n19208;
  assign n19283 = ~n19281 & ~n19282;
  assign n19284 = n19281 & n19282;
  assign n19285 = ~n19283 & ~n19284;
  assign n19286 = pi118  & n2976;
  assign n19287 = pi116  & n3182;
  assign n19288 = pi117  & n2971;
  assign n19289 = ~n19287 & ~n19288;
  assign n19290 = ~n19286 & n19289;
  assign n19291 = n2979 & n9716;
  assign n19292 = n19290 & ~n19291;
  assign n19293 = pi29  & ~n19292;
  assign n19294 = pi29  & ~n19293;
  assign n19295 = ~n19292 & ~n19293;
  assign n19296 = ~n19294 & ~n19295;
  assign n19297 = ~n18997 & ~n19203;
  assign n19298 = n19296 & n19297;
  assign n19299 = ~n19296 & ~n19297;
  assign n19300 = ~n19298 & ~n19299;
  assign n19301 = ~n19182 & ~n19196;
  assign n19302 = ~n19170 & ~n19173;
  assign n19303 = pi106  & n5636;
  assign n19304 = pi104  & n5909;
  assign n19305 = pi105  & n5631;
  assign n19306 = ~n19304 & ~n19305;
  assign n19307 = ~n19303 & n19306;
  assign n19308 = n5639 & n6090;
  assign n19309 = n19307 & ~n19308;
  assign n19310 = pi41  & ~n19309;
  assign n19311 = pi41  & ~n19310;
  assign n19312 = ~n19309 & ~n19310;
  assign n19313 = ~n19311 & ~n19312;
  assign n19314 = ~n19165 & ~n19167;
  assign n19315 = ~n19148 & ~n19161;
  assign n19316 = ~n19123 & ~n19137;
  assign n19317 = ~n19101 & ~n19115;
  assign n19318 = pi88  & n11193;
  assign n19319 = pi86  & n11567;
  assign n19320 = pi87  & n11188;
  assign n19321 = ~n19319 & ~n19320;
  assign n19322 = ~n19318 & n19321;
  assign n19323 = n2277 & n11196;
  assign n19324 = n19322 & ~n19323;
  assign n19325 = pi59  & ~n19324;
  assign n19326 = pi59  & ~n19325;
  assign n19327 = ~n19324 & ~n19325;
  assign n19328 = ~n19326 & ~n19327;
  assign n19329 = pi85  & n12295;
  assign n19330 = pi83  & n12693;
  assign n19331 = pi84  & n12290;
  assign n19332 = ~n19330 & ~n19331;
  assign n19333 = ~n19329 & n19332;
  assign n19334 = n1943 & n12298;
  assign n19335 = n19333 & ~n19334;
  assign n19336 = pi62  & ~n19335;
  assign n19337 = pi62  & ~n19336;
  assign n19338 = ~n19335 & ~n19336;
  assign n19339 = ~n19337 & ~n19338;
  assign n19340 = pi81  & n13477;
  assign n19341 = pi82  & ~n13122;
  assign n19342 = ~n19340 & ~n19341;
  assign n19343 = ~pi17  & ~n19342;
  assign n19344 = pi17  & n19342;
  assign n19345 = ~n19343 & ~n19344;
  assign n19346 = ~n19090 & n19345;
  assign n19347 = n19090 & ~n19345;
  assign n19348 = ~n19346 & ~n19347;
  assign n19349 = ~n19339 & n19348;
  assign n19350 = n19339 & ~n19348;
  assign n19351 = ~n19349 & ~n19350;
  assign n19352 = ~n19096 & n19351;
  assign n19353 = n19096 & ~n19351;
  assign n19354 = ~n19352 & ~n19353;
  assign n19355 = n19328 & ~n19354;
  assign n19356 = ~n19328 & n19354;
  assign n19357 = ~n19355 & ~n19356;
  assign n19358 = ~n19317 & n19357;
  assign n19359 = n19317 & ~n19357;
  assign n19360 = ~n19358 & ~n19359;
  assign n19361 = pi91  & n10135;
  assign n19362 = pi89  & n10478;
  assign n19363 = pi90  & n10130;
  assign n19364 = ~n19362 & ~n19363;
  assign n19365 = ~n19361 & n19364;
  assign n19366 = n2926 & n10138;
  assign n19367 = n19365 & ~n19366;
  assign n19368 = pi56  & ~n19367;
  assign n19369 = pi56  & ~n19368;
  assign n19370 = ~n19367 & ~n19368;
  assign n19371 = ~n19369 & ~n19370;
  assign n19372 = n19360 & ~n19371;
  assign n19373 = n19360 & ~n19372;
  assign n19374 = ~n19371 & ~n19372;
  assign n19375 = ~n19373 & ~n19374;
  assign n19376 = ~n19117 & ~n19120;
  assign n19377 = n19375 & n19376;
  assign n19378 = ~n19375 & ~n19376;
  assign n19379 = ~n19377 & ~n19378;
  assign n19380 = pi94  & n9096;
  assign n19381 = pi92  & n9453;
  assign n19382 = pi93  & n9091;
  assign n19383 = ~n19381 & ~n19382;
  assign n19384 = ~n19380 & n19383;
  assign n19385 = n3499 & n9099;
  assign n19386 = n19384 & ~n19385;
  assign n19387 = pi53  & ~n19386;
  assign n19388 = pi53  & ~n19387;
  assign n19389 = ~n19386 & ~n19387;
  assign n19390 = ~n19388 & ~n19389;
  assign n19391 = n19379 & ~n19390;
  assign n19392 = ~n19379 & n19390;
  assign n19393 = ~n19391 & ~n19392;
  assign n19394 = n19316 & ~n19393;
  assign n19395 = ~n19316 & n19393;
  assign n19396 = ~n19394 & ~n19395;
  assign n19397 = pi97  & n8137;
  assign n19398 = pi95  & n8471;
  assign n19399 = pi96  & n8132;
  assign n19400 = ~n19398 & ~n19399;
  assign n19401 = ~n19397 & n19400;
  assign n19402 = n3946 & n8140;
  assign n19403 = n19401 & ~n19402;
  assign n19404 = pi50  & ~n19403;
  assign n19405 = pi50  & ~n19404;
  assign n19406 = ~n19403 & ~n19404;
  assign n19407 = ~n19405 & ~n19406;
  assign n19408 = ~n19141 & ~n19143;
  assign n19409 = ~n19407 & n19408;
  assign n19410 = n19407 & ~n19408;
  assign n19411 = ~n19409 & ~n19410;
  assign n19412 = ~n19396 & n19411;
  assign n19413 = n19396 & ~n19411;
  assign n19414 = ~n19412 & ~n19413;
  assign n19415 = pi100  & n7239;
  assign n19416 = pi98  & n7556;
  assign n19417 = pi99  & n7234;
  assign n19418 = ~n19416 & ~n19417;
  assign n19419 = ~n19415 & n19418;
  assign n19420 = n4808 & n7242;
  assign n19421 = n19419 & ~n19420;
  assign n19422 = pi47  & ~n19421;
  assign n19423 = pi47  & ~n19422;
  assign n19424 = ~n19421 & ~n19422;
  assign n19425 = ~n19423 & ~n19424;
  assign n19426 = ~n19414 & ~n19425;
  assign n19427 = n19414 & n19425;
  assign n19428 = ~n19426 & ~n19427;
  assign n19429 = n19315 & ~n19428;
  assign n19430 = ~n19315 & n19428;
  assign n19431 = ~n19429 & ~n19430;
  assign n19432 = pi103  & n6396;
  assign n19433 = pi101  & n6735;
  assign n19434 = pi102  & n6391;
  assign n19435 = ~n19433 & ~n19434;
  assign n19436 = ~n19432 & n19435;
  assign n19437 = n5540 & n6399;
  assign n19438 = n19436 & ~n19437;
  assign n19439 = pi44  & ~n19438;
  assign n19440 = pi44  & ~n19439;
  assign n19441 = ~n19438 & ~n19439;
  assign n19442 = ~n19440 & ~n19441;
  assign n19443 = n19431 & ~n19442;
  assign n19444 = ~n19431 & n19442;
  assign n19445 = ~n19443 & ~n19444;
  assign n19446 = n19314 & n19445;
  assign n19447 = ~n19314 & ~n19445;
  assign n19448 = ~n19446 & ~n19447;
  assign n19449 = ~n19313 & n19448;
  assign n19450 = n19313 & ~n19448;
  assign n19451 = ~n19449 & ~n19450;
  assign n19452 = n19302 & ~n19451;
  assign n19453 = ~n19302 & n19451;
  assign n19454 = ~n19452 & ~n19453;
  assign n19455 = pi109  & n4896;
  assign n19456 = pi107  & n5148;
  assign n19457 = pi108  & n4891;
  assign n19458 = ~n19456 & ~n19457;
  assign n19459 = ~n19455 & n19458;
  assign n19460 = n4899 & n7170;
  assign n19461 = n19459 & ~n19460;
  assign n19462 = pi38  & ~n19461;
  assign n19463 = pi38  & ~n19462;
  assign n19464 = ~n19461 & ~n19462;
  assign n19465 = ~n19463 & ~n19464;
  assign n19466 = n19454 & ~n19465;
  assign n19467 = n19454 & ~n19466;
  assign n19468 = ~n19465 & ~n19466;
  assign n19469 = ~n19467 & ~n19468;
  assign n19470 = ~n19176 & ~n19179;
  assign n19471 = n19469 & n19470;
  assign n19472 = ~n19469 & ~n19470;
  assign n19473 = ~n19471 & ~n19472;
  assign n19474 = pi112  & n4182;
  assign n19475 = pi110  & n4416;
  assign n19476 = pi111  & n4177;
  assign n19477 = ~n19475 & ~n19476;
  assign n19478 = ~n19474 & n19477;
  assign n19479 = n4185 & n7795;
  assign n19480 = n19478 & ~n19479;
  assign n19481 = pi35  & ~n19480;
  assign n19482 = pi35  & ~n19481;
  assign n19483 = ~n19480 & ~n19481;
  assign n19484 = ~n19482 & ~n19483;
  assign n19485 = n19473 & ~n19484;
  assign n19486 = ~n19473 & n19484;
  assign n19487 = ~n19485 & ~n19486;
  assign n19488 = n19301 & ~n19487;
  assign n19489 = ~n19301 & n19487;
  assign n19490 = ~n19488 & ~n19489;
  assign n19491 = pi115  & n3550;
  assign n19492 = pi113  & n3735;
  assign n19493 = pi114  & n3545;
  assign n19494 = ~n19492 & ~n19493;
  assign n19495 = ~n19491 & n19494;
  assign n19496 = n3553 & n8727;
  assign n19497 = n19495 & ~n19496;
  assign n19498 = pi32  & ~n19497;
  assign n19499 = pi32  & ~n19498;
  assign n19500 = ~n19497 & ~n19498;
  assign n19501 = ~n19499 & ~n19500;
  assign n19502 = ~n19013 & ~n19200;
  assign n19503 = ~n19501 & ~n19502;
  assign n19504 = n19501 & n19502;
  assign n19505 = ~n19503 & ~n19504;
  assign n19506 = n19490 & n19505;
  assign n19507 = ~n19490 & ~n19505;
  assign n19508 = ~n19506 & ~n19507;
  assign n19509 = n19300 & n19508;
  assign n19510 = ~n19300 & ~n19508;
  assign n19511 = ~n19509 & ~n19510;
  assign n19512 = n19285 & n19511;
  assign n19513 = ~n19285 & ~n19511;
  assign n19514 = ~n19512 & ~n19513;
  assign n19515 = n19270 & n19514;
  assign n19516 = ~n19270 & ~n19514;
  assign n19517 = ~n19515 & ~n19516;
  assign n19518 = n19255 & n19517;
  assign n19519 = ~n19255 & ~n19517;
  assign n19520 = ~n19518 & ~n19519;
  assign n19521 = ~n19240 & n19520;
  assign n19522 = n19240 & ~n19520;
  assign n19523 = ~n19521 & ~n19522;
  assign n19524 = ~n19239 & n19523;
  assign n19525 = n19239 & ~n19523;
  assign po81  = ~n19524 & ~n19525;
  assign n19527 = ~n19521 & ~n19524;
  assign n19528 = ~n19253 & ~n19518;
  assign n19529 = pi125  & n2004;
  assign n19530 = pi123  & n2141;
  assign n19531 = pi124  & n1999;
  assign n19532 = ~n19530 & ~n19531;
  assign n19533 = ~n19529 & n19532;
  assign n19534 = n2007 & n12591;
  assign n19535 = n19533 & ~n19534;
  assign n19536 = pi23  & ~n19535;
  assign n19537 = pi23  & ~n19536;
  assign n19538 = ~n19535 & ~n19536;
  assign n19539 = ~n19537 & ~n19538;
  assign n19540 = ~n19283 & ~n19512;
  assign n19541 = n19539 & n19540;
  assign n19542 = ~n19539 & ~n19540;
  assign n19543 = ~n19541 & ~n19542;
  assign n19544 = pi122  & n2486;
  assign n19545 = pi120  & n2644;
  assign n19546 = pi121  & n2481;
  assign n19547 = ~n19545 & ~n19546;
  assign n19548 = ~n19544 & n19547;
  assign n19549 = n2489 & n11463;
  assign n19550 = n19548 & ~n19549;
  assign n19551 = pi26  & ~n19550;
  assign n19552 = pi26  & ~n19551;
  assign n19553 = ~n19550 & ~n19551;
  assign n19554 = ~n19552 & ~n19553;
  assign n19555 = ~n19299 & ~n19509;
  assign n19556 = n19554 & n19555;
  assign n19557 = ~n19554 & ~n19555;
  assign n19558 = ~n19556 & ~n19557;
  assign n19559 = pi119  & n2976;
  assign n19560 = pi117  & n3182;
  assign n19561 = pi118  & n2971;
  assign n19562 = ~n19560 & ~n19561;
  assign n19563 = ~n19559 & n19562;
  assign n19564 = n2979 & n10048;
  assign n19565 = n19563 & ~n19564;
  assign n19566 = pi29  & ~n19565;
  assign n19567 = pi29  & ~n19566;
  assign n19568 = ~n19565 & ~n19566;
  assign n19569 = ~n19567 & ~n19568;
  assign n19570 = ~n19503 & ~n19506;
  assign n19571 = n19569 & n19570;
  assign n19572 = ~n19569 & ~n19570;
  assign n19573 = ~n19571 & ~n19572;
  assign n19574 = pi116  & n3550;
  assign n19575 = pi114  & n3735;
  assign n19576 = pi115  & n3545;
  assign n19577 = ~n19575 & ~n19576;
  assign n19578 = ~n19574 & n19577;
  assign n19579 = n3553 & n9042;
  assign n19580 = n19578 & ~n19579;
  assign n19581 = pi32  & ~n19580;
  assign n19582 = pi32  & ~n19581;
  assign n19583 = ~n19580 & ~n19581;
  assign n19584 = ~n19582 & ~n19583;
  assign n19585 = ~n19485 & ~n19489;
  assign n19586 = n19584 & n19585;
  assign n19587 = ~n19584 & ~n19585;
  assign n19588 = ~n19586 & ~n19587;
  assign n19589 = ~n19466 & ~n19472;
  assign n19590 = ~n19449 & ~n19453;
  assign n19591 = ~n19443 & ~n19446;
  assign n19592 = pi104  & n6396;
  assign n19593 = pi102  & n6735;
  assign n19594 = pi103  & n6391;
  assign n19595 = ~n19593 & ~n19594;
  assign n19596 = ~n19592 & n19595;
  assign n19597 = n5565 & n6399;
  assign n19598 = n19596 & ~n19597;
  assign n19599 = pi44  & ~n19598;
  assign n19600 = pi44  & ~n19599;
  assign n19601 = ~n19598 & ~n19599;
  assign n19602 = ~n19600 & ~n19601;
  assign n19603 = ~n19426 & ~n19430;
  assign n19604 = ~n19391 & ~n19395;
  assign n19605 = pi92  & n10135;
  assign n19606 = pi90  & n10478;
  assign n19607 = pi91  & n10130;
  assign n19608 = ~n19606 & ~n19607;
  assign n19609 = ~n19605 & n19608;
  assign n19610 = n3119 & n10138;
  assign n19611 = n19609 & ~n19610;
  assign n19612 = pi56  & ~n19611;
  assign n19613 = pi56  & ~n19612;
  assign n19614 = ~n19611 & ~n19612;
  assign n19615 = ~n19613 & ~n19614;
  assign n19616 = ~n19356 & ~n19358;
  assign n19617 = pi82  & n13477;
  assign n19618 = pi83  & ~n13122;
  assign n19619 = ~n19617 & ~n19618;
  assign n19620 = ~n19343 & ~n19346;
  assign n19621 = ~n19619 & n19620;
  assign n19622 = n19619 & ~n19620;
  assign n19623 = ~n19621 & ~n19622;
  assign n19624 = pi86  & n12295;
  assign n19625 = pi84  & n12693;
  assign n19626 = pi85  & n12290;
  assign n19627 = ~n19625 & ~n19626;
  assign n19628 = ~n19624 & n19627;
  assign n19629 = n2099 & n12298;
  assign n19630 = n19628 & ~n19629;
  assign n19631 = pi62  & ~n19630;
  assign n19632 = pi62  & ~n19631;
  assign n19633 = ~n19630 & ~n19631;
  assign n19634 = ~n19632 & ~n19633;
  assign n19635 = ~n19623 & n19634;
  assign n19636 = n19623 & ~n19634;
  assign n19637 = ~n19635 & ~n19636;
  assign n19638 = ~n19349 & ~n19352;
  assign n19639 = n19637 & ~n19638;
  assign n19640 = ~n19637 & n19638;
  assign n19641 = ~n19639 & ~n19640;
  assign n19642 = pi89  & n11193;
  assign n19643 = pi87  & n11567;
  assign n19644 = pi88  & n11188;
  assign n19645 = ~n19643 & ~n19644;
  assign n19646 = ~n19642 & n19645;
  assign n19647 = n2432 & n11196;
  assign n19648 = n19646 & ~n19647;
  assign n19649 = pi59  & ~n19648;
  assign n19650 = pi59  & ~n19649;
  assign n19651 = ~n19648 & ~n19649;
  assign n19652 = ~n19650 & ~n19651;
  assign n19653 = n19641 & ~n19652;
  assign n19654 = ~n19641 & n19652;
  assign n19655 = ~n19653 & ~n19654;
  assign n19656 = ~n19616 & n19655;
  assign n19657 = n19616 & ~n19655;
  assign n19658 = ~n19656 & ~n19657;
  assign n19659 = n19615 & ~n19658;
  assign n19660 = ~n19615 & n19658;
  assign n19661 = ~n19659 & ~n19660;
  assign n19662 = ~n19372 & ~n19378;
  assign n19663 = n19661 & ~n19662;
  assign n19664 = ~n19661 & n19662;
  assign n19665 = ~n19663 & ~n19664;
  assign n19666 = pi95  & n9096;
  assign n19667 = pi93  & n9453;
  assign n19668 = pi94  & n9091;
  assign n19669 = ~n19667 & ~n19668;
  assign n19670 = ~n19666 & n19669;
  assign n19671 = n3710 & n9099;
  assign n19672 = n19670 & ~n19671;
  assign n19673 = pi53  & ~n19672;
  assign n19674 = pi53  & ~n19673;
  assign n19675 = ~n19672 & ~n19673;
  assign n19676 = ~n19674 & ~n19675;
  assign n19677 = n19665 & ~n19676;
  assign n19678 = ~n19665 & n19676;
  assign n19679 = ~n19677 & ~n19678;
  assign n19680 = n19604 & ~n19679;
  assign n19681 = ~n19604 & n19679;
  assign n19682 = ~n19680 & ~n19681;
  assign n19683 = pi98  & n8137;
  assign n19684 = pi96  & n8471;
  assign n19685 = pi97  & n8132;
  assign n19686 = ~n19684 & ~n19685;
  assign n19687 = ~n19683 & n19686;
  assign n19688 = n4360 & n8140;
  assign n19689 = n19687 & ~n19688;
  assign n19690 = pi50  & ~n19689;
  assign n19691 = pi50  & ~n19690;
  assign n19692 = ~n19689 & ~n19690;
  assign n19693 = ~n19691 & ~n19692;
  assign n19694 = n19682 & ~n19693;
  assign n19695 = ~n19682 & n19693;
  assign n19696 = ~n19694 & ~n19695;
  assign n19697 = ~n19410 & ~n19412;
  assign n19698 = ~n19696 & ~n19697;
  assign n19699 = n19696 & n19697;
  assign n19700 = ~n19698 & ~n19699;
  assign n19701 = pi101  & n7239;
  assign n19702 = pi99  & n7556;
  assign n19703 = pi100  & n7234;
  assign n19704 = ~n19702 & ~n19703;
  assign n19705 = ~n19701 & n19704;
  assign n19706 = n5056 & n7242;
  assign n19707 = n19705 & ~n19706;
  assign n19708 = pi47  & ~n19707;
  assign n19709 = pi47  & ~n19708;
  assign n19710 = ~n19707 & ~n19708;
  assign n19711 = ~n19709 & ~n19710;
  assign n19712 = ~n19700 & n19711;
  assign n19713 = n19700 & ~n19711;
  assign n19714 = ~n19712 & ~n19713;
  assign n19715 = ~n19603 & n19714;
  assign n19716 = n19603 & ~n19714;
  assign n19717 = ~n19715 & ~n19716;
  assign n19718 = ~n19602 & n19717;
  assign n19719 = n19602 & ~n19717;
  assign n19720 = ~n19718 & ~n19719;
  assign n19721 = ~n19591 & n19720;
  assign n19722 = n19591 & ~n19720;
  assign n19723 = ~n19721 & ~n19722;
  assign n19724 = pi107  & n5636;
  assign n19725 = pi105  & n5909;
  assign n19726 = pi106  & n5631;
  assign n19727 = ~n19725 & ~n19726;
  assign n19728 = ~n19724 & n19727;
  assign n19729 = n5639 & n6614;
  assign n19730 = n19728 & ~n19729;
  assign n19731 = pi41  & ~n19730;
  assign n19732 = pi41  & ~n19731;
  assign n19733 = ~n19730 & ~n19731;
  assign n19734 = ~n19732 & ~n19733;
  assign n19735 = n19723 & ~n19734;
  assign n19736 = ~n19723 & n19734;
  assign n19737 = ~n19735 & ~n19736;
  assign n19738 = n19590 & ~n19737;
  assign n19739 = ~n19590 & n19737;
  assign n19740 = ~n19738 & ~n19739;
  assign n19741 = pi110  & n4896;
  assign n19742 = pi108  & n5148;
  assign n19743 = pi109  & n4891;
  assign n19744 = ~n19742 & ~n19743;
  assign n19745 = ~n19741 & n19744;
  assign n19746 = n4899 & n7474;
  assign n19747 = n19745 & ~n19746;
  assign n19748 = pi38  & ~n19747;
  assign n19749 = pi38  & ~n19748;
  assign n19750 = ~n19747 & ~n19748;
  assign n19751 = ~n19749 & ~n19750;
  assign n19752 = n19740 & ~n19751;
  assign n19753 = ~n19740 & n19751;
  assign n19754 = ~n19752 & ~n19753;
  assign n19755 = n19589 & ~n19754;
  assign n19756 = ~n19589 & n19754;
  assign n19757 = ~n19755 & ~n19756;
  assign n19758 = pi113  & n4182;
  assign n19759 = pi111  & n4416;
  assign n19760 = pi112  & n4177;
  assign n19761 = ~n19759 & ~n19760;
  assign n19762 = ~n19758 & n19761;
  assign n19763 = n4185 & n8387;
  assign n19764 = n19762 & ~n19763;
  assign n19765 = pi35  & ~n19764;
  assign n19766 = pi35  & ~n19765;
  assign n19767 = ~n19764 & ~n19765;
  assign n19768 = ~n19766 & ~n19767;
  assign n19769 = n19757 & ~n19768;
  assign n19770 = ~n19757 & n19768;
  assign n19771 = ~n19769 & ~n19770;
  assign n19772 = n19588 & n19771;
  assign n19773 = ~n19588 & ~n19771;
  assign n19774 = n19573 & ~n19773;
  assign n19775 = ~n19772 & n19774;
  assign n19776 = n19573 & ~n19775;
  assign n19777 = ~n19773 & ~n19775;
  assign n19778 = ~n19772 & n19777;
  assign n19779 = ~n19776 & ~n19778;
  assign n19780 = n19558 & ~n19779;
  assign n19781 = ~n19558 & n19779;
  assign n19782 = n19543 & ~n19781;
  assign n19783 = ~n19780 & n19782;
  assign n19784 = n19543 & ~n19783;
  assign n19785 = ~n19781 & ~n19783;
  assign n19786 = ~n19780 & n19785;
  assign n19787 = ~n19784 & ~n19786;
  assign n19788 = ~n19269 & ~n19515;
  assign n19789 = pi126  & n1713;
  assign n19790 = pi127  & n1577;
  assign n19791 = ~n19789 & ~n19790;
  assign n19792 = ~n1585 & n19791;
  assign n19793 = ~n13389 & n19791;
  assign n19794 = ~n19792 & ~n19793;
  assign n19795 = pi20  & ~n19794;
  assign n19796 = ~pi20  & n19794;
  assign n19797 = ~n19795 & ~n19796;
  assign n19798 = ~n19788 & ~n19797;
  assign n19799 = n19788 & n19797;
  assign n19800 = ~n19798 & ~n19799;
  assign n19801 = ~n19787 & n19800;
  assign n19802 = n19787 & ~n19800;
  assign n19803 = ~n19801 & ~n19802;
  assign n19804 = ~n19528 & n19803;
  assign n19805 = n19528 & ~n19803;
  assign n19806 = ~n19804 & ~n19805;
  assign n19807 = ~n19527 & n19806;
  assign n19808 = n19527 & ~n19806;
  assign po82  = ~n19807 & ~n19808;
  assign n19810 = ~n19804 & ~n19807;
  assign n19811 = ~n19798 & ~n19801;
  assign n19812 = pi126  & n2004;
  assign n19813 = pi124  & n2141;
  assign n19814 = pi125  & n1999;
  assign n19815 = ~n19813 & ~n19814;
  assign n19816 = ~n19812 & n19815;
  assign n19817 = n2007 & n12979;
  assign n19818 = n19816 & ~n19817;
  assign n19819 = pi23  & ~n19818;
  assign n19820 = pi23  & ~n19819;
  assign n19821 = ~n19818 & ~n19819;
  assign n19822 = ~n19820 & ~n19821;
  assign n19823 = ~n19557 & ~n19780;
  assign n19824 = ~n19822 & ~n19823;
  assign n19825 = n19822 & n19823;
  assign n19826 = ~n19824 & ~n19825;
  assign n19827 = pi123  & n2486;
  assign n19828 = pi121  & n2644;
  assign n19829 = pi122  & n2481;
  assign n19830 = ~n19828 & ~n19829;
  assign n19831 = ~n19827 & n19830;
  assign n19832 = n2489 & n11489;
  assign n19833 = n19831 & ~n19832;
  assign n19834 = pi26  & ~n19833;
  assign n19835 = pi26  & ~n19834;
  assign n19836 = ~n19833 & ~n19834;
  assign n19837 = ~n19835 & ~n19836;
  assign n19838 = ~n19572 & ~n19775;
  assign n19839 = n19837 & n19838;
  assign n19840 = ~n19837 & ~n19838;
  assign n19841 = ~n19839 & ~n19840;
  assign n19842 = pi117  & n3550;
  assign n19843 = pi115  & n3735;
  assign n19844 = pi116  & n3545;
  assign n19845 = ~n19843 & ~n19844;
  assign n19846 = ~n19842 & n19845;
  assign n19847 = n3553 & n9691;
  assign n19848 = n19846 & ~n19847;
  assign n19849 = pi32  & ~n19848;
  assign n19850 = pi32  & ~n19849;
  assign n19851 = ~n19848 & ~n19849;
  assign n19852 = ~n19850 & ~n19851;
  assign n19853 = ~n19756 & ~n19769;
  assign n19854 = n19852 & n19853;
  assign n19855 = ~n19852 & ~n19853;
  assign n19856 = ~n19854 & ~n19855;
  assign n19857 = ~n19721 & ~n19735;
  assign n19858 = pi108  & n5636;
  assign n19859 = pi106  & n5909;
  assign n19860 = pi107  & n5631;
  assign n19861 = ~n19859 & ~n19860;
  assign n19862 = ~n19858 & n19861;
  assign n19863 = n5639 & n6639;
  assign n19864 = n19862 & ~n19863;
  assign n19865 = pi41  & ~n19864;
  assign n19866 = pi41  & ~n19865;
  assign n19867 = ~n19864 & ~n19865;
  assign n19868 = ~n19866 & ~n19867;
  assign n19869 = ~n19715 & ~n19718;
  assign n19870 = pi105  & n6396;
  assign n19871 = pi103  & n6735;
  assign n19872 = pi104  & n6391;
  assign n19873 = ~n19871 & ~n19872;
  assign n19874 = ~n19870 & n19873;
  assign n19875 = n6065 & n6399;
  assign n19876 = n19874 & ~n19875;
  assign n19877 = pi44  & ~n19876;
  assign n19878 = pi44  & ~n19877;
  assign n19879 = ~n19876 & ~n19877;
  assign n19880 = ~n19878 & ~n19879;
  assign n19881 = ~n19699 & ~n19713;
  assign n19882 = pi102  & n7239;
  assign n19883 = pi100  & n7556;
  assign n19884 = pi101  & n7234;
  assign n19885 = ~n19883 & ~n19884;
  assign n19886 = ~n19882 & n19885;
  assign n19887 = n5296 & n7242;
  assign n19888 = n19886 & ~n19887;
  assign n19889 = pi47  & ~n19888;
  assign n19890 = pi47  & ~n19889;
  assign n19891 = ~n19888 & ~n19889;
  assign n19892 = ~n19890 & ~n19891;
  assign n19893 = ~n19681 & ~n19694;
  assign n19894 = pi99  & n8137;
  assign n19895 = pi97  & n8471;
  assign n19896 = pi98  & n8132;
  assign n19897 = ~n19895 & ~n19896;
  assign n19898 = ~n19894 & n19897;
  assign n19899 = n4584 & n8140;
  assign n19900 = n19898 & ~n19899;
  assign n19901 = pi50  & ~n19900;
  assign n19902 = pi50  & ~n19901;
  assign n19903 = ~n19900 & ~n19901;
  assign n19904 = ~n19902 & ~n19903;
  assign n19905 = ~n19663 & ~n19677;
  assign n19906 = pi96  & n9096;
  assign n19907 = pi94  & n9453;
  assign n19908 = pi95  & n9091;
  assign n19909 = ~n19907 & ~n19908;
  assign n19910 = ~n19906 & n19909;
  assign n19911 = n3921 & n9099;
  assign n19912 = n19910 & ~n19911;
  assign n19913 = pi53  & ~n19912;
  assign n19914 = pi53  & ~n19913;
  assign n19915 = ~n19912 & ~n19913;
  assign n19916 = ~n19914 & ~n19915;
  assign n19917 = ~n19639 & ~n19653;
  assign n19918 = pi90  & n11193;
  assign n19919 = pi88  & n11567;
  assign n19920 = pi89  & n11188;
  assign n19921 = ~n19919 & ~n19920;
  assign n19922 = ~n19918 & n19921;
  assign n19923 = n2606 & n11196;
  assign n19924 = n19922 & ~n19923;
  assign n19925 = pi59  & ~n19924;
  assign n19926 = pi59  & ~n19925;
  assign n19927 = ~n19924 & ~n19925;
  assign n19928 = ~n19926 & ~n19927;
  assign n19929 = ~n19622 & ~n19636;
  assign n19930 = pi83  & n13477;
  assign n19931 = pi84  & ~n13122;
  assign n19932 = ~n19930 & ~n19931;
  assign n19933 = ~n19619 & n19932;
  assign n19934 = n19619 & ~n19932;
  assign n19935 = ~n19933 & ~n19934;
  assign n19936 = pi87  & n12295;
  assign n19937 = pi85  & n12693;
  assign n19938 = pi86  & n12290;
  assign n19939 = ~n19937 & ~n19938;
  assign n19940 = ~n19936 & n19939;
  assign n19941 = ~n12298 & n19940;
  assign n19942 = ~n2252 & n19940;
  assign n19943 = ~n19941 & ~n19942;
  assign n19944 = pi62  & ~n19943;
  assign n19945 = ~pi62  & n19943;
  assign n19946 = ~n19944 & ~n19945;
  assign n19947 = n19935 & ~n19946;
  assign n19948 = ~n19935 & n19946;
  assign n19949 = ~n19947 & ~n19948;
  assign n19950 = ~n19929 & n19949;
  assign n19951 = n19929 & ~n19949;
  assign n19952 = ~n19950 & ~n19951;
  assign n19953 = ~n19928 & n19952;
  assign n19954 = n19928 & ~n19952;
  assign n19955 = ~n19953 & ~n19954;
  assign n19956 = ~n19917 & n19955;
  assign n19957 = n19917 & ~n19955;
  assign n19958 = ~n19956 & ~n19957;
  assign n19959 = pi93  & n10135;
  assign n19960 = pi91  & n10478;
  assign n19961 = pi92  & n10130;
  assign n19962 = ~n19960 & ~n19961;
  assign n19963 = ~n19959 & n19962;
  assign n19964 = n3144 & n10138;
  assign n19965 = n19963 & ~n19964;
  assign n19966 = pi56  & ~n19965;
  assign n19967 = pi56  & ~n19966;
  assign n19968 = ~n19965 & ~n19966;
  assign n19969 = ~n19967 & ~n19968;
  assign n19970 = n19958 & ~n19969;
  assign n19971 = n19958 & ~n19970;
  assign n19972 = ~n19969 & ~n19970;
  assign n19973 = ~n19971 & ~n19972;
  assign n19974 = ~n19656 & ~n19660;
  assign n19975 = ~n19973 & ~n19974;
  assign n19976 = n19973 & n19974;
  assign n19977 = ~n19975 & ~n19976;
  assign n19978 = n19916 & n19977;
  assign n19979 = ~n19916 & ~n19977;
  assign n19980 = ~n19978 & ~n19979;
  assign n19981 = ~n19905 & ~n19980;
  assign n19982 = n19905 & n19980;
  assign n19983 = ~n19981 & ~n19982;
  assign n19984 = ~n19904 & n19983;
  assign n19985 = n19904 & ~n19983;
  assign n19986 = ~n19984 & ~n19985;
  assign n19987 = ~n19893 & n19986;
  assign n19988 = n19893 & ~n19986;
  assign n19989 = ~n19987 & ~n19988;
  assign n19990 = ~n19892 & n19989;
  assign n19991 = n19892 & ~n19989;
  assign n19992 = ~n19990 & ~n19991;
  assign n19993 = ~n19881 & n19992;
  assign n19994 = n19881 & ~n19992;
  assign n19995 = ~n19993 & ~n19994;
  assign n19996 = ~n19880 & n19995;
  assign n19997 = n19880 & ~n19995;
  assign n19998 = ~n19996 & ~n19997;
  assign n19999 = ~n19869 & n19998;
  assign n20000 = n19869 & ~n19998;
  assign n20001 = ~n19999 & ~n20000;
  assign n20002 = ~n19868 & n20001;
  assign n20003 = n19868 & ~n20001;
  assign n20004 = ~n20002 & ~n20003;
  assign n20005 = ~n19857 & n20004;
  assign n20006 = n19857 & ~n20004;
  assign n20007 = ~n20005 & ~n20006;
  assign n20008 = pi111  & n4896;
  assign n20009 = pi109  & n5148;
  assign n20010 = pi110  & n4891;
  assign n20011 = ~n20009 & ~n20010;
  assign n20012 = ~n20008 & n20011;
  assign n20013 = n4899 & n7770;
  assign n20014 = n20012 & ~n20013;
  assign n20015 = pi38  & ~n20014;
  assign n20016 = pi38  & ~n20015;
  assign n20017 = ~n20014 & ~n20015;
  assign n20018 = ~n20016 & ~n20017;
  assign n20019 = n20007 & ~n20018;
  assign n20020 = n20007 & ~n20019;
  assign n20021 = ~n20018 & ~n20019;
  assign n20022 = ~n20020 & ~n20021;
  assign n20023 = ~n19739 & ~n19752;
  assign n20024 = n20022 & n20023;
  assign n20025 = ~n20022 & ~n20023;
  assign n20026 = ~n20024 & ~n20025;
  assign n20027 = pi114  & n4182;
  assign n20028 = pi112  & n4416;
  assign n20029 = pi113  & n4177;
  assign n20030 = ~n20028 & ~n20029;
  assign n20031 = ~n20027 & n20030;
  assign n20032 = n4185 & n8702;
  assign n20033 = n20031 & ~n20032;
  assign n20034 = pi35  & ~n20033;
  assign n20035 = pi35  & ~n20034;
  assign n20036 = ~n20033 & ~n20034;
  assign n20037 = ~n20035 & ~n20036;
  assign n20038 = n20026 & ~n20037;
  assign n20039 = ~n20026 & n20037;
  assign n20040 = n19856 & ~n20039;
  assign n20041 = ~n20038 & n20040;
  assign n20042 = n19856 & ~n20041;
  assign n20043 = ~n20039 & ~n20041;
  assign n20044 = ~n20038 & n20043;
  assign n20045 = ~n20042 & ~n20044;
  assign n20046 = pi120  & n2976;
  assign n20047 = pi118  & n3182;
  assign n20048 = pi119  & n2971;
  assign n20049 = ~n20047 & ~n20048;
  assign n20050 = ~n20046 & n20049;
  assign n20051 = n2979 & n10734;
  assign n20052 = n20050 & ~n20051;
  assign n20053 = pi29  & ~n20052;
  assign n20054 = pi29  & ~n20053;
  assign n20055 = ~n20052 & ~n20053;
  assign n20056 = ~n20054 & ~n20055;
  assign n20057 = ~n19587 & ~n19772;
  assign n20058 = ~n20056 & ~n20057;
  assign n20059 = n20056 & n20057;
  assign n20060 = ~n20058 & ~n20059;
  assign n20061 = ~n20045 & n20060;
  assign n20062 = n20045 & ~n20060;
  assign n20063 = ~n20061 & ~n20062;
  assign n20064 = n19841 & n20063;
  assign n20065 = ~n19841 & ~n20063;
  assign n20066 = ~n20064 & ~n20065;
  assign n20067 = n19826 & n20066;
  assign n20068 = ~n19826 & ~n20066;
  assign n20069 = ~n20067 & ~n20068;
  assign n20070 = ~n19542 & ~n19783;
  assign n20071 = pi127  & n1713;
  assign n20072 = n1585 & n13387;
  assign n20073 = ~n20071 & ~n20072;
  assign n20074 = pi20  & ~n20073;
  assign n20075 = pi20  & ~n20074;
  assign n20076 = ~n20073 & ~n20074;
  assign n20077 = ~n20075 & ~n20076;
  assign n20078 = ~n20070 & ~n20077;
  assign n20079 = n20070 & n20077;
  assign n20080 = ~n20078 & ~n20079;
  assign n20081 = n20069 & n20080;
  assign n20082 = ~n20069 & ~n20080;
  assign n20083 = ~n20081 & ~n20082;
  assign n20084 = ~n19811 & n20083;
  assign n20085 = n19811 & ~n20083;
  assign n20086 = ~n20084 & ~n20085;
  assign n20087 = ~n19810 & n20086;
  assign n20088 = n19810 & ~n20086;
  assign po83  = ~n20087 & ~n20088;
  assign n20090 = ~n19824 & ~n20067;
  assign n20091 = pi127  & n2004;
  assign n20092 = pi125  & n2141;
  assign n20093 = pi126  & n1999;
  assign n20094 = ~n20092 & ~n20093;
  assign n20095 = ~n20091 & n20094;
  assign n20096 = n2007 & n13365;
  assign n20097 = n20095 & ~n20096;
  assign n20098 = pi23  & ~n20097;
  assign n20099 = pi23  & ~n20098;
  assign n20100 = ~n20097 & ~n20098;
  assign n20101 = ~n20099 & ~n20100;
  assign n20102 = ~n20090 & ~n20101;
  assign n20103 = ~n20090 & ~n20102;
  assign n20104 = ~n20101 & ~n20102;
  assign n20105 = ~n20103 & ~n20104;
  assign n20106 = pi124  & n2486;
  assign n20107 = pi122  & n2644;
  assign n20108 = pi123  & n2481;
  assign n20109 = ~n20107 & ~n20108;
  assign n20110 = ~n20106 & n20109;
  assign n20111 = n2489 & n11858;
  assign n20112 = n20110 & ~n20111;
  assign n20113 = pi26  & ~n20112;
  assign n20114 = pi26  & ~n20113;
  assign n20115 = ~n20112 & ~n20113;
  assign n20116 = ~n20114 & ~n20115;
  assign n20117 = ~n19840 & ~n20064;
  assign n20118 = n20116 & n20117;
  assign n20119 = ~n20116 & ~n20117;
  assign n20120 = ~n20118 & ~n20119;
  assign n20121 = ~n20058 & ~n20061;
  assign n20122 = pi121  & n2976;
  assign n20123 = pi119  & n3182;
  assign n20124 = pi120  & n2971;
  assign n20125 = ~n20123 & ~n20124;
  assign n20126 = ~n20122 & n20125;
  assign n20127 = n2979 & n11086;
  assign n20128 = n20126 & ~n20127;
  assign n20129 = pi29  & ~n20128;
  assign n20130 = pi29  & ~n20129;
  assign n20131 = ~n20128 & ~n20129;
  assign n20132 = ~n20130 & ~n20131;
  assign n20133 = ~n20121 & ~n20132;
  assign n20134 = n20121 & n20132;
  assign n20135 = ~n20133 & ~n20134;
  assign n20136 = pi118  & n3550;
  assign n20137 = pi116  & n3735;
  assign n20138 = pi117  & n3545;
  assign n20139 = ~n20137 & ~n20138;
  assign n20140 = ~n20136 & n20139;
  assign n20141 = n3553 & n9716;
  assign n20142 = n20140 & ~n20141;
  assign n20143 = pi32  & ~n20142;
  assign n20144 = pi32  & ~n20143;
  assign n20145 = ~n20142 & ~n20143;
  assign n20146 = ~n20144 & ~n20145;
  assign n20147 = ~n19855 & ~n20041;
  assign n20148 = n20146 & n20147;
  assign n20149 = ~n20146 & ~n20147;
  assign n20150 = ~n20148 & ~n20149;
  assign n20151 = ~n20025 & ~n20038;
  assign n20152 = ~n20005 & ~n20019;
  assign n20153 = ~n19999 & ~n20002;
  assign n20154 = ~n19987 & ~n19990;
  assign n20155 = ~n19981 & ~n19984;
  assign n20156 = ~n19956 & ~n19970;
  assign n20157 = ~n19950 & ~n19953;
  assign n20158 = pi84  & n13477;
  assign n20159 = pi85  & ~n13122;
  assign n20160 = ~n20158 & ~n20159;
  assign n20161 = ~pi20  & ~n20160;
  assign n20162 = pi20  & n20160;
  assign n20163 = ~n20161 & ~n20162;
  assign n20164 = ~n19932 & n20163;
  assign n20165 = n19932 & ~n20163;
  assign n20166 = ~n20164 & ~n20165;
  assign n20167 = pi88  & n12295;
  assign n20168 = pi86  & n12693;
  assign n20169 = pi87  & n12290;
  assign n20170 = ~n20168 & ~n20169;
  assign n20171 = ~n20167 & n20170;
  assign n20172 = n2277 & n12298;
  assign n20173 = n20171 & ~n20172;
  assign n20174 = pi62  & ~n20173;
  assign n20175 = pi62  & ~n20174;
  assign n20176 = ~n20173 & ~n20174;
  assign n20177 = ~n20175 & ~n20176;
  assign n20178 = n20166 & ~n20177;
  assign n20179 = ~n20166 & n20177;
  assign n20180 = ~n20178 & ~n20179;
  assign n20181 = ~n19933 & ~n19947;
  assign n20182 = n20180 & ~n20181;
  assign n20183 = n20180 & ~n20182;
  assign n20184 = ~n20181 & ~n20182;
  assign n20185 = ~n20183 & ~n20184;
  assign n20186 = pi91  & n11193;
  assign n20187 = pi89  & n11567;
  assign n20188 = pi90  & n11188;
  assign n20189 = ~n20187 & ~n20188;
  assign n20190 = ~n20186 & n20189;
  assign n20191 = n2926 & n11196;
  assign n20192 = n20190 & ~n20191;
  assign n20193 = pi59  & ~n20192;
  assign n20194 = pi59  & ~n20193;
  assign n20195 = ~n20192 & ~n20193;
  assign n20196 = ~n20194 & ~n20195;
  assign n20197 = ~n20185 & ~n20196;
  assign n20198 = n20185 & n20196;
  assign n20199 = ~n20197 & ~n20198;
  assign n20200 = n20157 & ~n20199;
  assign n20201 = ~n20157 & n20199;
  assign n20202 = ~n20200 & ~n20201;
  assign n20203 = pi94  & n10135;
  assign n20204 = pi92  & n10478;
  assign n20205 = pi93  & n10130;
  assign n20206 = ~n20204 & ~n20205;
  assign n20207 = ~n20203 & n20206;
  assign n20208 = n3499 & n10138;
  assign n20209 = n20207 & ~n20208;
  assign n20210 = pi56  & ~n20209;
  assign n20211 = pi56  & ~n20210;
  assign n20212 = ~n20209 & ~n20210;
  assign n20213 = ~n20211 & ~n20212;
  assign n20214 = n20202 & ~n20213;
  assign n20215 = ~n20202 & n20213;
  assign n20216 = ~n20214 & ~n20215;
  assign n20217 = n20156 & ~n20216;
  assign n20218 = ~n20156 & n20216;
  assign n20219 = ~n20217 & ~n20218;
  assign n20220 = pi97  & n9096;
  assign n20221 = pi95  & n9453;
  assign n20222 = pi96  & n9091;
  assign n20223 = ~n20221 & ~n20222;
  assign n20224 = ~n20220 & n20223;
  assign n20225 = n3946 & n9099;
  assign n20226 = n20224 & ~n20225;
  assign n20227 = pi53  & ~n20226;
  assign n20228 = pi53  & ~n20227;
  assign n20229 = ~n20226 & ~n20227;
  assign n20230 = ~n20228 & ~n20229;
  assign n20231 = ~n19976 & ~n19978;
  assign n20232 = ~n20230 & n20231;
  assign n20233 = n20230 & ~n20231;
  assign n20234 = ~n20232 & ~n20233;
  assign n20235 = ~n20219 & n20234;
  assign n20236 = n20219 & ~n20234;
  assign n20237 = ~n20235 & ~n20236;
  assign n20238 = pi100  & n8137;
  assign n20239 = pi98  & n8471;
  assign n20240 = pi99  & n8132;
  assign n20241 = ~n20239 & ~n20240;
  assign n20242 = ~n20238 & n20241;
  assign n20243 = n4808 & n8140;
  assign n20244 = n20242 & ~n20243;
  assign n20245 = pi50  & ~n20244;
  assign n20246 = pi50  & ~n20245;
  assign n20247 = ~n20244 & ~n20245;
  assign n20248 = ~n20246 & ~n20247;
  assign n20249 = ~n20237 & ~n20248;
  assign n20250 = n20237 & n20248;
  assign n20251 = ~n20249 & ~n20250;
  assign n20252 = n20155 & ~n20251;
  assign n20253 = ~n20155 & n20251;
  assign n20254 = ~n20252 & ~n20253;
  assign n20255 = pi103  & n7239;
  assign n20256 = pi101  & n7556;
  assign n20257 = pi102  & n7234;
  assign n20258 = ~n20256 & ~n20257;
  assign n20259 = ~n20255 & n20258;
  assign n20260 = n5540 & n7242;
  assign n20261 = n20259 & ~n20260;
  assign n20262 = pi47  & ~n20261;
  assign n20263 = pi47  & ~n20262;
  assign n20264 = ~n20261 & ~n20262;
  assign n20265 = ~n20263 & ~n20264;
  assign n20266 = n20254 & ~n20265;
  assign n20267 = ~n20254 & n20265;
  assign n20268 = ~n20266 & ~n20267;
  assign n20269 = n20154 & ~n20268;
  assign n20270 = ~n20154 & n20268;
  assign n20271 = ~n20269 & ~n20270;
  assign n20272 = pi106  & n6396;
  assign n20273 = pi104  & n6735;
  assign n20274 = pi105  & n6391;
  assign n20275 = ~n20273 & ~n20274;
  assign n20276 = ~n20272 & n20275;
  assign n20277 = n6090 & n6399;
  assign n20278 = n20276 & ~n20277;
  assign n20279 = pi44  & ~n20278;
  assign n20280 = pi44  & ~n20279;
  assign n20281 = ~n20278 & ~n20279;
  assign n20282 = ~n20280 & ~n20281;
  assign n20283 = n20271 & ~n20282;
  assign n20284 = n20271 & ~n20283;
  assign n20285 = ~n20282 & ~n20283;
  assign n20286 = ~n20284 & ~n20285;
  assign n20287 = ~n19993 & ~n19996;
  assign n20288 = n20286 & n20287;
  assign n20289 = ~n20286 & ~n20287;
  assign n20290 = ~n20288 & ~n20289;
  assign n20291 = pi109  & n5636;
  assign n20292 = pi107  & n5909;
  assign n20293 = pi108  & n5631;
  assign n20294 = ~n20292 & ~n20293;
  assign n20295 = ~n20291 & n20294;
  assign n20296 = n5639 & n7170;
  assign n20297 = n20295 & ~n20296;
  assign n20298 = pi41  & ~n20297;
  assign n20299 = pi41  & ~n20298;
  assign n20300 = ~n20297 & ~n20298;
  assign n20301 = ~n20299 & ~n20300;
  assign n20302 = n20290 & ~n20301;
  assign n20303 = ~n20290 & n20301;
  assign n20304 = ~n20302 & ~n20303;
  assign n20305 = n20153 & ~n20304;
  assign n20306 = ~n20153 & n20304;
  assign n20307 = ~n20305 & ~n20306;
  assign n20308 = pi112  & n4896;
  assign n20309 = pi110  & n5148;
  assign n20310 = pi111  & n4891;
  assign n20311 = ~n20309 & ~n20310;
  assign n20312 = ~n20308 & n20311;
  assign n20313 = n4899 & n7795;
  assign n20314 = n20312 & ~n20313;
  assign n20315 = pi38  & ~n20314;
  assign n20316 = pi38  & ~n20315;
  assign n20317 = ~n20314 & ~n20315;
  assign n20318 = ~n20316 & ~n20317;
  assign n20319 = n20307 & ~n20318;
  assign n20320 = ~n20307 & n20318;
  assign n20321 = ~n20319 & ~n20320;
  assign n20322 = n20152 & ~n20321;
  assign n20323 = ~n20152 & n20321;
  assign n20324 = ~n20322 & ~n20323;
  assign n20325 = pi115  & n4182;
  assign n20326 = pi113  & n4416;
  assign n20327 = pi114  & n4177;
  assign n20328 = ~n20326 & ~n20327;
  assign n20329 = ~n20325 & n20328;
  assign n20330 = n4185 & n8727;
  assign n20331 = n20329 & ~n20330;
  assign n20332 = pi35  & ~n20331;
  assign n20333 = pi35  & ~n20332;
  assign n20334 = ~n20331 & ~n20332;
  assign n20335 = ~n20333 & ~n20334;
  assign n20336 = n20324 & ~n20335;
  assign n20337 = ~n20324 & n20335;
  assign n20338 = ~n20151 & ~n20337;
  assign n20339 = ~n20336 & n20338;
  assign n20340 = ~n20151 & ~n20339;
  assign n20341 = ~n20336 & ~n20339;
  assign n20342 = ~n20337 & n20341;
  assign n20343 = ~n20340 & ~n20342;
  assign n20344 = n20150 & ~n20343;
  assign n20345 = ~n20150 & n20343;
  assign n20346 = n20135 & ~n20345;
  assign n20347 = ~n20344 & n20346;
  assign n20348 = n20135 & ~n20347;
  assign n20349 = ~n20345 & ~n20347;
  assign n20350 = ~n20344 & n20349;
  assign n20351 = ~n20348 & ~n20350;
  assign n20352 = n20120 & ~n20351;
  assign n20353 = ~n20120 & n20351;
  assign n20354 = ~n20105 & ~n20353;
  assign n20355 = ~n20352 & n20354;
  assign n20356 = ~n20105 & ~n20355;
  assign n20357 = ~n20353 & ~n20355;
  assign n20358 = ~n20352 & n20357;
  assign n20359 = ~n20356 & ~n20358;
  assign n20360 = ~n20078 & ~n20081;
  assign n20361 = n20359 & n20360;
  assign n20362 = ~n20359 & ~n20360;
  assign n20363 = ~n20361 & ~n20362;
  assign n20364 = ~n20084 & ~n20087;
  assign n20365 = n20363 & ~n20364;
  assign n20366 = ~n20363 & n20364;
  assign po84  = ~n20365 & ~n20366;
  assign n20368 = ~n20119 & ~n20352;
  assign n20369 = pi126  & n2141;
  assign n20370 = pi127  & n1999;
  assign n20371 = ~n20369 & ~n20370;
  assign n20372 = ~n2007 & n20371;
  assign n20373 = ~n13389 & n20371;
  assign n20374 = ~n20372 & ~n20373;
  assign n20375 = pi23  & ~n20374;
  assign n20376 = ~pi23  & n20374;
  assign n20377 = ~n20375 & ~n20376;
  assign n20378 = ~n20368 & ~n20377;
  assign n20379 = n20368 & n20377;
  assign n20380 = ~n20378 & ~n20379;
  assign n20381 = pi125  & n2486;
  assign n20382 = pi123  & n2644;
  assign n20383 = pi124  & n2481;
  assign n20384 = ~n20382 & ~n20383;
  assign n20385 = ~n20381 & n20384;
  assign n20386 = n2489 & n12591;
  assign n20387 = n20385 & ~n20386;
  assign n20388 = pi26  & ~n20387;
  assign n20389 = pi26  & ~n20388;
  assign n20390 = ~n20387 & ~n20388;
  assign n20391 = ~n20389 & ~n20390;
  assign n20392 = ~n20133 & ~n20347;
  assign n20393 = n20391 & n20392;
  assign n20394 = ~n20391 & ~n20392;
  assign n20395 = ~n20393 & ~n20394;
  assign n20396 = ~n20149 & ~n20344;
  assign n20397 = pi122  & n2976;
  assign n20398 = pi120  & n3182;
  assign n20399 = pi121  & n2971;
  assign n20400 = ~n20398 & ~n20399;
  assign n20401 = ~n20397 & n20400;
  assign n20402 = ~n2979 & n20401;
  assign n20403 = ~n11463 & n20401;
  assign n20404 = ~n20402 & ~n20403;
  assign n20405 = pi29  & ~n20404;
  assign n20406 = ~pi29  & n20404;
  assign n20407 = ~n20405 & ~n20406;
  assign n20408 = ~n20396 & ~n20407;
  assign n20409 = n20396 & n20407;
  assign n20410 = ~n20408 & ~n20409;
  assign n20411 = pi119  & n3550;
  assign n20412 = pi117  & n3735;
  assign n20413 = pi118  & n3545;
  assign n20414 = ~n20412 & ~n20413;
  assign n20415 = ~n20411 & n20414;
  assign n20416 = n3553 & n10048;
  assign n20417 = n20415 & ~n20416;
  assign n20418 = pi32  & ~n20417;
  assign n20419 = pi32  & ~n20418;
  assign n20420 = ~n20417 & ~n20418;
  assign n20421 = ~n20419 & ~n20420;
  assign n20422 = ~n20341 & ~n20421;
  assign n20423 = n20341 & n20421;
  assign n20424 = ~n20422 & ~n20423;
  assign n20425 = ~n20319 & ~n20323;
  assign n20426 = ~n20302 & ~n20306;
  assign n20427 = ~n20283 & ~n20289;
  assign n20428 = ~n20266 & ~n20270;
  assign n20429 = pi104  & n7239;
  assign n20430 = pi102  & n7556;
  assign n20431 = pi103  & n7234;
  assign n20432 = ~n20430 & ~n20431;
  assign n20433 = ~n20429 & n20432;
  assign n20434 = n5565 & n7242;
  assign n20435 = n20433 & ~n20434;
  assign n20436 = pi47  & ~n20435;
  assign n20437 = pi47  & ~n20436;
  assign n20438 = ~n20435 & ~n20436;
  assign n20439 = ~n20437 & ~n20438;
  assign n20440 = ~n20249 & ~n20253;
  assign n20441 = ~n20214 & ~n20218;
  assign n20442 = ~n20197 & ~n20201;
  assign n20443 = pi92  & n11193;
  assign n20444 = pi90  & n11567;
  assign n20445 = pi91  & n11188;
  assign n20446 = ~n20444 & ~n20445;
  assign n20447 = ~n20443 & n20446;
  assign n20448 = n3119 & n11196;
  assign n20449 = n20447 & ~n20448;
  assign n20450 = pi59  & ~n20449;
  assign n20451 = pi59  & ~n20450;
  assign n20452 = ~n20449 & ~n20450;
  assign n20453 = ~n20451 & ~n20452;
  assign n20454 = ~n20178 & ~n20182;
  assign n20455 = pi85  & n13477;
  assign n20456 = pi86  & ~n13122;
  assign n20457 = ~n20455 & ~n20456;
  assign n20458 = ~n20161 & ~n20164;
  assign n20459 = ~n20457 & n20458;
  assign n20460 = n20457 & ~n20458;
  assign n20461 = ~n20459 & ~n20460;
  assign n20462 = pi89  & n12295;
  assign n20463 = pi87  & n12693;
  assign n20464 = pi88  & n12290;
  assign n20465 = ~n20463 & ~n20464;
  assign n20466 = ~n20462 & n20465;
  assign n20467 = ~n12298 & n20466;
  assign n20468 = ~n2432 & n20466;
  assign n20469 = ~n20467 & ~n20468;
  assign n20470 = pi62  & ~n20469;
  assign n20471 = ~pi62  & n20469;
  assign n20472 = ~n20470 & ~n20471;
  assign n20473 = n20461 & ~n20472;
  assign n20474 = ~n20461 & n20472;
  assign n20475 = ~n20473 & ~n20474;
  assign n20476 = ~n20454 & n20475;
  assign n20477 = n20454 & ~n20475;
  assign n20478 = ~n20476 & ~n20477;
  assign n20479 = ~n20453 & n20478;
  assign n20480 = n20453 & ~n20478;
  assign n20481 = ~n20479 & ~n20480;
  assign n20482 = ~n20442 & n20481;
  assign n20483 = n20442 & ~n20481;
  assign n20484 = ~n20482 & ~n20483;
  assign n20485 = pi95  & n10135;
  assign n20486 = pi93  & n10478;
  assign n20487 = pi94  & n10130;
  assign n20488 = ~n20486 & ~n20487;
  assign n20489 = ~n20485 & n20488;
  assign n20490 = n3710 & n10138;
  assign n20491 = n20489 & ~n20490;
  assign n20492 = pi56  & ~n20491;
  assign n20493 = pi56  & ~n20492;
  assign n20494 = ~n20491 & ~n20492;
  assign n20495 = ~n20493 & ~n20494;
  assign n20496 = n20484 & ~n20495;
  assign n20497 = ~n20484 & n20495;
  assign n20498 = ~n20496 & ~n20497;
  assign n20499 = n20441 & ~n20498;
  assign n20500 = ~n20441 & n20498;
  assign n20501 = ~n20499 & ~n20500;
  assign n20502 = pi98  & n9096;
  assign n20503 = pi96  & n9453;
  assign n20504 = pi97  & n9091;
  assign n20505 = ~n20503 & ~n20504;
  assign n20506 = ~n20502 & n20505;
  assign n20507 = n4360 & n9099;
  assign n20508 = n20506 & ~n20507;
  assign n20509 = pi53  & ~n20508;
  assign n20510 = pi53  & ~n20509;
  assign n20511 = ~n20508 & ~n20509;
  assign n20512 = ~n20510 & ~n20511;
  assign n20513 = n20501 & ~n20512;
  assign n20514 = ~n20501 & n20512;
  assign n20515 = ~n20513 & ~n20514;
  assign n20516 = ~n20233 & ~n20235;
  assign n20517 = ~n20515 & ~n20516;
  assign n20518 = n20515 & n20516;
  assign n20519 = ~n20517 & ~n20518;
  assign n20520 = pi101  & n8137;
  assign n20521 = pi99  & n8471;
  assign n20522 = pi100  & n8132;
  assign n20523 = ~n20521 & ~n20522;
  assign n20524 = ~n20520 & n20523;
  assign n20525 = n5056 & n8140;
  assign n20526 = n20524 & ~n20525;
  assign n20527 = pi50  & ~n20526;
  assign n20528 = pi50  & ~n20527;
  assign n20529 = ~n20526 & ~n20527;
  assign n20530 = ~n20528 & ~n20529;
  assign n20531 = ~n20519 & n20530;
  assign n20532 = n20519 & ~n20530;
  assign n20533 = ~n20531 & ~n20532;
  assign n20534 = ~n20440 & n20533;
  assign n20535 = n20440 & ~n20533;
  assign n20536 = ~n20534 & ~n20535;
  assign n20537 = ~n20439 & n20536;
  assign n20538 = n20439 & ~n20536;
  assign n20539 = ~n20537 & ~n20538;
  assign n20540 = ~n20428 & n20539;
  assign n20541 = n20428 & ~n20539;
  assign n20542 = ~n20540 & ~n20541;
  assign n20543 = pi107  & n6396;
  assign n20544 = pi105  & n6735;
  assign n20545 = pi106  & n6391;
  assign n20546 = ~n20544 & ~n20545;
  assign n20547 = ~n20543 & n20546;
  assign n20548 = n6399 & n6614;
  assign n20549 = n20547 & ~n20548;
  assign n20550 = pi44  & ~n20549;
  assign n20551 = pi44  & ~n20550;
  assign n20552 = ~n20549 & ~n20550;
  assign n20553 = ~n20551 & ~n20552;
  assign n20554 = n20542 & ~n20553;
  assign n20555 = ~n20542 & n20553;
  assign n20556 = ~n20554 & ~n20555;
  assign n20557 = n20427 & ~n20556;
  assign n20558 = ~n20427 & n20556;
  assign n20559 = ~n20557 & ~n20558;
  assign n20560 = pi110  & n5636;
  assign n20561 = pi108  & n5909;
  assign n20562 = pi109  & n5631;
  assign n20563 = ~n20561 & ~n20562;
  assign n20564 = ~n20560 & n20563;
  assign n20565 = n5639 & n7474;
  assign n20566 = n20564 & ~n20565;
  assign n20567 = pi41  & ~n20566;
  assign n20568 = pi41  & ~n20567;
  assign n20569 = ~n20566 & ~n20567;
  assign n20570 = ~n20568 & ~n20569;
  assign n20571 = n20559 & ~n20570;
  assign n20572 = ~n20559 & n20570;
  assign n20573 = ~n20571 & ~n20572;
  assign n20574 = n20426 & ~n20573;
  assign n20575 = ~n20426 & n20573;
  assign n20576 = ~n20574 & ~n20575;
  assign n20577 = pi113  & n4896;
  assign n20578 = pi111  & n5148;
  assign n20579 = pi112  & n4891;
  assign n20580 = ~n20578 & ~n20579;
  assign n20581 = ~n20577 & n20580;
  assign n20582 = n4899 & n8387;
  assign n20583 = n20581 & ~n20582;
  assign n20584 = pi38  & ~n20583;
  assign n20585 = pi38  & ~n20584;
  assign n20586 = ~n20583 & ~n20584;
  assign n20587 = ~n20585 & ~n20586;
  assign n20588 = n20576 & ~n20587;
  assign n20589 = ~n20576 & n20587;
  assign n20590 = ~n20588 & ~n20589;
  assign n20591 = n20425 & ~n20590;
  assign n20592 = ~n20425 & n20590;
  assign n20593 = ~n20591 & ~n20592;
  assign n20594 = pi116  & n4182;
  assign n20595 = pi114  & n4416;
  assign n20596 = pi115  & n4177;
  assign n20597 = ~n20595 & ~n20596;
  assign n20598 = ~n20594 & n20597;
  assign n20599 = n4185 & n9042;
  assign n20600 = n20598 & ~n20599;
  assign n20601 = pi35  & ~n20600;
  assign n20602 = pi35  & ~n20601;
  assign n20603 = ~n20600 & ~n20601;
  assign n20604 = ~n20602 & ~n20603;
  assign n20605 = n20593 & ~n20604;
  assign n20606 = ~n20593 & n20604;
  assign n20607 = ~n20605 & ~n20606;
  assign n20608 = n20424 & n20607;
  assign n20609 = ~n20424 & ~n20607;
  assign n20610 = n20410 & ~n20609;
  assign n20611 = ~n20608 & n20610;
  assign n20612 = n20410 & ~n20611;
  assign n20613 = ~n20609 & ~n20611;
  assign n20614 = ~n20608 & n20613;
  assign n20615 = ~n20612 & ~n20614;
  assign n20616 = n20395 & ~n20615;
  assign n20617 = ~n20395 & n20615;
  assign n20618 = n20380 & ~n20617;
  assign n20619 = ~n20616 & n20618;
  assign n20620 = n20380 & ~n20619;
  assign n20621 = ~n20617 & ~n20619;
  assign n20622 = ~n20616 & n20621;
  assign n20623 = ~n20620 & ~n20622;
  assign n20624 = ~n20102 & ~n20355;
  assign n20625 = n20623 & n20624;
  assign n20626 = ~n20623 & ~n20624;
  assign n20627 = ~n20625 & ~n20626;
  assign n20628 = ~n20362 & ~n20365;
  assign n20629 = n20627 & ~n20628;
  assign n20630 = ~n20627 & n20628;
  assign po85  = ~n20629 & ~n20630;
  assign n20632 = ~n20626 & ~n20629;
  assign n20633 = ~n20378 & ~n20619;
  assign n20634 = ~n20394 & ~n20616;
  assign n20635 = pi127  & n2141;
  assign n20636 = n2007 & n13387;
  assign n20637 = ~n20635 & ~n20636;
  assign n20638 = pi23  & ~n20637;
  assign n20639 = pi23  & ~n20638;
  assign n20640 = ~n20637 & ~n20638;
  assign n20641 = ~n20639 & ~n20640;
  assign n20642 = ~n20634 & ~n20641;
  assign n20643 = n20634 & n20641;
  assign n20644 = ~n20642 & ~n20643;
  assign n20645 = pi126  & n2486;
  assign n20646 = pi124  & n2644;
  assign n20647 = pi125  & n2481;
  assign n20648 = ~n20646 & ~n20647;
  assign n20649 = ~n20645 & n20648;
  assign n20650 = n2489 & n12979;
  assign n20651 = n20649 & ~n20650;
  assign n20652 = pi26  & ~n20651;
  assign n20653 = pi26  & ~n20652;
  assign n20654 = ~n20651 & ~n20652;
  assign n20655 = ~n20653 & ~n20654;
  assign n20656 = ~n20408 & ~n20611;
  assign n20657 = n20655 & n20656;
  assign n20658 = ~n20655 & ~n20656;
  assign n20659 = ~n20657 & ~n20658;
  assign n20660 = pi123  & n2976;
  assign n20661 = pi121  & n3182;
  assign n20662 = pi122  & n2971;
  assign n20663 = ~n20661 & ~n20662;
  assign n20664 = ~n20660 & n20663;
  assign n20665 = n2979 & n11489;
  assign n20666 = n20664 & ~n20665;
  assign n20667 = pi29  & ~n20666;
  assign n20668 = pi29  & ~n20667;
  assign n20669 = ~n20666 & ~n20667;
  assign n20670 = ~n20668 & ~n20669;
  assign n20671 = ~n20422 & ~n20608;
  assign n20672 = ~n20670 & ~n20671;
  assign n20673 = n20670 & n20671;
  assign n20674 = ~n20672 & ~n20673;
  assign n20675 = pi120  & n3550;
  assign n20676 = pi118  & n3735;
  assign n20677 = pi119  & n3545;
  assign n20678 = ~n20676 & ~n20677;
  assign n20679 = ~n20675 & n20678;
  assign n20680 = n3553 & n10734;
  assign n20681 = n20679 & ~n20680;
  assign n20682 = pi32  & ~n20681;
  assign n20683 = pi32  & ~n20682;
  assign n20684 = ~n20681 & ~n20682;
  assign n20685 = ~n20683 & ~n20684;
  assign n20686 = ~n20592 & ~n20605;
  assign n20687 = n20685 & n20686;
  assign n20688 = ~n20685 & ~n20686;
  assign n20689 = ~n20687 & ~n20688;
  assign n20690 = pi117  & n4182;
  assign n20691 = pi115  & n4416;
  assign n20692 = pi116  & n4177;
  assign n20693 = ~n20691 & ~n20692;
  assign n20694 = ~n20690 & n20693;
  assign n20695 = n4185 & n9691;
  assign n20696 = n20694 & ~n20695;
  assign n20697 = pi35  & ~n20696;
  assign n20698 = pi35  & ~n20697;
  assign n20699 = ~n20696 & ~n20697;
  assign n20700 = ~n20698 & ~n20699;
  assign n20701 = ~n20575 & ~n20588;
  assign n20702 = ~n20540 & ~n20554;
  assign n20703 = pi108  & n6396;
  assign n20704 = pi106  & n6735;
  assign n20705 = pi107  & n6391;
  assign n20706 = ~n20704 & ~n20705;
  assign n20707 = ~n20703 & n20706;
  assign n20708 = n6399 & n6639;
  assign n20709 = n20707 & ~n20708;
  assign n20710 = pi44  & ~n20709;
  assign n20711 = pi44  & ~n20710;
  assign n20712 = ~n20709 & ~n20710;
  assign n20713 = ~n20711 & ~n20712;
  assign n20714 = ~n20534 & ~n20537;
  assign n20715 = pi105  & n7239;
  assign n20716 = pi103  & n7556;
  assign n20717 = pi104  & n7234;
  assign n20718 = ~n20716 & ~n20717;
  assign n20719 = ~n20715 & n20718;
  assign n20720 = n6065 & n7242;
  assign n20721 = n20719 & ~n20720;
  assign n20722 = pi47  & ~n20721;
  assign n20723 = pi47  & ~n20722;
  assign n20724 = ~n20721 & ~n20722;
  assign n20725 = ~n20723 & ~n20724;
  assign n20726 = ~n20500 & ~n20513;
  assign n20727 = pi99  & n9096;
  assign n20728 = pi97  & n9453;
  assign n20729 = pi98  & n9091;
  assign n20730 = ~n20728 & ~n20729;
  assign n20731 = ~n20727 & n20730;
  assign n20732 = n4584 & n9099;
  assign n20733 = n20731 & ~n20732;
  assign n20734 = pi53  & ~n20733;
  assign n20735 = pi53  & ~n20734;
  assign n20736 = ~n20733 & ~n20734;
  assign n20737 = ~n20735 & ~n20736;
  assign n20738 = ~n20482 & ~n20496;
  assign n20739 = ~n20460 & ~n20473;
  assign n20740 = pi86  & n13477;
  assign n20741 = pi87  & ~n13122;
  assign n20742 = ~n20740 & ~n20741;
  assign n20743 = ~n20457 & n20742;
  assign n20744 = n20457 & ~n20742;
  assign n20745 = ~n20743 & ~n20744;
  assign n20746 = pi90  & n12295;
  assign n20747 = pi88  & n12693;
  assign n20748 = pi89  & n12290;
  assign n20749 = ~n20747 & ~n20748;
  assign n20750 = ~n20746 & n20749;
  assign n20751 = ~n12298 & n20750;
  assign n20752 = ~n2606 & n20750;
  assign n20753 = ~n20751 & ~n20752;
  assign n20754 = pi62  & ~n20753;
  assign n20755 = ~pi62  & n20753;
  assign n20756 = ~n20754 & ~n20755;
  assign n20757 = n20745 & ~n20756;
  assign n20758 = ~n20745 & n20756;
  assign n20759 = ~n20757 & ~n20758;
  assign n20760 = ~n20739 & n20759;
  assign n20761 = n20739 & ~n20759;
  assign n20762 = ~n20760 & ~n20761;
  assign n20763 = pi93  & n11193;
  assign n20764 = pi91  & n11567;
  assign n20765 = pi92  & n11188;
  assign n20766 = ~n20764 & ~n20765;
  assign n20767 = ~n20763 & n20766;
  assign n20768 = n3144 & n11196;
  assign n20769 = n20767 & ~n20768;
  assign n20770 = pi59  & ~n20769;
  assign n20771 = pi59  & ~n20770;
  assign n20772 = ~n20769 & ~n20770;
  assign n20773 = ~n20771 & ~n20772;
  assign n20774 = n20762 & ~n20773;
  assign n20775 = n20762 & ~n20774;
  assign n20776 = ~n20773 & ~n20774;
  assign n20777 = ~n20775 & ~n20776;
  assign n20778 = ~n20476 & ~n20479;
  assign n20779 = n20777 & n20778;
  assign n20780 = ~n20777 & ~n20778;
  assign n20781 = ~n20779 & ~n20780;
  assign n20782 = pi96  & n10135;
  assign n20783 = pi94  & n10478;
  assign n20784 = pi95  & n10130;
  assign n20785 = ~n20783 & ~n20784;
  assign n20786 = ~n20782 & n20785;
  assign n20787 = n3921 & n10138;
  assign n20788 = n20786 & ~n20787;
  assign n20789 = pi56  & ~n20788;
  assign n20790 = pi56  & ~n20789;
  assign n20791 = ~n20788 & ~n20789;
  assign n20792 = ~n20790 & ~n20791;
  assign n20793 = ~n20781 & n20792;
  assign n20794 = n20781 & ~n20792;
  assign n20795 = ~n20793 & ~n20794;
  assign n20796 = ~n20738 & n20795;
  assign n20797 = n20738 & ~n20795;
  assign n20798 = ~n20796 & ~n20797;
  assign n20799 = ~n20737 & n20798;
  assign n20800 = n20737 & ~n20798;
  assign n20801 = ~n20799 & ~n20800;
  assign n20802 = ~n20726 & n20801;
  assign n20803 = n20726 & ~n20801;
  assign n20804 = ~n20802 & ~n20803;
  assign n20805 = pi102  & n8137;
  assign n20806 = pi100  & n8471;
  assign n20807 = pi101  & n8132;
  assign n20808 = ~n20806 & ~n20807;
  assign n20809 = ~n20805 & n20808;
  assign n20810 = n5296 & n8140;
  assign n20811 = n20809 & ~n20810;
  assign n20812 = pi50  & ~n20811;
  assign n20813 = pi50  & ~n20812;
  assign n20814 = ~n20811 & ~n20812;
  assign n20815 = ~n20813 & ~n20814;
  assign n20816 = n20804 & ~n20815;
  assign n20817 = n20804 & ~n20816;
  assign n20818 = ~n20815 & ~n20816;
  assign n20819 = ~n20817 & ~n20818;
  assign n20820 = ~n20518 & ~n20532;
  assign n20821 = ~n20819 & ~n20820;
  assign n20822 = n20819 & n20820;
  assign n20823 = ~n20821 & ~n20822;
  assign n20824 = n20725 & n20823;
  assign n20825 = ~n20725 & ~n20823;
  assign n20826 = ~n20824 & ~n20825;
  assign n20827 = ~n20714 & ~n20826;
  assign n20828 = n20714 & n20826;
  assign n20829 = ~n20827 & ~n20828;
  assign n20830 = ~n20713 & n20829;
  assign n20831 = n20713 & ~n20829;
  assign n20832 = ~n20830 & ~n20831;
  assign n20833 = ~n20702 & n20832;
  assign n20834 = n20702 & ~n20832;
  assign n20835 = ~n20833 & ~n20834;
  assign n20836 = pi111  & n5636;
  assign n20837 = pi109  & n5909;
  assign n20838 = pi110  & n5631;
  assign n20839 = ~n20837 & ~n20838;
  assign n20840 = ~n20836 & n20839;
  assign n20841 = n5639 & n7770;
  assign n20842 = n20840 & ~n20841;
  assign n20843 = pi41  & ~n20842;
  assign n20844 = pi41  & ~n20843;
  assign n20845 = ~n20842 & ~n20843;
  assign n20846 = ~n20844 & ~n20845;
  assign n20847 = n20835 & ~n20846;
  assign n20848 = n20835 & ~n20847;
  assign n20849 = ~n20846 & ~n20847;
  assign n20850 = ~n20848 & ~n20849;
  assign n20851 = ~n20558 & ~n20571;
  assign n20852 = n20850 & n20851;
  assign n20853 = ~n20850 & ~n20851;
  assign n20854 = ~n20852 & ~n20853;
  assign n20855 = pi114  & n4896;
  assign n20856 = pi112  & n5148;
  assign n20857 = pi113  & n4891;
  assign n20858 = ~n20856 & ~n20857;
  assign n20859 = ~n20855 & n20858;
  assign n20860 = n4899 & n8702;
  assign n20861 = n20859 & ~n20860;
  assign n20862 = pi38  & ~n20861;
  assign n20863 = pi38  & ~n20862;
  assign n20864 = ~n20861 & ~n20862;
  assign n20865 = ~n20863 & ~n20864;
  assign n20866 = ~n20854 & n20865;
  assign n20867 = n20854 & ~n20865;
  assign n20868 = ~n20866 & ~n20867;
  assign n20869 = ~n20701 & n20868;
  assign n20870 = n20701 & ~n20868;
  assign n20871 = ~n20869 & ~n20870;
  assign n20872 = ~n20700 & n20871;
  assign n20873 = n20700 & ~n20871;
  assign n20874 = ~n20872 & ~n20873;
  assign n20875 = n20689 & n20874;
  assign n20876 = ~n20689 & ~n20874;
  assign n20877 = ~n20875 & ~n20876;
  assign n20878 = n20674 & n20877;
  assign n20879 = ~n20674 & ~n20877;
  assign n20880 = ~n20878 & ~n20879;
  assign n20881 = n20659 & n20880;
  assign n20882 = ~n20659 & ~n20880;
  assign n20883 = ~n20881 & ~n20882;
  assign n20884 = n20644 & n20883;
  assign n20885 = ~n20644 & ~n20883;
  assign n20886 = ~n20884 & ~n20885;
  assign n20887 = ~n20633 & n20886;
  assign n20888 = n20633 & ~n20886;
  assign n20889 = ~n20887 & ~n20888;
  assign n20890 = ~n20632 & n20889;
  assign n20891 = n20632 & ~n20889;
  assign po86  = ~n20890 & ~n20891;
  assign n20893 = ~n20887 & ~n20890;
  assign n20894 = ~n20642 & ~n20884;
  assign n20895 = ~n20658 & ~n20881;
  assign n20896 = pi127  & n2486;
  assign n20897 = pi125  & n2644;
  assign n20898 = pi126  & n2481;
  assign n20899 = ~n20897 & ~n20898;
  assign n20900 = ~n20896 & n20899;
  assign n20901 = n2489 & n13365;
  assign n20902 = n20900 & ~n20901;
  assign n20903 = pi26  & ~n20902;
  assign n20904 = pi26  & ~n20903;
  assign n20905 = ~n20902 & ~n20903;
  assign n20906 = ~n20904 & ~n20905;
  assign n20907 = ~n20895 & ~n20906;
  assign n20908 = ~n20895 & ~n20907;
  assign n20909 = ~n20906 & ~n20907;
  assign n20910 = ~n20908 & ~n20909;
  assign n20911 = ~n20672 & ~n20878;
  assign n20912 = pi124  & n2976;
  assign n20913 = pi122  & n3182;
  assign n20914 = pi123  & n2971;
  assign n20915 = ~n20913 & ~n20914;
  assign n20916 = ~n20912 & n20915;
  assign n20917 = n2979 & n11858;
  assign n20918 = n20916 & ~n20917;
  assign n20919 = pi29  & ~n20918;
  assign n20920 = pi29  & ~n20919;
  assign n20921 = ~n20918 & ~n20919;
  assign n20922 = ~n20920 & ~n20921;
  assign n20923 = ~n20911 & n20922;
  assign n20924 = n20911 & ~n20922;
  assign n20925 = ~n20923 & ~n20924;
  assign n20926 = pi121  & n3550;
  assign n20927 = pi119  & n3735;
  assign n20928 = pi120  & n3545;
  assign n20929 = ~n20927 & ~n20928;
  assign n20930 = ~n20926 & n20929;
  assign n20931 = n3553 & n11086;
  assign n20932 = n20930 & ~n20931;
  assign n20933 = pi32  & ~n20932;
  assign n20934 = pi32  & ~n20933;
  assign n20935 = ~n20932 & ~n20933;
  assign n20936 = ~n20934 & ~n20935;
  assign n20937 = ~n20688 & ~n20875;
  assign n20938 = n20936 & n20937;
  assign n20939 = ~n20936 & ~n20937;
  assign n20940 = ~n20938 & ~n20939;
  assign n20941 = ~n20869 & ~n20872;
  assign n20942 = ~n20853 & ~n20867;
  assign n20943 = ~n20833 & ~n20847;
  assign n20944 = ~n20827 & ~n20830;
  assign n20945 = ~n20822 & ~n20824;
  assign n20946 = ~n20802 & ~n20816;
  assign n20947 = ~n20796 & ~n20799;
  assign n20948 = ~n20760 & ~n20774;
  assign n20949 = ~n20743 & ~n20757;
  assign n20950 = pi87  & n13477;
  assign n20951 = pi88  & ~n13122;
  assign n20952 = ~n20950 & ~n20951;
  assign n20953 = ~pi23  & ~n20952;
  assign n20954 = pi23  & n20952;
  assign n20955 = ~n20953 & ~n20954;
  assign n20956 = ~n20742 & n20955;
  assign n20957 = n20742 & ~n20955;
  assign n20958 = ~n20956 & ~n20957;
  assign n20959 = pi91  & n12295;
  assign n20960 = pi89  & n12693;
  assign n20961 = pi90  & n12290;
  assign n20962 = ~n20960 & ~n20961;
  assign n20963 = ~n20959 & n20962;
  assign n20964 = n2926 & n12298;
  assign n20965 = n20963 & ~n20964;
  assign n20966 = pi62  & ~n20965;
  assign n20967 = pi62  & ~n20966;
  assign n20968 = ~n20965 & ~n20966;
  assign n20969 = ~n20967 & ~n20968;
  assign n20970 = n20958 & ~n20969;
  assign n20971 = ~n20958 & n20969;
  assign n20972 = ~n20970 & ~n20971;
  assign n20973 = ~n20949 & ~n20972;
  assign n20974 = n20949 & n20972;
  assign n20975 = ~n20973 & ~n20974;
  assign n20976 = pi94  & n11193;
  assign n20977 = pi92  & n11567;
  assign n20978 = pi93  & n11188;
  assign n20979 = ~n20977 & ~n20978;
  assign n20980 = ~n20976 & n20979;
  assign n20981 = n3499 & n11196;
  assign n20982 = n20980 & ~n20981;
  assign n20983 = pi59  & ~n20982;
  assign n20984 = pi59  & ~n20983;
  assign n20985 = ~n20982 & ~n20983;
  assign n20986 = ~n20984 & ~n20985;
  assign n20987 = ~n20975 & ~n20986;
  assign n20988 = n20975 & n20986;
  assign n20989 = ~n20987 & ~n20988;
  assign n20990 = n20948 & ~n20989;
  assign n20991 = ~n20948 & n20989;
  assign n20992 = ~n20990 & ~n20991;
  assign n20993 = pi97  & n10135;
  assign n20994 = pi95  & n10478;
  assign n20995 = pi96  & n10130;
  assign n20996 = ~n20994 & ~n20995;
  assign n20997 = ~n20993 & n20996;
  assign n20998 = n3946 & n10138;
  assign n20999 = n20997 & ~n20998;
  assign n21000 = pi56  & ~n20999;
  assign n21001 = pi56  & ~n21000;
  assign n21002 = ~n20999 & ~n21000;
  assign n21003 = ~n21001 & ~n21002;
  assign n21004 = ~n20780 & ~n20794;
  assign n21005 = ~n21003 & ~n21004;
  assign n21006 = n21003 & n21004;
  assign n21007 = ~n21005 & ~n21006;
  assign n21008 = n20992 & n21007;
  assign n21009 = ~n20992 & ~n21007;
  assign n21010 = ~n21008 & ~n21009;
  assign n21011 = pi100  & n9096;
  assign n21012 = pi98  & n9453;
  assign n21013 = pi99  & n9091;
  assign n21014 = ~n21012 & ~n21013;
  assign n21015 = ~n21011 & n21014;
  assign n21016 = n4808 & n9099;
  assign n21017 = n21015 & ~n21016;
  assign n21018 = pi53  & ~n21017;
  assign n21019 = pi53  & ~n21018;
  assign n21020 = ~n21017 & ~n21018;
  assign n21021 = ~n21019 & ~n21020;
  assign n21022 = n21010 & ~n21021;
  assign n21023 = ~n21010 & n21021;
  assign n21024 = ~n21022 & ~n21023;
  assign n21025 = n20947 & ~n21024;
  assign n21026 = ~n20947 & n21024;
  assign n21027 = ~n21025 & ~n21026;
  assign n21028 = pi103  & n8137;
  assign n21029 = pi101  & n8471;
  assign n21030 = pi102  & n8132;
  assign n21031 = ~n21029 & ~n21030;
  assign n21032 = ~n21028 & n21031;
  assign n21033 = n5540 & n8140;
  assign n21034 = n21032 & ~n21033;
  assign n21035 = pi50  & ~n21034;
  assign n21036 = pi50  & ~n21035;
  assign n21037 = ~n21034 & ~n21035;
  assign n21038 = ~n21036 & ~n21037;
  assign n21039 = n21027 & ~n21038;
  assign n21040 = ~n21027 & n21038;
  assign n21041 = ~n21039 & ~n21040;
  assign n21042 = n20946 & ~n21041;
  assign n21043 = ~n20946 & n21041;
  assign n21044 = ~n21042 & ~n21043;
  assign n21045 = pi106  & n7239;
  assign n21046 = pi104  & n7556;
  assign n21047 = pi105  & n7234;
  assign n21048 = ~n21046 & ~n21047;
  assign n21049 = ~n21045 & n21048;
  assign n21050 = n6090 & n7242;
  assign n21051 = n21049 & ~n21050;
  assign n21052 = pi47  & ~n21051;
  assign n21053 = pi47  & ~n21052;
  assign n21054 = ~n21051 & ~n21052;
  assign n21055 = ~n21053 & ~n21054;
  assign n21056 = n21044 & ~n21055;
  assign n21057 = ~n21044 & n21055;
  assign n21058 = ~n21056 & ~n21057;
  assign n21059 = n20945 & ~n21058;
  assign n21060 = ~n20945 & n21058;
  assign n21061 = ~n21059 & ~n21060;
  assign n21062 = pi109  & n6396;
  assign n21063 = pi107  & n6735;
  assign n21064 = pi108  & n6391;
  assign n21065 = ~n21063 & ~n21064;
  assign n21066 = ~n21062 & n21065;
  assign n21067 = n6399 & n7170;
  assign n21068 = n21066 & ~n21067;
  assign n21069 = pi44  & ~n21068;
  assign n21070 = pi44  & ~n21069;
  assign n21071 = ~n21068 & ~n21069;
  assign n21072 = ~n21070 & ~n21071;
  assign n21073 = ~n21061 & ~n21072;
  assign n21074 = n21061 & n21072;
  assign n21075 = ~n21073 & ~n21074;
  assign n21076 = n20944 & ~n21075;
  assign n21077 = ~n20944 & n21075;
  assign n21078 = ~n21076 & ~n21077;
  assign n21079 = pi112  & n5636;
  assign n21080 = pi110  & n5909;
  assign n21081 = pi111  & n5631;
  assign n21082 = ~n21080 & ~n21081;
  assign n21083 = ~n21079 & n21082;
  assign n21084 = n5639 & n7795;
  assign n21085 = n21083 & ~n21084;
  assign n21086 = pi41  & ~n21085;
  assign n21087 = pi41  & ~n21086;
  assign n21088 = ~n21085 & ~n21086;
  assign n21089 = ~n21087 & ~n21088;
  assign n21090 = n21078 & ~n21089;
  assign n21091 = ~n21078 & n21089;
  assign n21092 = ~n21090 & ~n21091;
  assign n21093 = n20943 & ~n21092;
  assign n21094 = ~n20943 & n21092;
  assign n21095 = ~n21093 & ~n21094;
  assign n21096 = pi115  & n4896;
  assign n21097 = pi113  & n5148;
  assign n21098 = pi114  & n4891;
  assign n21099 = ~n21097 & ~n21098;
  assign n21100 = ~n21096 & n21099;
  assign n21101 = n4899 & n8727;
  assign n21102 = n21100 & ~n21101;
  assign n21103 = pi38  & ~n21102;
  assign n21104 = pi38  & ~n21103;
  assign n21105 = ~n21102 & ~n21103;
  assign n21106 = ~n21104 & ~n21105;
  assign n21107 = n21095 & ~n21106;
  assign n21108 = ~n21095 & n21106;
  assign n21109 = ~n20942 & ~n21108;
  assign n21110 = ~n21107 & n21109;
  assign n21111 = ~n20942 & ~n21110;
  assign n21112 = ~n21107 & ~n21110;
  assign n21113 = ~n21108 & n21112;
  assign n21114 = ~n21111 & ~n21113;
  assign n21115 = pi118  & n4182;
  assign n21116 = pi116  & n4416;
  assign n21117 = pi117  & n4177;
  assign n21118 = ~n21116 & ~n21117;
  assign n21119 = ~n21115 & n21118;
  assign n21120 = n4185 & n9716;
  assign n21121 = n21119 & ~n21120;
  assign n21122 = pi35  & ~n21121;
  assign n21123 = pi35  & ~n21122;
  assign n21124 = ~n21121 & ~n21122;
  assign n21125 = ~n21123 & ~n21124;
  assign n21126 = n21114 & n21125;
  assign n21127 = ~n21114 & ~n21125;
  assign n21128 = ~n21126 & ~n21127;
  assign n21129 = ~n20941 & n21128;
  assign n21130 = n20941 & ~n21128;
  assign n21131 = ~n21129 & ~n21130;
  assign n21132 = n20940 & n21131;
  assign n21133 = ~n20940 & ~n21131;
  assign n21134 = ~n20925 & ~n21133;
  assign n21135 = ~n21132 & n21134;
  assign n21136 = ~n20925 & ~n21135;
  assign n21137 = ~n21133 & ~n21135;
  assign n21138 = ~n21132 & n21137;
  assign n21139 = ~n21136 & ~n21138;
  assign n21140 = ~n20910 & ~n21139;
  assign n21141 = n20910 & n21139;
  assign n21142 = ~n21140 & ~n21141;
  assign n21143 = ~n20894 & n21142;
  assign n21144 = n20894 & ~n21142;
  assign n21145 = ~n21143 & ~n21144;
  assign n21146 = ~n20893 & n21145;
  assign n21147 = n20893 & ~n21145;
  assign po87  = ~n21146 & ~n21147;
  assign n21149 = ~n21143 & ~n21146;
  assign n21150 = ~n20907 & ~n21140;
  assign n21151 = ~n21127 & ~n21129;
  assign n21152 = pi122  & n3550;
  assign n21153 = pi120  & n3735;
  assign n21154 = pi121  & n3545;
  assign n21155 = ~n21153 & ~n21154;
  assign n21156 = ~n21152 & n21155;
  assign n21157 = ~n3553 & n21156;
  assign n21158 = ~n11463 & n21156;
  assign n21159 = ~n21157 & ~n21158;
  assign n21160 = pi32  & ~n21159;
  assign n21161 = ~pi32  & n21159;
  assign n21162 = ~n21160 & ~n21161;
  assign n21163 = ~n21151 & ~n21162;
  assign n21164 = n21151 & n21162;
  assign n21165 = ~n21163 & ~n21164;
  assign n21166 = pi119  & n4182;
  assign n21167 = pi117  & n4416;
  assign n21168 = pi118  & n4177;
  assign n21169 = ~n21167 & ~n21168;
  assign n21170 = ~n21166 & n21169;
  assign n21171 = n4185 & n10048;
  assign n21172 = n21170 & ~n21171;
  assign n21173 = pi35  & ~n21172;
  assign n21174 = pi35  & ~n21173;
  assign n21175 = ~n21172 & ~n21173;
  assign n21176 = ~n21174 & ~n21175;
  assign n21177 = ~n21090 & ~n21094;
  assign n21178 = ~n21073 & ~n21077;
  assign n21179 = ~n21039 & ~n21043;
  assign n21180 = pi104  & n8137;
  assign n21181 = pi102  & n8471;
  assign n21182 = pi103  & n8132;
  assign n21183 = ~n21181 & ~n21182;
  assign n21184 = ~n21180 & n21183;
  assign n21185 = n5565 & n8140;
  assign n21186 = n21184 & ~n21185;
  assign n21187 = pi50  & ~n21186;
  assign n21188 = pi50  & ~n21187;
  assign n21189 = ~n21186 & ~n21187;
  assign n21190 = ~n21188 & ~n21189;
  assign n21191 = ~n21022 & ~n21026;
  assign n21192 = ~n21005 & ~n21008;
  assign n21193 = ~n20987 & ~n20991;
  assign n21194 = pi88  & n13477;
  assign n21195 = pi89  & ~n13122;
  assign n21196 = ~n21194 & ~n21195;
  assign n21197 = ~n20953 & ~n20956;
  assign n21198 = ~n21196 & n21197;
  assign n21199 = n21196 & ~n21197;
  assign n21200 = ~n21198 & ~n21199;
  assign n21201 = pi92  & n12295;
  assign n21202 = pi90  & n12693;
  assign n21203 = pi91  & n12290;
  assign n21204 = ~n21202 & ~n21203;
  assign n21205 = ~n21201 & n21204;
  assign n21206 = ~n12298 & n21205;
  assign n21207 = ~n3119 & n21205;
  assign n21208 = ~n21206 & ~n21207;
  assign n21209 = pi62  & ~n21208;
  assign n21210 = ~pi62  & n21208;
  assign n21211 = ~n21209 & ~n21210;
  assign n21212 = n21200 & ~n21211;
  assign n21213 = ~n21200 & n21211;
  assign n21214 = ~n21212 & ~n21213;
  assign n21215 = ~n20971 & ~n20974;
  assign n21216 = n21214 & n21215;
  assign n21217 = ~n21214 & ~n21215;
  assign n21218 = ~n21216 & ~n21217;
  assign n21219 = pi95  & n11193;
  assign n21220 = pi93  & n11567;
  assign n21221 = pi94  & n11188;
  assign n21222 = ~n21220 & ~n21221;
  assign n21223 = ~n21219 & n21222;
  assign n21224 = n3710 & n11196;
  assign n21225 = n21223 & ~n21224;
  assign n21226 = pi59  & ~n21225;
  assign n21227 = pi59  & ~n21226;
  assign n21228 = ~n21225 & ~n21226;
  assign n21229 = ~n21227 & ~n21228;
  assign n21230 = n21218 & ~n21229;
  assign n21231 = ~n21218 & n21229;
  assign n21232 = ~n21230 & ~n21231;
  assign n21233 = n21193 & ~n21232;
  assign n21234 = ~n21193 & n21232;
  assign n21235 = ~n21233 & ~n21234;
  assign n21236 = pi98  & n10135;
  assign n21237 = pi96  & n10478;
  assign n21238 = pi97  & n10130;
  assign n21239 = ~n21237 & ~n21238;
  assign n21240 = ~n21236 & n21239;
  assign n21241 = n4360 & n10138;
  assign n21242 = n21240 & ~n21241;
  assign n21243 = pi56  & ~n21242;
  assign n21244 = pi56  & ~n21243;
  assign n21245 = ~n21242 & ~n21243;
  assign n21246 = ~n21244 & ~n21245;
  assign n21247 = n21235 & ~n21246;
  assign n21248 = ~n21235 & n21246;
  assign n21249 = ~n21247 & ~n21248;
  assign n21250 = n21192 & ~n21249;
  assign n21251 = ~n21192 & n21249;
  assign n21252 = ~n21250 & ~n21251;
  assign n21253 = pi101  & n9096;
  assign n21254 = pi99  & n9453;
  assign n21255 = pi100  & n9091;
  assign n21256 = ~n21254 & ~n21255;
  assign n21257 = ~n21253 & n21256;
  assign n21258 = n5056 & n9099;
  assign n21259 = n21257 & ~n21258;
  assign n21260 = pi53  & ~n21259;
  assign n21261 = pi53  & ~n21260;
  assign n21262 = ~n21259 & ~n21260;
  assign n21263 = ~n21261 & ~n21262;
  assign n21264 = ~n21252 & n21263;
  assign n21265 = n21252 & ~n21263;
  assign n21266 = ~n21264 & ~n21265;
  assign n21267 = ~n21191 & n21266;
  assign n21268 = n21191 & ~n21266;
  assign n21269 = ~n21267 & ~n21268;
  assign n21270 = ~n21190 & n21269;
  assign n21271 = n21190 & ~n21269;
  assign n21272 = ~n21270 & ~n21271;
  assign n21273 = ~n21179 & n21272;
  assign n21274 = n21179 & ~n21272;
  assign n21275 = ~n21273 & ~n21274;
  assign n21276 = pi107  & n7239;
  assign n21277 = pi105  & n7556;
  assign n21278 = pi106  & n7234;
  assign n21279 = ~n21277 & ~n21278;
  assign n21280 = ~n21276 & n21279;
  assign n21281 = n6614 & n7242;
  assign n21282 = n21280 & ~n21281;
  assign n21283 = pi47  & ~n21282;
  assign n21284 = pi47  & ~n21283;
  assign n21285 = ~n21282 & ~n21283;
  assign n21286 = ~n21284 & ~n21285;
  assign n21287 = n21275 & ~n21286;
  assign n21288 = ~n21275 & n21286;
  assign n21289 = ~n21287 & ~n21288;
  assign n21290 = ~n21057 & ~n21060;
  assign n21291 = ~n21289 & ~n21290;
  assign n21292 = n21289 & n21290;
  assign n21293 = ~n21291 & ~n21292;
  assign n21294 = pi110  & n6396;
  assign n21295 = pi108  & n6735;
  assign n21296 = pi109  & n6391;
  assign n21297 = ~n21295 & ~n21296;
  assign n21298 = ~n21294 & n21297;
  assign n21299 = n6399 & n7474;
  assign n21300 = n21298 & ~n21299;
  assign n21301 = pi44  & ~n21300;
  assign n21302 = pi44  & ~n21301;
  assign n21303 = ~n21300 & ~n21301;
  assign n21304 = ~n21302 & ~n21303;
  assign n21305 = n21293 & ~n21304;
  assign n21306 = ~n21293 & n21304;
  assign n21307 = ~n21305 & ~n21306;
  assign n21308 = n21178 & ~n21307;
  assign n21309 = ~n21178 & n21307;
  assign n21310 = ~n21308 & ~n21309;
  assign n21311 = pi113  & n5636;
  assign n21312 = pi111  & n5909;
  assign n21313 = pi112  & n5631;
  assign n21314 = ~n21312 & ~n21313;
  assign n21315 = ~n21311 & n21314;
  assign n21316 = n5639 & n8387;
  assign n21317 = n21315 & ~n21316;
  assign n21318 = pi41  & ~n21317;
  assign n21319 = pi41  & ~n21318;
  assign n21320 = ~n21317 & ~n21318;
  assign n21321 = ~n21319 & ~n21320;
  assign n21322 = n21310 & ~n21321;
  assign n21323 = ~n21310 & n21321;
  assign n21324 = ~n21322 & ~n21323;
  assign n21325 = n21177 & ~n21324;
  assign n21326 = ~n21177 & n21324;
  assign n21327 = ~n21325 & ~n21326;
  assign n21328 = pi116  & n4896;
  assign n21329 = pi114  & n5148;
  assign n21330 = pi115  & n4891;
  assign n21331 = ~n21329 & ~n21330;
  assign n21332 = ~n21328 & n21331;
  assign n21333 = n4899 & n9042;
  assign n21334 = n21332 & ~n21333;
  assign n21335 = pi38  & ~n21334;
  assign n21336 = pi38  & ~n21335;
  assign n21337 = ~n21334 & ~n21335;
  assign n21338 = ~n21336 & ~n21337;
  assign n21339 = n21327 & ~n21338;
  assign n21340 = ~n21327 & n21338;
  assign n21341 = ~n21339 & ~n21340;
  assign n21342 = ~n21112 & n21341;
  assign n21343 = n21112 & ~n21341;
  assign n21344 = ~n21342 & ~n21343;
  assign n21345 = ~n21176 & n21344;
  assign n21346 = n21176 & ~n21344;
  assign n21347 = ~n21345 & ~n21346;
  assign n21348 = n21165 & n21347;
  assign n21349 = ~n21165 & ~n21347;
  assign n21350 = ~n21348 & ~n21349;
  assign n21351 = pi125  & n2976;
  assign n21352 = pi123  & n3182;
  assign n21353 = pi124  & n2971;
  assign n21354 = ~n21352 & ~n21353;
  assign n21355 = ~n21351 & n21354;
  assign n21356 = n2979 & n12591;
  assign n21357 = n21355 & ~n21356;
  assign n21358 = pi29  & ~n21357;
  assign n21359 = pi29  & ~n21358;
  assign n21360 = ~n21357 & ~n21358;
  assign n21361 = ~n21359 & ~n21360;
  assign n21362 = ~n20939 & ~n21132;
  assign n21363 = ~n21361 & ~n21362;
  assign n21364 = n21361 & n21362;
  assign n21365 = ~n21363 & ~n21364;
  assign n21366 = n21350 & n21365;
  assign n21367 = ~n21350 & ~n21365;
  assign n21368 = ~n21366 & ~n21367;
  assign n21369 = ~n20911 & ~n20922;
  assign n21370 = ~n21135 & ~n21369;
  assign n21371 = pi126  & n2644;
  assign n21372 = pi127  & n2481;
  assign n21373 = ~n21371 & ~n21372;
  assign n21374 = ~n2489 & n21373;
  assign n21375 = ~n13389 & n21373;
  assign n21376 = ~n21374 & ~n21375;
  assign n21377 = pi26  & ~n21376;
  assign n21378 = ~pi26  & n21376;
  assign n21379 = ~n21377 & ~n21378;
  assign n21380 = ~n21370 & ~n21379;
  assign n21381 = n21370 & n21379;
  assign n21382 = ~n21380 & ~n21381;
  assign n21383 = n21368 & n21382;
  assign n21384 = ~n21368 & ~n21382;
  assign n21385 = ~n21383 & ~n21384;
  assign n21386 = ~n21150 & n21385;
  assign n21387 = n21150 & ~n21385;
  assign n21388 = ~n21386 & ~n21387;
  assign n21389 = ~n21149 & n21388;
  assign n21390 = n21149 & ~n21388;
  assign po88  = ~n21389 & ~n21390;
  assign n21392 = ~n21386 & ~n21389;
  assign n21393 = ~n21380 & ~n21383;
  assign n21394 = pi126  & n2976;
  assign n21395 = pi124  & n3182;
  assign n21396 = pi125  & n2971;
  assign n21397 = ~n21395 & ~n21396;
  assign n21398 = ~n21394 & n21397;
  assign n21399 = n2979 & n12979;
  assign n21400 = n21398 & ~n21399;
  assign n21401 = pi29  & ~n21400;
  assign n21402 = pi29  & ~n21401;
  assign n21403 = ~n21400 & ~n21401;
  assign n21404 = ~n21402 & ~n21403;
  assign n21405 = ~n21163 & ~n21348;
  assign n21406 = n21404 & n21405;
  assign n21407 = ~n21404 & ~n21405;
  assign n21408 = ~n21406 & ~n21407;
  assign n21409 = pi123  & n3550;
  assign n21410 = pi121  & n3735;
  assign n21411 = pi122  & n3545;
  assign n21412 = ~n21410 & ~n21411;
  assign n21413 = ~n21409 & n21412;
  assign n21414 = n3553 & n11489;
  assign n21415 = n21413 & ~n21414;
  assign n21416 = pi32  & ~n21415;
  assign n21417 = pi32  & ~n21416;
  assign n21418 = ~n21415 & ~n21416;
  assign n21419 = ~n21417 & ~n21418;
  assign n21420 = ~n21342 & ~n21345;
  assign n21421 = n21419 & n21420;
  assign n21422 = ~n21419 & ~n21420;
  assign n21423 = ~n21421 & ~n21422;
  assign n21424 = pi120  & n4182;
  assign n21425 = pi118  & n4416;
  assign n21426 = pi119  & n4177;
  assign n21427 = ~n21425 & ~n21426;
  assign n21428 = ~n21424 & n21427;
  assign n21429 = n4185 & n10734;
  assign n21430 = n21428 & ~n21429;
  assign n21431 = pi35  & ~n21430;
  assign n21432 = pi35  & ~n21431;
  assign n21433 = ~n21430 & ~n21431;
  assign n21434 = ~n21432 & ~n21433;
  assign n21435 = ~n21326 & ~n21339;
  assign n21436 = pi117  & n4896;
  assign n21437 = pi115  & n5148;
  assign n21438 = pi116  & n4891;
  assign n21439 = ~n21437 & ~n21438;
  assign n21440 = ~n21436 & n21439;
  assign n21441 = n4899 & n9691;
  assign n21442 = n21440 & ~n21441;
  assign n21443 = pi38  & ~n21442;
  assign n21444 = pi38  & ~n21443;
  assign n21445 = ~n21442 & ~n21443;
  assign n21446 = ~n21444 & ~n21445;
  assign n21447 = ~n21309 & ~n21322;
  assign n21448 = ~n21273 & ~n21287;
  assign n21449 = pi108  & n7239;
  assign n21450 = pi106  & n7556;
  assign n21451 = pi107  & n7234;
  assign n21452 = ~n21450 & ~n21451;
  assign n21453 = ~n21449 & n21452;
  assign n21454 = n6639 & n7242;
  assign n21455 = n21453 & ~n21454;
  assign n21456 = pi47  & ~n21455;
  assign n21457 = pi47  & ~n21456;
  assign n21458 = ~n21455 & ~n21456;
  assign n21459 = ~n21457 & ~n21458;
  assign n21460 = ~n21267 & ~n21270;
  assign n21461 = pi105  & n8137;
  assign n21462 = pi103  & n8471;
  assign n21463 = pi104  & n8132;
  assign n21464 = ~n21462 & ~n21463;
  assign n21465 = ~n21461 & n21464;
  assign n21466 = n6065 & n8140;
  assign n21467 = n21465 & ~n21466;
  assign n21468 = pi50  & ~n21467;
  assign n21469 = pi50  & ~n21468;
  assign n21470 = ~n21467 & ~n21468;
  assign n21471 = ~n21469 & ~n21470;
  assign n21472 = ~n21234 & ~n21247;
  assign n21473 = pi99  & n10135;
  assign n21474 = pi97  & n10478;
  assign n21475 = pi98  & n10130;
  assign n21476 = ~n21474 & ~n21475;
  assign n21477 = ~n21473 & n21476;
  assign n21478 = n4584 & n10138;
  assign n21479 = n21477 & ~n21478;
  assign n21480 = pi56  & ~n21479;
  assign n21481 = pi56  & ~n21480;
  assign n21482 = ~n21479 & ~n21480;
  assign n21483 = ~n21481 & ~n21482;
  assign n21484 = ~n21216 & ~n21230;
  assign n21485 = pi96  & n11193;
  assign n21486 = pi94  & n11567;
  assign n21487 = pi95  & n11188;
  assign n21488 = ~n21486 & ~n21487;
  assign n21489 = ~n21485 & n21488;
  assign n21490 = n3921 & n11196;
  assign n21491 = n21489 & ~n21490;
  assign n21492 = pi59  & ~n21491;
  assign n21493 = pi59  & ~n21492;
  assign n21494 = ~n21491 & ~n21492;
  assign n21495 = ~n21493 & ~n21494;
  assign n21496 = ~n21199 & ~n21212;
  assign n21497 = pi89  & n13477;
  assign n21498 = pi90  & ~n13122;
  assign n21499 = ~n21497 & ~n21498;
  assign n21500 = ~n21196 & n21499;
  assign n21501 = n21196 & ~n21499;
  assign n21502 = ~n21500 & ~n21501;
  assign n21503 = pi93  & n12295;
  assign n21504 = pi91  & n12693;
  assign n21505 = pi92  & n12290;
  assign n21506 = ~n21504 & ~n21505;
  assign n21507 = ~n21503 & n21506;
  assign n21508 = ~n12298 & n21507;
  assign n21509 = ~n3144 & n21507;
  assign n21510 = ~n21508 & ~n21509;
  assign n21511 = pi62  & ~n21510;
  assign n21512 = ~pi62  & n21510;
  assign n21513 = ~n21511 & ~n21512;
  assign n21514 = n21502 & ~n21513;
  assign n21515 = ~n21502 & n21513;
  assign n21516 = ~n21514 & ~n21515;
  assign n21517 = ~n21496 & n21516;
  assign n21518 = n21496 & ~n21516;
  assign n21519 = ~n21517 & ~n21518;
  assign n21520 = ~n21495 & n21519;
  assign n21521 = n21495 & ~n21519;
  assign n21522 = ~n21520 & ~n21521;
  assign n21523 = ~n21484 & n21522;
  assign n21524 = n21484 & ~n21522;
  assign n21525 = ~n21523 & ~n21524;
  assign n21526 = ~n21483 & n21525;
  assign n21527 = n21483 & ~n21525;
  assign n21528 = ~n21526 & ~n21527;
  assign n21529 = ~n21472 & n21528;
  assign n21530 = n21472 & ~n21528;
  assign n21531 = ~n21529 & ~n21530;
  assign n21532 = pi102  & n9096;
  assign n21533 = pi100  & n9453;
  assign n21534 = pi101  & n9091;
  assign n21535 = ~n21533 & ~n21534;
  assign n21536 = ~n21532 & n21535;
  assign n21537 = n5296 & n9099;
  assign n21538 = n21536 & ~n21537;
  assign n21539 = pi53  & ~n21538;
  assign n21540 = pi53  & ~n21539;
  assign n21541 = ~n21538 & ~n21539;
  assign n21542 = ~n21540 & ~n21541;
  assign n21543 = n21531 & ~n21542;
  assign n21544 = n21531 & ~n21543;
  assign n21545 = ~n21542 & ~n21543;
  assign n21546 = ~n21544 & ~n21545;
  assign n21547 = ~n21251 & ~n21265;
  assign n21548 = ~n21546 & ~n21547;
  assign n21549 = n21546 & n21547;
  assign n21550 = ~n21548 & ~n21549;
  assign n21551 = n21471 & n21550;
  assign n21552 = ~n21471 & ~n21550;
  assign n21553 = ~n21551 & ~n21552;
  assign n21554 = ~n21460 & ~n21553;
  assign n21555 = n21460 & n21553;
  assign n21556 = ~n21554 & ~n21555;
  assign n21557 = ~n21459 & n21556;
  assign n21558 = n21459 & ~n21556;
  assign n21559 = ~n21557 & ~n21558;
  assign n21560 = ~n21448 & n21559;
  assign n21561 = n21448 & ~n21559;
  assign n21562 = ~n21560 & ~n21561;
  assign n21563 = pi111  & n6396;
  assign n21564 = pi109  & n6735;
  assign n21565 = pi110  & n6391;
  assign n21566 = ~n21564 & ~n21565;
  assign n21567 = ~n21563 & n21566;
  assign n21568 = n6399 & n7770;
  assign n21569 = n21567 & ~n21568;
  assign n21570 = pi44  & ~n21569;
  assign n21571 = pi44  & ~n21570;
  assign n21572 = ~n21569 & ~n21570;
  assign n21573 = ~n21571 & ~n21572;
  assign n21574 = n21562 & ~n21573;
  assign n21575 = n21562 & ~n21574;
  assign n21576 = ~n21573 & ~n21574;
  assign n21577 = ~n21575 & ~n21576;
  assign n21578 = ~n21292 & ~n21305;
  assign n21579 = n21577 & n21578;
  assign n21580 = ~n21577 & ~n21578;
  assign n21581 = ~n21579 & ~n21580;
  assign n21582 = pi114  & n5636;
  assign n21583 = pi112  & n5909;
  assign n21584 = pi113  & n5631;
  assign n21585 = ~n21583 & ~n21584;
  assign n21586 = ~n21582 & n21585;
  assign n21587 = n5639 & n8702;
  assign n21588 = n21586 & ~n21587;
  assign n21589 = pi41  & ~n21588;
  assign n21590 = pi41  & ~n21589;
  assign n21591 = ~n21588 & ~n21589;
  assign n21592 = ~n21590 & ~n21591;
  assign n21593 = ~n21581 & n21592;
  assign n21594 = n21581 & ~n21592;
  assign n21595 = ~n21593 & ~n21594;
  assign n21596 = ~n21447 & n21595;
  assign n21597 = n21447 & ~n21595;
  assign n21598 = ~n21596 & ~n21597;
  assign n21599 = ~n21446 & n21598;
  assign n21600 = n21446 & ~n21598;
  assign n21601 = ~n21599 & ~n21600;
  assign n21602 = ~n21435 & n21601;
  assign n21603 = n21435 & ~n21601;
  assign n21604 = ~n21602 & ~n21603;
  assign n21605 = ~n21434 & n21604;
  assign n21606 = n21434 & ~n21604;
  assign n21607 = ~n21605 & ~n21606;
  assign n21608 = n21423 & n21607;
  assign n21609 = ~n21423 & ~n21607;
  assign n21610 = ~n21608 & ~n21609;
  assign n21611 = ~n21408 & ~n21610;
  assign n21612 = n21408 & n21610;
  assign n21613 = ~n21611 & ~n21612;
  assign n21614 = ~n21363 & ~n21366;
  assign n21615 = pi127  & n2644;
  assign n21616 = n2489 & n13387;
  assign n21617 = ~n21615 & ~n21616;
  assign n21618 = pi26  & ~n21617;
  assign n21619 = pi26  & ~n21618;
  assign n21620 = ~n21617 & ~n21618;
  assign n21621 = ~n21619 & ~n21620;
  assign n21622 = ~n21614 & ~n21621;
  assign n21623 = n21614 & n21621;
  assign n21624 = ~n21622 & ~n21623;
  assign n21625 = n21613 & n21624;
  assign n21626 = ~n21613 & ~n21624;
  assign n21627 = ~n21625 & ~n21626;
  assign n21628 = ~n21393 & n21627;
  assign n21629 = n21393 & ~n21627;
  assign n21630 = ~n21628 & ~n21629;
  assign n21631 = ~n21392 & n21630;
  assign n21632 = n21392 & ~n21630;
  assign po89  = ~n21631 & ~n21632;
  assign n21634 = ~n21622 & ~n21625;
  assign n21635 = ~n21407 & ~n21612;
  assign n21636 = pi127  & n2976;
  assign n21637 = pi125  & n3182;
  assign n21638 = pi126  & n2971;
  assign n21639 = ~n21637 & ~n21638;
  assign n21640 = ~n21636 & n21639;
  assign n21641 = n2979 & n13365;
  assign n21642 = n21640 & ~n21641;
  assign n21643 = pi29  & ~n21642;
  assign n21644 = pi29  & ~n21643;
  assign n21645 = ~n21642 & ~n21643;
  assign n21646 = ~n21644 & ~n21645;
  assign n21647 = ~n21635 & ~n21646;
  assign n21648 = ~n21635 & ~n21647;
  assign n21649 = ~n21646 & ~n21647;
  assign n21650 = ~n21648 & ~n21649;
  assign n21651 = ~n21602 & ~n21605;
  assign n21652 = ~n21596 & ~n21599;
  assign n21653 = ~n21580 & ~n21594;
  assign n21654 = ~n21560 & ~n21574;
  assign n21655 = ~n21554 & ~n21557;
  assign n21656 = pi109  & n7239;
  assign n21657 = pi107  & n7556;
  assign n21658 = pi108  & n7234;
  assign n21659 = ~n21657 & ~n21658;
  assign n21660 = ~n21656 & n21659;
  assign n21661 = n7170 & n7242;
  assign n21662 = n21660 & ~n21661;
  assign n21663 = pi47  & ~n21662;
  assign n21664 = pi47  & ~n21663;
  assign n21665 = ~n21662 & ~n21663;
  assign n21666 = ~n21664 & ~n21665;
  assign n21667 = ~n21549 & ~n21551;
  assign n21668 = ~n21523 & ~n21526;
  assign n21669 = pi97  & n11193;
  assign n21670 = pi95  & n11567;
  assign n21671 = pi96  & n11188;
  assign n21672 = ~n21670 & ~n21671;
  assign n21673 = ~n21669 & n21672;
  assign n21674 = n3946 & n11196;
  assign n21675 = n21673 & ~n21674;
  assign n21676 = pi59  & ~n21675;
  assign n21677 = pi59  & ~n21676;
  assign n21678 = ~n21675 & ~n21676;
  assign n21679 = ~n21677 & ~n21678;
  assign n21680 = ~n21517 & ~n21520;
  assign n21681 = n21679 & n21680;
  assign n21682 = ~n21679 & ~n21680;
  assign n21683 = ~n21681 & ~n21682;
  assign n21684 = ~n21500 & ~n21514;
  assign n21685 = pi90  & n13477;
  assign n21686 = pi91  & ~n13122;
  assign n21687 = ~n21685 & ~n21686;
  assign n21688 = ~pi26  & ~n21687;
  assign n21689 = pi26  & n21687;
  assign n21690 = ~n21688 & ~n21689;
  assign n21691 = ~n21499 & n21690;
  assign n21692 = n21499 & ~n21690;
  assign n21693 = ~n21691 & ~n21692;
  assign n21694 = ~n21684 & n21693;
  assign n21695 = n21684 & ~n21693;
  assign n21696 = ~n21694 & ~n21695;
  assign n21697 = pi94  & n12295;
  assign n21698 = pi92  & n12693;
  assign n21699 = pi93  & n12290;
  assign n21700 = ~n21698 & ~n21699;
  assign n21701 = ~n21697 & n21700;
  assign n21702 = n3499 & n12298;
  assign n21703 = n21701 & ~n21702;
  assign n21704 = pi62  & ~n21703;
  assign n21705 = pi62  & ~n21704;
  assign n21706 = ~n21703 & ~n21704;
  assign n21707 = ~n21705 & ~n21706;
  assign n21708 = n21696 & ~n21707;
  assign n21709 = n21696 & ~n21708;
  assign n21710 = ~n21707 & ~n21708;
  assign n21711 = ~n21709 & ~n21710;
  assign n21712 = ~n21683 & n21711;
  assign n21713 = n21683 & ~n21711;
  assign n21714 = ~n21712 & ~n21713;
  assign n21715 = pi100  & n10135;
  assign n21716 = pi98  & n10478;
  assign n21717 = pi99  & n10130;
  assign n21718 = ~n21716 & ~n21717;
  assign n21719 = ~n21715 & n21718;
  assign n21720 = n4808 & n10138;
  assign n21721 = n21719 & ~n21720;
  assign n21722 = pi56  & ~n21721;
  assign n21723 = pi56  & ~n21722;
  assign n21724 = ~n21721 & ~n21722;
  assign n21725 = ~n21723 & ~n21724;
  assign n21726 = n21714 & ~n21725;
  assign n21727 = ~n21714 & n21725;
  assign n21728 = ~n21726 & ~n21727;
  assign n21729 = n21668 & ~n21728;
  assign n21730 = ~n21668 & n21728;
  assign n21731 = ~n21729 & ~n21730;
  assign n21732 = pi103  & n9096;
  assign n21733 = pi101  & n9453;
  assign n21734 = pi102  & n9091;
  assign n21735 = ~n21733 & ~n21734;
  assign n21736 = ~n21732 & n21735;
  assign n21737 = n5540 & n9099;
  assign n21738 = n21736 & ~n21737;
  assign n21739 = pi53  & ~n21738;
  assign n21740 = pi53  & ~n21739;
  assign n21741 = ~n21738 & ~n21739;
  assign n21742 = ~n21740 & ~n21741;
  assign n21743 = n21731 & ~n21742;
  assign n21744 = n21731 & ~n21743;
  assign n21745 = ~n21742 & ~n21743;
  assign n21746 = ~n21744 & ~n21745;
  assign n21747 = ~n21529 & ~n21543;
  assign n21748 = n21746 & n21747;
  assign n21749 = ~n21746 & ~n21747;
  assign n21750 = ~n21748 & ~n21749;
  assign n21751 = pi106  & n8137;
  assign n21752 = pi104  & n8471;
  assign n21753 = pi105  & n8132;
  assign n21754 = ~n21752 & ~n21753;
  assign n21755 = ~n21751 & n21754;
  assign n21756 = n6090 & n8140;
  assign n21757 = n21755 & ~n21756;
  assign n21758 = pi50  & ~n21757;
  assign n21759 = pi50  & ~n21758;
  assign n21760 = ~n21757 & ~n21758;
  assign n21761 = ~n21759 & ~n21760;
  assign n21762 = n21750 & ~n21761;
  assign n21763 = ~n21750 & n21761;
  assign n21764 = ~n21762 & ~n21763;
  assign n21765 = n21667 & n21764;
  assign n21766 = ~n21667 & ~n21764;
  assign n21767 = ~n21765 & ~n21766;
  assign n21768 = ~n21666 & n21767;
  assign n21769 = n21666 & ~n21767;
  assign n21770 = ~n21768 & ~n21769;
  assign n21771 = n21655 & ~n21770;
  assign n21772 = ~n21655 & n21770;
  assign n21773 = ~n21771 & ~n21772;
  assign n21774 = pi112  & n6396;
  assign n21775 = pi110  & n6735;
  assign n21776 = pi111  & n6391;
  assign n21777 = ~n21775 & ~n21776;
  assign n21778 = ~n21774 & n21777;
  assign n21779 = n6399 & n7795;
  assign n21780 = n21778 & ~n21779;
  assign n21781 = pi44  & ~n21780;
  assign n21782 = pi44  & ~n21781;
  assign n21783 = ~n21780 & ~n21781;
  assign n21784 = ~n21782 & ~n21783;
  assign n21785 = n21773 & ~n21784;
  assign n21786 = ~n21773 & n21784;
  assign n21787 = ~n21785 & ~n21786;
  assign n21788 = n21654 & ~n21787;
  assign n21789 = ~n21654 & n21787;
  assign n21790 = ~n21788 & ~n21789;
  assign n21791 = pi115  & n5636;
  assign n21792 = pi113  & n5909;
  assign n21793 = pi114  & n5631;
  assign n21794 = ~n21792 & ~n21793;
  assign n21795 = ~n21791 & n21794;
  assign n21796 = n5639 & n8727;
  assign n21797 = n21795 & ~n21796;
  assign n21798 = pi41  & ~n21797;
  assign n21799 = pi41  & ~n21798;
  assign n21800 = ~n21797 & ~n21798;
  assign n21801 = ~n21799 & ~n21800;
  assign n21802 = n21790 & ~n21801;
  assign n21803 = ~n21790 & n21801;
  assign n21804 = ~n21653 & ~n21803;
  assign n21805 = ~n21802 & n21804;
  assign n21806 = ~n21653 & ~n21805;
  assign n21807 = ~n21802 & ~n21805;
  assign n21808 = ~n21803 & n21807;
  assign n21809 = ~n21806 & ~n21808;
  assign n21810 = pi118  & n4896;
  assign n21811 = pi116  & n5148;
  assign n21812 = pi117  & n4891;
  assign n21813 = ~n21811 & ~n21812;
  assign n21814 = ~n21810 & n21813;
  assign n21815 = n4899 & n9716;
  assign n21816 = n21814 & ~n21815;
  assign n21817 = pi38  & ~n21816;
  assign n21818 = pi38  & ~n21817;
  assign n21819 = ~n21816 & ~n21817;
  assign n21820 = ~n21818 & ~n21819;
  assign n21821 = n21809 & n21820;
  assign n21822 = ~n21809 & ~n21820;
  assign n21823 = ~n21821 & ~n21822;
  assign n21824 = ~n21652 & n21823;
  assign n21825 = n21652 & ~n21823;
  assign n21826 = ~n21824 & ~n21825;
  assign n21827 = pi121  & n4182;
  assign n21828 = pi119  & n4416;
  assign n21829 = pi120  & n4177;
  assign n21830 = ~n21828 & ~n21829;
  assign n21831 = ~n21827 & n21830;
  assign n21832 = n4185 & n11086;
  assign n21833 = n21831 & ~n21832;
  assign n21834 = pi35  & ~n21833;
  assign n21835 = pi35  & ~n21834;
  assign n21836 = ~n21833 & ~n21834;
  assign n21837 = ~n21835 & ~n21836;
  assign n21838 = n21826 & ~n21837;
  assign n21839 = ~n21826 & n21837;
  assign n21840 = ~n21838 & ~n21839;
  assign n21841 = n21651 & ~n21840;
  assign n21842 = ~n21651 & n21840;
  assign n21843 = ~n21841 & ~n21842;
  assign n21844 = pi124  & n3550;
  assign n21845 = pi122  & n3735;
  assign n21846 = pi123  & n3545;
  assign n21847 = ~n21845 & ~n21846;
  assign n21848 = ~n21844 & n21847;
  assign n21849 = n3553 & n11858;
  assign n21850 = n21848 & ~n21849;
  assign n21851 = pi32  & ~n21850;
  assign n21852 = pi32  & ~n21851;
  assign n21853 = ~n21850 & ~n21851;
  assign n21854 = ~n21852 & ~n21853;
  assign n21855 = ~n21422 & ~n21608;
  assign n21856 = n21854 & n21855;
  assign n21857 = ~n21854 & ~n21855;
  assign n21858 = ~n21856 & ~n21857;
  assign n21859 = n21843 & n21858;
  assign n21860 = ~n21843 & ~n21858;
  assign n21861 = ~n21859 & ~n21860;
  assign n21862 = ~n21650 & n21861;
  assign n21863 = n21650 & ~n21861;
  assign n21864 = ~n21862 & ~n21863;
  assign n21865 = n21634 & ~n21864;
  assign n21866 = ~n21634 & n21864;
  assign n21867 = ~n21865 & ~n21866;
  assign n21868 = ~n21628 & ~n21631;
  assign n21869 = n21867 & ~n21868;
  assign n21870 = ~n21867 & n21868;
  assign po90  = ~n21869 & ~n21870;
  assign n21872 = ~n21857 & ~n21859;
  assign n21873 = pi126  & n3182;
  assign n21874 = pi127  & n2971;
  assign n21875 = ~n21873 & ~n21874;
  assign n21876 = ~n2979 & n21875;
  assign n21877 = ~n13389 & n21875;
  assign n21878 = ~n21876 & ~n21877;
  assign n21879 = pi29  & ~n21878;
  assign n21880 = ~pi29  & n21878;
  assign n21881 = ~n21879 & ~n21880;
  assign n21882 = ~n21872 & ~n21881;
  assign n21883 = n21872 & n21881;
  assign n21884 = ~n21882 & ~n21883;
  assign n21885 = pi125  & n3550;
  assign n21886 = pi123  & n3735;
  assign n21887 = pi124  & n3545;
  assign n21888 = ~n21886 & ~n21887;
  assign n21889 = ~n21885 & n21888;
  assign n21890 = n3553 & n12591;
  assign n21891 = n21889 & ~n21890;
  assign n21892 = pi32  & ~n21891;
  assign n21893 = pi32  & ~n21892;
  assign n21894 = ~n21891 & ~n21892;
  assign n21895 = ~n21893 & ~n21894;
  assign n21896 = ~n21838 & ~n21842;
  assign n21897 = n21895 & n21896;
  assign n21898 = ~n21895 & ~n21896;
  assign n21899 = ~n21897 & ~n21898;
  assign n21900 = ~n21822 & ~n21824;
  assign n21901 = pi119  & n4896;
  assign n21902 = pi117  & n5148;
  assign n21903 = pi118  & n4891;
  assign n21904 = ~n21902 & ~n21903;
  assign n21905 = ~n21901 & n21904;
  assign n21906 = n4899 & n10048;
  assign n21907 = n21905 & ~n21906;
  assign n21908 = pi38  & ~n21907;
  assign n21909 = pi38  & ~n21908;
  assign n21910 = ~n21907 & ~n21908;
  assign n21911 = ~n21909 & ~n21910;
  assign n21912 = ~n21785 & ~n21789;
  assign n21913 = ~n21768 & ~n21772;
  assign n21914 = ~n21762 & ~n21765;
  assign n21915 = ~n21743 & ~n21749;
  assign n21916 = pi104  & n9096;
  assign n21917 = pi102  & n9453;
  assign n21918 = pi103  & n9091;
  assign n21919 = ~n21917 & ~n21918;
  assign n21920 = ~n21916 & n21919;
  assign n21921 = n5565 & n9099;
  assign n21922 = n21920 & ~n21921;
  assign n21923 = pi53  & ~n21922;
  assign n21924 = pi53  & ~n21923;
  assign n21925 = ~n21922 & ~n21923;
  assign n21926 = ~n21924 & ~n21925;
  assign n21927 = ~n21726 & ~n21730;
  assign n21928 = pi101  & n10135;
  assign n21929 = pi99  & n10478;
  assign n21930 = pi100  & n10130;
  assign n21931 = ~n21929 & ~n21930;
  assign n21932 = ~n21928 & n21931;
  assign n21933 = n5056 & n10138;
  assign n21934 = n21932 & ~n21933;
  assign n21935 = pi56  & ~n21934;
  assign n21936 = pi56  & ~n21935;
  assign n21937 = ~n21934 & ~n21935;
  assign n21938 = ~n21936 & ~n21937;
  assign n21939 = pi91  & n13477;
  assign n21940 = pi92  & ~n13122;
  assign n21941 = ~n21939 & ~n21940;
  assign n21942 = ~n21688 & ~n21691;
  assign n21943 = ~n21941 & n21942;
  assign n21944 = n21941 & ~n21942;
  assign n21945 = ~n21943 & ~n21944;
  assign n21946 = pi95  & n12295;
  assign n21947 = pi93  & n12693;
  assign n21948 = pi94  & n12290;
  assign n21949 = ~n21947 & ~n21948;
  assign n21950 = ~n21946 & n21949;
  assign n21951 = n3710 & n12298;
  assign n21952 = n21950 & ~n21951;
  assign n21953 = pi62  & ~n21952;
  assign n21954 = pi62  & ~n21953;
  assign n21955 = ~n21952 & ~n21953;
  assign n21956 = ~n21954 & ~n21955;
  assign n21957 = ~n21945 & n21956;
  assign n21958 = n21945 & ~n21956;
  assign n21959 = ~n21957 & ~n21958;
  assign n21960 = ~n21694 & ~n21708;
  assign n21961 = n21959 & ~n21960;
  assign n21962 = ~n21959 & n21960;
  assign n21963 = ~n21961 & ~n21962;
  assign n21964 = pi98  & n11193;
  assign n21965 = pi96  & n11567;
  assign n21966 = pi97  & n11188;
  assign n21967 = ~n21965 & ~n21966;
  assign n21968 = ~n21964 & n21967;
  assign n21969 = n4360 & n11196;
  assign n21970 = n21968 & ~n21969;
  assign n21971 = pi59  & ~n21970;
  assign n21972 = pi59  & ~n21971;
  assign n21973 = ~n21970 & ~n21971;
  assign n21974 = ~n21972 & ~n21973;
  assign n21975 = n21963 & ~n21974;
  assign n21976 = n21963 & ~n21975;
  assign n21977 = ~n21974 & ~n21975;
  assign n21978 = ~n21976 & ~n21977;
  assign n21979 = ~n21682 & ~n21713;
  assign n21980 = ~n21978 & ~n21979;
  assign n21981 = n21978 & n21979;
  assign n21982 = ~n21980 & ~n21981;
  assign n21983 = n21938 & n21982;
  assign n21984 = ~n21938 & ~n21982;
  assign n21985 = ~n21983 & ~n21984;
  assign n21986 = ~n21927 & ~n21985;
  assign n21987 = n21927 & n21985;
  assign n21988 = ~n21986 & ~n21987;
  assign n21989 = ~n21926 & n21988;
  assign n21990 = n21926 & ~n21988;
  assign n21991 = ~n21989 & ~n21990;
  assign n21992 = ~n21915 & n21991;
  assign n21993 = n21915 & ~n21991;
  assign n21994 = ~n21992 & ~n21993;
  assign n21995 = pi107  & n8137;
  assign n21996 = pi105  & n8471;
  assign n21997 = pi106  & n8132;
  assign n21998 = ~n21996 & ~n21997;
  assign n21999 = ~n21995 & n21998;
  assign n22000 = n6614 & n8140;
  assign n22001 = n21999 & ~n22000;
  assign n22002 = pi50  & ~n22001;
  assign n22003 = pi50  & ~n22002;
  assign n22004 = ~n22001 & ~n22002;
  assign n22005 = ~n22003 & ~n22004;
  assign n22006 = n21994 & ~n22005;
  assign n22007 = ~n21994 & n22005;
  assign n22008 = ~n22006 & ~n22007;
  assign n22009 = n21914 & ~n22008;
  assign n22010 = ~n21914 & n22008;
  assign n22011 = ~n22009 & ~n22010;
  assign n22012 = pi110  & n7239;
  assign n22013 = pi108  & n7556;
  assign n22014 = pi109  & n7234;
  assign n22015 = ~n22013 & ~n22014;
  assign n22016 = ~n22012 & n22015;
  assign n22017 = n7242 & n7474;
  assign n22018 = n22016 & ~n22017;
  assign n22019 = pi47  & ~n22018;
  assign n22020 = pi47  & ~n22019;
  assign n22021 = ~n22018 & ~n22019;
  assign n22022 = ~n22020 & ~n22021;
  assign n22023 = n22011 & ~n22022;
  assign n22024 = ~n22011 & n22022;
  assign n22025 = ~n22023 & ~n22024;
  assign n22026 = n21913 & ~n22025;
  assign n22027 = ~n21913 & n22025;
  assign n22028 = ~n22026 & ~n22027;
  assign n22029 = pi113  & n6396;
  assign n22030 = pi111  & n6735;
  assign n22031 = pi112  & n6391;
  assign n22032 = ~n22030 & ~n22031;
  assign n22033 = ~n22029 & n22032;
  assign n22034 = n6399 & n8387;
  assign n22035 = n22033 & ~n22034;
  assign n22036 = pi44  & ~n22035;
  assign n22037 = pi44  & ~n22036;
  assign n22038 = ~n22035 & ~n22036;
  assign n22039 = ~n22037 & ~n22038;
  assign n22040 = n22028 & ~n22039;
  assign n22041 = ~n22028 & n22039;
  assign n22042 = ~n22040 & ~n22041;
  assign n22043 = n21912 & ~n22042;
  assign n22044 = ~n21912 & n22042;
  assign n22045 = ~n22043 & ~n22044;
  assign n22046 = pi116  & n5636;
  assign n22047 = pi114  & n5909;
  assign n22048 = pi115  & n5631;
  assign n22049 = ~n22047 & ~n22048;
  assign n22050 = ~n22046 & n22049;
  assign n22051 = n5639 & n9042;
  assign n22052 = n22050 & ~n22051;
  assign n22053 = pi41  & ~n22052;
  assign n22054 = pi41  & ~n22053;
  assign n22055 = ~n22052 & ~n22053;
  assign n22056 = ~n22054 & ~n22055;
  assign n22057 = n22045 & ~n22056;
  assign n22058 = ~n22045 & n22056;
  assign n22059 = ~n22057 & ~n22058;
  assign n22060 = ~n21807 & n22059;
  assign n22061 = n21807 & ~n22059;
  assign n22062 = ~n22060 & ~n22061;
  assign n22063 = ~n21911 & n22062;
  assign n22064 = n21911 & ~n22062;
  assign n22065 = ~n22063 & ~n22064;
  assign n22066 = ~n21900 & n22065;
  assign n22067 = n21900 & ~n22065;
  assign n22068 = ~n22066 & ~n22067;
  assign n22069 = pi122  & n4182;
  assign n22070 = pi120  & n4416;
  assign n22071 = pi121  & n4177;
  assign n22072 = ~n22070 & ~n22071;
  assign n22073 = ~n22069 & n22072;
  assign n22074 = n4185 & n11463;
  assign n22075 = n22073 & ~n22074;
  assign n22076 = pi35  & ~n22075;
  assign n22077 = pi35  & ~n22076;
  assign n22078 = ~n22075 & ~n22076;
  assign n22079 = ~n22077 & ~n22078;
  assign n22080 = n22068 & ~n22079;
  assign n22081 = n22068 & ~n22080;
  assign n22082 = ~n22079 & ~n22080;
  assign n22083 = ~n22081 & ~n22082;
  assign n22084 = n21899 & ~n22083;
  assign n22085 = ~n21899 & n22083;
  assign n22086 = n21884 & ~n22085;
  assign n22087 = ~n22084 & n22086;
  assign n22088 = n21884 & ~n22087;
  assign n22089 = ~n22085 & ~n22087;
  assign n22090 = ~n22084 & n22089;
  assign n22091 = ~n22088 & ~n22090;
  assign n22092 = ~n21647 & ~n21862;
  assign n22093 = n22091 & n22092;
  assign n22094 = ~n22091 & ~n22092;
  assign n22095 = ~n22093 & ~n22094;
  assign n22096 = ~n21866 & ~n21869;
  assign n22097 = n22095 & ~n22096;
  assign n22098 = ~n22095 & n22096;
  assign po91  = ~n22097 & ~n22098;
  assign n22100 = ~n22094 & ~n22097;
  assign n22101 = ~n21882 & ~n22087;
  assign n22102 = pi126  & n3550;
  assign n22103 = pi124  & n3735;
  assign n22104 = pi125  & n3545;
  assign n22105 = ~n22103 & ~n22104;
  assign n22106 = ~n22102 & n22105;
  assign n22107 = n3553 & n12979;
  assign n22108 = n22106 & ~n22107;
  assign n22109 = pi32  & ~n22108;
  assign n22110 = pi32  & ~n22109;
  assign n22111 = ~n22108 & ~n22109;
  assign n22112 = ~n22110 & ~n22111;
  assign n22113 = ~n22066 & ~n22080;
  assign n22114 = n22112 & n22113;
  assign n22115 = ~n22112 & ~n22113;
  assign n22116 = ~n22114 & ~n22115;
  assign n22117 = ~n22060 & ~n22063;
  assign n22118 = pi120  & n4896;
  assign n22119 = pi118  & n5148;
  assign n22120 = pi119  & n4891;
  assign n22121 = ~n22119 & ~n22120;
  assign n22122 = ~n22118 & n22121;
  assign n22123 = n4899 & n10734;
  assign n22124 = n22122 & ~n22123;
  assign n22125 = pi38  & ~n22124;
  assign n22126 = pi38  & ~n22125;
  assign n22127 = ~n22124 & ~n22125;
  assign n22128 = ~n22126 & ~n22127;
  assign n22129 = ~n22044 & ~n22057;
  assign n22130 = pi117  & n5636;
  assign n22131 = pi115  & n5909;
  assign n22132 = pi116  & n5631;
  assign n22133 = ~n22131 & ~n22132;
  assign n22134 = ~n22130 & n22133;
  assign n22135 = n5639 & n9691;
  assign n22136 = n22134 & ~n22135;
  assign n22137 = pi41  & ~n22136;
  assign n22138 = pi41  & ~n22137;
  assign n22139 = ~n22136 & ~n22137;
  assign n22140 = ~n22138 & ~n22139;
  assign n22141 = ~n22027 & ~n22040;
  assign n22142 = ~n21992 & ~n22006;
  assign n22143 = pi108  & n8137;
  assign n22144 = pi106  & n8471;
  assign n22145 = pi107  & n8132;
  assign n22146 = ~n22144 & ~n22145;
  assign n22147 = ~n22143 & n22146;
  assign n22148 = n6639 & n8140;
  assign n22149 = n22147 & ~n22148;
  assign n22150 = pi50  & ~n22149;
  assign n22151 = pi50  & ~n22150;
  assign n22152 = ~n22149 & ~n22150;
  assign n22153 = ~n22151 & ~n22152;
  assign n22154 = ~n21986 & ~n21989;
  assign n22155 = ~n21961 & ~n21975;
  assign n22156 = pi99  & n11193;
  assign n22157 = pi97  & n11567;
  assign n22158 = pi98  & n11188;
  assign n22159 = ~n22157 & ~n22158;
  assign n22160 = ~n22156 & n22159;
  assign n22161 = n4584 & n11196;
  assign n22162 = n22160 & ~n22161;
  assign n22163 = pi59  & ~n22162;
  assign n22164 = pi59  & ~n22163;
  assign n22165 = ~n22162 & ~n22163;
  assign n22166 = ~n22164 & ~n22165;
  assign n22167 = ~n21944 & ~n21958;
  assign n22168 = pi92  & n13477;
  assign n22169 = pi93  & ~n13122;
  assign n22170 = ~n22168 & ~n22169;
  assign n22171 = n21941 & ~n22170;
  assign n22172 = ~n21941 & n22170;
  assign n22173 = ~n22167 & ~n22172;
  assign n22174 = ~n22171 & n22173;
  assign n22175 = ~n22167 & ~n22174;
  assign n22176 = ~n22172 & ~n22174;
  assign n22177 = ~n22171 & n22176;
  assign n22178 = ~n22175 & ~n22177;
  assign n22179 = pi96  & n12295;
  assign n22180 = pi94  & n12693;
  assign n22181 = pi95  & n12290;
  assign n22182 = ~n22180 & ~n22181;
  assign n22183 = ~n22179 & n22182;
  assign n22184 = n3921 & n12298;
  assign n22185 = n22183 & ~n22184;
  assign n22186 = pi62  & ~n22185;
  assign n22187 = pi62  & ~n22186;
  assign n22188 = ~n22185 & ~n22186;
  assign n22189 = ~n22187 & ~n22188;
  assign n22190 = ~n22178 & ~n22189;
  assign n22191 = n22178 & n22189;
  assign n22192 = ~n22190 & ~n22191;
  assign n22193 = ~n22166 & n22192;
  assign n22194 = n22166 & ~n22192;
  assign n22195 = ~n22193 & ~n22194;
  assign n22196 = ~n22155 & n22195;
  assign n22197 = n22155 & ~n22195;
  assign n22198 = ~n22196 & ~n22197;
  assign n22199 = pi102  & n10135;
  assign n22200 = pi100  & n10478;
  assign n22201 = pi101  & n10130;
  assign n22202 = ~n22200 & ~n22201;
  assign n22203 = ~n22199 & n22202;
  assign n22204 = n5296 & n10138;
  assign n22205 = n22203 & ~n22204;
  assign n22206 = pi56  & ~n22205;
  assign n22207 = pi56  & ~n22206;
  assign n22208 = ~n22205 & ~n22206;
  assign n22209 = ~n22207 & ~n22208;
  assign n22210 = n22198 & ~n22209;
  assign n22211 = ~n22198 & n22209;
  assign n22212 = ~n22210 & ~n22211;
  assign n22213 = ~n21981 & ~n21983;
  assign n22214 = n22212 & n22213;
  assign n22215 = n22212 & ~n22214;
  assign n22216 = n22213 & ~n22214;
  assign n22217 = ~n22215 & ~n22216;
  assign n22218 = pi105  & n9096;
  assign n22219 = pi103  & n9453;
  assign n22220 = pi104  & n9091;
  assign n22221 = ~n22219 & ~n22220;
  assign n22222 = ~n22218 & n22221;
  assign n22223 = n6065 & n9099;
  assign n22224 = n22222 & ~n22223;
  assign n22225 = pi53  & ~n22224;
  assign n22226 = pi53  & ~n22225;
  assign n22227 = ~n22224 & ~n22225;
  assign n22228 = ~n22226 & ~n22227;
  assign n22229 = ~n22217 & ~n22228;
  assign n22230 = n22217 & n22228;
  assign n22231 = ~n22229 & ~n22230;
  assign n22232 = ~n22154 & n22231;
  assign n22233 = n22154 & ~n22231;
  assign n22234 = ~n22232 & ~n22233;
  assign n22235 = ~n22153 & n22234;
  assign n22236 = n22153 & ~n22234;
  assign n22237 = ~n22235 & ~n22236;
  assign n22238 = ~n22142 & n22237;
  assign n22239 = n22142 & ~n22237;
  assign n22240 = ~n22238 & ~n22239;
  assign n22241 = pi111  & n7239;
  assign n22242 = pi109  & n7556;
  assign n22243 = pi110  & n7234;
  assign n22244 = ~n22242 & ~n22243;
  assign n22245 = ~n22241 & n22244;
  assign n22246 = n7242 & n7770;
  assign n22247 = n22245 & ~n22246;
  assign n22248 = pi47  & ~n22247;
  assign n22249 = pi47  & ~n22248;
  assign n22250 = ~n22247 & ~n22248;
  assign n22251 = ~n22249 & ~n22250;
  assign n22252 = n22240 & ~n22251;
  assign n22253 = n22240 & ~n22252;
  assign n22254 = ~n22251 & ~n22252;
  assign n22255 = ~n22253 & ~n22254;
  assign n22256 = ~n22010 & ~n22023;
  assign n22257 = n22255 & n22256;
  assign n22258 = ~n22255 & ~n22256;
  assign n22259 = ~n22257 & ~n22258;
  assign n22260 = pi114  & n6396;
  assign n22261 = pi112  & n6735;
  assign n22262 = pi113  & n6391;
  assign n22263 = ~n22261 & ~n22262;
  assign n22264 = ~n22260 & n22263;
  assign n22265 = n6399 & n8702;
  assign n22266 = n22264 & ~n22265;
  assign n22267 = pi44  & ~n22266;
  assign n22268 = pi44  & ~n22267;
  assign n22269 = ~n22266 & ~n22267;
  assign n22270 = ~n22268 & ~n22269;
  assign n22271 = ~n22259 & n22270;
  assign n22272 = n22259 & ~n22270;
  assign n22273 = ~n22271 & ~n22272;
  assign n22274 = ~n22141 & n22273;
  assign n22275 = n22141 & ~n22273;
  assign n22276 = ~n22274 & ~n22275;
  assign n22277 = ~n22140 & n22276;
  assign n22278 = n22140 & ~n22276;
  assign n22279 = ~n22277 & ~n22278;
  assign n22280 = ~n22129 & n22279;
  assign n22281 = n22129 & ~n22279;
  assign n22282 = ~n22280 & ~n22281;
  assign n22283 = ~n22128 & n22282;
  assign n22284 = n22128 & ~n22282;
  assign n22285 = ~n22283 & ~n22284;
  assign n22286 = ~n22117 & n22285;
  assign n22287 = n22117 & ~n22285;
  assign n22288 = ~n22286 & ~n22287;
  assign n22289 = pi123  & n4182;
  assign n22290 = pi121  & n4416;
  assign n22291 = pi122  & n4177;
  assign n22292 = ~n22290 & ~n22291;
  assign n22293 = ~n22289 & n22292;
  assign n22294 = n4185 & n11489;
  assign n22295 = n22293 & ~n22294;
  assign n22296 = pi35  & ~n22295;
  assign n22297 = pi35  & ~n22296;
  assign n22298 = ~n22295 & ~n22296;
  assign n22299 = ~n22297 & ~n22298;
  assign n22300 = n22288 & ~n22299;
  assign n22301 = n22288 & ~n22300;
  assign n22302 = ~n22299 & ~n22300;
  assign n22303 = ~n22301 & ~n22302;
  assign n22304 = ~n22116 & n22303;
  assign n22305 = n22116 & ~n22303;
  assign n22306 = ~n22304 & ~n22305;
  assign n22307 = ~n21898 & ~n22084;
  assign n22308 = pi127  & n3182;
  assign n22309 = n2979 & n13387;
  assign n22310 = ~n22308 & ~n22309;
  assign n22311 = pi29  & ~n22310;
  assign n22312 = pi29  & ~n22311;
  assign n22313 = ~n22310 & ~n22311;
  assign n22314 = ~n22312 & ~n22313;
  assign n22315 = ~n22307 & ~n22314;
  assign n22316 = n22307 & n22314;
  assign n22317 = ~n22315 & ~n22316;
  assign n22318 = n22306 & n22317;
  assign n22319 = ~n22306 & ~n22317;
  assign n22320 = ~n22318 & ~n22319;
  assign n22321 = ~n22101 & n22320;
  assign n22322 = n22101 & ~n22320;
  assign n22323 = ~n22321 & ~n22322;
  assign n22324 = ~n22100 & n22323;
  assign n22325 = n22100 & ~n22323;
  assign po92  = ~n22324 & ~n22325;
  assign n22327 = ~n22321 & ~n22324;
  assign n22328 = ~n22315 & ~n22318;
  assign n22329 = ~n22280 & ~n22283;
  assign n22330 = ~n22274 & ~n22277;
  assign n22331 = ~n22258 & ~n22272;
  assign n22332 = ~n22238 & ~n22252;
  assign n22333 = ~n22232 & ~n22235;
  assign n22334 = pi109  & n8137;
  assign n22335 = pi107  & n8471;
  assign n22336 = pi108  & n8132;
  assign n22337 = ~n22335 & ~n22336;
  assign n22338 = ~n22334 & n22337;
  assign n22339 = n7170 & n8140;
  assign n22340 = n22338 & ~n22339;
  assign n22341 = pi50  & ~n22340;
  assign n22342 = pi50  & ~n22341;
  assign n22343 = ~n22340 & ~n22341;
  assign n22344 = ~n22342 & ~n22343;
  assign n22345 = ~n22214 & ~n22229;
  assign n22346 = ~n22196 & ~n22210;
  assign n22347 = ~n22190 & ~n22193;
  assign n22348 = pi100  & n11193;
  assign n22349 = pi98  & n11567;
  assign n22350 = pi99  & n11188;
  assign n22351 = ~n22349 & ~n22350;
  assign n22352 = ~n22348 & n22351;
  assign n22353 = n4808 & n11196;
  assign n22354 = n22352 & ~n22353;
  assign n22355 = pi59  & ~n22354;
  assign n22356 = pi59  & ~n22355;
  assign n22357 = ~n22354 & ~n22355;
  assign n22358 = ~n22356 & ~n22357;
  assign n22359 = pi97  & n12295;
  assign n22360 = pi95  & n12693;
  assign n22361 = pi96  & n12290;
  assign n22362 = ~n22360 & ~n22361;
  assign n22363 = ~n22359 & n22362;
  assign n22364 = n3946 & n12298;
  assign n22365 = n22363 & ~n22364;
  assign n22366 = pi62  & ~n22365;
  assign n22367 = pi62  & ~n22366;
  assign n22368 = ~n22365 & ~n22366;
  assign n22369 = ~n22367 & ~n22368;
  assign n22370 = pi93  & n13477;
  assign n22371 = pi94  & ~n13122;
  assign n22372 = ~n22370 & ~n22371;
  assign n22373 = ~pi29  & ~n22372;
  assign n22374 = pi29  & n22372;
  assign n22375 = ~n22373 & ~n22374;
  assign n22376 = ~n22170 & n22375;
  assign n22377 = n22170 & ~n22375;
  assign n22378 = ~n22376 & ~n22377;
  assign n22379 = ~n22176 & n22378;
  assign n22380 = n22176 & ~n22378;
  assign n22381 = ~n22379 & ~n22380;
  assign n22382 = ~n22369 & n22381;
  assign n22383 = n22369 & ~n22381;
  assign n22384 = ~n22382 & ~n22383;
  assign n22385 = ~n22358 & n22384;
  assign n22386 = n22358 & ~n22384;
  assign n22387 = ~n22385 & ~n22386;
  assign n22388 = ~n22347 & n22387;
  assign n22389 = n22347 & ~n22387;
  assign n22390 = ~n22388 & ~n22389;
  assign n22391 = pi103  & n10135;
  assign n22392 = pi101  & n10478;
  assign n22393 = pi102  & n10130;
  assign n22394 = ~n22392 & ~n22393;
  assign n22395 = ~n22391 & n22394;
  assign n22396 = n5540 & n10138;
  assign n22397 = n22395 & ~n22396;
  assign n22398 = pi56  & ~n22397;
  assign n22399 = pi56  & ~n22398;
  assign n22400 = ~n22397 & ~n22398;
  assign n22401 = ~n22399 & ~n22400;
  assign n22402 = n22390 & ~n22401;
  assign n22403 = ~n22390 & n22401;
  assign n22404 = ~n22402 & ~n22403;
  assign n22405 = n22346 & ~n22404;
  assign n22406 = ~n22346 & n22404;
  assign n22407 = ~n22405 & ~n22406;
  assign n22408 = pi106  & n9096;
  assign n22409 = pi104  & n9453;
  assign n22410 = pi105  & n9091;
  assign n22411 = ~n22409 & ~n22410;
  assign n22412 = ~n22408 & n22411;
  assign n22413 = n6090 & n9099;
  assign n22414 = n22412 & ~n22413;
  assign n22415 = pi53  & ~n22414;
  assign n22416 = pi53  & ~n22415;
  assign n22417 = ~n22414 & ~n22415;
  assign n22418 = ~n22416 & ~n22417;
  assign n22419 = n22407 & ~n22418;
  assign n22420 = ~n22407 & n22418;
  assign n22421 = ~n22419 & ~n22420;
  assign n22422 = ~n22345 & n22421;
  assign n22423 = n22345 & ~n22421;
  assign n22424 = ~n22422 & ~n22423;
  assign n22425 = ~n22344 & n22424;
  assign n22426 = n22344 & ~n22424;
  assign n22427 = ~n22425 & ~n22426;
  assign n22428 = n22333 & ~n22427;
  assign n22429 = ~n22333 & n22427;
  assign n22430 = ~n22428 & ~n22429;
  assign n22431 = pi112  & n7239;
  assign n22432 = pi110  & n7556;
  assign n22433 = pi111  & n7234;
  assign n22434 = ~n22432 & ~n22433;
  assign n22435 = ~n22431 & n22434;
  assign n22436 = n7242 & n7795;
  assign n22437 = n22435 & ~n22436;
  assign n22438 = pi47  & ~n22437;
  assign n22439 = pi47  & ~n22438;
  assign n22440 = ~n22437 & ~n22438;
  assign n22441 = ~n22439 & ~n22440;
  assign n22442 = n22430 & ~n22441;
  assign n22443 = ~n22430 & n22441;
  assign n22444 = ~n22442 & ~n22443;
  assign n22445 = n22332 & ~n22444;
  assign n22446 = ~n22332 & n22444;
  assign n22447 = ~n22445 & ~n22446;
  assign n22448 = pi115  & n6396;
  assign n22449 = pi113  & n6735;
  assign n22450 = pi114  & n6391;
  assign n22451 = ~n22449 & ~n22450;
  assign n22452 = ~n22448 & n22451;
  assign n22453 = n6399 & n8727;
  assign n22454 = n22452 & ~n22453;
  assign n22455 = pi44  & ~n22454;
  assign n22456 = pi44  & ~n22455;
  assign n22457 = ~n22454 & ~n22455;
  assign n22458 = ~n22456 & ~n22457;
  assign n22459 = n22447 & ~n22458;
  assign n22460 = ~n22447 & n22458;
  assign n22461 = ~n22331 & ~n22460;
  assign n22462 = ~n22459 & n22461;
  assign n22463 = ~n22331 & ~n22462;
  assign n22464 = ~n22459 & ~n22462;
  assign n22465 = ~n22460 & n22464;
  assign n22466 = ~n22463 & ~n22465;
  assign n22467 = pi118  & n5636;
  assign n22468 = pi116  & n5909;
  assign n22469 = pi117  & n5631;
  assign n22470 = ~n22468 & ~n22469;
  assign n22471 = ~n22467 & n22470;
  assign n22472 = n5639 & n9716;
  assign n22473 = n22471 & ~n22472;
  assign n22474 = pi41  & ~n22473;
  assign n22475 = pi41  & ~n22474;
  assign n22476 = ~n22473 & ~n22474;
  assign n22477 = ~n22475 & ~n22476;
  assign n22478 = n22466 & n22477;
  assign n22479 = ~n22466 & ~n22477;
  assign n22480 = ~n22478 & ~n22479;
  assign n22481 = ~n22330 & n22480;
  assign n22482 = n22330 & ~n22480;
  assign n22483 = ~n22481 & ~n22482;
  assign n22484 = pi121  & n4896;
  assign n22485 = pi119  & n5148;
  assign n22486 = pi120  & n4891;
  assign n22487 = ~n22485 & ~n22486;
  assign n22488 = ~n22484 & n22487;
  assign n22489 = n4899 & n11086;
  assign n22490 = n22488 & ~n22489;
  assign n22491 = pi38  & ~n22490;
  assign n22492 = pi38  & ~n22491;
  assign n22493 = ~n22490 & ~n22491;
  assign n22494 = ~n22492 & ~n22493;
  assign n22495 = n22483 & ~n22494;
  assign n22496 = ~n22483 & n22494;
  assign n22497 = ~n22495 & ~n22496;
  assign n22498 = n22329 & ~n22497;
  assign n22499 = ~n22329 & n22497;
  assign n22500 = ~n22498 & ~n22499;
  assign n22501 = pi124  & n4182;
  assign n22502 = pi122  & n4416;
  assign n22503 = pi123  & n4177;
  assign n22504 = ~n22502 & ~n22503;
  assign n22505 = ~n22501 & n22504;
  assign n22506 = n4185 & n11858;
  assign n22507 = n22505 & ~n22506;
  assign n22508 = pi35  & ~n22507;
  assign n22509 = pi35  & ~n22508;
  assign n22510 = ~n22507 & ~n22508;
  assign n22511 = ~n22509 & ~n22510;
  assign n22512 = n22500 & ~n22511;
  assign n22513 = n22500 & ~n22512;
  assign n22514 = ~n22511 & ~n22512;
  assign n22515 = ~n22513 & ~n22514;
  assign n22516 = ~n22286 & ~n22300;
  assign n22517 = n22515 & n22516;
  assign n22518 = ~n22515 & ~n22516;
  assign n22519 = ~n22517 & ~n22518;
  assign n22520 = ~n22115 & ~n22305;
  assign n22521 = pi127  & n3550;
  assign n22522 = pi125  & n3735;
  assign n22523 = pi126  & n3545;
  assign n22524 = ~n22522 & ~n22523;
  assign n22525 = ~n22521 & n22524;
  assign n22526 = n3553 & n13365;
  assign n22527 = n22525 & ~n22526;
  assign n22528 = pi32  & ~n22527;
  assign n22529 = pi32  & ~n22528;
  assign n22530 = ~n22527 & ~n22528;
  assign n22531 = ~n22529 & ~n22530;
  assign n22532 = ~n22520 & ~n22531;
  assign n22533 = ~n22520 & ~n22532;
  assign n22534 = ~n22531 & ~n22532;
  assign n22535 = ~n22533 & ~n22534;
  assign n22536 = ~n22519 & n22535;
  assign n22537 = n22519 & ~n22535;
  assign n22538 = ~n22536 & ~n22537;
  assign n22539 = ~n22328 & n22538;
  assign n22540 = n22328 & ~n22538;
  assign n22541 = ~n22539 & ~n22540;
  assign n22542 = ~n22327 & n22541;
  assign n22543 = n22327 & ~n22541;
  assign po93  = ~n22542 & ~n22543;
  assign n22545 = ~n22539 & ~n22542;
  assign n22546 = ~n22512 & ~n22518;
  assign n22547 = pi126  & n3735;
  assign n22548 = pi127  & n3545;
  assign n22549 = ~n22547 & ~n22548;
  assign n22550 = ~n3553 & n22549;
  assign n22551 = ~n13389 & n22549;
  assign n22552 = ~n22550 & ~n22551;
  assign n22553 = pi32  & ~n22552;
  assign n22554 = ~pi32  & n22552;
  assign n22555 = ~n22553 & ~n22554;
  assign n22556 = ~n22546 & ~n22555;
  assign n22557 = n22546 & n22555;
  assign n22558 = ~n22556 & ~n22557;
  assign n22559 = ~n22479 & ~n22481;
  assign n22560 = pi119  & n5636;
  assign n22561 = pi117  & n5909;
  assign n22562 = pi118  & n5631;
  assign n22563 = ~n22561 & ~n22562;
  assign n22564 = ~n22560 & n22563;
  assign n22565 = n5639 & n10048;
  assign n22566 = n22564 & ~n22565;
  assign n22567 = pi41  & ~n22566;
  assign n22568 = pi41  & ~n22567;
  assign n22569 = ~n22566 & ~n22567;
  assign n22570 = ~n22568 & ~n22569;
  assign n22571 = ~n22442 & ~n22446;
  assign n22572 = ~n22425 & ~n22429;
  assign n22573 = ~n22419 & ~n22422;
  assign n22574 = ~n22402 & ~n22406;
  assign n22575 = pi104  & n10135;
  assign n22576 = pi102  & n10478;
  assign n22577 = pi103  & n10130;
  assign n22578 = ~n22576 & ~n22577;
  assign n22579 = ~n22575 & n22578;
  assign n22580 = n5565 & n10138;
  assign n22581 = n22579 & ~n22580;
  assign n22582 = pi56  & ~n22581;
  assign n22583 = pi56  & ~n22582;
  assign n22584 = ~n22581 & ~n22582;
  assign n22585 = ~n22583 & ~n22584;
  assign n22586 = ~n22385 & ~n22388;
  assign n22587 = pi101  & n11193;
  assign n22588 = pi99  & n11567;
  assign n22589 = pi100  & n11188;
  assign n22590 = ~n22588 & ~n22589;
  assign n22591 = ~n22587 & n22590;
  assign n22592 = n5056 & n11196;
  assign n22593 = n22591 & ~n22592;
  assign n22594 = pi59  & ~n22593;
  assign n22595 = pi59  & ~n22594;
  assign n22596 = ~n22593 & ~n22594;
  assign n22597 = ~n22595 & ~n22596;
  assign n22598 = ~n22379 & ~n22382;
  assign n22599 = pi94  & n13477;
  assign n22600 = pi95  & ~n13122;
  assign n22601 = ~n22599 & ~n22600;
  assign n22602 = ~n22373 & ~n22376;
  assign n22603 = ~n22601 & n22602;
  assign n22604 = n22601 & ~n22602;
  assign n22605 = ~n22603 & ~n22604;
  assign n22606 = pi98  & n12295;
  assign n22607 = pi96  & n12693;
  assign n22608 = pi97  & n12290;
  assign n22609 = ~n22607 & ~n22608;
  assign n22610 = ~n22606 & n22609;
  assign n22611 = n4360 & n12298;
  assign n22612 = n22610 & ~n22611;
  assign n22613 = pi62  & ~n22612;
  assign n22614 = pi62  & ~n22613;
  assign n22615 = ~n22612 & ~n22613;
  assign n22616 = ~n22614 & ~n22615;
  assign n22617 = ~n22605 & n22616;
  assign n22618 = n22605 & ~n22616;
  assign n22619 = ~n22617 & ~n22618;
  assign n22620 = ~n22598 & n22619;
  assign n22621 = n22598 & ~n22619;
  assign n22622 = ~n22620 & ~n22621;
  assign n22623 = ~n22597 & n22622;
  assign n22624 = n22597 & ~n22622;
  assign n22625 = ~n22623 & ~n22624;
  assign n22626 = ~n22586 & n22625;
  assign n22627 = n22586 & ~n22625;
  assign n22628 = ~n22626 & ~n22627;
  assign n22629 = ~n22585 & n22628;
  assign n22630 = n22585 & ~n22628;
  assign n22631 = ~n22629 & ~n22630;
  assign n22632 = ~n22574 & n22631;
  assign n22633 = n22574 & ~n22631;
  assign n22634 = ~n22632 & ~n22633;
  assign n22635 = pi107  & n9096;
  assign n22636 = pi105  & n9453;
  assign n22637 = pi106  & n9091;
  assign n22638 = ~n22636 & ~n22637;
  assign n22639 = ~n22635 & n22638;
  assign n22640 = n6614 & n9099;
  assign n22641 = n22639 & ~n22640;
  assign n22642 = pi53  & ~n22641;
  assign n22643 = pi53  & ~n22642;
  assign n22644 = ~n22641 & ~n22642;
  assign n22645 = ~n22643 & ~n22644;
  assign n22646 = n22634 & ~n22645;
  assign n22647 = ~n22634 & n22645;
  assign n22648 = ~n22646 & ~n22647;
  assign n22649 = n22573 & ~n22648;
  assign n22650 = ~n22573 & n22648;
  assign n22651 = ~n22649 & ~n22650;
  assign n22652 = pi110  & n8137;
  assign n22653 = pi108  & n8471;
  assign n22654 = pi109  & n8132;
  assign n22655 = ~n22653 & ~n22654;
  assign n22656 = ~n22652 & n22655;
  assign n22657 = n7474 & n8140;
  assign n22658 = n22656 & ~n22657;
  assign n22659 = pi50  & ~n22658;
  assign n22660 = pi50  & ~n22659;
  assign n22661 = ~n22658 & ~n22659;
  assign n22662 = ~n22660 & ~n22661;
  assign n22663 = n22651 & ~n22662;
  assign n22664 = ~n22651 & n22662;
  assign n22665 = ~n22663 & ~n22664;
  assign n22666 = n22572 & ~n22665;
  assign n22667 = ~n22572 & n22665;
  assign n22668 = ~n22666 & ~n22667;
  assign n22669 = pi113  & n7239;
  assign n22670 = pi111  & n7556;
  assign n22671 = pi112  & n7234;
  assign n22672 = ~n22670 & ~n22671;
  assign n22673 = ~n22669 & n22672;
  assign n22674 = n7242 & n8387;
  assign n22675 = n22673 & ~n22674;
  assign n22676 = pi47  & ~n22675;
  assign n22677 = pi47  & ~n22676;
  assign n22678 = ~n22675 & ~n22676;
  assign n22679 = ~n22677 & ~n22678;
  assign n22680 = n22668 & ~n22679;
  assign n22681 = ~n22668 & n22679;
  assign n22682 = ~n22680 & ~n22681;
  assign n22683 = n22571 & ~n22682;
  assign n22684 = ~n22571 & n22682;
  assign n22685 = ~n22683 & ~n22684;
  assign n22686 = pi116  & n6396;
  assign n22687 = pi114  & n6735;
  assign n22688 = pi115  & n6391;
  assign n22689 = ~n22687 & ~n22688;
  assign n22690 = ~n22686 & n22689;
  assign n22691 = n6399 & n9042;
  assign n22692 = n22690 & ~n22691;
  assign n22693 = pi44  & ~n22692;
  assign n22694 = pi44  & ~n22693;
  assign n22695 = ~n22692 & ~n22693;
  assign n22696 = ~n22694 & ~n22695;
  assign n22697 = n22685 & ~n22696;
  assign n22698 = ~n22685 & n22696;
  assign n22699 = ~n22697 & ~n22698;
  assign n22700 = ~n22464 & n22699;
  assign n22701 = n22464 & ~n22699;
  assign n22702 = ~n22700 & ~n22701;
  assign n22703 = ~n22570 & n22702;
  assign n22704 = n22570 & ~n22702;
  assign n22705 = ~n22703 & ~n22704;
  assign n22706 = ~n22559 & n22705;
  assign n22707 = n22559 & ~n22705;
  assign n22708 = ~n22706 & ~n22707;
  assign n22709 = pi122  & n4896;
  assign n22710 = pi120  & n5148;
  assign n22711 = pi121  & n4891;
  assign n22712 = ~n22710 & ~n22711;
  assign n22713 = ~n22709 & n22712;
  assign n22714 = n4899 & n11463;
  assign n22715 = n22713 & ~n22714;
  assign n22716 = pi38  & ~n22715;
  assign n22717 = pi38  & ~n22716;
  assign n22718 = ~n22715 & ~n22716;
  assign n22719 = ~n22717 & ~n22718;
  assign n22720 = n22708 & ~n22719;
  assign n22721 = n22708 & ~n22720;
  assign n22722 = ~n22719 & ~n22720;
  assign n22723 = ~n22721 & ~n22722;
  assign n22724 = ~n22495 & ~n22499;
  assign n22725 = n22723 & n22724;
  assign n22726 = ~n22723 & ~n22724;
  assign n22727 = ~n22725 & ~n22726;
  assign n22728 = pi125  & n4182;
  assign n22729 = pi123  & n4416;
  assign n22730 = pi124  & n4177;
  assign n22731 = ~n22729 & ~n22730;
  assign n22732 = ~n22728 & n22731;
  assign n22733 = n4185 & n12591;
  assign n22734 = n22732 & ~n22733;
  assign n22735 = pi35  & ~n22734;
  assign n22736 = pi35  & ~n22735;
  assign n22737 = ~n22734 & ~n22735;
  assign n22738 = ~n22736 & ~n22737;
  assign n22739 = n22727 & ~n22738;
  assign n22740 = ~n22727 & n22738;
  assign n22741 = n22558 & ~n22740;
  assign n22742 = ~n22739 & n22741;
  assign n22743 = n22558 & ~n22742;
  assign n22744 = ~n22740 & ~n22742;
  assign n22745 = ~n22739 & n22744;
  assign n22746 = ~n22743 & ~n22745;
  assign n22747 = ~n22532 & ~n22537;
  assign n22748 = ~n22746 & ~n22747;
  assign n22749 = n22746 & n22747;
  assign n22750 = ~n22748 & ~n22749;
  assign n22751 = ~n22545 & n22750;
  assign n22752 = n22545 & ~n22750;
  assign po94  = ~n22751 & ~n22752;
  assign n22754 = ~n22748 & ~n22751;
  assign n22755 = ~n22556 & ~n22742;
  assign n22756 = ~n22726 & ~n22739;
  assign n22757 = pi127  & n3735;
  assign n22758 = n3553 & n13387;
  assign n22759 = ~n22757 & ~n22758;
  assign n22760 = pi32  & ~n22759;
  assign n22761 = pi32  & ~n22760;
  assign n22762 = ~n22759 & ~n22760;
  assign n22763 = ~n22761 & ~n22762;
  assign n22764 = ~n22756 & ~n22763;
  assign n22765 = n22756 & n22763;
  assign n22766 = ~n22764 & ~n22765;
  assign n22767 = ~n22700 & ~n22703;
  assign n22768 = pi120  & n5636;
  assign n22769 = pi118  & n5909;
  assign n22770 = pi119  & n5631;
  assign n22771 = ~n22769 & ~n22770;
  assign n22772 = ~n22768 & n22771;
  assign n22773 = n5639 & n10734;
  assign n22774 = n22772 & ~n22773;
  assign n22775 = pi41  & ~n22774;
  assign n22776 = pi41  & ~n22775;
  assign n22777 = ~n22774 & ~n22775;
  assign n22778 = ~n22776 & ~n22777;
  assign n22779 = ~n22684 & ~n22697;
  assign n22780 = pi117  & n6396;
  assign n22781 = pi115  & n6735;
  assign n22782 = pi116  & n6391;
  assign n22783 = ~n22781 & ~n22782;
  assign n22784 = ~n22780 & n22783;
  assign n22785 = n6399 & n9691;
  assign n22786 = n22784 & ~n22785;
  assign n22787 = pi44  & ~n22786;
  assign n22788 = pi44  & ~n22787;
  assign n22789 = ~n22786 & ~n22787;
  assign n22790 = ~n22788 & ~n22789;
  assign n22791 = ~n22667 & ~n22680;
  assign n22792 = ~n22632 & ~n22646;
  assign n22793 = pi108  & n9096;
  assign n22794 = pi106  & n9453;
  assign n22795 = pi107  & n9091;
  assign n22796 = ~n22794 & ~n22795;
  assign n22797 = ~n22793 & n22796;
  assign n22798 = n6639 & n9099;
  assign n22799 = n22797 & ~n22798;
  assign n22800 = pi53  & ~n22799;
  assign n22801 = pi53  & ~n22800;
  assign n22802 = ~n22799 & ~n22800;
  assign n22803 = ~n22801 & ~n22802;
  assign n22804 = ~n22626 & ~n22629;
  assign n22805 = pi105  & n10135;
  assign n22806 = pi103  & n10478;
  assign n22807 = pi104  & n10130;
  assign n22808 = ~n22806 & ~n22807;
  assign n22809 = ~n22805 & n22808;
  assign n22810 = n6065 & n10138;
  assign n22811 = n22809 & ~n22810;
  assign n22812 = pi56  & ~n22811;
  assign n22813 = pi56  & ~n22812;
  assign n22814 = ~n22811 & ~n22812;
  assign n22815 = ~n22813 & ~n22814;
  assign n22816 = ~n22620 & ~n22623;
  assign n22817 = pi102  & n11193;
  assign n22818 = pi100  & n11567;
  assign n22819 = pi101  & n11188;
  assign n22820 = ~n22818 & ~n22819;
  assign n22821 = ~n22817 & n22820;
  assign n22822 = n5296 & n11196;
  assign n22823 = n22821 & ~n22822;
  assign n22824 = pi59  & ~n22823;
  assign n22825 = pi59  & ~n22824;
  assign n22826 = ~n22823 & ~n22824;
  assign n22827 = ~n22825 & ~n22826;
  assign n22828 = ~n22604 & ~n22618;
  assign n22829 = pi95  & n13477;
  assign n22830 = pi96  & ~n13122;
  assign n22831 = ~n22829 & ~n22830;
  assign n22832 = ~n22601 & n22831;
  assign n22833 = n22601 & ~n22831;
  assign n22834 = ~n22828 & ~n22833;
  assign n22835 = ~n22832 & n22834;
  assign n22836 = ~n22828 & ~n22835;
  assign n22837 = ~n22832 & ~n22835;
  assign n22838 = ~n22833 & n22837;
  assign n22839 = ~n22836 & ~n22838;
  assign n22840 = pi99  & n12295;
  assign n22841 = pi97  & n12693;
  assign n22842 = pi98  & n12290;
  assign n22843 = ~n22841 & ~n22842;
  assign n22844 = ~n22840 & n22843;
  assign n22845 = n4584 & n12298;
  assign n22846 = n22844 & ~n22845;
  assign n22847 = pi62  & ~n22846;
  assign n22848 = pi62  & ~n22847;
  assign n22849 = ~n22846 & ~n22847;
  assign n22850 = ~n22848 & ~n22849;
  assign n22851 = ~n22839 & ~n22850;
  assign n22852 = n22839 & n22850;
  assign n22853 = ~n22851 & ~n22852;
  assign n22854 = n22827 & n22853;
  assign n22855 = ~n22827 & ~n22853;
  assign n22856 = ~n22854 & ~n22855;
  assign n22857 = ~n22816 & ~n22856;
  assign n22858 = n22816 & n22856;
  assign n22859 = ~n22857 & ~n22858;
  assign n22860 = ~n22815 & n22859;
  assign n22861 = n22815 & ~n22859;
  assign n22862 = ~n22860 & ~n22861;
  assign n22863 = ~n22804 & n22862;
  assign n22864 = n22804 & ~n22862;
  assign n22865 = ~n22863 & ~n22864;
  assign n22866 = ~n22803 & n22865;
  assign n22867 = n22803 & ~n22865;
  assign n22868 = ~n22866 & ~n22867;
  assign n22869 = ~n22792 & n22868;
  assign n22870 = n22792 & ~n22868;
  assign n22871 = ~n22869 & ~n22870;
  assign n22872 = pi111  & n8137;
  assign n22873 = pi109  & n8471;
  assign n22874 = pi110  & n8132;
  assign n22875 = ~n22873 & ~n22874;
  assign n22876 = ~n22872 & n22875;
  assign n22877 = n7770 & n8140;
  assign n22878 = n22876 & ~n22877;
  assign n22879 = pi50  & ~n22878;
  assign n22880 = pi50  & ~n22879;
  assign n22881 = ~n22878 & ~n22879;
  assign n22882 = ~n22880 & ~n22881;
  assign n22883 = n22871 & ~n22882;
  assign n22884 = n22871 & ~n22883;
  assign n22885 = ~n22882 & ~n22883;
  assign n22886 = ~n22884 & ~n22885;
  assign n22887 = ~n22650 & ~n22663;
  assign n22888 = n22886 & n22887;
  assign n22889 = ~n22886 & ~n22887;
  assign n22890 = ~n22888 & ~n22889;
  assign n22891 = pi114  & n7239;
  assign n22892 = pi112  & n7556;
  assign n22893 = pi113  & n7234;
  assign n22894 = ~n22892 & ~n22893;
  assign n22895 = ~n22891 & n22894;
  assign n22896 = n7242 & n8702;
  assign n22897 = n22895 & ~n22896;
  assign n22898 = pi47  & ~n22897;
  assign n22899 = pi47  & ~n22898;
  assign n22900 = ~n22897 & ~n22898;
  assign n22901 = ~n22899 & ~n22900;
  assign n22902 = ~n22890 & n22901;
  assign n22903 = n22890 & ~n22901;
  assign n22904 = ~n22902 & ~n22903;
  assign n22905 = ~n22791 & n22904;
  assign n22906 = n22791 & ~n22904;
  assign n22907 = ~n22905 & ~n22906;
  assign n22908 = ~n22790 & n22907;
  assign n22909 = n22790 & ~n22907;
  assign n22910 = ~n22908 & ~n22909;
  assign n22911 = ~n22779 & n22910;
  assign n22912 = n22779 & ~n22910;
  assign n22913 = ~n22911 & ~n22912;
  assign n22914 = ~n22778 & n22913;
  assign n22915 = n22778 & ~n22913;
  assign n22916 = ~n22914 & ~n22915;
  assign n22917 = ~n22767 & n22916;
  assign n22918 = n22767 & ~n22916;
  assign n22919 = ~n22917 & ~n22918;
  assign n22920 = pi123  & n4896;
  assign n22921 = pi121  & n5148;
  assign n22922 = pi122  & n4891;
  assign n22923 = ~n22921 & ~n22922;
  assign n22924 = ~n22920 & n22923;
  assign n22925 = n4899 & n11489;
  assign n22926 = n22924 & ~n22925;
  assign n22927 = pi38  & ~n22926;
  assign n22928 = pi38  & ~n22927;
  assign n22929 = ~n22926 & ~n22927;
  assign n22930 = ~n22928 & ~n22929;
  assign n22931 = n22919 & ~n22930;
  assign n22932 = n22919 & ~n22931;
  assign n22933 = ~n22930 & ~n22931;
  assign n22934 = ~n22932 & ~n22933;
  assign n22935 = ~n22706 & ~n22720;
  assign n22936 = n22934 & n22935;
  assign n22937 = ~n22934 & ~n22935;
  assign n22938 = ~n22936 & ~n22937;
  assign n22939 = pi126  & n4182;
  assign n22940 = pi124  & n4416;
  assign n22941 = pi125  & n4177;
  assign n22942 = ~n22940 & ~n22941;
  assign n22943 = ~n22939 & n22942;
  assign n22944 = n4185 & n12979;
  assign n22945 = n22943 & ~n22944;
  assign n22946 = pi35  & ~n22945;
  assign n22947 = pi35  & ~n22946;
  assign n22948 = ~n22945 & ~n22946;
  assign n22949 = ~n22947 & ~n22948;
  assign n22950 = n22938 & ~n22949;
  assign n22951 = ~n22938 & n22949;
  assign n22952 = ~n22950 & ~n22951;
  assign n22953 = n22766 & ~n22952;
  assign n22954 = ~n22766 & n22952;
  assign n22955 = ~n22953 & ~n22954;
  assign n22956 = ~n22755 & ~n22955;
  assign n22957 = ~n22755 & ~n22956;
  assign n22958 = ~n22955 & ~n22956;
  assign n22959 = ~n22957 & ~n22958;
  assign n22960 = ~n22754 & ~n22959;
  assign n22961 = n22754 & n22959;
  assign po95  = ~n22960 & ~n22961;
  assign n22963 = ~n22956 & ~n22960;
  assign n22964 = ~n22911 & ~n22914;
  assign n22965 = ~n22905 & ~n22908;
  assign n22966 = ~n22889 & ~n22903;
  assign n22967 = ~n22869 & ~n22883;
  assign n22968 = ~n22863 & ~n22866;
  assign n22969 = ~n22857 & ~n22860;
  assign n22970 = pi103  & n11193;
  assign n22971 = pi101  & n11567;
  assign n22972 = pi102  & n11188;
  assign n22973 = ~n22971 & ~n22972;
  assign n22974 = ~n22970 & n22973;
  assign n22975 = n5540 & n11196;
  assign n22976 = n22974 & ~n22975;
  assign n22977 = pi59  & ~n22976;
  assign n22978 = pi59  & ~n22977;
  assign n22979 = ~n22976 & ~n22977;
  assign n22980 = ~n22978 & ~n22979;
  assign n22981 = pi100  & n12295;
  assign n22982 = pi98  & n12693;
  assign n22983 = pi99  & n12290;
  assign n22984 = ~n22982 & ~n22983;
  assign n22985 = ~n22981 & n22984;
  assign n22986 = n4808 & n12298;
  assign n22987 = n22985 & ~n22986;
  assign n22988 = pi62  & ~n22987;
  assign n22989 = pi62  & ~n22988;
  assign n22990 = ~n22987 & ~n22988;
  assign n22991 = ~n22989 & ~n22990;
  assign n22992 = pi96  & n13477;
  assign n22993 = pi97  & ~n13122;
  assign n22994 = ~n22992 & ~n22993;
  assign n22995 = ~pi32  & ~n22994;
  assign n22996 = pi32  & n22994;
  assign n22997 = ~n22995 & ~n22996;
  assign n22998 = ~n22831 & n22997;
  assign n22999 = n22831 & ~n22997;
  assign n23000 = ~n22998 & ~n22999;
  assign n23001 = ~n22837 & n23000;
  assign n23002 = n22837 & ~n23000;
  assign n23003 = ~n23001 & ~n23002;
  assign n23004 = ~n22991 & n23003;
  assign n23005 = n22991 & ~n23003;
  assign n23006 = ~n23004 & ~n23005;
  assign n23007 = ~n22980 & n23006;
  assign n23008 = n22980 & ~n23006;
  assign n23009 = ~n23007 & ~n23008;
  assign n23010 = ~n22852 & ~n22854;
  assign n23011 = n23009 & n23010;
  assign n23012 = ~n23009 & ~n23010;
  assign n23013 = ~n23011 & ~n23012;
  assign n23014 = pi106  & n10135;
  assign n23015 = pi104  & n10478;
  assign n23016 = pi105  & n10130;
  assign n23017 = ~n23015 & ~n23016;
  assign n23018 = ~n23014 & n23017;
  assign n23019 = n6090 & n10138;
  assign n23020 = n23018 & ~n23019;
  assign n23021 = pi56  & ~n23020;
  assign n23022 = pi56  & ~n23021;
  assign n23023 = ~n23020 & ~n23021;
  assign n23024 = ~n23022 & ~n23023;
  assign n23025 = n23013 & ~n23024;
  assign n23026 = ~n23013 & n23024;
  assign n23027 = ~n23025 & ~n23026;
  assign n23028 = n22969 & ~n23027;
  assign n23029 = ~n22969 & n23027;
  assign n23030 = ~n23028 & ~n23029;
  assign n23031 = pi109  & n9096;
  assign n23032 = pi107  & n9453;
  assign n23033 = pi108  & n9091;
  assign n23034 = ~n23032 & ~n23033;
  assign n23035 = ~n23031 & n23034;
  assign n23036 = n7170 & n9099;
  assign n23037 = n23035 & ~n23036;
  assign n23038 = pi53  & ~n23037;
  assign n23039 = pi53  & ~n23038;
  assign n23040 = ~n23037 & ~n23038;
  assign n23041 = ~n23039 & ~n23040;
  assign n23042 = n23030 & ~n23041;
  assign n23043 = ~n23030 & n23041;
  assign n23044 = ~n23042 & ~n23043;
  assign n23045 = n22968 & ~n23044;
  assign n23046 = ~n22968 & n23044;
  assign n23047 = ~n23045 & ~n23046;
  assign n23048 = pi112  & n8137;
  assign n23049 = pi110  & n8471;
  assign n23050 = pi111  & n8132;
  assign n23051 = ~n23049 & ~n23050;
  assign n23052 = ~n23048 & n23051;
  assign n23053 = n7795 & n8140;
  assign n23054 = n23052 & ~n23053;
  assign n23055 = pi50  & ~n23054;
  assign n23056 = pi50  & ~n23055;
  assign n23057 = ~n23054 & ~n23055;
  assign n23058 = ~n23056 & ~n23057;
  assign n23059 = n23047 & ~n23058;
  assign n23060 = ~n23047 & n23058;
  assign n23061 = ~n23059 & ~n23060;
  assign n23062 = n22967 & ~n23061;
  assign n23063 = ~n22967 & n23061;
  assign n23064 = ~n23062 & ~n23063;
  assign n23065 = pi115  & n7239;
  assign n23066 = pi113  & n7556;
  assign n23067 = pi114  & n7234;
  assign n23068 = ~n23066 & ~n23067;
  assign n23069 = ~n23065 & n23068;
  assign n23070 = n7242 & n8727;
  assign n23071 = n23069 & ~n23070;
  assign n23072 = pi47  & ~n23071;
  assign n23073 = pi47  & ~n23072;
  assign n23074 = ~n23071 & ~n23072;
  assign n23075 = ~n23073 & ~n23074;
  assign n23076 = n23064 & ~n23075;
  assign n23077 = ~n23064 & n23075;
  assign n23078 = ~n22966 & ~n23077;
  assign n23079 = ~n23076 & n23078;
  assign n23080 = ~n22966 & ~n23079;
  assign n23081 = ~n23076 & ~n23079;
  assign n23082 = ~n23077 & n23081;
  assign n23083 = ~n23080 & ~n23082;
  assign n23084 = pi118  & n6396;
  assign n23085 = pi116  & n6735;
  assign n23086 = pi117  & n6391;
  assign n23087 = ~n23085 & ~n23086;
  assign n23088 = ~n23084 & n23087;
  assign n23089 = n6399 & n9716;
  assign n23090 = n23088 & ~n23089;
  assign n23091 = pi44  & ~n23090;
  assign n23092 = pi44  & ~n23091;
  assign n23093 = ~n23090 & ~n23091;
  assign n23094 = ~n23092 & ~n23093;
  assign n23095 = n23083 & n23094;
  assign n23096 = ~n23083 & ~n23094;
  assign n23097 = ~n23095 & ~n23096;
  assign n23098 = ~n22965 & n23097;
  assign n23099 = n22965 & ~n23097;
  assign n23100 = ~n23098 & ~n23099;
  assign n23101 = pi121  & n5636;
  assign n23102 = pi119  & n5909;
  assign n23103 = pi120  & n5631;
  assign n23104 = ~n23102 & ~n23103;
  assign n23105 = ~n23101 & n23104;
  assign n23106 = n5639 & n11086;
  assign n23107 = n23105 & ~n23106;
  assign n23108 = pi41  & ~n23107;
  assign n23109 = pi41  & ~n23108;
  assign n23110 = ~n23107 & ~n23108;
  assign n23111 = ~n23109 & ~n23110;
  assign n23112 = n23100 & ~n23111;
  assign n23113 = ~n23100 & n23111;
  assign n23114 = ~n23112 & ~n23113;
  assign n23115 = n22964 & ~n23114;
  assign n23116 = ~n22964 & n23114;
  assign n23117 = ~n23115 & ~n23116;
  assign n23118 = pi124  & n4896;
  assign n23119 = pi122  & n5148;
  assign n23120 = pi123  & n4891;
  assign n23121 = ~n23119 & ~n23120;
  assign n23122 = ~n23118 & n23121;
  assign n23123 = n4899 & n11858;
  assign n23124 = n23122 & ~n23123;
  assign n23125 = pi38  & ~n23124;
  assign n23126 = pi38  & ~n23125;
  assign n23127 = ~n23124 & ~n23125;
  assign n23128 = ~n23126 & ~n23127;
  assign n23129 = n23117 & ~n23128;
  assign n23130 = n23117 & ~n23129;
  assign n23131 = ~n23128 & ~n23129;
  assign n23132 = ~n23130 & ~n23131;
  assign n23133 = ~n22917 & ~n22931;
  assign n23134 = n23132 & n23133;
  assign n23135 = ~n23132 & ~n23133;
  assign n23136 = ~n23134 & ~n23135;
  assign n23137 = ~n22937 & ~n22950;
  assign n23138 = pi127  & n4182;
  assign n23139 = pi125  & n4416;
  assign n23140 = pi126  & n4177;
  assign n23141 = ~n23139 & ~n23140;
  assign n23142 = ~n23138 & n23141;
  assign n23143 = n4185 & n13365;
  assign n23144 = n23142 & ~n23143;
  assign n23145 = pi35  & ~n23144;
  assign n23146 = pi35  & ~n23145;
  assign n23147 = ~n23144 & ~n23145;
  assign n23148 = ~n23146 & ~n23147;
  assign n23149 = ~n23137 & ~n23148;
  assign n23150 = ~n23137 & ~n23149;
  assign n23151 = ~n23148 & ~n23149;
  assign n23152 = ~n23150 & ~n23151;
  assign n23153 = ~n23136 & n23152;
  assign n23154 = n23136 & ~n23152;
  assign n23155 = ~n23153 & ~n23154;
  assign n23156 = ~n22765 & ~n22953;
  assign n23157 = n23155 & n23156;
  assign n23158 = ~n23155 & ~n23156;
  assign n23159 = ~n23157 & ~n23158;
  assign n23160 = ~n22963 & n23159;
  assign n23161 = n22963 & ~n23159;
  assign po96  = ~n23160 & ~n23161;
  assign n23163 = ~n23157 & ~n23160;
  assign n23164 = ~n23129 & ~n23135;
  assign n23165 = pi126  & n4416;
  assign n23166 = pi127  & n4177;
  assign n23167 = ~n23165 & ~n23166;
  assign n23168 = ~n4185 & n23167;
  assign n23169 = ~n13389 & n23167;
  assign n23170 = ~n23168 & ~n23169;
  assign n23171 = pi35  & ~n23170;
  assign n23172 = ~pi35  & n23170;
  assign n23173 = ~n23171 & ~n23172;
  assign n23174 = ~n23164 & ~n23173;
  assign n23175 = n23164 & n23173;
  assign n23176 = ~n23174 & ~n23175;
  assign n23177 = ~n23096 & ~n23098;
  assign n23178 = pi119  & n6396;
  assign n23179 = pi117  & n6735;
  assign n23180 = pi118  & n6391;
  assign n23181 = ~n23179 & ~n23180;
  assign n23182 = ~n23178 & n23181;
  assign n23183 = n6399 & n10048;
  assign n23184 = n23182 & ~n23183;
  assign n23185 = pi44  & ~n23184;
  assign n23186 = pi44  & ~n23185;
  assign n23187 = ~n23184 & ~n23185;
  assign n23188 = ~n23186 & ~n23187;
  assign n23189 = ~n23059 & ~n23063;
  assign n23190 = ~n23042 & ~n23046;
  assign n23191 = ~n23025 & ~n23029;
  assign n23192 = ~n23007 & ~n23011;
  assign n23193 = pi104  & n11193;
  assign n23194 = pi102  & n11567;
  assign n23195 = pi103  & n11188;
  assign n23196 = ~n23194 & ~n23195;
  assign n23197 = ~n23193 & n23196;
  assign n23198 = n5565 & n11196;
  assign n23199 = n23197 & ~n23198;
  assign n23200 = pi59  & ~n23199;
  assign n23201 = pi59  & ~n23200;
  assign n23202 = ~n23199 & ~n23200;
  assign n23203 = ~n23201 & ~n23202;
  assign n23204 = ~n23001 & ~n23004;
  assign n23205 = pi97  & n13477;
  assign n23206 = pi98  & ~n13122;
  assign n23207 = ~n23205 & ~n23206;
  assign n23208 = ~n22995 & ~n22998;
  assign n23209 = ~n23207 & n23208;
  assign n23210 = n23207 & ~n23208;
  assign n23211 = ~n23209 & ~n23210;
  assign n23212 = pi101  & n12295;
  assign n23213 = pi99  & n12693;
  assign n23214 = pi100  & n12290;
  assign n23215 = ~n23213 & ~n23214;
  assign n23216 = ~n23212 & n23215;
  assign n23217 = n5056 & n12298;
  assign n23218 = n23216 & ~n23217;
  assign n23219 = pi62  & ~n23218;
  assign n23220 = pi62  & ~n23219;
  assign n23221 = ~n23218 & ~n23219;
  assign n23222 = ~n23220 & ~n23221;
  assign n23223 = ~n23211 & n23222;
  assign n23224 = n23211 & ~n23222;
  assign n23225 = ~n23223 & ~n23224;
  assign n23226 = ~n23204 & n23225;
  assign n23227 = n23204 & ~n23225;
  assign n23228 = ~n23226 & ~n23227;
  assign n23229 = ~n23203 & n23228;
  assign n23230 = n23203 & ~n23228;
  assign n23231 = ~n23229 & ~n23230;
  assign n23232 = ~n23192 & n23231;
  assign n23233 = n23192 & ~n23231;
  assign n23234 = ~n23232 & ~n23233;
  assign n23235 = pi107  & n10135;
  assign n23236 = pi105  & n10478;
  assign n23237 = pi106  & n10130;
  assign n23238 = ~n23236 & ~n23237;
  assign n23239 = ~n23235 & n23238;
  assign n23240 = n6614 & n10138;
  assign n23241 = n23239 & ~n23240;
  assign n23242 = pi56  & ~n23241;
  assign n23243 = pi56  & ~n23242;
  assign n23244 = ~n23241 & ~n23242;
  assign n23245 = ~n23243 & ~n23244;
  assign n23246 = n23234 & ~n23245;
  assign n23247 = ~n23234 & n23245;
  assign n23248 = ~n23246 & ~n23247;
  assign n23249 = n23191 & ~n23248;
  assign n23250 = ~n23191 & n23248;
  assign n23251 = ~n23249 & ~n23250;
  assign n23252 = pi110  & n9096;
  assign n23253 = pi108  & n9453;
  assign n23254 = pi109  & n9091;
  assign n23255 = ~n23253 & ~n23254;
  assign n23256 = ~n23252 & n23255;
  assign n23257 = n7474 & n9099;
  assign n23258 = n23256 & ~n23257;
  assign n23259 = pi53  & ~n23258;
  assign n23260 = pi53  & ~n23259;
  assign n23261 = ~n23258 & ~n23259;
  assign n23262 = ~n23260 & ~n23261;
  assign n23263 = n23251 & ~n23262;
  assign n23264 = ~n23251 & n23262;
  assign n23265 = ~n23263 & ~n23264;
  assign n23266 = n23190 & ~n23265;
  assign n23267 = ~n23190 & n23265;
  assign n23268 = ~n23266 & ~n23267;
  assign n23269 = pi113  & n8137;
  assign n23270 = pi111  & n8471;
  assign n23271 = pi112  & n8132;
  assign n23272 = ~n23270 & ~n23271;
  assign n23273 = ~n23269 & n23272;
  assign n23274 = n8140 & n8387;
  assign n23275 = n23273 & ~n23274;
  assign n23276 = pi50  & ~n23275;
  assign n23277 = pi50  & ~n23276;
  assign n23278 = ~n23275 & ~n23276;
  assign n23279 = ~n23277 & ~n23278;
  assign n23280 = n23268 & ~n23279;
  assign n23281 = ~n23268 & n23279;
  assign n23282 = ~n23280 & ~n23281;
  assign n23283 = n23189 & ~n23282;
  assign n23284 = ~n23189 & n23282;
  assign n23285 = ~n23283 & ~n23284;
  assign n23286 = pi116  & n7239;
  assign n23287 = pi114  & n7556;
  assign n23288 = pi115  & n7234;
  assign n23289 = ~n23287 & ~n23288;
  assign n23290 = ~n23286 & n23289;
  assign n23291 = n7242 & n9042;
  assign n23292 = n23290 & ~n23291;
  assign n23293 = pi47  & ~n23292;
  assign n23294 = pi47  & ~n23293;
  assign n23295 = ~n23292 & ~n23293;
  assign n23296 = ~n23294 & ~n23295;
  assign n23297 = n23285 & ~n23296;
  assign n23298 = ~n23285 & n23296;
  assign n23299 = ~n23297 & ~n23298;
  assign n23300 = ~n23081 & n23299;
  assign n23301 = n23081 & ~n23299;
  assign n23302 = ~n23300 & ~n23301;
  assign n23303 = ~n23188 & n23302;
  assign n23304 = n23188 & ~n23302;
  assign n23305 = ~n23303 & ~n23304;
  assign n23306 = ~n23177 & n23305;
  assign n23307 = n23177 & ~n23305;
  assign n23308 = ~n23306 & ~n23307;
  assign n23309 = pi122  & n5636;
  assign n23310 = pi120  & n5909;
  assign n23311 = pi121  & n5631;
  assign n23312 = ~n23310 & ~n23311;
  assign n23313 = ~n23309 & n23312;
  assign n23314 = n5639 & n11463;
  assign n23315 = n23313 & ~n23314;
  assign n23316 = pi41  & ~n23315;
  assign n23317 = pi41  & ~n23316;
  assign n23318 = ~n23315 & ~n23316;
  assign n23319 = ~n23317 & ~n23318;
  assign n23320 = n23308 & ~n23319;
  assign n23321 = n23308 & ~n23320;
  assign n23322 = ~n23319 & ~n23320;
  assign n23323 = ~n23321 & ~n23322;
  assign n23324 = ~n23112 & ~n23116;
  assign n23325 = n23323 & n23324;
  assign n23326 = ~n23323 & ~n23324;
  assign n23327 = ~n23325 & ~n23326;
  assign n23328 = pi125  & n4896;
  assign n23329 = pi123  & n5148;
  assign n23330 = pi124  & n4891;
  assign n23331 = ~n23329 & ~n23330;
  assign n23332 = ~n23328 & n23331;
  assign n23333 = n4899 & n12591;
  assign n23334 = n23332 & ~n23333;
  assign n23335 = pi38  & ~n23334;
  assign n23336 = pi38  & ~n23335;
  assign n23337 = ~n23334 & ~n23335;
  assign n23338 = ~n23336 & ~n23337;
  assign n23339 = n23327 & ~n23338;
  assign n23340 = ~n23327 & n23338;
  assign n23341 = n23176 & ~n23340;
  assign n23342 = ~n23339 & n23341;
  assign n23343 = n23176 & ~n23342;
  assign n23344 = ~n23340 & ~n23342;
  assign n23345 = ~n23339 & n23344;
  assign n23346 = ~n23343 & ~n23345;
  assign n23347 = ~n23149 & ~n23154;
  assign n23348 = ~n23346 & ~n23347;
  assign n23349 = n23346 & n23347;
  assign n23350 = ~n23348 & ~n23349;
  assign n23351 = ~n23163 & n23350;
  assign n23352 = n23163 & ~n23350;
  assign po97  = ~n23351 & ~n23352;
  assign n23354 = ~n23348 & ~n23351;
  assign n23355 = ~n23174 & ~n23342;
  assign n23356 = ~n23326 & ~n23339;
  assign n23357 = pi127  & n4416;
  assign n23358 = n4185 & n13387;
  assign n23359 = ~n23357 & ~n23358;
  assign n23360 = pi35  & ~n23359;
  assign n23361 = pi35  & ~n23360;
  assign n23362 = ~n23359 & ~n23360;
  assign n23363 = ~n23361 & ~n23362;
  assign n23364 = ~n23356 & ~n23363;
  assign n23365 = n23356 & n23363;
  assign n23366 = ~n23364 & ~n23365;
  assign n23367 = ~n23300 & ~n23303;
  assign n23368 = pi120  & n6396;
  assign n23369 = pi118  & n6735;
  assign n23370 = pi119  & n6391;
  assign n23371 = ~n23369 & ~n23370;
  assign n23372 = ~n23368 & n23371;
  assign n23373 = n6399 & n10734;
  assign n23374 = n23372 & ~n23373;
  assign n23375 = pi44  & ~n23374;
  assign n23376 = pi44  & ~n23375;
  assign n23377 = ~n23374 & ~n23375;
  assign n23378 = ~n23376 & ~n23377;
  assign n23379 = ~n23284 & ~n23297;
  assign n23380 = pi117  & n7239;
  assign n23381 = pi115  & n7556;
  assign n23382 = pi116  & n7234;
  assign n23383 = ~n23381 & ~n23382;
  assign n23384 = ~n23380 & n23383;
  assign n23385 = n7242 & n9691;
  assign n23386 = n23384 & ~n23385;
  assign n23387 = pi47  & ~n23386;
  assign n23388 = pi47  & ~n23387;
  assign n23389 = ~n23386 & ~n23387;
  assign n23390 = ~n23388 & ~n23389;
  assign n23391 = ~n23267 & ~n23280;
  assign n23392 = ~n23250 & ~n23263;
  assign n23393 = ~n23232 & ~n23246;
  assign n23394 = pi108  & n10135;
  assign n23395 = pi106  & n10478;
  assign n23396 = pi107  & n10130;
  assign n23397 = ~n23395 & ~n23396;
  assign n23398 = ~n23394 & n23397;
  assign n23399 = n6639 & n10138;
  assign n23400 = n23398 & ~n23399;
  assign n23401 = pi56  & ~n23400;
  assign n23402 = pi56  & ~n23401;
  assign n23403 = ~n23400 & ~n23401;
  assign n23404 = ~n23402 & ~n23403;
  assign n23405 = ~n23226 & ~n23229;
  assign n23406 = pi105  & n11193;
  assign n23407 = pi103  & n11567;
  assign n23408 = pi104  & n11188;
  assign n23409 = ~n23407 & ~n23408;
  assign n23410 = ~n23406 & n23409;
  assign n23411 = n6065 & n11196;
  assign n23412 = n23410 & ~n23411;
  assign n23413 = pi59  & ~n23412;
  assign n23414 = pi59  & ~n23413;
  assign n23415 = ~n23412 & ~n23413;
  assign n23416 = ~n23414 & ~n23415;
  assign n23417 = ~n23210 & ~n23224;
  assign n23418 = pi98  & n13477;
  assign n23419 = pi99  & ~n13122;
  assign n23420 = ~n23418 & ~n23419;
  assign n23421 = ~n23207 & n23420;
  assign n23422 = n23207 & ~n23420;
  assign n23423 = ~n23417 & ~n23422;
  assign n23424 = ~n23421 & n23423;
  assign n23425 = ~n23417 & ~n23424;
  assign n23426 = ~n23421 & ~n23424;
  assign n23427 = ~n23422 & n23426;
  assign n23428 = ~n23425 & ~n23427;
  assign n23429 = pi102  & n12295;
  assign n23430 = pi100  & n12693;
  assign n23431 = pi101  & n12290;
  assign n23432 = ~n23430 & ~n23431;
  assign n23433 = ~n23429 & n23432;
  assign n23434 = n5296 & n12298;
  assign n23435 = n23433 & ~n23434;
  assign n23436 = pi62  & ~n23435;
  assign n23437 = pi62  & ~n23436;
  assign n23438 = ~n23435 & ~n23436;
  assign n23439 = ~n23437 & ~n23438;
  assign n23440 = ~n23428 & ~n23439;
  assign n23441 = n23428 & n23439;
  assign n23442 = ~n23440 & ~n23441;
  assign n23443 = n23416 & n23442;
  assign n23444 = ~n23416 & ~n23442;
  assign n23445 = ~n23443 & ~n23444;
  assign n23446 = ~n23405 & ~n23445;
  assign n23447 = n23405 & n23445;
  assign n23448 = ~n23446 & ~n23447;
  assign n23449 = ~n23404 & n23448;
  assign n23450 = n23404 & ~n23448;
  assign n23451 = ~n23449 & ~n23450;
  assign n23452 = ~n23393 & n23451;
  assign n23453 = n23393 & ~n23451;
  assign n23454 = ~n23452 & ~n23453;
  assign n23455 = pi111  & n9096;
  assign n23456 = pi109  & n9453;
  assign n23457 = pi110  & n9091;
  assign n23458 = ~n23456 & ~n23457;
  assign n23459 = ~n23455 & n23458;
  assign n23460 = n7770 & n9099;
  assign n23461 = n23459 & ~n23460;
  assign n23462 = pi53  & ~n23461;
  assign n23463 = pi53  & ~n23462;
  assign n23464 = ~n23461 & ~n23462;
  assign n23465 = ~n23463 & ~n23464;
  assign n23466 = n23454 & ~n23465;
  assign n23467 = ~n23454 & n23465;
  assign n23468 = ~n23466 & ~n23467;
  assign n23469 = n23392 & ~n23468;
  assign n23470 = ~n23392 & n23468;
  assign n23471 = ~n23469 & ~n23470;
  assign n23472 = pi114  & n8137;
  assign n23473 = pi112  & n8471;
  assign n23474 = pi113  & n8132;
  assign n23475 = ~n23473 & ~n23474;
  assign n23476 = ~n23472 & n23475;
  assign n23477 = n8140 & n8702;
  assign n23478 = n23476 & ~n23477;
  assign n23479 = pi50  & ~n23478;
  assign n23480 = pi50  & ~n23479;
  assign n23481 = ~n23478 & ~n23479;
  assign n23482 = ~n23480 & ~n23481;
  assign n23483 = ~n23471 & n23482;
  assign n23484 = n23471 & ~n23482;
  assign n23485 = ~n23483 & ~n23484;
  assign n23486 = ~n23391 & n23485;
  assign n23487 = n23391 & ~n23485;
  assign n23488 = ~n23486 & ~n23487;
  assign n23489 = ~n23390 & n23488;
  assign n23490 = n23390 & ~n23488;
  assign n23491 = ~n23489 & ~n23490;
  assign n23492 = ~n23379 & n23491;
  assign n23493 = n23379 & ~n23491;
  assign n23494 = ~n23492 & ~n23493;
  assign n23495 = ~n23378 & n23494;
  assign n23496 = n23378 & ~n23494;
  assign n23497 = ~n23495 & ~n23496;
  assign n23498 = ~n23367 & n23497;
  assign n23499 = n23367 & ~n23497;
  assign n23500 = ~n23498 & ~n23499;
  assign n23501 = pi123  & n5636;
  assign n23502 = pi121  & n5909;
  assign n23503 = pi122  & n5631;
  assign n23504 = ~n23502 & ~n23503;
  assign n23505 = ~n23501 & n23504;
  assign n23506 = n5639 & n11489;
  assign n23507 = n23505 & ~n23506;
  assign n23508 = pi41  & ~n23507;
  assign n23509 = pi41  & ~n23508;
  assign n23510 = ~n23507 & ~n23508;
  assign n23511 = ~n23509 & ~n23510;
  assign n23512 = n23500 & ~n23511;
  assign n23513 = n23500 & ~n23512;
  assign n23514 = ~n23511 & ~n23512;
  assign n23515 = ~n23513 & ~n23514;
  assign n23516 = ~n23306 & ~n23320;
  assign n23517 = n23515 & n23516;
  assign n23518 = ~n23515 & ~n23516;
  assign n23519 = ~n23517 & ~n23518;
  assign n23520 = pi126  & n4896;
  assign n23521 = pi124  & n5148;
  assign n23522 = pi125  & n4891;
  assign n23523 = ~n23521 & ~n23522;
  assign n23524 = ~n23520 & n23523;
  assign n23525 = n4899 & n12979;
  assign n23526 = n23524 & ~n23525;
  assign n23527 = pi38  & ~n23526;
  assign n23528 = pi38  & ~n23527;
  assign n23529 = ~n23526 & ~n23527;
  assign n23530 = ~n23528 & ~n23529;
  assign n23531 = n23519 & ~n23530;
  assign n23532 = ~n23519 & n23530;
  assign n23533 = ~n23531 & ~n23532;
  assign n23534 = n23366 & ~n23533;
  assign n23535 = ~n23366 & n23533;
  assign n23536 = ~n23534 & ~n23535;
  assign n23537 = ~n23355 & ~n23536;
  assign n23538 = n23355 & n23536;
  assign n23539 = ~n23537 & ~n23538;
  assign n23540 = ~n23354 & n23539;
  assign n23541 = n23354 & ~n23539;
  assign po98  = ~n23540 & ~n23541;
  assign n23543 = ~n23537 & ~n23540;
  assign n23544 = ~n23518 & ~n23531;
  assign n23545 = ~n23498 & ~n23512;
  assign n23546 = ~n23486 & ~n23489;
  assign n23547 = pi118  & n7239;
  assign n23548 = pi116  & n7556;
  assign n23549 = pi117  & n7234;
  assign n23550 = ~n23548 & ~n23549;
  assign n23551 = ~n23547 & n23550;
  assign n23552 = n7242 & n9716;
  assign n23553 = n23551 & ~n23552;
  assign n23554 = pi47  & ~n23553;
  assign n23555 = pi47  & ~n23554;
  assign n23556 = ~n23553 & ~n23554;
  assign n23557 = ~n23555 & ~n23556;
  assign n23558 = ~n23470 & ~n23484;
  assign n23559 = ~n23452 & ~n23466;
  assign n23560 = ~n23446 & ~n23449;
  assign n23561 = pi109  & n10135;
  assign n23562 = pi107  & n10478;
  assign n23563 = pi108  & n10130;
  assign n23564 = ~n23562 & ~n23563;
  assign n23565 = ~n23561 & n23564;
  assign n23566 = n7170 & n10138;
  assign n23567 = n23565 & ~n23566;
  assign n23568 = pi56  & ~n23567;
  assign n23569 = pi56  & ~n23568;
  assign n23570 = ~n23567 & ~n23568;
  assign n23571 = ~n23569 & ~n23570;
  assign n23572 = pi99  & n13477;
  assign n23573 = pi100  & ~n13122;
  assign n23574 = ~n23572 & ~n23573;
  assign n23575 = ~pi35  & ~n23420;
  assign n23576 = pi35  & n23420;
  assign n23577 = ~n23575 & ~n23576;
  assign n23578 = ~n23574 & n23577;
  assign n23579 = n23574 & ~n23577;
  assign n23580 = ~n23578 & ~n23579;
  assign n23581 = ~n23426 & n23580;
  assign n23582 = n23426 & ~n23580;
  assign n23583 = ~n23581 & ~n23582;
  assign n23584 = pi103  & n12295;
  assign n23585 = pi101  & n12693;
  assign n23586 = pi102  & n12290;
  assign n23587 = ~n23585 & ~n23586;
  assign n23588 = ~n23584 & n23587;
  assign n23589 = n5540 & n12298;
  assign n23590 = n23588 & ~n23589;
  assign n23591 = pi62  & ~n23590;
  assign n23592 = pi62  & ~n23591;
  assign n23593 = ~n23590 & ~n23591;
  assign n23594 = ~n23592 & ~n23593;
  assign n23595 = ~n23583 & n23594;
  assign n23596 = n23583 & ~n23594;
  assign n23597 = ~n23595 & ~n23596;
  assign n23598 = pi106  & n11193;
  assign n23599 = pi104  & n11567;
  assign n23600 = pi105  & n11188;
  assign n23601 = ~n23599 & ~n23600;
  assign n23602 = ~n23598 & n23601;
  assign n23603 = n6090 & n11196;
  assign n23604 = n23602 & ~n23603;
  assign n23605 = pi59  & ~n23604;
  assign n23606 = pi59  & ~n23605;
  assign n23607 = ~n23604 & ~n23605;
  assign n23608 = ~n23606 & ~n23607;
  assign n23609 = n23597 & ~n23608;
  assign n23610 = ~n23597 & n23608;
  assign n23611 = ~n23609 & ~n23610;
  assign n23612 = ~n23441 & ~n23443;
  assign n23613 = n23611 & n23612;
  assign n23614 = ~n23611 & ~n23612;
  assign n23615 = ~n23613 & ~n23614;
  assign n23616 = ~n23571 & n23615;
  assign n23617 = n23571 & ~n23615;
  assign n23618 = ~n23616 & ~n23617;
  assign n23619 = n23560 & ~n23618;
  assign n23620 = ~n23560 & n23618;
  assign n23621 = ~n23619 & ~n23620;
  assign n23622 = pi112  & n9096;
  assign n23623 = pi110  & n9453;
  assign n23624 = pi111  & n9091;
  assign n23625 = ~n23623 & ~n23624;
  assign n23626 = ~n23622 & n23625;
  assign n23627 = n7795 & n9099;
  assign n23628 = n23626 & ~n23627;
  assign n23629 = pi53  & ~n23628;
  assign n23630 = pi53  & ~n23629;
  assign n23631 = ~n23628 & ~n23629;
  assign n23632 = ~n23630 & ~n23631;
  assign n23633 = n23621 & ~n23632;
  assign n23634 = ~n23621 & n23632;
  assign n23635 = ~n23633 & ~n23634;
  assign n23636 = n23559 & ~n23635;
  assign n23637 = ~n23559 & n23635;
  assign n23638 = ~n23636 & ~n23637;
  assign n23639 = pi115  & n8137;
  assign n23640 = pi113  & n8471;
  assign n23641 = pi114  & n8132;
  assign n23642 = ~n23640 & ~n23641;
  assign n23643 = ~n23639 & n23642;
  assign n23644 = n8140 & n8727;
  assign n23645 = n23643 & ~n23644;
  assign n23646 = pi50  & ~n23645;
  assign n23647 = pi50  & ~n23646;
  assign n23648 = ~n23645 & ~n23646;
  assign n23649 = ~n23647 & ~n23648;
  assign n23650 = ~n23638 & n23649;
  assign n23651 = n23638 & ~n23649;
  assign n23652 = ~n23650 & ~n23651;
  assign n23653 = ~n23558 & n23652;
  assign n23654 = n23558 & ~n23652;
  assign n23655 = ~n23653 & ~n23654;
  assign n23656 = ~n23557 & n23655;
  assign n23657 = n23557 & ~n23655;
  assign n23658 = ~n23656 & ~n23657;
  assign n23659 = ~n23546 & n23658;
  assign n23660 = n23546 & ~n23658;
  assign n23661 = ~n23659 & ~n23660;
  assign n23662 = pi121  & n6396;
  assign n23663 = pi119  & n6735;
  assign n23664 = pi120  & n6391;
  assign n23665 = ~n23663 & ~n23664;
  assign n23666 = ~n23662 & n23665;
  assign n23667 = n6399 & n11086;
  assign n23668 = n23666 & ~n23667;
  assign n23669 = pi44  & ~n23668;
  assign n23670 = pi44  & ~n23669;
  assign n23671 = ~n23668 & ~n23669;
  assign n23672 = ~n23670 & ~n23671;
  assign n23673 = n23661 & ~n23672;
  assign n23674 = n23661 & ~n23673;
  assign n23675 = ~n23672 & ~n23673;
  assign n23676 = ~n23674 & ~n23675;
  assign n23677 = ~n23492 & ~n23495;
  assign n23678 = n23676 & n23677;
  assign n23679 = ~n23676 & ~n23677;
  assign n23680 = ~n23678 & ~n23679;
  assign n23681 = pi124  & n5636;
  assign n23682 = pi122  & n5909;
  assign n23683 = pi123  & n5631;
  assign n23684 = ~n23682 & ~n23683;
  assign n23685 = ~n23681 & n23684;
  assign n23686 = n5639 & n11858;
  assign n23687 = n23685 & ~n23686;
  assign n23688 = pi41  & ~n23687;
  assign n23689 = pi41  & ~n23688;
  assign n23690 = ~n23687 & ~n23688;
  assign n23691 = ~n23689 & ~n23690;
  assign n23692 = n23680 & ~n23691;
  assign n23693 = ~n23680 & n23691;
  assign n23694 = ~n23692 & ~n23693;
  assign n23695 = n23545 & ~n23694;
  assign n23696 = ~n23545 & n23694;
  assign n23697 = ~n23695 & ~n23696;
  assign n23698 = pi127  & n4896;
  assign n23699 = pi125  & n5148;
  assign n23700 = pi126  & n4891;
  assign n23701 = ~n23699 & ~n23700;
  assign n23702 = ~n23698 & n23701;
  assign n23703 = n4899 & n13365;
  assign n23704 = n23702 & ~n23703;
  assign n23705 = pi38  & ~n23704;
  assign n23706 = pi38  & ~n23705;
  assign n23707 = ~n23704 & ~n23705;
  assign n23708 = ~n23706 & ~n23707;
  assign n23709 = n23697 & ~n23708;
  assign n23710 = ~n23697 & n23708;
  assign n23711 = ~n23709 & ~n23710;
  assign n23712 = n23544 & ~n23711;
  assign n23713 = ~n23544 & n23711;
  assign n23714 = ~n23712 & ~n23713;
  assign n23715 = ~n23365 & ~n23534;
  assign n23716 = n23714 & n23715;
  assign n23717 = ~n23714 & ~n23715;
  assign n23718 = ~n23716 & ~n23717;
  assign n23719 = ~n23543 & n23718;
  assign n23720 = n23543 & ~n23718;
  assign po99  = ~n23719 & ~n23720;
  assign n23722 = ~n23692 & ~n23696;
  assign n23723 = pi126  & n5148;
  assign n23724 = pi127  & n4891;
  assign n23725 = ~n23723 & ~n23724;
  assign n23726 = ~n4899 & n23725;
  assign n23727 = ~n13389 & n23725;
  assign n23728 = ~n23726 & ~n23727;
  assign n23729 = pi38  & ~n23728;
  assign n23730 = ~pi38  & n23728;
  assign n23731 = ~n23729 & ~n23730;
  assign n23732 = ~n23722 & ~n23731;
  assign n23733 = n23722 & n23731;
  assign n23734 = ~n23732 & ~n23733;
  assign n23735 = ~n23673 & ~n23679;
  assign n23736 = ~n23656 & ~n23659;
  assign n23737 = pi119  & n7239;
  assign n23738 = pi117  & n7556;
  assign n23739 = pi118  & n7234;
  assign n23740 = ~n23738 & ~n23739;
  assign n23741 = ~n23737 & n23740;
  assign n23742 = n7242 & n10048;
  assign n23743 = n23741 & ~n23742;
  assign n23744 = pi47  & ~n23743;
  assign n23745 = pi47  & ~n23744;
  assign n23746 = ~n23743 & ~n23744;
  assign n23747 = ~n23745 & ~n23746;
  assign n23748 = ~n23651 & ~n23653;
  assign n23749 = ~n23633 & ~n23637;
  assign n23750 = ~n23609 & ~n23613;
  assign n23751 = ~n23581 & ~n23596;
  assign n23752 = pi104  & n12295;
  assign n23753 = pi102  & n12693;
  assign n23754 = pi103  & n12290;
  assign n23755 = ~n23753 & ~n23754;
  assign n23756 = ~n23752 & n23755;
  assign n23757 = n5565 & n12298;
  assign n23758 = n23756 & ~n23757;
  assign n23759 = pi62  & ~n23758;
  assign n23760 = pi62  & ~n23759;
  assign n23761 = ~n23758 & ~n23759;
  assign n23762 = ~n23760 & ~n23761;
  assign n23763 = pi100  & n13477;
  assign n23764 = pi101  & ~n13122;
  assign n23765 = ~n23763 & ~n23764;
  assign n23766 = ~n23575 & ~n23578;
  assign n23767 = n23765 & ~n23766;
  assign n23768 = ~n23765 & n23766;
  assign n23769 = ~n23767 & ~n23768;
  assign n23770 = ~n23762 & n23769;
  assign n23771 = n23762 & ~n23769;
  assign n23772 = ~n23770 & ~n23771;
  assign n23773 = n23751 & ~n23772;
  assign n23774 = ~n23751 & n23772;
  assign n23775 = ~n23773 & ~n23774;
  assign n23776 = pi107  & n11193;
  assign n23777 = pi105  & n11567;
  assign n23778 = pi106  & n11188;
  assign n23779 = ~n23777 & ~n23778;
  assign n23780 = ~n23776 & n23779;
  assign n23781 = n6614 & n11196;
  assign n23782 = n23780 & ~n23781;
  assign n23783 = pi59  & ~n23782;
  assign n23784 = pi59  & ~n23783;
  assign n23785 = ~n23782 & ~n23783;
  assign n23786 = ~n23784 & ~n23785;
  assign n23787 = n23775 & ~n23786;
  assign n23788 = ~n23775 & n23786;
  assign n23789 = ~n23787 & ~n23788;
  assign n23790 = n23750 & ~n23789;
  assign n23791 = ~n23750 & n23789;
  assign n23792 = ~n23790 & ~n23791;
  assign n23793 = pi110  & n10135;
  assign n23794 = pi108  & n10478;
  assign n23795 = pi109  & n10130;
  assign n23796 = ~n23794 & ~n23795;
  assign n23797 = ~n23793 & n23796;
  assign n23798 = n7474 & n10138;
  assign n23799 = n23797 & ~n23798;
  assign n23800 = pi56  & ~n23799;
  assign n23801 = pi56  & ~n23800;
  assign n23802 = ~n23799 & ~n23800;
  assign n23803 = ~n23801 & ~n23802;
  assign n23804 = n23792 & ~n23803;
  assign n23805 = n23792 & ~n23804;
  assign n23806 = ~n23803 & ~n23804;
  assign n23807 = ~n23805 & ~n23806;
  assign n23808 = ~n23616 & ~n23620;
  assign n23809 = n23807 & n23808;
  assign n23810 = ~n23807 & ~n23808;
  assign n23811 = ~n23809 & ~n23810;
  assign n23812 = pi113  & n9096;
  assign n23813 = pi111  & n9453;
  assign n23814 = pi112  & n9091;
  assign n23815 = ~n23813 & ~n23814;
  assign n23816 = ~n23812 & n23815;
  assign n23817 = n8387 & n9099;
  assign n23818 = n23816 & ~n23817;
  assign n23819 = pi53  & ~n23818;
  assign n23820 = pi53  & ~n23819;
  assign n23821 = ~n23818 & ~n23819;
  assign n23822 = ~n23820 & ~n23821;
  assign n23823 = n23811 & ~n23822;
  assign n23824 = ~n23811 & n23822;
  assign n23825 = ~n23823 & ~n23824;
  assign n23826 = n23749 & ~n23825;
  assign n23827 = ~n23749 & n23825;
  assign n23828 = ~n23826 & ~n23827;
  assign n23829 = pi116  & n8137;
  assign n23830 = pi114  & n8471;
  assign n23831 = pi115  & n8132;
  assign n23832 = ~n23830 & ~n23831;
  assign n23833 = ~n23829 & n23832;
  assign n23834 = n8140 & n9042;
  assign n23835 = n23833 & ~n23834;
  assign n23836 = pi50  & ~n23835;
  assign n23837 = pi50  & ~n23836;
  assign n23838 = ~n23835 & ~n23836;
  assign n23839 = ~n23837 & ~n23838;
  assign n23840 = n23828 & ~n23839;
  assign n23841 = ~n23828 & n23839;
  assign n23842 = ~n23840 & ~n23841;
  assign n23843 = ~n23748 & n23842;
  assign n23844 = n23748 & ~n23842;
  assign n23845 = ~n23843 & ~n23844;
  assign n23846 = ~n23747 & n23845;
  assign n23847 = n23747 & ~n23845;
  assign n23848 = ~n23846 & ~n23847;
  assign n23849 = n23736 & ~n23848;
  assign n23850 = ~n23736 & n23848;
  assign n23851 = ~n23849 & ~n23850;
  assign n23852 = pi122  & n6396;
  assign n23853 = pi120  & n6735;
  assign n23854 = pi121  & n6391;
  assign n23855 = ~n23853 & ~n23854;
  assign n23856 = ~n23852 & n23855;
  assign n23857 = n6399 & n11463;
  assign n23858 = n23856 & ~n23857;
  assign n23859 = pi44  & ~n23858;
  assign n23860 = pi44  & ~n23859;
  assign n23861 = ~n23858 & ~n23859;
  assign n23862 = ~n23860 & ~n23861;
  assign n23863 = n23851 & ~n23862;
  assign n23864 = ~n23851 & n23862;
  assign n23865 = ~n23863 & ~n23864;
  assign n23866 = n23735 & ~n23865;
  assign n23867 = ~n23735 & n23865;
  assign n23868 = ~n23866 & ~n23867;
  assign n23869 = pi125  & n5636;
  assign n23870 = pi123  & n5909;
  assign n23871 = pi124  & n5631;
  assign n23872 = ~n23870 & ~n23871;
  assign n23873 = ~n23869 & n23872;
  assign n23874 = n5639 & n12591;
  assign n23875 = n23873 & ~n23874;
  assign n23876 = pi41  & ~n23875;
  assign n23877 = pi41  & ~n23876;
  assign n23878 = ~n23875 & ~n23876;
  assign n23879 = ~n23877 & ~n23878;
  assign n23880 = n23868 & ~n23879;
  assign n23881 = ~n23868 & n23879;
  assign n23882 = n23734 & ~n23881;
  assign n23883 = ~n23880 & n23882;
  assign n23884 = n23734 & ~n23883;
  assign n23885 = ~n23881 & ~n23883;
  assign n23886 = ~n23880 & n23885;
  assign n23887 = ~n23884 & ~n23886;
  assign n23888 = ~n23709 & ~n23713;
  assign n23889 = n23887 & n23888;
  assign n23890 = ~n23887 & ~n23888;
  assign n23891 = ~n23889 & ~n23890;
  assign n23892 = ~n23716 & ~n23719;
  assign n23893 = n23891 & ~n23892;
  assign n23894 = ~n23891 & n23892;
  assign po100  = ~n23893 & ~n23894;
  assign n23896 = ~n23890 & ~n23893;
  assign n23897 = ~n23732 & ~n23883;
  assign n23898 = ~n23867 & ~n23880;
  assign n23899 = pi127  & n5148;
  assign n23900 = n4899 & n13387;
  assign n23901 = ~n23899 & ~n23900;
  assign n23902 = pi38  & ~n23901;
  assign n23903 = pi38  & ~n23902;
  assign n23904 = ~n23901 & ~n23902;
  assign n23905 = ~n23903 & ~n23904;
  assign n23906 = ~n23898 & ~n23905;
  assign n23907 = n23898 & n23905;
  assign n23908 = ~n23906 & ~n23907;
  assign n23909 = ~n23843 & ~n23846;
  assign n23910 = pi120  & n7239;
  assign n23911 = pi118  & n7556;
  assign n23912 = pi119  & n7234;
  assign n23913 = ~n23911 & ~n23912;
  assign n23914 = ~n23910 & n23913;
  assign n23915 = n7242 & n10734;
  assign n23916 = n23914 & ~n23915;
  assign n23917 = pi47  & ~n23916;
  assign n23918 = pi47  & ~n23917;
  assign n23919 = ~n23916 & ~n23917;
  assign n23920 = ~n23918 & ~n23919;
  assign n23921 = ~n23827 & ~n23840;
  assign n23922 = pi117  & n8137;
  assign n23923 = pi115  & n8471;
  assign n23924 = pi116  & n8132;
  assign n23925 = ~n23923 & ~n23924;
  assign n23926 = ~n23922 & n23925;
  assign n23927 = n8140 & n9691;
  assign n23928 = n23926 & ~n23927;
  assign n23929 = pi50  & ~n23928;
  assign n23930 = pi50  & ~n23929;
  assign n23931 = ~n23928 & ~n23929;
  assign n23932 = ~n23930 & ~n23931;
  assign n23933 = ~n23810 & ~n23823;
  assign n23934 = ~n23791 & ~n23804;
  assign n23935 = ~n23774 & ~n23787;
  assign n23936 = ~n23767 & ~n23770;
  assign n23937 = pi101  & n13477;
  assign n23938 = pi102  & ~n13122;
  assign n23939 = ~n23937 & ~n23938;
  assign n23940 = n23765 & ~n23939;
  assign n23941 = ~n23765 & n23939;
  assign n23942 = ~n23940 & ~n23941;
  assign n23943 = ~n23936 & n23942;
  assign n23944 = n23936 & ~n23942;
  assign n23945 = ~n23943 & ~n23944;
  assign n23946 = pi105  & n12295;
  assign n23947 = pi103  & n12693;
  assign n23948 = pi104  & n12290;
  assign n23949 = ~n23947 & ~n23948;
  assign n23950 = ~n23946 & n23949;
  assign n23951 = n6065 & n12298;
  assign n23952 = n23950 & ~n23951;
  assign n23953 = pi62  & ~n23952;
  assign n23954 = pi62  & ~n23953;
  assign n23955 = ~n23952 & ~n23953;
  assign n23956 = ~n23954 & ~n23955;
  assign n23957 = n23945 & ~n23956;
  assign n23958 = n23945 & ~n23957;
  assign n23959 = ~n23956 & ~n23957;
  assign n23960 = ~n23958 & ~n23959;
  assign n23961 = pi108  & n11193;
  assign n23962 = pi106  & n11567;
  assign n23963 = pi107  & n11188;
  assign n23964 = ~n23962 & ~n23963;
  assign n23965 = ~n23961 & n23964;
  assign n23966 = n6639 & n11196;
  assign n23967 = n23965 & ~n23966;
  assign n23968 = pi59  & ~n23967;
  assign n23969 = pi59  & ~n23968;
  assign n23970 = ~n23967 & ~n23968;
  assign n23971 = ~n23969 & ~n23970;
  assign n23972 = ~n23960 & ~n23971;
  assign n23973 = n23960 & n23971;
  assign n23974 = ~n23972 & ~n23973;
  assign n23975 = n23935 & ~n23974;
  assign n23976 = ~n23935 & n23974;
  assign n23977 = ~n23975 & ~n23976;
  assign n23978 = pi111  & n10135;
  assign n23979 = pi109  & n10478;
  assign n23980 = pi110  & n10130;
  assign n23981 = ~n23979 & ~n23980;
  assign n23982 = ~n23978 & n23981;
  assign n23983 = n7770 & n10138;
  assign n23984 = n23982 & ~n23983;
  assign n23985 = pi56  & ~n23984;
  assign n23986 = pi56  & ~n23985;
  assign n23987 = ~n23984 & ~n23985;
  assign n23988 = ~n23986 & ~n23987;
  assign n23989 = n23977 & ~n23988;
  assign n23990 = ~n23977 & n23988;
  assign n23991 = ~n23989 & ~n23990;
  assign n23992 = n23934 & ~n23991;
  assign n23993 = ~n23934 & n23991;
  assign n23994 = ~n23992 & ~n23993;
  assign n23995 = pi114  & n9096;
  assign n23996 = pi112  & n9453;
  assign n23997 = pi113  & n9091;
  assign n23998 = ~n23996 & ~n23997;
  assign n23999 = ~n23995 & n23998;
  assign n24000 = n8702 & n9099;
  assign n24001 = n23999 & ~n24000;
  assign n24002 = pi53  & ~n24001;
  assign n24003 = pi53  & ~n24002;
  assign n24004 = ~n24001 & ~n24002;
  assign n24005 = ~n24003 & ~n24004;
  assign n24006 = ~n23994 & n24005;
  assign n24007 = n23994 & ~n24005;
  assign n24008 = ~n24006 & ~n24007;
  assign n24009 = ~n23933 & n24008;
  assign n24010 = ~n23933 & ~n24009;
  assign n24011 = n24008 & ~n24009;
  assign n24012 = ~n24010 & ~n24011;
  assign n24013 = ~n23932 & ~n24012;
  assign n24014 = n23932 & n24012;
  assign n24015 = ~n24013 & ~n24014;
  assign n24016 = ~n23921 & n24015;
  assign n24017 = n23921 & ~n24015;
  assign n24018 = ~n24016 & ~n24017;
  assign n24019 = ~n23920 & n24018;
  assign n24020 = n23920 & ~n24018;
  assign n24021 = ~n24019 & ~n24020;
  assign n24022 = ~n23909 & n24021;
  assign n24023 = n23909 & ~n24021;
  assign n24024 = ~n24022 & ~n24023;
  assign n24025 = pi123  & n6396;
  assign n24026 = pi121  & n6735;
  assign n24027 = pi122  & n6391;
  assign n24028 = ~n24026 & ~n24027;
  assign n24029 = ~n24025 & n24028;
  assign n24030 = n6399 & n11489;
  assign n24031 = n24029 & ~n24030;
  assign n24032 = pi44  & ~n24031;
  assign n24033 = pi44  & ~n24032;
  assign n24034 = ~n24031 & ~n24032;
  assign n24035 = ~n24033 & ~n24034;
  assign n24036 = n24024 & ~n24035;
  assign n24037 = n24024 & ~n24036;
  assign n24038 = ~n24035 & ~n24036;
  assign n24039 = ~n24037 & ~n24038;
  assign n24040 = ~n23850 & ~n23863;
  assign n24041 = n24039 & n24040;
  assign n24042 = ~n24039 & ~n24040;
  assign n24043 = ~n24041 & ~n24042;
  assign n24044 = pi126  & n5636;
  assign n24045 = pi124  & n5909;
  assign n24046 = pi125  & n5631;
  assign n24047 = ~n24045 & ~n24046;
  assign n24048 = ~n24044 & n24047;
  assign n24049 = n5639 & n12979;
  assign n24050 = n24048 & ~n24049;
  assign n24051 = pi41  & ~n24050;
  assign n24052 = pi41  & ~n24051;
  assign n24053 = ~n24050 & ~n24051;
  assign n24054 = ~n24052 & ~n24053;
  assign n24055 = n24043 & ~n24054;
  assign n24056 = ~n24043 & n24054;
  assign n24057 = ~n24055 & ~n24056;
  assign n24058 = n23908 & ~n24057;
  assign n24059 = ~n23908 & n24057;
  assign n24060 = ~n24058 & ~n24059;
  assign n24061 = ~n23897 & ~n24060;
  assign n24062 = n23897 & n24060;
  assign n24063 = ~n24061 & ~n24062;
  assign n24064 = ~n23896 & n24063;
  assign n24065 = n23896 & ~n24063;
  assign po101  = ~n24064 & ~n24065;
  assign n24067 = ~n24061 & ~n24064;
  assign n24068 = ~n24042 & ~n24055;
  assign n24069 = ~n24022 & ~n24036;
  assign n24070 = ~n24009 & ~n24013;
  assign n24071 = pi118  & n8137;
  assign n24072 = pi116  & n8471;
  assign n24073 = pi117  & n8132;
  assign n24074 = ~n24072 & ~n24073;
  assign n24075 = ~n24071 & n24074;
  assign n24076 = n8140 & n9716;
  assign n24077 = n24075 & ~n24076;
  assign n24078 = pi50  & ~n24077;
  assign n24079 = pi50  & ~n24078;
  assign n24080 = ~n24077 & ~n24078;
  assign n24081 = ~n24079 & ~n24080;
  assign n24082 = ~n23993 & ~n24007;
  assign n24083 = ~n23976 & ~n23989;
  assign n24084 = pi112  & n10135;
  assign n24085 = pi110  & n10478;
  assign n24086 = pi111  & n10130;
  assign n24087 = ~n24085 & ~n24086;
  assign n24088 = ~n24084 & n24087;
  assign n24089 = n7795 & n10138;
  assign n24090 = n24088 & ~n24089;
  assign n24091 = pi56  & ~n24090;
  assign n24092 = pi56  & ~n24091;
  assign n24093 = ~n24090 & ~n24091;
  assign n24094 = ~n24092 & ~n24093;
  assign n24095 = ~n23957 & ~n23972;
  assign n24096 = ~n23940 & ~n23943;
  assign n24097 = pi102  & n13477;
  assign n24098 = pi103  & ~n13122;
  assign n24099 = ~n24097 & ~n24098;
  assign n24100 = ~pi38  & ~n23765;
  assign n24101 = pi38  & n23765;
  assign n24102 = ~n24100 & ~n24101;
  assign n24103 = ~n24099 & n24102;
  assign n24104 = n24099 & ~n24102;
  assign n24105 = ~n24103 & ~n24104;
  assign n24106 = ~n24096 & n24105;
  assign n24107 = n24096 & ~n24105;
  assign n24108 = ~n24106 & ~n24107;
  assign n24109 = pi106  & n12295;
  assign n24110 = pi104  & n12693;
  assign n24111 = pi105  & n12290;
  assign n24112 = ~n24110 & ~n24111;
  assign n24113 = ~n24109 & n24112;
  assign n24114 = n6090 & n12298;
  assign n24115 = n24113 & ~n24114;
  assign n24116 = pi62  & ~n24115;
  assign n24117 = pi62  & ~n24116;
  assign n24118 = ~n24115 & ~n24116;
  assign n24119 = ~n24117 & ~n24118;
  assign n24120 = n24108 & ~n24119;
  assign n24121 = n24108 & ~n24120;
  assign n24122 = ~n24119 & ~n24120;
  assign n24123 = ~n24121 & ~n24122;
  assign n24124 = pi109  & n11193;
  assign n24125 = pi107  & n11567;
  assign n24126 = pi108  & n11188;
  assign n24127 = ~n24125 & ~n24126;
  assign n24128 = ~n24124 & n24127;
  assign n24129 = n7170 & n11196;
  assign n24130 = n24128 & ~n24129;
  assign n24131 = pi59  & ~n24130;
  assign n24132 = pi59  & ~n24131;
  assign n24133 = ~n24130 & ~n24131;
  assign n24134 = ~n24132 & ~n24133;
  assign n24135 = ~n24123 & ~n24134;
  assign n24136 = n24123 & n24134;
  assign n24137 = ~n24135 & ~n24136;
  assign n24138 = ~n24095 & n24137;
  assign n24139 = n24095 & ~n24137;
  assign n24140 = ~n24138 & ~n24139;
  assign n24141 = ~n24094 & n24140;
  assign n24142 = n24094 & ~n24140;
  assign n24143 = ~n24141 & ~n24142;
  assign n24144 = n24083 & ~n24143;
  assign n24145 = ~n24083 & n24143;
  assign n24146 = ~n24144 & ~n24145;
  assign n24147 = pi115  & n9096;
  assign n24148 = pi113  & n9453;
  assign n24149 = pi114  & n9091;
  assign n24150 = ~n24148 & ~n24149;
  assign n24151 = ~n24147 & n24150;
  assign n24152 = n8727 & n9099;
  assign n24153 = n24151 & ~n24152;
  assign n24154 = pi53  & ~n24153;
  assign n24155 = pi53  & ~n24154;
  assign n24156 = ~n24153 & ~n24154;
  assign n24157 = ~n24155 & ~n24156;
  assign n24158 = ~n24146 & n24157;
  assign n24159 = n24146 & ~n24157;
  assign n24160 = ~n24158 & ~n24159;
  assign n24161 = ~n24082 & n24160;
  assign n24162 = n24082 & ~n24160;
  assign n24163 = ~n24161 & ~n24162;
  assign n24164 = ~n24081 & n24163;
  assign n24165 = n24081 & ~n24163;
  assign n24166 = ~n24164 & ~n24165;
  assign n24167 = ~n24070 & n24166;
  assign n24168 = n24070 & ~n24166;
  assign n24169 = ~n24167 & ~n24168;
  assign n24170 = pi121  & n7239;
  assign n24171 = pi119  & n7556;
  assign n24172 = pi120  & n7234;
  assign n24173 = ~n24171 & ~n24172;
  assign n24174 = ~n24170 & n24173;
  assign n24175 = n7242 & n11086;
  assign n24176 = n24174 & ~n24175;
  assign n24177 = pi47  & ~n24176;
  assign n24178 = pi47  & ~n24177;
  assign n24179 = ~n24176 & ~n24177;
  assign n24180 = ~n24178 & ~n24179;
  assign n24181 = n24169 & ~n24180;
  assign n24182 = n24169 & ~n24181;
  assign n24183 = ~n24180 & ~n24181;
  assign n24184 = ~n24182 & ~n24183;
  assign n24185 = ~n24016 & ~n24019;
  assign n24186 = n24184 & n24185;
  assign n24187 = ~n24184 & ~n24185;
  assign n24188 = ~n24186 & ~n24187;
  assign n24189 = pi124  & n6396;
  assign n24190 = pi122  & n6735;
  assign n24191 = pi123  & n6391;
  assign n24192 = ~n24190 & ~n24191;
  assign n24193 = ~n24189 & n24192;
  assign n24194 = n6399 & n11858;
  assign n24195 = n24193 & ~n24194;
  assign n24196 = pi44  & ~n24195;
  assign n24197 = pi44  & ~n24196;
  assign n24198 = ~n24195 & ~n24196;
  assign n24199 = ~n24197 & ~n24198;
  assign n24200 = n24188 & ~n24199;
  assign n24201 = ~n24188 & n24199;
  assign n24202 = ~n24200 & ~n24201;
  assign n24203 = n24069 & ~n24202;
  assign n24204 = ~n24069 & n24202;
  assign n24205 = ~n24203 & ~n24204;
  assign n24206 = pi127  & n5636;
  assign n24207 = pi125  & n5909;
  assign n24208 = pi126  & n5631;
  assign n24209 = ~n24207 & ~n24208;
  assign n24210 = ~n24206 & n24209;
  assign n24211 = n5639 & n13365;
  assign n24212 = n24210 & ~n24211;
  assign n24213 = pi41  & ~n24212;
  assign n24214 = pi41  & ~n24213;
  assign n24215 = ~n24212 & ~n24213;
  assign n24216 = ~n24214 & ~n24215;
  assign n24217 = n24205 & ~n24216;
  assign n24218 = ~n24205 & n24216;
  assign n24219 = ~n24217 & ~n24218;
  assign n24220 = n24068 & ~n24219;
  assign n24221 = ~n24068 & n24219;
  assign n24222 = ~n24220 & ~n24221;
  assign n24223 = ~n23907 & ~n24058;
  assign n24224 = n24222 & n24223;
  assign n24225 = ~n24222 & ~n24223;
  assign n24226 = ~n24224 & ~n24225;
  assign n24227 = ~n24067 & n24226;
  assign n24228 = n24067 & ~n24226;
  assign po102  = ~n24227 & ~n24228;
  assign n24230 = ~n24200 & ~n24204;
  assign n24231 = pi126  & n5909;
  assign n24232 = pi127  & n5631;
  assign n24233 = ~n24231 & ~n24232;
  assign n24234 = ~n5639 & n24233;
  assign n24235 = ~n13389 & n24233;
  assign n24236 = ~n24234 & ~n24235;
  assign n24237 = pi41  & ~n24236;
  assign n24238 = ~pi41  & n24236;
  assign n24239 = ~n24237 & ~n24238;
  assign n24240 = ~n24230 & ~n24239;
  assign n24241 = n24230 & n24239;
  assign n24242 = ~n24240 & ~n24241;
  assign n24243 = ~n24181 & ~n24187;
  assign n24244 = ~n24164 & ~n24167;
  assign n24245 = pi119  & n8137;
  assign n24246 = pi117  & n8471;
  assign n24247 = pi118  & n8132;
  assign n24248 = ~n24246 & ~n24247;
  assign n24249 = ~n24245 & n24248;
  assign n24250 = n8140 & n10048;
  assign n24251 = n24249 & ~n24250;
  assign n24252 = pi50  & ~n24251;
  assign n24253 = pi50  & ~n24252;
  assign n24254 = ~n24251 & ~n24252;
  assign n24255 = ~n24253 & ~n24254;
  assign n24256 = ~n24159 & ~n24161;
  assign n24257 = ~n24141 & ~n24145;
  assign n24258 = ~n24106 & ~n24120;
  assign n24259 = pi103  & n13477;
  assign n24260 = pi104  & ~n13122;
  assign n24261 = ~n24259 & ~n24260;
  assign n24262 = ~n24100 & ~n24103;
  assign n24263 = n24261 & ~n24262;
  assign n24264 = ~n24261 & n24262;
  assign n24265 = ~n24263 & ~n24264;
  assign n24266 = pi107  & n12295;
  assign n24267 = pi105  & n12693;
  assign n24268 = pi106  & n12290;
  assign n24269 = ~n24267 & ~n24268;
  assign n24270 = ~n24266 & n24269;
  assign n24271 = ~n12298 & n24270;
  assign n24272 = ~n6614 & n24270;
  assign n24273 = ~n24271 & ~n24272;
  assign n24274 = pi62  & ~n24273;
  assign n24275 = ~pi62  & n24273;
  assign n24276 = ~n24274 & ~n24275;
  assign n24277 = n24265 & ~n24276;
  assign n24278 = ~n24265 & n24276;
  assign n24279 = ~n24277 & ~n24278;
  assign n24280 = ~n24258 & n24279;
  assign n24281 = n24258 & ~n24279;
  assign n24282 = ~n24280 & ~n24281;
  assign n24283 = pi110  & n11193;
  assign n24284 = pi108  & n11567;
  assign n24285 = pi109  & n11188;
  assign n24286 = ~n24284 & ~n24285;
  assign n24287 = ~n24283 & n24286;
  assign n24288 = n7474 & n11196;
  assign n24289 = n24287 & ~n24288;
  assign n24290 = pi59  & ~n24289;
  assign n24291 = pi59  & ~n24290;
  assign n24292 = ~n24289 & ~n24290;
  assign n24293 = ~n24291 & ~n24292;
  assign n24294 = n24282 & ~n24293;
  assign n24295 = n24282 & ~n24294;
  assign n24296 = ~n24293 & ~n24294;
  assign n24297 = ~n24295 & ~n24296;
  assign n24298 = ~n24135 & ~n24138;
  assign n24299 = n24297 & n24298;
  assign n24300 = ~n24297 & ~n24298;
  assign n24301 = ~n24299 & ~n24300;
  assign n24302 = pi113  & n10135;
  assign n24303 = pi111  & n10478;
  assign n24304 = pi112  & n10130;
  assign n24305 = ~n24303 & ~n24304;
  assign n24306 = ~n24302 & n24305;
  assign n24307 = n8387 & n10138;
  assign n24308 = n24306 & ~n24307;
  assign n24309 = pi56  & ~n24308;
  assign n24310 = pi56  & ~n24309;
  assign n24311 = ~n24308 & ~n24309;
  assign n24312 = ~n24310 & ~n24311;
  assign n24313 = n24301 & ~n24312;
  assign n24314 = ~n24301 & n24312;
  assign n24315 = ~n24313 & ~n24314;
  assign n24316 = n24257 & ~n24315;
  assign n24317 = ~n24257 & n24315;
  assign n24318 = ~n24316 & ~n24317;
  assign n24319 = pi116  & n9096;
  assign n24320 = pi114  & n9453;
  assign n24321 = pi115  & n9091;
  assign n24322 = ~n24320 & ~n24321;
  assign n24323 = ~n24319 & n24322;
  assign n24324 = n9042 & n9099;
  assign n24325 = n24323 & ~n24324;
  assign n24326 = pi53  & ~n24325;
  assign n24327 = pi53  & ~n24326;
  assign n24328 = ~n24325 & ~n24326;
  assign n24329 = ~n24327 & ~n24328;
  assign n24330 = n24318 & ~n24329;
  assign n24331 = ~n24318 & n24329;
  assign n24332 = ~n24330 & ~n24331;
  assign n24333 = ~n24256 & n24332;
  assign n24334 = n24256 & ~n24332;
  assign n24335 = ~n24333 & ~n24334;
  assign n24336 = ~n24255 & n24335;
  assign n24337 = n24255 & ~n24335;
  assign n24338 = ~n24336 & ~n24337;
  assign n24339 = n24244 & ~n24338;
  assign n24340 = ~n24244 & n24338;
  assign n24341 = ~n24339 & ~n24340;
  assign n24342 = pi122  & n7239;
  assign n24343 = pi120  & n7556;
  assign n24344 = pi121  & n7234;
  assign n24345 = ~n24343 & ~n24344;
  assign n24346 = ~n24342 & n24345;
  assign n24347 = n7242 & n11463;
  assign n24348 = n24346 & ~n24347;
  assign n24349 = pi47  & ~n24348;
  assign n24350 = pi47  & ~n24349;
  assign n24351 = ~n24348 & ~n24349;
  assign n24352 = ~n24350 & ~n24351;
  assign n24353 = n24341 & ~n24352;
  assign n24354 = ~n24341 & n24352;
  assign n24355 = ~n24353 & ~n24354;
  assign n24356 = n24243 & ~n24355;
  assign n24357 = ~n24243 & n24355;
  assign n24358 = ~n24356 & ~n24357;
  assign n24359 = pi125  & n6396;
  assign n24360 = pi123  & n6735;
  assign n24361 = pi124  & n6391;
  assign n24362 = ~n24360 & ~n24361;
  assign n24363 = ~n24359 & n24362;
  assign n24364 = n6399 & n12591;
  assign n24365 = n24363 & ~n24364;
  assign n24366 = pi44  & ~n24365;
  assign n24367 = pi44  & ~n24366;
  assign n24368 = ~n24365 & ~n24366;
  assign n24369 = ~n24367 & ~n24368;
  assign n24370 = n24358 & ~n24369;
  assign n24371 = ~n24358 & n24369;
  assign n24372 = n24242 & ~n24371;
  assign n24373 = ~n24370 & n24372;
  assign n24374 = n24242 & ~n24373;
  assign n24375 = ~n24371 & ~n24373;
  assign n24376 = ~n24370 & n24375;
  assign n24377 = ~n24374 & ~n24376;
  assign n24378 = ~n24217 & ~n24221;
  assign n24379 = n24377 & n24378;
  assign n24380 = ~n24377 & ~n24378;
  assign n24381 = ~n24379 & ~n24380;
  assign n24382 = ~n24224 & ~n24227;
  assign n24383 = n24381 & ~n24382;
  assign n24384 = ~n24381 & n24382;
  assign po103  = ~n24383 & ~n24384;
  assign n24386 = ~n24380 & ~n24383;
  assign n24387 = ~n24240 & ~n24373;
  assign n24388 = ~n24357 & ~n24370;
  assign n24389 = pi127  & n5909;
  assign n24390 = n5639 & n13387;
  assign n24391 = ~n24389 & ~n24390;
  assign n24392 = pi41  & ~n24391;
  assign n24393 = pi41  & ~n24392;
  assign n24394 = ~n24391 & ~n24392;
  assign n24395 = ~n24393 & ~n24394;
  assign n24396 = ~n24388 & ~n24395;
  assign n24397 = n24388 & n24395;
  assign n24398 = ~n24396 & ~n24397;
  assign n24399 = ~n24340 & ~n24353;
  assign n24400 = ~n24333 & ~n24336;
  assign n24401 = pi120  & n8137;
  assign n24402 = pi118  & n8471;
  assign n24403 = pi119  & n8132;
  assign n24404 = ~n24402 & ~n24403;
  assign n24405 = ~n24401 & n24404;
  assign n24406 = n8140 & n10734;
  assign n24407 = n24405 & ~n24406;
  assign n24408 = pi50  & ~n24407;
  assign n24409 = pi50  & ~n24408;
  assign n24410 = ~n24407 & ~n24408;
  assign n24411 = ~n24409 & ~n24410;
  assign n24412 = ~n24317 & ~n24330;
  assign n24413 = pi117  & n9096;
  assign n24414 = pi115  & n9453;
  assign n24415 = pi116  & n9091;
  assign n24416 = ~n24414 & ~n24415;
  assign n24417 = ~n24413 & n24416;
  assign n24418 = n9099 & n9691;
  assign n24419 = n24417 & ~n24418;
  assign n24420 = pi53  & ~n24419;
  assign n24421 = pi53  & ~n24420;
  assign n24422 = ~n24419 & ~n24420;
  assign n24423 = ~n24421 & ~n24422;
  assign n24424 = ~n24300 & ~n24313;
  assign n24425 = ~n24280 & ~n24294;
  assign n24426 = pi108  & n12295;
  assign n24427 = pi106  & n12693;
  assign n24428 = pi107  & n12290;
  assign n24429 = ~n24427 & ~n24428;
  assign n24430 = ~n24426 & n24429;
  assign n24431 = n6639 & n12298;
  assign n24432 = n24430 & ~n24431;
  assign n24433 = pi62  & ~n24432;
  assign n24434 = pi62  & ~n24433;
  assign n24435 = ~n24432 & ~n24433;
  assign n24436 = ~n24434 & ~n24435;
  assign n24437 = ~n24263 & ~n24277;
  assign n24438 = pi104  & n13477;
  assign n24439 = pi105  & ~n13122;
  assign n24440 = ~n24438 & ~n24439;
  assign n24441 = n24261 & ~n24440;
  assign n24442 = ~n24261 & n24440;
  assign n24443 = ~n24441 & ~n24442;
  assign n24444 = ~n24437 & n24443;
  assign n24445 = n24437 & ~n24443;
  assign n24446 = ~n24444 & ~n24445;
  assign n24447 = n24436 & n24446;
  assign n24448 = ~n24436 & ~n24446;
  assign n24449 = ~n24447 & ~n24448;
  assign n24450 = pi111  & n11193;
  assign n24451 = pi109  & n11567;
  assign n24452 = pi110  & n11188;
  assign n24453 = ~n24451 & ~n24452;
  assign n24454 = ~n24450 & n24453;
  assign n24455 = n7770 & n11196;
  assign n24456 = n24454 & ~n24455;
  assign n24457 = pi59  & ~n24456;
  assign n24458 = pi59  & ~n24457;
  assign n24459 = ~n24456 & ~n24457;
  assign n24460 = ~n24458 & ~n24459;
  assign n24461 = ~n24449 & ~n24460;
  assign n24462 = n24449 & n24460;
  assign n24463 = ~n24461 & ~n24462;
  assign n24464 = n24425 & ~n24463;
  assign n24465 = ~n24425 & n24463;
  assign n24466 = ~n24464 & ~n24465;
  assign n24467 = pi114  & n10135;
  assign n24468 = pi112  & n10478;
  assign n24469 = pi113  & n10130;
  assign n24470 = ~n24468 & ~n24469;
  assign n24471 = ~n24467 & n24470;
  assign n24472 = n8702 & n10138;
  assign n24473 = n24471 & ~n24472;
  assign n24474 = pi56  & ~n24473;
  assign n24475 = pi56  & ~n24474;
  assign n24476 = ~n24473 & ~n24474;
  assign n24477 = ~n24475 & ~n24476;
  assign n24478 = ~n24466 & n24477;
  assign n24479 = n24466 & ~n24477;
  assign n24480 = ~n24478 & ~n24479;
  assign n24481 = ~n24424 & n24480;
  assign n24482 = n24424 & ~n24480;
  assign n24483 = ~n24481 & ~n24482;
  assign n24484 = ~n24423 & n24483;
  assign n24485 = n24423 & ~n24483;
  assign n24486 = ~n24484 & ~n24485;
  assign n24487 = ~n24412 & n24486;
  assign n24488 = n24412 & ~n24486;
  assign n24489 = ~n24487 & ~n24488;
  assign n24490 = ~n24411 & n24489;
  assign n24491 = n24411 & ~n24489;
  assign n24492 = ~n24490 & ~n24491;
  assign n24493 = ~n24400 & n24492;
  assign n24494 = n24400 & ~n24492;
  assign n24495 = ~n24493 & ~n24494;
  assign n24496 = pi123  & n7239;
  assign n24497 = pi121  & n7556;
  assign n24498 = pi122  & n7234;
  assign n24499 = ~n24497 & ~n24498;
  assign n24500 = ~n24496 & n24499;
  assign n24501 = n7242 & n11489;
  assign n24502 = n24500 & ~n24501;
  assign n24503 = pi47  & ~n24502;
  assign n24504 = pi47  & ~n24503;
  assign n24505 = ~n24502 & ~n24503;
  assign n24506 = ~n24504 & ~n24505;
  assign n24507 = n24495 & ~n24506;
  assign n24508 = ~n24495 & n24506;
  assign n24509 = ~n24507 & ~n24508;
  assign n24510 = n24399 & ~n24509;
  assign n24511 = ~n24399 & n24509;
  assign n24512 = ~n24510 & ~n24511;
  assign n24513 = pi126  & n6396;
  assign n24514 = pi124  & n6735;
  assign n24515 = pi125  & n6391;
  assign n24516 = ~n24514 & ~n24515;
  assign n24517 = ~n24513 & n24516;
  assign n24518 = n6399 & n12979;
  assign n24519 = n24517 & ~n24518;
  assign n24520 = pi44  & ~n24519;
  assign n24521 = pi44  & ~n24520;
  assign n24522 = ~n24519 & ~n24520;
  assign n24523 = ~n24521 & ~n24522;
  assign n24524 = n24512 & ~n24523;
  assign n24525 = ~n24512 & n24523;
  assign n24526 = ~n24524 & ~n24525;
  assign n24527 = n24398 & ~n24526;
  assign n24528 = ~n24398 & n24526;
  assign n24529 = ~n24527 & ~n24528;
  assign n24530 = ~n24387 & ~n24529;
  assign n24531 = n24387 & n24529;
  assign n24532 = ~n24530 & ~n24531;
  assign n24533 = ~n24386 & n24532;
  assign n24534 = n24386 & ~n24532;
  assign po104  = ~n24533 & ~n24534;
  assign n24536 = ~n24530 & ~n24533;
  assign n24537 = ~n24511 & ~n24524;
  assign n24538 = ~n24487 & ~n24490;
  assign n24539 = pi121  & n8137;
  assign n24540 = pi119  & n8471;
  assign n24541 = pi120  & n8132;
  assign n24542 = ~n24540 & ~n24541;
  assign n24543 = ~n24539 & n24542;
  assign n24544 = n8140 & n11086;
  assign n24545 = n24543 & ~n24544;
  assign n24546 = pi50  & ~n24545;
  assign n24547 = pi50  & ~n24546;
  assign n24548 = ~n24545 & ~n24546;
  assign n24549 = ~n24547 & ~n24548;
  assign n24550 = ~n24481 & ~n24484;
  assign n24551 = pi118  & n9096;
  assign n24552 = pi116  & n9453;
  assign n24553 = pi117  & n9091;
  assign n24554 = ~n24552 & ~n24553;
  assign n24555 = ~n24551 & n24554;
  assign n24556 = n9099 & n9716;
  assign n24557 = n24555 & ~n24556;
  assign n24558 = pi53  & ~n24557;
  assign n24559 = pi53  & ~n24558;
  assign n24560 = ~n24557 & ~n24558;
  assign n24561 = ~n24559 & ~n24560;
  assign n24562 = ~n24465 & ~n24479;
  assign n24563 = pi115  & n10135;
  assign n24564 = pi113  & n10478;
  assign n24565 = pi114  & n10130;
  assign n24566 = ~n24564 & ~n24565;
  assign n24567 = ~n24563 & n24566;
  assign n24568 = n8727 & n10138;
  assign n24569 = n24567 & ~n24568;
  assign n24570 = pi56  & ~n24569;
  assign n24571 = pi56  & ~n24570;
  assign n24572 = ~n24569 & ~n24570;
  assign n24573 = ~n24571 & ~n24572;
  assign n24574 = ~n24436 & n24446;
  assign n24575 = ~n24461 & ~n24574;
  assign n24576 = ~n24441 & ~n24444;
  assign n24577 = pi105  & n13477;
  assign n24578 = pi106  & ~n13122;
  assign n24579 = ~n24577 & ~n24578;
  assign n24580 = ~pi41  & ~n24261;
  assign n24581 = pi41  & n24261;
  assign n24582 = ~n24580 & ~n24581;
  assign n24583 = n24579 & ~n24582;
  assign n24584 = ~n24579 & n24582;
  assign n24585 = ~n24583 & ~n24584;
  assign n24586 = pi109  & n12295;
  assign n24587 = pi107  & n12693;
  assign n24588 = pi108  & n12290;
  assign n24589 = ~n24587 & ~n24588;
  assign n24590 = ~n24586 & n24589;
  assign n24591 = n7170 & n12298;
  assign n24592 = n24590 & ~n24591;
  assign n24593 = pi62  & ~n24592;
  assign n24594 = pi62  & ~n24593;
  assign n24595 = ~n24592 & ~n24593;
  assign n24596 = ~n24594 & ~n24595;
  assign n24597 = n24585 & ~n24596;
  assign n24598 = ~n24585 & n24596;
  assign n24599 = ~n24597 & ~n24598;
  assign n24600 = n24576 & ~n24599;
  assign n24601 = ~n24576 & n24599;
  assign n24602 = ~n24600 & ~n24601;
  assign n24603 = pi112  & n11193;
  assign n24604 = pi110  & n11567;
  assign n24605 = pi111  & n11188;
  assign n24606 = ~n24604 & ~n24605;
  assign n24607 = ~n24603 & n24606;
  assign n24608 = n7795 & n11196;
  assign n24609 = n24607 & ~n24608;
  assign n24610 = pi59  & ~n24609;
  assign n24611 = pi59  & ~n24610;
  assign n24612 = ~n24609 & ~n24610;
  assign n24613 = ~n24611 & ~n24612;
  assign n24614 = n24602 & ~n24613;
  assign n24615 = ~n24602 & n24613;
  assign n24616 = ~n24614 & ~n24615;
  assign n24617 = ~n24575 & n24616;
  assign n24618 = n24575 & ~n24616;
  assign n24619 = ~n24617 & ~n24618;
  assign n24620 = ~n24573 & n24619;
  assign n24621 = n24573 & ~n24619;
  assign n24622 = ~n24620 & ~n24621;
  assign n24623 = ~n24562 & n24622;
  assign n24624 = n24562 & ~n24622;
  assign n24625 = ~n24623 & ~n24624;
  assign n24626 = n24561 & ~n24625;
  assign n24627 = ~n24561 & n24625;
  assign n24628 = ~n24626 & ~n24627;
  assign n24629 = ~n24550 & n24628;
  assign n24630 = n24550 & ~n24628;
  assign n24631 = ~n24629 & ~n24630;
  assign n24632 = n24549 & ~n24631;
  assign n24633 = ~n24549 & n24631;
  assign n24634 = ~n24632 & ~n24633;
  assign n24635 = ~n24538 & n24634;
  assign n24636 = n24538 & ~n24634;
  assign n24637 = ~n24635 & ~n24636;
  assign n24638 = pi124  & n7239;
  assign n24639 = pi122  & n7556;
  assign n24640 = pi123  & n7234;
  assign n24641 = ~n24639 & ~n24640;
  assign n24642 = ~n24638 & n24641;
  assign n24643 = n7242 & n11858;
  assign n24644 = n24642 & ~n24643;
  assign n24645 = pi47  & ~n24644;
  assign n24646 = pi47  & ~n24645;
  assign n24647 = ~n24644 & ~n24645;
  assign n24648 = ~n24646 & ~n24647;
  assign n24649 = n24637 & ~n24648;
  assign n24650 = n24637 & ~n24649;
  assign n24651 = ~n24648 & ~n24649;
  assign n24652 = ~n24650 & ~n24651;
  assign n24653 = ~n24493 & ~n24507;
  assign n24654 = n24652 & n24653;
  assign n24655 = ~n24652 & ~n24653;
  assign n24656 = ~n24654 & ~n24655;
  assign n24657 = pi127  & n6396;
  assign n24658 = pi125  & n6735;
  assign n24659 = pi126  & n6391;
  assign n24660 = ~n24658 & ~n24659;
  assign n24661 = ~n24657 & n24660;
  assign n24662 = n6399 & n13365;
  assign n24663 = n24661 & ~n24662;
  assign n24664 = pi44  & ~n24663;
  assign n24665 = pi44  & ~n24664;
  assign n24666 = ~n24663 & ~n24664;
  assign n24667 = ~n24665 & ~n24666;
  assign n24668 = n24656 & ~n24667;
  assign n24669 = ~n24656 & n24667;
  assign n24670 = ~n24668 & ~n24669;
  assign n24671 = n24537 & ~n24670;
  assign n24672 = ~n24537 & n24670;
  assign n24673 = ~n24671 & ~n24672;
  assign n24674 = ~n24397 & ~n24527;
  assign n24675 = n24673 & n24674;
  assign n24676 = ~n24673 & ~n24674;
  assign n24677 = ~n24675 & ~n24676;
  assign n24678 = ~n24536 & n24677;
  assign n24679 = n24536 & ~n24677;
  assign po105  = ~n24678 & ~n24679;
  assign n24681 = ~n24668 & ~n24672;
  assign n24682 = ~n24649 & ~n24655;
  assign n24683 = pi126  & n6735;
  assign n24684 = pi127  & n6391;
  assign n24685 = ~n24683 & ~n24684;
  assign n24686 = ~n6399 & n24685;
  assign n24687 = ~n13389 & n24685;
  assign n24688 = ~n24686 & ~n24687;
  assign n24689 = pi44  & ~n24688;
  assign n24690 = ~pi44  & n24688;
  assign n24691 = ~n24689 & ~n24690;
  assign n24692 = ~n24682 & ~n24691;
  assign n24693 = n24682 & n24691;
  assign n24694 = ~n24692 & ~n24693;
  assign n24695 = pi125  & n7239;
  assign n24696 = pi123  & n7556;
  assign n24697 = pi124  & n7234;
  assign n24698 = ~n24696 & ~n24697;
  assign n24699 = ~n24695 & n24698;
  assign n24700 = n7242 & n12591;
  assign n24701 = n24699 & ~n24700;
  assign n24702 = pi47  & ~n24701;
  assign n24703 = pi47  & ~n24702;
  assign n24704 = ~n24701 & ~n24702;
  assign n24705 = ~n24703 & ~n24704;
  assign n24706 = ~n24633 & ~n24635;
  assign n24707 = pi122  & n8137;
  assign n24708 = pi120  & n8471;
  assign n24709 = pi121  & n8132;
  assign n24710 = ~n24708 & ~n24709;
  assign n24711 = ~n24707 & n24710;
  assign n24712 = n8140 & n11463;
  assign n24713 = n24711 & ~n24712;
  assign n24714 = pi50  & ~n24713;
  assign n24715 = pi50  & ~n24714;
  assign n24716 = ~n24713 & ~n24714;
  assign n24717 = ~n24715 & ~n24716;
  assign n24718 = ~n24627 & ~n24629;
  assign n24719 = ~n24620 & ~n24623;
  assign n24720 = ~n24614 & ~n24617;
  assign n24721 = ~n24597 & ~n24601;
  assign n24722 = pi110  & n12295;
  assign n24723 = pi108  & n12693;
  assign n24724 = pi109  & n12290;
  assign n24725 = ~n24723 & ~n24724;
  assign n24726 = ~n24722 & n24725;
  assign n24727 = ~n12298 & n24726;
  assign n24728 = ~n7474 & n24726;
  assign n24729 = ~n24727 & ~n24728;
  assign n24730 = pi62  & ~n24729;
  assign n24731 = ~pi62  & n24729;
  assign n24732 = ~n24730 & ~n24731;
  assign n24733 = pi106  & n13477;
  assign n24734 = pi107  & ~n13122;
  assign n24735 = ~n24733 & ~n24734;
  assign n24736 = ~n24580 & ~n24584;
  assign n24737 = n24735 & ~n24736;
  assign n24738 = ~n24735 & n24736;
  assign n24739 = ~n24737 & ~n24738;
  assign n24740 = ~n24732 & n24739;
  assign n24741 = n24732 & ~n24739;
  assign n24742 = ~n24740 & ~n24741;
  assign n24743 = ~n24721 & n24742;
  assign n24744 = n24721 & ~n24742;
  assign n24745 = ~n24743 & ~n24744;
  assign n24746 = pi113  & n11193;
  assign n24747 = pi111  & n11567;
  assign n24748 = pi112  & n11188;
  assign n24749 = ~n24747 & ~n24748;
  assign n24750 = ~n24746 & n24749;
  assign n24751 = n8387 & n11196;
  assign n24752 = n24750 & ~n24751;
  assign n24753 = pi59  & ~n24752;
  assign n24754 = pi59  & ~n24753;
  assign n24755 = ~n24752 & ~n24753;
  assign n24756 = ~n24754 & ~n24755;
  assign n24757 = n24745 & ~n24756;
  assign n24758 = ~n24745 & n24756;
  assign n24759 = ~n24757 & ~n24758;
  assign n24760 = n24720 & ~n24759;
  assign n24761 = ~n24720 & n24759;
  assign n24762 = ~n24760 & ~n24761;
  assign n24763 = pi116  & n10135;
  assign n24764 = pi114  & n10478;
  assign n24765 = pi115  & n10130;
  assign n24766 = ~n24764 & ~n24765;
  assign n24767 = ~n24763 & n24766;
  assign n24768 = n9042 & n10138;
  assign n24769 = n24767 & ~n24768;
  assign n24770 = pi56  & ~n24769;
  assign n24771 = pi56  & ~n24770;
  assign n24772 = ~n24769 & ~n24770;
  assign n24773 = ~n24771 & ~n24772;
  assign n24774 = n24762 & ~n24773;
  assign n24775 = ~n24762 & n24773;
  assign n24776 = ~n24774 & ~n24775;
  assign n24777 = n24719 & ~n24776;
  assign n24778 = ~n24719 & n24776;
  assign n24779 = ~n24777 & ~n24778;
  assign n24780 = pi119  & n9096;
  assign n24781 = pi117  & n9453;
  assign n24782 = pi118  & n9091;
  assign n24783 = ~n24781 & ~n24782;
  assign n24784 = ~n24780 & n24783;
  assign n24785 = n9099 & n10048;
  assign n24786 = n24784 & ~n24785;
  assign n24787 = pi53  & ~n24786;
  assign n24788 = pi53  & ~n24787;
  assign n24789 = ~n24786 & ~n24787;
  assign n24790 = ~n24788 & ~n24789;
  assign n24791 = n24779 & ~n24790;
  assign n24792 = ~n24779 & n24790;
  assign n24793 = ~n24791 & ~n24792;
  assign n24794 = ~n24718 & n24793;
  assign n24795 = n24718 & ~n24793;
  assign n24796 = ~n24794 & ~n24795;
  assign n24797 = n24717 & ~n24796;
  assign n24798 = ~n24717 & n24796;
  assign n24799 = ~n24797 & ~n24798;
  assign n24800 = ~n24706 & n24799;
  assign n24801 = n24706 & ~n24799;
  assign n24802 = ~n24800 & ~n24801;
  assign n24803 = ~n24705 & n24802;
  assign n24804 = ~n24705 & ~n24803;
  assign n24805 = n24802 & ~n24803;
  assign n24806 = ~n24804 & ~n24805;
  assign n24807 = n24694 & ~n24806;
  assign n24808 = ~n24694 & n24806;
  assign n24809 = ~n24807 & ~n24808;
  assign n24810 = n24681 & ~n24809;
  assign n24811 = ~n24681 & n24809;
  assign n24812 = ~n24810 & ~n24811;
  assign n24813 = ~n24675 & ~n24678;
  assign n24814 = n24812 & ~n24813;
  assign n24815 = ~n24812 & n24813;
  assign po106  = ~n24814 & ~n24815;
  assign n24817 = ~n24811 & ~n24814;
  assign n24818 = ~n24692 & ~n24807;
  assign n24819 = ~n24794 & ~n24798;
  assign n24820 = ~n24778 & ~n24791;
  assign n24821 = pi120  & n9096;
  assign n24822 = pi118  & n9453;
  assign n24823 = pi119  & n9091;
  assign n24824 = ~n24822 & ~n24823;
  assign n24825 = ~n24821 & n24824;
  assign n24826 = n9099 & n10734;
  assign n24827 = n24825 & ~n24826;
  assign n24828 = pi53  & ~n24827;
  assign n24829 = pi53  & ~n24828;
  assign n24830 = ~n24827 & ~n24828;
  assign n24831 = ~n24829 & ~n24830;
  assign n24832 = ~n24761 & ~n24774;
  assign n24833 = pi117  & n10135;
  assign n24834 = pi115  & n10478;
  assign n24835 = pi116  & n10130;
  assign n24836 = ~n24834 & ~n24835;
  assign n24837 = ~n24833 & n24836;
  assign n24838 = n9691 & n10138;
  assign n24839 = n24837 & ~n24838;
  assign n24840 = pi56  & ~n24839;
  assign n24841 = pi56  & ~n24840;
  assign n24842 = ~n24839 & ~n24840;
  assign n24843 = ~n24841 & ~n24842;
  assign n24844 = ~n24743 & ~n24757;
  assign n24845 = pi114  & n11193;
  assign n24846 = pi112  & n11567;
  assign n24847 = pi113  & n11188;
  assign n24848 = ~n24846 & ~n24847;
  assign n24849 = ~n24845 & n24848;
  assign n24850 = n8702 & n11196;
  assign n24851 = n24849 & ~n24850;
  assign n24852 = pi59  & ~n24851;
  assign n24853 = pi59  & ~n24852;
  assign n24854 = ~n24851 & ~n24852;
  assign n24855 = ~n24853 & ~n24854;
  assign n24856 = ~n24737 & ~n24740;
  assign n24857 = pi107  & n13477;
  assign n24858 = pi108  & ~n13122;
  assign n24859 = ~n24857 & ~n24858;
  assign n24860 = n24735 & ~n24859;
  assign n24861 = ~n24735 & n24859;
  assign n24862 = ~n24860 & ~n24861;
  assign n24863 = pi111  & n12295;
  assign n24864 = pi109  & n12693;
  assign n24865 = pi110  & n12290;
  assign n24866 = ~n24864 & ~n24865;
  assign n24867 = ~n24863 & n24866;
  assign n24868 = ~n12298 & n24867;
  assign n24869 = ~n7770 & n24867;
  assign n24870 = ~n24868 & ~n24869;
  assign n24871 = pi62  & ~n24870;
  assign n24872 = ~pi62  & n24870;
  assign n24873 = ~n24871 & ~n24872;
  assign n24874 = n24862 & ~n24873;
  assign n24875 = ~n24862 & n24873;
  assign n24876 = ~n24874 & ~n24875;
  assign n24877 = ~n24856 & n24876;
  assign n24878 = ~n24856 & ~n24877;
  assign n24879 = n24876 & ~n24877;
  assign n24880 = ~n24878 & ~n24879;
  assign n24881 = ~n24855 & ~n24880;
  assign n24882 = n24855 & n24880;
  assign n24883 = ~n24881 & ~n24882;
  assign n24884 = ~n24844 & n24883;
  assign n24885 = n24844 & ~n24883;
  assign n24886 = ~n24884 & ~n24885;
  assign n24887 = ~n24843 & n24886;
  assign n24888 = n24843 & ~n24886;
  assign n24889 = ~n24887 & ~n24888;
  assign n24890 = ~n24832 & n24889;
  assign n24891 = n24832 & ~n24889;
  assign n24892 = ~n24890 & ~n24891;
  assign n24893 = ~n24831 & n24892;
  assign n24894 = n24831 & ~n24892;
  assign n24895 = ~n24893 & ~n24894;
  assign n24896 = ~n24820 & n24895;
  assign n24897 = n24820 & ~n24895;
  assign n24898 = ~n24896 & ~n24897;
  assign n24899 = pi123  & n8137;
  assign n24900 = pi121  & n8471;
  assign n24901 = pi122  & n8132;
  assign n24902 = ~n24900 & ~n24901;
  assign n24903 = ~n24899 & n24902;
  assign n24904 = n8140 & n11489;
  assign n24905 = n24903 & ~n24904;
  assign n24906 = pi50  & ~n24905;
  assign n24907 = pi50  & ~n24906;
  assign n24908 = ~n24905 & ~n24906;
  assign n24909 = ~n24907 & ~n24908;
  assign n24910 = n24898 & ~n24909;
  assign n24911 = ~n24898 & n24909;
  assign n24912 = ~n24910 & ~n24911;
  assign n24913 = ~n24819 & n24912;
  assign n24914 = n24819 & ~n24912;
  assign n24915 = ~n24913 & ~n24914;
  assign n24916 = pi126  & n7239;
  assign n24917 = pi124  & n7556;
  assign n24918 = pi125  & n7234;
  assign n24919 = ~n24917 & ~n24918;
  assign n24920 = ~n24916 & n24919;
  assign n24921 = n7242 & n12979;
  assign n24922 = n24920 & ~n24921;
  assign n24923 = pi47  & ~n24922;
  assign n24924 = pi47  & ~n24923;
  assign n24925 = ~n24922 & ~n24923;
  assign n24926 = ~n24924 & ~n24925;
  assign n24927 = n24915 & ~n24926;
  assign n24928 = n24915 & ~n24927;
  assign n24929 = ~n24926 & ~n24927;
  assign n24930 = ~n24928 & ~n24929;
  assign n24931 = ~n24800 & ~n24803;
  assign n24932 = pi127  & n6735;
  assign n24933 = n6399 & n13387;
  assign n24934 = ~n24932 & ~n24933;
  assign n24935 = pi44  & ~n24934;
  assign n24936 = pi44  & ~n24935;
  assign n24937 = ~n24934 & ~n24935;
  assign n24938 = ~n24936 & ~n24937;
  assign n24939 = ~n24931 & ~n24938;
  assign n24940 = n24931 & n24938;
  assign n24941 = ~n24939 & ~n24940;
  assign n24942 = n24930 & n24941;
  assign n24943 = ~n24930 & ~n24941;
  assign n24944 = ~n24942 & ~n24943;
  assign n24945 = ~n24818 & ~n24944;
  assign n24946 = n24818 & n24944;
  assign n24947 = ~n24945 & ~n24946;
  assign n24948 = ~n24817 & n24947;
  assign n24949 = n24817 & ~n24947;
  assign po107  = ~n24948 & ~n24949;
  assign n24951 = ~n24945 & ~n24948;
  assign n24952 = ~n24896 & ~n24910;
  assign n24953 = pi124  & n8137;
  assign n24954 = pi122  & n8471;
  assign n24955 = pi123  & n8132;
  assign n24956 = ~n24954 & ~n24955;
  assign n24957 = ~n24953 & n24956;
  assign n24958 = n8140 & n11858;
  assign n24959 = n24957 & ~n24958;
  assign n24960 = pi50  & ~n24959;
  assign n24961 = pi50  & ~n24960;
  assign n24962 = ~n24959 & ~n24960;
  assign n24963 = ~n24961 & ~n24962;
  assign n24964 = ~n24890 & ~n24893;
  assign n24965 = pi121  & n9096;
  assign n24966 = pi119  & n9453;
  assign n24967 = pi120  & n9091;
  assign n24968 = ~n24966 & ~n24967;
  assign n24969 = ~n24965 & n24968;
  assign n24970 = n9099 & n11086;
  assign n24971 = n24969 & ~n24970;
  assign n24972 = pi53  & ~n24971;
  assign n24973 = pi53  & ~n24972;
  assign n24974 = ~n24971 & ~n24972;
  assign n24975 = ~n24973 & ~n24974;
  assign n24976 = ~n24884 & ~n24887;
  assign n24977 = pi118  & n10135;
  assign n24978 = pi116  & n10478;
  assign n24979 = pi117  & n10130;
  assign n24980 = ~n24978 & ~n24979;
  assign n24981 = ~n24977 & n24980;
  assign n24982 = n9716 & n10138;
  assign n24983 = n24981 & ~n24982;
  assign n24984 = pi56  & ~n24983;
  assign n24985 = pi56  & ~n24984;
  assign n24986 = ~n24983 & ~n24984;
  assign n24987 = ~n24985 & ~n24986;
  assign n24988 = ~n24877 & ~n24881;
  assign n24989 = ~n24860 & ~n24874;
  assign n24990 = pi108  & n13477;
  assign n24991 = pi109  & ~n13122;
  assign n24992 = ~n24990 & ~n24991;
  assign n24993 = ~pi44  & ~n24992;
  assign n24994 = pi44  & n24992;
  assign n24995 = ~n24993 & ~n24994;
  assign n24996 = ~n24735 & n24995;
  assign n24997 = n24735 & ~n24995;
  assign n24998 = ~n24996 & ~n24997;
  assign n24999 = ~n24989 & n24998;
  assign n25000 = n24989 & ~n24998;
  assign n25001 = ~n24999 & ~n25000;
  assign n25002 = pi112  & n12295;
  assign n25003 = pi110  & n12693;
  assign n25004 = pi111  & n12290;
  assign n25005 = ~n25003 & ~n25004;
  assign n25006 = ~n25002 & n25005;
  assign n25007 = n7795 & n12298;
  assign n25008 = n25006 & ~n25007;
  assign n25009 = pi62  & ~n25008;
  assign n25010 = pi62  & ~n25009;
  assign n25011 = ~n25008 & ~n25009;
  assign n25012 = ~n25010 & ~n25011;
  assign n25013 = n25001 & ~n25012;
  assign n25014 = n25001 & ~n25013;
  assign n25015 = ~n25012 & ~n25013;
  assign n25016 = ~n25014 & ~n25015;
  assign n25017 = pi115  & n11193;
  assign n25018 = pi113  & n11567;
  assign n25019 = pi114  & n11188;
  assign n25020 = ~n25018 & ~n25019;
  assign n25021 = ~n25017 & n25020;
  assign n25022 = n8727 & n11196;
  assign n25023 = n25021 & ~n25022;
  assign n25024 = pi59  & ~n25023;
  assign n25025 = pi59  & ~n25024;
  assign n25026 = ~n25023 & ~n25024;
  assign n25027 = ~n25025 & ~n25026;
  assign n25028 = n25016 & n25027;
  assign n25029 = ~n25016 & ~n25027;
  assign n25030 = ~n25028 & ~n25029;
  assign n25031 = ~n24988 & n25030;
  assign n25032 = n24988 & ~n25030;
  assign n25033 = ~n25031 & ~n25032;
  assign n25034 = n24987 & ~n25033;
  assign n25035 = ~n24987 & n25033;
  assign n25036 = ~n25034 & ~n25035;
  assign n25037 = ~n24976 & n25036;
  assign n25038 = n24976 & ~n25036;
  assign n25039 = ~n25037 & ~n25038;
  assign n25040 = n24975 & ~n25039;
  assign n25041 = ~n24975 & n25039;
  assign n25042 = ~n25040 & ~n25041;
  assign n25043 = ~n24964 & n25042;
  assign n25044 = n24964 & ~n25042;
  assign n25045 = ~n25043 & ~n25044;
  assign n25046 = n24963 & ~n25045;
  assign n25047 = ~n24963 & n25045;
  assign n25048 = ~n25046 & ~n25047;
  assign n25049 = ~n24952 & n25048;
  assign n25050 = n24952 & ~n25048;
  assign n25051 = ~n25049 & ~n25050;
  assign n25052 = pi127  & n7239;
  assign n25053 = pi125  & n7556;
  assign n25054 = pi126  & n7234;
  assign n25055 = ~n25053 & ~n25054;
  assign n25056 = ~n25052 & n25055;
  assign n25057 = n7242 & n13365;
  assign n25058 = n25056 & ~n25057;
  assign n25059 = pi47  & ~n25058;
  assign n25060 = pi47  & ~n25059;
  assign n25061 = ~n25058 & ~n25059;
  assign n25062 = ~n25060 & ~n25061;
  assign n25063 = n25051 & ~n25062;
  assign n25064 = n25051 & ~n25063;
  assign n25065 = ~n25062 & ~n25063;
  assign n25066 = ~n25064 & ~n25065;
  assign n25067 = ~n24913 & ~n24927;
  assign n25068 = n25066 & n25067;
  assign n25069 = ~n25066 & ~n25067;
  assign n25070 = ~n25068 & ~n25069;
  assign n25071 = ~n24940 & ~n24942;
  assign n25072 = n25070 & n25071;
  assign n25073 = ~n25070 & ~n25071;
  assign n25074 = ~n25072 & ~n25073;
  assign n25075 = ~n24951 & n25074;
  assign n25076 = n24951 & ~n25074;
  assign po108  = ~n25075 & ~n25076;
  assign n25078 = ~n25063 & ~n25069;
  assign n25079 = ~n25047 & ~n25049;
  assign n25080 = pi126  & n7556;
  assign n25081 = pi127  & n7234;
  assign n25082 = ~n25080 & ~n25081;
  assign n25083 = ~n7242 & n25082;
  assign n25084 = ~n13389 & n25082;
  assign n25085 = ~n25083 & ~n25084;
  assign n25086 = pi47  & ~n25085;
  assign n25087 = ~pi47  & n25085;
  assign n25088 = ~n25086 & ~n25087;
  assign n25089 = ~n25079 & ~n25088;
  assign n25090 = n25079 & n25088;
  assign n25091 = ~n25089 & ~n25090;
  assign n25092 = pi125  & n8137;
  assign n25093 = pi123  & n8471;
  assign n25094 = pi124  & n8132;
  assign n25095 = ~n25093 & ~n25094;
  assign n25096 = ~n25092 & n25095;
  assign n25097 = n8140 & n12591;
  assign n25098 = n25096 & ~n25097;
  assign n25099 = pi50  & ~n25098;
  assign n25100 = pi50  & ~n25099;
  assign n25101 = ~n25098 & ~n25099;
  assign n25102 = ~n25100 & ~n25101;
  assign n25103 = ~n25041 & ~n25043;
  assign n25104 = pi122  & n9096;
  assign n25105 = pi120  & n9453;
  assign n25106 = pi121  & n9091;
  assign n25107 = ~n25105 & ~n25106;
  assign n25108 = ~n25104 & n25107;
  assign n25109 = n9099 & n11463;
  assign n25110 = n25108 & ~n25109;
  assign n25111 = pi53  & ~n25110;
  assign n25112 = pi53  & ~n25111;
  assign n25113 = ~n25110 & ~n25111;
  assign n25114 = ~n25112 & ~n25113;
  assign n25115 = ~n25035 & ~n25037;
  assign n25116 = ~n25029 & ~n25031;
  assign n25117 = pi116  & n11193;
  assign n25118 = pi114  & n11567;
  assign n25119 = pi115  & n11188;
  assign n25120 = ~n25118 & ~n25119;
  assign n25121 = ~n25117 & n25120;
  assign n25122 = n9042 & n11196;
  assign n25123 = n25121 & ~n25122;
  assign n25124 = pi59  & ~n25123;
  assign n25125 = pi59  & ~n25124;
  assign n25126 = ~n25123 & ~n25124;
  assign n25127 = ~n25125 & ~n25126;
  assign n25128 = ~n24999 & ~n25013;
  assign n25129 = pi109  & n13477;
  assign n25130 = pi110  & ~n13122;
  assign n25131 = ~n25129 & ~n25130;
  assign n25132 = ~n24993 & ~n24996;
  assign n25133 = ~n25131 & n25132;
  assign n25134 = n25131 & ~n25132;
  assign n25135 = ~n25133 & ~n25134;
  assign n25136 = pi113  & n12295;
  assign n25137 = pi111  & n12693;
  assign n25138 = pi112  & n12290;
  assign n25139 = ~n25137 & ~n25138;
  assign n25140 = ~n25136 & n25139;
  assign n25141 = n8387 & n12298;
  assign n25142 = n25140 & ~n25141;
  assign n25143 = pi62  & ~n25142;
  assign n25144 = pi62  & ~n25143;
  assign n25145 = ~n25142 & ~n25143;
  assign n25146 = ~n25144 & ~n25145;
  assign n25147 = ~n25135 & n25146;
  assign n25148 = n25135 & ~n25146;
  assign n25149 = ~n25147 & ~n25148;
  assign n25150 = ~n25128 & n25149;
  assign n25151 = n25128 & ~n25149;
  assign n25152 = ~n25150 & ~n25151;
  assign n25153 = ~n25127 & n25152;
  assign n25154 = n25127 & ~n25152;
  assign n25155 = ~n25153 & ~n25154;
  assign n25156 = ~n25116 & n25155;
  assign n25157 = n25116 & ~n25155;
  assign n25158 = ~n25156 & ~n25157;
  assign n25159 = pi119  & n10135;
  assign n25160 = pi117  & n10478;
  assign n25161 = pi118  & n10130;
  assign n25162 = ~n25160 & ~n25161;
  assign n25163 = ~n25159 & n25162;
  assign n25164 = n10048 & n10138;
  assign n25165 = n25163 & ~n25164;
  assign n25166 = pi56  & ~n25165;
  assign n25167 = pi56  & ~n25166;
  assign n25168 = ~n25165 & ~n25166;
  assign n25169 = ~n25167 & ~n25168;
  assign n25170 = n25158 & ~n25169;
  assign n25171 = ~n25158 & n25169;
  assign n25172 = ~n25170 & ~n25171;
  assign n25173 = ~n25115 & n25172;
  assign n25174 = n25115 & ~n25172;
  assign n25175 = ~n25173 & ~n25174;
  assign n25176 = n25114 & ~n25175;
  assign n25177 = ~n25114 & n25175;
  assign n25178 = ~n25176 & ~n25177;
  assign n25179 = ~n25103 & n25178;
  assign n25180 = n25103 & ~n25178;
  assign n25181 = ~n25179 & ~n25180;
  assign n25182 = ~n25102 & n25181;
  assign n25183 = ~n25102 & ~n25182;
  assign n25184 = n25181 & ~n25182;
  assign n25185 = ~n25183 & ~n25184;
  assign n25186 = n25091 & ~n25185;
  assign n25187 = ~n25091 & n25185;
  assign n25188 = ~n25186 & ~n25187;
  assign n25189 = n25078 & ~n25188;
  assign n25190 = ~n25078 & n25188;
  assign n25191 = ~n25189 & ~n25190;
  assign n25192 = ~n25072 & ~n25075;
  assign n25193 = n25191 & ~n25192;
  assign n25194 = ~n25191 & n25192;
  assign po109  = ~n25193 & ~n25194;
  assign n25196 = ~n25089 & ~n25186;
  assign n25197 = ~n25173 & ~n25177;
  assign n25198 = ~n25156 & ~n25170;
  assign n25199 = pi120  & n10135;
  assign n25200 = pi118  & n10478;
  assign n25201 = pi119  & n10130;
  assign n25202 = ~n25200 & ~n25201;
  assign n25203 = ~n25199 & n25202;
  assign n25204 = n10138 & n10734;
  assign n25205 = n25203 & ~n25204;
  assign n25206 = pi56  & ~n25205;
  assign n25207 = pi56  & ~n25206;
  assign n25208 = ~n25205 & ~n25206;
  assign n25209 = ~n25207 & ~n25208;
  assign n25210 = ~n25150 & ~n25153;
  assign n25211 = pi117  & n11193;
  assign n25212 = pi115  & n11567;
  assign n25213 = pi116  & n11188;
  assign n25214 = ~n25212 & ~n25213;
  assign n25215 = ~n25211 & n25214;
  assign n25216 = n9691 & n11196;
  assign n25217 = n25215 & ~n25216;
  assign n25218 = pi59  & ~n25217;
  assign n25219 = pi59  & ~n25218;
  assign n25220 = ~n25217 & ~n25218;
  assign n25221 = ~n25219 & ~n25220;
  assign n25222 = ~n25134 & ~n25148;
  assign n25223 = pi110  & n13477;
  assign n25224 = pi111  & ~n13122;
  assign n25225 = ~n25223 & ~n25224;
  assign n25226 = n25131 & ~n25225;
  assign n25227 = ~n25131 & n25225;
  assign n25228 = ~n25222 & ~n25227;
  assign n25229 = ~n25226 & n25228;
  assign n25230 = ~n25222 & ~n25229;
  assign n25231 = ~n25227 & ~n25229;
  assign n25232 = ~n25226 & n25231;
  assign n25233 = ~n25230 & ~n25232;
  assign n25234 = pi114  & n12295;
  assign n25235 = pi112  & n12693;
  assign n25236 = pi113  & n12290;
  assign n25237 = ~n25235 & ~n25236;
  assign n25238 = ~n25234 & n25237;
  assign n25239 = n8702 & n12298;
  assign n25240 = n25238 & ~n25239;
  assign n25241 = pi62  & ~n25240;
  assign n25242 = pi62  & ~n25241;
  assign n25243 = ~n25240 & ~n25241;
  assign n25244 = ~n25242 & ~n25243;
  assign n25245 = ~n25233 & ~n25244;
  assign n25246 = n25233 & n25244;
  assign n25247 = ~n25245 & ~n25246;
  assign n25248 = ~n25221 & n25247;
  assign n25249 = n25221 & ~n25247;
  assign n25250 = ~n25248 & ~n25249;
  assign n25251 = ~n25210 & n25250;
  assign n25252 = n25210 & ~n25250;
  assign n25253 = ~n25251 & ~n25252;
  assign n25254 = ~n25209 & n25253;
  assign n25255 = n25209 & ~n25253;
  assign n25256 = ~n25254 & ~n25255;
  assign n25257 = ~n25198 & n25256;
  assign n25258 = n25198 & ~n25256;
  assign n25259 = ~n25257 & ~n25258;
  assign n25260 = pi123  & n9096;
  assign n25261 = pi121  & n9453;
  assign n25262 = pi122  & n9091;
  assign n25263 = ~n25261 & ~n25262;
  assign n25264 = ~n25260 & n25263;
  assign n25265 = n9099 & n11489;
  assign n25266 = n25264 & ~n25265;
  assign n25267 = pi53  & ~n25266;
  assign n25268 = pi53  & ~n25267;
  assign n25269 = ~n25266 & ~n25267;
  assign n25270 = ~n25268 & ~n25269;
  assign n25271 = n25259 & ~n25270;
  assign n25272 = ~n25259 & n25270;
  assign n25273 = ~n25271 & ~n25272;
  assign n25274 = ~n25197 & n25273;
  assign n25275 = n25197 & ~n25273;
  assign n25276 = ~n25274 & ~n25275;
  assign n25277 = pi126  & n8137;
  assign n25278 = pi124  & n8471;
  assign n25279 = pi125  & n8132;
  assign n25280 = ~n25278 & ~n25279;
  assign n25281 = ~n25277 & n25280;
  assign n25282 = n8140 & n12979;
  assign n25283 = n25281 & ~n25282;
  assign n25284 = pi50  & ~n25283;
  assign n25285 = pi50  & ~n25284;
  assign n25286 = ~n25283 & ~n25284;
  assign n25287 = ~n25285 & ~n25286;
  assign n25288 = n25276 & ~n25287;
  assign n25289 = n25276 & ~n25288;
  assign n25290 = ~n25287 & ~n25288;
  assign n25291 = ~n25289 & ~n25290;
  assign n25292 = ~n25179 & ~n25182;
  assign n25293 = pi127  & n7556;
  assign n25294 = ~n7242 & ~n25293;
  assign n25295 = ~n13387 & ~n25293;
  assign n25296 = ~n25294 & ~n25295;
  assign n25297 = pi47  & ~n25296;
  assign n25298 = ~pi47  & n25296;
  assign n25299 = ~n25297 & ~n25298;
  assign n25300 = ~n25292 & ~n25299;
  assign n25301 = n25292 & n25299;
  assign n25302 = ~n25300 & ~n25301;
  assign n25303 = ~n25291 & n25302;
  assign n25304 = n25291 & ~n25302;
  assign n25305 = ~n25303 & ~n25304;
  assign n25306 = n25196 & ~n25305;
  assign n25307 = ~n25196 & n25305;
  assign n25308 = ~n25306 & ~n25307;
  assign n25309 = ~n25190 & ~n25193;
  assign n25310 = n25308 & ~n25309;
  assign n25311 = ~n25308 & n25309;
  assign po110  = ~n25310 & ~n25311;
  assign n25313 = ~n25257 & ~n25271;
  assign n25314 = pi124  & n9096;
  assign n25315 = pi122  & n9453;
  assign n25316 = pi123  & n9091;
  assign n25317 = ~n25315 & ~n25316;
  assign n25318 = ~n25314 & n25317;
  assign n25319 = n9099 & n11858;
  assign n25320 = n25318 & ~n25319;
  assign n25321 = pi53  & ~n25320;
  assign n25322 = pi53  & ~n25321;
  assign n25323 = ~n25320 & ~n25321;
  assign n25324 = ~n25322 & ~n25323;
  assign n25325 = ~n25251 & ~n25254;
  assign n25326 = pi121  & n10135;
  assign n25327 = pi119  & n10478;
  assign n25328 = pi120  & n10130;
  assign n25329 = ~n25327 & ~n25328;
  assign n25330 = ~n25326 & n25329;
  assign n25331 = n10138 & n11086;
  assign n25332 = n25330 & ~n25331;
  assign n25333 = pi56  & ~n25332;
  assign n25334 = pi56  & ~n25333;
  assign n25335 = ~n25332 & ~n25333;
  assign n25336 = ~n25334 & ~n25335;
  assign n25337 = ~n25245 & ~n25248;
  assign n25338 = pi118  & n11193;
  assign n25339 = pi116  & n11567;
  assign n25340 = pi117  & n11188;
  assign n25341 = ~n25339 & ~n25340;
  assign n25342 = ~n25338 & n25341;
  assign n25343 = n9716 & n11196;
  assign n25344 = n25342 & ~n25343;
  assign n25345 = pi59  & ~n25344;
  assign n25346 = pi59  & ~n25345;
  assign n25347 = ~n25344 & ~n25345;
  assign n25348 = ~n25346 & ~n25347;
  assign n25349 = pi115  & n12295;
  assign n25350 = pi113  & n12693;
  assign n25351 = pi114  & n12290;
  assign n25352 = ~n25350 & ~n25351;
  assign n25353 = ~n25349 & n25352;
  assign n25354 = n8727 & n12298;
  assign n25355 = n25353 & ~n25354;
  assign n25356 = pi62  & ~n25355;
  assign n25357 = pi62  & ~n25356;
  assign n25358 = ~n25355 & ~n25356;
  assign n25359 = ~n25357 & ~n25358;
  assign n25360 = pi111  & n13477;
  assign n25361 = pi112  & ~n13122;
  assign n25362 = ~n25360 & ~n25361;
  assign n25363 = ~pi47  & ~n25225;
  assign n25364 = pi47  & n25225;
  assign n25365 = ~n25363 & ~n25364;
  assign n25366 = ~n25362 & n25365;
  assign n25367 = n25362 & ~n25365;
  assign n25368 = ~n25366 & ~n25367;
  assign n25369 = ~n25359 & n25368;
  assign n25370 = n25359 & ~n25368;
  assign n25371 = ~n25369 & ~n25370;
  assign n25372 = ~n25231 & n25371;
  assign n25373 = n25231 & ~n25371;
  assign n25374 = ~n25372 & ~n25373;
  assign n25375 = n25348 & ~n25374;
  assign n25376 = ~n25348 & n25374;
  assign n25377 = ~n25375 & ~n25376;
  assign n25378 = ~n25337 & n25377;
  assign n25379 = n25337 & ~n25377;
  assign n25380 = ~n25378 & ~n25379;
  assign n25381 = n25336 & ~n25380;
  assign n25382 = ~n25336 & n25380;
  assign n25383 = ~n25381 & ~n25382;
  assign n25384 = ~n25325 & n25383;
  assign n25385 = n25325 & ~n25383;
  assign n25386 = ~n25384 & ~n25385;
  assign n25387 = n25324 & ~n25386;
  assign n25388 = ~n25324 & n25386;
  assign n25389 = ~n25387 & ~n25388;
  assign n25390 = ~n25313 & n25389;
  assign n25391 = n25313 & ~n25389;
  assign n25392 = ~n25390 & ~n25391;
  assign n25393 = pi127  & n8137;
  assign n25394 = pi125  & n8471;
  assign n25395 = pi126  & n8132;
  assign n25396 = ~n25394 & ~n25395;
  assign n25397 = ~n25393 & n25396;
  assign n25398 = n8140 & n13365;
  assign n25399 = n25397 & ~n25398;
  assign n25400 = pi50  & ~n25399;
  assign n25401 = pi50  & ~n25400;
  assign n25402 = ~n25399 & ~n25400;
  assign n25403 = ~n25401 & ~n25402;
  assign n25404 = n25392 & ~n25403;
  assign n25405 = n25392 & ~n25404;
  assign n25406 = ~n25403 & ~n25404;
  assign n25407 = ~n25405 & ~n25406;
  assign n25408 = ~n25274 & ~n25288;
  assign n25409 = n25407 & n25408;
  assign n25410 = ~n25407 & ~n25408;
  assign n25411 = ~n25409 & ~n25410;
  assign n25412 = ~n25300 & ~n25303;
  assign n25413 = ~n25411 & n25412;
  assign n25414 = n25411 & ~n25412;
  assign n25415 = ~n25413 & ~n25414;
  assign n25416 = ~n25307 & ~n25310;
  assign n25417 = n25415 & ~n25416;
  assign n25418 = ~n25415 & n25416;
  assign po111  = ~n25417 & ~n25418;
  assign n25420 = ~n25388 & ~n25390;
  assign n25421 = pi125  & n9096;
  assign n25422 = pi123  & n9453;
  assign n25423 = pi124  & n9091;
  assign n25424 = ~n25422 & ~n25423;
  assign n25425 = ~n25421 & n25424;
  assign n25426 = n9099 & n12591;
  assign n25427 = n25425 & ~n25426;
  assign n25428 = pi53  & ~n25427;
  assign n25429 = pi53  & ~n25428;
  assign n25430 = ~n25427 & ~n25428;
  assign n25431 = ~n25429 & ~n25430;
  assign n25432 = ~n25382 & ~n25384;
  assign n25433 = pi122  & n10135;
  assign n25434 = pi120  & n10478;
  assign n25435 = pi121  & n10130;
  assign n25436 = ~n25434 & ~n25435;
  assign n25437 = ~n25433 & n25436;
  assign n25438 = n10138 & n11463;
  assign n25439 = n25437 & ~n25438;
  assign n25440 = pi56  & ~n25439;
  assign n25441 = pi56  & ~n25440;
  assign n25442 = ~n25439 & ~n25440;
  assign n25443 = ~n25441 & ~n25442;
  assign n25444 = ~n25376 & ~n25378;
  assign n25445 = pi119  & n11193;
  assign n25446 = pi117  & n11567;
  assign n25447 = pi118  & n11188;
  assign n25448 = ~n25446 & ~n25447;
  assign n25449 = ~n25445 & n25448;
  assign n25450 = n10048 & n11196;
  assign n25451 = n25449 & ~n25450;
  assign n25452 = pi59  & ~n25451;
  assign n25453 = pi59  & ~n25452;
  assign n25454 = ~n25451 & ~n25452;
  assign n25455 = ~n25453 & ~n25454;
  assign n25456 = ~n25369 & ~n25372;
  assign n25457 = pi112  & n13477;
  assign n25458 = pi113  & ~n13122;
  assign n25459 = ~n25457 & ~n25458;
  assign n25460 = ~n25363 & ~n25366;
  assign n25461 = n25459 & ~n25460;
  assign n25462 = ~n25459 & n25460;
  assign n25463 = ~n25461 & ~n25462;
  assign n25464 = pi116  & n12295;
  assign n25465 = pi114  & n12693;
  assign n25466 = pi115  & n12290;
  assign n25467 = ~n25465 & ~n25466;
  assign n25468 = ~n25464 & n25467;
  assign n25469 = ~n12298 & n25468;
  assign n25470 = ~n9042 & n25468;
  assign n25471 = ~n25469 & ~n25470;
  assign n25472 = pi62  & ~n25471;
  assign n25473 = ~pi62  & n25471;
  assign n25474 = ~n25472 & ~n25473;
  assign n25475 = n25463 & ~n25474;
  assign n25476 = ~n25463 & n25474;
  assign n25477 = ~n25475 & ~n25476;
  assign n25478 = ~n25456 & n25477;
  assign n25479 = n25456 & ~n25477;
  assign n25480 = ~n25478 & ~n25479;
  assign n25481 = ~n25455 & n25480;
  assign n25482 = n25455 & ~n25480;
  assign n25483 = ~n25481 & ~n25482;
  assign n25484 = ~n25444 & n25483;
  assign n25485 = n25444 & ~n25483;
  assign n25486 = ~n25484 & ~n25485;
  assign n25487 = ~n25443 & n25486;
  assign n25488 = n25443 & ~n25486;
  assign n25489 = ~n25487 & ~n25488;
  assign n25490 = ~n25432 & n25489;
  assign n25491 = n25432 & ~n25489;
  assign n25492 = ~n25490 & ~n25491;
  assign n25493 = ~n25431 & n25492;
  assign n25494 = n25431 & ~n25492;
  assign n25495 = ~n25493 & ~n25494;
  assign n25496 = ~n25420 & n25495;
  assign n25497 = n25420 & ~n25495;
  assign n25498 = ~n25496 & ~n25497;
  assign n25499 = pi126  & n8471;
  assign n25500 = pi127  & n8132;
  assign n25501 = ~n25499 & ~n25500;
  assign n25502 = n8140 & n13389;
  assign n25503 = n25501 & ~n25502;
  assign n25504 = pi50  & ~n25503;
  assign n25505 = pi50  & ~n25504;
  assign n25506 = ~n25503 & ~n25504;
  assign n25507 = ~n25505 & ~n25506;
  assign n25508 = n25498 & ~n25507;
  assign n25509 = n25498 & ~n25508;
  assign n25510 = ~n25507 & ~n25508;
  assign n25511 = ~n25509 & ~n25510;
  assign n25512 = ~n25404 & ~n25410;
  assign n25513 = n25511 & n25512;
  assign n25514 = ~n25511 & ~n25512;
  assign n25515 = ~n25513 & ~n25514;
  assign n25516 = ~n25414 & ~n25417;
  assign n25517 = n25515 & ~n25516;
  assign n25518 = ~n25515 & n25516;
  assign po112  = ~n25517 & ~n25518;
  assign n25520 = ~n25496 & ~n25508;
  assign n25521 = ~n25490 & ~n25493;
  assign n25522 = pi127  & n8471;
  assign n25523 = ~n8140 & ~n25522;
  assign n25524 = ~n13387 & ~n25522;
  assign n25525 = ~n25523 & ~n25524;
  assign n25526 = pi50  & ~n25525;
  assign n25527 = ~pi50  & n25525;
  assign n25528 = ~n25526 & ~n25527;
  assign n25529 = ~n25521 & ~n25528;
  assign n25530 = n25521 & n25528;
  assign n25531 = ~n25529 & ~n25530;
  assign n25532 = ~n25478 & ~n25481;
  assign n25533 = ~n25461 & ~n25475;
  assign n25534 = pi117  & n12295;
  assign n25535 = pi115  & n12693;
  assign n25536 = pi116  & n12290;
  assign n25537 = ~n25535 & ~n25536;
  assign n25538 = ~n25534 & n25537;
  assign n25539 = n9691 & n12298;
  assign n25540 = n25538 & ~n25539;
  assign n25541 = pi62  & ~n25540;
  assign n25542 = pi62  & ~n25541;
  assign n25543 = ~n25540 & ~n25541;
  assign n25544 = ~n25542 & ~n25543;
  assign n25545 = pi113  & n13477;
  assign n25546 = pi114  & ~n13122;
  assign n25547 = ~n25545 & ~n25546;
  assign n25548 = n25459 & ~n25547;
  assign n25549 = ~n25459 & n25547;
  assign n25550 = ~n25548 & ~n25549;
  assign n25551 = ~n25544 & n25550;
  assign n25552 = n25544 & ~n25550;
  assign n25553 = ~n25551 & ~n25552;
  assign n25554 = n25533 & ~n25553;
  assign n25555 = ~n25533 & n25553;
  assign n25556 = ~n25554 & ~n25555;
  assign n25557 = pi120  & n11193;
  assign n25558 = pi118  & n11567;
  assign n25559 = pi119  & n11188;
  assign n25560 = ~n25558 & ~n25559;
  assign n25561 = ~n25557 & n25560;
  assign n25562 = n10734 & n11196;
  assign n25563 = n25561 & ~n25562;
  assign n25564 = pi59  & ~n25563;
  assign n25565 = pi59  & ~n25564;
  assign n25566 = ~n25563 & ~n25564;
  assign n25567 = ~n25565 & ~n25566;
  assign n25568 = ~n25556 & n25567;
  assign n25569 = n25556 & ~n25567;
  assign n25570 = ~n25568 & ~n25569;
  assign n25571 = ~n25532 & n25570;
  assign n25572 = n25532 & ~n25570;
  assign n25573 = ~n25571 & ~n25572;
  assign n25574 = pi123  & n10135;
  assign n25575 = pi121  & n10478;
  assign n25576 = pi122  & n10130;
  assign n25577 = ~n25575 & ~n25576;
  assign n25578 = ~n25574 & n25577;
  assign n25579 = n10138 & n11489;
  assign n25580 = n25578 & ~n25579;
  assign n25581 = pi56  & ~n25580;
  assign n25582 = pi56  & ~n25581;
  assign n25583 = ~n25580 & ~n25581;
  assign n25584 = ~n25582 & ~n25583;
  assign n25585 = n25573 & ~n25584;
  assign n25586 = n25573 & ~n25585;
  assign n25587 = ~n25584 & ~n25585;
  assign n25588 = ~n25586 & ~n25587;
  assign n25589 = ~n25484 & ~n25487;
  assign n25590 = n25588 & n25589;
  assign n25591 = ~n25588 & ~n25589;
  assign n25592 = ~n25590 & ~n25591;
  assign n25593 = pi126  & n9096;
  assign n25594 = pi124  & n9453;
  assign n25595 = pi125  & n9091;
  assign n25596 = ~n25594 & ~n25595;
  assign n25597 = ~n25593 & n25596;
  assign n25598 = n9099 & n12979;
  assign n25599 = n25597 & ~n25598;
  assign n25600 = pi53  & ~n25599;
  assign n25601 = pi53  & ~n25600;
  assign n25602 = ~n25599 & ~n25600;
  assign n25603 = ~n25601 & ~n25602;
  assign n25604 = n25592 & ~n25603;
  assign n25605 = ~n25592 & n25603;
  assign n25606 = ~n25604 & ~n25605;
  assign n25607 = n25531 & n25606;
  assign n25608 = ~n25531 & ~n25606;
  assign n25609 = ~n25607 & ~n25608;
  assign n25610 = n25520 & ~n25609;
  assign n25611 = ~n25520 & n25609;
  assign n25612 = ~n25610 & ~n25611;
  assign n25613 = ~n25514 & ~n25517;
  assign n25614 = n25612 & ~n25613;
  assign n25615 = ~n25612 & n25613;
  assign po113  = ~n25614 & ~n25615;
  assign n25617 = ~n25591 & ~n25604;
  assign n25618 = ~n25571 & ~n25585;
  assign n25619 = pi124  & n10135;
  assign n25620 = pi122  & n10478;
  assign n25621 = pi123  & n10130;
  assign n25622 = ~n25620 & ~n25621;
  assign n25623 = ~n25619 & n25622;
  assign n25624 = n10138 & n11858;
  assign n25625 = n25623 & ~n25624;
  assign n25626 = pi56  & ~n25625;
  assign n25627 = pi56  & ~n25626;
  assign n25628 = ~n25625 & ~n25626;
  assign n25629 = ~n25627 & ~n25628;
  assign n25630 = ~n25555 & ~n25569;
  assign n25631 = pi121  & n11193;
  assign n25632 = pi119  & n11567;
  assign n25633 = pi120  & n11188;
  assign n25634 = ~n25632 & ~n25633;
  assign n25635 = ~n25631 & n25634;
  assign n25636 = n11086 & n11196;
  assign n25637 = n25635 & ~n25636;
  assign n25638 = pi59  & ~n25637;
  assign n25639 = pi59  & ~n25638;
  assign n25640 = ~n25637 & ~n25638;
  assign n25641 = ~n25639 & ~n25640;
  assign n25642 = pi118  & n12295;
  assign n25643 = pi116  & n12693;
  assign n25644 = pi117  & n12290;
  assign n25645 = ~n25643 & ~n25644;
  assign n25646 = ~n25642 & n25645;
  assign n25647 = n9716 & n12298;
  assign n25648 = n25646 & ~n25647;
  assign n25649 = pi62  & ~n25648;
  assign n25650 = pi62  & ~n25649;
  assign n25651 = ~n25648 & ~n25649;
  assign n25652 = ~n25650 & ~n25651;
  assign n25653 = ~n25548 & ~n25551;
  assign n25654 = pi114  & n13477;
  assign n25655 = pi115  & ~n13122;
  assign n25656 = ~n25654 & ~n25655;
  assign n25657 = ~pi50  & ~n25656;
  assign n25658 = pi50  & n25656;
  assign n25659 = ~n25657 & ~n25658;
  assign n25660 = ~n25459 & n25659;
  assign n25661 = n25459 & ~n25659;
  assign n25662 = ~n25660 & ~n25661;
  assign n25663 = ~n25653 & n25662;
  assign n25664 = n25653 & ~n25662;
  assign n25665 = ~n25663 & ~n25664;
  assign n25666 = ~n25652 & n25665;
  assign n25667 = n25652 & ~n25665;
  assign n25668 = ~n25666 & ~n25667;
  assign n25669 = ~n25641 & n25668;
  assign n25670 = n25641 & ~n25668;
  assign n25671 = ~n25669 & ~n25670;
  assign n25672 = ~n25630 & n25671;
  assign n25673 = n25630 & ~n25671;
  assign n25674 = ~n25672 & ~n25673;
  assign n25675 = ~n25629 & n25674;
  assign n25676 = n25629 & ~n25674;
  assign n25677 = ~n25675 & ~n25676;
  assign n25678 = ~n25618 & n25677;
  assign n25679 = n25618 & ~n25677;
  assign n25680 = ~n25678 & ~n25679;
  assign n25681 = pi127  & n9096;
  assign n25682 = pi125  & n9453;
  assign n25683 = pi126  & n9091;
  assign n25684 = ~n25682 & ~n25683;
  assign n25685 = ~n25681 & n25684;
  assign n25686 = n9099 & n13365;
  assign n25687 = n25685 & ~n25686;
  assign n25688 = pi53  & ~n25687;
  assign n25689 = pi53  & ~n25688;
  assign n25690 = ~n25687 & ~n25688;
  assign n25691 = ~n25689 & ~n25690;
  assign n25692 = n25680 & ~n25691;
  assign n25693 = ~n25680 & n25691;
  assign n25694 = ~n25692 & ~n25693;
  assign n25695 = n25617 & ~n25694;
  assign n25696 = ~n25617 & n25694;
  assign n25697 = ~n25695 & ~n25696;
  assign n25698 = ~n25529 & ~n25607;
  assign n25699 = ~n25697 & n25698;
  assign n25700 = n25697 & ~n25698;
  assign n25701 = ~n25699 & ~n25700;
  assign n25702 = ~n25611 & ~n25614;
  assign n25703 = n25701 & ~n25702;
  assign n25704 = ~n25701 & n25702;
  assign po114  = ~n25703 & ~n25704;
  assign n25706 = ~n25692 & ~n25696;
  assign n25707 = ~n25675 & ~n25678;
  assign n25708 = pi125  & n10135;
  assign n25709 = pi123  & n10478;
  assign n25710 = pi124  & n10130;
  assign n25711 = ~n25709 & ~n25710;
  assign n25712 = ~n25708 & n25711;
  assign n25713 = n10138 & n12591;
  assign n25714 = n25712 & ~n25713;
  assign n25715 = pi56  & ~n25714;
  assign n25716 = pi56  & ~n25715;
  assign n25717 = ~n25714 & ~n25715;
  assign n25718 = ~n25716 & ~n25717;
  assign n25719 = ~n25669 & ~n25672;
  assign n25720 = pi122  & n11193;
  assign n25721 = pi120  & n11567;
  assign n25722 = pi121  & n11188;
  assign n25723 = ~n25721 & ~n25722;
  assign n25724 = ~n25720 & n25723;
  assign n25725 = n11196 & n11463;
  assign n25726 = n25724 & ~n25725;
  assign n25727 = pi59  & ~n25726;
  assign n25728 = pi59  & ~n25727;
  assign n25729 = ~n25726 & ~n25727;
  assign n25730 = ~n25728 & ~n25729;
  assign n25731 = ~n25663 & ~n25666;
  assign n25732 = pi115  & n13477;
  assign n25733 = pi116  & ~n13122;
  assign n25734 = ~n25732 & ~n25733;
  assign n25735 = ~n25657 & ~n25660;
  assign n25736 = ~n25734 & n25735;
  assign n25737 = n25734 & ~n25735;
  assign n25738 = ~n25736 & ~n25737;
  assign n25739 = pi119  & n12295;
  assign n25740 = pi117  & n12693;
  assign n25741 = pi118  & n12290;
  assign n25742 = ~n25740 & ~n25741;
  assign n25743 = ~n25739 & n25742;
  assign n25744 = n10048 & n12298;
  assign n25745 = n25743 & ~n25744;
  assign n25746 = pi62  & ~n25745;
  assign n25747 = pi62  & ~n25746;
  assign n25748 = ~n25745 & ~n25746;
  assign n25749 = ~n25747 & ~n25748;
  assign n25750 = ~n25738 & n25749;
  assign n25751 = n25738 & ~n25749;
  assign n25752 = ~n25750 & ~n25751;
  assign n25753 = ~n25731 & n25752;
  assign n25754 = n25731 & ~n25752;
  assign n25755 = ~n25753 & ~n25754;
  assign n25756 = ~n25730 & n25755;
  assign n25757 = n25730 & ~n25755;
  assign n25758 = ~n25756 & ~n25757;
  assign n25759 = ~n25719 & n25758;
  assign n25760 = ~n25719 & ~n25759;
  assign n25761 = n25758 & ~n25759;
  assign n25762 = ~n25760 & ~n25761;
  assign n25763 = ~n25718 & ~n25762;
  assign n25764 = n25718 & n25762;
  assign n25765 = ~n25763 & ~n25764;
  assign n25766 = ~n25707 & n25765;
  assign n25767 = n25707 & ~n25765;
  assign n25768 = ~n25766 & ~n25767;
  assign n25769 = pi126  & n9453;
  assign n25770 = pi127  & n9091;
  assign n25771 = ~n25769 & ~n25770;
  assign n25772 = n9099 & n13389;
  assign n25773 = n25771 & ~n25772;
  assign n25774 = pi53  & ~n25773;
  assign n25775 = pi53  & ~n25774;
  assign n25776 = ~n25773 & ~n25774;
  assign n25777 = ~n25775 & ~n25776;
  assign n25778 = n25768 & ~n25777;
  assign n25779 = ~n25768 & n25777;
  assign n25780 = ~n25778 & ~n25779;
  assign n25781 = n25706 & ~n25780;
  assign n25782 = ~n25706 & n25780;
  assign n25783 = ~n25781 & ~n25782;
  assign n25784 = ~n25700 & ~n25703;
  assign n25785 = n25783 & ~n25784;
  assign n25786 = ~n25783 & n25784;
  assign po115  = ~n25785 & ~n25786;
  assign n25788 = ~n25766 & ~n25778;
  assign n25789 = ~n25759 & ~n25763;
  assign n25790 = pi127  & n9453;
  assign n25791 = ~n9099 & ~n25790;
  assign n25792 = ~n13387 & ~n25790;
  assign n25793 = ~n25791 & ~n25792;
  assign n25794 = pi53  & ~n25793;
  assign n25795 = ~pi53  & n25793;
  assign n25796 = ~n25794 & ~n25795;
  assign n25797 = ~n25789 & ~n25796;
  assign n25798 = n25789 & n25796;
  assign n25799 = ~n25797 & ~n25798;
  assign n25800 = ~n25753 & ~n25756;
  assign n25801 = pi123  & n11193;
  assign n25802 = pi121  & n11567;
  assign n25803 = pi122  & n11188;
  assign n25804 = ~n25802 & ~n25803;
  assign n25805 = ~n25801 & n25804;
  assign n25806 = n11196 & n11489;
  assign n25807 = n25805 & ~n25806;
  assign n25808 = pi59  & ~n25807;
  assign n25809 = pi59  & ~n25808;
  assign n25810 = ~n25807 & ~n25808;
  assign n25811 = ~n25809 & ~n25810;
  assign n25812 = ~n25737 & ~n25751;
  assign n25813 = pi116  & n13477;
  assign n25814 = pi117  & ~n13122;
  assign n25815 = ~n25813 & ~n25814;
  assign n25816 = n25734 & ~n25815;
  assign n25817 = ~n25734 & n25815;
  assign n25818 = ~n25812 & ~n25817;
  assign n25819 = ~n25816 & n25818;
  assign n25820 = ~n25812 & ~n25819;
  assign n25821 = ~n25817 & ~n25819;
  assign n25822 = ~n25816 & n25821;
  assign n25823 = ~n25820 & ~n25822;
  assign n25824 = pi120  & n12295;
  assign n25825 = pi118  & n12693;
  assign n25826 = pi119  & n12290;
  assign n25827 = ~n25825 & ~n25826;
  assign n25828 = ~n25824 & n25827;
  assign n25829 = n10734 & n12298;
  assign n25830 = n25828 & ~n25829;
  assign n25831 = pi62  & ~n25830;
  assign n25832 = pi62  & ~n25831;
  assign n25833 = ~n25830 & ~n25831;
  assign n25834 = ~n25832 & ~n25833;
  assign n25835 = ~n25823 & ~n25834;
  assign n25836 = n25823 & n25834;
  assign n25837 = ~n25835 & ~n25836;
  assign n25838 = ~n25811 & n25837;
  assign n25839 = n25811 & ~n25837;
  assign n25840 = ~n25838 & ~n25839;
  assign n25841 = n25800 & ~n25840;
  assign n25842 = ~n25800 & n25840;
  assign n25843 = ~n25841 & ~n25842;
  assign n25844 = pi126  & n10135;
  assign n25845 = pi124  & n10478;
  assign n25846 = pi125  & n10130;
  assign n25847 = ~n25845 & ~n25846;
  assign n25848 = ~n25844 & n25847;
  assign n25849 = n10138 & n12979;
  assign n25850 = n25848 & ~n25849;
  assign n25851 = pi56  & ~n25850;
  assign n25852 = pi56  & ~n25851;
  assign n25853 = ~n25850 & ~n25851;
  assign n25854 = ~n25852 & ~n25853;
  assign n25855 = n25843 & ~n25854;
  assign n25856 = ~n25843 & n25854;
  assign n25857 = ~n25855 & ~n25856;
  assign n25858 = n25799 & n25857;
  assign n25859 = ~n25799 & ~n25857;
  assign n25860 = ~n25858 & ~n25859;
  assign n25861 = n25788 & ~n25860;
  assign n25862 = ~n25788 & n25860;
  assign n25863 = ~n25861 & ~n25862;
  assign n25864 = ~n25782 & ~n25785;
  assign n25865 = n25863 & ~n25864;
  assign n25866 = ~n25863 & n25864;
  assign po116  = ~n25865 & ~n25866;
  assign n25868 = ~n25862 & ~n25865;
  assign n25869 = ~n25797 & ~n25858;
  assign n25870 = ~n25842 & ~n25855;
  assign n25871 = pi127  & n10135;
  assign n25872 = pi125  & n10478;
  assign n25873 = pi126  & n10130;
  assign n25874 = ~n25872 & ~n25873;
  assign n25875 = ~n25871 & n25874;
  assign n25876 = n10138 & n13365;
  assign n25877 = n25875 & ~n25876;
  assign n25878 = pi56  & ~n25877;
  assign n25879 = pi56  & ~n25878;
  assign n25880 = ~n25877 & ~n25878;
  assign n25881 = ~n25879 & ~n25880;
  assign n25882 = ~n25870 & ~n25881;
  assign n25883 = ~n25870 & ~n25882;
  assign n25884 = ~n25881 & ~n25882;
  assign n25885 = ~n25883 & ~n25884;
  assign n25886 = ~n25835 & ~n25838;
  assign n25887 = pi124  & n11193;
  assign n25888 = pi122  & n11567;
  assign n25889 = pi123  & n11188;
  assign n25890 = ~n25888 & ~n25889;
  assign n25891 = ~n25887 & n25890;
  assign n25892 = n11196 & n11858;
  assign n25893 = n25891 & ~n25892;
  assign n25894 = pi59  & ~n25893;
  assign n25895 = pi59  & ~n25894;
  assign n25896 = ~n25893 & ~n25894;
  assign n25897 = ~n25895 & ~n25896;
  assign n25898 = pi117  & n13477;
  assign n25899 = pi118  & ~n13122;
  assign n25900 = ~n25898 & ~n25899;
  assign n25901 = ~pi53  & ~n25815;
  assign n25902 = pi53  & n25815;
  assign n25903 = ~n25901 & ~n25902;
  assign n25904 = n25900 & ~n25903;
  assign n25905 = ~n25900 & n25903;
  assign n25906 = ~n25904 & ~n25905;
  assign n25907 = pi121  & n12295;
  assign n25908 = pi119  & n12693;
  assign n25909 = pi120  & n12290;
  assign n25910 = ~n25908 & ~n25909;
  assign n25911 = ~n25907 & n25910;
  assign n25912 = n11086 & n12298;
  assign n25913 = n25911 & ~n25912;
  assign n25914 = pi62  & ~n25913;
  assign n25915 = pi62  & ~n25914;
  assign n25916 = ~n25913 & ~n25914;
  assign n25917 = ~n25915 & ~n25916;
  assign n25918 = n25906 & ~n25917;
  assign n25919 = ~n25906 & n25917;
  assign n25920 = ~n25918 & ~n25919;
  assign n25921 = ~n25821 & n25920;
  assign n25922 = n25821 & ~n25920;
  assign n25923 = ~n25921 & ~n25922;
  assign n25924 = ~n25897 & n25923;
  assign n25925 = n25897 & ~n25923;
  assign n25926 = ~n25924 & ~n25925;
  assign n25927 = ~n25886 & n25926;
  assign n25928 = n25886 & ~n25926;
  assign n25929 = ~n25927 & ~n25928;
  assign n25930 = ~n25885 & n25929;
  assign n25931 = n25885 & ~n25929;
  assign n25932 = ~n25930 & ~n25931;
  assign n25933 = ~n25869 & n25932;
  assign n25934 = n25869 & ~n25932;
  assign n25935 = ~n25933 & ~n25934;
  assign n25936 = ~n25868 & n25935;
  assign n25937 = n25868 & ~n25935;
  assign po117  = ~n25936 & ~n25937;
  assign n25939 = ~n25933 & ~n25936;
  assign n25940 = ~n25882 & ~n25930;
  assign n25941 = ~n25924 & ~n25927;
  assign n25942 = pi125  & n11193;
  assign n25943 = pi123  & n11567;
  assign n25944 = pi124  & n11188;
  assign n25945 = ~n25943 & ~n25944;
  assign n25946 = ~n25942 & n25945;
  assign n25947 = n11196 & n12591;
  assign n25948 = n25946 & ~n25947;
  assign n25949 = pi59  & ~n25948;
  assign n25950 = pi59  & ~n25949;
  assign n25951 = ~n25948 & ~n25949;
  assign n25952 = ~n25950 & ~n25951;
  assign n25953 = ~n25918 & ~n25921;
  assign n25954 = pi118  & n13477;
  assign n25955 = pi119  & ~n13122;
  assign n25956 = ~n25954 & ~n25955;
  assign n25957 = ~n25901 & ~n25905;
  assign n25958 = n25956 & ~n25957;
  assign n25959 = ~n25956 & n25957;
  assign n25960 = ~n25958 & ~n25959;
  assign n25961 = pi122  & n12295;
  assign n25962 = pi120  & n12693;
  assign n25963 = pi121  & n12290;
  assign n25964 = ~n25962 & ~n25963;
  assign n25965 = ~n25961 & n25964;
  assign n25966 = ~n12298 & n25965;
  assign n25967 = ~n11463 & n25965;
  assign n25968 = ~n25966 & ~n25967;
  assign n25969 = pi62  & ~n25968;
  assign n25970 = ~pi62  & n25968;
  assign n25971 = ~n25969 & ~n25970;
  assign n25972 = n25960 & ~n25971;
  assign n25973 = ~n25960 & n25971;
  assign n25974 = ~n25972 & ~n25973;
  assign n25975 = ~n25953 & n25974;
  assign n25976 = n25953 & ~n25974;
  assign n25977 = ~n25975 & ~n25976;
  assign n25978 = ~n25952 & n25977;
  assign n25979 = n25952 & ~n25977;
  assign n25980 = ~n25978 & ~n25979;
  assign n25981 = ~n25941 & n25980;
  assign n25982 = n25941 & ~n25980;
  assign n25983 = ~n25981 & ~n25982;
  assign n25984 = pi126  & n10478;
  assign n25985 = pi127  & n10130;
  assign n25986 = ~n25984 & ~n25985;
  assign n25987 = n10138 & n13389;
  assign n25988 = n25986 & ~n25987;
  assign n25989 = pi56  & ~n25988;
  assign n25990 = pi56  & ~n25989;
  assign n25991 = ~n25988 & ~n25989;
  assign n25992 = ~n25990 & ~n25991;
  assign n25993 = n25983 & ~n25992;
  assign n25994 = ~n25983 & n25992;
  assign n25995 = ~n25993 & ~n25994;
  assign n25996 = ~n25940 & n25995;
  assign n25997 = n25940 & ~n25995;
  assign n25998 = ~n25996 & ~n25997;
  assign n25999 = ~n25939 & n25998;
  assign n26000 = n25939 & ~n25998;
  assign po118  = ~n25999 & ~n26000;
  assign n26002 = ~n25981 & ~n25993;
  assign n26003 = ~n25975 & ~n25978;
  assign n26004 = pi127  & n10478;
  assign n26005 = ~n10138 & ~n26004;
  assign n26006 = ~n13387 & ~n26004;
  assign n26007 = ~n26005 & ~n26006;
  assign n26008 = pi56  & ~n26007;
  assign n26009 = ~pi56  & n26007;
  assign n26010 = ~n26008 & ~n26009;
  assign n26011 = ~n26003 & ~n26010;
  assign n26012 = n26003 & n26010;
  assign n26013 = ~n26011 & ~n26012;
  assign n26014 = ~n25958 & ~n25972;
  assign n26015 = pi123  & n12295;
  assign n26016 = pi121  & n12693;
  assign n26017 = pi122  & n12290;
  assign n26018 = ~n26016 & ~n26017;
  assign n26019 = ~n26015 & n26018;
  assign n26020 = n11489 & n12298;
  assign n26021 = n26019 & ~n26020;
  assign n26022 = pi62  & ~n26021;
  assign n26023 = pi62  & ~n26022;
  assign n26024 = ~n26021 & ~n26022;
  assign n26025 = ~n26023 & ~n26024;
  assign n26026 = pi119  & n13477;
  assign n26027 = pi120  & ~n13122;
  assign n26028 = ~n26026 & ~n26027;
  assign n26029 = n25956 & ~n26028;
  assign n26030 = ~n25956 & n26028;
  assign n26031 = ~n26029 & ~n26030;
  assign n26032 = ~n26025 & n26031;
  assign n26033 = n26025 & ~n26031;
  assign n26034 = ~n26032 & ~n26033;
  assign n26035 = n26014 & ~n26034;
  assign n26036 = ~n26014 & n26034;
  assign n26037 = ~n26035 & ~n26036;
  assign n26038 = pi126  & n11193;
  assign n26039 = pi124  & n11567;
  assign n26040 = pi125  & n11188;
  assign n26041 = ~n26039 & ~n26040;
  assign n26042 = ~n26038 & n26041;
  assign n26043 = n11196 & n12979;
  assign n26044 = n26042 & ~n26043;
  assign n26045 = pi59  & ~n26044;
  assign n26046 = pi59  & ~n26045;
  assign n26047 = ~n26044 & ~n26045;
  assign n26048 = ~n26046 & ~n26047;
  assign n26049 = n26037 & ~n26048;
  assign n26050 = ~n26037 & n26048;
  assign n26051 = ~n26049 & ~n26050;
  assign n26052 = n26013 & n26051;
  assign n26053 = ~n26013 & ~n26051;
  assign n26054 = ~n26052 & ~n26053;
  assign n26055 = n26002 & ~n26054;
  assign n26056 = ~n26002 & n26054;
  assign n26057 = ~n26055 & ~n26056;
  assign n26058 = ~n25996 & ~n25999;
  assign n26059 = n26057 & ~n26058;
  assign n26060 = ~n26057 & n26058;
  assign po119  = ~n26059 & ~n26060;
  assign n26062 = ~n26036 & ~n26049;
  assign n26063 = pi127  & n11193;
  assign n26064 = pi125  & n11567;
  assign n26065 = pi126  & n11188;
  assign n26066 = ~n26064 & ~n26065;
  assign n26067 = ~n26063 & n26066;
  assign n26068 = n11196 & n13365;
  assign n26069 = n26067 & ~n26068;
  assign n26070 = pi59  & ~n26069;
  assign n26071 = pi59  & ~n26070;
  assign n26072 = ~n26069 & ~n26070;
  assign n26073 = ~n26071 & ~n26072;
  assign n26074 = ~n26062 & ~n26073;
  assign n26075 = ~n26062 & ~n26074;
  assign n26076 = ~n26073 & ~n26074;
  assign n26077 = ~n26075 & ~n26076;
  assign n26078 = ~n26029 & ~n26032;
  assign n26079 = pi120  & n13477;
  assign n26080 = pi121  & ~n13122;
  assign n26081 = ~n26079 & ~n26080;
  assign n26082 = ~pi56  & ~n26081;
  assign n26083 = pi56  & n26081;
  assign n26084 = ~n26082 & ~n26083;
  assign n26085 = ~n25956 & n26084;
  assign n26086 = n25956 & ~n26084;
  assign n26087 = ~n26085 & ~n26086;
  assign n26088 = n26078 & ~n26087;
  assign n26089 = ~n26078 & n26087;
  assign n26090 = ~n26088 & ~n26089;
  assign n26091 = pi124  & n12295;
  assign n26092 = pi122  & n12693;
  assign n26093 = pi123  & n12290;
  assign n26094 = ~n26092 & ~n26093;
  assign n26095 = ~n26091 & n26094;
  assign n26096 = n11858 & n12298;
  assign n26097 = n26095 & ~n26096;
  assign n26098 = pi62  & ~n26097;
  assign n26099 = pi62  & ~n26098;
  assign n26100 = ~n26097 & ~n26098;
  assign n26101 = ~n26099 & ~n26100;
  assign n26102 = n26090 & ~n26101;
  assign n26103 = ~n26090 & n26101;
  assign n26104 = ~n26077 & ~n26103;
  assign n26105 = ~n26102 & n26104;
  assign n26106 = ~n26077 & ~n26105;
  assign n26107 = ~n26103 & ~n26105;
  assign n26108 = ~n26102 & n26107;
  assign n26109 = ~n26106 & ~n26108;
  assign n26110 = ~n26011 & ~n26052;
  assign n26111 = n26109 & n26110;
  assign n26112 = ~n26109 & ~n26110;
  assign n26113 = ~n26111 & ~n26112;
  assign n26114 = ~n26056 & ~n26059;
  assign n26115 = n26113 & ~n26114;
  assign n26116 = ~n26113 & n26114;
  assign po120  = ~n26115 & ~n26116;
  assign n26118 = ~n26089 & ~n26102;
  assign n26119 = pi121  & n13477;
  assign n26120 = pi122  & ~n13122;
  assign n26121 = ~n26119 & ~n26120;
  assign n26122 = ~n26082 & ~n26085;
  assign n26123 = ~n26121 & n26122;
  assign n26124 = n26121 & ~n26122;
  assign n26125 = ~n26123 & ~n26124;
  assign n26126 = pi125  & n12295;
  assign n26127 = pi123  & n12693;
  assign n26128 = pi124  & n12290;
  assign n26129 = ~n26127 & ~n26128;
  assign n26130 = ~n26126 & n26129;
  assign n26131 = ~n12298 & n26130;
  assign n26132 = ~n12591 & n26130;
  assign n26133 = ~n26131 & ~n26132;
  assign n26134 = pi62  & ~n26133;
  assign n26135 = ~pi62  & n26133;
  assign n26136 = ~n26134 & ~n26135;
  assign n26137 = n26125 & ~n26136;
  assign n26138 = ~n26125 & n26136;
  assign n26139 = ~n26137 & ~n26138;
  assign n26140 = ~n26118 & n26139;
  assign n26141 = n26118 & ~n26139;
  assign n26142 = ~n26140 & ~n26141;
  assign n26143 = pi126  & n11567;
  assign n26144 = pi127  & n11188;
  assign n26145 = ~n26143 & ~n26144;
  assign n26146 = n11196 & n13389;
  assign n26147 = n26145 & ~n26146;
  assign n26148 = pi59  & ~n26147;
  assign n26149 = pi59  & ~n26148;
  assign n26150 = ~n26147 & ~n26148;
  assign n26151 = ~n26149 & ~n26150;
  assign n26152 = n26142 & ~n26151;
  assign n26153 = n26142 & ~n26152;
  assign n26154 = ~n26151 & ~n26152;
  assign n26155 = ~n26153 & ~n26154;
  assign n26156 = ~n26074 & ~n26105;
  assign n26157 = n26155 & n26156;
  assign n26158 = ~n26155 & ~n26156;
  assign n26159 = ~n26157 & ~n26158;
  assign n26160 = ~n26112 & ~n26115;
  assign n26161 = n26159 & ~n26160;
  assign n26162 = ~n26159 & n26160;
  assign po121  = ~n26161 & ~n26162;
  assign n26164 = ~n26158 & ~n26161;
  assign n26165 = ~n26140 & ~n26152;
  assign n26166 = ~n26124 & ~n26137;
  assign n26167 = pi122  & n13477;
  assign n26168 = pi123  & ~n13122;
  assign n26169 = ~n26167 & ~n26168;
  assign n26170 = n26121 & ~n26169;
  assign n26171 = ~n26121 & n26169;
  assign n26172 = ~n26166 & ~n26171;
  assign n26173 = ~n26170 & n26172;
  assign n26174 = ~n26166 & ~n26173;
  assign n26175 = ~n26171 & ~n26173;
  assign n26176 = ~n26170 & n26175;
  assign n26177 = ~n26174 & ~n26176;
  assign n26178 = pi126  & n12295;
  assign n26179 = pi124  & n12693;
  assign n26180 = pi125  & n12290;
  assign n26181 = ~n26179 & ~n26180;
  assign n26182 = ~n26178 & n26181;
  assign n26183 = n12298 & n12979;
  assign n26184 = n26182 & ~n26183;
  assign n26185 = pi62  & ~n26184;
  assign n26186 = pi62  & ~n26185;
  assign n26187 = ~n26184 & ~n26185;
  assign n26188 = ~n26186 & ~n26187;
  assign n26189 = pi127  & n11567;
  assign n26190 = n11196 & n13387;
  assign n26191 = ~n26189 & ~n26190;
  assign n26192 = pi59  & ~n26191;
  assign n26193 = pi59  & ~n26192;
  assign n26194 = ~n26191 & ~n26192;
  assign n26195 = ~n26193 & ~n26194;
  assign n26196 = ~n26188 & ~n26195;
  assign n26197 = n26188 & n26195;
  assign n26198 = ~n26196 & ~n26197;
  assign n26199 = ~n26177 & n26198;
  assign n26200 = n26177 & ~n26198;
  assign n26201 = ~n26199 & ~n26200;
  assign n26202 = ~n26165 & n26201;
  assign n26203 = n26165 & ~n26201;
  assign n26204 = ~n26202 & ~n26203;
  assign n26205 = ~n26164 & n26204;
  assign n26206 = n26164 & ~n26204;
  assign po122  = ~n26205 & ~n26206;
  assign n26208 = ~n26202 & ~n26205;
  assign n26209 = ~n26196 & ~n26199;
  assign n26210 = pi123  & n13477;
  assign n26211 = pi124  & ~n13122;
  assign n26212 = ~n26210 & ~n26211;
  assign n26213 = ~pi59  & ~n26169;
  assign n26214 = pi59  & n26169;
  assign n26215 = ~n26213 & ~n26214;
  assign n26216 = n26212 & ~n26215;
  assign n26217 = ~n26212 & n26215;
  assign n26218 = ~n26216 & ~n26217;
  assign n26219 = pi127  & n12295;
  assign n26220 = pi125  & n12693;
  assign n26221 = pi126  & n12290;
  assign n26222 = ~n26220 & ~n26221;
  assign n26223 = ~n26219 & n26222;
  assign n26224 = n12298 & n13365;
  assign n26225 = n26223 & ~n26224;
  assign n26226 = pi62  & ~n26225;
  assign n26227 = pi62  & ~n26226;
  assign n26228 = ~n26225 & ~n26226;
  assign n26229 = ~n26227 & ~n26228;
  assign n26230 = n26218 & ~n26229;
  assign n26231 = ~n26218 & n26229;
  assign n26232 = ~n26230 & ~n26231;
  assign n26233 = ~n26175 & n26232;
  assign n26234 = n26175 & ~n26232;
  assign n26235 = ~n26233 & ~n26234;
  assign n26236 = ~n26209 & n26235;
  assign n26237 = ~n26209 & ~n26236;
  assign n26238 = n26235 & ~n26236;
  assign n26239 = ~n26237 & ~n26238;
  assign n26240 = ~n26208 & ~n26239;
  assign n26241 = n26208 & n26239;
  assign po123  = ~n26240 & ~n26241;
  assign n26243 = ~n26236 & ~n26240;
  assign n26244 = ~n26230 & ~n26233;
  assign n26245 = pi124  & n13477;
  assign n26246 = pi125  & ~n13122;
  assign n26247 = ~n26245 & ~n26246;
  assign n26248 = ~n26213 & ~n26217;
  assign n26249 = n26247 & ~n26248;
  assign n26250 = ~n26247 & n26248;
  assign n26251 = ~n26249 & ~n26250;
  assign n26252 = pi126  & n12693;
  assign n26253 = pi127  & n12290;
  assign n26254 = ~n26252 & ~n26253;
  assign n26255 = ~n12298 & n26254;
  assign n26256 = ~n13389 & n26254;
  assign n26257 = ~n26255 & ~n26256;
  assign n26258 = pi62  & ~n26257;
  assign n26259 = ~pi62  & n26257;
  assign n26260 = ~n26258 & ~n26259;
  assign n26261 = n26251 & ~n26260;
  assign n26262 = ~n26251 & n26260;
  assign n26263 = ~n26261 & ~n26262;
  assign n26264 = ~n26244 & n26263;
  assign n26265 = n26244 & ~n26263;
  assign n26266 = ~n26264 & ~n26265;
  assign n26267 = ~n26243 & n26266;
  assign n26268 = n26243 & ~n26266;
  assign po124  = ~n26267 & ~n26268;
  assign n26270 = ~n26264 & ~n26267;
  assign n26271 = ~n26249 & ~n26261;
  assign n26272 = pi125  & n13477;
  assign n26273 = pi126  & ~n13122;
  assign n26274 = ~n26272 & ~n26273;
  assign n26275 = n26247 & ~n26274;
  assign n26276 = ~n26247 & n26274;
  assign n26277 = ~n26275 & ~n26276;
  assign n26278 = pi127  & n12693;
  assign n26279 = ~n12298 & ~n26278;
  assign n26280 = ~n13387 & ~n26278;
  assign n26281 = ~n26279 & ~n26280;
  assign n26282 = pi62  & ~n26281;
  assign n26283 = ~pi62  & n26281;
  assign n26284 = ~n26282 & ~n26283;
  assign n26285 = n26277 & ~n26284;
  assign n26286 = ~n26277 & n26284;
  assign n26287 = ~n26285 & ~n26286;
  assign n26288 = ~n26271 & n26287;
  assign n26289 = n26271 & ~n26287;
  assign n26290 = ~n26288 & ~n26289;
  assign n26291 = ~n26270 & n26290;
  assign n26292 = n26270 & ~n26290;
  assign po125  = ~n26291 & ~n26292;
  assign n26294 = ~n26288 & ~n26291;
  assign n26295 = ~n26275 & ~n26285;
  assign n26296 = pi126  & n13477;
  assign n26297 = pi127  & ~n13122;
  assign n26298 = ~n26296 & ~n26297;
  assign n26299 = ~pi62  & ~n26298;
  assign n26300 = pi62  & n26298;
  assign n26301 = ~n26299 & ~n26300;
  assign n26302 = ~n26247 & n26301;
  assign n26303 = n26247 & ~n26301;
  assign n26304 = ~n26302 & ~n26303;
  assign n26305 = ~n26295 & n26304;
  assign n26306 = n26295 & ~n26304;
  assign n26307 = ~n26305 & ~n26306;
  assign n26308 = ~n26294 & n26307;
  assign n26309 = n26294 & ~n26307;
  assign po126  = ~n26308 & ~n26309;
  assign n26311 = ~n26299 & ~n26302;
  assign n26312 = pi127  & n13477;
  assign n26313 = ~n26311 & n26312;
  assign n26314 = n26311 & ~n26312;
  assign n26315 = ~n26313 & ~n26314;
  assign n26316 = ~n26305 & ~n26308;
  assign n26317 = n26315 & n26316;
  assign n26318 = ~n26315 & ~n26316;
  assign po127  = ~n26317 & ~n26318;
endmodule
