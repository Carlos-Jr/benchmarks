module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 , pi128 , pi129 , pi130 ,
    pi131 , pi132 , pi133 , pi134 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 , pi128 , pi129 ,
    pi130 , pi131 , pi132 , pi133 , pi134 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ;
  wire n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132,
    n1133, n1134, n1135, n1136, n1137, n1138,
    n1139, n1140, n1141, n1142, n1143, n1144,
    n1145, n1146, n1147, n1148, n1149, n1150,
    n1151, n1152, n1153, n1154, n1155, n1156,
    n1157, n1158, n1159, n1160, n1161, n1162,
    n1163, n1164, n1165, n1166, n1167, n1168,
    n1169, n1170, n1171, n1172, n1173, n1174,
    n1175, n1176, n1177, n1178, n1179, n1180,
    n1181, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198,
    n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1206, n1207, n1208, n1209, n1210,
    n1211, n1212, n1213, n1214, n1215, n1216,
    n1217, n1218, n1219, n1220, n1221, n1222,
    n1223, n1224, n1225, n1226, n1227, n1228,
    n1229, n1230, n1231, n1232, n1233, n1234,
    n1235, n1236, n1237, n1238, n1239, n1240,
    n1241, n1242, n1243, n1244, n1245, n1246,
    n1247, n1248, n1249, n1250, n1251, n1252,
    n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264,
    n1265, n1266, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294,
    n1295, n1296, n1297, n1298, n1299, n1300,
    n1301, n1302, n1303, n1304, n1305, n1306,
    n1307, n1308, n1309, n1310, n1311, n1312,
    n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324,
    n1325, n1326, n1327, n1328, n1329, n1330,
    n1331, n1332, n1333, n1334, n1335, n1336,
    n1337, n1338, n1339, n1340, n1341, n1342,
    n1343, n1344, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1362, n1363, n1364, n1365, n1366,
    n1367, n1368, n1369, n1370, n1371, n1372,
    n1373, n1374, n1375, n1376, n1377, n1378,
    n1379, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396,
    n1397, n1398, n1399, n1400, n1401, n1402,
    n1403, n1404, n1405, n1406, n1407, n1408,
    n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1419, n1420, n1421,
    n1422, n1423, n1424, n1425, n1426, n1427,
    n1428, n1429, n1430, n1431, n1432, n1433,
    n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445,
    n1446, n1447, n1448, n1449, n1450, n1451,
    n1452, n1453, n1454, n1455, n1456, n1457,
    n1458, n1459, n1460, n1461, n1462, n1463,
    n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481,
    n1482, n1483, n1484, n1485, n1486, n1487,
    n1488, n1489, n1490, n1491, n1492, n1493,
    n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517,
    n1518, n1519, n1520, n1521, n1522, n1523,
    n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541,
    n1542, n1543, n1544, n1545, n1546, n1547,
    n1548, n1549, n1550, n1551, n1552, n1553,
    n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571,
    n1572, n1573, n1574, n1575, n1576, n1577,
    n1578, n1579, n1580, n1581, n1582, n1583,
    n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1598, n1599, n1600, n1601,
    n1602, n1603, n1604, n1605, n1606, n1607,
    n1608, n1609, n1610, n1611, n1612, n1613,
    n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625,
    n1626, n1627, n1628, n1629, n1630, n1631,
    n1632, n1633, n1634, n1635, n1636, n1637,
    n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661,
    n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1716,
    n1717, n1718, n1719, n1720, n1721, n1722,
    n1723, n1724, n1725, n1726, n1727, n1728,
    n1729, n1730, n1731, n1732, n1733, n1734,
    n1735, n1736, n1737, n1738, n1739, n1740,
    n1741, n1742, n1743, n1744, n1745, n1746,
    n1747, n1748, n1749, n1750, n1751, n1752,
    n1753, n1754, n1755, n1756, n1757, n1758,
    n1759, n1760, n1761, n1762, n1763, n1764,
    n1765, n1766, n1767, n1768, n1769, n1770,
    n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782,
    n1783, n1784, n1785, n1786, n1787, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795,
    n1796, n1797, n1798, n1799, n1800, n1801,
    n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813,
    n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825,
    n1826, n1827, n1828, n1829, n1830, n1831,
    n1832, n1833, n1834, n1835, n1836, n1837,
    n1838, n1839, n1840, n1841, n1842, n1843,
    n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855,
    n1856, n1857, n1858, n1859, n1860, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2008,
    n2009, n2010, n2011, n2012, n2013, n2014,
    n2015, n2016, n2017, n2018, n2019, n2020,
    n2021, n2022, n2023, n2024, n2025, n2026,
    n2027, n2028, n2029, n2030, n2031, n2032,
    n2033, n2034, n2035, n2036, n2037, n2038,
    n2039, n2040, n2041, n2042, n2043, n2044,
    n2045, n2046, n2047, n2048, n2049, n2050,
    n2051, n2052, n2053, n2054, n2055, n2056,
    n2057, n2058, n2059, n2060, n2061, n2062,
    n2063, n2064, n2065, n2066, n2067, n2068,
    n2069, n2070, n2071, n2072, n2073, n2074,
    n2075, n2076, n2077, n2078, n2079, n2081,
    n2082, n2083, n2084, n2085, n2086, n2087,
    n2088, n2089, n2090, n2091, n2092, n2093,
    n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105,
    n2106, n2107, n2108, n2109, n2110, n2111,
    n2112, n2113, n2114, n2115, n2116, n2117,
    n2118, n2119, n2120, n2121, n2122, n2123,
    n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135,
    n2136, n2137, n2138, n2139, n2140, n2141,
    n2142, n2143, n2144, n2145, n2146, n2147,
    n2148, n2149, n2150, n2151, n2152, n2154,
    n2155, n2156, n2157, n2158, n2159, n2160,
    n2161, n2162, n2163, n2164, n2165, n2166,
    n2167, n2168, n2169, n2170, n2171, n2172,
    n2173, n2174, n2175, n2176, n2177, n2178,
    n2179, n2180, n2181, n2182, n2183, n2184,
    n2185, n2186, n2187, n2188, n2189, n2190,
    n2191, n2192, n2193, n2194, n2195, n2196,
    n2197, n2198, n2199, n2200, n2201, n2202,
    n2203, n2204, n2205, n2206, n2207, n2208,
    n2209, n2210, n2211, n2212, n2213, n2214,
    n2215, n2216, n2217, n2218, n2219, n2220,
    n2221, n2222, n2223, n2224, n2225, n2227,
    n2228, n2229, n2230, n2231, n2232, n2233,
    n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245,
    n2246, n2247, n2248, n2249, n2250, n2251,
    n2252, n2253, n2254, n2255, n2256, n2257,
    n2258, n2259, n2260, n2261, n2262, n2263,
    n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275,
    n2276, n2277, n2278, n2279, n2280, n2281,
    n2282, n2283, n2284, n2285, n2286, n2287,
    n2288, n2289, n2290, n2291, n2292, n2293,
    n2294, n2295, n2296, n2297, n2298, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2446,
    n2447, n2448, n2449, n2450, n2451, n2452,
    n2453, n2454, n2455, n2456, n2457, n2458,
    n2459, n2460, n2461, n2462, n2463, n2464,
    n2465, n2466, n2467, n2468, n2469, n2470,
    n2471, n2472, n2473, n2474, n2475, n2476,
    n2477, n2478, n2479, n2480, n2481, n2482,
    n2483, n2484, n2485, n2486, n2487, n2488,
    n2489, n2490, n2491, n2492, n2493, n2494,
    n2495, n2496, n2497, n2498, n2499, n2500,
    n2501, n2502, n2503, n2504, n2505, n2506,
    n2507, n2508, n2509, n2510, n2511, n2512,
    n2513, n2514, n2515, n2516, n2517, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525,
    n2526, n2527, n2528, n2529, n2530, n2531,
    n2532, n2533, n2534, n2535, n2536, n2537,
    n2538, n2539, n2540, n2541, n2542, n2543,
    n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555,
    n2556, n2557, n2558, n2559, n2560, n2561,
    n2562, n2563, n2564, n2565, n2566, n2567,
    n2568, n2569, n2570, n2571, n2572, n2573,
    n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585,
    n2586, n2587, n2588, n2589, n2590, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2609, n2610, n2611,
    n2612, n2613, n2614, n2615, n2616, n2617,
    n2618, n2619, n2620, n2621, n2622, n2623,
    n2624, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2677, n2678, n2679, n2680, n2681,
    n2682, n2683, n2684, n2685, n2686, n2687,
    n2688, n2689, n2690, n2691, n2692, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2711, n2712, n2713,
    n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725,
    n2726, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2762, n2763, n2764,
    n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2779, n2780, n2781, n2782, n2783,
    n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2813, n2814, n2815,
    n2816, n2817, n2818, n2819, n2820, n2821,
    n2822, n2823, n2824, n2825, n2826, n2827,
    n2828, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2864, n2865, n2866,
    n2867, n2868, n2869, n2870, n2871, n2872,
    n2873, n2874, n2875, n2876, n2877, n2878,
    n2879, n2881, n2882, n2883, n2884, n2885,
    n2886, n2887, n2888, n2889, n2890, n2891,
    n2892, n2893, n2894, n2895, n2896, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2915, n2916, n2917,
    n2918, n2919, n2920, n2921, n2922, n2923,
    n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2966, n2967, n2968,
    n2969, n2970, n2971, n2972, n2973, n2974,
    n2975, n2976, n2977, n2978, n2979, n2980,
    n2981, n2983, n2984, n2985, n2986, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025,
    n3026, n3027, n3028, n3029, n3030, n3031,
    n3032, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3068, n3069, n3070,
    n3071, n3072, n3073, n3074, n3075, n3076,
    n3077, n3078, n3079, n3080, n3081, n3082,
    n3083, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095,
    n3096, n3097, n3098, n3099, n3100, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3119, n3120, n3121,
    n3122, n3123, n3124, n3125, n3126, n3127,
    n3128, n3129, n3130, n3131, n3132, n3133,
    n3134, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3170, n3171, n3172,
    n3173, n3174, n3175, n3176, n3177, n3178,
    n3179, n3180, n3181, n3182, n3183, n3184,
    n3185, n3187, n3188, n3189, n3190, n3191,
    n3192, n3193, n3194, n3195, n3196, n3197,
    n3198, n3199, n3200, n3201, n3202, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3221, n3222, n3223,
    n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235,
    n3236, n3238, n3239, n3240, n3241, n3242,
    n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3272, n3273, n3274,
    n3275, n3276, n3277, n3278, n3279, n3280,
    n3281, n3282, n3283, n3284, n3285, n3286,
    n3287, n3289, n3290, n3291, n3292, n3293,
    n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3306,
    n3307, n3308, n3309, n3310, n3311, n3312,
    n3313, n3314, n3315, n3316, n3317, n3318,
    n3319, n3320, n3321, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3374, n3375, n3376,
    n3377, n3378, n3379, n3380, n3381, n3382,
    n3383, n3384, n3385, n3386, n3387, n3388,
    n3389, n3391, n3392, n3393, n3394, n3395,
    n3396, n3397, n3398, n3399, n3400, n3401,
    n3402, n3403, n3404, n3405, n3406, n3408,
    n3409, n3411, n3412, n3414, n3415, n3417,
    n3418, n3420, n3421, n3423, n3424, n3426,
    n3427, n3429, n3430, n3432, n3433, n3435,
    n3436, n3438, n3439, n3441, n3442, n3444,
    n3445, n3447, n3448, n3450, n3451, n3453,
    n3454, n3456, n3457, n3459, n3460, n3462,
    n3463, n3465, n3466, n3468, n3469, n3471,
    n3472, n3474, n3475, n3477, n3478, n3480,
    n3481, n3483, n3484, n3486, n3487, n3489,
    n3490, n3492, n3493, n3495, n3496, n3498,
    n3499, n3501, n3502, n3504, n3505, n3507,
    n3508, n3510, n3511, n3513, n3514, n3516,
    n3517, n3519, n3520, n3522, n3523, n3525,
    n3526, n3528, n3529, n3531, n3532, n3534,
    n3535, n3537, n3538, n3540, n3541, n3543,
    n3544, n3546, n3547, n3549, n3550, n3552,
    n3553, n3555, n3556, n3558, n3559, n3561,
    n3562, n3564, n3565, n3567, n3568, n3570,
    n3571, n3573, n3574, n3576, n3577, n3579,
    n3580, n3582, n3583, n3585, n3586, n3588,
    n3589, n3591, n3592, n3594, n3595, n3597,
    n3598;
  assign n264 = pi77  & pi128 ;
  assign n265 = pi129  & n264;
  assign n266 = pi78  & ~pi128 ;
  assign n267 = pi129  & n266;
  assign n268 = pi80  & ~pi128 ;
  assign n269 = ~pi129  & n268;
  assign n270 = pi79  & pi128 ;
  assign n271 = ~pi129  & n270;
  assign n272 = ~n265 & ~n267;
  assign n273 = ~n269 & ~n271;
  assign n274 = n272 & n273;
  assign n275 = ~pi130  & ~pi131 ;
  assign n276 = ~n274 & n275;
  assign n277 = pi73  & pi128 ;
  assign n278 = pi129  & n277;
  assign n279 = pi74  & ~pi128 ;
  assign n280 = pi129  & n279;
  assign n281 = pi76  & ~pi128 ;
  assign n282 = ~pi129  & n281;
  assign n283 = pi75  & pi128 ;
  assign n284 = ~pi129  & n283;
  assign n285 = ~n278 & ~n280;
  assign n286 = ~n282 & ~n284;
  assign n287 = n285 & n286;
  assign n288 = pi130  & ~pi131 ;
  assign n289 = ~n287 & n288;
  assign n290 = pi65  & pi128 ;
  assign n291 = pi129  & n290;
  assign n292 = pi66  & ~pi128 ;
  assign n293 = pi129  & n292;
  assign n294 = pi68  & ~pi128 ;
  assign n295 = ~pi129  & n294;
  assign n296 = pi67  & pi128 ;
  assign n297 = ~pi129  & n296;
  assign n298 = ~n291 & ~n293;
  assign n299 = ~n295 & ~n297;
  assign n300 = n298 & n299;
  assign n301 = pi130  & pi131 ;
  assign n302 = ~n300 & n301;
  assign n303 = pi69  & pi128 ;
  assign n304 = pi129  & n303;
  assign n305 = pi70  & ~pi128 ;
  assign n306 = pi129  & n305;
  assign n307 = pi72  & ~pi128 ;
  assign n308 = ~pi129  & n307;
  assign n309 = pi71  & pi128 ;
  assign n310 = ~pi129  & n309;
  assign n311 = ~n304 & ~n306;
  assign n312 = ~n308 & ~n310;
  assign n313 = n311 & n312;
  assign n314 = ~pi130  & pi131 ;
  assign n315 = ~n313 & n314;
  assign n316 = ~n276 & ~n289;
  assign n317 = ~n302 & ~n315;
  assign n318 = n316 & n317;
  assign n319 = pi132  & pi133 ;
  assign n320 = ~n318 & n319;
  assign n321 = pi93  & pi128 ;
  assign n322 = pi129  & n321;
  assign n323 = pi94  & ~pi128 ;
  assign n324 = pi129  & n323;
  assign n325 = pi96  & ~pi128 ;
  assign n326 = ~pi129  & n325;
  assign n327 = pi95  & pi128 ;
  assign n328 = ~pi129  & n327;
  assign n329 = ~n322 & ~n324;
  assign n330 = ~n326 & ~n328;
  assign n331 = n329 & n330;
  assign n332 = n275 & ~n331;
  assign n333 = pi89  & pi128 ;
  assign n334 = pi129  & n333;
  assign n335 = pi90  & ~pi128 ;
  assign n336 = pi129  & n335;
  assign n337 = pi92  & ~pi128 ;
  assign n338 = ~pi129  & n337;
  assign n339 = pi91  & pi128 ;
  assign n340 = ~pi129  & n339;
  assign n341 = ~n334 & ~n336;
  assign n342 = ~n338 & ~n340;
  assign n343 = n341 & n342;
  assign n344 = n288 & ~n343;
  assign n345 = pi81  & pi128 ;
  assign n346 = pi129  & n345;
  assign n347 = pi82  & ~pi128 ;
  assign n348 = pi129  & n347;
  assign n349 = pi84  & ~pi128 ;
  assign n350 = ~pi129  & n349;
  assign n351 = pi83  & pi128 ;
  assign n352 = ~pi129  & n351;
  assign n353 = ~n346 & ~n348;
  assign n354 = ~n350 & ~n352;
  assign n355 = n353 & n354;
  assign n356 = n301 & ~n355;
  assign n357 = pi85  & pi128 ;
  assign n358 = pi129  & n357;
  assign n359 = pi86  & ~pi128 ;
  assign n360 = pi129  & n359;
  assign n361 = pi88  & ~pi128 ;
  assign n362 = ~pi129  & n361;
  assign n363 = pi87  & pi128 ;
  assign n364 = ~pi129  & n363;
  assign n365 = ~n358 & ~n360;
  assign n366 = ~n362 & ~n364;
  assign n367 = n365 & n366;
  assign n368 = n314 & ~n367;
  assign n369 = ~n332 & ~n344;
  assign n370 = ~n356 & ~n368;
  assign n371 = n369 & n370;
  assign n372 = ~pi132  & pi133 ;
  assign n373 = ~n371 & n372;
  assign n374 = pi125  & pi128 ;
  assign n375 = pi129  & n374;
  assign n376 = pi126  & ~pi128 ;
  assign n377 = pi129  & n376;
  assign n378 = pi0  & ~pi128 ;
  assign n379 = ~pi129  & n378;
  assign n380 = pi127  & pi128 ;
  assign n381 = ~pi129  & n380;
  assign n382 = ~n375 & ~n377;
  assign n383 = ~n379 & ~n381;
  assign n384 = n382 & n383;
  assign n385 = n275 & ~n384;
  assign n386 = pi121  & pi128 ;
  assign n387 = pi129  & n386;
  assign n388 = pi122  & ~pi128 ;
  assign n389 = pi129  & n388;
  assign n390 = pi124  & ~pi128 ;
  assign n391 = ~pi129  & n390;
  assign n392 = pi123  & pi128 ;
  assign n393 = ~pi129  & n392;
  assign n394 = ~n387 & ~n389;
  assign n395 = ~n391 & ~n393;
  assign n396 = n394 & n395;
  assign n397 = n288 & ~n396;
  assign n398 = pi113  & pi128 ;
  assign n399 = pi129  & n398;
  assign n400 = pi114  & ~pi128 ;
  assign n401 = pi129  & n400;
  assign n402 = pi116  & ~pi128 ;
  assign n403 = ~pi129  & n402;
  assign n404 = pi115  & pi128 ;
  assign n405 = ~pi129  & n404;
  assign n406 = ~n399 & ~n401;
  assign n407 = ~n403 & ~n405;
  assign n408 = n406 & n407;
  assign n409 = n301 & ~n408;
  assign n410 = pi117  & pi128 ;
  assign n411 = pi129  & n410;
  assign n412 = pi118  & ~pi128 ;
  assign n413 = pi129  & n412;
  assign n414 = pi120  & ~pi128 ;
  assign n415 = ~pi129  & n414;
  assign n416 = pi119  & pi128 ;
  assign n417 = ~pi129  & n416;
  assign n418 = ~n411 & ~n413;
  assign n419 = ~n415 & ~n417;
  assign n420 = n418 & n419;
  assign n421 = n314 & ~n420;
  assign n422 = ~n385 & ~n397;
  assign n423 = ~n409 & ~n421;
  assign n424 = n422 & n423;
  assign n425 = ~pi132  & ~pi133 ;
  assign n426 = ~n424 & n425;
  assign n427 = pi109  & pi128 ;
  assign n428 = pi129  & n427;
  assign n429 = pi110  & ~pi128 ;
  assign n430 = pi129  & n429;
  assign n431 = pi112  & ~pi128 ;
  assign n432 = ~pi129  & n431;
  assign n433 = pi111  & pi128 ;
  assign n434 = ~pi129  & n433;
  assign n435 = ~n428 & ~n430;
  assign n436 = ~n432 & ~n434;
  assign n437 = n435 & n436;
  assign n438 = n275 & ~n437;
  assign n439 = pi105  & pi128 ;
  assign n440 = pi129  & n439;
  assign n441 = pi106  & ~pi128 ;
  assign n442 = pi129  & n441;
  assign n443 = pi108  & ~pi128 ;
  assign n444 = ~pi129  & n443;
  assign n445 = pi107  & pi128 ;
  assign n446 = ~pi129  & n445;
  assign n447 = ~n440 & ~n442;
  assign n448 = ~n444 & ~n446;
  assign n449 = n447 & n448;
  assign n450 = n288 & ~n449;
  assign n451 = pi97  & pi128 ;
  assign n452 = pi129  & n451;
  assign n453 = pi98  & ~pi128 ;
  assign n454 = pi129  & n453;
  assign n455 = pi100  & ~pi128 ;
  assign n456 = ~pi129  & n455;
  assign n457 = pi99  & pi128 ;
  assign n458 = ~pi129  & n457;
  assign n459 = ~n452 & ~n454;
  assign n460 = ~n456 & ~n458;
  assign n461 = n459 & n460;
  assign n462 = n301 & ~n461;
  assign n463 = pi101  & pi128 ;
  assign n464 = pi129  & n463;
  assign n465 = pi102  & ~pi128 ;
  assign n466 = pi129  & n465;
  assign n467 = pi104  & ~pi128 ;
  assign n468 = ~pi129  & n467;
  assign n469 = pi103  & pi128 ;
  assign n470 = ~pi129  & n469;
  assign n471 = ~n464 & ~n466;
  assign n472 = ~n468 & ~n470;
  assign n473 = n471 & n472;
  assign n474 = n314 & ~n473;
  assign n475 = ~n438 & ~n450;
  assign n476 = ~n462 & ~n474;
  assign n477 = n475 & n476;
  assign n478 = pi132  & ~pi133 ;
  assign n479 = ~n477 & n478;
  assign n480 = ~n320 & ~n373;
  assign n481 = ~n426 & ~n479;
  assign n482 = n480 & n481;
  assign n483 = ~pi134  & ~n482;
  assign n484 = pi13  & pi128 ;
  assign n485 = pi129  & n484;
  assign n486 = pi14  & ~pi128 ;
  assign n487 = pi129  & n486;
  assign n488 = pi16  & ~pi128 ;
  assign n489 = ~pi129  & n488;
  assign n490 = pi15  & pi128 ;
  assign n491 = ~pi129  & n490;
  assign n492 = ~n485 & ~n487;
  assign n493 = ~n489 & ~n491;
  assign n494 = n492 & n493;
  assign n495 = n275 & ~n494;
  assign n496 = pi9  & pi128 ;
  assign n497 = pi129  & n496;
  assign n498 = pi10  & ~pi128 ;
  assign n499 = pi129  & n498;
  assign n500 = pi12  & ~pi128 ;
  assign n501 = ~pi129  & n500;
  assign n502 = pi11  & pi128 ;
  assign n503 = ~pi129  & n502;
  assign n504 = ~n497 & ~n499;
  assign n505 = ~n501 & ~n503;
  assign n506 = n504 & n505;
  assign n507 = n288 & ~n506;
  assign n508 = pi1  & pi128 ;
  assign n509 = pi129  & n508;
  assign n510 = pi2  & ~pi128 ;
  assign n511 = pi129  & n510;
  assign n512 = pi4  & ~pi128 ;
  assign n513 = ~pi129  & n512;
  assign n514 = pi3  & pi128 ;
  assign n515 = ~pi129  & n514;
  assign n516 = ~n509 & ~n511;
  assign n517 = ~n513 & ~n515;
  assign n518 = n516 & n517;
  assign n519 = n301 & ~n518;
  assign n520 = pi5  & pi128 ;
  assign n521 = pi129  & n520;
  assign n522 = pi6  & ~pi128 ;
  assign n523 = pi129  & n522;
  assign n524 = pi8  & ~pi128 ;
  assign n525 = ~pi129  & n524;
  assign n526 = pi7  & pi128 ;
  assign n527 = ~pi129  & n526;
  assign n528 = ~n521 & ~n523;
  assign n529 = ~n525 & ~n527;
  assign n530 = n528 & n529;
  assign n531 = n314 & ~n530;
  assign n532 = ~n495 & ~n507;
  assign n533 = ~n519 & ~n531;
  assign n534 = n532 & n533;
  assign n535 = n319 & ~n534;
  assign n536 = pi29  & pi128 ;
  assign n537 = pi129  & n536;
  assign n538 = pi30  & ~pi128 ;
  assign n539 = pi129  & n538;
  assign n540 = pi32  & ~pi128 ;
  assign n541 = ~pi129  & n540;
  assign n542 = pi31  & pi128 ;
  assign n543 = ~pi129  & n542;
  assign n544 = ~n537 & ~n539;
  assign n545 = ~n541 & ~n543;
  assign n546 = n544 & n545;
  assign n547 = n275 & ~n546;
  assign n548 = pi25  & pi128 ;
  assign n549 = pi129  & n548;
  assign n550 = pi26  & ~pi128 ;
  assign n551 = pi129  & n550;
  assign n552 = pi28  & ~pi128 ;
  assign n553 = ~pi129  & n552;
  assign n554 = pi27  & pi128 ;
  assign n555 = ~pi129  & n554;
  assign n556 = ~n549 & ~n551;
  assign n557 = ~n553 & ~n555;
  assign n558 = n556 & n557;
  assign n559 = n288 & ~n558;
  assign n560 = pi17  & pi128 ;
  assign n561 = pi129  & n560;
  assign n562 = pi18  & ~pi128 ;
  assign n563 = pi129  & n562;
  assign n564 = pi20  & ~pi128 ;
  assign n565 = ~pi129  & n564;
  assign n566 = pi19  & pi128 ;
  assign n567 = ~pi129  & n566;
  assign n568 = ~n561 & ~n563;
  assign n569 = ~n565 & ~n567;
  assign n570 = n568 & n569;
  assign n571 = n301 & ~n570;
  assign n572 = pi21  & pi128 ;
  assign n573 = pi129  & n572;
  assign n574 = pi22  & ~pi128 ;
  assign n575 = pi129  & n574;
  assign n576 = pi24  & ~pi128 ;
  assign n577 = ~pi129  & n576;
  assign n578 = pi23  & pi128 ;
  assign n579 = ~pi129  & n578;
  assign n580 = ~n573 & ~n575;
  assign n581 = ~n577 & ~n579;
  assign n582 = n580 & n581;
  assign n583 = n314 & ~n582;
  assign n584 = ~n547 & ~n559;
  assign n585 = ~n571 & ~n583;
  assign n586 = n584 & n585;
  assign n587 = n372 & ~n586;
  assign n588 = pi61  & pi128 ;
  assign n589 = pi129  & n588;
  assign n590 = pi62  & ~pi128 ;
  assign n591 = pi129  & n590;
  assign n592 = pi64  & ~pi128 ;
  assign n593 = ~pi129  & n592;
  assign n594 = pi63  & pi128 ;
  assign n595 = ~pi129  & n594;
  assign n596 = ~n589 & ~n591;
  assign n597 = ~n593 & ~n595;
  assign n598 = n596 & n597;
  assign n599 = n275 & ~n598;
  assign n600 = pi57  & pi128 ;
  assign n601 = pi129  & n600;
  assign n602 = pi58  & ~pi128 ;
  assign n603 = pi129  & n602;
  assign n604 = pi60  & ~pi128 ;
  assign n605 = ~pi129  & n604;
  assign n606 = pi59  & pi128 ;
  assign n607 = ~pi129  & n606;
  assign n608 = ~n601 & ~n603;
  assign n609 = ~n605 & ~n607;
  assign n610 = n608 & n609;
  assign n611 = n288 & ~n610;
  assign n612 = pi49  & pi128 ;
  assign n613 = pi129  & n612;
  assign n614 = pi50  & ~pi128 ;
  assign n615 = pi129  & n614;
  assign n616 = pi52  & ~pi128 ;
  assign n617 = ~pi129  & n616;
  assign n618 = pi51  & pi128 ;
  assign n619 = ~pi129  & n618;
  assign n620 = ~n613 & ~n615;
  assign n621 = ~n617 & ~n619;
  assign n622 = n620 & n621;
  assign n623 = n301 & ~n622;
  assign n624 = pi53  & pi128 ;
  assign n625 = pi129  & n624;
  assign n626 = pi54  & ~pi128 ;
  assign n627 = pi129  & n626;
  assign n628 = pi56  & ~pi128 ;
  assign n629 = ~pi129  & n628;
  assign n630 = pi55  & pi128 ;
  assign n631 = ~pi129  & n630;
  assign n632 = ~n625 & ~n627;
  assign n633 = ~n629 & ~n631;
  assign n634 = n632 & n633;
  assign n635 = n314 & ~n634;
  assign n636 = ~n599 & ~n611;
  assign n637 = ~n623 & ~n635;
  assign n638 = n636 & n637;
  assign n639 = n425 & ~n638;
  assign n640 = pi45  & pi128 ;
  assign n641 = pi129  & n640;
  assign n642 = pi46  & ~pi128 ;
  assign n643 = pi129  & n642;
  assign n644 = pi48  & ~pi128 ;
  assign n645 = ~pi129  & n644;
  assign n646 = pi47  & pi128 ;
  assign n647 = ~pi129  & n646;
  assign n648 = ~n641 & ~n643;
  assign n649 = ~n645 & ~n647;
  assign n650 = n648 & n649;
  assign n651 = n275 & ~n650;
  assign n652 = pi41  & pi128 ;
  assign n653 = pi129  & n652;
  assign n654 = pi42  & ~pi128 ;
  assign n655 = pi129  & n654;
  assign n656 = pi44  & ~pi128 ;
  assign n657 = ~pi129  & n656;
  assign n658 = pi43  & pi128 ;
  assign n659 = ~pi129  & n658;
  assign n660 = ~n653 & ~n655;
  assign n661 = ~n657 & ~n659;
  assign n662 = n660 & n661;
  assign n663 = n288 & ~n662;
  assign n664 = pi33  & pi128 ;
  assign n665 = pi129  & n664;
  assign n666 = pi34  & ~pi128 ;
  assign n667 = pi129  & n666;
  assign n668 = pi36  & ~pi128 ;
  assign n669 = ~pi129  & n668;
  assign n670 = pi35  & pi128 ;
  assign n671 = ~pi129  & n670;
  assign n672 = ~n665 & ~n667;
  assign n673 = ~n669 & ~n671;
  assign n674 = n672 & n673;
  assign n675 = n301 & ~n674;
  assign n676 = pi40  & ~pi128 ;
  assign n677 = ~pi129  & n676;
  assign n678 = pi37  & pi128 ;
  assign n679 = pi129  & n678;
  assign n680 = pi39  & pi128 ;
  assign n681 = ~pi129  & n680;
  assign n682 = pi38  & ~pi128 ;
  assign n683 = pi129  & n682;
  assign n684 = ~n677 & ~n679;
  assign n685 = ~n681 & ~n683;
  assign n686 = n684 & n685;
  assign n687 = n314 & ~n686;
  assign n688 = ~n651 & ~n663;
  assign n689 = ~n675 & ~n687;
  assign n690 = n688 & n689;
  assign n691 = n478 & ~n690;
  assign n692 = ~n535 & ~n587;
  assign n693 = ~n639 & ~n691;
  assign n694 = n692 & n693;
  assign n695 = pi134  & ~n694;
  assign po0  = n483 | n695;
  assign n697 = pi81  & ~pi128 ;
  assign n698 = ~pi129  & n697;
  assign n699 = pi78  & pi128 ;
  assign n700 = pi129  & n699;
  assign n701 = pi80  & pi128 ;
  assign n702 = ~pi129  & n701;
  assign n703 = pi79  & ~pi128 ;
  assign n704 = pi129  & n703;
  assign n705 = ~n698 & ~n700;
  assign n706 = ~n702 & ~n704;
  assign n707 = n705 & n706;
  assign n708 = n275 & ~n707;
  assign n709 = pi77  & ~pi128 ;
  assign n710 = ~pi129  & n709;
  assign n711 = pi74  & pi128 ;
  assign n712 = pi129  & n711;
  assign n713 = pi76  & pi128 ;
  assign n714 = ~pi129  & n713;
  assign n715 = pi75  & ~pi128 ;
  assign n716 = pi129  & n715;
  assign n717 = ~n710 & ~n712;
  assign n718 = ~n714 & ~n716;
  assign n719 = n717 & n718;
  assign n720 = n288 & ~n719;
  assign n721 = pi69  & ~pi128 ;
  assign n722 = ~pi129  & n721;
  assign n723 = pi66  & pi128 ;
  assign n724 = pi129  & n723;
  assign n725 = pi68  & pi128 ;
  assign n726 = ~pi129  & n725;
  assign n727 = pi67  & ~pi128 ;
  assign n728 = pi129  & n727;
  assign n729 = ~n722 & ~n724;
  assign n730 = ~n726 & ~n728;
  assign n731 = n729 & n730;
  assign n732 = n301 & ~n731;
  assign n733 = pi73  & ~pi128 ;
  assign n734 = ~pi129  & n733;
  assign n735 = pi70  & pi128 ;
  assign n736 = pi129  & n735;
  assign n737 = pi72  & pi128 ;
  assign n738 = ~pi129  & n737;
  assign n739 = pi71  & ~pi128 ;
  assign n740 = pi129  & n739;
  assign n741 = ~n734 & ~n736;
  assign n742 = ~n738 & ~n740;
  assign n743 = n741 & n742;
  assign n744 = n314 & ~n743;
  assign n745 = ~n708 & ~n720;
  assign n746 = ~n732 & ~n744;
  assign n747 = n745 & n746;
  assign n748 = n319 & ~n747;
  assign n749 = pi97  & ~pi128 ;
  assign n750 = ~pi129  & n749;
  assign n751 = pi94  & pi128 ;
  assign n752 = pi129  & n751;
  assign n753 = pi96  & pi128 ;
  assign n754 = ~pi129  & n753;
  assign n755 = pi95  & ~pi128 ;
  assign n756 = pi129  & n755;
  assign n757 = ~n750 & ~n752;
  assign n758 = ~n754 & ~n756;
  assign n759 = n757 & n758;
  assign n760 = n275 & ~n759;
  assign n761 = pi93  & ~pi128 ;
  assign n762 = ~pi129  & n761;
  assign n763 = pi90  & pi128 ;
  assign n764 = pi129  & n763;
  assign n765 = pi92  & pi128 ;
  assign n766 = ~pi129  & n765;
  assign n767 = pi91  & ~pi128 ;
  assign n768 = pi129  & n767;
  assign n769 = ~n762 & ~n764;
  assign n770 = ~n766 & ~n768;
  assign n771 = n769 & n770;
  assign n772 = n288 & ~n771;
  assign n773 = pi85  & ~pi128 ;
  assign n774 = ~pi129  & n773;
  assign n775 = pi82  & pi128 ;
  assign n776 = pi129  & n775;
  assign n777 = pi84  & pi128 ;
  assign n778 = ~pi129  & n777;
  assign n779 = pi83  & ~pi128 ;
  assign n780 = pi129  & n779;
  assign n781 = ~n774 & ~n776;
  assign n782 = ~n778 & ~n780;
  assign n783 = n781 & n782;
  assign n784 = n301 & ~n783;
  assign n785 = pi89  & ~pi128 ;
  assign n786 = ~pi129  & n785;
  assign n787 = pi86  & pi128 ;
  assign n788 = pi129  & n787;
  assign n789 = pi88  & pi128 ;
  assign n790 = ~pi129  & n789;
  assign n791 = pi87  & ~pi128 ;
  assign n792 = pi129  & n791;
  assign n793 = ~n786 & ~n788;
  assign n794 = ~n790 & ~n792;
  assign n795 = n793 & n794;
  assign n796 = n314 & ~n795;
  assign n797 = ~n760 & ~n772;
  assign n798 = ~n784 & ~n796;
  assign n799 = n797 & n798;
  assign n800 = n372 & ~n799;
  assign n801 = pi1  & ~pi128 ;
  assign n802 = ~pi129  & n801;
  assign n803 = pi126  & pi128 ;
  assign n804 = pi129  & n803;
  assign n805 = pi0  & pi128 ;
  assign n806 = ~pi129  & n805;
  assign n807 = pi127  & ~pi128 ;
  assign n808 = pi129  & n807;
  assign n809 = ~n802 & ~n804;
  assign n810 = ~n806 & ~n808;
  assign n811 = n809 & n810;
  assign n812 = n275 & ~n811;
  assign n813 = pi125  & ~pi128 ;
  assign n814 = ~pi129  & n813;
  assign n815 = pi122  & pi128 ;
  assign n816 = pi129  & n815;
  assign n817 = pi124  & pi128 ;
  assign n818 = ~pi129  & n817;
  assign n819 = pi123  & ~pi128 ;
  assign n820 = pi129  & n819;
  assign n821 = ~n814 & ~n816;
  assign n822 = ~n818 & ~n820;
  assign n823 = n821 & n822;
  assign n824 = n288 & ~n823;
  assign n825 = pi117  & ~pi128 ;
  assign n826 = ~pi129  & n825;
  assign n827 = pi114  & pi128 ;
  assign n828 = pi129  & n827;
  assign n829 = pi116  & pi128 ;
  assign n830 = ~pi129  & n829;
  assign n831 = pi115  & ~pi128 ;
  assign n832 = pi129  & n831;
  assign n833 = ~n826 & ~n828;
  assign n834 = ~n830 & ~n832;
  assign n835 = n833 & n834;
  assign n836 = n301 & ~n835;
  assign n837 = pi121  & ~pi128 ;
  assign n838 = ~pi129  & n837;
  assign n839 = pi118  & pi128 ;
  assign n840 = pi129  & n839;
  assign n841 = pi120  & pi128 ;
  assign n842 = ~pi129  & n841;
  assign n843 = pi119  & ~pi128 ;
  assign n844 = pi129  & n843;
  assign n845 = ~n838 & ~n840;
  assign n846 = ~n842 & ~n844;
  assign n847 = n845 & n846;
  assign n848 = n314 & ~n847;
  assign n849 = ~n812 & ~n824;
  assign n850 = ~n836 & ~n848;
  assign n851 = n849 & n850;
  assign n852 = n425 & ~n851;
  assign n853 = pi113  & ~pi128 ;
  assign n854 = ~pi129  & n853;
  assign n855 = pi110  & pi128 ;
  assign n856 = pi129  & n855;
  assign n857 = pi112  & pi128 ;
  assign n858 = ~pi129  & n857;
  assign n859 = pi111  & ~pi128 ;
  assign n860 = pi129  & n859;
  assign n861 = ~n854 & ~n856;
  assign n862 = ~n858 & ~n860;
  assign n863 = n861 & n862;
  assign n864 = n275 & ~n863;
  assign n865 = pi109  & ~pi128 ;
  assign n866 = ~pi129  & n865;
  assign n867 = pi106  & pi128 ;
  assign n868 = pi129  & n867;
  assign n869 = pi108  & pi128 ;
  assign n870 = ~pi129  & n869;
  assign n871 = pi107  & ~pi128 ;
  assign n872 = pi129  & n871;
  assign n873 = ~n866 & ~n868;
  assign n874 = ~n870 & ~n872;
  assign n875 = n873 & n874;
  assign n876 = n288 & ~n875;
  assign n877 = pi101  & ~pi128 ;
  assign n878 = ~pi129  & n877;
  assign n879 = pi98  & pi128 ;
  assign n880 = pi129  & n879;
  assign n881 = pi100  & pi128 ;
  assign n882 = ~pi129  & n881;
  assign n883 = pi99  & ~pi128 ;
  assign n884 = pi129  & n883;
  assign n885 = ~n878 & ~n880;
  assign n886 = ~n882 & ~n884;
  assign n887 = n885 & n886;
  assign n888 = n301 & ~n887;
  assign n889 = pi105  & ~pi128 ;
  assign n890 = ~pi129  & n889;
  assign n891 = pi102  & pi128 ;
  assign n892 = pi129  & n891;
  assign n893 = pi104  & pi128 ;
  assign n894 = ~pi129  & n893;
  assign n895 = pi103  & ~pi128 ;
  assign n896 = pi129  & n895;
  assign n897 = ~n890 & ~n892;
  assign n898 = ~n894 & ~n896;
  assign n899 = n897 & n898;
  assign n900 = n314 & ~n899;
  assign n901 = ~n864 & ~n876;
  assign n902 = ~n888 & ~n900;
  assign n903 = n901 & n902;
  assign n904 = n478 & ~n903;
  assign n905 = ~n748 & ~n800;
  assign n906 = ~n852 & ~n904;
  assign n907 = n905 & n906;
  assign n908 = ~pi134  & ~n907;
  assign n909 = pi65  & ~pi128 ;
  assign n910 = ~pi129  & n909;
  assign n911 = pi62  & pi128 ;
  assign n912 = pi129  & n911;
  assign n913 = pi64  & pi128 ;
  assign n914 = ~pi129  & n913;
  assign n915 = pi63  & ~pi128 ;
  assign n916 = pi129  & n915;
  assign n917 = ~n910 & ~n912;
  assign n918 = ~n914 & ~n916;
  assign n919 = n917 & n918;
  assign n920 = n275 & ~n919;
  assign n921 = pi61  & ~pi128 ;
  assign n922 = ~pi129  & n921;
  assign n923 = pi58  & pi128 ;
  assign n924 = pi129  & n923;
  assign n925 = pi60  & pi128 ;
  assign n926 = ~pi129  & n925;
  assign n927 = pi59  & ~pi128 ;
  assign n928 = pi129  & n927;
  assign n929 = ~n922 & ~n924;
  assign n930 = ~n926 & ~n928;
  assign n931 = n929 & n930;
  assign n932 = n288 & ~n931;
  assign n933 = pi53  & ~pi128 ;
  assign n934 = ~pi129  & n933;
  assign n935 = pi50  & pi128 ;
  assign n936 = pi129  & n935;
  assign n937 = pi52  & pi128 ;
  assign n938 = ~pi129  & n937;
  assign n939 = pi51  & ~pi128 ;
  assign n940 = pi129  & n939;
  assign n941 = ~n934 & ~n936;
  assign n942 = ~n938 & ~n940;
  assign n943 = n941 & n942;
  assign n944 = n301 & ~n943;
  assign n945 = pi57  & ~pi128 ;
  assign n946 = ~pi129  & n945;
  assign n947 = pi54  & pi128 ;
  assign n948 = pi129  & n947;
  assign n949 = pi56  & pi128 ;
  assign n950 = ~pi129  & n949;
  assign n951 = pi55  & ~pi128 ;
  assign n952 = pi129  & n951;
  assign n953 = ~n946 & ~n948;
  assign n954 = ~n950 & ~n952;
  assign n955 = n953 & n954;
  assign n956 = n314 & ~n955;
  assign n957 = ~n920 & ~n932;
  assign n958 = ~n944 & ~n956;
  assign n959 = n957 & n958;
  assign n960 = n425 & ~n959;
  assign n961 = pi17  & ~pi128 ;
  assign n962 = ~pi129  & n961;
  assign n963 = pi14  & pi128 ;
  assign n964 = pi129  & n963;
  assign n965 = pi16  & pi128 ;
  assign n966 = ~pi129  & n965;
  assign n967 = pi15  & ~pi128 ;
  assign n968 = pi129  & n967;
  assign n969 = ~n962 & ~n964;
  assign n970 = ~n966 & ~n968;
  assign n971 = n969 & n970;
  assign n972 = n275 & ~n971;
  assign n973 = pi13  & ~pi128 ;
  assign n974 = ~pi129  & n973;
  assign n975 = pi10  & pi128 ;
  assign n976 = pi129  & n975;
  assign n977 = pi12  & pi128 ;
  assign n978 = ~pi129  & n977;
  assign n979 = pi11  & ~pi128 ;
  assign n980 = pi129  & n979;
  assign n981 = ~n974 & ~n976;
  assign n982 = ~n978 & ~n980;
  assign n983 = n981 & n982;
  assign n984 = n288 & ~n983;
  assign n985 = pi5  & ~pi128 ;
  assign n986 = ~pi129  & n985;
  assign n987 = pi2  & pi128 ;
  assign n988 = pi129  & n987;
  assign n989 = pi4  & pi128 ;
  assign n990 = ~pi129  & n989;
  assign n991 = pi3  & ~pi128 ;
  assign n992 = pi129  & n991;
  assign n993 = ~n986 & ~n988;
  assign n994 = ~n990 & ~n992;
  assign n995 = n993 & n994;
  assign n996 = n301 & ~n995;
  assign n997 = pi9  & ~pi128 ;
  assign n998 = ~pi129  & n997;
  assign n999 = pi6  & pi128 ;
  assign n1000 = pi129  & n999;
  assign n1001 = pi8  & pi128 ;
  assign n1002 = ~pi129  & n1001;
  assign n1003 = pi7  & ~pi128 ;
  assign n1004 = pi129  & n1003;
  assign n1005 = ~n998 & ~n1000;
  assign n1006 = ~n1002 & ~n1004;
  assign n1007 = n1005 & n1006;
  assign n1008 = n314 & ~n1007;
  assign n1009 = ~n972 & ~n984;
  assign n1010 = ~n996 & ~n1008;
  assign n1011 = n1009 & n1010;
  assign n1012 = n319 & ~n1011;
  assign n1013 = pi49  & ~pi128 ;
  assign n1014 = ~pi129  & n1013;
  assign n1015 = pi46  & pi128 ;
  assign n1016 = pi129  & n1015;
  assign n1017 = pi48  & pi128 ;
  assign n1018 = ~pi129  & n1017;
  assign n1019 = pi47  & ~pi128 ;
  assign n1020 = pi129  & n1019;
  assign n1021 = ~n1014 & ~n1016;
  assign n1022 = ~n1018 & ~n1020;
  assign n1023 = n1021 & n1022;
  assign n1024 = n275 & ~n1023;
  assign n1025 = pi42  & pi128 ;
  assign n1026 = pi129  & n1025;
  assign n1027 = pi43  & ~pi128 ;
  assign n1028 = pi129  & n1027;
  assign n1029 = pi45  & ~pi128 ;
  assign n1030 = ~pi129  & n1029;
  assign n1031 = pi44  & pi128 ;
  assign n1032 = ~pi129  & n1031;
  assign n1033 = ~n1026 & ~n1028;
  assign n1034 = ~n1030 & ~n1032;
  assign n1035 = n1033 & n1034;
  assign n1036 = n288 & ~n1035;
  assign n1037 = pi37  & ~pi128 ;
  assign n1038 = ~pi129  & n1037;
  assign n1039 = pi34  & pi128 ;
  assign n1040 = pi129  & n1039;
  assign n1041 = pi36  & pi128 ;
  assign n1042 = ~pi129  & n1041;
  assign n1043 = pi35  & ~pi128 ;
  assign n1044 = pi129  & n1043;
  assign n1045 = ~n1038 & ~n1040;
  assign n1046 = ~n1042 & ~n1044;
  assign n1047 = n1045 & n1046;
  assign n1048 = n301 & ~n1047;
  assign n1049 = pi41  & ~pi128 ;
  assign n1050 = ~pi129  & n1049;
  assign n1051 = pi40  & pi128 ;
  assign n1052 = ~pi129  & n1051;
  assign n1053 = pi39  & ~pi128 ;
  assign n1054 = pi129  & n1053;
  assign n1055 = pi38  & pi128 ;
  assign n1056 = pi129  & n1055;
  assign n1057 = ~n1050 & ~n1052;
  assign n1058 = ~n1054 & ~n1056;
  assign n1059 = n1057 & n1058;
  assign n1060 = n314 & ~n1059;
  assign n1061 = ~n1024 & ~n1036;
  assign n1062 = ~n1048 & ~n1060;
  assign n1063 = n1061 & n1062;
  assign n1064 = n478 & ~n1063;
  assign n1065 = pi33  & ~pi128 ;
  assign n1066 = ~pi129  & n1065;
  assign n1067 = pi30  & pi128 ;
  assign n1068 = pi129  & n1067;
  assign n1069 = pi32  & pi128 ;
  assign n1070 = ~pi129  & n1069;
  assign n1071 = pi31  & ~pi128 ;
  assign n1072 = pi129  & n1071;
  assign n1073 = ~n1066 & ~n1068;
  assign n1074 = ~n1070 & ~n1072;
  assign n1075 = n1073 & n1074;
  assign n1076 = n275 & ~n1075;
  assign n1077 = pi29  & ~pi128 ;
  assign n1078 = ~pi129  & n1077;
  assign n1079 = pi26  & pi128 ;
  assign n1080 = pi129  & n1079;
  assign n1081 = pi28  & pi128 ;
  assign n1082 = ~pi129  & n1081;
  assign n1083 = pi27  & ~pi128 ;
  assign n1084 = pi129  & n1083;
  assign n1085 = ~n1078 & ~n1080;
  assign n1086 = ~n1082 & ~n1084;
  assign n1087 = n1085 & n1086;
  assign n1088 = n288 & ~n1087;
  assign n1089 = pi21  & ~pi128 ;
  assign n1090 = ~pi129  & n1089;
  assign n1091 = pi18  & pi128 ;
  assign n1092 = pi129  & n1091;
  assign n1093 = pi20  & pi128 ;
  assign n1094 = ~pi129  & n1093;
  assign n1095 = pi19  & ~pi128 ;
  assign n1096 = pi129  & n1095;
  assign n1097 = ~n1090 & ~n1092;
  assign n1098 = ~n1094 & ~n1096;
  assign n1099 = n1097 & n1098;
  assign n1100 = n301 & ~n1099;
  assign n1101 = pi25  & ~pi128 ;
  assign n1102 = ~pi129  & n1101;
  assign n1103 = pi22  & pi128 ;
  assign n1104 = pi129  & n1103;
  assign n1105 = pi24  & pi128 ;
  assign n1106 = ~pi129  & n1105;
  assign n1107 = pi23  & ~pi128 ;
  assign n1108 = pi129  & n1107;
  assign n1109 = ~n1102 & ~n1104;
  assign n1110 = ~n1106 & ~n1108;
  assign n1111 = n1109 & n1110;
  assign n1112 = n314 & ~n1111;
  assign n1113 = ~n1076 & ~n1088;
  assign n1114 = ~n1100 & ~n1112;
  assign n1115 = n1113 & n1114;
  assign n1116 = n372 & ~n1115;
  assign n1117 = ~n960 & ~n1012;
  assign n1118 = ~n1064 & ~n1116;
  assign n1119 = n1117 & n1118;
  assign n1120 = pi134  & ~n1119;
  assign po1  = n908 | n1120;
  assign n1122 = ~pi129  & n345;
  assign n1123 = ~pi129  & n347;
  assign n1124 = pi129  & n268;
  assign n1125 = pi129  & n270;
  assign n1126 = ~n1122 & ~n1123;
  assign n1127 = ~n1124 & ~n1125;
  assign n1128 = n1126 & n1127;
  assign n1129 = n275 & ~n1128;
  assign n1130 = ~pi129  & n264;
  assign n1131 = ~pi129  & n266;
  assign n1132 = pi129  & n281;
  assign n1133 = pi129  & n283;
  assign n1134 = ~n1130 & ~n1131;
  assign n1135 = ~n1132 & ~n1133;
  assign n1136 = n1134 & n1135;
  assign n1137 = n288 & ~n1136;
  assign n1138 = ~pi129  & n303;
  assign n1139 = ~pi129  & n305;
  assign n1140 = pi129  & n294;
  assign n1141 = pi129  & n296;
  assign n1142 = ~n1138 & ~n1139;
  assign n1143 = ~n1140 & ~n1141;
  assign n1144 = n1142 & n1143;
  assign n1145 = n301 & ~n1144;
  assign n1146 = ~pi129  & n277;
  assign n1147 = ~pi129  & n279;
  assign n1148 = pi129  & n307;
  assign n1149 = pi129  & n309;
  assign n1150 = ~n1146 & ~n1147;
  assign n1151 = ~n1148 & ~n1149;
  assign n1152 = n1150 & n1151;
  assign n1153 = n314 & ~n1152;
  assign n1154 = ~n1129 & ~n1137;
  assign n1155 = ~n1145 & ~n1153;
  assign n1156 = n1154 & n1155;
  assign n1157 = n319 & ~n1156;
  assign n1158 = ~pi129  & n451;
  assign n1159 = ~pi129  & n453;
  assign n1160 = pi129  & n325;
  assign n1161 = pi129  & n327;
  assign n1162 = ~n1158 & ~n1159;
  assign n1163 = ~n1160 & ~n1161;
  assign n1164 = n1162 & n1163;
  assign n1165 = n275 & ~n1164;
  assign n1166 = ~pi129  & n321;
  assign n1167 = ~pi129  & n323;
  assign n1168 = pi129  & n337;
  assign n1169 = pi129  & n339;
  assign n1170 = ~n1166 & ~n1167;
  assign n1171 = ~n1168 & ~n1169;
  assign n1172 = n1170 & n1171;
  assign n1173 = n288 & ~n1172;
  assign n1174 = ~pi129  & n357;
  assign n1175 = ~pi129  & n359;
  assign n1176 = pi129  & n349;
  assign n1177 = pi129  & n351;
  assign n1178 = ~n1174 & ~n1175;
  assign n1179 = ~n1176 & ~n1177;
  assign n1180 = n1178 & n1179;
  assign n1181 = n301 & ~n1180;
  assign n1182 = ~pi129  & n333;
  assign n1183 = ~pi129  & n335;
  assign n1184 = pi129  & n361;
  assign n1185 = pi129  & n363;
  assign n1186 = ~n1182 & ~n1183;
  assign n1187 = ~n1184 & ~n1185;
  assign n1188 = n1186 & n1187;
  assign n1189 = n314 & ~n1188;
  assign n1190 = ~n1165 & ~n1173;
  assign n1191 = ~n1181 & ~n1189;
  assign n1192 = n1190 & n1191;
  assign n1193 = n372 & ~n1192;
  assign n1194 = ~pi129  & n508;
  assign n1195 = ~pi129  & n510;
  assign n1196 = pi129  & n378;
  assign n1197 = pi129  & n380;
  assign n1198 = ~n1194 & ~n1195;
  assign n1199 = ~n1196 & ~n1197;
  assign n1200 = n1198 & n1199;
  assign n1201 = n275 & ~n1200;
  assign n1202 = ~pi129  & n374;
  assign n1203 = ~pi129  & n376;
  assign n1204 = pi129  & n390;
  assign n1205 = pi129  & n392;
  assign n1206 = ~n1202 & ~n1203;
  assign n1207 = ~n1204 & ~n1205;
  assign n1208 = n1206 & n1207;
  assign n1209 = n288 & ~n1208;
  assign n1210 = ~pi129  & n410;
  assign n1211 = ~pi129  & n412;
  assign n1212 = pi129  & n402;
  assign n1213 = pi129  & n404;
  assign n1214 = ~n1210 & ~n1211;
  assign n1215 = ~n1212 & ~n1213;
  assign n1216 = n1214 & n1215;
  assign n1217 = n301 & ~n1216;
  assign n1218 = ~pi129  & n386;
  assign n1219 = ~pi129  & n388;
  assign n1220 = pi129  & n414;
  assign n1221 = pi129  & n416;
  assign n1222 = ~n1218 & ~n1219;
  assign n1223 = ~n1220 & ~n1221;
  assign n1224 = n1222 & n1223;
  assign n1225 = n314 & ~n1224;
  assign n1226 = ~n1201 & ~n1209;
  assign n1227 = ~n1217 & ~n1225;
  assign n1228 = n1226 & n1227;
  assign n1229 = n425 & ~n1228;
  assign n1230 = ~pi129  & n398;
  assign n1231 = ~pi129  & n400;
  assign n1232 = pi129  & n431;
  assign n1233 = pi129  & n433;
  assign n1234 = ~n1230 & ~n1231;
  assign n1235 = ~n1232 & ~n1233;
  assign n1236 = n1234 & n1235;
  assign n1237 = n275 & ~n1236;
  assign n1238 = ~pi129  & n427;
  assign n1239 = ~pi129  & n429;
  assign n1240 = pi129  & n443;
  assign n1241 = pi129  & n445;
  assign n1242 = ~n1238 & ~n1239;
  assign n1243 = ~n1240 & ~n1241;
  assign n1244 = n1242 & n1243;
  assign n1245 = n288 & ~n1244;
  assign n1246 = ~pi129  & n463;
  assign n1247 = ~pi129  & n465;
  assign n1248 = pi129  & n455;
  assign n1249 = pi129  & n457;
  assign n1250 = ~n1246 & ~n1247;
  assign n1251 = ~n1248 & ~n1249;
  assign n1252 = n1250 & n1251;
  assign n1253 = n301 & ~n1252;
  assign n1254 = ~pi129  & n439;
  assign n1255 = ~pi129  & n441;
  assign n1256 = pi129  & n467;
  assign n1257 = pi129  & n469;
  assign n1258 = ~n1254 & ~n1255;
  assign n1259 = ~n1256 & ~n1257;
  assign n1260 = n1258 & n1259;
  assign n1261 = n314 & ~n1260;
  assign n1262 = ~n1237 & ~n1245;
  assign n1263 = ~n1253 & ~n1261;
  assign n1264 = n1262 & n1263;
  assign n1265 = n478 & ~n1264;
  assign n1266 = ~n1157 & ~n1193;
  assign n1267 = ~n1229 & ~n1265;
  assign n1268 = n1266 & n1267;
  assign n1269 = ~pi134  & ~n1268;
  assign n1270 = ~pi129  & n290;
  assign n1271 = ~pi129  & n292;
  assign n1272 = pi129  & n592;
  assign n1273 = pi129  & n594;
  assign n1274 = ~n1270 & ~n1271;
  assign n1275 = ~n1272 & ~n1273;
  assign n1276 = n1274 & n1275;
  assign n1277 = n275 & ~n1276;
  assign n1278 = ~pi129  & n588;
  assign n1279 = ~pi129  & n590;
  assign n1280 = pi129  & n604;
  assign n1281 = pi129  & n606;
  assign n1282 = ~n1278 & ~n1279;
  assign n1283 = ~n1280 & ~n1281;
  assign n1284 = n1282 & n1283;
  assign n1285 = n288 & ~n1284;
  assign n1286 = ~pi129  & n624;
  assign n1287 = ~pi129  & n626;
  assign n1288 = pi129  & n616;
  assign n1289 = pi129  & n618;
  assign n1290 = ~n1286 & ~n1287;
  assign n1291 = ~n1288 & ~n1289;
  assign n1292 = n1290 & n1291;
  assign n1293 = n301 & ~n1292;
  assign n1294 = ~pi129  & n600;
  assign n1295 = ~pi129  & n602;
  assign n1296 = pi129  & n628;
  assign n1297 = pi129  & n630;
  assign n1298 = ~n1294 & ~n1295;
  assign n1299 = ~n1296 & ~n1297;
  assign n1300 = n1298 & n1299;
  assign n1301 = n314 & ~n1300;
  assign n1302 = ~n1277 & ~n1285;
  assign n1303 = ~n1293 & ~n1301;
  assign n1304 = n1302 & n1303;
  assign n1305 = n425 & ~n1304;
  assign n1306 = ~pi129  & n560;
  assign n1307 = ~pi129  & n562;
  assign n1308 = pi129  & n488;
  assign n1309 = pi129  & n490;
  assign n1310 = ~n1306 & ~n1307;
  assign n1311 = ~n1308 & ~n1309;
  assign n1312 = n1310 & n1311;
  assign n1313 = n275 & ~n1312;
  assign n1314 = ~pi129  & n484;
  assign n1315 = ~pi129  & n486;
  assign n1316 = pi129  & n500;
  assign n1317 = pi129  & n502;
  assign n1318 = ~n1314 & ~n1315;
  assign n1319 = ~n1316 & ~n1317;
  assign n1320 = n1318 & n1319;
  assign n1321 = n288 & ~n1320;
  assign n1322 = ~pi129  & n520;
  assign n1323 = ~pi129  & n522;
  assign n1324 = pi129  & n512;
  assign n1325 = pi129  & n514;
  assign n1326 = ~n1322 & ~n1323;
  assign n1327 = ~n1324 & ~n1325;
  assign n1328 = n1326 & n1327;
  assign n1329 = n301 & ~n1328;
  assign n1330 = ~pi129  & n496;
  assign n1331 = ~pi129  & n498;
  assign n1332 = pi129  & n524;
  assign n1333 = pi129  & n526;
  assign n1334 = ~n1330 & ~n1331;
  assign n1335 = ~n1332 & ~n1333;
  assign n1336 = n1334 & n1335;
  assign n1337 = n314 & ~n1336;
  assign n1338 = ~n1313 & ~n1321;
  assign n1339 = ~n1329 & ~n1337;
  assign n1340 = n1338 & n1339;
  assign n1341 = n319 & ~n1340;
  assign n1342 = ~pi129  & n612;
  assign n1343 = ~pi129  & n614;
  assign n1344 = pi129  & n644;
  assign n1345 = pi129  & n646;
  assign n1346 = ~n1342 & ~n1343;
  assign n1347 = ~n1344 & ~n1345;
  assign n1348 = n1346 & n1347;
  assign n1349 = n275 & ~n1348;
  assign n1350 = pi129  & n658;
  assign n1351 = pi129  & n656;
  assign n1352 = ~pi129  & n642;
  assign n1353 = ~pi129  & n640;
  assign n1354 = ~n1350 & ~n1351;
  assign n1355 = ~n1352 & ~n1353;
  assign n1356 = n1354 & n1355;
  assign n1357 = n288 & ~n1356;
  assign n1358 = ~pi129  & n678;
  assign n1359 = ~pi129  & n682;
  assign n1360 = pi129  & n668;
  assign n1361 = pi129  & n670;
  assign n1362 = ~n1358 & ~n1359;
  assign n1363 = ~n1360 & ~n1361;
  assign n1364 = n1362 & n1363;
  assign n1365 = n301 & ~n1364;
  assign n1366 = ~pi129  & n652;
  assign n1367 = ~pi129  & n654;
  assign n1368 = pi129  & n680;
  assign n1369 = pi129  & n676;
  assign n1370 = ~n1366 & ~n1367;
  assign n1371 = ~n1368 & ~n1369;
  assign n1372 = n1370 & n1371;
  assign n1373 = n314 & ~n1372;
  assign n1374 = ~n1349 & ~n1357;
  assign n1375 = ~n1365 & ~n1373;
  assign n1376 = n1374 & n1375;
  assign n1377 = n478 & ~n1376;
  assign n1378 = ~pi129  & n664;
  assign n1379 = ~pi129  & n666;
  assign n1380 = pi129  & n540;
  assign n1381 = pi129  & n542;
  assign n1382 = ~n1378 & ~n1379;
  assign n1383 = ~n1380 & ~n1381;
  assign n1384 = n1382 & n1383;
  assign n1385 = n275 & ~n1384;
  assign n1386 = ~pi129  & n536;
  assign n1387 = ~pi129  & n538;
  assign n1388 = pi129  & n552;
  assign n1389 = pi129  & n554;
  assign n1390 = ~n1386 & ~n1387;
  assign n1391 = ~n1388 & ~n1389;
  assign n1392 = n1390 & n1391;
  assign n1393 = n288 & ~n1392;
  assign n1394 = ~pi129  & n572;
  assign n1395 = ~pi129  & n574;
  assign n1396 = pi129  & n564;
  assign n1397 = pi129  & n566;
  assign n1398 = ~n1394 & ~n1395;
  assign n1399 = ~n1396 & ~n1397;
  assign n1400 = n1398 & n1399;
  assign n1401 = n301 & ~n1400;
  assign n1402 = ~pi129  & n548;
  assign n1403 = ~pi129  & n550;
  assign n1404 = pi129  & n576;
  assign n1405 = pi129  & n578;
  assign n1406 = ~n1402 & ~n1403;
  assign n1407 = ~n1404 & ~n1405;
  assign n1408 = n1406 & n1407;
  assign n1409 = n314 & ~n1408;
  assign n1410 = ~n1385 & ~n1393;
  assign n1411 = ~n1401 & ~n1409;
  assign n1412 = n1410 & n1411;
  assign n1413 = n372 & ~n1412;
  assign n1414 = ~n1305 & ~n1341;
  assign n1415 = ~n1377 & ~n1413;
  assign n1416 = n1414 & n1415;
  assign n1417 = pi134  & ~n1416;
  assign po2  = n1269 | n1417;
  assign n1419 = pi129  & n853;
  assign n1420 = ~pi129  & n827;
  assign n1421 = pi129  & n857;
  assign n1422 = ~pi129  & n831;
  assign n1423 = ~n1419 & ~n1420;
  assign n1424 = ~n1421 & ~n1422;
  assign n1425 = n1423 & n1424;
  assign n1426 = n275 & ~n1425;
  assign n1427 = pi129  & n865;
  assign n1428 = ~pi129  & n855;
  assign n1429 = pi129  & n869;
  assign n1430 = ~pi129  & n859;
  assign n1431 = ~n1427 & ~n1428;
  assign n1432 = ~n1429 & ~n1430;
  assign n1433 = n1431 & n1432;
  assign n1434 = n288 & ~n1433;
  assign n1435 = pi129  & n877;
  assign n1436 = ~pi129  & n891;
  assign n1437 = pi129  & n881;
  assign n1438 = ~pi129  & n895;
  assign n1439 = ~n1435 & ~n1436;
  assign n1440 = ~n1437 & ~n1438;
  assign n1441 = n1439 & n1440;
  assign n1442 = n301 & ~n1441;
  assign n1443 = pi129  & n889;
  assign n1444 = ~pi129  & n867;
  assign n1445 = pi129  & n893;
  assign n1446 = ~pi129  & n871;
  assign n1447 = ~n1443 & ~n1444;
  assign n1448 = ~n1445 & ~n1446;
  assign n1449 = n1447 & n1448;
  assign n1450 = n314 & ~n1449;
  assign n1451 = ~n1426 & ~n1434;
  assign n1452 = ~n1442 & ~n1450;
  assign n1453 = n1451 & n1452;
  assign n1454 = n478 & ~n1453;
  assign n1455 = pi129  & n749;
  assign n1456 = ~pi129  & n879;
  assign n1457 = pi129  & n753;
  assign n1458 = ~pi129  & n883;
  assign n1459 = ~n1455 & ~n1456;
  assign n1460 = ~n1457 & ~n1458;
  assign n1461 = n1459 & n1460;
  assign n1462 = n275 & ~n1461;
  assign n1463 = pi129  & n761;
  assign n1464 = ~pi129  & n751;
  assign n1465 = pi129  & n765;
  assign n1466 = ~pi129  & n755;
  assign n1467 = ~n1463 & ~n1464;
  assign n1468 = ~n1465 & ~n1466;
  assign n1469 = n1467 & n1468;
  assign n1470 = n288 & ~n1469;
  assign n1471 = pi129  & n773;
  assign n1472 = ~pi129  & n787;
  assign n1473 = pi129  & n777;
  assign n1474 = ~pi129  & n791;
  assign n1475 = ~n1471 & ~n1472;
  assign n1476 = ~n1473 & ~n1474;
  assign n1477 = n1475 & n1476;
  assign n1478 = n301 & ~n1477;
  assign n1479 = pi129  & n785;
  assign n1480 = ~pi129  & n763;
  assign n1481 = pi129  & n789;
  assign n1482 = ~pi129  & n767;
  assign n1483 = ~n1479 & ~n1480;
  assign n1484 = ~n1481 & ~n1482;
  assign n1485 = n1483 & n1484;
  assign n1486 = n314 & ~n1485;
  assign n1487 = ~n1462 & ~n1470;
  assign n1488 = ~n1478 & ~n1486;
  assign n1489 = n1487 & n1488;
  assign n1490 = n372 & ~n1489;
  assign n1491 = pi129  & n801;
  assign n1492 = ~pi129  & n987;
  assign n1493 = pi129  & n805;
  assign n1494 = ~pi129  & n991;
  assign n1495 = ~n1491 & ~n1492;
  assign n1496 = ~n1493 & ~n1494;
  assign n1497 = n1495 & n1496;
  assign n1498 = n275 & ~n1497;
  assign n1499 = pi129  & n813;
  assign n1500 = ~pi129  & n803;
  assign n1501 = pi129  & n817;
  assign n1502 = ~pi129  & n807;
  assign n1503 = ~n1499 & ~n1500;
  assign n1504 = ~n1501 & ~n1502;
  assign n1505 = n1503 & n1504;
  assign n1506 = n288 & ~n1505;
  assign n1507 = pi129  & n825;
  assign n1508 = ~pi129  & n839;
  assign n1509 = pi129  & n829;
  assign n1510 = ~pi129  & n843;
  assign n1511 = ~n1507 & ~n1508;
  assign n1512 = ~n1509 & ~n1510;
  assign n1513 = n1511 & n1512;
  assign n1514 = n301 & ~n1513;
  assign n1515 = pi129  & n837;
  assign n1516 = ~pi129  & n815;
  assign n1517 = pi129  & n841;
  assign n1518 = ~pi129  & n819;
  assign n1519 = ~n1515 & ~n1516;
  assign n1520 = ~n1517 & ~n1518;
  assign n1521 = n1519 & n1520;
  assign n1522 = n314 & ~n1521;
  assign n1523 = ~n1498 & ~n1506;
  assign n1524 = ~n1514 & ~n1522;
  assign n1525 = n1523 & n1524;
  assign n1526 = n425 & ~n1525;
  assign n1527 = pi129  & n697;
  assign n1528 = ~pi129  & n775;
  assign n1529 = pi129  & n701;
  assign n1530 = ~pi129  & n779;
  assign n1531 = ~n1527 & ~n1528;
  assign n1532 = ~n1529 & ~n1530;
  assign n1533 = n1531 & n1532;
  assign n1534 = n275 & ~n1533;
  assign n1535 = pi129  & n709;
  assign n1536 = ~pi129  & n699;
  assign n1537 = pi129  & n713;
  assign n1538 = ~pi129  & n703;
  assign n1539 = ~n1535 & ~n1536;
  assign n1540 = ~n1537 & ~n1538;
  assign n1541 = n1539 & n1540;
  assign n1542 = n288 & ~n1541;
  assign n1543 = pi129  & n721;
  assign n1544 = ~pi129  & n735;
  assign n1545 = pi129  & n725;
  assign n1546 = ~pi129  & n739;
  assign n1547 = ~n1543 & ~n1544;
  assign n1548 = ~n1545 & ~n1546;
  assign n1549 = n1547 & n1548;
  assign n1550 = n301 & ~n1549;
  assign n1551 = pi129  & n733;
  assign n1552 = ~pi129  & n711;
  assign n1553 = pi129  & n737;
  assign n1554 = ~pi129  & n715;
  assign n1555 = ~n1551 & ~n1552;
  assign n1556 = ~n1553 & ~n1554;
  assign n1557 = n1555 & n1556;
  assign n1558 = n314 & ~n1557;
  assign n1559 = ~n1534 & ~n1542;
  assign n1560 = ~n1550 & ~n1558;
  assign n1561 = n1559 & n1560;
  assign n1562 = n319 & ~n1561;
  assign n1563 = ~n1454 & ~n1490;
  assign n1564 = ~n1526 & ~n1562;
  assign n1565 = n1563 & n1564;
  assign n1566 = ~pi134  & ~n1565;
  assign n1567 = pi129  & n909;
  assign n1568 = ~pi129  & n723;
  assign n1569 = pi129  & n913;
  assign n1570 = ~pi129  & n727;
  assign n1571 = ~n1567 & ~n1568;
  assign n1572 = ~n1569 & ~n1570;
  assign n1573 = n1571 & n1572;
  assign n1574 = n275 & ~n1573;
  assign n1575 = pi129  & n921;
  assign n1576 = ~pi129  & n911;
  assign n1577 = pi129  & n925;
  assign n1578 = ~pi129  & n915;
  assign n1579 = ~n1575 & ~n1576;
  assign n1580 = ~n1577 & ~n1578;
  assign n1581 = n1579 & n1580;
  assign n1582 = n288 & ~n1581;
  assign n1583 = pi129  & n933;
  assign n1584 = ~pi129  & n947;
  assign n1585 = pi129  & n937;
  assign n1586 = ~pi129  & n951;
  assign n1587 = ~n1583 & ~n1584;
  assign n1588 = ~n1585 & ~n1586;
  assign n1589 = n1587 & n1588;
  assign n1590 = n301 & ~n1589;
  assign n1591 = pi129  & n945;
  assign n1592 = ~pi129  & n923;
  assign n1593 = pi129  & n949;
  assign n1594 = ~pi129  & n927;
  assign n1595 = ~n1591 & ~n1592;
  assign n1596 = ~n1593 & ~n1594;
  assign n1597 = n1595 & n1596;
  assign n1598 = n314 & ~n1597;
  assign n1599 = ~n1574 & ~n1582;
  assign n1600 = ~n1590 & ~n1598;
  assign n1601 = n1599 & n1600;
  assign n1602 = n425 & ~n1601;
  assign n1603 = pi129  & n1013;
  assign n1604 = ~pi129  & n935;
  assign n1605 = pi129  & n1017;
  assign n1606 = ~pi129  & n939;
  assign n1607 = ~n1603 & ~n1604;
  assign n1608 = ~n1605 & ~n1606;
  assign n1609 = n1607 & n1608;
  assign n1610 = n275 & ~n1609;
  assign n1611 = pi129  & n1031;
  assign n1612 = pi129  & n1029;
  assign n1613 = ~pi129  & n1019;
  assign n1614 = ~pi129  & n1015;
  assign n1615 = ~n1611 & ~n1612;
  assign n1616 = ~n1613 & ~n1614;
  assign n1617 = n1615 & n1616;
  assign n1618 = n288 & ~n1617;
  assign n1619 = pi129  & n1037;
  assign n1620 = ~pi129  & n1055;
  assign n1621 = pi129  & n1041;
  assign n1622 = ~pi129  & n1053;
  assign n1623 = ~n1619 & ~n1620;
  assign n1624 = ~n1621 & ~n1622;
  assign n1625 = n1623 & n1624;
  assign n1626 = n301 & ~n1625;
  assign n1627 = pi129  & n1049;
  assign n1628 = ~pi129  & n1025;
  assign n1629 = pi129  & n1051;
  assign n1630 = ~pi129  & n1027;
  assign n1631 = ~n1627 & ~n1628;
  assign n1632 = ~n1629 & ~n1630;
  assign n1633 = n1631 & n1632;
  assign n1634 = n314 & ~n1633;
  assign n1635 = ~n1610 & ~n1618;
  assign n1636 = ~n1626 & ~n1634;
  assign n1637 = n1635 & n1636;
  assign n1638 = n478 & ~n1637;
  assign n1639 = pi129  & n961;
  assign n1640 = ~pi129  & n1091;
  assign n1641 = pi129  & n965;
  assign n1642 = ~pi129  & n1095;
  assign n1643 = ~n1639 & ~n1640;
  assign n1644 = ~n1641 & ~n1642;
  assign n1645 = n1643 & n1644;
  assign n1646 = n275 & ~n1645;
  assign n1647 = pi129  & n973;
  assign n1648 = ~pi129  & n963;
  assign n1649 = pi129  & n977;
  assign n1650 = ~pi129  & n967;
  assign n1651 = ~n1647 & ~n1648;
  assign n1652 = ~n1649 & ~n1650;
  assign n1653 = n1651 & n1652;
  assign n1654 = n288 & ~n1653;
  assign n1655 = pi129  & n985;
  assign n1656 = ~pi129  & n999;
  assign n1657 = pi129  & n989;
  assign n1658 = ~pi129  & n1003;
  assign n1659 = ~n1655 & ~n1656;
  assign n1660 = ~n1657 & ~n1658;
  assign n1661 = n1659 & n1660;
  assign n1662 = n301 & ~n1661;
  assign n1663 = pi129  & n997;
  assign n1664 = ~pi129  & n975;
  assign n1665 = pi129  & n1001;
  assign n1666 = ~pi129  & n979;
  assign n1667 = ~n1663 & ~n1664;
  assign n1668 = ~n1665 & ~n1666;
  assign n1669 = n1667 & n1668;
  assign n1670 = n314 & ~n1669;
  assign n1671 = ~n1646 & ~n1654;
  assign n1672 = ~n1662 & ~n1670;
  assign n1673 = n1671 & n1672;
  assign n1674 = n319 & ~n1673;
  assign n1675 = pi129  & n1065;
  assign n1676 = ~pi129  & n1039;
  assign n1677 = pi129  & n1069;
  assign n1678 = ~pi129  & n1043;
  assign n1679 = ~n1675 & ~n1676;
  assign n1680 = ~n1677 & ~n1678;
  assign n1681 = n1679 & n1680;
  assign n1682 = n275 & ~n1681;
  assign n1683 = pi129  & n1077;
  assign n1684 = ~pi129  & n1067;
  assign n1685 = pi129  & n1081;
  assign n1686 = ~pi129  & n1071;
  assign n1687 = ~n1683 & ~n1684;
  assign n1688 = ~n1685 & ~n1686;
  assign n1689 = n1687 & n1688;
  assign n1690 = n288 & ~n1689;
  assign n1691 = pi129  & n1089;
  assign n1692 = ~pi129  & n1103;
  assign n1693 = pi129  & n1093;
  assign n1694 = ~pi129  & n1107;
  assign n1695 = ~n1691 & ~n1692;
  assign n1696 = ~n1693 & ~n1694;
  assign n1697 = n1695 & n1696;
  assign n1698 = n301 & ~n1697;
  assign n1699 = pi129  & n1101;
  assign n1700 = ~pi129  & n1079;
  assign n1701 = pi129  & n1105;
  assign n1702 = ~pi129  & n1083;
  assign n1703 = ~n1699 & ~n1700;
  assign n1704 = ~n1701 & ~n1702;
  assign n1705 = n1703 & n1704;
  assign n1706 = n314 & ~n1705;
  assign n1707 = ~n1682 & ~n1690;
  assign n1708 = ~n1698 & ~n1706;
  assign n1709 = n1707 & n1708;
  assign n1710 = n372 & ~n1709;
  assign n1711 = ~n1602 & ~n1638;
  assign n1712 = ~n1674 & ~n1710;
  assign n1713 = n1711 & n1712;
  assign n1714 = pi134  & ~n1713;
  assign po3  = n1566 | n1714;
  assign n1716 = n275 & ~n355;
  assign n1717 = ~n274 & n288;
  assign n1718 = n301 & ~n313;
  assign n1719 = ~n287 & n314;
  assign n1720 = ~n1716 & ~n1717;
  assign n1721 = ~n1718 & ~n1719;
  assign n1722 = n1720 & n1721;
  assign n1723 = n319 & ~n1722;
  assign n1724 = n275 & ~n461;
  assign n1725 = n288 & ~n331;
  assign n1726 = n301 & ~n367;
  assign n1727 = n314 & ~n343;
  assign n1728 = ~n1724 & ~n1725;
  assign n1729 = ~n1726 & ~n1727;
  assign n1730 = n1728 & n1729;
  assign n1731 = n372 & ~n1730;
  assign n1732 = n275 & ~n518;
  assign n1733 = n288 & ~n384;
  assign n1734 = n301 & ~n420;
  assign n1735 = n314 & ~n396;
  assign n1736 = ~n1732 & ~n1733;
  assign n1737 = ~n1734 & ~n1735;
  assign n1738 = n1736 & n1737;
  assign n1739 = n425 & ~n1738;
  assign n1740 = n275 & ~n408;
  assign n1741 = n288 & ~n437;
  assign n1742 = n301 & ~n473;
  assign n1743 = n314 & ~n449;
  assign n1744 = ~n1740 & ~n1741;
  assign n1745 = ~n1742 & ~n1743;
  assign n1746 = n1744 & n1745;
  assign n1747 = n478 & ~n1746;
  assign n1748 = ~n1723 & ~n1731;
  assign n1749 = ~n1739 & ~n1747;
  assign n1750 = n1748 & n1749;
  assign n1751 = ~pi134  & ~n1750;
  assign n1752 = n275 & ~n622;
  assign n1753 = n288 & ~n650;
  assign n1754 = n301 & ~n686;
  assign n1755 = n314 & ~n662;
  assign n1756 = ~n1752 & ~n1753;
  assign n1757 = ~n1754 & ~n1755;
  assign n1758 = n1756 & n1757;
  assign n1759 = n478 & ~n1758;
  assign n1760 = n275 & ~n300;
  assign n1761 = n288 & ~n598;
  assign n1762 = n301 & ~n634;
  assign n1763 = n314 & ~n610;
  assign n1764 = ~n1760 & ~n1761;
  assign n1765 = ~n1762 & ~n1763;
  assign n1766 = n1764 & n1765;
  assign n1767 = n425 & ~n1766;
  assign n1768 = n275 & ~n674;
  assign n1769 = n288 & ~n546;
  assign n1770 = n301 & ~n582;
  assign n1771 = n314 & ~n558;
  assign n1772 = ~n1768 & ~n1769;
  assign n1773 = ~n1770 & ~n1771;
  assign n1774 = n1772 & n1773;
  assign n1775 = n372 & ~n1774;
  assign n1776 = n275 & ~n570;
  assign n1777 = n288 & ~n494;
  assign n1778 = n301 & ~n530;
  assign n1779 = n314 & ~n506;
  assign n1780 = ~n1776 & ~n1777;
  assign n1781 = ~n1778 & ~n1779;
  assign n1782 = n1780 & n1781;
  assign n1783 = n319 & ~n1782;
  assign n1784 = ~n1759 & ~n1767;
  assign n1785 = ~n1775 & ~n1783;
  assign n1786 = n1784 & n1785;
  assign n1787 = pi134  & ~n1786;
  assign po4  = n1751 | n1787;
  assign n1789 = n275 & ~n783;
  assign n1790 = n288 & ~n707;
  assign n1791 = n301 & ~n743;
  assign n1792 = n314 & ~n719;
  assign n1793 = ~n1789 & ~n1790;
  assign n1794 = ~n1791 & ~n1792;
  assign n1795 = n1793 & n1794;
  assign n1796 = n319 & ~n1795;
  assign n1797 = n275 & ~n887;
  assign n1798 = n288 & ~n759;
  assign n1799 = n301 & ~n795;
  assign n1800 = n314 & ~n771;
  assign n1801 = ~n1797 & ~n1798;
  assign n1802 = ~n1799 & ~n1800;
  assign n1803 = n1801 & n1802;
  assign n1804 = n372 & ~n1803;
  assign n1805 = n275 & ~n995;
  assign n1806 = n288 & ~n811;
  assign n1807 = n301 & ~n847;
  assign n1808 = n314 & ~n823;
  assign n1809 = ~n1805 & ~n1806;
  assign n1810 = ~n1807 & ~n1808;
  assign n1811 = n1809 & n1810;
  assign n1812 = n425 & ~n1811;
  assign n1813 = n275 & ~n835;
  assign n1814 = n288 & ~n863;
  assign n1815 = n301 & ~n899;
  assign n1816 = n314 & ~n875;
  assign n1817 = ~n1813 & ~n1814;
  assign n1818 = ~n1815 & ~n1816;
  assign n1819 = n1817 & n1818;
  assign n1820 = n478 & ~n1819;
  assign n1821 = ~n1796 & ~n1804;
  assign n1822 = ~n1812 & ~n1820;
  assign n1823 = n1821 & n1822;
  assign n1824 = ~pi134  & ~n1823;
  assign n1825 = n275 & ~n943;
  assign n1826 = n288 & ~n1023;
  assign n1827 = n301 & ~n1059;
  assign n1828 = n314 & ~n1035;
  assign n1829 = ~n1825 & ~n1826;
  assign n1830 = ~n1827 & ~n1828;
  assign n1831 = n1829 & n1830;
  assign n1832 = n478 & ~n1831;
  assign n1833 = n275 & ~n731;
  assign n1834 = n288 & ~n919;
  assign n1835 = n301 & ~n955;
  assign n1836 = n314 & ~n931;
  assign n1837 = ~n1833 & ~n1834;
  assign n1838 = ~n1835 & ~n1836;
  assign n1839 = n1837 & n1838;
  assign n1840 = n425 & ~n1839;
  assign n1841 = n275 & ~n1047;
  assign n1842 = n288 & ~n1075;
  assign n1843 = n301 & ~n1111;
  assign n1844 = n314 & ~n1087;
  assign n1845 = ~n1841 & ~n1842;
  assign n1846 = ~n1843 & ~n1844;
  assign n1847 = n1845 & n1846;
  assign n1848 = n372 & ~n1847;
  assign n1849 = n275 & ~n1099;
  assign n1850 = n288 & ~n971;
  assign n1851 = n301 & ~n1007;
  assign n1852 = n314 & ~n983;
  assign n1853 = ~n1849 & ~n1850;
  assign n1854 = ~n1851 & ~n1852;
  assign n1855 = n1853 & n1854;
  assign n1856 = n319 & ~n1855;
  assign n1857 = ~n1832 & ~n1840;
  assign n1858 = ~n1848 & ~n1856;
  assign n1859 = n1857 & n1858;
  assign n1860 = pi134  & ~n1859;
  assign po5  = n1824 | n1860;
  assign n1862 = n275 & ~n1180;
  assign n1863 = n288 & ~n1128;
  assign n1864 = n301 & ~n1152;
  assign n1865 = n314 & ~n1136;
  assign n1866 = ~n1862 & ~n1863;
  assign n1867 = ~n1864 & ~n1865;
  assign n1868 = n1866 & n1867;
  assign n1869 = n319 & ~n1868;
  assign n1870 = n275 & ~n1252;
  assign n1871 = n288 & ~n1164;
  assign n1872 = n301 & ~n1188;
  assign n1873 = n314 & ~n1172;
  assign n1874 = ~n1870 & ~n1871;
  assign n1875 = ~n1872 & ~n1873;
  assign n1876 = n1874 & n1875;
  assign n1877 = n372 & ~n1876;
  assign n1878 = n275 & ~n1328;
  assign n1879 = n288 & ~n1200;
  assign n1880 = n301 & ~n1224;
  assign n1881 = n314 & ~n1208;
  assign n1882 = ~n1878 & ~n1879;
  assign n1883 = ~n1880 & ~n1881;
  assign n1884 = n1882 & n1883;
  assign n1885 = n425 & ~n1884;
  assign n1886 = n275 & ~n1216;
  assign n1887 = n288 & ~n1236;
  assign n1888 = n301 & ~n1260;
  assign n1889 = n314 & ~n1244;
  assign n1890 = ~n1886 & ~n1887;
  assign n1891 = ~n1888 & ~n1889;
  assign n1892 = n1890 & n1891;
  assign n1893 = n478 & ~n1892;
  assign n1894 = ~n1869 & ~n1877;
  assign n1895 = ~n1885 & ~n1893;
  assign n1896 = n1894 & n1895;
  assign n1897 = ~pi134  & ~n1896;
  assign n1898 = n275 & ~n1292;
  assign n1899 = n288 & ~n1348;
  assign n1900 = n301 & ~n1372;
  assign n1901 = n314 & ~n1356;
  assign n1902 = ~n1898 & ~n1899;
  assign n1903 = ~n1900 & ~n1901;
  assign n1904 = n1902 & n1903;
  assign n1905 = n478 & ~n1904;
  assign n1906 = n275 & ~n1144;
  assign n1907 = n288 & ~n1276;
  assign n1908 = n301 & ~n1300;
  assign n1909 = n314 & ~n1284;
  assign n1910 = ~n1906 & ~n1907;
  assign n1911 = ~n1908 & ~n1909;
  assign n1912 = n1910 & n1911;
  assign n1913 = n425 & ~n1912;
  assign n1914 = n275 & ~n1364;
  assign n1915 = n288 & ~n1384;
  assign n1916 = n301 & ~n1408;
  assign n1917 = n314 & ~n1392;
  assign n1918 = ~n1914 & ~n1915;
  assign n1919 = ~n1916 & ~n1917;
  assign n1920 = n1918 & n1919;
  assign n1921 = n372 & ~n1920;
  assign n1922 = n275 & ~n1400;
  assign n1923 = n288 & ~n1312;
  assign n1924 = n301 & ~n1336;
  assign n1925 = n314 & ~n1320;
  assign n1926 = ~n1922 & ~n1923;
  assign n1927 = ~n1924 & ~n1925;
  assign n1928 = n1926 & n1927;
  assign n1929 = n319 & ~n1928;
  assign n1930 = ~n1905 & ~n1913;
  assign n1931 = ~n1921 & ~n1929;
  assign n1932 = n1930 & n1931;
  assign n1933 = pi134  & ~n1932;
  assign po6  = n1897 | n1933;
  assign n1935 = n275 & ~n1477;
  assign n1936 = n288 & ~n1533;
  assign n1937 = n301 & ~n1557;
  assign n1938 = n314 & ~n1541;
  assign n1939 = ~n1935 & ~n1936;
  assign n1940 = ~n1937 & ~n1938;
  assign n1941 = n1939 & n1940;
  assign n1942 = n319 & ~n1941;
  assign n1943 = n275 & ~n1441;
  assign n1944 = n288 & ~n1461;
  assign n1945 = n301 & ~n1485;
  assign n1946 = n314 & ~n1469;
  assign n1947 = ~n1943 & ~n1944;
  assign n1948 = ~n1945 & ~n1946;
  assign n1949 = n1947 & n1948;
  assign n1950 = n372 & ~n1949;
  assign n1951 = n275 & ~n1661;
  assign n1952 = n288 & ~n1497;
  assign n1953 = n301 & ~n1521;
  assign n1954 = n314 & ~n1505;
  assign n1955 = ~n1951 & ~n1952;
  assign n1956 = ~n1953 & ~n1954;
  assign n1957 = n1955 & n1956;
  assign n1958 = n425 & ~n1957;
  assign n1959 = n275 & ~n1513;
  assign n1960 = n288 & ~n1425;
  assign n1961 = n301 & ~n1449;
  assign n1962 = n314 & ~n1433;
  assign n1963 = ~n1959 & ~n1960;
  assign n1964 = ~n1961 & ~n1962;
  assign n1965 = n1963 & n1964;
  assign n1966 = n478 & ~n1965;
  assign n1967 = ~n1942 & ~n1950;
  assign n1968 = ~n1958 & ~n1966;
  assign n1969 = n1967 & n1968;
  assign n1970 = ~pi134  & ~n1969;
  assign n1971 = n288 & ~n1609;
  assign n1972 = n314 & ~n1617;
  assign n1973 = n301 & ~n1633;
  assign n1974 = n275 & ~n1589;
  assign n1975 = ~n1971 & ~n1972;
  assign n1976 = ~n1973 & ~n1974;
  assign n1977 = n1975 & n1976;
  assign n1978 = n478 & ~n1977;
  assign n1979 = n275 & ~n1549;
  assign n1980 = n288 & ~n1573;
  assign n1981 = n301 & ~n1597;
  assign n1982 = n314 & ~n1581;
  assign n1983 = ~n1979 & ~n1980;
  assign n1984 = ~n1981 & ~n1982;
  assign n1985 = n1983 & n1984;
  assign n1986 = n425 & ~n1985;
  assign n1987 = n275 & ~n1625;
  assign n1988 = n288 & ~n1681;
  assign n1989 = n301 & ~n1705;
  assign n1990 = n314 & ~n1689;
  assign n1991 = ~n1987 & ~n1988;
  assign n1992 = ~n1989 & ~n1990;
  assign n1993 = n1991 & n1992;
  assign n1994 = n372 & ~n1993;
  assign n1995 = n275 & ~n1697;
  assign n1996 = n288 & ~n1645;
  assign n1997 = n301 & ~n1669;
  assign n1998 = n314 & ~n1653;
  assign n1999 = ~n1995 & ~n1996;
  assign n2000 = ~n1997 & ~n1998;
  assign n2001 = n1999 & n2000;
  assign n2002 = n319 & ~n2001;
  assign n2003 = ~n1978 & ~n1986;
  assign n2004 = ~n1994 & ~n2002;
  assign n2005 = n2003 & n2004;
  assign n2006 = pi134  & ~n2005;
  assign po7  = n1970 | n2006;
  assign n2008 = n275 & ~n367;
  assign n2009 = n288 & ~n355;
  assign n2010 = ~n287 & n301;
  assign n2011 = ~n274 & n314;
  assign n2012 = ~n2008 & ~n2009;
  assign n2013 = ~n2010 & ~n2011;
  assign n2014 = n2012 & n2013;
  assign n2015 = n319 & ~n2014;
  assign n2016 = n275 & ~n473;
  assign n2017 = n288 & ~n461;
  assign n2018 = n301 & ~n343;
  assign n2019 = n314 & ~n331;
  assign n2020 = ~n2016 & ~n2017;
  assign n2021 = ~n2018 & ~n2019;
  assign n2022 = n2020 & n2021;
  assign n2023 = n372 & ~n2022;
  assign n2024 = n275 & ~n530;
  assign n2025 = n288 & ~n518;
  assign n2026 = n301 & ~n396;
  assign n2027 = n314 & ~n384;
  assign n2028 = ~n2024 & ~n2025;
  assign n2029 = ~n2026 & ~n2027;
  assign n2030 = n2028 & n2029;
  assign n2031 = n425 & ~n2030;
  assign n2032 = n275 & ~n420;
  assign n2033 = n288 & ~n408;
  assign n2034 = n301 & ~n449;
  assign n2035 = n314 & ~n437;
  assign n2036 = ~n2032 & ~n2033;
  assign n2037 = ~n2034 & ~n2035;
  assign n2038 = n2036 & n2037;
  assign n2039 = n478 & ~n2038;
  assign n2040 = ~n2015 & ~n2023;
  assign n2041 = ~n2031 & ~n2039;
  assign n2042 = n2040 & n2041;
  assign n2043 = ~pi134  & ~n2042;
  assign n2044 = n275 & ~n634;
  assign n2045 = n288 & ~n622;
  assign n2046 = n301 & ~n662;
  assign n2047 = n314 & ~n650;
  assign n2048 = ~n2044 & ~n2045;
  assign n2049 = ~n2046 & ~n2047;
  assign n2050 = n2048 & n2049;
  assign n2051 = n478 & ~n2050;
  assign n2052 = n275 & ~n313;
  assign n2053 = n288 & ~n300;
  assign n2054 = n301 & ~n610;
  assign n2055 = n314 & ~n598;
  assign n2056 = ~n2052 & ~n2053;
  assign n2057 = ~n2054 & ~n2055;
  assign n2058 = n2056 & n2057;
  assign n2059 = n425 & ~n2058;
  assign n2060 = n275 & ~n686;
  assign n2061 = n288 & ~n674;
  assign n2062 = n301 & ~n558;
  assign n2063 = n314 & ~n546;
  assign n2064 = ~n2060 & ~n2061;
  assign n2065 = ~n2062 & ~n2063;
  assign n2066 = n2064 & n2065;
  assign n2067 = n372 & ~n2066;
  assign n2068 = n275 & ~n582;
  assign n2069 = n288 & ~n570;
  assign n2070 = n301 & ~n506;
  assign n2071 = n314 & ~n494;
  assign n2072 = ~n2068 & ~n2069;
  assign n2073 = ~n2070 & ~n2071;
  assign n2074 = n2072 & n2073;
  assign n2075 = n319 & ~n2074;
  assign n2076 = ~n2051 & ~n2059;
  assign n2077 = ~n2067 & ~n2075;
  assign n2078 = n2076 & n2077;
  assign n2079 = pi134  & ~n2078;
  assign po8  = n2043 | n2079;
  assign n2081 = n275 & ~n795;
  assign n2082 = n288 & ~n783;
  assign n2083 = n301 & ~n719;
  assign n2084 = n314 & ~n707;
  assign n2085 = ~n2081 & ~n2082;
  assign n2086 = ~n2083 & ~n2084;
  assign n2087 = n2085 & n2086;
  assign n2088 = n319 & ~n2087;
  assign n2089 = n275 & ~n899;
  assign n2090 = n288 & ~n887;
  assign n2091 = n301 & ~n771;
  assign n2092 = n314 & ~n759;
  assign n2093 = ~n2089 & ~n2090;
  assign n2094 = ~n2091 & ~n2092;
  assign n2095 = n2093 & n2094;
  assign n2096 = n372 & ~n2095;
  assign n2097 = n275 & ~n1007;
  assign n2098 = n288 & ~n995;
  assign n2099 = n301 & ~n823;
  assign n2100 = n314 & ~n811;
  assign n2101 = ~n2097 & ~n2098;
  assign n2102 = ~n2099 & ~n2100;
  assign n2103 = n2101 & n2102;
  assign n2104 = n425 & ~n2103;
  assign n2105 = n275 & ~n847;
  assign n2106 = n288 & ~n835;
  assign n2107 = n301 & ~n875;
  assign n2108 = n314 & ~n863;
  assign n2109 = ~n2105 & ~n2106;
  assign n2110 = ~n2107 & ~n2108;
  assign n2111 = n2109 & n2110;
  assign n2112 = n478 & ~n2111;
  assign n2113 = ~n2088 & ~n2096;
  assign n2114 = ~n2104 & ~n2112;
  assign n2115 = n2113 & n2114;
  assign n2116 = ~pi134  & ~n2115;
  assign n2117 = n275 & ~n955;
  assign n2118 = n288 & ~n943;
  assign n2119 = n301 & ~n1035;
  assign n2120 = n314 & ~n1023;
  assign n2121 = ~n2117 & ~n2118;
  assign n2122 = ~n2119 & ~n2120;
  assign n2123 = n2121 & n2122;
  assign n2124 = n478 & ~n2123;
  assign n2125 = n275 & ~n743;
  assign n2126 = n288 & ~n731;
  assign n2127 = n301 & ~n931;
  assign n2128 = n314 & ~n919;
  assign n2129 = ~n2125 & ~n2126;
  assign n2130 = ~n2127 & ~n2128;
  assign n2131 = n2129 & n2130;
  assign n2132 = n425 & ~n2131;
  assign n2133 = n275 & ~n1059;
  assign n2134 = n288 & ~n1047;
  assign n2135 = n301 & ~n1087;
  assign n2136 = n314 & ~n1075;
  assign n2137 = ~n2133 & ~n2134;
  assign n2138 = ~n2135 & ~n2136;
  assign n2139 = n2137 & n2138;
  assign n2140 = n372 & ~n2139;
  assign n2141 = n275 & ~n1111;
  assign n2142 = n288 & ~n1099;
  assign n2143 = n301 & ~n983;
  assign n2144 = n314 & ~n971;
  assign n2145 = ~n2141 & ~n2142;
  assign n2146 = ~n2143 & ~n2144;
  assign n2147 = n2145 & n2146;
  assign n2148 = n319 & ~n2147;
  assign n2149 = ~n2124 & ~n2132;
  assign n2150 = ~n2140 & ~n2148;
  assign n2151 = n2149 & n2150;
  assign n2152 = pi134  & ~n2151;
  assign po9  = n2116 | n2152;
  assign n2154 = n275 & ~n1188;
  assign n2155 = n288 & ~n1180;
  assign n2156 = n301 & ~n1136;
  assign n2157 = n314 & ~n1128;
  assign n2158 = ~n2154 & ~n2155;
  assign n2159 = ~n2156 & ~n2157;
  assign n2160 = n2158 & n2159;
  assign n2161 = n319 & ~n2160;
  assign n2162 = n275 & ~n1260;
  assign n2163 = n288 & ~n1252;
  assign n2164 = n301 & ~n1172;
  assign n2165 = n314 & ~n1164;
  assign n2166 = ~n2162 & ~n2163;
  assign n2167 = ~n2164 & ~n2165;
  assign n2168 = n2166 & n2167;
  assign n2169 = n372 & ~n2168;
  assign n2170 = n275 & ~n1336;
  assign n2171 = n288 & ~n1328;
  assign n2172 = n301 & ~n1208;
  assign n2173 = n314 & ~n1200;
  assign n2174 = ~n2170 & ~n2171;
  assign n2175 = ~n2172 & ~n2173;
  assign n2176 = n2174 & n2175;
  assign n2177 = n425 & ~n2176;
  assign n2178 = n275 & ~n1224;
  assign n2179 = n288 & ~n1216;
  assign n2180 = n301 & ~n1244;
  assign n2181 = n314 & ~n1236;
  assign n2182 = ~n2178 & ~n2179;
  assign n2183 = ~n2180 & ~n2181;
  assign n2184 = n2182 & n2183;
  assign n2185 = n478 & ~n2184;
  assign n2186 = ~n2161 & ~n2169;
  assign n2187 = ~n2177 & ~n2185;
  assign n2188 = n2186 & n2187;
  assign n2189 = ~pi134  & ~n2188;
  assign n2190 = n275 & ~n1300;
  assign n2191 = n288 & ~n1292;
  assign n2192 = n301 & ~n1356;
  assign n2193 = n314 & ~n1348;
  assign n2194 = ~n2190 & ~n2191;
  assign n2195 = ~n2192 & ~n2193;
  assign n2196 = n2194 & n2195;
  assign n2197 = n478 & ~n2196;
  assign n2198 = n275 & ~n1152;
  assign n2199 = n288 & ~n1144;
  assign n2200 = n301 & ~n1284;
  assign n2201 = n314 & ~n1276;
  assign n2202 = ~n2198 & ~n2199;
  assign n2203 = ~n2200 & ~n2201;
  assign n2204 = n2202 & n2203;
  assign n2205 = n425 & ~n2204;
  assign n2206 = n275 & ~n1372;
  assign n2207 = n288 & ~n1364;
  assign n2208 = n301 & ~n1392;
  assign n2209 = n314 & ~n1384;
  assign n2210 = ~n2206 & ~n2207;
  assign n2211 = ~n2208 & ~n2209;
  assign n2212 = n2210 & n2211;
  assign n2213 = n372 & ~n2212;
  assign n2214 = n275 & ~n1408;
  assign n2215 = n288 & ~n1400;
  assign n2216 = n301 & ~n1320;
  assign n2217 = n314 & ~n1312;
  assign n2218 = ~n2214 & ~n2215;
  assign n2219 = ~n2216 & ~n2217;
  assign n2220 = n2218 & n2219;
  assign n2221 = n319 & ~n2220;
  assign n2222 = ~n2197 & ~n2205;
  assign n2223 = ~n2213 & ~n2221;
  assign n2224 = n2222 & n2223;
  assign n2225 = pi134  & ~n2224;
  assign po10  = n2189 | n2225;
  assign n2227 = n275 & ~n1485;
  assign n2228 = n288 & ~n1477;
  assign n2229 = n301 & ~n1541;
  assign n2230 = n314 & ~n1533;
  assign n2231 = ~n2227 & ~n2228;
  assign n2232 = ~n2229 & ~n2230;
  assign n2233 = n2231 & n2232;
  assign n2234 = n319 & ~n2233;
  assign n2235 = n275 & ~n1449;
  assign n2236 = n288 & ~n1441;
  assign n2237 = n301 & ~n1469;
  assign n2238 = n314 & ~n1461;
  assign n2239 = ~n2235 & ~n2236;
  assign n2240 = ~n2237 & ~n2238;
  assign n2241 = n2239 & n2240;
  assign n2242 = n372 & ~n2241;
  assign n2243 = n275 & ~n1669;
  assign n2244 = n288 & ~n1661;
  assign n2245 = n301 & ~n1505;
  assign n2246 = n314 & ~n1497;
  assign n2247 = ~n2243 & ~n2244;
  assign n2248 = ~n2245 & ~n2246;
  assign n2249 = n2247 & n2248;
  assign n2250 = n425 & ~n2249;
  assign n2251 = n275 & ~n1521;
  assign n2252 = n288 & ~n1513;
  assign n2253 = n301 & ~n1433;
  assign n2254 = n314 & ~n1425;
  assign n2255 = ~n2251 & ~n2252;
  assign n2256 = ~n2253 & ~n2254;
  assign n2257 = n2255 & n2256;
  assign n2258 = n478 & ~n2257;
  assign n2259 = ~n2234 & ~n2242;
  assign n2260 = ~n2250 & ~n2258;
  assign n2261 = n2259 & n2260;
  assign n2262 = ~pi134  & ~n2261;
  assign n2263 = n275 & ~n1597;
  assign n2264 = n314 & ~n1609;
  assign n2265 = n301 & ~n1617;
  assign n2266 = n288 & ~n1589;
  assign n2267 = ~n2263 & ~n2264;
  assign n2268 = ~n2265 & ~n2266;
  assign n2269 = n2267 & n2268;
  assign n2270 = n478 & ~n2269;
  assign n2271 = n275 & ~n1557;
  assign n2272 = n288 & ~n1549;
  assign n2273 = n301 & ~n1581;
  assign n2274 = n314 & ~n1573;
  assign n2275 = ~n2271 & ~n2272;
  assign n2276 = ~n2273 & ~n2274;
  assign n2277 = n2275 & n2276;
  assign n2278 = n425 & ~n2277;
  assign n2279 = n275 & ~n1633;
  assign n2280 = n288 & ~n1625;
  assign n2281 = n301 & ~n1689;
  assign n2282 = n314 & ~n1681;
  assign n2283 = ~n2279 & ~n2280;
  assign n2284 = ~n2281 & ~n2282;
  assign n2285 = n2283 & n2284;
  assign n2286 = n372 & ~n2285;
  assign n2287 = n275 & ~n1705;
  assign n2288 = n288 & ~n1697;
  assign n2289 = n301 & ~n1653;
  assign n2290 = n314 & ~n1645;
  assign n2291 = ~n2287 & ~n2288;
  assign n2292 = ~n2289 & ~n2290;
  assign n2293 = n2291 & n2292;
  assign n2294 = n319 & ~n2293;
  assign n2295 = ~n2270 & ~n2278;
  assign n2296 = ~n2286 & ~n2294;
  assign n2297 = n2295 & n2296;
  assign n2298 = pi134  & ~n2297;
  assign po11  = n2262 | n2298;
  assign n2300 = n275 & ~n343;
  assign n2301 = n288 & ~n367;
  assign n2302 = ~n274 & n301;
  assign n2303 = n314 & ~n355;
  assign n2304 = ~n2300 & ~n2301;
  assign n2305 = ~n2302 & ~n2303;
  assign n2306 = n2304 & n2305;
  assign n2307 = n319 & ~n2306;
  assign n2308 = n275 & ~n449;
  assign n2309 = n288 & ~n473;
  assign n2310 = n301 & ~n331;
  assign n2311 = n314 & ~n461;
  assign n2312 = ~n2308 & ~n2309;
  assign n2313 = ~n2310 & ~n2311;
  assign n2314 = n2312 & n2313;
  assign n2315 = n372 & ~n2314;
  assign n2316 = n275 & ~n506;
  assign n2317 = n288 & ~n530;
  assign n2318 = n301 & ~n384;
  assign n2319 = n314 & ~n518;
  assign n2320 = ~n2316 & ~n2317;
  assign n2321 = ~n2318 & ~n2319;
  assign n2322 = n2320 & n2321;
  assign n2323 = n425 & ~n2322;
  assign n2324 = n275 & ~n396;
  assign n2325 = n288 & ~n420;
  assign n2326 = n301 & ~n437;
  assign n2327 = n314 & ~n408;
  assign n2328 = ~n2324 & ~n2325;
  assign n2329 = ~n2326 & ~n2327;
  assign n2330 = n2328 & n2329;
  assign n2331 = n478 & ~n2330;
  assign n2332 = ~n2307 & ~n2315;
  assign n2333 = ~n2323 & ~n2331;
  assign n2334 = n2332 & n2333;
  assign n2335 = ~pi134  & ~n2334;
  assign n2336 = n275 & ~n610;
  assign n2337 = n288 & ~n634;
  assign n2338 = n301 & ~n650;
  assign n2339 = n314 & ~n622;
  assign n2340 = ~n2336 & ~n2337;
  assign n2341 = ~n2338 & ~n2339;
  assign n2342 = n2340 & n2341;
  assign n2343 = n478 & ~n2342;
  assign n2344 = n275 & ~n287;
  assign n2345 = n288 & ~n313;
  assign n2346 = n301 & ~n598;
  assign n2347 = ~n300 & n314;
  assign n2348 = ~n2344 & ~n2345;
  assign n2349 = ~n2346 & ~n2347;
  assign n2350 = n2348 & n2349;
  assign n2351 = n425 & ~n2350;
  assign n2352 = n275 & ~n662;
  assign n2353 = n288 & ~n686;
  assign n2354 = n301 & ~n546;
  assign n2355 = n314 & ~n674;
  assign n2356 = ~n2352 & ~n2353;
  assign n2357 = ~n2354 & ~n2355;
  assign n2358 = n2356 & n2357;
  assign n2359 = n372 & ~n2358;
  assign n2360 = n275 & ~n558;
  assign n2361 = n288 & ~n582;
  assign n2362 = n301 & ~n494;
  assign n2363 = n314 & ~n570;
  assign n2364 = ~n2360 & ~n2361;
  assign n2365 = ~n2362 & ~n2363;
  assign n2366 = n2364 & n2365;
  assign n2367 = n319 & ~n2366;
  assign n2368 = ~n2343 & ~n2351;
  assign n2369 = ~n2359 & ~n2367;
  assign n2370 = n2368 & n2369;
  assign n2371 = pi134  & ~n2370;
  assign po12  = n2335 | n2371;
  assign n2373 = n275 & ~n771;
  assign n2374 = n288 & ~n795;
  assign n2375 = n301 & ~n707;
  assign n2376 = n314 & ~n783;
  assign n2377 = ~n2373 & ~n2374;
  assign n2378 = ~n2375 & ~n2376;
  assign n2379 = n2377 & n2378;
  assign n2380 = n319 & ~n2379;
  assign n2381 = n275 & ~n875;
  assign n2382 = n288 & ~n899;
  assign n2383 = n301 & ~n759;
  assign n2384 = n314 & ~n887;
  assign n2385 = ~n2381 & ~n2382;
  assign n2386 = ~n2383 & ~n2384;
  assign n2387 = n2385 & n2386;
  assign n2388 = n372 & ~n2387;
  assign n2389 = n275 & ~n983;
  assign n2390 = n288 & ~n1007;
  assign n2391 = n301 & ~n811;
  assign n2392 = n314 & ~n995;
  assign n2393 = ~n2389 & ~n2390;
  assign n2394 = ~n2391 & ~n2392;
  assign n2395 = n2393 & n2394;
  assign n2396 = n425 & ~n2395;
  assign n2397 = n275 & ~n823;
  assign n2398 = n288 & ~n847;
  assign n2399 = n301 & ~n863;
  assign n2400 = n314 & ~n835;
  assign n2401 = ~n2397 & ~n2398;
  assign n2402 = ~n2399 & ~n2400;
  assign n2403 = n2401 & n2402;
  assign n2404 = n478 & ~n2403;
  assign n2405 = ~n2380 & ~n2388;
  assign n2406 = ~n2396 & ~n2404;
  assign n2407 = n2405 & n2406;
  assign n2408 = ~pi134  & ~n2407;
  assign n2409 = n275 & ~n931;
  assign n2410 = n288 & ~n955;
  assign n2411 = n301 & ~n1023;
  assign n2412 = n314 & ~n943;
  assign n2413 = ~n2409 & ~n2410;
  assign n2414 = ~n2411 & ~n2412;
  assign n2415 = n2413 & n2414;
  assign n2416 = n478 & ~n2415;
  assign n2417 = n275 & ~n719;
  assign n2418 = n288 & ~n743;
  assign n2419 = n301 & ~n919;
  assign n2420 = n314 & ~n731;
  assign n2421 = ~n2417 & ~n2418;
  assign n2422 = ~n2419 & ~n2420;
  assign n2423 = n2421 & n2422;
  assign n2424 = n425 & ~n2423;
  assign n2425 = n275 & ~n1035;
  assign n2426 = n288 & ~n1059;
  assign n2427 = n301 & ~n1075;
  assign n2428 = n314 & ~n1047;
  assign n2429 = ~n2425 & ~n2426;
  assign n2430 = ~n2427 & ~n2428;
  assign n2431 = n2429 & n2430;
  assign n2432 = n372 & ~n2431;
  assign n2433 = n275 & ~n1087;
  assign n2434 = n288 & ~n1111;
  assign n2435 = n301 & ~n971;
  assign n2436 = n314 & ~n1099;
  assign n2437 = ~n2433 & ~n2434;
  assign n2438 = ~n2435 & ~n2436;
  assign n2439 = n2437 & n2438;
  assign n2440 = n319 & ~n2439;
  assign n2441 = ~n2416 & ~n2424;
  assign n2442 = ~n2432 & ~n2440;
  assign n2443 = n2441 & n2442;
  assign n2444 = pi134  & ~n2443;
  assign po13  = n2408 | n2444;
  assign n2446 = n275 & ~n1172;
  assign n2447 = n288 & ~n1188;
  assign n2448 = n301 & ~n1128;
  assign n2449 = n314 & ~n1180;
  assign n2450 = ~n2446 & ~n2447;
  assign n2451 = ~n2448 & ~n2449;
  assign n2452 = n2450 & n2451;
  assign n2453 = n319 & ~n2452;
  assign n2454 = n275 & ~n1244;
  assign n2455 = n288 & ~n1260;
  assign n2456 = n301 & ~n1164;
  assign n2457 = n314 & ~n1252;
  assign n2458 = ~n2454 & ~n2455;
  assign n2459 = ~n2456 & ~n2457;
  assign n2460 = n2458 & n2459;
  assign n2461 = n372 & ~n2460;
  assign n2462 = n275 & ~n1320;
  assign n2463 = n288 & ~n1336;
  assign n2464 = n301 & ~n1200;
  assign n2465 = n314 & ~n1328;
  assign n2466 = ~n2462 & ~n2463;
  assign n2467 = ~n2464 & ~n2465;
  assign n2468 = n2466 & n2467;
  assign n2469 = n425 & ~n2468;
  assign n2470 = n275 & ~n1208;
  assign n2471 = n288 & ~n1224;
  assign n2472 = n301 & ~n1236;
  assign n2473 = n314 & ~n1216;
  assign n2474 = ~n2470 & ~n2471;
  assign n2475 = ~n2472 & ~n2473;
  assign n2476 = n2474 & n2475;
  assign n2477 = n478 & ~n2476;
  assign n2478 = ~n2453 & ~n2461;
  assign n2479 = ~n2469 & ~n2477;
  assign n2480 = n2478 & n2479;
  assign n2481 = ~pi134  & ~n2480;
  assign n2482 = n275 & ~n1284;
  assign n2483 = n288 & ~n1300;
  assign n2484 = n301 & ~n1348;
  assign n2485 = n314 & ~n1292;
  assign n2486 = ~n2482 & ~n2483;
  assign n2487 = ~n2484 & ~n2485;
  assign n2488 = n2486 & n2487;
  assign n2489 = n478 & ~n2488;
  assign n2490 = n275 & ~n1136;
  assign n2491 = n288 & ~n1152;
  assign n2492 = n301 & ~n1276;
  assign n2493 = n314 & ~n1144;
  assign n2494 = ~n2490 & ~n2491;
  assign n2495 = ~n2492 & ~n2493;
  assign n2496 = n2494 & n2495;
  assign n2497 = n425 & ~n2496;
  assign n2498 = n275 & ~n1356;
  assign n2499 = n288 & ~n1372;
  assign n2500 = n301 & ~n1384;
  assign n2501 = n314 & ~n1364;
  assign n2502 = ~n2498 & ~n2499;
  assign n2503 = ~n2500 & ~n2501;
  assign n2504 = n2502 & n2503;
  assign n2505 = n372 & ~n2504;
  assign n2506 = n275 & ~n1392;
  assign n2507 = n288 & ~n1408;
  assign n2508 = n301 & ~n1312;
  assign n2509 = n314 & ~n1400;
  assign n2510 = ~n2506 & ~n2507;
  assign n2511 = ~n2508 & ~n2509;
  assign n2512 = n2510 & n2511;
  assign n2513 = n319 & ~n2512;
  assign n2514 = ~n2489 & ~n2497;
  assign n2515 = ~n2505 & ~n2513;
  assign n2516 = n2514 & n2515;
  assign n2517 = pi134  & ~n2516;
  assign po14  = n2481 | n2517;
  assign n2519 = n275 & ~n1469;
  assign n2520 = n288 & ~n1485;
  assign n2521 = n301 & ~n1533;
  assign n2522 = n314 & ~n1477;
  assign n2523 = ~n2519 & ~n2520;
  assign n2524 = ~n2521 & ~n2522;
  assign n2525 = n2523 & n2524;
  assign n2526 = n319 & ~n2525;
  assign n2527 = n275 & ~n1433;
  assign n2528 = n288 & ~n1449;
  assign n2529 = n301 & ~n1461;
  assign n2530 = n314 & ~n1441;
  assign n2531 = ~n2527 & ~n2528;
  assign n2532 = ~n2529 & ~n2530;
  assign n2533 = n2531 & n2532;
  assign n2534 = n372 & ~n2533;
  assign n2535 = n275 & ~n1653;
  assign n2536 = n288 & ~n1669;
  assign n2537 = n301 & ~n1497;
  assign n2538 = n314 & ~n1661;
  assign n2539 = ~n2535 & ~n2536;
  assign n2540 = ~n2537 & ~n2538;
  assign n2541 = n2539 & n2540;
  assign n2542 = n425 & ~n2541;
  assign n2543 = n275 & ~n1505;
  assign n2544 = n288 & ~n1521;
  assign n2545 = n301 & ~n1425;
  assign n2546 = n314 & ~n1513;
  assign n2547 = ~n2543 & ~n2544;
  assign n2548 = ~n2545 & ~n2546;
  assign n2549 = n2547 & n2548;
  assign n2550 = n478 & ~n2549;
  assign n2551 = ~n2526 & ~n2534;
  assign n2552 = ~n2542 & ~n2550;
  assign n2553 = n2551 & n2552;
  assign n2554 = ~pi134  & ~n2553;
  assign n2555 = n275 & ~n1581;
  assign n2556 = n288 & ~n1597;
  assign n2557 = n301 & ~n1609;
  assign n2558 = n314 & ~n1589;
  assign n2559 = ~n2555 & ~n2556;
  assign n2560 = ~n2557 & ~n2558;
  assign n2561 = n2559 & n2560;
  assign n2562 = n478 & ~n2561;
  assign n2563 = n275 & ~n1541;
  assign n2564 = n288 & ~n1557;
  assign n2565 = n301 & ~n1573;
  assign n2566 = n314 & ~n1549;
  assign n2567 = ~n2563 & ~n2564;
  assign n2568 = ~n2565 & ~n2566;
  assign n2569 = n2567 & n2568;
  assign n2570 = n425 & ~n2569;
  assign n2571 = n275 & ~n1617;
  assign n2572 = n288 & ~n1633;
  assign n2573 = n301 & ~n1681;
  assign n2574 = n314 & ~n1625;
  assign n2575 = ~n2571 & ~n2572;
  assign n2576 = ~n2573 & ~n2574;
  assign n2577 = n2575 & n2576;
  assign n2578 = n372 & ~n2577;
  assign n2579 = n275 & ~n1689;
  assign n2580 = n288 & ~n1705;
  assign n2581 = n301 & ~n1645;
  assign n2582 = n314 & ~n1697;
  assign n2583 = ~n2579 & ~n2580;
  assign n2584 = ~n2581 & ~n2582;
  assign n2585 = n2583 & n2584;
  assign n2586 = n319 & ~n2585;
  assign n2587 = ~n2562 & ~n2570;
  assign n2588 = ~n2578 & ~n2586;
  assign n2589 = n2587 & n2588;
  assign n2590 = pi134  & ~n2589;
  assign po15  = n2554 | n2590;
  assign n2592 = n319 & ~n371;
  assign n2593 = n372 & ~n477;
  assign n2594 = n425 & ~n534;
  assign n2595 = ~n424 & n478;
  assign n2596 = ~n2592 & ~n2593;
  assign n2597 = ~n2594 & ~n2595;
  assign n2598 = n2596 & n2597;
  assign n2599 = ~pi134  & ~n2598;
  assign n2600 = ~n318 & n425;
  assign n2601 = n319 & ~n586;
  assign n2602 = n478 & ~n638;
  assign n2603 = n372 & ~n690;
  assign n2604 = ~n2600 & ~n2601;
  assign n2605 = ~n2602 & ~n2603;
  assign n2606 = n2604 & n2605;
  assign n2607 = pi134  & ~n2606;
  assign po16  = n2599 | n2607;
  assign n2609 = n319 & ~n799;
  assign n2610 = n372 & ~n903;
  assign n2611 = n425 & ~n1011;
  assign n2612 = n478 & ~n851;
  assign n2613 = ~n2609 & ~n2610;
  assign n2614 = ~n2611 & ~n2612;
  assign n2615 = n2613 & n2614;
  assign n2616 = ~pi134  & ~n2615;
  assign n2617 = n478 & ~n959;
  assign n2618 = n425 & ~n747;
  assign n2619 = n372 & ~n1063;
  assign n2620 = n319 & ~n1115;
  assign n2621 = ~n2617 & ~n2618;
  assign n2622 = ~n2619 & ~n2620;
  assign n2623 = n2621 & n2622;
  assign n2624 = pi134  & ~n2623;
  assign po17  = n2616 | n2624;
  assign n2626 = n319 & ~n1192;
  assign n2627 = n372 & ~n1264;
  assign n2628 = n425 & ~n1340;
  assign n2629 = n478 & ~n1228;
  assign n2630 = ~n2626 & ~n2627;
  assign n2631 = ~n2628 & ~n2629;
  assign n2632 = n2630 & n2631;
  assign n2633 = ~pi134  & ~n2632;
  assign n2634 = n478 & ~n1304;
  assign n2635 = n425 & ~n1156;
  assign n2636 = n372 & ~n1376;
  assign n2637 = n319 & ~n1412;
  assign n2638 = ~n2634 & ~n2635;
  assign n2639 = ~n2636 & ~n2637;
  assign n2640 = n2638 & n2639;
  assign n2641 = pi134  & ~n2640;
  assign po18  = n2633 | n2641;
  assign n2643 = n372 & ~n1453;
  assign n2644 = n319 & ~n1489;
  assign n2645 = n478 & ~n1525;
  assign n2646 = n425 & ~n1673;
  assign n2647 = ~n2643 & ~n2644;
  assign n2648 = ~n2645 & ~n2646;
  assign n2649 = n2647 & n2648;
  assign n2650 = ~pi134  & ~n2649;
  assign n2651 = n478 & ~n1601;
  assign n2652 = n425 & ~n1561;
  assign n2653 = n319 & ~n1709;
  assign n2654 = n372 & ~n1637;
  assign n2655 = ~n2651 & ~n2652;
  assign n2656 = ~n2653 & ~n2654;
  assign n2657 = n2655 & n2656;
  assign n2658 = pi134  & ~n2657;
  assign po19  = n2650 | n2658;
  assign n2660 = n319 & ~n1730;
  assign n2661 = n372 & ~n1746;
  assign n2662 = n425 & ~n1782;
  assign n2663 = n478 & ~n1738;
  assign n2664 = ~n2660 & ~n2661;
  assign n2665 = ~n2662 & ~n2663;
  assign n2666 = n2664 & n2665;
  assign n2667 = ~pi134  & ~n2666;
  assign n2668 = n425 & ~n1722;
  assign n2669 = n372 & ~n1758;
  assign n2670 = n319 & ~n1774;
  assign n2671 = n478 & ~n1766;
  assign n2672 = ~n2668 & ~n2669;
  assign n2673 = ~n2670 & ~n2671;
  assign n2674 = n2672 & n2673;
  assign n2675 = pi134  & ~n2674;
  assign po20  = n2667 | n2675;
  assign n2677 = n319 & ~n1803;
  assign n2678 = n372 & ~n1819;
  assign n2679 = n425 & ~n1855;
  assign n2680 = n478 & ~n1811;
  assign n2681 = ~n2677 & ~n2678;
  assign n2682 = ~n2679 & ~n2680;
  assign n2683 = n2681 & n2682;
  assign n2684 = ~pi134  & ~n2683;
  assign n2685 = n425 & ~n1795;
  assign n2686 = n372 & ~n1831;
  assign n2687 = n319 & ~n1847;
  assign n2688 = n478 & ~n1839;
  assign n2689 = ~n2685 & ~n2686;
  assign n2690 = ~n2687 & ~n2688;
  assign n2691 = n2689 & n2690;
  assign n2692 = pi134  & ~n2691;
  assign po21  = n2684 | n2692;
  assign n2694 = n319 & ~n1876;
  assign n2695 = n372 & ~n1892;
  assign n2696 = n425 & ~n1928;
  assign n2697 = n478 & ~n1884;
  assign n2698 = ~n2694 & ~n2695;
  assign n2699 = ~n2696 & ~n2697;
  assign n2700 = n2698 & n2699;
  assign n2701 = ~pi134  & ~n2700;
  assign n2702 = n425 & ~n1868;
  assign n2703 = n372 & ~n1904;
  assign n2704 = n319 & ~n1920;
  assign n2705 = n478 & ~n1912;
  assign n2706 = ~n2702 & ~n2703;
  assign n2707 = ~n2704 & ~n2705;
  assign n2708 = n2706 & n2707;
  assign n2709 = pi134  & ~n2708;
  assign po22  = n2701 | n2709;
  assign n2711 = n319 & ~n1949;
  assign n2712 = n425 & ~n2001;
  assign n2713 = n478 & ~n1957;
  assign n2714 = n372 & ~n1965;
  assign n2715 = ~n2711 & ~n2712;
  assign n2716 = ~n2713 & ~n2714;
  assign n2717 = n2715 & n2716;
  assign n2718 = ~pi134  & ~n2717;
  assign n2719 = n372 & ~n1977;
  assign n2720 = n478 & ~n1985;
  assign n2721 = n319 & ~n1993;
  assign n2722 = n425 & ~n1941;
  assign n2723 = ~n2719 & ~n2720;
  assign n2724 = ~n2721 & ~n2722;
  assign n2725 = n2723 & n2724;
  assign n2726 = pi134  & ~n2725;
  assign po23  = n2718 | n2726;
  assign n2728 = n319 & ~n2022;
  assign n2729 = n425 & ~n2074;
  assign n2730 = n478 & ~n2030;
  assign n2731 = n372 & ~n2038;
  assign n2732 = ~n2728 & ~n2729;
  assign n2733 = ~n2730 & ~n2731;
  assign n2734 = n2732 & n2733;
  assign n2735 = ~pi134  & ~n2734;
  assign n2736 = n372 & ~n2050;
  assign n2737 = n478 & ~n2058;
  assign n2738 = n319 & ~n2066;
  assign n2739 = n425 & ~n2014;
  assign n2740 = ~n2736 & ~n2737;
  assign n2741 = ~n2738 & ~n2739;
  assign n2742 = n2740 & n2741;
  assign n2743 = pi134  & ~n2742;
  assign po24  = n2735 | n2743;
  assign n2745 = n319 & ~n2095;
  assign n2746 = n425 & ~n2147;
  assign n2747 = n478 & ~n2103;
  assign n2748 = n372 & ~n2111;
  assign n2749 = ~n2745 & ~n2746;
  assign n2750 = ~n2747 & ~n2748;
  assign n2751 = n2749 & n2750;
  assign n2752 = ~pi134  & ~n2751;
  assign n2753 = n372 & ~n2123;
  assign n2754 = n478 & ~n2131;
  assign n2755 = n319 & ~n2139;
  assign n2756 = n425 & ~n2087;
  assign n2757 = ~n2753 & ~n2754;
  assign n2758 = ~n2755 & ~n2756;
  assign n2759 = n2757 & n2758;
  assign n2760 = pi134  & ~n2759;
  assign po25  = n2752 | n2760;
  assign n2762 = n319 & ~n2168;
  assign n2763 = n372 & ~n2184;
  assign n2764 = n425 & ~n2220;
  assign n2765 = n478 & ~n2176;
  assign n2766 = ~n2762 & ~n2763;
  assign n2767 = ~n2764 & ~n2765;
  assign n2768 = n2766 & n2767;
  assign n2769 = ~pi134  & ~n2768;
  assign n2770 = n372 & ~n2196;
  assign n2771 = n478 & ~n2204;
  assign n2772 = n319 & ~n2212;
  assign n2773 = n425 & ~n2160;
  assign n2774 = ~n2770 & ~n2771;
  assign n2775 = ~n2772 & ~n2773;
  assign n2776 = n2774 & n2775;
  assign n2777 = pi134  & ~n2776;
  assign po26  = n2769 | n2777;
  assign n2779 = n319 & ~n2241;
  assign n2780 = n372 & ~n2257;
  assign n2781 = n425 & ~n2293;
  assign n2782 = n478 & ~n2249;
  assign n2783 = ~n2779 & ~n2780;
  assign n2784 = ~n2781 & ~n2782;
  assign n2785 = n2783 & n2784;
  assign n2786 = ~pi134  & ~n2785;
  assign n2787 = n372 & ~n2269;
  assign n2788 = n478 & ~n2277;
  assign n2789 = n319 & ~n2285;
  assign n2790 = n425 & ~n2233;
  assign n2791 = ~n2787 & ~n2788;
  assign n2792 = ~n2789 & ~n2790;
  assign n2793 = n2791 & n2792;
  assign n2794 = pi134  & ~n2793;
  assign po27  = n2786 | n2794;
  assign n2796 = n319 & ~n2314;
  assign n2797 = n372 & ~n2330;
  assign n2798 = n425 & ~n2366;
  assign n2799 = n478 & ~n2322;
  assign n2800 = ~n2796 & ~n2797;
  assign n2801 = ~n2798 & ~n2799;
  assign n2802 = n2800 & n2801;
  assign n2803 = ~pi134  & ~n2802;
  assign n2804 = n372 & ~n2342;
  assign n2805 = n478 & ~n2350;
  assign n2806 = n319 & ~n2358;
  assign n2807 = n425 & ~n2306;
  assign n2808 = ~n2804 & ~n2805;
  assign n2809 = ~n2806 & ~n2807;
  assign n2810 = n2808 & n2809;
  assign n2811 = pi134  & ~n2810;
  assign po28  = n2803 | n2811;
  assign n2813 = n319 & ~n2387;
  assign n2814 = n372 & ~n2403;
  assign n2815 = n425 & ~n2439;
  assign n2816 = n478 & ~n2395;
  assign n2817 = ~n2813 & ~n2814;
  assign n2818 = ~n2815 & ~n2816;
  assign n2819 = n2817 & n2818;
  assign n2820 = ~pi134  & ~n2819;
  assign n2821 = n372 & ~n2415;
  assign n2822 = n478 & ~n2423;
  assign n2823 = n319 & ~n2431;
  assign n2824 = n425 & ~n2379;
  assign n2825 = ~n2821 & ~n2822;
  assign n2826 = ~n2823 & ~n2824;
  assign n2827 = n2825 & n2826;
  assign n2828 = pi134  & ~n2827;
  assign po29  = n2820 | n2828;
  assign n2830 = n319 & ~n2460;
  assign n2831 = n372 & ~n2476;
  assign n2832 = n425 & ~n2512;
  assign n2833 = n478 & ~n2468;
  assign n2834 = ~n2830 & ~n2831;
  assign n2835 = ~n2832 & ~n2833;
  assign n2836 = n2834 & n2835;
  assign n2837 = ~pi134  & ~n2836;
  assign n2838 = n372 & ~n2488;
  assign n2839 = n478 & ~n2496;
  assign n2840 = n319 & ~n2504;
  assign n2841 = n425 & ~n2452;
  assign n2842 = ~n2838 & ~n2839;
  assign n2843 = ~n2840 & ~n2841;
  assign n2844 = n2842 & n2843;
  assign n2845 = pi134  & ~n2844;
  assign po30  = n2837 | n2845;
  assign n2847 = n319 & ~n2533;
  assign n2848 = n372 & ~n2549;
  assign n2849 = n425 & ~n2585;
  assign n2850 = n478 & ~n2541;
  assign n2851 = ~n2847 & ~n2848;
  assign n2852 = ~n2849 & ~n2850;
  assign n2853 = n2851 & n2852;
  assign n2854 = ~pi134  & ~n2853;
  assign n2855 = n372 & ~n2561;
  assign n2856 = n478 & ~n2569;
  assign n2857 = n319 & ~n2577;
  assign n2858 = n425 & ~n2525;
  assign n2859 = ~n2855 & ~n2856;
  assign n2860 = ~n2857 & ~n2858;
  assign n2861 = n2859 & n2860;
  assign n2862 = pi134  & ~n2861;
  assign po31  = n2854 | n2862;
  assign n2864 = n319 & ~n477;
  assign n2865 = n372 & ~n424;
  assign n2866 = n425 & ~n586;
  assign n2867 = n478 & ~n534;
  assign n2868 = ~n2864 & ~n2865;
  assign n2869 = ~n2866 & ~n2867;
  assign n2870 = n2868 & n2869;
  assign n2871 = ~pi134  & ~n2870;
  assign n2872 = ~n318 & n478;
  assign n2873 = ~n371 & n425;
  assign n2874 = n372 & ~n638;
  assign n2875 = n319 & ~n690;
  assign n2876 = ~n2872 & ~n2873;
  assign n2877 = ~n2874 & ~n2875;
  assign n2878 = n2876 & n2877;
  assign n2879 = pi134  & ~n2878;
  assign po32  = n2871 | n2879;
  assign n2881 = n319 & ~n903;
  assign n2882 = n372 & ~n851;
  assign n2883 = n425 & ~n1115;
  assign n2884 = n478 & ~n1011;
  assign n2885 = ~n2881 & ~n2882;
  assign n2886 = ~n2883 & ~n2884;
  assign n2887 = n2885 & n2886;
  assign n2888 = ~pi134  & ~n2887;
  assign n2889 = n372 & ~n959;
  assign n2890 = n478 & ~n747;
  assign n2891 = n319 & ~n1063;
  assign n2892 = n425 & ~n799;
  assign n2893 = ~n2889 & ~n2890;
  assign n2894 = ~n2891 & ~n2892;
  assign n2895 = n2893 & n2894;
  assign n2896 = pi134  & ~n2895;
  assign po33  = n2888 | n2896;
  assign n2898 = n319 & ~n1264;
  assign n2899 = n372 & ~n1228;
  assign n2900 = n425 & ~n1412;
  assign n2901 = n478 & ~n1340;
  assign n2902 = ~n2898 & ~n2899;
  assign n2903 = ~n2900 & ~n2901;
  assign n2904 = n2902 & n2903;
  assign n2905 = ~pi134  & ~n2904;
  assign n2906 = n372 & ~n1304;
  assign n2907 = n478 & ~n1156;
  assign n2908 = n319 & ~n1376;
  assign n2909 = n425 & ~n1192;
  assign n2910 = ~n2906 & ~n2907;
  assign n2911 = ~n2908 & ~n2909;
  assign n2912 = n2910 & n2911;
  assign n2913 = pi134  & ~n2912;
  assign po34  = n2905 | n2913;
  assign n2915 = n319 & ~n1453;
  assign n2916 = n425 & ~n1709;
  assign n2917 = n372 & ~n1525;
  assign n2918 = n478 & ~n1673;
  assign n2919 = ~n2915 & ~n2916;
  assign n2920 = ~n2917 & ~n2918;
  assign n2921 = n2919 & n2920;
  assign n2922 = ~pi134  & ~n2921;
  assign n2923 = n372 & ~n1601;
  assign n2924 = n425 & ~n1489;
  assign n2925 = n319 & ~n1637;
  assign n2926 = n478 & ~n1561;
  assign n2927 = ~n2923 & ~n2924;
  assign n2928 = ~n2925 & ~n2926;
  assign n2929 = n2927 & n2928;
  assign n2930 = pi134  & ~n2929;
  assign po35  = n2922 | n2930;
  assign n2932 = n319 & ~n1746;
  assign n2933 = n372 & ~n1738;
  assign n2934 = n425 & ~n1774;
  assign n2935 = n478 & ~n1782;
  assign n2936 = ~n2932 & ~n2933;
  assign n2937 = ~n2934 & ~n2935;
  assign n2938 = n2936 & n2937;
  assign n2939 = ~pi134  & ~n2938;
  assign n2940 = n478 & ~n1722;
  assign n2941 = n425 & ~n1730;
  assign n2942 = n372 & ~n1766;
  assign n2943 = n319 & ~n1758;
  assign n2944 = ~n2940 & ~n2941;
  assign n2945 = ~n2942 & ~n2943;
  assign n2946 = n2944 & n2945;
  assign n2947 = pi134  & ~n2946;
  assign po36  = n2939 | n2947;
  assign n2949 = n319 & ~n1819;
  assign n2950 = n372 & ~n1811;
  assign n2951 = n425 & ~n1847;
  assign n2952 = n478 & ~n1855;
  assign n2953 = ~n2949 & ~n2950;
  assign n2954 = ~n2951 & ~n2952;
  assign n2955 = n2953 & n2954;
  assign n2956 = ~pi134  & ~n2955;
  assign n2957 = n478 & ~n1795;
  assign n2958 = n425 & ~n1803;
  assign n2959 = n372 & ~n1839;
  assign n2960 = n319 & ~n1831;
  assign n2961 = ~n2957 & ~n2958;
  assign n2962 = ~n2959 & ~n2960;
  assign n2963 = n2961 & n2962;
  assign n2964 = pi134  & ~n2963;
  assign po37  = n2956 | n2964;
  assign n2966 = n319 & ~n1892;
  assign n2967 = n372 & ~n1884;
  assign n2968 = n425 & ~n1920;
  assign n2969 = n478 & ~n1928;
  assign n2970 = ~n2966 & ~n2967;
  assign n2971 = ~n2968 & ~n2969;
  assign n2972 = n2970 & n2971;
  assign n2973 = ~pi134  & ~n2972;
  assign n2974 = n478 & ~n1868;
  assign n2975 = n425 & ~n1876;
  assign n2976 = n372 & ~n1912;
  assign n2977 = n319 & ~n1904;
  assign n2978 = ~n2974 & ~n2975;
  assign n2979 = ~n2976 & ~n2977;
  assign n2980 = n2978 & n2979;
  assign n2981 = pi134  & ~n2980;
  assign po38  = n2973 | n2981;
  assign n2983 = n478 & ~n2001;
  assign n2984 = n425 & ~n1993;
  assign n2985 = n372 & ~n1957;
  assign n2986 = n319 & ~n1965;
  assign n2987 = ~n2983 & ~n2984;
  assign n2988 = ~n2985 & ~n2986;
  assign n2989 = n2987 & n2988;
  assign n2990 = ~pi134  & ~n2989;
  assign n2991 = n319 & ~n1977;
  assign n2992 = n372 & ~n1985;
  assign n2993 = n425 & ~n1949;
  assign n2994 = n478 & ~n1941;
  assign n2995 = ~n2991 & ~n2992;
  assign n2996 = ~n2993 & ~n2994;
  assign n2997 = n2995 & n2996;
  assign n2998 = pi134  & ~n2997;
  assign po39  = n2990 | n2998;
  assign n3000 = n478 & ~n2074;
  assign n3001 = n425 & ~n2066;
  assign n3002 = n372 & ~n2030;
  assign n3003 = n319 & ~n2038;
  assign n3004 = ~n3000 & ~n3001;
  assign n3005 = ~n3002 & ~n3003;
  assign n3006 = n3004 & n3005;
  assign n3007 = ~pi134  & ~n3006;
  assign n3008 = n319 & ~n2050;
  assign n3009 = n372 & ~n2058;
  assign n3010 = n425 & ~n2022;
  assign n3011 = n478 & ~n2014;
  assign n3012 = ~n3008 & ~n3009;
  assign n3013 = ~n3010 & ~n3011;
  assign n3014 = n3012 & n3013;
  assign n3015 = pi134  & ~n3014;
  assign po40  = n3007 | n3015;
  assign n3017 = n478 & ~n2147;
  assign n3018 = n425 & ~n2139;
  assign n3019 = n372 & ~n2103;
  assign n3020 = n319 & ~n2111;
  assign n3021 = ~n3017 & ~n3018;
  assign n3022 = ~n3019 & ~n3020;
  assign n3023 = n3021 & n3022;
  assign n3024 = ~pi134  & ~n3023;
  assign n3025 = n319 & ~n2123;
  assign n3026 = n372 & ~n2131;
  assign n3027 = n425 & ~n2095;
  assign n3028 = n478 & ~n2087;
  assign n3029 = ~n3025 & ~n3026;
  assign n3030 = ~n3027 & ~n3028;
  assign n3031 = n3029 & n3030;
  assign n3032 = pi134  & ~n3031;
  assign po41  = n3024 | n3032;
  assign n3034 = n319 & ~n2184;
  assign n3035 = n372 & ~n2176;
  assign n3036 = n425 & ~n2212;
  assign n3037 = n478 & ~n2220;
  assign n3038 = ~n3034 & ~n3035;
  assign n3039 = ~n3036 & ~n3037;
  assign n3040 = n3038 & n3039;
  assign n3041 = ~pi134  & ~n3040;
  assign n3042 = n319 & ~n2196;
  assign n3043 = n372 & ~n2204;
  assign n3044 = n425 & ~n2168;
  assign n3045 = n478 & ~n2160;
  assign n3046 = ~n3042 & ~n3043;
  assign n3047 = ~n3044 & ~n3045;
  assign n3048 = n3046 & n3047;
  assign n3049 = pi134  & ~n3048;
  assign po42  = n3041 | n3049;
  assign n3051 = n319 & ~n2257;
  assign n3052 = n372 & ~n2249;
  assign n3053 = n425 & ~n2285;
  assign n3054 = n478 & ~n2293;
  assign n3055 = ~n3051 & ~n3052;
  assign n3056 = ~n3053 & ~n3054;
  assign n3057 = n3055 & n3056;
  assign n3058 = ~pi134  & ~n3057;
  assign n3059 = n319 & ~n2269;
  assign n3060 = n372 & ~n2277;
  assign n3061 = n425 & ~n2241;
  assign n3062 = n478 & ~n2233;
  assign n3063 = ~n3059 & ~n3060;
  assign n3064 = ~n3061 & ~n3062;
  assign n3065 = n3063 & n3064;
  assign n3066 = pi134  & ~n3065;
  assign po43  = n3058 | n3066;
  assign n3068 = n319 & ~n2330;
  assign n3069 = n372 & ~n2322;
  assign n3070 = n425 & ~n2358;
  assign n3071 = n478 & ~n2366;
  assign n3072 = ~n3068 & ~n3069;
  assign n3073 = ~n3070 & ~n3071;
  assign n3074 = n3072 & n3073;
  assign n3075 = ~pi134  & ~n3074;
  assign n3076 = n319 & ~n2342;
  assign n3077 = n372 & ~n2350;
  assign n3078 = n425 & ~n2314;
  assign n3079 = n478 & ~n2306;
  assign n3080 = ~n3076 & ~n3077;
  assign n3081 = ~n3078 & ~n3079;
  assign n3082 = n3080 & n3081;
  assign n3083 = pi134  & ~n3082;
  assign po44  = n3075 | n3083;
  assign n3085 = n319 & ~n2403;
  assign n3086 = n372 & ~n2395;
  assign n3087 = n425 & ~n2431;
  assign n3088 = n478 & ~n2439;
  assign n3089 = ~n3085 & ~n3086;
  assign n3090 = ~n3087 & ~n3088;
  assign n3091 = n3089 & n3090;
  assign n3092 = ~pi134  & ~n3091;
  assign n3093 = n319 & ~n2415;
  assign n3094 = n372 & ~n2423;
  assign n3095 = n425 & ~n2387;
  assign n3096 = n478 & ~n2379;
  assign n3097 = ~n3093 & ~n3094;
  assign n3098 = ~n3095 & ~n3096;
  assign n3099 = n3097 & n3098;
  assign n3100 = pi134  & ~n3099;
  assign po45  = n3092 | n3100;
  assign n3102 = n319 & ~n2476;
  assign n3103 = n372 & ~n2468;
  assign n3104 = n425 & ~n2504;
  assign n3105 = n478 & ~n2512;
  assign n3106 = ~n3102 & ~n3103;
  assign n3107 = ~n3104 & ~n3105;
  assign n3108 = n3106 & n3107;
  assign n3109 = ~pi134  & ~n3108;
  assign n3110 = n319 & ~n2488;
  assign n3111 = n372 & ~n2496;
  assign n3112 = n425 & ~n2460;
  assign n3113 = n478 & ~n2452;
  assign n3114 = ~n3110 & ~n3111;
  assign n3115 = ~n3112 & ~n3113;
  assign n3116 = n3114 & n3115;
  assign n3117 = pi134  & ~n3116;
  assign po46  = n3109 | n3117;
  assign n3119 = n319 & ~n2549;
  assign n3120 = n372 & ~n2541;
  assign n3121 = n425 & ~n2577;
  assign n3122 = n478 & ~n2585;
  assign n3123 = ~n3119 & ~n3120;
  assign n3124 = ~n3121 & ~n3122;
  assign n3125 = n3123 & n3124;
  assign n3126 = ~pi134  & ~n3125;
  assign n3127 = n319 & ~n2561;
  assign n3128 = n372 & ~n2569;
  assign n3129 = n425 & ~n2533;
  assign n3130 = n478 & ~n2525;
  assign n3131 = ~n3127 & ~n3128;
  assign n3132 = ~n3129 & ~n3130;
  assign n3133 = n3131 & n3132;
  assign n3134 = pi134  & ~n3133;
  assign po47  = n3126 | n3134;
  assign n3136 = n319 & ~n424;
  assign n3137 = n372 & ~n534;
  assign n3138 = n425 & ~n690;
  assign n3139 = n478 & ~n586;
  assign n3140 = ~n3136 & ~n3137;
  assign n3141 = ~n3138 & ~n3139;
  assign n3142 = n3140 & n3141;
  assign n3143 = ~pi134  & ~n3142;
  assign n3144 = ~n318 & n372;
  assign n3145 = ~n371 & n478;
  assign n3146 = n319 & ~n638;
  assign n3147 = n425 & ~n477;
  assign n3148 = ~n3144 & ~n3145;
  assign n3149 = ~n3146 & ~n3147;
  assign n3150 = n3148 & n3149;
  assign n3151 = pi134  & ~n3150;
  assign po48  = n3143 | n3151;
  assign n3153 = n319 & ~n851;
  assign n3154 = n372 & ~n1011;
  assign n3155 = n425 & ~n1063;
  assign n3156 = n478 & ~n1115;
  assign n3157 = ~n3153 & ~n3154;
  assign n3158 = ~n3155 & ~n3156;
  assign n3159 = n3157 & n3158;
  assign n3160 = ~pi134  & ~n3159;
  assign n3161 = n319 & ~n959;
  assign n3162 = n372 & ~n747;
  assign n3163 = n425 & ~n903;
  assign n3164 = n478 & ~n799;
  assign n3165 = ~n3161 & ~n3162;
  assign n3166 = ~n3163 & ~n3164;
  assign n3167 = n3165 & n3166;
  assign n3168 = pi134  & ~n3167;
  assign po49  = n3160 | n3168;
  assign n3170 = n319 & ~n1228;
  assign n3171 = n372 & ~n1340;
  assign n3172 = n425 & ~n1376;
  assign n3173 = n478 & ~n1412;
  assign n3174 = ~n3170 & ~n3171;
  assign n3175 = ~n3172 & ~n3173;
  assign n3176 = n3174 & n3175;
  assign n3177 = ~pi134  & ~n3176;
  assign n3178 = n319 & ~n1304;
  assign n3179 = n372 & ~n1156;
  assign n3180 = n425 & ~n1264;
  assign n3181 = n478 & ~n1192;
  assign n3182 = ~n3178 & ~n3179;
  assign n3183 = ~n3180 & ~n3181;
  assign n3184 = n3182 & n3183;
  assign n3185 = pi134  & ~n3184;
  assign po50  = n3177 | n3185;
  assign n3187 = n425 & ~n1637;
  assign n3188 = n478 & ~n1709;
  assign n3189 = n319 & ~n1525;
  assign n3190 = n372 & ~n1673;
  assign n3191 = ~n3187 & ~n3188;
  assign n3192 = ~n3189 & ~n3190;
  assign n3193 = n3191 & n3192;
  assign n3194 = ~pi134  & ~n3193;
  assign n3195 = n319 & ~n1601;
  assign n3196 = n425 & ~n1453;
  assign n3197 = n372 & ~n1561;
  assign n3198 = n478 & ~n1489;
  assign n3199 = ~n3195 & ~n3196;
  assign n3200 = ~n3197 & ~n3198;
  assign n3201 = n3199 & n3200;
  assign n3202 = pi134  & ~n3201;
  assign po51  = n3194 | n3202;
  assign n3204 = n425 & ~n1758;
  assign n3205 = n319 & ~n1738;
  assign n3206 = n478 & ~n1774;
  assign n3207 = n372 & ~n1782;
  assign n3208 = ~n3204 & ~n3205;
  assign n3209 = ~n3206 & ~n3207;
  assign n3210 = n3208 & n3209;
  assign n3211 = ~pi134  & ~n3210;
  assign n3212 = n372 & ~n1722;
  assign n3213 = n478 & ~n1730;
  assign n3214 = n425 & ~n1746;
  assign n3215 = n319 & ~n1766;
  assign n3216 = ~n3212 & ~n3213;
  assign n3217 = ~n3214 & ~n3215;
  assign n3218 = n3216 & n3217;
  assign n3219 = pi134  & ~n3218;
  assign po52  = n3211 | n3219;
  assign n3221 = n425 & ~n1831;
  assign n3222 = n319 & ~n1811;
  assign n3223 = n478 & ~n1847;
  assign n3224 = n372 & ~n1855;
  assign n3225 = ~n3221 & ~n3222;
  assign n3226 = ~n3223 & ~n3224;
  assign n3227 = n3225 & n3226;
  assign n3228 = ~pi134  & ~n3227;
  assign n3229 = n372 & ~n1795;
  assign n3230 = n478 & ~n1803;
  assign n3231 = n425 & ~n1819;
  assign n3232 = n319 & ~n1839;
  assign n3233 = ~n3229 & ~n3230;
  assign n3234 = ~n3231 & ~n3232;
  assign n3235 = n3233 & n3234;
  assign n3236 = pi134  & ~n3235;
  assign po53  = n3228 | n3236;
  assign n3238 = n425 & ~n1904;
  assign n3239 = n319 & ~n1884;
  assign n3240 = n478 & ~n1920;
  assign n3241 = n372 & ~n1928;
  assign n3242 = ~n3238 & ~n3239;
  assign n3243 = ~n3240 & ~n3241;
  assign n3244 = n3242 & n3243;
  assign n3245 = ~pi134  & ~n3244;
  assign n3246 = n372 & ~n1868;
  assign n3247 = n478 & ~n1876;
  assign n3248 = n425 & ~n1892;
  assign n3249 = n319 & ~n1912;
  assign n3250 = ~n3246 & ~n3247;
  assign n3251 = ~n3248 & ~n3249;
  assign n3252 = n3250 & n3251;
  assign n3253 = pi134  & ~n3252;
  assign po54  = n3245 | n3253;
  assign n3255 = n425 & ~n1977;
  assign n3256 = n372 & ~n2001;
  assign n3257 = n319 & ~n1957;
  assign n3258 = n478 & ~n1993;
  assign n3259 = ~n3255 & ~n3256;
  assign n3260 = ~n3257 & ~n3258;
  assign n3261 = n3259 & n3260;
  assign n3262 = ~pi134  & ~n3261;
  assign n3263 = n319 & ~n1985;
  assign n3264 = n372 & ~n1941;
  assign n3265 = n425 & ~n1965;
  assign n3266 = n478 & ~n1949;
  assign n3267 = ~n3263 & ~n3264;
  assign n3268 = ~n3265 & ~n3266;
  assign n3269 = n3267 & n3268;
  assign n3270 = pi134  & ~n3269;
  assign po55  = n3262 | n3270;
  assign n3272 = n425 & ~n2050;
  assign n3273 = n372 & ~n2074;
  assign n3274 = n319 & ~n2030;
  assign n3275 = n478 & ~n2066;
  assign n3276 = ~n3272 & ~n3273;
  assign n3277 = ~n3274 & ~n3275;
  assign n3278 = n3276 & n3277;
  assign n3279 = ~pi134  & ~n3278;
  assign n3280 = n319 & ~n2058;
  assign n3281 = n372 & ~n2014;
  assign n3282 = n425 & ~n2038;
  assign n3283 = n478 & ~n2022;
  assign n3284 = ~n3280 & ~n3281;
  assign n3285 = ~n3282 & ~n3283;
  assign n3286 = n3284 & n3285;
  assign n3287 = pi134  & ~n3286;
  assign po56  = n3279 | n3287;
  assign n3289 = n425 & ~n2123;
  assign n3290 = n372 & ~n2147;
  assign n3291 = n319 & ~n2103;
  assign n3292 = n478 & ~n2139;
  assign n3293 = ~n3289 & ~n3290;
  assign n3294 = ~n3291 & ~n3292;
  assign n3295 = n3293 & n3294;
  assign n3296 = ~pi134  & ~n3295;
  assign n3297 = n319 & ~n2131;
  assign n3298 = n372 & ~n2087;
  assign n3299 = n425 & ~n2111;
  assign n3300 = n478 & ~n2095;
  assign n3301 = ~n3297 & ~n3298;
  assign n3302 = ~n3299 & ~n3300;
  assign n3303 = n3301 & n3302;
  assign n3304 = pi134  & ~n3303;
  assign po57  = n3296 | n3304;
  assign n3306 = n425 & ~n2196;
  assign n3307 = n319 & ~n2176;
  assign n3308 = n478 & ~n2212;
  assign n3309 = n372 & ~n2220;
  assign n3310 = ~n3306 & ~n3307;
  assign n3311 = ~n3308 & ~n3309;
  assign n3312 = n3310 & n3311;
  assign n3313 = ~pi134  & ~n3312;
  assign n3314 = n319 & ~n2204;
  assign n3315 = n372 & ~n2160;
  assign n3316 = n425 & ~n2184;
  assign n3317 = n478 & ~n2168;
  assign n3318 = ~n3314 & ~n3315;
  assign n3319 = ~n3316 & ~n3317;
  assign n3320 = n3318 & n3319;
  assign n3321 = pi134  & ~n3320;
  assign po58  = n3313 | n3321;
  assign n3323 = n425 & ~n2269;
  assign n3324 = n319 & ~n2249;
  assign n3325 = n478 & ~n2285;
  assign n3326 = n372 & ~n2293;
  assign n3327 = ~n3323 & ~n3324;
  assign n3328 = ~n3325 & ~n3326;
  assign n3329 = n3327 & n3328;
  assign n3330 = ~pi134  & ~n3329;
  assign n3331 = n319 & ~n2277;
  assign n3332 = n372 & ~n2233;
  assign n3333 = n425 & ~n2257;
  assign n3334 = n478 & ~n2241;
  assign n3335 = ~n3331 & ~n3332;
  assign n3336 = ~n3333 & ~n3334;
  assign n3337 = n3335 & n3336;
  assign n3338 = pi134  & ~n3337;
  assign po59  = n3330 | n3338;
  assign n3340 = n425 & ~n2342;
  assign n3341 = n319 & ~n2322;
  assign n3342 = n478 & ~n2358;
  assign n3343 = n372 & ~n2366;
  assign n3344 = ~n3340 & ~n3341;
  assign n3345 = ~n3342 & ~n3343;
  assign n3346 = n3344 & n3345;
  assign n3347 = ~pi134  & ~n3346;
  assign n3348 = n319 & ~n2350;
  assign n3349 = n372 & ~n2306;
  assign n3350 = n425 & ~n2330;
  assign n3351 = n478 & ~n2314;
  assign n3352 = ~n3348 & ~n3349;
  assign n3353 = ~n3350 & ~n3351;
  assign n3354 = n3352 & n3353;
  assign n3355 = pi134  & ~n3354;
  assign po60  = n3347 | n3355;
  assign n3357 = n425 & ~n2415;
  assign n3358 = n319 & ~n2395;
  assign n3359 = n478 & ~n2431;
  assign n3360 = n372 & ~n2439;
  assign n3361 = ~n3357 & ~n3358;
  assign n3362 = ~n3359 & ~n3360;
  assign n3363 = n3361 & n3362;
  assign n3364 = ~pi134  & ~n3363;
  assign n3365 = n319 & ~n2423;
  assign n3366 = n372 & ~n2379;
  assign n3367 = n425 & ~n2403;
  assign n3368 = n478 & ~n2387;
  assign n3369 = ~n3365 & ~n3366;
  assign n3370 = ~n3367 & ~n3368;
  assign n3371 = n3369 & n3370;
  assign n3372 = pi134  & ~n3371;
  assign po61  = n3364 | n3372;
  assign n3374 = n425 & ~n2488;
  assign n3375 = n319 & ~n2468;
  assign n3376 = n478 & ~n2504;
  assign n3377 = n372 & ~n2512;
  assign n3378 = ~n3374 & ~n3375;
  assign n3379 = ~n3376 & ~n3377;
  assign n3380 = n3378 & n3379;
  assign n3381 = ~pi134  & ~n3380;
  assign n3382 = n319 & ~n2496;
  assign n3383 = n372 & ~n2452;
  assign n3384 = n425 & ~n2476;
  assign n3385 = n478 & ~n2460;
  assign n3386 = ~n3382 & ~n3383;
  assign n3387 = ~n3384 & ~n3385;
  assign n3388 = n3386 & n3387;
  assign n3389 = pi134  & ~n3388;
  assign po62  = n3381 | n3389;
  assign n3391 = n425 & ~n2561;
  assign n3392 = n319 & ~n2541;
  assign n3393 = n478 & ~n2577;
  assign n3394 = n372 & ~n2585;
  assign n3395 = ~n3391 & ~n3392;
  assign n3396 = ~n3393 & ~n3394;
  assign n3397 = n3395 & n3396;
  assign n3398 = ~pi134  & ~n3397;
  assign n3399 = n319 & ~n2569;
  assign n3400 = n372 & ~n2525;
  assign n3401 = n425 & ~n2549;
  assign n3402 = n478 & ~n2533;
  assign n3403 = ~n3399 & ~n3400;
  assign n3404 = ~n3401 & ~n3402;
  assign n3405 = n3403 & n3404;
  assign n3406 = pi134  & ~n3405;
  assign po63  = n3398 | n3406;
  assign n3408 = ~pi134  & ~n694;
  assign n3409 = pi134  & ~n482;
  assign po64  = n3408 | n3409;
  assign n3411 = ~pi134  & ~n1119;
  assign n3412 = pi134  & ~n907;
  assign po65  = n3411 | n3412;
  assign n3414 = ~pi134  & ~n1416;
  assign n3415 = pi134  & ~n1268;
  assign po66  = n3414 | n3415;
  assign n3417 = ~pi134  & ~n1713;
  assign n3418 = pi134  & ~n1565;
  assign po67  = n3417 | n3418;
  assign n3420 = ~pi134  & ~n1786;
  assign n3421 = pi134  & ~n1750;
  assign po68  = n3420 | n3421;
  assign n3423 = ~pi134  & ~n1859;
  assign n3424 = pi134  & ~n1823;
  assign po69  = n3423 | n3424;
  assign n3426 = ~pi134  & ~n1932;
  assign n3427 = pi134  & ~n1896;
  assign po70  = n3426 | n3427;
  assign n3429 = ~pi134  & ~n2005;
  assign n3430 = pi134  & ~n1969;
  assign po71  = n3429 | n3430;
  assign n3432 = ~pi134  & ~n2078;
  assign n3433 = pi134  & ~n2042;
  assign po72  = n3432 | n3433;
  assign n3435 = ~pi134  & ~n2151;
  assign n3436 = pi134  & ~n2115;
  assign po73  = n3435 | n3436;
  assign n3438 = ~pi134  & ~n2224;
  assign n3439 = pi134  & ~n2188;
  assign po74  = n3438 | n3439;
  assign n3441 = ~pi134  & ~n2297;
  assign n3442 = pi134  & ~n2261;
  assign po75  = n3441 | n3442;
  assign n3444 = ~pi134  & ~n2370;
  assign n3445 = pi134  & ~n2334;
  assign po76  = n3444 | n3445;
  assign n3447 = ~pi134  & ~n2443;
  assign n3448 = pi134  & ~n2407;
  assign po77  = n3447 | n3448;
  assign n3450 = ~pi134  & ~n2516;
  assign n3451 = pi134  & ~n2480;
  assign po78  = n3450 | n3451;
  assign n3453 = ~pi134  & ~n2589;
  assign n3454 = pi134  & ~n2553;
  assign po79  = n3453 | n3454;
  assign n3456 = ~pi134  & ~n2606;
  assign n3457 = pi134  & ~n2598;
  assign po80  = n3456 | n3457;
  assign n3459 = ~pi134  & ~n2623;
  assign n3460 = pi134  & ~n2615;
  assign po81  = n3459 | n3460;
  assign n3462 = ~pi134  & ~n2640;
  assign n3463 = pi134  & ~n2632;
  assign po82  = n3462 | n3463;
  assign n3465 = ~pi134  & ~n2657;
  assign n3466 = pi134  & ~n2649;
  assign po83  = n3465 | n3466;
  assign n3468 = ~pi134  & ~n2674;
  assign n3469 = pi134  & ~n2666;
  assign po84  = n3468 | n3469;
  assign n3471 = ~pi134  & ~n2691;
  assign n3472 = pi134  & ~n2683;
  assign po85  = n3471 | n3472;
  assign n3474 = ~pi134  & ~n2708;
  assign n3475 = pi134  & ~n2700;
  assign po86  = n3474 | n3475;
  assign n3477 = ~pi134  & ~n2725;
  assign n3478 = pi134  & ~n2717;
  assign po87  = n3477 | n3478;
  assign n3480 = ~pi134  & ~n2742;
  assign n3481 = pi134  & ~n2734;
  assign po88  = n3480 | n3481;
  assign n3483 = ~pi134  & ~n2759;
  assign n3484 = pi134  & ~n2751;
  assign po89  = n3483 | n3484;
  assign n3486 = ~pi134  & ~n2776;
  assign n3487 = pi134  & ~n2768;
  assign po90  = n3486 | n3487;
  assign n3489 = ~pi134  & ~n2793;
  assign n3490 = pi134  & ~n2785;
  assign po91  = n3489 | n3490;
  assign n3492 = ~pi134  & ~n2810;
  assign n3493 = pi134  & ~n2802;
  assign po92  = n3492 | n3493;
  assign n3495 = ~pi134  & ~n2827;
  assign n3496 = pi134  & ~n2819;
  assign po93  = n3495 | n3496;
  assign n3498 = ~pi134  & ~n2844;
  assign n3499 = pi134  & ~n2836;
  assign po94  = n3498 | n3499;
  assign n3501 = ~pi134  & ~n2861;
  assign n3502 = pi134  & ~n2853;
  assign po95  = n3501 | n3502;
  assign n3504 = ~pi134  & ~n2878;
  assign n3505 = pi134  & ~n2870;
  assign po96  = n3504 | n3505;
  assign n3507 = ~pi134  & ~n2895;
  assign n3508 = pi134  & ~n2887;
  assign po97  = n3507 | n3508;
  assign n3510 = ~pi134  & ~n2912;
  assign n3511 = pi134  & ~n2904;
  assign po98  = n3510 | n3511;
  assign n3513 = ~pi134  & ~n2929;
  assign n3514 = pi134  & ~n2921;
  assign po99  = n3513 | n3514;
  assign n3516 = ~pi134  & ~n2946;
  assign n3517 = pi134  & ~n2938;
  assign po100  = n3516 | n3517;
  assign n3519 = ~pi134  & ~n2963;
  assign n3520 = pi134  & ~n2955;
  assign po101  = n3519 | n3520;
  assign n3522 = ~pi134  & ~n2980;
  assign n3523 = pi134  & ~n2972;
  assign po102  = n3522 | n3523;
  assign n3525 = ~pi134  & ~n2997;
  assign n3526 = pi134  & ~n2989;
  assign po103  = n3525 | n3526;
  assign n3528 = ~pi134  & ~n3014;
  assign n3529 = pi134  & ~n3006;
  assign po104  = n3528 | n3529;
  assign n3531 = ~pi134  & ~n3031;
  assign n3532 = pi134  & ~n3023;
  assign po105  = n3531 | n3532;
  assign n3534 = ~pi134  & ~n3048;
  assign n3535 = pi134  & ~n3040;
  assign po106  = n3534 | n3535;
  assign n3537 = ~pi134  & ~n3065;
  assign n3538 = pi134  & ~n3057;
  assign po107  = n3537 | n3538;
  assign n3540 = ~pi134  & ~n3082;
  assign n3541 = pi134  & ~n3074;
  assign po108  = n3540 | n3541;
  assign n3543 = ~pi134  & ~n3099;
  assign n3544 = pi134  & ~n3091;
  assign po109  = n3543 | n3544;
  assign n3546 = ~pi134  & ~n3116;
  assign n3547 = pi134  & ~n3108;
  assign po110  = n3546 | n3547;
  assign n3549 = ~pi134  & ~n3133;
  assign n3550 = pi134  & ~n3125;
  assign po111  = n3549 | n3550;
  assign n3552 = ~pi134  & ~n3150;
  assign n3553 = pi134  & ~n3142;
  assign po112  = n3552 | n3553;
  assign n3555 = ~pi134  & ~n3167;
  assign n3556 = pi134  & ~n3159;
  assign po113  = n3555 | n3556;
  assign n3558 = ~pi134  & ~n3184;
  assign n3559 = pi134  & ~n3176;
  assign po114  = n3558 | n3559;
  assign n3561 = ~pi134  & ~n3201;
  assign n3562 = pi134  & ~n3193;
  assign po115  = n3561 | n3562;
  assign n3564 = ~pi134  & ~n3218;
  assign n3565 = pi134  & ~n3210;
  assign po116  = n3564 | n3565;
  assign n3567 = ~pi134  & ~n3235;
  assign n3568 = pi134  & ~n3227;
  assign po117  = n3567 | n3568;
  assign n3570 = ~pi134  & ~n3252;
  assign n3571 = pi134  & ~n3244;
  assign po118  = n3570 | n3571;
  assign n3573 = ~pi134  & ~n3269;
  assign n3574 = pi134  & ~n3261;
  assign po119  = n3573 | n3574;
  assign n3576 = ~pi134  & ~n3286;
  assign n3577 = pi134  & ~n3278;
  assign po120  = n3576 | n3577;
  assign n3579 = ~pi134  & ~n3303;
  assign n3580 = pi134  & ~n3295;
  assign po121  = n3579 | n3580;
  assign n3582 = ~pi134  & ~n3320;
  assign n3583 = pi134  & ~n3312;
  assign po122  = n3582 | n3583;
  assign n3585 = ~pi134  & ~n3337;
  assign n3586 = pi134  & ~n3329;
  assign po123  = n3585 | n3586;
  assign n3588 = ~pi134  & ~n3354;
  assign n3589 = pi134  & ~n3346;
  assign po124  = n3588 | n3589;
  assign n3591 = ~pi134  & ~n3371;
  assign n3592 = pi134  & ~n3363;
  assign po125  = n3591 | n3592;
  assign n3594 = ~pi134  & ~n3388;
  assign n3595 = pi134  & ~n3380;
  assign po126  = n3594 | n3595;
  assign n3597 = ~pi134  & ~n3405;
  assign n3598 = pi134  & ~n3397;
  assign po127  = n3597 | n3598;
endmodule
