module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 , pi32 ,
    pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 , pi40 ,
    pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 , pi56 ,
    pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 , pi64 ,
    pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 , pi80 ,
    pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 , pi88 ,
    pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 , pi103 ,
    pi104 , pi105 , pi106 , pi107 , pi108 , pi109 , pi110 ,
    pi111 , pi112 , pi113 , pi114 , pi115 , pi116 , pi117 ,
    pi118 , pi119 , pi120 , pi121 , pi122 , pi123 , pi124 ,
    pi125 , pi126 , pi127 ,
    po0 , po1 , po2 , po3 , po4 , po5 ,
    po6 , po7 , po8 , po9 , po10 ,
    po11 , po12 , po13 , po14 , po15 ,
    po16 , po17 , po18 , po19 , po20 ,
    po21 , po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 , po30 ,
    po31 , po32 , po33 , po34 , po35 ,
    po36 , po37 , po38 , po39 , po40 ,
    po41 , po42 , po43 , po44 , po45 ,
    po46 , po47 , po48 , po49 , po50 ,
    po51 , po52 , po53 , po54 , po55 ,
    po56 , po57 , po58 , po59 , po60 ,
    po61 , po62 , po63   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    pi32 , pi33 , pi34 , pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 , pi54 , pi55 ,
    pi56 , pi57 , pi58 , pi59 , pi60 , pi61 , pi62 , pi63 ,
    pi64 , pi65 , pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 , pi78 , pi79 ,
    pi80 , pi81 , pi82 , pi83 , pi84 , pi85 , pi86 , pi87 ,
    pi88 , pi89 , pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 , pi109 ,
    pi110 , pi111 , pi112 , pi113 , pi114 , pi115 , pi116 ,
    pi117 , pi118 , pi119 , pi120 , pi121 , pi122 , pi123 ,
    pi124 , pi125 , pi126 , pi127 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 ;
  wire n194, n195, n196, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n214, n215, n216,
    n217, n218, n219, n220, n221, n222, n223,
    n224, n225, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237,
    n238, n240, n241, n242, n243, n244, n245,
    n246, n247, n248, n249, n250, n251, n252,
    n253, n254, n255, n256, n257, n258, n259,
    n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273,
    n274, n275, n277, n278, n279, n280, n281,
    n282, n283, n284, n285, n286, n287, n288,
    n289, n290, n291, n292, n293, n294, n295,
    n296, n297, n298, n299, n300, n301, n302,
    n303, n304, n305, n306, n307, n308, n309,
    n310, n311, n312, n313, n314, n315, n316,
    n317, n318, n319, n320, n321, n322, n323,
    n325, n326, n327, n328, n329, n330, n331,
    n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395,
    n396, n397, n398, n399, n400, n401, n402,
    n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416,
    n417, n418, n419, n420, n421, n422, n423,
    n424, n425, n426, n427, n428, n429, n430,
    n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n452, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n642, n643,
    n644, n645, n646, n647, n648, n649, n650,
    n651, n652, n653, n654, n655, n656, n657,
    n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671,
    n672, n673, n674, n675, n676, n677, n678,
    n679, n680, n681, n682, n683, n684, n685,
    n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699,
    n700, n701, n702, n703, n704, n705, n706,
    n707, n708, n710, n711, n712, n713, n714,
    n715, n716, n717, n718, n719, n720, n721,
    n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735,
    n736, n737, n738, n739, n740, n741, n742,
    n743, n744, n745, n746, n747, n748, n749,
    n750, n751, n752, n753, n754, n755, n756,
    n757, n758, n759, n760, n761, n762, n763,
    n764, n765, n766, n767, n768, n769, n770,
    n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791,
    n792, n793, n794, n795, n796, n797, n798,
    n799, n800, n801, n802, n803, n804, n805,
    n806, n807, n808, n809, n810, n811, n812,
    n813, n814, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827,
    n828, n829, n830, n831, n832, n833, n834,
    n835, n836, n837, n838, n839, n840, n841,
    n842, n843, n844, n845, n846, n847, n848,
    n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n876,
    n877, n878, n879, n880, n881, n882, n883,
    n884, n885, n886, n887, n888, n889, n890,
    n891, n892, n893, n894, n895, n896, n897,
    n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911,
    n912, n913, n914, n915, n916, n917, n918,
    n919, n920, n921, n922, n923, n924, n925,
    n926, n927, n928, n930, n931, n932, n933,
    n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954,
    n955, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968,
    n969, n970, n971, n972, n973, n974, n975,
    n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989,
    n990, n991, n992, n993, n994, n995, n996,
    n997, n998, n999, n1000, n1001, n1002,
    n1003, n1004, n1005, n1006, n1007, n1008,
    n1009, n1010, n1011, n1012, n1013, n1014,
    n1015, n1016, n1017, n1018, n1019, n1020,
    n1021, n1022, n1023, n1024, n1025, n1026,
    n1027, n1028, n1029, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1038,
    n1039, n1040, n1041, n1042, n1043, n1044,
    n1045, n1046, n1047, n1048, n1049, n1050,
    n1051, n1053, n1054, n1055, n1056, n1057,
    n1058, n1059, n1060, n1061, n1062, n1063,
    n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075,
    n1076, n1077, n1078, n1079, n1080, n1081,
    n1082, n1083, n1084, n1085, n1086, n1087,
    n1088, n1089, n1090, n1091, n1092, n1093,
    n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105,
    n1106, n1107, n1108, n1109, n1110, n1111,
    n1112, n1113, n1114, n1115, n1116, n1117,
    n1118, n1119, n1120, n1121, n1122, n1123,
    n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1139, n1140, n1141,
    n1142, n1143, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153,
    n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165,
    n1166, n1167, n1168, n1169, n1170, n1171,
    n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183,
    n1184, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486,
    n1487, n1488, n1489, n1490, n1491, n1492,
    n1493, n1494, n1495, n1496, n1497, n1498,
    n1499, n1500, n1501, n1502, n1503, n1504,
    n1505, n1506, n1507, n1508, n1509, n1510,
    n1511, n1512, n1513, n1514, n1515, n1516,
    n1517, n1518, n1519, n1520, n1521, n1522,
    n1523, n1524, n1525, n1526, n1527, n1528,
    n1529, n1530, n1531, n1532, n1533, n1534,
    n1535, n1536, n1537, n1538, n1539, n1540,
    n1541, n1542, n1543, n1544, n1545, n1546,
    n1547, n1548, n1549, n1550, n1551, n1552,
    n1553, n1554, n1555, n1556, n1557, n1558,
    n1559, n1560, n1561, n1562, n1563, n1564,
    n1565, n1566, n1567, n1568, n1569, n1570,
    n1571, n1572, n1573, n1574, n1575, n1576,
    n1577, n1578, n1579, n1580, n1581, n1582,
    n1583, n1584, n1585, n1586, n1587, n1588,
    n1589, n1590, n1591, n1592, n1593, n1594,
    n1595, n1596, n1597, n1598, n1599, n1600,
    n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612,
    n1613, n1614, n1615, n1616, n1617, n1618,
    n1619, n1620, n1621, n1622, n1623, n1624,
    n1625, n1626, n1627, n1628, n1629, n1630,
    n1631, n1632, n1633, n1634, n1635, n1636,
    n1637, n1638, n1639, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655,
    n1656, n1657, n1658, n1659, n1660, n1661,
    n1662, n1663, n1664, n1665, n1666, n1667,
    n1668, n1669, n1670, n1671, n1672, n1673,
    n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685,
    n1686, n1687, n1688, n1689, n1690, n1691,
    n1692, n1693, n1694, n1695, n1696, n1697,
    n1698, n1699, n1700, n1701, n1702, n1703,
    n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715,
    n1716, n1717, n1718, n1719, n1720, n1721,
    n1722, n1723, n1724, n1725, n1726, n1727,
    n1728, n1729, n1730, n1731, n1732, n1733,
    n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751,
    n1752, n1753, n1754, n1755, n1756, n1757,
    n1758, n1759, n1760, n1761, n1762, n1763,
    n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775,
    n1776, n1777, n1778, n1779, n1780, n1781,
    n1782, n1783, n1784, n1785, n1786, n1787,
    n1788, n1789, n1790, n1791, n1792, n1793,
    n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805,
    n1806, n1807, n1808, n1809, n1810, n1812,
    n1813, n1814, n1815, n1816, n1817, n1818,
    n1819, n1820, n1821, n1822, n1823, n1824,
    n1825, n1826, n1827, n1828, n1829, n1830,
    n1831, n1832, n1833, n1834, n1835, n1836,
    n1837, n1838, n1839, n1840, n1841, n1842,
    n1843, n1844, n1845, n1846, n1847, n1848,
    n1849, n1850, n1851, n1852, n1853, n1854,
    n1855, n1856, n1857, n1858, n1859, n1860,
    n1861, n1862, n1863, n1864, n1865, n1866,
    n1867, n1868, n1869, n1870, n1871, n1872,
    n1873, n1874, n1875, n1876, n1877, n1878,
    n1879, n1880, n1881, n1882, n1883, n1884,
    n1885, n1886, n1887, n1888, n1889, n1890,
    n1891, n1892, n1893, n1894, n1895, n1896,
    n1897, n1898, n1899, n1900, n1901, n1902,
    n1903, n1904, n1905, n1906, n1907, n1908,
    n1909, n1910, n1911, n1912, n1913, n1914,
    n1915, n1916, n1917, n1918, n1919, n1920,
    n1921, n1922, n1923, n1924, n1925, n1926,
    n1927, n1928, n1929, n1930, n1931, n1932,
    n1933, n1934, n1935, n1936, n1937, n1938,
    n1939, n1940, n1941, n1942, n1943, n1944,
    n1945, n1946, n1947, n1948, n1949, n1950,
    n1951, n1952, n1953, n1954, n1955, n1956,
    n1957, n1958, n1959, n1960, n1961, n1962,
    n1963, n1964, n1965, n1966, n1967, n1968,
    n1969, n1970, n1971, n1972, n1973, n1974,
    n1975, n1976, n1977, n1978, n1979, n1980,
    n1981, n1982, n1983, n1984, n1985, n1986,
    n1987, n1988, n1989, n1990, n1991, n1992,
    n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005,
    n2006, n2007, n2008, n2009, n2010, n2011,
    n2012, n2013, n2014, n2015, n2016, n2017,
    n2018, n2019, n2020, n2021, n2022, n2023,
    n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035,
    n2036, n2037, n2038, n2039, n2040, n2041,
    n2042, n2043, n2044, n2045, n2046, n2047,
    n2048, n2049, n2050, n2051, n2052, n2053,
    n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065,
    n2066, n2067, n2068, n2069, n2070, n2071,
    n2072, n2073, n2074, n2075, n2076, n2077,
    n2078, n2079, n2080, n2081, n2082, n2083,
    n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095,
    n2096, n2097, n2098, n2099, n2100, n2101,
    n2102, n2103, n2104, n2105, n2106, n2107,
    n2108, n2109, n2110, n2111, n2112, n2113,
    n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125,
    n2126, n2127, n2128, n2129, n2130, n2131,
    n2132, n2133, n2134, n2135, n2136, n2137,
    n2138, n2139, n2140, n2141, n2142, n2143,
    n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155,
    n2156, n2157, n2158, n2159, n2160, n2161,
    n2162, n2163, n2164, n2165, n2166, n2167,
    n2168, n2169, n2170, n2171, n2172, n2173,
    n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2592, n2593, n2594, n2595, n2596,
    n2597, n2598, n2599, n2600, n2601, n2602,
    n2603, n2604, n2605, n2606, n2607, n2608,
    n2609, n2610, n2611, n2612, n2613, n2614,
    n2615, n2616, n2617, n2618, n2619, n2620,
    n2621, n2622, n2623, n2624, n2625, n2626,
    n2627, n2628, n2629, n2630, n2631, n2632,
    n2633, n2634, n2635, n2636, n2637, n2638,
    n2639, n2640, n2641, n2642, n2643, n2644,
    n2645, n2646, n2647, n2648, n2649, n2650,
    n2651, n2652, n2653, n2654, n2655, n2656,
    n2657, n2658, n2659, n2660, n2661, n2662,
    n2663, n2664, n2665, n2666, n2667, n2668,
    n2669, n2670, n2671, n2672, n2673, n2674,
    n2675, n2676, n2677, n2678, n2679, n2680,
    n2681, n2682, n2683, n2684, n2685, n2686,
    n2687, n2688, n2689, n2690, n2691, n2692,
    n2693, n2694, n2695, n2696, n2697, n2698,
    n2699, n2700, n2701, n2702, n2703, n2704,
    n2705, n2706, n2707, n2708, n2709, n2710,
    n2711, n2712, n2713, n2714, n2715, n2716,
    n2717, n2718, n2719, n2720, n2721, n2722,
    n2723, n2724, n2725, n2726, n2727, n2728,
    n2729, n2730, n2731, n2732, n2733, n2734,
    n2735, n2736, n2737, n2738, n2739, n2740,
    n2741, n2742, n2743, n2744, n2745, n2746,
    n2747, n2748, n2749, n2750, n2751, n2752,
    n2753, n2754, n2755, n2756, n2757, n2758,
    n2759, n2760, n2761, n2762, n2763, n2764,
    n2765, n2766, n2767, n2768, n2769, n2770,
    n2771, n2772, n2773, n2774, n2775, n2776,
    n2777, n2778, n2779, n2780, n2781, n2782,
    n2783, n2784, n2785, n2786, n2787, n2788,
    n2789, n2790, n2791, n2792, n2793, n2794,
    n2795, n2796, n2797, n2798, n2799, n2800,
    n2801, n2802, n2803, n2804, n2805, n2806,
    n2807, n2808, n2809, n2810, n2812, n2813,
    n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825,
    n2826, n2827, n2828, n2829, n2830, n2831,
    n2832, n2833, n2834, n2835, n2836, n2837,
    n2838, n2839, n2840, n2841, n2842, n2843,
    n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855,
    n2856, n2857, n2858, n2859, n2860, n2861,
    n2862, n2863, n2864, n2865, n2866, n2867,
    n2868, n2869, n2870, n2871, n2872, n2873,
    n2874, n2875, n2876, n2877, n2878, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885,
    n2886, n2887, n2888, n2889, n2890, n2891,
    n2892, n2893, n2894, n2895, n2896, n2897,
    n2898, n2899, n2900, n2901, n2902, n2903,
    n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915,
    n2916, n2917, n2918, n2919, n2920, n2921,
    n2922, n2923, n2924, n2925, n2926, n2927,
    n2928, n2929, n2930, n2931, n2932, n2933,
    n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945,
    n2946, n2947, n2948, n2949, n2950, n2951,
    n2952, n2953, n2954, n2955, n2956, n2957,
    n2958, n2959, n2960, n2961, n2962, n2963,
    n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975,
    n2976, n2977, n2978, n2979, n2980, n2981,
    n2982, n2983, n2984, n2985, n2986, n2987,
    n2988, n2989, n2990, n2991, n2992, n2993,
    n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005,
    n3006, n3007, n3008, n3009, n3010, n3011,
    n3012, n3013, n3014, n3015, n3016, n3017,
    n3018, n3019, n3020, n3021, n3022, n3023,
    n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035,
    n3036, n3037, n3038, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3277,
    n3278, n3279, n3280, n3281, n3282, n3283,
    n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505,
    n3506, n3507, n3508, n3509, n3510, n3511,
    n3512, n3513, n3514, n3515, n3516, n3517,
    n3518, n3519, n3520, n3521, n3522, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722,
    n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927,
    n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951,
    n3952, n3953, n3954, n3955, n3956, n3957,
    n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987,
    n3988, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4017,
    n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4134, n4135, n4136, n4137, n4138,
    n4139, n4140, n4141, n4142, n4143, n4144,
    n4145, n4146, n4147, n4148, n4149, n4150,
    n4151, n4152, n4153, n4154, n4155, n4156,
    n4157, n4158, n4159, n4160, n4161, n4162,
    n4163, n4164, n4165, n4166, n4167, n4168,
    n4169, n4170, n4171, n4172, n4173, n4174,
    n4175, n4176, n4177, n4178, n4179, n4180,
    n4181, n4182, n4183, n4184, n4185, n4186,
    n4187, n4188, n4189, n4190, n4191, n4192,
    n4193, n4194, n4195, n4196, n4197, n4198,
    n4199, n4200, n4201, n4202, n4203, n4204,
    n4205, n4206, n4207, n4208, n4209, n4210,
    n4211, n4212, n4213, n4214, n4215, n4216,
    n4217, n4218, n4219, n4220, n4221, n4222,
    n4223, n4224, n4225, n4226, n4227, n4228,
    n4229, n4230, n4231, n4232, n4233, n4234,
    n4235, n4236, n4237, n4238, n4239, n4240,
    n4241, n4242, n4243, n4244, n4245, n4246,
    n4247, n4248, n4249, n4250, n4251, n4252,
    n4253, n4254, n4255, n4256, n4257, n4258,
    n4259, n4260, n4261, n4262, n4263, n4264,
    n4265, n4266, n4267, n4268, n4269, n4270,
    n4271, n4272, n4273, n4274, n4275, n4276,
    n4277, n4278, n4279, n4280, n4281, n4282,
    n4283, n4284, n4285, n4286, n4287, n4288,
    n4289, n4290, n4291, n4292, n4293, n4294,
    n4295, n4296, n4297, n4298, n4299, n4300,
    n4301, n4302, n4303, n4304, n4305, n4306,
    n4307, n4308, n4309, n4310, n4311, n4312,
    n4313, n4314, n4315, n4316, n4317, n4318,
    n4319, n4320, n4321, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355,
    n4356, n4357, n4358, n4359, n4360, n4361,
    n4362, n4363, n4364, n4365, n4366, n4367,
    n4368, n4369, n4370, n4371, n4372, n4373,
    n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385,
    n4386, n4387, n4388, n4389, n4390, n4391,
    n4392, n4393, n4394, n4395, n4396, n4397,
    n4398, n4399, n4400, n4401, n4402, n4403,
    n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415,
    n4416, n4417, n4418, n4419, n4420, n4421,
    n4422, n4423, n4424, n4425, n4426, n4427,
    n4428, n4429, n4430, n4431, n4432, n4433,
    n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445,
    n4446, n4447, n4448, n4449, n4450, n4451,
    n4452, n4453, n4454, n4455, n4456, n4457,
    n4458, n4459, n4460, n4461, n4462, n4463,
    n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481,
    n4482, n4483, n4484, n4485, n4486, n4487,
    n4488, n4489, n4490, n4491, n4492, n4493,
    n4494, n4495, n4496, n4497, n4498, n4499,
    n4500, n4501, n4502, n4503, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511,
    n4512, n4513, n4514, n4515, n4516, n4517,
    n4518, n4519, n4520, n4521, n4522, n4523,
    n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535,
    n4536, n4537, n4538, n4539, n4540, n4541,
    n4542, n4543, n4544, n4545, n4546, n4547,
    n4548, n4549, n4550, n4551, n4552, n4553,
    n4554, n4555, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4563, n4564, n4565,
    n4566, n4567, n4568, n4569, n4570, n4571,
    n4572, n4573, n4574, n4575, n4576, n4577,
    n4578, n4579, n4580, n4581, n4582, n4583,
    n4584, n4585, n4586, n4587, n4588, n4589,
    n4590, n4591, n4592, n4593, n4594, n4595,
    n4596, n4597, n4598, n4599, n4600, n4601,
    n4602, n4603, n4604, n4605, n4606, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4643, n4644,
    n4645, n4646, n4647, n4648, n4649, n4650,
    n4651, n4652, n4653, n4654, n4655, n4656,
    n4657, n4658, n4659, n4660, n4661, n4662,
    n4663, n4664, n4665, n4666, n4667, n4668,
    n4669, n4670, n4671, n4672, n4673, n4674,
    n4675, n4676, n4677, n4678, n4679, n4680,
    n4681, n4682, n4683, n4684, n4685, n4686,
    n4687, n4688, n4689, n4690, n4691, n4692,
    n4693, n4694, n4695, n4696, n4697, n4698,
    n4699, n4700, n4701, n4702, n4703, n4704,
    n4705, n4706, n4707, n4708, n4709, n4710,
    n4711, n4712, n4713, n4714, n4715, n4716,
    n4717, n4718, n4719, n4720, n4721, n4722,
    n4723, n4724, n4725, n4726, n4727, n4728,
    n4729, n4730, n4731, n4732, n4733, n4734,
    n4735, n4736, n4737, n4738, n4739, n4740,
    n4741, n4742, n4743, n4744, n4745, n4746,
    n4747, n4748, n4749, n4750, n4751, n4752,
    n4753, n4754, n4755, n4756, n4757, n4758,
    n4759, n4760, n4761, n4762, n4763, n4764,
    n4765, n4766, n4767, n4768, n4769, n4770,
    n4771, n4772, n4773, n4774, n4775, n4776,
    n4777, n4778, n4779, n4780, n4781, n4782,
    n4783, n4784, n4785, n4786, n4787, n4788,
    n4789, n4790, n4791, n4792, n4793, n4794,
    n4795, n4796, n4797, n4798, n4799, n4800,
    n4801, n4802, n4803, n4804, n4805, n4806,
    n4807, n4808, n4809, n4810, n4811, n4812,
    n4813, n4814, n4815, n4816, n4817, n4818,
    n4819, n4820, n4821, n4822, n4823, n4824,
    n4825, n4826, n4827, n4828, n4829, n4830,
    n4831, n4832, n4833, n4834, n4835, n4836,
    n4837, n4838, n4839, n4840, n4841, n4842,
    n4843, n4844, n4845, n4846, n4847, n4848,
    n4849, n4850, n4851, n4852, n4853, n4854,
    n4855, n4856, n4857, n4858, n4859, n4860,
    n4861, n4862, n4863, n4864, n4865, n4866,
    n4867, n4868, n4869, n4870, n4871, n4872,
    n4873, n4874, n4875, n4876, n4877, n4878,
    n4879, n4880, n4881, n4882, n4883, n4884,
    n4885, n4886, n4887, n4888, n4889, n4890,
    n4891, n4892, n4893, n4894, n4895, n4896,
    n4897, n4898, n4899, n4900, n4902, n4903,
    n4904, n4905, n4906, n4907, n4908, n4909,
    n4910, n4911, n4912, n4913, n4914, n4915,
    n4916, n4917, n4918, n4919, n4920, n4921,
    n4922, n4923, n4924, n4925, n4926, n4927,
    n4928, n4929, n4930, n4931, n4932, n4933,
    n4934, n4935, n4936, n4937, n4938, n4939,
    n4940, n4941, n4942, n4943, n4944, n4945,
    n4946, n4947, n4948, n4949, n4950, n4951,
    n4952, n4953, n4954, n4955, n4956, n4957,
    n4958, n4959, n4960, n4961, n4962, n4963,
    n4964, n4965, n4966, n4967, n4968, n4969,
    n4970, n4971, n4972, n4973, n4974, n4975,
    n4976, n4977, n4978, n4979, n4980, n4981,
    n4982, n4983, n4984, n4985, n4986, n4987,
    n4988, n4989, n4990, n4991, n4992, n4993,
    n4994, n4995, n4996, n4997, n4998, n4999,
    n5000, n5001, n5002, n5003, n5004, n5005,
    n5006, n5007, n5008, n5009, n5010, n5011,
    n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5050, n5051, n5052, n5053,
    n5054, n5055, n5056, n5057, n5058, n5059,
    n5060, n5061, n5062, n5063, n5064, n5065,
    n5066, n5067, n5068, n5069, n5070, n5071,
    n5072, n5073, n5074, n5075, n5076, n5077,
    n5078, n5079, n5080, n5081, n5082, n5083,
    n5084, n5085, n5086, n5087, n5088, n5089,
    n5090, n5091, n5092, n5093, n5094, n5095,
    n5096, n5097, n5098, n5099, n5100, n5101,
    n5102, n5103, n5104, n5105, n5106, n5107,
    n5108, n5109, n5110, n5111, n5112, n5113,
    n5114, n5115, n5116, n5117, n5118, n5119,
    n5120, n5121, n5122, n5123, n5124, n5125,
    n5126, n5127, n5128, n5129, n5130, n5131,
    n5132, n5133, n5134, n5135, n5136, n5137,
    n5138, n5139, n5140, n5141, n5142, n5143,
    n5144, n5145, n5146, n5147, n5148, n5149,
    n5150, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5160, n5161,
    n5162, n5163, n5164, n5165, n5166, n5167,
    n5168, n5169, n5170, n5171, n5172, n5173,
    n5174, n5175, n5176, n5177, n5178, n5179,
    n5180, n5181, n5182, n5183, n5184, n5185,
    n5186, n5187, n5188, n5189, n5190, n5191,
    n5192, n5193, n5194, n5195, n5196, n5197,
    n5198, n5199, n5200, n5201, n5202, n5203,
    n5204, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372,
    n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390,
    n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402,
    n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414,
    n5415, n5416, n5417, n5418, n5419, n5420,
    n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5436, n5437, n5438,
    n5439, n5440, n5441, n5442, n5443, n5444,
    n5445, n5446, n5447, n5448, n5449, n5450,
    n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5460, n5461, n5462,
    n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5470, n5471, n5472, n5473, n5474,
    n5475, n5476, n5477, n5478, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541,
    n5542, n5543, n5544, n5545, n5546, n5547,
    n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571,
    n5572, n5573, n5574, n5575, n5576, n5577,
    n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601,
    n5602, n5603, n5604, n5605, n5606, n5607,
    n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619,
    n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631,
    n5632, n5633, n5634, n5635, n5636, n5637,
    n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649,
    n5650, n5651, n5652, n5653, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661,
    n5662, n5663, n5664, n5665, n5666, n5667,
    n5668, n5669, n5670, n5671, n5672, n5673,
    n5674, n5675, n5676, n5677, n5678, n5679,
    n5680, n5681, n5682, n5683, n5684, n5685,
    n5686, n5687, n5688, n5689, n5690, n5691,
    n5692, n5693, n5694, n5695, n5696, n5697,
    n5698, n5699, n5700, n5701, n5702, n5703,
    n5704, n5705, n5706, n5707, n5708, n5709,
    n5710, n5711, n5712, n5713, n5714, n5715,
    n5716, n5717, n5718, n5719, n5720, n5721,
    n5722, n5723, n5724, n5725, n5726, n5727,
    n5728, n5729, n5730, n5731, n5732, n5733,
    n5734, n5735, n5736, n5737, n5738, n5739,
    n5740, n5741, n5742, n5743, n5744, n5745,
    n5746, n5747, n5748, n5749, n5750, n5751,
    n5752, n5753, n5754, n5755, n5756, n5757,
    n5758, n5759, n5760, n5761, n5762, n5763,
    n5764, n5765, n5766, n5767, n5768, n5769,
    n5770, n5771, n5772, n5773, n5774, n5775,
    n5776, n5777, n5778, n5779, n5780, n5781,
    n5782, n5783, n5784, n5785, n5786, n5787,
    n5788, n5789, n5790, n5791, n5792, n5793,
    n5794, n5795, n5796, n5797, n5798, n5799,
    n5800, n5801, n5802, n5803, n5804, n5805,
    n5806, n5807, n5808, n5809, n5810, n5811,
    n5812, n5813, n5814, n5815, n5816, n5817,
    n5818, n5819, n5820, n5821, n5822, n5823,
    n5824, n5825, n5826, n5827, n5828, n5829,
    n5830, n5831, n5832, n5833, n5834, n5835,
    n5836, n5837, n5838, n5839, n5840, n5842,
    n5843, n5844, n5845, n5846, n5847, n5848,
    n5849, n5850, n5851, n5852, n5853, n5854,
    n5855, n5856, n5857, n5858, n5859, n5860,
    n5861, n5862, n5863, n5864, n5865, n5866,
    n5867, n5868, n5869, n5870, n5871, n5872,
    n5873, n5874, n5875, n5876, n5877, n5878,
    n5879, n5880, n5881, n5882, n5883, n5884,
    n5885, n5886, n5887, n5888, n5889, n5890,
    n5891, n5892, n5893, n5894, n5895, n5896,
    n5897, n5898, n5899, n5900, n5901, n5902,
    n5903, n5904, n5905, n5906, n5907, n5908,
    n5909, n5910, n5911, n5912, n5913, n5914,
    n5915, n5916, n5917, n5918, n5919, n5920,
    n5921, n5922, n5923, n5924, n5925, n5926,
    n5927, n5928, n5929, n5930, n5931, n5932,
    n5933, n5934, n5935, n5936, n5937, n5938,
    n5939, n5940, n5941, n5942, n5943, n5944,
    n5945, n5946, n5947, n5948, n5949, n5950,
    n5951, n5952, n5953, n5954, n5955, n5956,
    n5957, n5958, n5959, n5960, n5961, n5962,
    n5963, n5964, n5965, n5966, n5967, n5968,
    n5969, n5970, n5971, n5972, n5973, n5974,
    n5975, n5976, n5977, n5978, n5979, n5980,
    n5981, n5982, n5983, n5984, n5985, n5986,
    n5987, n5988, n5989, n5990, n5991, n5992,
    n5993, n5994, n5995, n5996, n5997, n5998,
    n5999, n6000, n6001, n6002, n6003, n6004,
    n6005, n6006, n6007, n6008, n6009, n6010,
    n6011, n6012, n6013, n6014, n6015, n6016,
    n6017, n6018, n6019, n6020, n6021, n6022,
    n6023, n6024, n6025, n6026, n6027, n6028,
    n6029, n6030, n6031, n6032, n6033, n6034,
    n6035, n6036, n6037, n6038, n6039, n6040,
    n6041, n6042, n6043, n6044, n6045, n6046,
    n6047, n6048, n6049, n6050, n6051, n6052,
    n6053, n6054, n6055, n6056, n6057, n6058,
    n6059, n6060, n6061, n6062, n6063, n6064,
    n6065, n6066, n6067, n6068, n6069, n6070,
    n6071, n6072, n6073, n6074, n6075, n6076,
    n6077, n6078, n6079, n6080, n6081, n6082,
    n6083, n6084, n6085, n6086, n6087, n6088,
    n6089, n6090, n6091, n6092, n6093, n6094,
    n6095, n6096, n6097, n6098, n6099, n6100,
    n6101, n6102, n6103, n6104, n6105, n6106,
    n6107, n6108, n6109, n6110, n6111, n6112,
    n6113, n6114, n6115, n6116, n6117, n6118,
    n6119, n6120, n6121, n6122, n6123, n6124,
    n6125, n6126, n6127, n6128, n6129, n6130,
    n6131, n6132, n6133, n6134, n6135, n6136,
    n6137, n6138, n6139, n6140, n6141, n6142,
    n6143, n6144, n6145, n6146, n6147, n6148,
    n6149, n6150, n6151, n6152, n6153, n6154,
    n6155, n6156, n6157, n6158, n6159, n6160,
    n6161, n6162, n6163, n6164, n6165, n6166,
    n6167, n6168, n6169, n6170, n6171, n6172,
    n6173, n6174, n6176, n6177, n6178, n6179,
    n6180, n6181, n6182, n6183, n6184, n6185,
    n6186, n6187, n6188, n6189, n6190, n6191,
    n6192, n6193, n6194, n6195, n6196, n6197,
    n6198, n6199, n6200, n6201, n6202, n6203,
    n6204, n6205, n6206, n6207, n6208, n6209,
    n6210, n6211, n6212, n6213, n6214, n6215,
    n6216, n6217, n6218, n6219, n6220, n6221,
    n6222, n6223, n6224, n6225, n6226, n6227,
    n6228, n6229, n6230, n6231, n6232, n6233,
    n6234, n6235, n6236, n6237, n6238, n6239,
    n6240, n6241, n6242, n6243, n6244, n6245,
    n6246, n6247, n6248, n6249, n6250, n6251,
    n6252, n6253, n6254, n6255, n6256, n6257,
    n6258, n6259, n6260, n6261, n6262, n6263,
    n6264, n6265, n6266, n6267, n6268, n6269,
    n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6277, n6278, n6279, n6280, n6281,
    n6282, n6283, n6284, n6285, n6286, n6287,
    n6288, n6289, n6290, n6291, n6292, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311,
    n6312, n6313, n6314, n6315, n6316, n6317,
    n6318, n6319, n6320, n6321, n6322, n6323,
    n6324, n6325, n6326, n6327, n6328, n6329,
    n6330, n6331, n6332, n6333, n6334, n6335,
    n6336, n6337, n6338, n6339, n6340, n6341,
    n6342, n6343, n6344, n6345, n6346, n6347,
    n6348, n6349, n6350, n6351, n6352, n6353,
    n6354, n6355, n6356, n6357, n6358, n6359,
    n6360, n6361, n6362, n6363, n6364, n6365,
    n6366, n6367, n6368, n6369, n6370, n6371,
    n6372, n6373, n6374, n6375, n6376, n6377,
    n6378, n6379, n6380, n6381, n6382, n6383,
    n6384, n6385, n6386, n6387, n6388, n6389,
    n6390, n6391, n6392, n6393, n6394, n6395,
    n6396, n6397, n6398, n6399, n6400, n6401,
    n6402, n6403, n6404, n6405, n6406, n6407,
    n6408, n6409, n6410, n6411, n6412, n6413,
    n6414, n6415, n6416, n6417, n6418, n6419,
    n6420, n6421, n6422, n6423, n6424, n6425,
    n6426, n6427, n6428, n6429, n6430, n6431,
    n6432, n6433, n6434, n6435, n6436, n6437,
    n6438, n6439, n6440, n6441, n6442, n6443,
    n6444, n6445, n6446, n6447, n6448, n6449,
    n6450, n6451, n6452, n6453, n6454, n6455,
    n6456, n6457, n6458, n6459, n6460, n6461,
    n6462, n6463, n6464, n6465, n6466, n6467,
    n6468, n6469, n6470, n6471, n6472, n6473,
    n6474, n6475, n6476, n6477, n6478, n6479,
    n6480, n6481, n6482, n6483, n6484, n6485,
    n6486, n6487, n6488, n6489, n6490, n6491,
    n6492, n6493, n6494, n6495, n6496, n6497,
    n6498, n6499, n6500, n6501, n6502, n6503,
    n6504, n6505, n6506, n6507, n6508, n6509,
    n6510, n6511, n6512, n6513, n6514, n6515,
    n6516, n6518, n6519, n6520, n6521, n6522,
    n6523, n6524, n6525, n6526, n6527, n6528,
    n6529, n6530, n6531, n6532, n6533, n6534,
    n6535, n6536, n6537, n6538, n6539, n6540,
    n6541, n6542, n6543, n6544, n6545, n6546,
    n6547, n6548, n6549, n6550, n6551, n6552,
    n6553, n6554, n6555, n6556, n6557, n6558,
    n6559, n6560, n6561, n6562, n6563, n6564,
    n6565, n6566, n6567, n6568, n6569, n6570,
    n6571, n6572, n6573, n6574, n6575, n6576,
    n6577, n6578, n6579, n6580, n6581, n6582,
    n6583, n6584, n6585, n6586, n6587, n6588,
    n6589, n6590, n6591, n6592, n6593, n6594,
    n6595, n6596, n6597, n6598, n6599, n6600,
    n6601, n6602, n6603, n6604, n6605, n6606,
    n6607, n6608, n6609, n6610, n6611, n6612,
    n6613, n6614, n6615, n6616, n6617, n6618,
    n6619, n6620, n6621, n6622, n6623, n6624,
    n6625, n6626, n6627, n6628, n6629, n6630,
    n6631, n6632, n6633, n6634, n6635, n6636,
    n6637, n6638, n6639, n6640, n6641, n6642,
    n6643, n6644, n6645, n6646, n6647, n6648,
    n6649, n6650, n6651, n6652, n6653, n6654,
    n6655, n6656, n6657, n6658, n6659, n6660,
    n6661, n6662, n6663, n6664, n6665, n6666,
    n6667, n6668, n6669, n6670, n6671, n6672,
    n6673, n6674, n6675, n6676, n6677, n6678,
    n6679, n6680, n6681, n6682, n6683, n6684,
    n6685, n6686, n6687, n6688, n6689, n6690,
    n6691, n6692, n6693, n6694, n6695, n6696,
    n6697, n6698, n6699, n6700, n6701, n6702,
    n6703, n6704, n6705, n6706, n6707, n6708,
    n6709, n6710, n6711, n6712, n6713, n6714,
    n6715, n6716, n6717, n6718, n6719, n6720,
    n6721, n6722, n6723, n6724, n6725, n6726,
    n6727, n6728, n6729, n6730, n6731, n6732,
    n6733, n6734, n6735, n6736, n6737, n6738,
    n6739, n6740, n6741, n6742, n6743, n6744,
    n6745, n6746, n6747, n6748, n6749, n6750,
    n6751, n6752, n6753, n6754, n6755, n6756,
    n6757, n6758, n6759, n6760, n6761, n6762,
    n6763, n6764, n6765, n6766, n6767, n6768,
    n6769, n6770, n6771, n6772, n6773, n6774,
    n6775, n6776, n6777, n6778, n6779, n6780,
    n6781, n6782, n6783, n6784, n6785, n6786,
    n6787, n6788, n6789, n6790, n6791, n6792,
    n6793, n6794, n6795, n6796, n6797, n6798,
    n6799, n6800, n6801, n6802, n6803, n6804,
    n6805, n6806, n6807, n6808, n6809, n6810,
    n6811, n6812, n6813, n6814, n6815, n6816,
    n6817, n6818, n6819, n6820, n6821, n6822,
    n6823, n6824, n6825, n6826, n6827, n6828,
    n6829, n6830, n6831, n6832, n6833, n6834,
    n6835, n6836, n6837, n6838, n6839, n6840,
    n6841, n6842, n6843, n6844, n6845, n6846,
    n6847, n6848, n6849, n6850, n6851, n6852,
    n6853, n6854, n6855, n6856, n6857, n6858,
    n6859, n6860, n6861, n6862, n6863, n6864,
    n6865, n6866, n6867, n6869, n6870, n6871,
    n6872, n6873, n6874, n6875, n6876, n6877,
    n6878, n6879, n6880, n6881, n6882, n6883,
    n6884, n6885, n6886, n6887, n6888, n6889,
    n6890, n6891, n6892, n6893, n6894, n6895,
    n6896, n6897, n6898, n6899, n6900, n6901,
    n6902, n6903, n6904, n6905, n6906, n6907,
    n6908, n6909, n6910, n6911, n6912, n6913,
    n6914, n6915, n6916, n6917, n6918, n6919,
    n6920, n6921, n6922, n6923, n6924, n6925,
    n6926, n6927, n6928, n6929, n6930, n6931,
    n6932, n6933, n6934, n6935, n6936, n6937,
    n6938, n6939, n6940, n6941, n6942, n6943,
    n6944, n6945, n6946, n6947, n6948, n6949,
    n6950, n6951, n6952, n6953, n6954, n6955,
    n6956, n6957, n6958, n6959, n6960, n6961,
    n6962, n6963, n6964, n6965, n6966, n6967,
    n6968, n6969, n6970, n6971, n6972, n6973,
    n6974, n6975, n6976, n6977, n6978, n6979,
    n6980, n6981, n6982, n6983, n6984, n6985,
    n6986, n6987, n6988, n6989, n6990, n6991,
    n6992, n6993, n6994, n6995, n6996, n6997,
    n6998, n6999, n7000, n7001, n7002, n7003,
    n7004, n7005, n7006, n7007, n7008, n7009,
    n7010, n7011, n7012, n7013, n7014, n7015,
    n7016, n7017, n7018, n7019, n7020, n7021,
    n7022, n7023, n7024, n7025, n7026, n7027,
    n7028, n7029, n7030, n7031, n7032, n7033,
    n7034, n7035, n7036, n7037, n7038, n7039,
    n7040, n7041, n7042, n7043, n7044, n7045,
    n7046, n7047, n7048, n7049, n7050, n7051,
    n7052, n7053, n7054, n7055, n7056, n7057,
    n7058, n7059, n7060, n7061, n7062, n7063,
    n7064, n7065, n7066, n7067, n7068, n7069,
    n7070, n7071, n7072, n7073, n7074, n7075,
    n7076, n7077, n7078, n7079, n7080, n7081,
    n7082, n7083, n7084, n7085, n7086, n7087,
    n7088, n7089, n7090, n7091, n7092, n7093,
    n7094, n7095, n7096, n7097, n7098, n7099,
    n7100, n7101, n7102, n7103, n7104, n7105,
    n7106, n7107, n7108, n7109, n7110, n7111,
    n7112, n7113, n7114, n7115, n7116, n7117,
    n7118, n7119, n7120, n7121, n7122, n7123,
    n7124, n7125, n7126, n7127, n7128, n7129,
    n7130, n7131, n7132, n7133, n7134, n7135,
    n7136, n7137, n7138, n7139, n7140, n7141,
    n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153,
    n7154, n7155, n7156, n7157, n7158, n7159,
    n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171,
    n7172, n7173, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7227, n7228, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370,
    n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400,
    n7401, n7402, n7403, n7404, n7405, n7406,
    n7407, n7408, n7409, n7410, n7411, n7412,
    n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430,
    n7431, n7432, n7433, n7434, n7435, n7436,
    n7437, n7438, n7439, n7440, n7441, n7442,
    n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472,
    n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496,
    n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562,
    n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580,
    n7581, n7582, n7583, n7584, n7585, n7586,
    n7587, n7588, n7589, n7590, n7591, n7592,
    n7593, n7594, n7595, n7596, n7597, n7598,
    n7599, n7600, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7620, n7621, n7622, n7623,
    n7624, n7625, n7626, n7627, n7628, n7629,
    n7630, n7631, n7632, n7633, n7634, n7635,
    n7636, n7637, n7638, n7639, n7640, n7641,
    n7642, n7643, n7644, n7645, n7646, n7647,
    n7648, n7649, n7650, n7651, n7652, n7653,
    n7654, n7655, n7656, n7657, n7658, n7659,
    n7660, n7661, n7662, n7663, n7664, n7665,
    n7666, n7667, n7668, n7669, n7670, n7671,
    n7672, n7673, n7674, n7675, n7676, n7677,
    n7678, n7679, n7680, n7681, n7682, n7683,
    n7684, n7685, n7686, n7687, n7688, n7689,
    n7690, n7691, n7692, n7693, n7694, n7695,
    n7696, n7697, n7698, n7699, n7700, n7701,
    n7702, n7703, n7704, n7705, n7706, n7707,
    n7708, n7709, n7710, n7711, n7712, n7713,
    n7714, n7715, n7716, n7717, n7718, n7719,
    n7720, n7721, n7722, n7723, n7724, n7725,
    n7726, n7727, n7728, n7729, n7730, n7731,
    n7732, n7733, n7734, n7735, n7736, n7737,
    n7738, n7739, n7740, n7741, n7742, n7743,
    n7744, n7745, n7746, n7747, n7748, n7749,
    n7750, n7751, n7752, n7753, n7754, n7755,
    n7756, n7757, n7758, n7759, n7760, n7761,
    n7762, n7763, n7764, n7765, n7766, n7767,
    n7768, n7769, n7770, n7771, n7772, n7773,
    n7774, n7775, n7776, n7777, n7778, n7779,
    n7780, n7781, n7782, n7783, n7784, n7785,
    n7786, n7787, n7788, n7789, n7790, n7791,
    n7792, n7793, n7794, n7795, n7796, n7797,
    n7798, n7799, n7800, n7801, n7802, n7803,
    n7804, n7805, n7806, n7807, n7808, n7809,
    n7810, n7811, n7812, n7813, n7814, n7815,
    n7816, n7817, n7818, n7819, n7820, n7821,
    n7822, n7823, n7824, n7825, n7826, n7827,
    n7828, n7829, n7830, n7831, n7832, n7833,
    n7834, n7835, n7836, n7837, n7838, n7839,
    n7840, n7841, n7842, n7843, n7844, n7845,
    n7846, n7847, n7848, n7849, n7850, n7851,
    n7852, n7853, n7854, n7855, n7856, n7857,
    n7858, n7859, n7860, n7861, n7862, n7863,
    n7864, n7865, n7866, n7867, n7868, n7869,
    n7870, n7871, n7872, n7873, n7874, n7875,
    n7876, n7877, n7878, n7879, n7880, n7881,
    n7882, n7883, n7884, n7885, n7886, n7887,
    n7888, n7889, n7890, n7891, n7892, n7893,
    n7894, n7895, n7896, n7897, n7898, n7899,
    n7900, n7901, n7902, n7903, n7904, n7905,
    n7906, n7907, n7908, n7909, n7910, n7911,
    n7912, n7913, n7914, n7915, n7916, n7917,
    n7918, n7919, n7920, n7921, n7922, n7923,
    n7924, n7925, n7926, n7927, n7928, n7929,
    n7930, n7931, n7932, n7933, n7934, n7935,
    n7936, n7937, n7938, n7939, n7940, n7941,
    n7942, n7943, n7944, n7945, n7946, n7947,
    n7948, n7949, n7950, n7951, n7952, n7953,
    n7954, n7955, n7956, n7957, n7958, n7959,
    n7960, n7961, n7962, n7963, n7964, n7965,
    n7966, n7967, n7968, n7969, n7970, n7971,
    n7972, n7973, n7974, n7975, n7976, n7977,
    n7978, n7979, n7980, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062,
    n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8090, n8091, n8092,
    n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104,
    n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116,
    n8117, n8118, n8119, n8120, n8121, n8122,
    n8123, n8124, n8125, n8126, n8127, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134,
    n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146,
    n8147, n8148, n8149, n8150, n8151, n8152,
    n8153, n8154, n8155, n8156, n8157, n8158,
    n8159, n8160, n8161, n8162, n8163, n8164,
    n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176,
    n8177, n8178, n8179, n8180, n8181, n8182,
    n8183, n8184, n8185, n8186, n8187, n8188,
    n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206,
    n8207, n8208, n8209, n8210, n8211, n8212,
    n8213, n8214, n8215, n8216, n8217, n8218,
    n8219, n8220, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236,
    n8237, n8238, n8239, n8240, n8241, n8242,
    n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8272,
    n8273, n8274, n8275, n8276, n8277, n8278,
    n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296,
    n8297, n8298, n8299, n8300, n8301, n8302,
    n8303, n8304, n8305, n8306, n8307, n8308,
    n8309, n8310, n8311, n8312, n8313, n8314,
    n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326,
    n8327, n8328, n8329, n8330, n8331, n8332,
    n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356,
    n8357, n8358, n8359, n8360, n8361, n8362,
    n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8371, n8372, n8373, n8374, n8375,
    n8376, n8377, n8378, n8379, n8380, n8381,
    n8382, n8383, n8384, n8385, n8386, n8387,
    n8388, n8389, n8390, n8391, n8392, n8393,
    n8394, n8395, n8396, n8397, n8398, n8399,
    n8400, n8401, n8402, n8403, n8404, n8405,
    n8406, n8407, n8408, n8409, n8410, n8411,
    n8412, n8413, n8414, n8415, n8416, n8417,
    n8418, n8419, n8420, n8421, n8422, n8423,
    n8424, n8425, n8426, n8427, n8428, n8429,
    n8430, n8431, n8432, n8433, n8434, n8435,
    n8436, n8437, n8438, n8439, n8440, n8441,
    n8442, n8443, n8444, n8445, n8446, n8447,
    n8448, n8449, n8450, n8451, n8452, n8453,
    n8454, n8455, n8456, n8457, n8458, n8459,
    n8460, n8461, n8462, n8463, n8464, n8465,
    n8466, n8467, n8468, n8469, n8470, n8471,
    n8472, n8473, n8474, n8475, n8476, n8477,
    n8478, n8479, n8480, n8481, n8482, n8483,
    n8484, n8485, n8486, n8487, n8488, n8489,
    n8490, n8491, n8492, n8493, n8494, n8495,
    n8496, n8497, n8498, n8499, n8500, n8501,
    n8502, n8503, n8504, n8505, n8506, n8507,
    n8508, n8509, n8510, n8511, n8512, n8513,
    n8514, n8515, n8516, n8517, n8518, n8519,
    n8520, n8521, n8522, n8523, n8524, n8525,
    n8526, n8527, n8528, n8529, n8530, n8531,
    n8532, n8533, n8534, n8535, n8536, n8537,
    n8538, n8539, n8540, n8541, n8542, n8543,
    n8544, n8545, n8546, n8547, n8548, n8549,
    n8550, n8551, n8552, n8553, n8554, n8555,
    n8556, n8557, n8558, n8559, n8560, n8561,
    n8562, n8563, n8564, n8565, n8566, n8567,
    n8568, n8569, n8570, n8571, n8572, n8573,
    n8574, n8575, n8576, n8577, n8578, n8579,
    n8580, n8581, n8582, n8583, n8584, n8585,
    n8586, n8587, n8588, n8589, n8590, n8591,
    n8592, n8593, n8594, n8595, n8596, n8597,
    n8598, n8599, n8600, n8601, n8602, n8603,
    n8604, n8605, n8606, n8607, n8608, n8609,
    n8610, n8611, n8612, n8613, n8614, n8615,
    n8616, n8617, n8618, n8619, n8620, n8621,
    n8622, n8623, n8624, n8625, n8626, n8627,
    n8628, n8629, n8630, n8631, n8632, n8633,
    n8634, n8635, n8636, n8637, n8638, n8639,
    n8640, n8641, n8642, n8643, n8644, n8645,
    n8646, n8647, n8648, n8649, n8650, n8651,
    n8652, n8653, n8654, n8655, n8656, n8657,
    n8658, n8659, n8660, n8661, n8662, n8663,
    n8664, n8665, n8666, n8667, n8668, n8669,
    n8670, n8671, n8672, n8673, n8674, n8675,
    n8676, n8677, n8678, n8679, n8680, n8681,
    n8682, n8683, n8684, n8685, n8686, n8687,
    n8688, n8689, n8690, n8691, n8692, n8693,
    n8694, n8695, n8696, n8697, n8698, n8699,
    n8700, n8701, n8702, n8703, n8704, n8705,
    n8706, n8707, n8708, n8709, n8710, n8711,
    n8712, n8713, n8714, n8715, n8716, n8717,
    n8718, n8719, n8720, n8721, n8722, n8723,
    n8724, n8725, n8726, n8727, n8728, n8729,
    n8730, n8731, n8732, n8733, n8734, n8735,
    n8736, n8737, n8738, n8739, n8740, n8741,
    n8742, n8743, n8744, n8745, n8746, n8747,
    n8748, n8749, n8750, n8751, n8752, n8753,
    n8754, n8755, n8756, n8757, n8758, n8759,
    n8760, n8761, n8762, n8763, n8764, n8765,
    n8766, n8767, n8768, n8770, n8771, n8772,
    n8773, n8774, n8775, n8776, n8777, n8778,
    n8779, n8780, n8781, n8782, n8783, n8784,
    n8785, n8786, n8787, n8788, n8789, n8790,
    n8791, n8792, n8793, n8794, n8795, n8796,
    n8797, n8798, n8799, n8800, n8801, n8802,
    n8803, n8804, n8805, n8806, n8807, n8808,
    n8809, n8810, n8811, n8812, n8813, n8814,
    n8815, n8816, n8817, n8818, n8819, n8820,
    n8821, n8822, n8823, n8824, n8825, n8826,
    n8827, n8828, n8829, n8830, n8831, n8832,
    n8833, n8834, n8835, n8836, n8837, n8838,
    n8839, n8840, n8841, n8842, n8843, n8844,
    n8845, n8846, n8847, n8848, n8849, n8850,
    n8851, n8852, n8853, n8854, n8855, n8856,
    n8857, n8858, n8859, n8860, n8861, n8862,
    n8863, n8864, n8865, n8866, n8867, n8868,
    n8869, n8870, n8871, n8872, n8873, n8874,
    n8875, n8876, n8877, n8878, n8879, n8880,
    n8881, n8882, n8883, n8884, n8885, n8886,
    n8887, n8888, n8889, n8890, n8891, n8892,
    n8893, n8894, n8895, n8896, n8897, n8898,
    n8899, n8900, n8901, n8902, n8903, n8904,
    n8905, n8906, n8907, n8908, n8909, n8910,
    n8911, n8912, n8913, n8914, n8915, n8916,
    n8917, n8918, n8919, n8920, n8921, n8922,
    n8923, n8924, n8925, n8926, n8927, n8928,
    n8929, n8930, n8931, n8932, n8933, n8934,
    n8935, n8936, n8937, n8938, n8939, n8940,
    n8941, n8942, n8943, n8944, n8945, n8946,
    n8947, n8948, n8949, n8950, n8951, n8952,
    n8953, n8954, n8955, n8956, n8957, n8958,
    n8959, n8960, n8961, n8962, n8963, n8964,
    n8965, n8966, n8967, n8968, n8969, n8970,
    n8971, n8972, n8973, n8974, n8975, n8976,
    n8977, n8978, n8979, n8980, n8981, n8982,
    n8983, n8984, n8985, n8986, n8987, n8988,
    n8989, n8990, n8991, n8992, n8993, n8994,
    n8995, n8996, n8997, n8998, n8999, n9000,
    n9001, n9002, n9003, n9004, n9005, n9006,
    n9007, n9008, n9009, n9010, n9011, n9012,
    n9013, n9014, n9015, n9016, n9017, n9018,
    n9019, n9020, n9021, n9022, n9023, n9024,
    n9025, n9026, n9027, n9028, n9029, n9030,
    n9031, n9032, n9033, n9034, n9035, n9036,
    n9037, n9038, n9039, n9040, n9041, n9042,
    n9043, n9044, n9045, n9046, n9047, n9048,
    n9049, n9050, n9051, n9052, n9053, n9054,
    n9055, n9056, n9057, n9058, n9059, n9060,
    n9061, n9062, n9063, n9064, n9065, n9066,
    n9067, n9068, n9069, n9070, n9071, n9072,
    n9073, n9074, n9075, n9076, n9077, n9078,
    n9079, n9080, n9081, n9082, n9083, n9084,
    n9085, n9086, n9087, n9088, n9089, n9090,
    n9091, n9092, n9093, n9094, n9095, n9096,
    n9097, n9098, n9099, n9100, n9101, n9102,
    n9103, n9104, n9105, n9106, n9107, n9108,
    n9109, n9110, n9111, n9112, n9113, n9114,
    n9115, n9116, n9117, n9118, n9119, n9120,
    n9121, n9122, n9123, n9124, n9125, n9126,
    n9127, n9128, n9129, n9130, n9131, n9132,
    n9133, n9134, n9135, n9136, n9137, n9138,
    n9139, n9140, n9141, n9142, n9143, n9144,
    n9145, n9146, n9147, n9148, n9149, n9150,
    n9151, n9152, n9153, n9154, n9155, n9156,
    n9157, n9158, n9159, n9160, n9161, n9162,
    n9163, n9164, n9165, n9166, n9167, n9168,
    n9169, n9170, n9171, n9172, n9173, n9174,
    n9175, n9176, n9177, n9178, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271,
    n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289,
    n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301,
    n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319,
    n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331,
    n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349,
    n9350, n9351, n9352, n9353, n9354, n9355,
    n9356, n9357, n9358, n9359, n9360, n9361,
    n9362, n9363, n9364, n9365, n9366, n9367,
    n9368, n9369, n9370, n9371, n9372, n9373,
    n9374, n9375, n9376, n9377, n9378, n9379,
    n9380, n9381, n9382, n9383, n9384, n9385,
    n9386, n9387, n9388, n9389, n9390, n9391,
    n9392, n9393, n9394, n9395, n9396, n9397,
    n9398, n9399, n9400, n9401, n9402, n9403,
    n9404, n9405, n9406, n9407, n9408, n9409,
    n9410, n9411, n9412, n9413, n9414, n9415,
    n9416, n9417, n9418, n9419, n9420, n9421,
    n9422, n9423, n9424, n9425, n9426, n9427,
    n9428, n9429, n9430, n9431, n9432, n9433,
    n9434, n9435, n9436, n9437, n9438, n9439,
    n9440, n9441, n9442, n9443, n9444, n9445,
    n9446, n9447, n9448, n9449, n9450, n9451,
    n9452, n9453, n9454, n9455, n9456, n9457,
    n9458, n9459, n9460, n9461, n9462, n9463,
    n9464, n9465, n9466, n9467, n9468, n9469,
    n9470, n9471, n9472, n9473, n9474, n9475,
    n9476, n9477, n9478, n9479, n9480, n9481,
    n9482, n9483, n9484, n9485, n9486, n9487,
    n9488, n9489, n9490, n9491, n9492, n9493,
    n9494, n9495, n9496, n9497, n9498, n9499,
    n9500, n9501, n9502, n9503, n9504, n9505,
    n9506, n9507, n9508, n9509, n9510, n9511,
    n9512, n9513, n9514, n9515, n9516, n9517,
    n9518, n9519, n9520, n9521, n9522, n9523,
    n9524, n9525, n9526, n9527, n9528, n9529,
    n9530, n9531, n9532, n9533, n9534, n9535,
    n9536, n9537, n9538, n9539, n9540, n9541,
    n9542, n9543, n9544, n9545, n9546, n9547,
    n9548, n9549, n9550, n9551, n9552, n9553,
    n9554, n9555, n9556, n9557, n9558, n9559,
    n9560, n9561, n9562, n9563, n9564, n9565,
    n9566, n9567, n9568, n9569, n9570, n9571,
    n9572, n9573, n9574, n9575, n9576, n9577,
    n9578, n9579, n9580, n9581, n9582, n9583,
    n9584, n9585, n9586, n9587, n9588, n9589,
    n9590, n9591, n9592, n9593, n9594, n9595,
    n9596, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10025, n10026, n10027, n10028, n10029,
    n10030, n10031, n10032, n10033, n10034, n10035,
    n10036, n10037, n10038, n10039, n10040, n10041,
    n10042, n10043, n10044, n10045, n10046, n10047,
    n10048, n10049, n10050, n10051, n10052, n10053,
    n10054, n10055, n10056, n10057, n10058, n10059,
    n10060, n10061, n10062, n10063, n10064, n10065,
    n10066, n10067, n10068, n10069, n10070, n10071,
    n10072, n10073, n10074, n10075, n10076, n10077,
    n10078, n10079, n10080, n10081, n10082, n10083,
    n10084, n10085, n10086, n10087, n10088, n10089,
    n10090, n10091, n10092, n10093, n10094, n10095,
    n10096, n10097, n10098, n10099, n10100, n10101,
    n10102, n10103, n10104, n10105, n10106, n10107,
    n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119,
    n10120, n10121, n10122, n10123, n10124, n10125,
    n10126, n10127, n10128, n10129, n10130, n10131,
    n10132, n10133, n10134, n10135, n10136, n10137,
    n10138, n10139, n10140, n10141, n10142, n10143,
    n10144, n10145, n10146, n10147, n10148, n10149,
    n10150, n10151, n10152, n10153, n10154, n10155,
    n10156, n10157, n10158, n10159, n10160, n10161,
    n10162, n10163, n10164, n10165, n10166, n10167,
    n10168, n10169, n10170, n10171, n10172, n10173,
    n10174, n10175, n10176, n10177, n10178, n10179,
    n10180, n10181, n10182, n10183, n10184, n10185,
    n10186, n10187, n10188, n10189, n10190, n10191,
    n10192, n10193, n10194, n10195, n10196, n10197,
    n10198, n10199, n10200, n10201, n10202, n10203,
    n10204, n10205, n10206, n10207, n10208, n10209,
    n10210, n10211, n10212, n10213, n10214, n10215,
    n10216, n10217, n10218, n10219, n10220, n10221,
    n10222, n10223, n10224, n10225, n10226, n10227,
    n10228, n10229, n10230, n10231, n10232, n10233,
    n10234, n10235, n10236, n10237, n10238, n10239,
    n10240, n10241, n10242, n10243, n10244, n10245,
    n10246, n10247, n10248, n10249, n10250, n10251,
    n10252, n10253, n10254, n10255, n10256, n10257,
    n10258, n10259, n10260, n10261, n10262, n10263,
    n10264, n10265, n10266, n10267, n10268, n10269,
    n10270, n10271, n10272, n10273, n10274, n10275,
    n10276, n10277, n10278, n10279, n10280, n10281,
    n10282, n10283, n10284, n10285, n10286, n10287,
    n10288, n10289, n10290, n10291, n10292, n10293,
    n10294, n10295, n10296, n10297, n10298, n10299,
    n10300, n10301, n10302, n10303, n10304, n10305,
    n10306, n10307, n10308, n10309, n10310, n10311,
    n10312, n10313, n10314, n10315, n10316, n10317,
    n10318, n10319, n10320, n10321, n10322, n10323,
    n10324, n10325, n10326, n10327, n10328, n10329,
    n10330, n10331, n10332, n10333, n10334, n10335,
    n10336, n10337, n10338, n10339, n10340, n10341,
    n10342, n10343, n10344, n10345, n10346, n10347,
    n10348, n10349, n10350, n10351, n10352, n10353,
    n10354, n10355, n10356, n10357, n10358, n10359,
    n10360, n10361, n10362, n10363, n10364, n10365,
    n10366, n10367, n10368, n10369, n10370, n10371,
    n10372, n10373, n10374, n10375, n10376, n10377,
    n10378, n10379, n10380, n10381, n10382, n10383,
    n10384, n10385, n10386, n10387, n10388, n10389,
    n10390, n10391, n10392, n10393, n10394, n10395,
    n10396, n10397, n10398, n10399, n10400, n10401,
    n10402, n10403, n10404, n10405, n10406, n10407,
    n10408, n10409, n10410, n10411, n10412, n10413,
    n10414, n10415, n10416, n10417, n10418, n10419,
    n10420, n10421, n10422, n10423, n10424, n10425,
    n10426, n10427, n10428, n10429, n10430, n10431,
    n10432, n10433, n10434, n10435, n10436, n10437,
    n10438, n10439, n10440, n10441, n10442, n10443,
    n10444, n10445, n10446, n10447, n10448, n10449,
    n10450, n10451, n10452, n10453, n10454, n10455,
    n10456, n10457, n10458, n10459, n10460, n10462,
    n10463, n10464, n10465, n10466, n10467, n10468,
    n10469, n10470, n10471, n10472, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10480,
    n10481, n10482, n10483, n10484, n10485, n10486,
    n10487, n10488, n10489, n10490, n10491, n10492,
    n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504,
    n10505, n10506, n10507, n10508, n10509, n10510,
    n10511, n10512, n10513, n10514, n10515, n10516,
    n10517, n10518, n10519, n10520, n10521, n10522,
    n10523, n10524, n10525, n10526, n10527, n10528,
    n10529, n10530, n10531, n10532, n10533, n10534,
    n10535, n10536, n10537, n10538, n10539, n10540,
    n10541, n10542, n10543, n10544, n10545, n10546,
    n10547, n10548, n10549, n10550, n10551, n10552,
    n10553, n10554, n10555, n10556, n10557, n10558,
    n10559, n10560, n10561, n10562, n10563, n10564,
    n10565, n10566, n10567, n10568, n10569, n10570,
    n10571, n10572, n10573, n10574, n10575, n10576,
    n10577, n10578, n10579, n10580, n10581, n10582,
    n10583, n10584, n10585, n10586, n10587, n10588,
    n10589, n10590, n10591, n10592, n10593, n10594,
    n10595, n10596, n10597, n10598, n10599, n10600,
    n10601, n10602, n10603, n10604, n10605, n10606,
    n10607, n10608, n10609, n10610, n10611, n10612,
    n10613, n10614, n10615, n10616, n10617, n10618,
    n10619, n10620, n10621, n10622, n10623, n10624,
    n10625, n10626, n10627, n10628, n10629, n10630,
    n10631, n10632, n10633, n10634, n10635, n10636,
    n10637, n10638, n10639, n10640, n10641, n10642,
    n10643, n10644, n10645, n10646, n10647, n10648,
    n10649, n10650, n10651, n10652, n10653, n10654,
    n10655, n10656, n10657, n10658, n10659, n10660,
    n10661, n10662, n10663, n10664, n10665, n10666,
    n10667, n10668, n10669, n10670, n10671, n10672,
    n10673, n10674, n10675, n10676, n10677, n10678,
    n10679, n10680, n10681, n10682, n10683, n10684,
    n10685, n10686, n10687, n10688, n10689, n10690,
    n10691, n10692, n10693, n10694, n10695, n10696,
    n10697, n10698, n10699, n10700, n10701, n10702,
    n10703, n10704, n10705, n10706, n10707, n10708,
    n10709, n10710, n10711, n10712, n10713, n10714,
    n10715, n10716, n10717, n10718, n10719, n10720,
    n10721, n10722, n10723, n10724, n10725, n10726,
    n10727, n10728, n10729, n10730, n10731, n10732,
    n10733, n10734, n10735, n10736, n10737, n10738,
    n10739, n10740, n10741, n10742, n10743, n10744,
    n10745, n10746, n10747, n10748, n10749, n10750,
    n10751, n10752, n10753, n10754, n10755, n10756,
    n10757, n10758, n10759, n10760, n10761, n10762,
    n10763, n10764, n10765, n10766, n10767, n10768,
    n10769, n10770, n10771, n10772, n10773, n10774,
    n10775, n10776, n10777, n10778, n10779, n10780,
    n10781, n10782, n10783, n10784, n10785, n10786,
    n10787, n10788, n10789, n10790, n10791, n10792,
    n10793, n10794, n10795, n10796, n10797, n10798,
    n10799, n10800, n10801, n10802, n10803, n10804,
    n10805, n10806, n10807, n10808, n10809, n10810,
    n10811, n10812, n10813, n10814, n10815, n10816,
    n10817, n10818, n10819, n10820, n10821, n10822,
    n10823, n10824, n10825, n10826, n10827, n10828,
    n10829, n10830, n10831, n10832, n10833, n10834,
    n10835, n10836, n10837, n10838, n10839, n10840,
    n10841, n10842, n10843, n10844, n10845, n10846,
    n10847, n10848, n10849, n10850, n10851, n10852,
    n10853, n10854, n10855, n10856, n10857, n10858,
    n10859, n10860, n10861, n10862, n10863, n10864,
    n10865, n10866, n10867, n10868, n10869, n10870,
    n10871, n10872, n10873, n10874, n10875, n10876,
    n10877, n10878, n10879, n10880, n10881, n10882,
    n10883, n10884, n10885, n10886, n10887, n10888,
    n10889, n10890, n10891, n10892, n10893, n10894,
    n10895, n10896, n10897, n10898, n10899, n10900,
    n10901, n10902, n10903, n10904, n10905, n10906,
    n10907, n10908, n10910, n10911, n10912, n10913,
    n10914, n10915, n10916, n10917, n10918, n10919,
    n10920, n10921, n10922, n10923, n10924, n10925,
    n10926, n10927, n10928, n10929, n10930, n10931,
    n10932, n10933, n10934, n10935, n10936, n10937,
    n10938, n10939, n10940, n10941, n10942, n10943,
    n10944, n10945, n10946, n10947, n10948, n10949,
    n10950, n10951, n10952, n10953, n10954, n10955,
    n10956, n10957, n10958, n10959, n10960, n10961,
    n10962, n10963, n10964, n10965, n10966, n10967,
    n10968, n10969, n10970, n10971, n10972, n10973,
    n10974, n10975, n10976, n10977, n10978, n10979,
    n10980, n10981, n10982, n10983, n10984, n10985,
    n10986, n10987, n10988, n10989, n10990, n10991,
    n10992, n10993, n10994, n10995, n10996, n10997,
    n10998, n10999, n11000, n11001, n11002, n11003,
    n11004, n11005, n11006, n11007, n11008, n11009,
    n11010, n11011, n11012, n11013, n11014, n11015,
    n11016, n11017, n11018, n11019, n11020, n11021,
    n11022, n11023, n11024, n11025, n11026, n11027,
    n11028, n11029, n11030, n11031, n11032, n11033,
    n11034, n11035, n11036, n11037, n11038, n11039,
    n11040, n11041, n11042, n11043, n11044, n11045,
    n11046, n11047, n11048, n11049, n11050, n11051,
    n11052, n11053, n11054, n11055, n11056, n11057,
    n11058, n11059, n11060, n11061, n11062, n11063,
    n11064, n11065, n11066, n11067, n11068, n11069,
    n11070, n11071, n11072, n11073, n11074, n11075,
    n11076, n11077, n11078, n11079, n11080, n11081,
    n11082, n11083, n11084, n11085, n11086, n11087,
    n11088, n11089, n11090, n11091, n11092, n11093,
    n11094, n11095, n11096, n11097, n11098, n11099,
    n11100, n11101, n11102, n11103, n11104, n11105,
    n11106, n11107, n11108, n11109, n11110, n11111,
    n11112, n11113, n11114, n11115, n11116, n11117,
    n11118, n11119, n11120, n11121, n11122, n11123,
    n11124, n11125, n11126, n11127, n11128, n11129,
    n11130, n11131, n11132, n11133, n11134, n11135,
    n11136, n11137, n11138, n11139, n11140, n11141,
    n11142, n11143, n11144, n11145, n11146, n11147,
    n11148, n11149, n11150, n11151, n11152, n11153,
    n11154, n11155, n11156, n11157, n11158, n11159,
    n11160, n11161, n11162, n11163, n11164, n11165,
    n11166, n11167, n11168, n11169, n11170, n11171,
    n11172, n11173, n11174, n11175, n11176, n11177,
    n11178, n11179, n11180, n11181, n11182, n11183,
    n11184, n11185, n11186, n11187, n11188, n11189,
    n11190, n11191, n11192, n11193, n11194, n11195,
    n11196, n11197, n11198, n11199, n11200, n11201,
    n11202, n11203, n11204, n11205, n11206, n11207,
    n11208, n11209, n11210, n11211, n11212, n11213,
    n11214, n11215, n11216, n11217, n11218, n11219,
    n11220, n11221, n11222, n11223, n11224, n11225,
    n11226, n11227, n11228, n11229, n11230, n11231,
    n11232, n11233, n11234, n11235, n11236, n11237,
    n11238, n11239, n11240, n11241, n11242, n11243,
    n11244, n11245, n11246, n11247, n11248, n11249,
    n11250, n11251, n11252, n11253, n11254, n11255,
    n11256, n11257, n11258, n11259, n11260, n11261,
    n11262, n11263, n11264, n11265, n11266, n11267,
    n11268, n11269, n11270, n11271, n11272, n11273,
    n11274, n11275, n11276, n11277, n11278, n11279,
    n11280, n11281, n11282, n11283, n11284, n11285,
    n11286, n11287, n11288, n11289, n11290, n11291,
    n11292, n11293, n11294, n11295, n11296, n11297,
    n11298, n11299, n11300, n11301, n11302, n11303,
    n11304, n11305, n11306, n11307, n11308, n11309,
    n11310, n11311, n11312, n11313, n11314, n11315,
    n11316, n11317, n11318, n11319, n11320, n11321,
    n11322, n11323, n11324, n11325, n11326, n11327,
    n11328, n11329, n11330, n11331, n11332, n11333,
    n11334, n11335, n11336, n11337, n11338, n11339,
    n11340, n11341, n11342, n11343, n11344, n11345,
    n11346, n11347, n11348, n11349, n11350, n11351,
    n11352, n11353, n11354, n11355, n11356, n11357,
    n11358, n11359, n11360, n11361, n11362, n11363,
    n11364, n11366, n11367, n11368, n11369, n11370,
    n11371, n11372, n11373, n11374, n11375, n11376,
    n11377, n11378, n11379, n11380, n11381, n11382,
    n11383, n11384, n11385, n11386, n11387, n11388,
    n11389, n11390, n11391, n11392, n11393, n11394,
    n11395, n11396, n11397, n11398, n11399, n11400,
    n11401, n11402, n11403, n11404, n11405, n11406,
    n11407, n11408, n11409, n11410, n11411, n11412,
    n11413, n11414, n11415, n11416, n11417, n11418,
    n11419, n11420, n11421, n11422, n11423, n11424,
    n11425, n11426, n11427, n11428, n11429, n11430,
    n11431, n11432, n11433, n11434, n11435, n11436,
    n11437, n11438, n11439, n11440, n11441, n11442,
    n11443, n11444, n11445, n11446, n11447, n11448,
    n11449, n11450, n11451, n11452, n11453, n11454,
    n11455, n11456, n11457, n11458, n11459, n11460,
    n11461, n11462, n11463, n11464, n11465, n11466,
    n11467, n11468, n11469, n11470, n11471, n11472,
    n11473, n11474, n11475, n11476, n11477, n11478,
    n11479, n11480, n11481, n11482, n11483, n11484,
    n11485, n11486, n11487, n11488, n11489, n11490,
    n11491, n11492, n11493, n11494, n11495, n11496,
    n11497, n11498, n11499, n11500, n11501, n11502,
    n11503, n11504, n11505, n11506, n11507, n11508,
    n11509, n11510, n11511, n11512, n11513, n11514,
    n11515, n11516, n11517, n11518, n11519, n11520,
    n11521, n11522, n11523, n11524, n11525, n11526,
    n11527, n11528, n11529, n11530, n11531, n11532,
    n11533, n11534, n11535, n11536, n11537, n11538,
    n11539, n11540, n11541, n11542, n11543, n11544,
    n11545, n11546, n11547, n11548, n11549, n11550,
    n11551, n11552, n11553, n11554, n11555, n11556,
    n11557, n11558, n11559, n11560, n11561, n11562,
    n11563, n11564, n11565, n11566, n11567, n11568,
    n11569, n11570, n11571, n11572, n11573, n11574,
    n11575, n11576, n11577, n11578, n11579, n11580,
    n11581, n11582, n11583, n11584, n11585, n11586,
    n11587, n11588, n11589, n11590, n11591, n11592,
    n11593, n11594, n11595, n11596, n11597, n11598,
    n11599, n11600, n11601, n11602, n11603, n11604,
    n11605, n11606, n11607, n11608, n11609, n11610,
    n11611, n11612, n11613, n11614, n11615, n11616,
    n11617, n11618, n11619, n11620, n11621, n11622,
    n11623, n11624, n11625, n11626, n11627, n11628,
    n11629, n11630, n11631, n11632, n11633, n11634,
    n11635, n11636, n11637, n11638, n11639, n11640,
    n11641, n11642, n11643, n11644, n11645, n11646,
    n11647, n11648, n11649, n11650, n11651, n11652,
    n11653, n11654, n11655, n11656, n11657, n11658,
    n11659, n11660, n11661, n11662, n11663, n11664,
    n11665, n11666, n11667, n11668, n11669, n11670,
    n11671, n11672, n11673, n11674, n11675, n11676,
    n11677, n11678, n11679, n11680, n11681, n11682,
    n11683, n11684, n11685, n11686, n11687, n11688,
    n11689, n11690, n11691, n11692, n11693, n11694,
    n11695, n11696, n11697, n11698, n11699, n11700,
    n11701, n11702, n11703, n11704, n11705, n11706,
    n11707, n11708, n11709, n11710, n11711, n11712,
    n11713, n11714, n11715, n11716, n11717, n11718,
    n11719, n11720, n11721, n11722, n11723, n11724,
    n11725, n11726, n11727, n11728, n11729, n11730,
    n11731, n11732, n11733, n11734, n11735, n11736,
    n11737, n11738, n11739, n11740, n11741, n11742,
    n11743, n11744, n11745, n11746, n11747, n11748,
    n11749, n11750, n11751, n11752, n11753, n11754,
    n11755, n11756, n11757, n11758, n11759, n11760,
    n11761, n11762, n11763, n11764, n11765, n11766,
    n11767, n11768, n11769, n11770, n11771, n11772,
    n11773, n11774, n11775, n11776, n11777, n11778,
    n11779, n11780, n11781, n11782, n11783, n11784,
    n11785, n11786, n11787, n11788, n11789, n11790,
    n11791, n11792, n11793, n11794, n11795, n11796,
    n11797, n11798, n11799, n11800, n11801, n11802,
    n11803, n11804, n11805, n11806, n11807, n11808,
    n11809, n11810, n11811, n11812, n11813, n11814,
    n11815, n11816, n11817, n11818, n11819, n11820,
    n11821, n11822, n11823, n11824, n11825, n11826,
    n11827, n11828, n11829, n11831, n11832, n11833,
    n11834, n11835, n11836, n11837, n11838, n11839,
    n11840, n11841, n11842, n11843, n11844, n11845,
    n11846, n11847, n11848, n11849, n11850, n11851,
    n11852, n11853, n11854, n11855, n11856, n11857,
    n11858, n11859, n11860, n11861, n11862, n11863,
    n11864, n11865, n11866, n11867, n11868, n11869,
    n11870, n11871, n11872, n11873, n11874, n11875,
    n11876, n11877, n11878, n11879, n11880, n11881,
    n11882, n11883, n11884, n11885, n11886, n11887,
    n11888, n11889, n11890, n11891, n11892, n11893,
    n11894, n11895, n11896, n11897, n11898, n11899,
    n11900, n11901, n11902, n11903, n11904, n11905,
    n11906, n11907, n11908, n11909, n11910, n11911,
    n11912, n11913, n11914, n11915, n11916, n11917,
    n11918, n11919, n11920, n11921, n11922, n11923,
    n11924, n11925, n11926, n11927, n11928, n11929,
    n11930, n11931, n11932, n11933, n11934, n11935,
    n11936, n11937, n11938, n11939, n11940, n11941,
    n11942, n11943, n11944, n11945, n11946, n11947,
    n11948, n11949, n11950, n11951, n11952, n11953,
    n11954, n11955, n11956, n11957, n11958, n11959,
    n11960, n11961, n11962, n11963, n11964, n11965,
    n11966, n11967, n11968, n11969, n11970, n11971,
    n11972, n11973, n11974, n11975, n11976, n11977,
    n11978, n11979, n11980, n11981, n11982, n11983,
    n11984, n11985, n11986, n11987, n11988, n11989,
    n11990, n11991, n11992, n11993, n11994, n11995,
    n11996, n11997, n11998, n11999, n12000, n12001,
    n12002, n12003, n12004, n12005, n12006, n12007,
    n12008, n12009, n12010, n12011, n12012, n12013,
    n12014, n12015, n12016, n12017, n12018, n12019,
    n12020, n12021, n12022, n12023, n12024, n12025,
    n12026, n12027, n12028, n12029, n12030, n12031,
    n12032, n12033, n12034, n12035, n12036, n12037,
    n12038, n12039, n12040, n12041, n12042, n12043,
    n12044, n12045, n12046, n12047, n12048, n12049,
    n12050, n12051, n12052, n12053, n12054, n12055,
    n12056, n12057, n12058, n12059, n12060, n12061,
    n12062, n12063, n12064, n12065, n12066, n12067,
    n12068, n12069, n12070, n12071, n12072, n12073,
    n12074, n12075, n12076, n12077, n12078, n12079,
    n12080, n12081, n12082, n12083, n12084, n12085,
    n12086, n12087, n12088, n12089, n12090, n12091,
    n12092, n12093, n12094, n12095, n12096, n12097,
    n12098, n12099, n12100, n12101, n12102, n12103,
    n12104, n12105, n12106, n12107, n12108, n12109,
    n12110, n12111, n12112, n12113, n12114, n12115,
    n12116, n12117, n12118, n12119, n12120, n12121,
    n12122, n12123, n12124, n12125, n12126, n12127,
    n12128, n12129, n12130, n12131, n12132, n12133,
    n12134, n12135, n12136, n12137, n12138, n12139,
    n12140, n12141, n12142, n12143, n12144, n12145,
    n12146, n12147, n12148, n12149, n12150, n12151,
    n12152, n12153, n12154, n12155, n12156, n12157,
    n12158, n12159, n12160, n12161, n12162, n12163,
    n12164, n12165, n12166, n12167, n12168, n12169,
    n12170, n12171, n12172, n12173, n12174, n12175,
    n12176, n12177, n12178, n12179, n12180, n12181,
    n12182, n12183, n12184, n12185, n12186, n12187,
    n12188, n12189, n12190, n12191, n12192, n12193,
    n12194, n12195, n12196, n12197, n12198, n12199,
    n12200, n12201, n12202, n12203, n12204, n12205,
    n12206, n12207, n12208, n12209, n12210, n12211,
    n12212, n12213, n12214, n12215, n12216, n12217,
    n12218, n12219, n12220, n12221, n12222, n12223,
    n12224, n12225, n12226, n12227, n12228, n12229,
    n12230, n12231, n12232, n12233, n12234, n12235,
    n12236, n12237, n12238, n12239, n12240, n12241,
    n12242, n12243, n12244, n12245, n12246, n12247,
    n12248, n12249, n12250, n12251, n12252, n12253,
    n12254, n12255, n12256, n12257, n12258, n12259,
    n12260, n12261, n12262, n12263, n12264, n12265,
    n12266, n12267, n12268, n12269, n12270, n12271,
    n12272, n12273, n12274, n12275, n12276, n12277,
    n12278, n12279, n12280, n12281, n12282, n12283,
    n12284, n12285, n12286, n12287, n12288, n12289,
    n12290, n12291, n12292, n12293, n12294, n12295,
    n12296, n12297, n12298, n12299, n12300, n12301,
    n12302, n12303, n12304, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314,
    n12315, n12316, n12317, n12318, n12319, n12320,
    n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12340, n12341, n12342, n12343, n12344,
    n12345, n12346, n12347, n12348, n12349, n12350,
    n12351, n12352, n12353, n12354, n12355, n12356,
    n12357, n12358, n12359, n12360, n12361, n12362,
    n12363, n12364, n12365, n12366, n12367, n12368,
    n12369, n12370, n12371, n12372, n12373, n12374,
    n12375, n12376, n12377, n12378, n12379, n12380,
    n12381, n12382, n12383, n12384, n12385, n12386,
    n12387, n12388, n12389, n12390, n12391, n12392,
    n12393, n12394, n12395, n12396, n12397, n12398,
    n12399, n12400, n12401, n12402, n12403, n12404,
    n12405, n12406, n12407, n12408, n12409, n12410,
    n12411, n12412, n12413, n12414, n12415, n12416,
    n12417, n12418, n12419, n12420, n12421, n12422,
    n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434,
    n12435, n12436, n12437, n12438, n12439, n12440,
    n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452,
    n12453, n12454, n12455, n12456, n12457, n12458,
    n12459, n12460, n12461, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470,
    n12471, n12472, n12473, n12474, n12475, n12476,
    n12477, n12478, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488,
    n12489, n12490, n12491, n12492, n12493, n12494,
    n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506,
    n12507, n12508, n12509, n12510, n12511, n12512,
    n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524,
    n12525, n12526, n12527, n12528, n12529, n12530,
    n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542,
    n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560,
    n12561, n12562, n12563, n12564, n12565, n12566,
    n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578,
    n12579, n12580, n12581, n12582, n12583, n12584,
    n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596,
    n12597, n12598, n12599, n12600, n12601, n12602,
    n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614,
    n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632,
    n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650,
    n12651, n12652, n12653, n12654, n12655, n12656,
    n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668,
    n12669, n12670, n12671, n12672, n12673, n12674,
    n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12691, n12692,
    n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704,
    n12705, n12706, n12707, n12708, n12709, n12710,
    n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722,
    n12723, n12724, n12725, n12726, n12727, n12728,
    n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740,
    n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758,
    n12759, n12760, n12761, n12762, n12763, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776,
    n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12792, n12793, n12794, n12795,
    n12796, n12797, n12798, n12799, n12800, n12801,
    n12802, n12803, n12804, n12805, n12806, n12807,
    n12808, n12809, n12810, n12811, n12812, n12813,
    n12814, n12815, n12816, n12817, n12818, n12819,
    n12820, n12821, n12822, n12823, n12824, n12825,
    n12826, n12827, n12828, n12829, n12830, n12831,
    n12832, n12833, n12834, n12835, n12836, n12837,
    n12838, n12839, n12840, n12841, n12842, n12843,
    n12844, n12845, n12846, n12847, n12848, n12849,
    n12850, n12851, n12852, n12853, n12854, n12855,
    n12856, n12857, n12858, n12859, n12860, n12861,
    n12862, n12863, n12864, n12865, n12866, n12867,
    n12868, n12869, n12870, n12871, n12872, n12873,
    n12874, n12875, n12876, n12877, n12878, n12879,
    n12880, n12881, n12882, n12883, n12884, n12885,
    n12886, n12887, n12888, n12889, n12890, n12891,
    n12892, n12893, n12894, n12895, n12896, n12897,
    n12898, n12899, n12900, n12901, n12902, n12903,
    n12904, n12905, n12906, n12907, n12908, n12909,
    n12910, n12911, n12912, n12913, n12914, n12915,
    n12916, n12917, n12918, n12919, n12920, n12921,
    n12922, n12923, n12924, n12925, n12926, n12927,
    n12928, n12929, n12930, n12931, n12932, n12933,
    n12934, n12935, n12936, n12937, n12938, n12939,
    n12940, n12941, n12942, n12943, n12944, n12945,
    n12946, n12947, n12948, n12949, n12950, n12951,
    n12952, n12953, n12954, n12955, n12956, n12957,
    n12958, n12959, n12960, n12961, n12962, n12963,
    n12964, n12965, n12966, n12967, n12968, n12969,
    n12970, n12971, n12972, n12973, n12974, n12975,
    n12976, n12977, n12978, n12979, n12980, n12981,
    n12982, n12983, n12984, n12985, n12986, n12987,
    n12988, n12989, n12990, n12991, n12992, n12993,
    n12994, n12995, n12996, n12997, n12998, n12999,
    n13000, n13001, n13002, n13003, n13004, n13005,
    n13006, n13007, n13008, n13009, n13010, n13011,
    n13012, n13013, n13014, n13015, n13016, n13017,
    n13018, n13019, n13020, n13021, n13022, n13023,
    n13024, n13025, n13026, n13027, n13028, n13029,
    n13030, n13031, n13032, n13033, n13034, n13035,
    n13036, n13037, n13038, n13039, n13040, n13041,
    n13042, n13043, n13044, n13045, n13046, n13047,
    n13048, n13049, n13050, n13051, n13052, n13053,
    n13054, n13055, n13056, n13057, n13058, n13059,
    n13060, n13061, n13062, n13063, n13064, n13065,
    n13066, n13067, n13068, n13069, n13070, n13071,
    n13072, n13073, n13074, n13075, n13076, n13077,
    n13078, n13079, n13080, n13081, n13082, n13083,
    n13084, n13085, n13086, n13087, n13088, n13089,
    n13090, n13091, n13092, n13093, n13094, n13095,
    n13096, n13097, n13098, n13099, n13100, n13101,
    n13102, n13103, n13104, n13105, n13106, n13107,
    n13108, n13109, n13110, n13111, n13112, n13113,
    n13114, n13115, n13116, n13117, n13118, n13119,
    n13120, n13121, n13122, n13123, n13124, n13125,
    n13126, n13127, n13128, n13129, n13130, n13131,
    n13132, n13133, n13134, n13135, n13136, n13137,
    n13138, n13139, n13140, n13141, n13142, n13143,
    n13144, n13145, n13146, n13147, n13148, n13149,
    n13150, n13151, n13152, n13153, n13154, n13155,
    n13156, n13157, n13158, n13159, n13160, n13161,
    n13162, n13163, n13164, n13165, n13166, n13167,
    n13168, n13169, n13170, n13171, n13172, n13173,
    n13174, n13175, n13176, n13177, n13178, n13179,
    n13180, n13181, n13182, n13183, n13184, n13185,
    n13186, n13187, n13188, n13189, n13190, n13191,
    n13192, n13193, n13194, n13195, n13196, n13197,
    n13198, n13199, n13200, n13201, n13202, n13203,
    n13204, n13205, n13206, n13207, n13208, n13209,
    n13210, n13211, n13212, n13213, n13214, n13215,
    n13216, n13217, n13218, n13219, n13220, n13221,
    n13222, n13223, n13224, n13225, n13226, n13227,
    n13228, n13229, n13230, n13231, n13232, n13233,
    n13234, n13235, n13236, n13237, n13238, n13239,
    n13240, n13241, n13242, n13243, n13244, n13245,
    n13246, n13247, n13248, n13249, n13250, n13251,
    n13252, n13253, n13254, n13255, n13256, n13257,
    n13258, n13259, n13260, n13261, n13262, n13263,
    n13264, n13265, n13266, n13267, n13268, n13269,
    n13270, n13271, n13272, n13273, n13274, n13275,
    n13276, n13277, n13278, n13279, n13280, n13281,
    n13282, n13283, n13284, n13286, n13287, n13288,
    n13289, n13290, n13291, n13292, n13293, n13294,
    n13295, n13296, n13297, n13298, n13299, n13300,
    n13301, n13302, n13303, n13304, n13305, n13306,
    n13307, n13308, n13309, n13310, n13311, n13312,
    n13313, n13314, n13315, n13316, n13317, n13318,
    n13319, n13320, n13321, n13322, n13323, n13324,
    n13325, n13326, n13327, n13328, n13329, n13330,
    n13331, n13332, n13333, n13334, n13335, n13336,
    n13337, n13338, n13339, n13340, n13341, n13342,
    n13343, n13344, n13345, n13346, n13347, n13348,
    n13349, n13350, n13351, n13352, n13353, n13354,
    n13355, n13356, n13357, n13358, n13359, n13360,
    n13361, n13362, n13363, n13364, n13365, n13366,
    n13367, n13368, n13369, n13370, n13371, n13372,
    n13373, n13374, n13375, n13376, n13377, n13378,
    n13379, n13380, n13381, n13382, n13383, n13384,
    n13385, n13386, n13387, n13388, n13389, n13390,
    n13391, n13392, n13393, n13394, n13395, n13396,
    n13397, n13398, n13399, n13400, n13401, n13402,
    n13403, n13404, n13405, n13406, n13407, n13408,
    n13409, n13410, n13411, n13412, n13413, n13414,
    n13415, n13416, n13417, n13418, n13419, n13420,
    n13421, n13422, n13423, n13424, n13425, n13426,
    n13427, n13428, n13429, n13430, n13431, n13432,
    n13433, n13434, n13435, n13436, n13437, n13438,
    n13439, n13440, n13441, n13442, n13443, n13444,
    n13445, n13446, n13447, n13448, n13449, n13450,
    n13451, n13452, n13453, n13454, n13455, n13456,
    n13457, n13458, n13459, n13460, n13461, n13462,
    n13463, n13464, n13465, n13466, n13467, n13468,
    n13469, n13470, n13471, n13472, n13473, n13474,
    n13475, n13476, n13477, n13478, n13479, n13480,
    n13481, n13482, n13483, n13484, n13485, n13486,
    n13487, n13488, n13489, n13490, n13491, n13492,
    n13493, n13494, n13495, n13496, n13497, n13498,
    n13499, n13500, n13501, n13502, n13503, n13504,
    n13505, n13506, n13507, n13508, n13509, n13510,
    n13511, n13512, n13513, n13514, n13515, n13516,
    n13517, n13518, n13519, n13520, n13521, n13522,
    n13523, n13524, n13525, n13526, n13527, n13528,
    n13529, n13530, n13531, n13532, n13533, n13534,
    n13535, n13536, n13537, n13538, n13539, n13540,
    n13541, n13542, n13543, n13544, n13545, n13546,
    n13547, n13548, n13549, n13550, n13551, n13552,
    n13553, n13554, n13555, n13556, n13557, n13558,
    n13559, n13560, n13561, n13562, n13563, n13564,
    n13565, n13566, n13567, n13568, n13569, n13570,
    n13571, n13572, n13573, n13574, n13575, n13576,
    n13577, n13578, n13579, n13580, n13581, n13582,
    n13583, n13584, n13585, n13586, n13587, n13588,
    n13589, n13590, n13591, n13592, n13593, n13594,
    n13595, n13596, n13597, n13598, n13599, n13600,
    n13601, n13602, n13603, n13604, n13605, n13606,
    n13607, n13608, n13609, n13610, n13611, n13612,
    n13613, n13614, n13615, n13616, n13617, n13618,
    n13619, n13620, n13621, n13622, n13623, n13624,
    n13625, n13626, n13627, n13628, n13629, n13630,
    n13631, n13632, n13633, n13634, n13635, n13636,
    n13637, n13638, n13639, n13640, n13641, n13642,
    n13643, n13644, n13645, n13646, n13647, n13648,
    n13649, n13650, n13651, n13652, n13653, n13654,
    n13655, n13656, n13657, n13658, n13659, n13660,
    n13661, n13662, n13663, n13664, n13665, n13666,
    n13667, n13668, n13669, n13670, n13671, n13672,
    n13673, n13674, n13675, n13676, n13677, n13678,
    n13679, n13680, n13681, n13682, n13683, n13684,
    n13685, n13686, n13687, n13688, n13689, n13690,
    n13691, n13692, n13693, n13694, n13695, n13696,
    n13697, n13698, n13699, n13700, n13701, n13702,
    n13703, n13704, n13705, n13706, n13707, n13708,
    n13709, n13710, n13711, n13712, n13713, n13714,
    n13715, n13716, n13717, n13718, n13719, n13720,
    n13721, n13722, n13723, n13724, n13725, n13726,
    n13727, n13728, n13729, n13730, n13731, n13732,
    n13733, n13734, n13735, n13736, n13737, n13738,
    n13739, n13740, n13741, n13742, n13743, n13744,
    n13745, n13746, n13747, n13748, n13749, n13750,
    n13751, n13752, n13753, n13754, n13755, n13756,
    n13757, n13758, n13759, n13760, n13761, n13762,
    n13763, n13764, n13765, n13766, n13767, n13768,
    n13769, n13770, n13771, n13772, n13773, n13774,
    n13775, n13776, n13777, n13778, n13779, n13780,
    n13781, n13782, n13783, n13784, n13785, n13786,
    n13787, n13789, n13790, n13791, n13792, n13793,
    n13794, n13795, n13796, n13797, n13798, n13799,
    n13800, n13801, n13802, n13803, n13804, n13805,
    n13806, n13807, n13808, n13809, n13810, n13811,
    n13812, n13813, n13814, n13815, n13816, n13817,
    n13818, n13819, n13820, n13821, n13822, n13823,
    n13824, n13825, n13826, n13827, n13828, n13829,
    n13830, n13831, n13832, n13833, n13834, n13835,
    n13836, n13837, n13838, n13839, n13840, n13841,
    n13842, n13843, n13844, n13845, n13846, n13847,
    n13848, n13849, n13850, n13851, n13852, n13853,
    n13854, n13855, n13856, n13857, n13858, n13859,
    n13860, n13861, n13862, n13863, n13864, n13865,
    n13866, n13867, n13868, n13869, n13870, n13871,
    n13872, n13873, n13874, n13875, n13876, n13877,
    n13878, n13879, n13880, n13881, n13882, n13883,
    n13884, n13885, n13886, n13887, n13888, n13889,
    n13890, n13891, n13892, n13893, n13894, n13895,
    n13896, n13897, n13898, n13899, n13900, n13901,
    n13902, n13903, n13904, n13905, n13906, n13907,
    n13908, n13909, n13910, n13911, n13912, n13913,
    n13914, n13915, n13916, n13917, n13918, n13919,
    n13920, n13921, n13922, n13923, n13924, n13925,
    n13926, n13927, n13928, n13929, n13930, n13931,
    n13932, n13933, n13934, n13935, n13936, n13937,
    n13938, n13939, n13940, n13941, n13942, n13943,
    n13944, n13945, n13946, n13947, n13948, n13949,
    n13950, n13951, n13952, n13953, n13954, n13955,
    n13956, n13957, n13958, n13959, n13960, n13961,
    n13962, n13963, n13964, n13965, n13966, n13967,
    n13968, n13969, n13970, n13971, n13972, n13973,
    n13974, n13975, n13976, n13977, n13978, n13979,
    n13980, n13981, n13982, n13983, n13984, n13985,
    n13986, n13987, n13988, n13989, n13990, n13991,
    n13992, n13993, n13994, n13995, n13996, n13997,
    n13998, n13999, n14000, n14001, n14002, n14003,
    n14004, n14005, n14006, n14007, n14008, n14009,
    n14010, n14011, n14012, n14013, n14014, n14015,
    n14016, n14017, n14018, n14019, n14020, n14021,
    n14022, n14023, n14024, n14025, n14026, n14027,
    n14028, n14029, n14030, n14031, n14032, n14033,
    n14034, n14035, n14036, n14037, n14038, n14039,
    n14040, n14041, n14042, n14043, n14044, n14045,
    n14046, n14047, n14048, n14049, n14050, n14051,
    n14052, n14053, n14054, n14055, n14056, n14057,
    n14058, n14059, n14060, n14061, n14062, n14063,
    n14064, n14065, n14066, n14067, n14068, n14069,
    n14070, n14071, n14072, n14073, n14074, n14075,
    n14076, n14077, n14078, n14079, n14080, n14081,
    n14082, n14083, n14084, n14085, n14086, n14087,
    n14088, n14089, n14090, n14091, n14092, n14093,
    n14094, n14095, n14096, n14097, n14098, n14099,
    n14100, n14101, n14102, n14103, n14104, n14105,
    n14106, n14107, n14108, n14109, n14110, n14111,
    n14112, n14113, n14114, n14115, n14116, n14117,
    n14118, n14119, n14120, n14121, n14122, n14123,
    n14124, n14125, n14126, n14127, n14128, n14129,
    n14130, n14131, n14132, n14133, n14134, n14135,
    n14136, n14137, n14138, n14139, n14140, n14141,
    n14142, n14143, n14144, n14145, n14146, n14147,
    n14148, n14149, n14150, n14151, n14152, n14153,
    n14154, n14155, n14156, n14157, n14158, n14159,
    n14160, n14161, n14162, n14163, n14164, n14165,
    n14166, n14167, n14168, n14169, n14170, n14171,
    n14172, n14173, n14174, n14175, n14176, n14177,
    n14178, n14179, n14180, n14181, n14182, n14183,
    n14184, n14185, n14186, n14187, n14188, n14189,
    n14190, n14191, n14192, n14193, n14194, n14195,
    n14196, n14197, n14198, n14199, n14200, n14201,
    n14202, n14203, n14204, n14205, n14206, n14207,
    n14208, n14209, n14210, n14211, n14212, n14213,
    n14214, n14215, n14216, n14217, n14218, n14219,
    n14220, n14221, n14222, n14223, n14224, n14225,
    n14226, n14227, n14228, n14229, n14230, n14231,
    n14232, n14233, n14234, n14235, n14236, n14237,
    n14238, n14239, n14240, n14241, n14242, n14243,
    n14244, n14245, n14246, n14247, n14248, n14249,
    n14250, n14251, n14252, n14253, n14254, n14255,
    n14256, n14257, n14258, n14259, n14260, n14261,
    n14262, n14263, n14264, n14265, n14266, n14267,
    n14268, n14269, n14270, n14271, n14272, n14273,
    n14274, n14275, n14276, n14277, n14278, n14279,
    n14280, n14281, n14282, n14283, n14284, n14285,
    n14286, n14287, n14288, n14289, n14290, n14291,
    n14292, n14293, n14294, n14295, n14296, n14297,
    n14298, n14299, n14300, n14302, n14303, n14304,
    n14305, n14306, n14307, n14308, n14309, n14310,
    n14311, n14312, n14313, n14314, n14315, n14316,
    n14317, n14318, n14319, n14320, n14321, n14322,
    n14323, n14324, n14325, n14326, n14327, n14328,
    n14329, n14330, n14331, n14332, n14333, n14334,
    n14335, n14336, n14337, n14338, n14339, n14340,
    n14341, n14342, n14343, n14344, n14345, n14346,
    n14347, n14348, n14349, n14350, n14351, n14352,
    n14353, n14354, n14355, n14356, n14357, n14358,
    n14359, n14360, n14361, n14362, n14363, n14364,
    n14365, n14366, n14367, n14368, n14369, n14370,
    n14371, n14372, n14373, n14374, n14375, n14376,
    n14377, n14378, n14379, n14380, n14381, n14382,
    n14383, n14384, n14385, n14386, n14387, n14388,
    n14389, n14390, n14391, n14392, n14393, n14394,
    n14395, n14396, n14397, n14398, n14399, n14400,
    n14401, n14402, n14403, n14404, n14405, n14406,
    n14407, n14408, n14409, n14410, n14411, n14412,
    n14413, n14414, n14415, n14416, n14417, n14418,
    n14419, n14420, n14421, n14422, n14423, n14424,
    n14425, n14426, n14427, n14428, n14429, n14430,
    n14431, n14432, n14433, n14434, n14435, n14436,
    n14437, n14438, n14439, n14440, n14441, n14442,
    n14443, n14444, n14445, n14446, n14447, n14448,
    n14449, n14450, n14451, n14452, n14453, n14454,
    n14455, n14456, n14457, n14458, n14459, n14460,
    n14461, n14462, n14463, n14464, n14465, n14466,
    n14467, n14468, n14469, n14470, n14471, n14472,
    n14473, n14474, n14475, n14476, n14477, n14478,
    n14479, n14480, n14481, n14482, n14483, n14484,
    n14485, n14486, n14487, n14488, n14489, n14490,
    n14491, n14492, n14493, n14494, n14495, n14496,
    n14497, n14498, n14499, n14500, n14501, n14502,
    n14503, n14504, n14505, n14506, n14507, n14508,
    n14509, n14510, n14511, n14512, n14513, n14514,
    n14515, n14516, n14517, n14518, n14519, n14520,
    n14521, n14522, n14523, n14524, n14525, n14526,
    n14527, n14528, n14529, n14530, n14531, n14532,
    n14533, n14534, n14535, n14536, n14537, n14538,
    n14539, n14540, n14541, n14542, n14543, n14544,
    n14545, n14546, n14547, n14548, n14549, n14550,
    n14551, n14552, n14553, n14554, n14555, n14556,
    n14557, n14558, n14559, n14560, n14561, n14562,
    n14563, n14564, n14565, n14566, n14567, n14568,
    n14569, n14570, n14571, n14572, n14573, n14574,
    n14575, n14576, n14577, n14578, n14579, n14580,
    n14581, n14582, n14583, n14584, n14585, n14586,
    n14587, n14588, n14589, n14590, n14591, n14592,
    n14593, n14594, n14595, n14596, n14597, n14598,
    n14599, n14600, n14601, n14602, n14603, n14604,
    n14605, n14606, n14607, n14608, n14609, n14610,
    n14611, n14612, n14613, n14614, n14615, n14616,
    n14617, n14618, n14619, n14620, n14621, n14622,
    n14623, n14624, n14625, n14626, n14627, n14628,
    n14629, n14630, n14631, n14632, n14633, n14634,
    n14635, n14636, n14637, n14638, n14639, n14640,
    n14641, n14642, n14643, n14644, n14645, n14646,
    n14647, n14648, n14649, n14650, n14651, n14652,
    n14653, n14654, n14655, n14656, n14657, n14658,
    n14659, n14660, n14661, n14662, n14663, n14664,
    n14665, n14666, n14667, n14668, n14669, n14670,
    n14671, n14672, n14673, n14674, n14675, n14676,
    n14677, n14678, n14679, n14680, n14681, n14682,
    n14683, n14684, n14685, n14686, n14687, n14688,
    n14689, n14690, n14691, n14692, n14693, n14694,
    n14695, n14696, n14697, n14698, n14699, n14700,
    n14701, n14702, n14703, n14704, n14705, n14706,
    n14707, n14708, n14709, n14710, n14711, n14712,
    n14713, n14714, n14715, n14716, n14717, n14718,
    n14719, n14720, n14721, n14722, n14723, n14724,
    n14725, n14726, n14727, n14728, n14729, n14730,
    n14731, n14732, n14733, n14734, n14735, n14736,
    n14737, n14738, n14739, n14740, n14741, n14742,
    n14743, n14744, n14745, n14746, n14747, n14748,
    n14749, n14750, n14751, n14752, n14753, n14754,
    n14755, n14756, n14757, n14758, n14759, n14760,
    n14761, n14762, n14763, n14764, n14765, n14766,
    n14767, n14768, n14769, n14770, n14771, n14772,
    n14773, n14774, n14775, n14776, n14777, n14778,
    n14779, n14780, n14781, n14782, n14783, n14784,
    n14785, n14786, n14787, n14788, n14789, n14790,
    n14791, n14792, n14793, n14794, n14795, n14796,
    n14797, n14798, n14799, n14800, n14801, n14802,
    n14803, n14804, n14805, n14806, n14807, n14808,
    n14809, n14810, n14811, n14812, n14813, n14814,
    n14815, n14816, n14817, n14818, n14819, n14820,
    n14821, n14822, n14823, n14824, n14826, n14827,
    n14828, n14829, n14830, n14831, n14832, n14833,
    n14834, n14835, n14836, n14837, n14838, n14839,
    n14840, n14841, n14842, n14843, n14844, n14845,
    n14846, n14847, n14848, n14849, n14850, n14851,
    n14852, n14853, n14854, n14855, n14856, n14857,
    n14858, n14859, n14860, n14861, n14862, n14863,
    n14864, n14865, n14866, n14867, n14868, n14869,
    n14870, n14871, n14872, n14873, n14874, n14875,
    n14876, n14877, n14878, n14879, n14880, n14881,
    n14882, n14883, n14884, n14885, n14886, n14887,
    n14888, n14889, n14890, n14891, n14892, n14893,
    n14894, n14895, n14896, n14897, n14898, n14899,
    n14900, n14901, n14902, n14903, n14904, n14905,
    n14906, n14907, n14908, n14909, n14910, n14911,
    n14912, n14913, n14914, n14915, n14916, n14917,
    n14918, n14919, n14920, n14921, n14922, n14923,
    n14924, n14925, n14926, n14927, n14928, n14929,
    n14930, n14931, n14932, n14933, n14934, n14935,
    n14936, n14937, n14938, n14939, n14940, n14941,
    n14942, n14943, n14944, n14945, n14946, n14947,
    n14948, n14949, n14950, n14951, n14952, n14953,
    n14954, n14955, n14956, n14957, n14958, n14959,
    n14960, n14961, n14962, n14963, n14964, n14965,
    n14966, n14967, n14968, n14969, n14970, n14971,
    n14972, n14973, n14974, n14975, n14976, n14977,
    n14978, n14979, n14980, n14981, n14982, n14983,
    n14984, n14985, n14986, n14987, n14988, n14989,
    n14990, n14991, n14992, n14993, n14994, n14995,
    n14996, n14997, n14998, n14999, n15000, n15001,
    n15002, n15003, n15004, n15005, n15006, n15007,
    n15008, n15009, n15010, n15011, n15012, n15013,
    n15014, n15015, n15016, n15017, n15018, n15019,
    n15020, n15021, n15022, n15023, n15024, n15025,
    n15026, n15027, n15028, n15029, n15030, n15031,
    n15032, n15033, n15034, n15035, n15036, n15037,
    n15038, n15039, n15040, n15041, n15042, n15043,
    n15044, n15045, n15046, n15047, n15048, n15049,
    n15050, n15051, n15052, n15053, n15054, n15055,
    n15056, n15057, n15058, n15059, n15060, n15061,
    n15062, n15063, n15064, n15065, n15066, n15067,
    n15068, n15069, n15070, n15071, n15072, n15073,
    n15074, n15075, n15076, n15077, n15078, n15079,
    n15080, n15081, n15082, n15083, n15084, n15085,
    n15086, n15087, n15088, n15089, n15090, n15091,
    n15092, n15093, n15094, n15095, n15096, n15097,
    n15098, n15099, n15100, n15101, n15102, n15103,
    n15104, n15105, n15106, n15107, n15108, n15109,
    n15110, n15111, n15112, n15113, n15114, n15115,
    n15116, n15117, n15118, n15119, n15120, n15121,
    n15122, n15123, n15124, n15125, n15126, n15127,
    n15128, n15129, n15130, n15131, n15132, n15133,
    n15134, n15135, n15136, n15137, n15138, n15139,
    n15140, n15141, n15142, n15143, n15144, n15145,
    n15146, n15147, n15148, n15149, n15150, n15151,
    n15152, n15153, n15154, n15155, n15156, n15157,
    n15158, n15159, n15160, n15161, n15162, n15163,
    n15164, n15165, n15166, n15167, n15168, n15169,
    n15170, n15171, n15172, n15173, n15174, n15175,
    n15176, n15177, n15178, n15179, n15180, n15181,
    n15182, n15183, n15184, n15185, n15186, n15187,
    n15188, n15189, n15190, n15191, n15192, n15193,
    n15194, n15195, n15196, n15197, n15198, n15199,
    n15200, n15201, n15202, n15203, n15204, n15205,
    n15206, n15207, n15208, n15209, n15210, n15211,
    n15212, n15213, n15214, n15215, n15216, n15217,
    n15218, n15219, n15220, n15221, n15222, n15223,
    n15224, n15225, n15226, n15227, n15228, n15229,
    n15230, n15231, n15232, n15233, n15234, n15235,
    n15236, n15237, n15238, n15239, n15240, n15241,
    n15242, n15243, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15252, n15253,
    n15254, n15255, n15256, n15257, n15258, n15259,
    n15260, n15261, n15262, n15263, n15264, n15265,
    n15266, n15267, n15268, n15269, n15270, n15271,
    n15272, n15273, n15274, n15275, n15276, n15277,
    n15278, n15279, n15280, n15281, n15282, n15283,
    n15284, n15285, n15286, n15287, n15288, n15289,
    n15290, n15291, n15292, n15293, n15294, n15295,
    n15296, n15297, n15298, n15299, n15300, n15301,
    n15302, n15303, n15304, n15305, n15306, n15307,
    n15308, n15309, n15310, n15311, n15312, n15313,
    n15314, n15315, n15316, n15317, n15318, n15319,
    n15320, n15321, n15322, n15323, n15324, n15325,
    n15326, n15327, n15328, n15329, n15330, n15331,
    n15332, n15333, n15334, n15335, n15336, n15337,
    n15338, n15339, n15340, n15341, n15342, n15343,
    n15344, n15345, n15346, n15347, n15348, n15349,
    n15350, n15351, n15352, n15353, n15354, n15355,
    n15356, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368,
    n15369, n15370, n15371, n15372, n15373, n15374,
    n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392,
    n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404,
    n15405, n15406, n15407, n15408, n15409, n15410,
    n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422,
    n15423, n15424, n15425, n15426, n15427, n15428,
    n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440,
    n15441, n15442, n15443, n15444, n15445, n15446,
    n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458,
    n15459, n15460, n15461, n15462, n15463, n15464,
    n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476,
    n15477, n15478, n15479, n15480, n15481, n15482,
    n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494,
    n15495, n15496, n15497, n15498, n15499, n15500,
    n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512,
    n15513, n15514, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530,
    n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15768, n15769, n15770,
    n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782,
    n15783, n15784, n15785, n15786, n15787, n15788,
    n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800,
    n15801, n15802, n15803, n15804, n15805, n15806,
    n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824,
    n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854,
    n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872,
    n15873, n15874, n15875, n15876, n15877, n15878,
    n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890,
    n15891, n15892, n15893, n15894, n15895, n15896,
    n15897, n15899, n15900, n15901, n15902, n15903,
    n15904, n15905, n15906, n15907, n15908, n15909,
    n15910, n15911, n15912, n15913, n15914, n15915,
    n15916, n15917, n15918, n15919, n15920, n15921,
    n15922, n15923, n15924, n15925, n15926, n15927,
    n15928, n15929, n15930, n15931, n15932, n15933,
    n15934, n15935, n15936, n15937, n15938, n15939,
    n15940, n15941, n15942, n15943, n15944, n15945,
    n15946, n15947, n15948, n15949, n15950, n15951,
    n15952, n15953, n15954, n15955, n15956, n15957,
    n15958, n15959, n15960, n15961, n15962, n15963,
    n15964, n15965, n15966, n15967, n15968, n15969,
    n15970, n15971, n15972, n15973, n15974, n15975,
    n15976, n15977, n15978, n15979, n15980, n15981,
    n15982, n15983, n15984, n15985, n15986, n15987,
    n15988, n15989, n15990, n15991, n15992, n15993,
    n15994, n15995, n15996, n15997, n15998, n15999,
    n16000, n16001, n16002, n16003, n16004, n16005,
    n16006, n16007, n16008, n16009, n16010, n16011,
    n16012, n16013, n16014, n16015, n16016, n16017,
    n16018, n16019, n16020, n16021, n16022, n16023,
    n16024, n16025, n16026, n16027, n16028, n16029,
    n16030, n16031, n16032, n16033, n16034, n16035,
    n16036, n16037, n16038, n16039, n16040, n16041,
    n16042, n16043, n16044, n16045, n16046, n16047,
    n16048, n16049, n16050, n16051, n16052, n16053,
    n16054, n16055, n16056, n16057, n16058, n16059,
    n16060, n16061, n16062, n16063, n16064, n16065,
    n16066, n16067, n16068, n16069, n16070, n16071,
    n16072, n16073, n16074, n16075, n16076, n16077,
    n16078, n16079, n16080, n16081, n16082, n16083,
    n16084, n16085, n16086, n16087, n16088, n16089,
    n16090, n16091, n16092, n16093, n16094, n16095,
    n16096, n16097, n16098, n16099, n16100, n16101,
    n16102, n16103, n16104, n16105, n16106, n16107,
    n16108, n16109, n16110, n16111, n16112, n16113,
    n16114, n16115, n16116, n16117, n16118, n16119,
    n16120, n16121, n16122, n16123, n16124, n16125,
    n16126, n16127, n16128, n16129, n16130, n16131,
    n16132, n16133, n16134, n16135, n16136, n16137,
    n16138, n16139, n16140, n16141, n16142, n16143,
    n16144, n16145, n16146, n16147, n16148, n16149,
    n16150, n16151, n16152, n16153, n16154, n16155,
    n16156, n16157, n16158, n16159, n16160, n16161,
    n16162, n16163, n16164, n16165, n16166, n16167,
    n16168, n16169, n16170, n16171, n16172, n16173,
    n16174, n16175, n16176, n16177, n16178, n16179,
    n16180, n16181, n16182, n16183, n16184, n16185,
    n16186, n16187, n16188, n16189, n16190, n16191,
    n16192, n16193, n16194, n16195, n16196, n16197,
    n16198, n16199, n16200, n16201, n16202, n16203,
    n16204, n16205, n16206, n16207, n16208, n16209,
    n16210, n16211, n16212, n16213, n16214, n16215,
    n16216, n16217, n16218, n16219, n16220, n16221,
    n16222, n16223, n16224, n16225, n16226, n16227,
    n16228, n16229, n16230, n16231, n16232, n16233,
    n16234, n16235, n16236, n16237, n16238, n16239,
    n16240, n16241, n16242, n16243, n16244, n16245,
    n16246, n16247, n16248, n16249, n16250, n16251,
    n16252, n16253, n16254, n16255, n16256, n16257,
    n16258, n16259, n16260, n16261, n16262, n16263,
    n16264, n16265, n16266, n16267, n16268, n16269,
    n16270, n16271, n16272, n16273, n16274, n16275,
    n16276, n16277, n16278, n16279, n16280, n16281,
    n16282, n16283, n16284, n16285, n16286, n16287,
    n16288, n16289, n16290, n16291, n16292, n16293,
    n16294, n16295, n16296, n16297, n16298, n16299,
    n16300, n16301, n16302, n16303, n16304, n16305,
    n16306, n16307, n16308, n16309, n16310, n16311,
    n16312, n16313, n16314, n16315, n16316, n16317,
    n16318, n16319, n16320, n16321, n16322, n16323,
    n16324, n16325, n16326, n16327, n16328, n16329,
    n16330, n16331, n16332, n16333, n16334, n16335,
    n16336, n16337, n16338, n16339, n16340, n16341,
    n16342, n16343, n16344, n16345, n16346, n16347,
    n16348, n16349, n16350, n16351, n16352, n16353,
    n16354, n16355, n16356, n16357, n16358, n16359,
    n16360, n16361, n16362, n16363, n16364, n16365,
    n16366, n16367, n16368, n16369, n16370, n16371,
    n16372, n16373, n16374, n16375, n16376, n16377,
    n16378, n16379, n16380, n16381, n16382, n16383,
    n16384, n16385, n16386, n16387, n16388, n16389,
    n16390, n16391, n16392, n16393, n16394, n16395,
    n16396, n16397, n16398, n16399, n16400, n16401,
    n16402, n16403, n16404, n16405, n16406, n16407,
    n16408, n16409, n16410, n16411, n16412, n16413,
    n16414, n16415, n16416, n16417, n16418, n16419,
    n16420, n16421, n16422, n16423, n16424, n16425,
    n16426, n16427, n16428, n16429, n16430, n16431,
    n16432, n16433, n16434, n16435, n16436, n16437,
    n16438, n16439, n16440, n16441, n16442, n16443,
    n16444, n16445, n16446, n16447, n16448, n16450,
    n16451, n16452, n16453, n16454, n16455, n16456,
    n16457, n16458, n16459, n16460, n16461, n16462,
    n16463, n16464, n16465, n16466, n16467, n16468,
    n16469, n16470, n16471, n16472, n16473, n16474,
    n16475, n16476, n16477, n16478, n16479, n16480,
    n16481, n16482, n16483, n16484, n16485, n16486,
    n16487, n16488, n16489, n16490, n16491, n16492,
    n16493, n16494, n16495, n16496, n16497, n16498,
    n16499, n16500, n16501, n16502, n16503, n16504,
    n16505, n16506, n16507, n16508, n16509, n16510,
    n16511, n16512, n16513, n16514, n16515, n16516,
    n16517, n16518, n16519, n16520, n16521, n16522,
    n16523, n16524, n16525, n16526, n16527, n16528,
    n16529, n16530, n16531, n16532, n16533, n16534,
    n16535, n16536, n16537, n16538, n16539, n16540,
    n16541, n16542, n16543, n16544, n16545, n16546,
    n16547, n16548, n16549, n16550, n16551, n16552,
    n16553, n16554, n16555, n16556, n16557, n16558,
    n16559, n16560, n16561, n16562, n16563, n16564,
    n16565, n16566, n16567, n16568, n16569, n16570,
    n16571, n16572, n16573, n16574, n16575, n16576,
    n16577, n16578, n16579, n16580, n16581, n16582,
    n16583, n16584, n16585, n16586, n16587, n16588,
    n16589, n16590, n16591, n16592, n16593, n16594,
    n16595, n16596, n16597, n16598, n16599, n16600,
    n16601, n16602, n16603, n16604, n16605, n16606,
    n16607, n16608, n16609, n16610, n16611, n16612,
    n16613, n16614, n16615, n16616, n16617, n16618,
    n16619, n16620, n16621, n16622, n16623, n16624,
    n16625, n16626, n16627, n16628, n16629, n16630,
    n16631, n16632, n16633, n16634, n16635, n16636,
    n16637, n16638, n16639, n16640, n16641, n16642,
    n16643, n16644, n16645, n16646, n16647, n16648,
    n16649, n16650, n16651, n16652, n16653, n16654,
    n16655, n16656, n16657, n16658, n16659, n16660,
    n16661, n16662, n16663, n16664, n16665, n16666,
    n16667, n16668, n16669, n16670, n16671, n16672,
    n16673, n16674, n16675, n16676, n16677, n16678,
    n16679, n16680, n16681, n16682, n16683, n16684,
    n16685, n16686, n16687, n16688, n16689, n16690,
    n16691, n16692, n16693, n16694, n16695, n16696,
    n16697, n16698, n16699, n16700, n16701, n16702,
    n16703, n16704, n16705, n16706, n16707, n16708,
    n16709, n16710, n16711, n16712, n16713, n16714,
    n16715, n16716, n16717, n16718, n16719, n16720,
    n16721, n16722, n16723, n16724, n16725, n16726,
    n16727, n16728, n16729, n16730, n16731, n16732,
    n16733, n16734, n16735, n16736, n16737, n16738,
    n16739, n16740, n16741, n16742, n16743, n16744,
    n16745, n16746, n16747, n16748, n16749, n16750,
    n16751, n16752, n16753, n16754, n16755, n16756,
    n16757, n16758, n16759, n16760, n16761, n16762,
    n16763, n16764, n16765, n16766, n16767, n16768,
    n16769, n16770, n16771, n16772, n16773, n16774,
    n16775, n16776, n16777, n16778, n16779, n16780,
    n16781, n16782, n16783, n16784, n16785, n16786,
    n16787, n16788, n16789, n16790, n16791, n16792,
    n16793, n16794, n16795, n16796, n16797, n16798,
    n16799, n16800, n16801, n16802, n16803, n16804,
    n16805, n16806, n16807, n16808, n16809, n16810,
    n16811, n16812, n16813, n16814, n16815, n16816,
    n16817, n16818, n16819, n16820, n16821, n16822,
    n16823, n16824, n16825, n16826, n16827, n16828,
    n16829, n16830, n16831, n16832, n16833, n16834,
    n16835, n16836, n16837, n16838, n16839, n16840,
    n16841, n16842, n16843, n16844, n16845, n16846,
    n16847, n16848, n16849, n16850, n16851, n16852,
    n16853, n16854, n16855, n16856, n16857, n16858,
    n16859, n16860, n16861, n16862, n16863, n16864,
    n16865, n16866, n16867, n16868, n16869, n16870,
    n16871, n16872, n16873, n16874, n16875, n16876,
    n16877, n16878, n16879, n16880, n16881, n16882,
    n16883, n16884, n16885, n16886, n16887, n16888,
    n16889, n16890, n16891, n16892, n16893, n16894,
    n16895, n16896, n16897, n16898, n16899, n16900,
    n16901, n16902, n16903, n16904, n16905, n16906,
    n16907, n16908, n16909, n16910, n16911, n16912,
    n16913, n16914, n16915, n16916, n16917, n16918,
    n16919, n16920, n16921, n16922, n16923, n16924,
    n16925, n16926, n16927, n16928, n16929, n16930,
    n16931, n16932, n16933, n16934, n16935, n16936,
    n16937, n16938, n16939, n16940, n16941, n16942,
    n16943, n16944, n16945, n16946, n16947, n16948,
    n16949, n16950, n16951, n16952, n16953, n16954,
    n16955, n16956, n16957, n16958, n16959, n16960,
    n16961, n16962, n16963, n16964, n16965, n16966,
    n16967, n16968, n16969, n16970, n16971, n16972,
    n16973, n16974, n16975, n16976, n16977, n16978,
    n16979, n16980, n16981, n16982, n16983, n16984,
    n16985, n16986, n16987, n16988, n16989, n16990,
    n16991, n16992, n16993, n16994, n16995, n16996,
    n16997, n16998, n16999, n17000, n17001, n17002,
    n17003, n17004, n17005, n17006, n17007, n17008,
    n17009, n17010, n17012, n17013, n17014, n17015,
    n17016, n17017, n17018, n17019, n17020, n17021,
    n17022, n17023, n17024, n17025, n17026, n17027,
    n17028, n17029, n17030, n17031, n17032, n17033,
    n17034, n17035, n17036, n17037, n17038, n17039,
    n17040, n17041, n17042, n17043, n17044, n17045,
    n17046, n17047, n17048, n17049, n17050, n17051,
    n17052, n17053, n17054, n17055, n17056, n17057,
    n17058, n17059, n17060, n17061, n17062, n17063,
    n17064, n17065, n17066, n17067, n17068, n17069,
    n17070, n17071, n17072, n17073, n17074, n17075,
    n17076, n17077, n17078, n17079, n17080, n17081,
    n17082, n17083, n17084, n17085, n17086, n17087,
    n17088, n17089, n17090, n17091, n17092, n17093,
    n17094, n17095, n17096, n17097, n17098, n17099,
    n17100, n17101, n17102, n17103, n17104, n17105,
    n17106, n17107, n17108, n17109, n17110, n17111,
    n17112, n17113, n17114, n17115, n17116, n17117,
    n17118, n17119, n17120, n17121, n17122, n17123,
    n17124, n17125, n17126, n17127, n17128, n17129,
    n17130, n17131, n17132, n17133, n17134, n17135,
    n17136, n17137, n17138, n17139, n17140, n17141,
    n17142, n17143, n17144, n17145, n17146, n17147,
    n17148, n17149, n17150, n17151, n17152, n17153,
    n17154, n17155, n17156, n17157, n17158, n17159,
    n17160, n17161, n17162, n17163, n17164, n17165,
    n17166, n17167, n17168, n17169, n17170, n17171,
    n17172, n17173, n17174, n17175, n17176, n17177,
    n17178, n17179, n17180, n17181, n17182, n17183,
    n17184, n17185, n17186, n17187, n17188, n17189,
    n17190, n17191, n17192, n17193, n17194, n17195,
    n17196, n17197, n17198, n17199, n17200, n17201,
    n17202, n17203, n17204, n17205, n17206, n17207,
    n17208, n17209, n17210, n17211, n17212, n17213,
    n17214, n17215, n17216, n17217, n17218, n17219,
    n17220, n17221, n17222, n17223, n17224, n17225,
    n17226, n17227, n17228, n17229, n17230, n17231,
    n17232, n17233, n17234, n17235, n17236, n17237,
    n17238, n17239, n17240, n17241, n17242, n17243,
    n17244, n17245, n17246, n17247, n17248, n17249,
    n17250, n17251, n17252, n17253, n17254, n17255,
    n17256, n17257, n17258, n17259, n17260, n17261,
    n17262, n17263, n17264, n17265, n17266, n17267,
    n17268, n17269, n17270, n17271, n17272, n17273,
    n17274, n17275, n17276, n17277, n17278, n17279,
    n17280, n17281, n17282, n17283, n17284, n17285,
    n17286, n17287, n17288, n17289, n17290, n17291,
    n17292, n17293, n17294, n17295, n17296, n17297,
    n17298, n17299, n17300, n17301, n17302, n17303,
    n17304, n17305, n17306, n17307, n17308, n17309,
    n17310, n17311, n17312, n17313, n17314, n17315,
    n17316, n17317, n17318, n17319, n17320, n17321,
    n17322, n17323, n17324, n17325, n17326, n17327,
    n17328, n17329, n17330, n17331, n17332, n17333,
    n17334, n17335, n17336, n17337, n17338, n17339,
    n17340, n17341, n17342, n17343, n17344, n17345,
    n17346, n17347, n17348, n17349, n17350, n17351,
    n17352, n17353, n17354, n17355, n17356, n17357,
    n17358, n17359, n17360, n17361, n17362, n17363,
    n17364, n17365, n17366, n17367, n17368, n17369,
    n17370, n17371, n17372, n17373, n17374, n17375,
    n17376, n17377, n17378, n17379, n17380, n17381,
    n17382, n17383, n17384, n17385, n17386, n17387,
    n17388, n17389, n17390, n17391, n17392, n17393,
    n17394, n17395, n17396, n17397, n17398, n17399,
    n17400, n17401, n17402, n17403, n17404, n17405,
    n17406, n17407, n17408, n17409, n17410, n17411,
    n17412, n17413, n17414, n17415, n17416, n17417,
    n17418, n17419, n17420, n17421, n17422, n17423,
    n17424, n17425, n17426, n17427, n17428, n17429,
    n17430, n17431, n17432, n17433, n17434, n17435,
    n17436, n17437, n17438, n17439, n17440, n17441,
    n17442, n17443, n17444, n17445, n17446, n17447,
    n17448, n17449, n17450, n17451, n17452, n17453,
    n17454, n17455, n17456, n17457, n17458, n17459,
    n17460, n17461, n17462, n17463, n17464, n17465,
    n17466, n17467, n17468, n17469, n17470, n17471,
    n17472, n17473, n17474, n17475, n17476, n17477,
    n17478, n17479, n17480, n17481, n17482, n17483,
    n17484, n17485, n17486, n17487, n17488, n17489,
    n17490, n17491, n17492, n17493, n17494, n17495,
    n17496, n17497, n17498, n17499, n17500, n17501,
    n17502, n17503, n17504, n17505, n17506, n17507,
    n17508, n17509, n17510, n17511, n17512, n17513,
    n17514, n17515, n17516, n17517, n17518, n17519,
    n17520, n17521, n17522, n17523, n17524, n17525,
    n17526, n17527, n17528, n17529, n17530, n17531,
    n17532, n17533, n17534, n17535, n17536, n17537,
    n17538, n17539, n17540, n17541, n17542, n17543,
    n17544, n17545, n17546, n17547, n17548, n17549,
    n17550, n17551, n17552, n17553, n17554, n17555,
    n17556, n17557, n17558, n17559, n17560, n17561,
    n17562, n17563, n17564, n17565, n17566, n17567,
    n17568, n17569, n17570, n17571, n17572, n17573,
    n17574, n17575, n17576, n17577, n17578, n17579,
    n17580, n17582, n17583, n17584, n17585, n17586,
    n17587, n17588, n17589, n17590, n17591, n17592,
    n17593, n17594, n17595, n17596, n17597, n17598,
    n17599, n17600, n17601, n17602, n17603, n17604,
    n17605, n17606, n17607, n17608, n17609, n17610,
    n17611, n17612, n17613, n17614, n17615, n17616,
    n17617, n17618, n17619, n17620, n17621, n17622,
    n17623, n17624, n17625, n17626, n17627, n17628,
    n17629, n17630, n17631, n17632, n17633, n17634,
    n17635, n17636, n17637, n17638, n17639, n17640,
    n17641, n17642, n17643, n17644, n17645, n17646,
    n17647, n17648, n17649, n17650, n17651, n17652,
    n17653, n17654, n17655, n17656, n17657, n17658,
    n17659, n17660, n17661, n17662, n17663, n17664,
    n17665, n17666, n17667, n17668, n17669, n17670,
    n17671, n17672, n17673, n17674, n17675, n17676,
    n17677, n17678, n17679, n17680, n17681, n17682,
    n17683, n17684, n17685, n17686, n17687, n17688,
    n17689, n17690, n17691, n17692, n17693, n17694,
    n17695, n17696, n17697, n17698, n17699, n17700,
    n17701, n17702, n17703, n17704, n17705, n17706,
    n17707, n17708, n17709, n17710, n17711, n17712,
    n17713, n17714, n17715, n17716, n17717, n17718,
    n17719, n17720, n17721, n17722, n17723, n17724,
    n17725, n17726, n17727, n17728, n17729, n17730,
    n17731, n17732, n17733, n17734, n17735, n17736,
    n17737, n17738, n17739, n17740, n17741, n17742,
    n17743, n17744, n17745, n17746, n17747, n17748,
    n17749, n17750, n17751, n17752, n17753, n17754,
    n17755, n17756, n17757, n17758, n17759, n17760,
    n17761, n17762, n17763, n17764, n17765, n17766,
    n17767, n17768, n17769, n17770, n17771, n17772,
    n17773, n17774, n17775, n17776, n17777, n17778,
    n17779, n17780, n17781, n17782, n17783, n17784,
    n17785, n17786, n17787, n17788, n17789, n17790,
    n17791, n17792, n17793, n17794, n17795, n17796,
    n17797, n17798, n17799, n17800, n17801, n17802,
    n17803, n17804, n17805, n17806, n17807, n17808,
    n17809, n17810, n17811, n17812, n17813, n17814,
    n17815, n17816, n17817, n17818, n17819, n17820,
    n17821, n17822, n17823, n17824, n17825, n17826,
    n17827, n17828, n17829, n17830, n17831, n17832,
    n17833, n17834, n17835, n17836, n17837, n17838,
    n17839, n17840, n17841, n17842, n17843, n17844,
    n17845, n17846, n17847, n17848, n17849, n17850,
    n17851, n17852, n17853, n17854, n17855, n17856,
    n17857, n17858, n17859, n17860, n17861, n17862,
    n17863, n17864, n17865, n17866, n17867, n17868,
    n17869, n17870, n17871, n17872, n17873, n17874,
    n17875, n17876, n17877, n17878, n17879, n17880,
    n17881, n17882, n17883, n17884, n17885, n17886,
    n17887, n17888, n17889, n17890, n17891, n17892,
    n17893, n17894, n17895, n17896, n17897, n17898,
    n17899, n17900, n17901, n17902, n17903, n17904,
    n17905, n17906, n17907, n17908, n17909, n17910,
    n17911, n17912, n17913, n17914, n17915, n17916,
    n17917, n17918, n17919, n17920, n17921, n17922,
    n17923, n17924, n17925, n17926, n17927, n17928,
    n17929, n17930, n17931, n17932, n17933, n17934,
    n17935, n17936, n17937, n17938, n17939, n17940,
    n17941, n17942, n17943, n17944, n17945, n17946,
    n17947, n17948, n17949, n17950, n17951, n17952,
    n17953, n17954, n17955, n17956, n17957, n17958,
    n17959, n17960, n17961, n17962, n17963, n17964,
    n17965, n17966, n17967, n17968, n17969, n17970,
    n17971, n17972, n17973, n17974, n17975, n17976,
    n17977, n17978, n17979, n17980, n17981, n17982,
    n17983, n17984, n17985, n17986, n17987, n17988,
    n17989, n17990, n17991, n17992, n17993, n17994,
    n17995, n17996, n17997, n17998, n17999, n18000,
    n18001, n18002, n18003, n18004, n18005, n18006,
    n18007, n18008, n18009, n18010, n18011, n18012,
    n18013, n18014, n18015, n18016, n18017, n18018,
    n18019, n18020, n18021, n18022, n18023, n18024,
    n18025, n18026, n18027, n18028, n18029, n18030,
    n18031, n18032, n18033, n18034, n18035, n18036,
    n18037, n18038, n18039, n18040, n18041, n18042,
    n18043, n18044, n18045, n18046, n18047, n18048,
    n18049, n18050, n18051, n18052, n18053, n18054,
    n18055, n18056, n18057, n18058, n18059, n18060,
    n18061, n18062, n18063, n18064, n18065, n18066,
    n18067, n18068, n18069, n18070, n18071, n18072,
    n18073, n18074, n18075, n18076, n18077, n18078,
    n18079, n18080, n18081, n18082, n18083, n18084,
    n18085, n18086, n18087, n18088, n18089, n18090,
    n18091, n18092, n18093, n18094, n18095, n18096,
    n18097, n18098, n18099, n18100, n18101, n18102,
    n18103, n18104, n18105, n18106, n18107, n18108,
    n18109, n18110, n18111, n18112, n18113, n18114,
    n18115, n18116, n18117, n18118, n18119, n18120,
    n18121, n18122, n18123, n18124, n18125, n18126,
    n18127, n18128, n18129, n18130, n18131, n18132,
    n18133, n18134, n18135, n18136, n18137, n18138,
    n18139, n18140, n18141, n18142, n18143, n18144,
    n18145, n18146, n18147, n18148, n18149, n18150,
    n18151, n18152, n18153, n18154, n18155, n18156,
    n18157, n18158, n18159, n18161, n18162, n18163,
    n18164, n18165, n18166, n18167, n18168, n18169,
    n18170, n18171, n18172, n18173, n18174, n18175,
    n18176, n18177, n18178, n18179, n18180, n18181,
    n18182, n18183, n18184, n18185, n18186, n18187,
    n18188, n18189, n18190, n18191, n18192, n18193,
    n18194, n18195, n18196, n18197, n18198, n18199,
    n18200, n18201, n18202, n18203, n18204, n18205,
    n18206, n18207, n18208, n18209, n18210, n18211,
    n18212, n18213, n18214, n18215, n18216, n18217,
    n18218, n18219, n18220, n18221, n18222, n18223,
    n18224, n18225, n18226, n18227, n18228, n18229,
    n18230, n18231, n18232, n18233, n18234, n18235,
    n18236, n18237, n18238, n18239, n18240, n18241,
    n18242, n18243, n18244, n18245, n18246, n18247,
    n18248, n18249, n18250, n18251, n18252, n18253,
    n18254, n18255, n18256, n18257, n18258, n18259,
    n18260, n18261, n18262, n18263, n18264, n18265,
    n18266, n18267, n18268, n18269, n18270, n18271,
    n18272, n18273, n18274, n18275, n18276, n18277,
    n18278, n18279, n18280, n18281, n18282, n18283,
    n18284, n18285, n18286, n18287, n18288, n18289,
    n18290, n18291, n18292, n18293, n18294, n18295,
    n18296, n18297, n18298, n18299, n18300, n18301,
    n18302, n18303, n18304, n18305, n18306, n18307,
    n18308, n18309, n18310, n18311, n18312, n18313,
    n18314, n18315, n18316, n18317, n18318, n18319,
    n18320, n18321, n18322, n18323, n18324, n18325,
    n18326, n18327, n18328, n18329, n18330, n18331,
    n18332, n18333, n18334, n18335, n18336, n18337,
    n18338, n18339, n18340, n18341, n18342, n18343,
    n18344, n18345, n18346, n18347, n18348, n18349,
    n18350, n18351, n18352, n18353, n18354, n18355,
    n18356, n18357, n18358, n18359, n18360, n18361,
    n18362, n18363, n18364, n18365, n18366, n18367,
    n18368, n18369, n18370, n18371, n18372, n18373,
    n18374, n18375, n18376, n18377, n18378, n18379,
    n18380, n18381, n18382, n18383, n18384, n18385,
    n18386, n18387, n18388, n18389, n18390, n18391,
    n18392, n18393, n18394, n18395, n18396, n18397,
    n18398, n18399, n18400, n18401, n18402, n18403,
    n18404, n18405, n18406, n18407, n18408, n18409,
    n18410, n18411, n18412, n18413, n18414, n18415,
    n18416, n18417, n18418, n18419, n18420, n18421,
    n18422, n18423, n18424, n18425, n18426, n18427,
    n18428, n18429, n18430, n18431, n18432, n18433,
    n18434, n18435, n18436, n18437, n18438, n18439,
    n18440, n18441, n18442, n18443, n18444, n18445,
    n18446, n18447, n18448, n18449, n18450, n18451,
    n18452, n18453, n18454, n18455, n18456, n18457,
    n18458, n18459, n18460, n18461, n18462, n18463,
    n18464, n18465, n18466, n18467, n18468, n18469,
    n18470, n18471, n18472, n18473, n18474, n18475,
    n18476, n18477, n18478, n18479, n18480, n18481,
    n18482, n18483, n18484, n18485, n18486, n18487,
    n18488, n18489, n18490, n18491, n18492, n18493,
    n18494, n18495, n18496, n18497, n18498, n18499,
    n18500, n18501, n18502, n18503, n18504, n18505,
    n18506, n18507, n18508, n18509, n18510, n18511,
    n18512, n18513, n18514, n18515, n18516, n18517,
    n18518, n18519, n18520, n18521, n18522, n18523,
    n18524, n18525, n18526, n18527, n18528, n18529,
    n18530, n18531, n18532, n18533, n18534, n18535,
    n18536, n18537, n18538, n18539, n18540, n18541,
    n18542, n18543, n18544, n18545, n18546, n18547,
    n18548, n18549, n18550, n18551, n18552, n18553,
    n18554, n18555, n18556, n18557, n18558, n18559,
    n18560, n18561, n18562, n18563, n18564, n18565,
    n18566, n18567, n18568, n18569, n18570, n18571,
    n18572, n18573, n18574, n18575, n18576, n18577,
    n18578, n18579, n18580, n18581, n18582, n18583,
    n18584, n18585, n18586, n18587, n18588, n18589,
    n18590, n18591, n18592, n18593, n18594, n18595,
    n18596, n18597, n18598, n18599, n18600, n18601,
    n18602, n18603, n18604, n18605, n18606, n18607,
    n18608, n18609, n18610, n18611, n18612, n18613,
    n18614, n18615, n18616, n18617, n18618, n18619,
    n18620, n18621, n18622, n18623, n18624, n18625,
    n18626, n18627, n18628, n18629, n18630, n18631,
    n18632, n18633, n18634, n18635, n18636, n18637,
    n18638, n18639, n18640, n18641, n18642, n18643,
    n18644, n18645, n18646, n18647, n18648, n18649,
    n18650, n18651, n18652, n18653, n18654, n18655,
    n18656, n18657, n18658, n18659, n18660, n18661,
    n18662, n18663, n18664, n18665, n18666, n18667,
    n18668, n18669, n18670, n18671, n18672, n18673,
    n18674, n18675, n18676, n18677, n18678, n18679,
    n18680, n18681, n18682, n18683, n18684, n18685,
    n18686, n18687, n18688, n18689, n18690, n18691,
    n18692, n18693, n18694, n18695, n18696, n18697,
    n18698, n18699, n18700, n18701, n18702, n18703,
    n18704, n18705, n18706, n18707, n18708, n18709,
    n18710, n18711, n18712, n18713, n18714, n18715,
    n18716, n18717, n18718, n18719, n18720, n18721,
    n18722, n18723, n18724, n18725, n18726, n18727,
    n18728, n18729, n18730, n18731, n18732, n18733,
    n18734, n18735, n18736, n18737, n18738, n18739,
    n18740, n18741, n18742, n18743, n18744, n18745,
    n18746, n18747, n18748, n18750, n18751, n18752,
    n18753, n18754, n18755, n18756, n18757, n18758,
    n18759, n18760, n18761, n18762, n18763, n18764,
    n18765, n18766, n18767, n18768, n18769, n18770,
    n18771, n18772, n18773, n18774, n18775, n18776,
    n18777, n18778, n18779, n18780, n18781, n18782,
    n18783, n18784, n18785, n18786, n18787, n18788,
    n18789, n18790, n18791, n18792, n18793, n18794,
    n18795, n18796, n18797, n18798, n18799, n18800,
    n18801, n18802, n18803, n18804, n18805, n18806,
    n18807, n18808, n18809, n18810, n18811, n18812,
    n18813, n18814, n18815, n18816, n18817, n18818,
    n18819, n18820, n18821, n18822, n18823, n18824,
    n18825, n18826, n18827, n18828, n18829, n18830,
    n18831, n18832, n18833, n18834, n18835, n18836,
    n18837, n18838, n18839, n18840, n18841, n18842,
    n18843, n18844, n18845, n18846, n18847, n18848,
    n18849, n18850, n18851, n18852, n18853, n18854,
    n18855, n18856, n18857, n18858, n18859, n18860,
    n18861, n18862, n18863, n18864, n18865, n18866,
    n18867, n18868, n18869, n18870, n18871, n18872,
    n18873, n18874, n18875, n18876, n18877, n18878,
    n18879, n18880, n18881, n18882, n18883, n18884,
    n18885, n18886, n18887, n18888, n18889, n18890,
    n18891, n18892, n18893, n18894, n18895, n18896,
    n18897, n18898, n18899, n18900, n18901, n18902,
    n18903, n18904, n18905, n18906, n18907, n18908,
    n18909, n18910, n18911, n18912, n18913, n18914,
    n18915, n18916, n18917, n18918, n18919, n18920,
    n18921, n18922, n18923, n18924, n18925, n18926,
    n18927, n18928, n18929, n18930, n18931, n18932,
    n18933, n18934, n18935, n18936, n18937, n18938,
    n18939, n18940, n18941, n18942, n18943, n18944,
    n18945, n18946, n18947, n18948, n18949, n18950,
    n18951, n18952, n18953, n18954, n18955, n18956,
    n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968,
    n18969, n18970, n18971, n18972, n18973, n18974,
    n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986,
    n18987, n18988, n18989, n18990, n18991, n18992,
    n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004,
    n19005, n19006, n19007, n19008, n19009, n19010,
    n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022,
    n19023, n19024, n19025, n19026, n19027, n19028,
    n19029, n19030, n19031, n19032, n19033, n19034,
    n19035, n19036, n19037, n19038, n19039, n19040,
    n19041, n19042, n19043, n19044, n19045, n19046,
    n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058,
    n19059, n19060, n19061, n19062, n19063, n19064,
    n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076,
    n19077, n19078, n19079, n19080, n19081, n19082,
    n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094,
    n19095, n19096, n19097, n19098, n19099, n19100,
    n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112,
    n19113, n19114, n19115, n19116, n19117, n19118,
    n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130,
    n19131, n19132, n19133, n19134, n19135, n19136,
    n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148,
    n19149, n19150, n19151, n19152, n19153, n19154,
    n19155, n19156, n19157, n19158, n19159, n19160,
    n19161, n19162, n19163, n19164, n19165, n19166,
    n19167, n19168, n19169, n19170, n19171, n19172,
    n19173, n19174, n19175, n19176, n19177, n19178,
    n19179, n19180, n19181, n19182, n19183, n19184,
    n19185, n19186, n19187, n19188, n19189, n19190,
    n19191, n19192, n19193, n19194, n19195, n19196,
    n19197, n19198, n19199, n19200, n19201, n19202,
    n19203, n19204, n19205, n19206, n19207, n19208,
    n19209, n19210, n19211, n19212, n19213, n19214,
    n19215, n19216, n19217, n19218, n19219, n19220,
    n19221, n19222, n19223, n19224, n19225, n19226,
    n19227, n19228, n19229, n19230, n19231, n19232,
    n19233, n19234, n19235, n19236, n19237, n19238,
    n19239, n19240, n19241, n19242, n19243, n19244,
    n19245, n19246, n19247, n19248, n19249, n19250,
    n19251, n19252, n19253, n19254, n19255, n19256,
    n19257, n19258, n19259, n19260, n19261, n19262,
    n19263, n19264, n19265, n19266, n19267, n19268,
    n19269, n19270, n19271, n19272, n19273, n19274,
    n19275, n19276, n19277, n19278, n19279, n19280,
    n19281, n19282, n19283, n19284, n19285, n19286,
    n19287, n19288, n19289, n19290, n19291, n19292,
    n19293, n19294, n19295, n19296, n19297, n19298,
    n19299, n19300, n19301, n19302, n19303, n19304,
    n19305, n19306, n19307, n19308, n19309, n19310,
    n19311, n19312, n19313, n19314, n19315, n19316;
  assign po63  = pi126  | pi127 ;
  assign n194 = pi126  & pi127 ;
  assign n195 = ~pi124  & ~pi125 ;
  assign n196 = ~pi126  & ~n195;
  assign po62  = n194 | n196;
  assign n198 = ~pi124  & po62 ;
  assign n199 = pi125  & ~n198;
  assign n200 = n194 & n195;
  assign n201 = ~n199 & ~n200;
  assign n202 = pi124  & po62 ;
  assign n203 = ~pi122  & ~pi123 ;
  assign n204 = ~pi124  & n203;
  assign n205 = ~n202 & ~n204;
  assign n206 = n201 & ~n205;
  assign n207 = ~po63  & ~n206;
  assign n208 = ~n201 & n205;
  assign n209 = pi126  & n195;
  assign n210 = pi127  & ~n196;
  assign n211 = ~n209 & n210;
  assign n212 = ~n208 & ~n211;
  assign po61  = n207 | ~n212;
  assign n214 = ~pi122  & po61 ;
  assign n215 = ~pi123  & n214;
  assign n216 = po62  & ~po61 ;
  assign n217 = ~n215 & ~n216;
  assign n218 = pi124  & ~n217;
  assign n219 = ~pi124  & n217;
  assign n220 = ~n218 & ~n219;
  assign n221 = pi122  & po61 ;
  assign n222 = ~pi120  & ~pi121 ;
  assign n223 = ~pi122  & n222;
  assign n224 = ~n221 & ~n223;
  assign n225 = ~po62  & n224;
  assign n226 = pi123  & ~n214;
  assign n227 = ~n215 & ~n226;
  assign n228 = po62  & ~n224;
  assign n229 = ~n227 & ~n228;
  assign n230 = ~n225 & ~n229;
  assign n231 = ~n220 & n230;
  assign n232 = ~po63  & ~n231;
  assign n233 = n220 & ~n230;
  assign n234 = n205 & ~po61 ;
  assign n235 = po63  & ~n206;
  assign n236 = ~n208 & n235;
  assign n237 = ~n234 & n236;
  assign n238 = ~n233 & ~n237;
  assign po60  = n232 | ~n238;
  assign n240 = ~n225 & po60 ;
  assign n241 = ~n228 & n240;
  assign n242 = n227 & ~n241;
  assign n243 = n229 & n240;
  assign n244 = ~n242 & ~n243;
  assign n245 = po63  & ~n231;
  assign n246 = ~n233 & n245;
  assign n247 = ~n238 & ~n246;
  assign n248 = pi120  & po60 ;
  assign n249 = ~pi118  & ~pi119 ;
  assign n250 = ~pi120  & n249;
  assign n251 = ~n248 & ~n250;
  assign n252 = po61  & ~n251;
  assign n253 = ~pi120  & po60 ;
  assign n254 = pi121  & ~n253;
  assign n255 = ~pi121  & n253;
  assign n256 = ~n254 & ~n255;
  assign n257 = ~po61  & n251;
  assign n258 = n256 & ~n257;
  assign n259 = ~n252 & ~n258;
  assign n260 = ~po62  & n259;
  assign n261 = po62  & ~n259;
  assign n262 = po61  & ~po60 ;
  assign n263 = ~n255 & ~n262;
  assign n264 = pi122  & ~n263;
  assign n265 = ~pi122  & n263;
  assign n266 = ~n264 & ~n265;
  assign n267 = ~n261 & n266;
  assign n268 = ~n260 & ~n267;
  assign n269 = ~n244 & ~n247;
  assign n270 = n268 & n269;
  assign n271 = ~po63  & ~n270;
  assign n272 = n244 & ~n268;
  assign n273 = ~n220 & ~po60 ;
  assign n274 = n246 & ~n273;
  assign n275 = ~n272 & ~n274;
  assign po59  = n271 | ~n275;
  assign n277 = pi118  & po59 ;
  assign n278 = ~pi116  & ~pi117 ;
  assign n279 = ~pi118  & n278;
  assign n280 = ~n277 & ~n279;
  assign n281 = ~po60  & n280;
  assign n282 = po60  & ~n280;
  assign n283 = ~pi118  & po59 ;
  assign n284 = pi119  & ~n283;
  assign n285 = ~pi119  & n283;
  assign n286 = ~n284 & ~n285;
  assign n287 = ~n282 & ~n286;
  assign n288 = ~n281 & ~n287;
  assign n289 = po61  & n288;
  assign n290 = po60  & ~po59 ;
  assign n291 = ~n285 & ~n290;
  assign n292 = pi120  & ~n291;
  assign n293 = ~pi120  & n291;
  assign n294 = ~n292 & ~n293;
  assign n295 = ~po61  & ~n288;
  assign n296 = ~n294 & ~n295;
  assign n297 = ~n289 & ~n296;
  assign n298 = po62  & ~n297;
  assign n299 = ~po62  & ~n289;
  assign n300 = ~n296 & n299;
  assign n301 = ~n252 & ~n257;
  assign n302 = po59  & n301;
  assign n303 = n256 & ~n302;
  assign n304 = ~n256 & n302;
  assign n305 = ~n303 & ~n304;
  assign n306 = ~n300 & ~n305;
  assign n307 = ~n298 & ~n306;
  assign n308 = ~n268 & po59 ;
  assign n309 = ~n244 & ~n308;
  assign n310 = po59  & n309;
  assign n311 = ~n260 & ~n261;
  assign n312 = po59  & n311;
  assign n313 = ~n266 & ~n312;
  assign n314 = n266 & n312;
  assign n315 = ~n313 & ~n314;
  assign n316 = ~n272 & ~n310;
  assign n317 = ~n315 & n316;
  assign n318 = ~n307 & n317;
  assign n319 = ~po63  & ~n318;
  assign n320 = n307 & n315;
  assign n321 = po63  & ~n272;
  assign n322 = ~n309 & n321;
  assign n323 = ~n320 & ~n322;
  assign po58  = n319 | ~n323;
  assign n325 = pi116  & po58 ;
  assign n326 = ~pi114  & ~pi115 ;
  assign n327 = ~pi116  & n326;
  assign n328 = ~n325 & ~n327;
  assign n329 = po59  & ~n328;
  assign n330 = ~pi116  & po58 ;
  assign n331 = pi117  & ~n330;
  assign n332 = ~pi117  & n330;
  assign n333 = ~n331 & ~n332;
  assign n334 = ~po59  & n328;
  assign n335 = n333 & ~n334;
  assign n336 = ~n329 & ~n335;
  assign n337 = po60  & ~n336;
  assign n338 = ~po60  & ~n329;
  assign n339 = ~n335 & n338;
  assign n340 = po59  & ~po58 ;
  assign n341 = ~n332 & ~n340;
  assign n342 = pi118  & ~n341;
  assign n343 = ~pi118  & n341;
  assign n344 = ~n342 & ~n343;
  assign n345 = ~n339 & ~n344;
  assign n346 = ~n337 & ~n345;
  assign n347 = po61  & ~n346;
  assign n348 = ~po61  & n346;
  assign n349 = ~n281 & ~n282;
  assign n350 = po58  & n349;
  assign n351 = n286 & ~n350;
  assign n352 = ~n286 & n350;
  assign n353 = ~n351 & ~n352;
  assign n354 = ~n348 & ~n353;
  assign n355 = ~n347 & ~n354;
  assign n356 = po62  & ~n355;
  assign n357 = ~po62  & ~n347;
  assign n358 = ~n354 & n357;
  assign n359 = ~n289 & po58 ;
  assign n360 = ~n295 & n359;
  assign n361 = n294 & ~n360;
  assign n362 = n296 & n359;
  assign n363 = ~n361 & ~n362;
  assign n364 = ~n358 & n363;
  assign n365 = ~n356 & ~n364;
  assign n366 = ~n315 & po58 ;
  assign n367 = ~n307 & n366;
  assign n368 = ~n298 & ~n300;
  assign n369 = po58  & n368;
  assign n370 = n305 & ~n369;
  assign n371 = ~n305 & n369;
  assign n372 = ~n370 & ~n371;
  assign n373 = ~n320 & ~n367;
  assign n374 = n372 & n373;
  assign n375 = ~n365 & n374;
  assign n376 = ~po63  & ~n375;
  assign n377 = n365 & ~n372;
  assign n378 = ~n307 & ~n315;
  assign n379 = n307 & ~n366;
  assign n380 = po63  & ~n378;
  assign n381 = ~n379 & n380;
  assign n382 = ~n377 & ~n381;
  assign po57  = n376 | ~n382;
  assign n384 = n244 & ~po59 ;
  assign n385 = pi114  & po57 ;
  assign n386 = ~pi112  & ~pi113 ;
  assign n387 = ~pi114  & n386;
  assign n388 = ~n385 & ~n387;
  assign n389 = ~po58  & ~n384;
  assign n390 = n388 & n389;
  assign n391 = po58  & ~n388;
  assign n392 = ~pi114  & po57 ;
  assign n393 = pi115  & ~n392;
  assign n394 = ~pi115  & n392;
  assign n395 = ~n393 & ~n394;
  assign n396 = ~n391 & ~n395;
  assign n397 = ~n390 & ~n396;
  assign n398 = po59  & n397;
  assign n399 = po58  & ~po57 ;
  assign n400 = ~n394 & ~n399;
  assign n401 = pi116  & ~n400;
  assign n402 = ~pi116  & n400;
  assign n403 = ~n401 & ~n402;
  assign n404 = ~po59  & ~n397;
  assign n405 = ~n403 & ~n404;
  assign n406 = ~n398 & ~n405;
  assign n407 = po60  & ~n406;
  assign n408 = ~po60  & ~n398;
  assign n409 = ~n405 & n408;
  assign n410 = ~n329 & ~n334;
  assign n411 = po57  & n410;
  assign n412 = n333 & ~n411;
  assign n413 = ~n333 & n411;
  assign n414 = ~n412 & ~n413;
  assign n415 = ~n409 & ~n414;
  assign n416 = ~n407 & ~n415;
  assign n417 = po61  & ~n416;
  assign n418 = ~n337 & ~n339;
  assign n419 = po57  & n418;
  assign n420 = ~n344 & ~n419;
  assign n421 = n344 & n419;
  assign n422 = ~n420 & ~n421;
  assign n423 = ~po61  & n416;
  assign n424 = ~n422 & ~n423;
  assign n425 = ~n417 & ~n424;
  assign n426 = po62  & ~n425;
  assign n427 = ~po62  & ~n417;
  assign n428 = ~n424 & n427;
  assign n429 = ~n347 & ~n348;
  assign n430 = po57  & n429;
  assign n431 = n353 & ~n430;
  assign n432 = ~n353 & n430;
  assign n433 = ~n431 & ~n432;
  assign n434 = ~n428 & n433;
  assign n435 = ~n426 & ~n434;
  assign n436 = n372 & po57 ;
  assign n437 = ~n365 & n436;
  assign n438 = ~n356 & ~n358;
  assign n439 = po57  & n438;
  assign n440 = n363 & ~n439;
  assign n441 = ~n363 & n439;
  assign n442 = ~n440 & ~n441;
  assign n443 = ~n377 & ~n437;
  assign n444 = ~n442 & n443;
  assign n445 = ~n435 & n444;
  assign n446 = ~po63  & ~n445;
  assign n447 = n435 & n442;
  assign n448 = n365 & ~n436;
  assign n449 = ~n365 & n372;
  assign n450 = po63  & ~n449;
  assign n451 = ~n448 & n450;
  assign n452 = ~n447 & ~n451;
  assign po56  = n446 | ~n452;
  assign n454 = pi112  & po56 ;
  assign n455 = ~pi110  & ~pi111 ;
  assign n456 = ~pi112  & n455;
  assign n457 = ~n454 & ~n456;
  assign n458 = po57  & ~n457;
  assign n459 = ~pi112  & po56 ;
  assign n460 = pi113  & ~n459;
  assign n461 = ~pi113  & n459;
  assign n462 = ~n460 & ~n461;
  assign n463 = ~po57  & n457;
  assign n464 = n462 & ~n463;
  assign n465 = ~n458 & ~n464;
  assign n466 = po58  & ~n465;
  assign n467 = ~po58  & ~n458;
  assign n468 = ~n464 & n467;
  assign n469 = po57  & ~po56 ;
  assign n470 = ~n461 & ~n469;
  assign n471 = pi114  & ~n470;
  assign n472 = ~pi114  & n470;
  assign n473 = ~n471 & ~n472;
  assign n474 = ~n468 & ~n473;
  assign n475 = ~n466 & ~n474;
  assign n476 = po59  & ~n475;
  assign n477 = ~po59  & n475;
  assign n478 = ~n390 & ~n391;
  assign n479 = po56  & n478;
  assign n480 = n395 & ~n479;
  assign n481 = ~n395 & n479;
  assign n482 = ~n480 & ~n481;
  assign n483 = ~n477 & ~n482;
  assign n484 = ~n476 & ~n483;
  assign n485 = po60  & ~n484;
  assign n486 = ~po60  & ~n476;
  assign n487 = ~n483 & n486;
  assign n488 = ~n398 & po56 ;
  assign n489 = ~n404 & n488;
  assign n490 = n403 & ~n489;
  assign n491 = n405 & n488;
  assign n492 = ~n490 & ~n491;
  assign n493 = ~n487 & n492;
  assign n494 = ~n485 & ~n493;
  assign n495 = po61  & ~n494;
  assign n496 = ~po61  & n494;
  assign n497 = ~n407 & ~n409;
  assign n498 = po56  & n497;
  assign n499 = n414 & ~n498;
  assign n500 = ~n414 & n498;
  assign n501 = ~n499 & ~n500;
  assign n502 = ~n496 & n501;
  assign n503 = ~n495 & ~n502;
  assign n504 = po62  & ~n503;
  assign n505 = ~po62  & ~n495;
  assign n506 = ~n502 & n505;
  assign n507 = ~n417 & po56 ;
  assign n508 = ~n423 & n507;
  assign n509 = n422 & ~n508;
  assign n510 = n424 & n507;
  assign n511 = ~n509 & ~n510;
  assign n512 = ~n506 & n511;
  assign n513 = ~n504 & ~n512;
  assign n514 = n435 & po56 ;
  assign n515 = ~n442 & ~n514;
  assign n516 = ~n447 & ~n515;
  assign n517 = po56  & ~n516;
  assign n518 = ~n426 & ~n428;
  assign n519 = po56  & n518;
  assign n520 = n433 & n519;
  assign n521 = ~n433 & ~n519;
  assign n522 = ~n520 & ~n521;
  assign n523 = ~n517 & n522;
  assign n524 = ~n513 & n523;
  assign n525 = ~po63  & ~n524;
  assign n526 = n513 & ~n522;
  assign n527 = po63  & n516;
  assign n528 = ~n526 & ~n527;
  assign po55  = n525 | ~n528;
  assign n530 = pi110  & po55 ;
  assign n531 = ~pi108  & ~pi109 ;
  assign n532 = ~pi110  & n531;
  assign n533 = ~n530 & ~n532;
  assign n534 = po56  & ~n533;
  assign n535 = ~po56  & n533;
  assign n536 = ~pi110  & po55 ;
  assign n537 = pi111  & ~n536;
  assign n538 = ~pi111  & n536;
  assign n539 = ~n537 & ~n538;
  assign n540 = ~n535 & n539;
  assign n541 = ~n534 & ~n540;
  assign n542 = po57  & ~n541;
  assign n543 = po56  & ~po55 ;
  assign n544 = ~n538 & ~n543;
  assign n545 = pi112  & ~n544;
  assign n546 = ~pi112  & n544;
  assign n547 = ~n545 & ~n546;
  assign n548 = ~po57  & n541;
  assign n549 = ~n547 & ~n548;
  assign n550 = ~n542 & ~n549;
  assign n551 = po58  & ~n550;
  assign n552 = ~po58  & ~n542;
  assign n553 = ~n549 & n552;
  assign n554 = ~n458 & ~n463;
  assign n555 = po55  & n554;
  assign n556 = n462 & ~n555;
  assign n557 = ~n462 & n555;
  assign n558 = ~n556 & ~n557;
  assign n559 = ~n553 & ~n558;
  assign n560 = ~n551 & ~n559;
  assign n561 = po59  & ~n560;
  assign n562 = ~n466 & ~n468;
  assign n563 = po55  & n562;
  assign n564 = ~n473 & ~n563;
  assign n565 = n473 & n563;
  assign n566 = ~n564 & ~n565;
  assign n567 = ~po59  & n560;
  assign n568 = ~n566 & ~n567;
  assign n569 = ~n561 & ~n568;
  assign n570 = po60  & ~n569;
  assign n571 = ~po60  & ~n561;
  assign n572 = ~n568 & n571;
  assign n573 = ~n476 & ~n477;
  assign n574 = po55  & n573;
  assign n575 = n482 & ~n574;
  assign n576 = ~n482 & n574;
  assign n577 = ~n575 & ~n576;
  assign n578 = ~n572 & n577;
  assign n579 = ~n570 & ~n578;
  assign n580 = po61  & ~n579;
  assign n581 = ~n485 & ~n487;
  assign n582 = po55  & n581;
  assign n583 = n492 & ~n582;
  assign n584 = ~n492 & n582;
  assign n585 = ~n583 & ~n584;
  assign n586 = ~po61  & n579;
  assign n587 = ~n585 & ~n586;
  assign n588 = ~n580 & ~n587;
  assign n589 = po62  & ~n588;
  assign n590 = ~po62  & ~n580;
  assign n591 = ~n587 & n590;
  assign n592 = ~n495 & ~n496;
  assign n593 = po55  & n592;
  assign n594 = n501 & n593;
  assign n595 = ~n501 & ~n593;
  assign n596 = ~n594 & ~n595;
  assign n597 = ~n591 & n596;
  assign n598 = ~n589 & ~n597;
  assign n599 = ~n504 & ~n506;
  assign n600 = po55  & n599;
  assign n601 = n511 & ~n600;
  assign n602 = ~n511 & n600;
  assign n603 = ~n601 & ~n602;
  assign n604 = n513 & po55 ;
  assign n605 = n522 & ~n604;
  assign n606 = ~n526 & ~n605;
  assign n607 = po55  & ~n606;
  assign n608 = ~n603 & ~n607;
  assign n609 = ~n598 & n608;
  assign n610 = ~po63  & ~n609;
  assign n611 = n598 & n603;
  assign n612 = po63  & n606;
  assign n613 = ~n611 & ~n612;
  assign po54  = n610 | ~n613;
  assign n615 = pi108  & po54 ;
  assign n616 = ~pi106  & ~pi107 ;
  assign n617 = ~pi108  & n616;
  assign n618 = ~n615 & ~n617;
  assign n619 = po55  & ~n618;
  assign n620 = ~pi108  & po54 ;
  assign n621 = pi109  & ~n620;
  assign n622 = ~pi109  & n620;
  assign n623 = ~n621 & ~n622;
  assign n624 = ~po55  & n618;
  assign n625 = n623 & ~n624;
  assign n626 = ~n619 & ~n625;
  assign n627 = po56  & ~n626;
  assign n628 = ~po56  & ~n619;
  assign n629 = ~n625 & n628;
  assign n630 = po55  & ~po54 ;
  assign n631 = ~n622 & ~n630;
  assign n632 = pi110  & ~n631;
  assign n633 = ~pi110  & n631;
  assign n634 = ~n632 & ~n633;
  assign n635 = ~n629 & ~n634;
  assign n636 = ~n627 & ~n635;
  assign n637 = po57  & ~n636;
  assign n638 = ~po57  & n636;
  assign n639 = ~n534 & ~n535;
  assign n640 = po54  & n639;
  assign n641 = n539 & ~n640;
  assign n642 = ~n539 & n640;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~n638 & ~n643;
  assign n645 = ~n637 & ~n644;
  assign n646 = po58  & ~n645;
  assign n647 = ~po58  & ~n637;
  assign n648 = ~n644 & n647;
  assign n649 = ~n542 & po54 ;
  assign n650 = ~n548 & n649;
  assign n651 = n547 & ~n650;
  assign n652 = n549 & n649;
  assign n653 = ~n651 & ~n652;
  assign n654 = ~n648 & n653;
  assign n655 = ~n646 & ~n654;
  assign n656 = po59  & ~n655;
  assign n657 = ~po59  & n655;
  assign n658 = ~n551 & ~n553;
  assign n659 = po54  & n658;
  assign n660 = n558 & ~n659;
  assign n661 = ~n558 & n659;
  assign n662 = ~n660 & ~n661;
  assign n663 = ~n657 & n662;
  assign n664 = ~n656 & ~n663;
  assign n665 = po60  & ~n664;
  assign n666 = ~po60  & ~n656;
  assign n667 = ~n663 & n666;
  assign n668 = ~n561 & po54 ;
  assign n669 = ~n567 & n668;
  assign n670 = n566 & ~n669;
  assign n671 = n568 & n668;
  assign n672 = ~n670 & ~n671;
  assign n673 = ~n667 & n672;
  assign n674 = ~n665 & ~n673;
  assign n675 = po61  & ~n674;
  assign n676 = ~po61  & n674;
  assign n677 = ~n570 & ~n572;
  assign n678 = po54  & n677;
  assign n679 = n577 & n678;
  assign n680 = ~n577 & ~n678;
  assign n681 = ~n679 & ~n680;
  assign n682 = ~n676 & n681;
  assign n683 = ~n675 & ~n682;
  assign n684 = po62  & ~n683;
  assign n685 = ~po62  & ~n675;
  assign n686 = ~n682 & n685;
  assign n687 = ~n580 & po54 ;
  assign n688 = ~n586 & n687;
  assign n689 = n585 & ~n688;
  assign n690 = n587 & n687;
  assign n691 = ~n689 & ~n690;
  assign n692 = ~n686 & n691;
  assign n693 = ~n684 & ~n692;
  assign n694 = ~n589 & ~n591;
  assign n695 = po54  & n694;
  assign n696 = ~n596 & ~n695;
  assign n697 = n596 & n695;
  assign n698 = ~n696 & ~n697;
  assign n699 = n598 & po54 ;
  assign n700 = ~n603 & ~n699;
  assign n701 = ~n611 & ~n700;
  assign n702 = po54  & ~n701;
  assign n703 = n698 & ~n702;
  assign n704 = ~n693 & n703;
  assign n705 = ~po63  & ~n704;
  assign n706 = n693 & ~n698;
  assign n707 = po63  & n701;
  assign n708 = ~n706 & ~n707;
  assign po53  = n705 | ~n708;
  assign n710 = pi106  & po53 ;
  assign n711 = ~pi104  & ~pi105 ;
  assign n712 = ~pi106  & n711;
  assign n713 = ~n710 & ~n712;
  assign n714 = po54  & ~n713;
  assign n715 = ~po54  & n713;
  assign n716 = ~pi106  & po53 ;
  assign n717 = pi107  & ~n716;
  assign n718 = ~pi107  & n716;
  assign n719 = ~n717 & ~n718;
  assign n720 = ~n715 & n719;
  assign n721 = ~n714 & ~n720;
  assign n722 = po55  & ~n721;
  assign n723 = po54  & ~po53 ;
  assign n724 = ~n718 & ~n723;
  assign n725 = pi108  & ~n724;
  assign n726 = ~pi108  & n724;
  assign n727 = ~n725 & ~n726;
  assign n728 = ~po55  & n721;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~n722 & ~n729;
  assign n731 = po56  & ~n730;
  assign n732 = ~po56  & ~n722;
  assign n733 = ~n729 & n732;
  assign n734 = ~n619 & ~n624;
  assign n735 = po53  & n734;
  assign n736 = n623 & ~n735;
  assign n737 = ~n623 & n735;
  assign n738 = ~n736 & ~n737;
  assign n739 = ~n733 & ~n738;
  assign n740 = ~n731 & ~n739;
  assign n741 = po57  & ~n740;
  assign n742 = ~n627 & ~n629;
  assign n743 = po53  & n742;
  assign n744 = ~n634 & ~n743;
  assign n745 = n634 & n743;
  assign n746 = ~n744 & ~n745;
  assign n747 = ~po57  & n740;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~n741 & ~n748;
  assign n750 = po58  & ~n749;
  assign n751 = ~po58  & ~n741;
  assign n752 = ~n748 & n751;
  assign n753 = ~n637 & ~n638;
  assign n754 = po53  & n753;
  assign n755 = n643 & ~n754;
  assign n756 = ~n643 & n754;
  assign n757 = ~n755 & ~n756;
  assign n758 = ~n752 & n757;
  assign n759 = ~n750 & ~n758;
  assign n760 = po59  & ~n759;
  assign n761 = ~n646 & ~n648;
  assign n762 = po53  & n761;
  assign n763 = n653 & ~n762;
  assign n764 = ~n653 & n762;
  assign n765 = ~n763 & ~n764;
  assign n766 = ~po59  & n759;
  assign n767 = ~n765 & ~n766;
  assign n768 = ~n760 & ~n767;
  assign n769 = po60  & ~n768;
  assign n770 = ~po60  & ~n760;
  assign n771 = ~n767 & n770;
  assign n772 = ~n656 & ~n657;
  assign n773 = po53  & n772;
  assign n774 = n662 & n773;
  assign n775 = ~n662 & ~n773;
  assign n776 = ~n774 & ~n775;
  assign n777 = ~n771 & n776;
  assign n778 = ~n769 & ~n777;
  assign n779 = po61  & ~n778;
  assign n780 = ~n665 & ~n667;
  assign n781 = po53  & n780;
  assign n782 = n672 & ~n781;
  assign n783 = ~n672 & n781;
  assign n784 = ~n782 & ~n783;
  assign n785 = ~po61  & n778;
  assign n786 = ~n784 & ~n785;
  assign n787 = ~n779 & ~n786;
  assign n788 = po62  & ~n787;
  assign n789 = ~po62  & ~n779;
  assign n790 = ~n786 & n789;
  assign n791 = ~n675 & ~n676;
  assign n792 = po53  & n791;
  assign n793 = ~n681 & ~n792;
  assign n794 = n681 & n792;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~n790 & n795;
  assign n797 = ~n788 & ~n796;
  assign n798 = n698 & po53 ;
  assign n799 = ~n693 & n798;
  assign n800 = ~n684 & ~n686;
  assign n801 = po53  & n800;
  assign n802 = n691 & ~n801;
  assign n803 = ~n691 & n801;
  assign n804 = ~n802 & ~n803;
  assign n805 = ~n706 & ~n799;
  assign n806 = ~n804 & n805;
  assign n807 = ~n797 & n806;
  assign n808 = ~po63  & ~n807;
  assign n809 = n797 & n804;
  assign n810 = n693 & ~n798;
  assign n811 = ~n693 & n698;
  assign n812 = po63  & ~n811;
  assign n813 = ~n810 & n812;
  assign n814 = ~n809 & ~n813;
  assign po52  = n808 | ~n814;
  assign n816 = pi104  & po52 ;
  assign n817 = ~pi102  & ~pi103 ;
  assign n818 = ~pi104  & n817;
  assign n819 = ~n816 & ~n818;
  assign n820 = po53  & ~n819;
  assign n821 = ~pi104  & po52 ;
  assign n822 = pi105  & ~n821;
  assign n823 = ~pi105  & n821;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~po53  & n819;
  assign n826 = n824 & ~n825;
  assign n827 = ~n820 & ~n826;
  assign n828 = po54  & ~n827;
  assign n829 = ~po54  & ~n820;
  assign n830 = ~n826 & n829;
  assign n831 = po53  & ~po52 ;
  assign n832 = ~n823 & ~n831;
  assign n833 = pi106  & ~n832;
  assign n834 = ~pi106  & n832;
  assign n835 = ~n833 & ~n834;
  assign n836 = ~n830 & ~n835;
  assign n837 = ~n828 & ~n836;
  assign n838 = po55  & ~n837;
  assign n839 = ~po55  & n837;
  assign n840 = ~n714 & ~n715;
  assign n841 = po52  & n840;
  assign n842 = n719 & ~n841;
  assign n843 = ~n719 & n841;
  assign n844 = ~n842 & ~n843;
  assign n845 = ~n839 & ~n844;
  assign n846 = ~n838 & ~n845;
  assign n847 = po56  & ~n846;
  assign n848 = ~po56  & ~n838;
  assign n849 = ~n845 & n848;
  assign n850 = ~n722 & po52 ;
  assign n851 = ~n728 & n850;
  assign n852 = n727 & ~n851;
  assign n853 = n729 & n850;
  assign n854 = ~n852 & ~n853;
  assign n855 = ~n849 & n854;
  assign n856 = ~n847 & ~n855;
  assign n857 = po57  & ~n856;
  assign n858 = ~po57  & n856;
  assign n859 = ~n731 & ~n733;
  assign n860 = po52  & n859;
  assign n861 = n738 & ~n860;
  assign n862 = ~n738 & n860;
  assign n863 = ~n861 & ~n862;
  assign n864 = ~n858 & n863;
  assign n865 = ~n857 & ~n864;
  assign n866 = po58  & ~n865;
  assign n867 = ~po58  & ~n857;
  assign n868 = ~n864 & n867;
  assign n869 = ~n741 & po52 ;
  assign n870 = ~n747 & n869;
  assign n871 = n746 & ~n870;
  assign n872 = n748 & n869;
  assign n873 = ~n871 & ~n872;
  assign n874 = ~n868 & n873;
  assign n875 = ~n866 & ~n874;
  assign n876 = po59  & ~n875;
  assign n877 = ~po59  & n875;
  assign n878 = ~n750 & ~n752;
  assign n879 = po52  & n878;
  assign n880 = n757 & n879;
  assign n881 = ~n757 & ~n879;
  assign n882 = ~n880 & ~n881;
  assign n883 = ~n877 & n882;
  assign n884 = ~n876 & ~n883;
  assign n885 = po60  & ~n884;
  assign n886 = ~po60  & ~n876;
  assign n887 = ~n883 & n886;
  assign n888 = ~n760 & po52 ;
  assign n889 = ~n766 & n888;
  assign n890 = n765 & ~n889;
  assign n891 = n767 & n888;
  assign n892 = ~n890 & ~n891;
  assign n893 = ~n887 & n892;
  assign n894 = ~n885 & ~n893;
  assign n895 = po61  & ~n894;
  assign n896 = ~po61  & n894;
  assign n897 = ~n769 & ~n771;
  assign n898 = po52  & n897;
  assign n899 = n776 & n898;
  assign n900 = ~n776 & ~n898;
  assign n901 = ~n899 & ~n900;
  assign n902 = ~n896 & n901;
  assign n903 = ~n895 & ~n902;
  assign n904 = po62  & ~n903;
  assign n905 = ~po62  & ~n895;
  assign n906 = ~n902 & n905;
  assign n907 = ~n779 & po52 ;
  assign n908 = ~n785 & n907;
  assign n909 = n784 & ~n908;
  assign n910 = n786 & n907;
  assign n911 = ~n909 & ~n910;
  assign n912 = ~n906 & n911;
  assign n913 = ~n904 & ~n912;
  assign n914 = ~n788 & ~n790;
  assign n915 = po52  & n914;
  assign n916 = n795 & ~n915;
  assign n917 = ~n795 & n915;
  assign n918 = ~n916 & ~n917;
  assign n919 = n797 & po52 ;
  assign n920 = ~n804 & ~n919;
  assign n921 = ~n809 & ~n920;
  assign n922 = po52  & ~n921;
  assign n923 = ~n918 & ~n922;
  assign n924 = ~n913 & n923;
  assign n925 = ~po63  & ~n924;
  assign n926 = n913 & n918;
  assign n927 = po63  & n921;
  assign n928 = ~n926 & ~n927;
  assign po51  = n925 | ~n928;
  assign n930 = pi102  & po51 ;
  assign n931 = ~pi100  & ~pi101 ;
  assign n932 = ~pi102  & n931;
  assign n933 = ~n930 & ~n932;
  assign n934 = po52  & ~n933;
  assign n935 = ~po52  & n933;
  assign n936 = ~pi102  & po51 ;
  assign n937 = pi103  & ~n936;
  assign n938 = ~pi103  & n936;
  assign n939 = ~n937 & ~n938;
  assign n940 = ~n935 & n939;
  assign n941 = ~n934 & ~n940;
  assign n942 = po53  & ~n941;
  assign n943 = po52  & ~po51 ;
  assign n944 = ~n938 & ~n943;
  assign n945 = pi104  & ~n944;
  assign n946 = ~pi104  & n944;
  assign n947 = ~n945 & ~n946;
  assign n948 = ~po53  & n941;
  assign n949 = ~n947 & ~n948;
  assign n950 = ~n942 & ~n949;
  assign n951 = po54  & ~n950;
  assign n952 = ~po54  & ~n942;
  assign n953 = ~n949 & n952;
  assign n954 = ~n820 & ~n825;
  assign n955 = po51  & n954;
  assign n956 = n824 & ~n955;
  assign n957 = ~n824 & n955;
  assign n958 = ~n956 & ~n957;
  assign n959 = ~n953 & ~n958;
  assign n960 = ~n951 & ~n959;
  assign n961 = po55  & ~n960;
  assign n962 = ~n828 & ~n830;
  assign n963 = po51  & n962;
  assign n964 = ~n835 & ~n963;
  assign n965 = n835 & n963;
  assign n966 = ~n964 & ~n965;
  assign n967 = ~po55  & n960;
  assign n968 = ~n966 & ~n967;
  assign n969 = ~n961 & ~n968;
  assign n970 = po56  & ~n969;
  assign n971 = ~po56  & ~n961;
  assign n972 = ~n968 & n971;
  assign n973 = ~n838 & ~n839;
  assign n974 = po51  & n973;
  assign n975 = n844 & ~n974;
  assign n976 = ~n844 & n974;
  assign n977 = ~n975 & ~n976;
  assign n978 = ~n972 & n977;
  assign n979 = ~n970 & ~n978;
  assign n980 = po57  & ~n979;
  assign n981 = ~n847 & ~n849;
  assign n982 = po51  & n981;
  assign n983 = n854 & ~n982;
  assign n984 = ~n854 & n982;
  assign n985 = ~n983 & ~n984;
  assign n986 = ~po57  & n979;
  assign n987 = ~n985 & ~n986;
  assign n988 = ~n980 & ~n987;
  assign n989 = po58  & ~n988;
  assign n990 = ~po58  & ~n980;
  assign n991 = ~n987 & n990;
  assign n992 = ~n857 & ~n858;
  assign n993 = po51  & n992;
  assign n994 = n863 & n993;
  assign n995 = ~n863 & ~n993;
  assign n996 = ~n994 & ~n995;
  assign n997 = ~n991 & n996;
  assign n998 = ~n989 & ~n997;
  assign n999 = po59  & ~n998;
  assign n1000 = ~n866 & ~n868;
  assign n1001 = po51  & n1000;
  assign n1002 = n873 & ~n1001;
  assign n1003 = ~n873 & n1001;
  assign n1004 = ~n1002 & ~n1003;
  assign n1005 = ~po59  & n998;
  assign n1006 = ~n1004 & ~n1005;
  assign n1007 = ~n999 & ~n1006;
  assign n1008 = po60  & ~n1007;
  assign n1009 = ~po60  & ~n999;
  assign n1010 = ~n1006 & n1009;
  assign n1011 = ~n876 & ~n877;
  assign n1012 = po51  & n1011;
  assign n1013 = ~n882 & ~n1012;
  assign n1014 = n882 & n1012;
  assign n1015 = ~n1013 & ~n1014;
  assign n1016 = ~n1010 & n1015;
  assign n1017 = ~n1008 & ~n1016;
  assign n1018 = po61  & ~n1017;
  assign n1019 = ~n885 & ~n887;
  assign n1020 = po51  & n1019;
  assign n1021 = n892 & ~n1020;
  assign n1022 = ~n892 & n1020;
  assign n1023 = ~n1021 & ~n1022;
  assign n1024 = ~po61  & n1017;
  assign n1025 = ~n1023 & ~n1024;
  assign n1026 = ~n1018 & ~n1025;
  assign n1027 = po62  & ~n1026;
  assign n1028 = ~po62  & ~n1018;
  assign n1029 = ~n1025 & n1028;
  assign n1030 = ~n895 & ~n896;
  assign n1031 = po51  & n1030;
  assign n1032 = ~n901 & ~n1031;
  assign n1033 = n901 & n1031;
  assign n1034 = ~n1032 & ~n1033;
  assign n1035 = ~n1029 & n1034;
  assign n1036 = ~n1027 & ~n1035;
  assign n1037 = ~n904 & ~n906;
  assign n1038 = po51  & n1037;
  assign n1039 = n911 & ~n1038;
  assign n1040 = ~n911 & n1038;
  assign n1041 = ~n1039 & ~n1040;
  assign n1042 = n913 & po51 ;
  assign n1043 = ~n918 & ~n1042;
  assign n1044 = ~n926 & ~n1043;
  assign n1045 = po51  & ~n1044;
  assign n1046 = ~n1041 & ~n1045;
  assign n1047 = ~n1036 & n1046;
  assign n1048 = ~po63  & ~n1047;
  assign n1049 = n1036 & n1041;
  assign n1050 = po63  & n1044;
  assign n1051 = ~n1049 & ~n1050;
  assign po50  = n1048 | ~n1051;
  assign n1053 = pi100  & po50 ;
  assign n1054 = ~pi98  & ~pi99 ;
  assign n1055 = ~pi100  & n1054;
  assign n1056 = ~n1053 & ~n1055;
  assign n1057 = po51  & ~n1056;
  assign n1058 = ~pi100  & po50 ;
  assign n1059 = pi101  & ~n1058;
  assign n1060 = ~pi101  & n1058;
  assign n1061 = ~n1059 & ~n1060;
  assign n1062 = ~po51  & n1056;
  assign n1063 = n1061 & ~n1062;
  assign n1064 = ~n1057 & ~n1063;
  assign n1065 = po52  & ~n1064;
  assign n1066 = ~po52  & ~n1057;
  assign n1067 = ~n1063 & n1066;
  assign n1068 = po51  & ~po50 ;
  assign n1069 = ~n1060 & ~n1068;
  assign n1070 = pi102  & ~n1069;
  assign n1071 = ~pi102  & n1069;
  assign n1072 = ~n1070 & ~n1071;
  assign n1073 = ~n1067 & ~n1072;
  assign n1074 = ~n1065 & ~n1073;
  assign n1075 = po53  & ~n1074;
  assign n1076 = ~po53  & n1074;
  assign n1077 = ~n934 & ~n935;
  assign n1078 = po50  & n1077;
  assign n1079 = n939 & ~n1078;
  assign n1080 = ~n939 & n1078;
  assign n1081 = ~n1079 & ~n1080;
  assign n1082 = ~n1076 & ~n1081;
  assign n1083 = ~n1075 & ~n1082;
  assign n1084 = po54  & ~n1083;
  assign n1085 = ~po54  & ~n1075;
  assign n1086 = ~n1082 & n1085;
  assign n1087 = ~n942 & po50 ;
  assign n1088 = ~n948 & n1087;
  assign n1089 = n947 & ~n1088;
  assign n1090 = n949 & n1087;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = ~n1086 & n1091;
  assign n1093 = ~n1084 & ~n1092;
  assign n1094 = po55  & ~n1093;
  assign n1095 = ~po55  & n1093;
  assign n1096 = ~n951 & ~n953;
  assign n1097 = po50  & n1096;
  assign n1098 = n958 & ~n1097;
  assign n1099 = ~n958 & n1097;
  assign n1100 = ~n1098 & ~n1099;
  assign n1101 = ~n1095 & n1100;
  assign n1102 = ~n1094 & ~n1101;
  assign n1103 = po56  & ~n1102;
  assign n1104 = ~po56  & ~n1094;
  assign n1105 = ~n1101 & n1104;
  assign n1106 = ~n961 & po50 ;
  assign n1107 = ~n967 & n1106;
  assign n1108 = n966 & ~n1107;
  assign n1109 = n968 & n1106;
  assign n1110 = ~n1108 & ~n1109;
  assign n1111 = ~n1105 & n1110;
  assign n1112 = ~n1103 & ~n1111;
  assign n1113 = po57  & ~n1112;
  assign n1114 = ~po57  & n1112;
  assign n1115 = ~n970 & ~n972;
  assign n1116 = po50  & n1115;
  assign n1117 = n977 & n1116;
  assign n1118 = ~n977 & ~n1116;
  assign n1119 = ~n1117 & ~n1118;
  assign n1120 = ~n1114 & n1119;
  assign n1121 = ~n1113 & ~n1120;
  assign n1122 = po58  & ~n1121;
  assign n1123 = ~po58  & ~n1113;
  assign n1124 = ~n1120 & n1123;
  assign n1125 = ~n980 & po50 ;
  assign n1126 = ~n986 & n1125;
  assign n1127 = n985 & ~n1126;
  assign n1128 = n987 & n1125;
  assign n1129 = ~n1127 & ~n1128;
  assign n1130 = ~n1124 & n1129;
  assign n1131 = ~n1122 & ~n1130;
  assign n1132 = po59  & ~n1131;
  assign n1133 = ~po59  & n1131;
  assign n1134 = ~n989 & ~n991;
  assign n1135 = po50  & n1134;
  assign n1136 = ~n996 & ~n1135;
  assign n1137 = n996 & n1135;
  assign n1138 = ~n1136 & ~n1137;
  assign n1139 = ~n1133 & n1138;
  assign n1140 = ~n1132 & ~n1139;
  assign n1141 = po60  & ~n1140;
  assign n1142 = ~po60  & ~n1132;
  assign n1143 = ~n1139 & n1142;
  assign n1144 = ~n999 & po50 ;
  assign n1145 = ~n1005 & n1144;
  assign n1146 = n1004 & ~n1145;
  assign n1147 = n1006 & n1144;
  assign n1148 = ~n1146 & ~n1147;
  assign n1149 = ~n1143 & n1148;
  assign n1150 = ~n1141 & ~n1149;
  assign n1151 = po61  & ~n1150;
  assign n1152 = ~n1008 & ~n1010;
  assign n1153 = po50  & n1152;
  assign n1154 = n1015 & ~n1153;
  assign n1155 = ~n1015 & n1153;
  assign n1156 = ~n1154 & ~n1155;
  assign n1157 = ~po61  & n1150;
  assign n1158 = ~n1156 & ~n1157;
  assign n1159 = ~n1151 & ~n1158;
  assign n1160 = po62  & ~n1159;
  assign n1161 = ~po62  & ~n1151;
  assign n1162 = ~n1158 & n1161;
  assign n1163 = ~n1018 & po50 ;
  assign n1164 = ~n1024 & n1163;
  assign n1165 = n1023 & ~n1164;
  assign n1166 = n1025 & n1163;
  assign n1167 = ~n1165 & ~n1166;
  assign n1168 = ~n1162 & n1167;
  assign n1169 = ~n1160 & ~n1168;
  assign n1170 = ~n1027 & ~n1029;
  assign n1171 = po50  & n1170;
  assign n1172 = n1034 & ~n1171;
  assign n1173 = ~n1034 & n1171;
  assign n1174 = ~n1172 & ~n1173;
  assign n1175 = n1036 & po50 ;
  assign n1176 = ~n1041 & ~n1175;
  assign n1177 = ~n1049 & ~n1176;
  assign n1178 = po50  & ~n1177;
  assign n1179 = ~n1174 & ~n1178;
  assign n1180 = ~n1169 & n1179;
  assign n1181 = ~po63  & ~n1180;
  assign n1182 = n1169 & n1174;
  assign n1183 = po63  & n1177;
  assign n1184 = ~n1182 & ~n1183;
  assign po49  = n1181 | ~n1184;
  assign n1186 = pi98  & po49 ;
  assign n1187 = ~pi96  & ~pi97 ;
  assign n1188 = ~pi98  & n1187;
  assign n1189 = ~n1186 & ~n1188;
  assign n1190 = po50  & ~n1189;
  assign n1191 = ~po50  & n1189;
  assign n1192 = ~pi98  & po49 ;
  assign n1193 = pi99  & ~n1192;
  assign n1194 = ~pi99  & n1192;
  assign n1195 = ~n1193 & ~n1194;
  assign n1196 = ~n1191 & n1195;
  assign n1197 = ~n1190 & ~n1196;
  assign n1198 = po51  & ~n1197;
  assign n1199 = po50  & ~po49 ;
  assign n1200 = ~n1194 & ~n1199;
  assign n1201 = pi100  & ~n1200;
  assign n1202 = ~pi100  & n1200;
  assign n1203 = ~n1201 & ~n1202;
  assign n1204 = ~po51  & n1197;
  assign n1205 = ~n1203 & ~n1204;
  assign n1206 = ~n1198 & ~n1205;
  assign n1207 = po52  & ~n1206;
  assign n1208 = ~po52  & ~n1198;
  assign n1209 = ~n1205 & n1208;
  assign n1210 = ~n1057 & ~n1062;
  assign n1211 = po49  & n1210;
  assign n1212 = n1061 & ~n1211;
  assign n1213 = ~n1061 & n1211;
  assign n1214 = ~n1212 & ~n1213;
  assign n1215 = ~n1209 & ~n1214;
  assign n1216 = ~n1207 & ~n1215;
  assign n1217 = po53  & ~n1216;
  assign n1218 = ~n1065 & ~n1067;
  assign n1219 = po49  & n1218;
  assign n1220 = ~n1072 & ~n1219;
  assign n1221 = n1072 & n1219;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = ~po53  & n1216;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = ~n1217 & ~n1224;
  assign n1226 = po54  & ~n1225;
  assign n1227 = ~po54  & ~n1217;
  assign n1228 = ~n1224 & n1227;
  assign n1229 = ~n1075 & ~n1076;
  assign n1230 = po49  & n1229;
  assign n1231 = n1081 & ~n1230;
  assign n1232 = ~n1081 & n1230;
  assign n1233 = ~n1231 & ~n1232;
  assign n1234 = ~n1228 & n1233;
  assign n1235 = ~n1226 & ~n1234;
  assign n1236 = po55  & ~n1235;
  assign n1237 = ~n1084 & ~n1086;
  assign n1238 = po49  & n1237;
  assign n1239 = n1091 & ~n1238;
  assign n1240 = ~n1091 & n1238;
  assign n1241 = ~n1239 & ~n1240;
  assign n1242 = ~po55  & n1235;
  assign n1243 = ~n1241 & ~n1242;
  assign n1244 = ~n1236 & ~n1243;
  assign n1245 = po56  & ~n1244;
  assign n1246 = ~po56  & ~n1236;
  assign n1247 = ~n1243 & n1246;
  assign n1248 = ~n1094 & ~n1095;
  assign n1249 = po49  & n1248;
  assign n1250 = n1100 & n1249;
  assign n1251 = ~n1100 & ~n1249;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = ~n1247 & n1252;
  assign n1254 = ~n1245 & ~n1253;
  assign n1255 = po57  & ~n1254;
  assign n1256 = ~n1103 & ~n1105;
  assign n1257 = po49  & n1256;
  assign n1258 = n1110 & ~n1257;
  assign n1259 = ~n1110 & n1257;
  assign n1260 = ~n1258 & ~n1259;
  assign n1261 = ~po57  & n1254;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = ~n1255 & ~n1262;
  assign n1264 = po58  & ~n1263;
  assign n1265 = ~po58  & ~n1255;
  assign n1266 = ~n1262 & n1265;
  assign n1267 = ~n1113 & ~n1114;
  assign n1268 = po49  & n1267;
  assign n1269 = ~n1119 & ~n1268;
  assign n1270 = n1119 & n1268;
  assign n1271 = ~n1269 & ~n1270;
  assign n1272 = ~n1266 & n1271;
  assign n1273 = ~n1264 & ~n1272;
  assign n1274 = po59  & ~n1273;
  assign n1275 = ~n1122 & ~n1124;
  assign n1276 = po49  & n1275;
  assign n1277 = n1129 & ~n1276;
  assign n1278 = ~n1129 & n1276;
  assign n1279 = ~n1277 & ~n1278;
  assign n1280 = ~po59  & n1273;
  assign n1281 = ~n1279 & ~n1280;
  assign n1282 = ~n1274 & ~n1281;
  assign n1283 = po60  & ~n1282;
  assign n1284 = ~n1132 & ~n1133;
  assign n1285 = po49  & n1284;
  assign n1286 = n1138 & ~n1285;
  assign n1287 = ~n1138 & n1285;
  assign n1288 = ~n1286 & ~n1287;
  assign n1289 = ~po60  & ~n1274;
  assign n1290 = ~n1281 & n1289;
  assign n1291 = ~n1288 & ~n1290;
  assign n1292 = ~n1283 & ~n1291;
  assign n1293 = po61  & ~n1292;
  assign n1294 = ~n1141 & ~n1143;
  assign n1295 = po49  & n1294;
  assign n1296 = n1148 & ~n1295;
  assign n1297 = ~n1148 & n1295;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = ~po61  & n1292;
  assign n1300 = ~n1298 & ~n1299;
  assign n1301 = ~n1293 & ~n1300;
  assign n1302 = po62  & ~n1301;
  assign n1303 = ~po62  & ~n1293;
  assign n1304 = ~n1300 & n1303;
  assign n1305 = ~n1151 & po49 ;
  assign n1306 = ~n1157 & n1305;
  assign n1307 = n1156 & ~n1306;
  assign n1308 = n1158 & n1305;
  assign n1309 = ~n1307 & ~n1308;
  assign n1310 = ~n1304 & n1309;
  assign n1311 = ~n1302 & ~n1310;
  assign n1312 = ~n1160 & ~n1162;
  assign n1313 = po49  & n1312;
  assign n1314 = n1167 & ~n1313;
  assign n1315 = ~n1167 & n1313;
  assign n1316 = ~n1314 & ~n1315;
  assign n1317 = n1169 & po49 ;
  assign n1318 = ~n1174 & ~n1317;
  assign n1319 = ~n1182 & ~n1318;
  assign n1320 = po49  & ~n1319;
  assign n1321 = ~n1316 & ~n1320;
  assign n1322 = ~n1311 & n1321;
  assign n1323 = ~po63  & ~n1322;
  assign n1324 = n1311 & n1316;
  assign n1325 = po63  & n1319;
  assign n1326 = ~n1324 & ~n1325;
  assign po48  = n1323 | ~n1326;
  assign n1328 = pi96  & po48 ;
  assign n1329 = ~pi94  & ~pi95 ;
  assign n1330 = ~pi96  & n1329;
  assign n1331 = ~n1328 & ~n1330;
  assign n1332 = po49  & ~n1331;
  assign n1333 = ~pi96  & po48 ;
  assign n1334 = pi97  & ~n1333;
  assign n1335 = ~pi97  & n1333;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = ~po49  & n1331;
  assign n1338 = n1336 & ~n1337;
  assign n1339 = ~n1332 & ~n1338;
  assign n1340 = po50  & ~n1339;
  assign n1341 = ~po50  & ~n1332;
  assign n1342 = ~n1338 & n1341;
  assign n1343 = po49  & ~po48 ;
  assign n1344 = ~n1335 & ~n1343;
  assign n1345 = pi98  & ~n1344;
  assign n1346 = ~pi98  & n1344;
  assign n1347 = ~n1345 & ~n1346;
  assign n1348 = ~n1342 & ~n1347;
  assign n1349 = ~n1340 & ~n1348;
  assign n1350 = po51  & ~n1349;
  assign n1351 = ~po51  & n1349;
  assign n1352 = ~n1190 & ~n1191;
  assign n1353 = po48  & n1352;
  assign n1354 = n1195 & ~n1353;
  assign n1355 = ~n1195 & n1353;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = ~n1351 & ~n1356;
  assign n1358 = ~n1350 & ~n1357;
  assign n1359 = po52  & ~n1358;
  assign n1360 = ~po52  & ~n1350;
  assign n1361 = ~n1357 & n1360;
  assign n1362 = ~n1198 & po48 ;
  assign n1363 = ~n1204 & n1362;
  assign n1364 = n1203 & ~n1363;
  assign n1365 = n1205 & n1362;
  assign n1366 = ~n1364 & ~n1365;
  assign n1367 = ~n1361 & n1366;
  assign n1368 = ~n1359 & ~n1367;
  assign n1369 = po53  & ~n1368;
  assign n1370 = ~po53  & n1368;
  assign n1371 = ~n1207 & ~n1209;
  assign n1372 = po48  & n1371;
  assign n1373 = n1214 & ~n1372;
  assign n1374 = ~n1214 & n1372;
  assign n1375 = ~n1373 & ~n1374;
  assign n1376 = ~n1370 & n1375;
  assign n1377 = ~n1369 & ~n1376;
  assign n1378 = po54  & ~n1377;
  assign n1379 = ~po54  & ~n1369;
  assign n1380 = ~n1376 & n1379;
  assign n1381 = ~n1217 & po48 ;
  assign n1382 = ~n1223 & n1381;
  assign n1383 = n1222 & ~n1382;
  assign n1384 = n1224 & n1381;
  assign n1385 = ~n1383 & ~n1384;
  assign n1386 = ~n1380 & n1385;
  assign n1387 = ~n1378 & ~n1386;
  assign n1388 = po55  & ~n1387;
  assign n1389 = ~po55  & n1387;
  assign n1390 = ~n1226 & ~n1228;
  assign n1391 = po48  & n1390;
  assign n1392 = n1233 & n1391;
  assign n1393 = ~n1233 & ~n1391;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = ~n1389 & n1394;
  assign n1396 = ~n1388 & ~n1395;
  assign n1397 = po56  & ~n1396;
  assign n1398 = ~po56  & ~n1388;
  assign n1399 = ~n1395 & n1398;
  assign n1400 = ~n1236 & po48 ;
  assign n1401 = ~n1242 & n1400;
  assign n1402 = n1241 & ~n1401;
  assign n1403 = n1243 & n1400;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = ~n1399 & n1404;
  assign n1406 = ~n1397 & ~n1405;
  assign n1407 = po57  & ~n1406;
  assign n1408 = ~po57  & n1406;
  assign n1409 = ~n1245 & ~n1247;
  assign n1410 = po48  & n1409;
  assign n1411 = ~n1252 & ~n1410;
  assign n1412 = n1252 & n1410;
  assign n1413 = ~n1411 & ~n1412;
  assign n1414 = ~n1408 & n1413;
  assign n1415 = ~n1407 & ~n1414;
  assign n1416 = po58  & ~n1415;
  assign n1417 = ~po58  & ~n1407;
  assign n1418 = ~n1414 & n1417;
  assign n1419 = ~n1255 & po48 ;
  assign n1420 = ~n1261 & n1419;
  assign n1421 = n1260 & ~n1420;
  assign n1422 = n1262 & n1419;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = ~n1418 & n1423;
  assign n1425 = ~n1416 & ~n1424;
  assign n1426 = po59  & ~n1425;
  assign n1427 = ~n1264 & ~n1266;
  assign n1428 = po48  & n1427;
  assign n1429 = n1271 & ~n1428;
  assign n1430 = ~n1271 & n1428;
  assign n1431 = ~n1429 & ~n1430;
  assign n1432 = ~po59  & n1425;
  assign n1433 = ~n1431 & ~n1432;
  assign n1434 = ~n1426 & ~n1433;
  assign n1435 = po60  & ~n1434;
  assign n1436 = ~po60  & ~n1426;
  assign n1437 = ~n1433 & n1436;
  assign n1438 = ~n1274 & po48 ;
  assign n1439 = ~n1280 & n1438;
  assign n1440 = n1279 & ~n1439;
  assign n1441 = n1281 & n1438;
  assign n1442 = ~n1440 & ~n1441;
  assign n1443 = ~n1437 & n1442;
  assign n1444 = ~n1435 & ~n1443;
  assign n1445 = po61  & ~n1444;
  assign n1446 = ~po61  & n1444;
  assign n1447 = ~n1283 & po48 ;
  assign n1448 = ~n1290 & n1447;
  assign n1449 = n1288 & ~n1448;
  assign n1450 = n1291 & n1447;
  assign n1451 = ~n1449 & ~n1450;
  assign n1452 = ~n1446 & n1451;
  assign n1453 = ~n1445 & ~n1452;
  assign n1454 = po62  & ~n1453;
  assign n1455 = ~po62  & ~n1445;
  assign n1456 = ~n1452 & n1455;
  assign n1457 = ~n1293 & po48 ;
  assign n1458 = ~n1299 & n1457;
  assign n1459 = n1298 & ~n1458;
  assign n1460 = n1300 & n1457;
  assign n1461 = ~n1459 & ~n1460;
  assign n1462 = ~n1456 & n1461;
  assign n1463 = ~n1454 & ~n1462;
  assign n1464 = ~n1302 & ~n1304;
  assign n1465 = po48  & n1464;
  assign n1466 = n1309 & ~n1465;
  assign n1467 = ~n1309 & n1465;
  assign n1468 = ~n1466 & ~n1467;
  assign n1469 = n1311 & po48 ;
  assign n1470 = ~n1316 & ~n1469;
  assign n1471 = ~n1324 & ~n1470;
  assign n1472 = po48  & ~n1471;
  assign n1473 = ~n1468 & ~n1472;
  assign n1474 = ~n1463 & n1473;
  assign n1475 = ~po63  & ~n1474;
  assign n1476 = n1463 & n1468;
  assign n1477 = po63  & n1471;
  assign n1478 = ~n1476 & ~n1477;
  assign po47  = n1475 | ~n1478;
  assign n1480 = pi94  & po47 ;
  assign n1481 = ~pi92  & ~pi93 ;
  assign n1482 = ~pi94  & n1481;
  assign n1483 = ~n1480 & ~n1482;
  assign n1484 = po48  & ~n1483;
  assign n1485 = ~po48  & n1483;
  assign n1486 = ~pi94  & po47 ;
  assign n1487 = pi95  & ~n1486;
  assign n1488 = ~pi95  & n1486;
  assign n1489 = ~n1487 & ~n1488;
  assign n1490 = ~n1485 & n1489;
  assign n1491 = ~n1484 & ~n1490;
  assign n1492 = po49  & ~n1491;
  assign n1493 = po48  & ~po47 ;
  assign n1494 = ~n1488 & ~n1493;
  assign n1495 = pi96  & ~n1494;
  assign n1496 = ~pi96  & n1494;
  assign n1497 = ~n1495 & ~n1496;
  assign n1498 = ~po49  & n1491;
  assign n1499 = ~n1497 & ~n1498;
  assign n1500 = ~n1492 & ~n1499;
  assign n1501 = po50  & ~n1500;
  assign n1502 = ~po50  & ~n1492;
  assign n1503 = ~n1499 & n1502;
  assign n1504 = ~n1332 & ~n1337;
  assign n1505 = po47  & n1504;
  assign n1506 = n1336 & ~n1505;
  assign n1507 = ~n1336 & n1505;
  assign n1508 = ~n1506 & ~n1507;
  assign n1509 = ~n1503 & ~n1508;
  assign n1510 = ~n1501 & ~n1509;
  assign n1511 = po51  & ~n1510;
  assign n1512 = ~n1340 & ~n1342;
  assign n1513 = po47  & n1512;
  assign n1514 = ~n1347 & ~n1513;
  assign n1515 = n1347 & n1513;
  assign n1516 = ~n1514 & ~n1515;
  assign n1517 = ~po51  & n1510;
  assign n1518 = ~n1516 & ~n1517;
  assign n1519 = ~n1511 & ~n1518;
  assign n1520 = po52  & ~n1519;
  assign n1521 = ~po52  & ~n1511;
  assign n1522 = ~n1518 & n1521;
  assign n1523 = ~n1350 & ~n1351;
  assign n1524 = po47  & n1523;
  assign n1525 = n1356 & ~n1524;
  assign n1526 = ~n1356 & n1524;
  assign n1527 = ~n1525 & ~n1526;
  assign n1528 = ~n1522 & n1527;
  assign n1529 = ~n1520 & ~n1528;
  assign n1530 = po53  & ~n1529;
  assign n1531 = ~n1359 & ~n1361;
  assign n1532 = po47  & n1531;
  assign n1533 = n1366 & ~n1532;
  assign n1534 = ~n1366 & n1532;
  assign n1535 = ~n1533 & ~n1534;
  assign n1536 = ~po53  & n1529;
  assign n1537 = ~n1535 & ~n1536;
  assign n1538 = ~n1530 & ~n1537;
  assign n1539 = po54  & ~n1538;
  assign n1540 = ~po54  & ~n1530;
  assign n1541 = ~n1537 & n1540;
  assign n1542 = ~n1369 & ~n1370;
  assign n1543 = po47  & n1542;
  assign n1544 = n1375 & n1543;
  assign n1545 = ~n1375 & ~n1543;
  assign n1546 = ~n1544 & ~n1545;
  assign n1547 = ~n1541 & n1546;
  assign n1548 = ~n1539 & ~n1547;
  assign n1549 = po55  & ~n1548;
  assign n1550 = ~n1378 & ~n1380;
  assign n1551 = po47  & n1550;
  assign n1552 = n1385 & ~n1551;
  assign n1553 = ~n1385 & n1551;
  assign n1554 = ~n1552 & ~n1553;
  assign n1555 = ~po55  & n1548;
  assign n1556 = ~n1554 & ~n1555;
  assign n1557 = ~n1549 & ~n1556;
  assign n1558 = po56  & ~n1557;
  assign n1559 = ~po56  & ~n1549;
  assign n1560 = ~n1556 & n1559;
  assign n1561 = ~n1388 & ~n1389;
  assign n1562 = po47  & n1561;
  assign n1563 = ~n1394 & ~n1562;
  assign n1564 = n1394 & n1562;
  assign n1565 = ~n1563 & ~n1564;
  assign n1566 = ~n1560 & n1565;
  assign n1567 = ~n1558 & ~n1566;
  assign n1568 = po57  & ~n1567;
  assign n1569 = ~n1397 & ~n1399;
  assign n1570 = po47  & n1569;
  assign n1571 = n1404 & ~n1570;
  assign n1572 = ~n1404 & n1570;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = ~po57  & n1567;
  assign n1575 = ~n1573 & ~n1574;
  assign n1576 = ~n1568 & ~n1575;
  assign n1577 = po58  & ~n1576;
  assign n1578 = ~n1407 & ~n1408;
  assign n1579 = po47  & n1578;
  assign n1580 = n1413 & ~n1579;
  assign n1581 = ~n1413 & n1579;
  assign n1582 = ~n1580 & ~n1581;
  assign n1583 = ~po58  & ~n1568;
  assign n1584 = ~n1575 & n1583;
  assign n1585 = ~n1582 & ~n1584;
  assign n1586 = ~n1577 & ~n1585;
  assign n1587 = po59  & ~n1586;
  assign n1588 = ~n1416 & ~n1418;
  assign n1589 = po47  & n1588;
  assign n1590 = n1423 & ~n1589;
  assign n1591 = ~n1423 & n1589;
  assign n1592 = ~n1590 & ~n1591;
  assign n1593 = ~po59  & n1586;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = ~n1587 & ~n1594;
  assign n1596 = po60  & ~n1595;
  assign n1597 = ~po60  & ~n1587;
  assign n1598 = ~n1594 & n1597;
  assign n1599 = ~n1426 & po47 ;
  assign n1600 = ~n1432 & n1599;
  assign n1601 = n1431 & ~n1600;
  assign n1602 = n1433 & n1599;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = ~n1598 & n1603;
  assign n1605 = ~n1596 & ~n1604;
  assign n1606 = po61  & ~n1605;
  assign n1607 = ~n1435 & ~n1437;
  assign n1608 = po47  & n1607;
  assign n1609 = n1442 & ~n1608;
  assign n1610 = ~n1442 & n1608;
  assign n1611 = ~n1609 & ~n1610;
  assign n1612 = ~po61  & n1605;
  assign n1613 = ~n1611 & ~n1612;
  assign n1614 = ~n1606 & ~n1613;
  assign n1615 = po62  & ~n1614;
  assign n1616 = ~n1445 & ~n1446;
  assign n1617 = po47  & n1616;
  assign n1618 = n1451 & ~n1617;
  assign n1619 = ~n1451 & n1617;
  assign n1620 = ~n1618 & ~n1619;
  assign n1621 = ~po62  & ~n1606;
  assign n1622 = ~n1613 & n1621;
  assign n1623 = ~n1620 & ~n1622;
  assign n1624 = ~n1615 & ~n1623;
  assign n1625 = ~n1454 & ~n1456;
  assign n1626 = po47  & n1625;
  assign n1627 = n1461 & ~n1626;
  assign n1628 = ~n1461 & n1626;
  assign n1629 = ~n1627 & ~n1628;
  assign n1630 = n1463 & po47 ;
  assign n1631 = ~n1468 & ~n1630;
  assign n1632 = ~n1476 & ~n1631;
  assign n1633 = po47  & ~n1632;
  assign n1634 = ~n1629 & ~n1633;
  assign n1635 = ~n1624 & n1634;
  assign n1636 = ~po63  & ~n1635;
  assign n1637 = n1624 & n1629;
  assign n1638 = po63  & n1632;
  assign n1639 = ~n1637 & ~n1638;
  assign po46  = n1636 | ~n1639;
  assign n1641 = pi92  & po46 ;
  assign n1642 = ~pi90  & ~pi91 ;
  assign n1643 = ~pi92  & n1642;
  assign n1644 = ~n1641 & ~n1643;
  assign n1645 = po47  & ~n1644;
  assign n1646 = ~pi92  & po46 ;
  assign n1647 = pi93  & ~n1646;
  assign n1648 = ~pi93  & n1646;
  assign n1649 = ~n1647 & ~n1648;
  assign n1650 = ~po47  & n1644;
  assign n1651 = n1649 & ~n1650;
  assign n1652 = ~n1645 & ~n1651;
  assign n1653 = po48  & ~n1652;
  assign n1654 = ~po48  & ~n1645;
  assign n1655 = ~n1651 & n1654;
  assign n1656 = po47  & ~po46 ;
  assign n1657 = ~n1648 & ~n1656;
  assign n1658 = pi94  & ~n1657;
  assign n1659 = ~pi94  & n1657;
  assign n1660 = ~n1658 & ~n1659;
  assign n1661 = ~n1655 & ~n1660;
  assign n1662 = ~n1653 & ~n1661;
  assign n1663 = po49  & ~n1662;
  assign n1664 = ~po49  & n1662;
  assign n1665 = ~n1484 & ~n1485;
  assign n1666 = po46  & n1665;
  assign n1667 = n1489 & ~n1666;
  assign n1668 = ~n1489 & n1666;
  assign n1669 = ~n1667 & ~n1668;
  assign n1670 = ~n1664 & ~n1669;
  assign n1671 = ~n1663 & ~n1670;
  assign n1672 = po50  & ~n1671;
  assign n1673 = ~po50  & ~n1663;
  assign n1674 = ~n1670 & n1673;
  assign n1675 = ~n1492 & po46 ;
  assign n1676 = ~n1498 & n1675;
  assign n1677 = n1497 & ~n1676;
  assign n1678 = n1499 & n1675;
  assign n1679 = ~n1677 & ~n1678;
  assign n1680 = ~n1674 & n1679;
  assign n1681 = ~n1672 & ~n1680;
  assign n1682 = po51  & ~n1681;
  assign n1683 = ~po51  & n1681;
  assign n1684 = ~n1501 & ~n1503;
  assign n1685 = po46  & n1684;
  assign n1686 = n1508 & ~n1685;
  assign n1687 = ~n1508 & n1685;
  assign n1688 = ~n1686 & ~n1687;
  assign n1689 = ~n1683 & n1688;
  assign n1690 = ~n1682 & ~n1689;
  assign n1691 = po52  & ~n1690;
  assign n1692 = ~po52  & ~n1682;
  assign n1693 = ~n1689 & n1692;
  assign n1694 = ~n1511 & po46 ;
  assign n1695 = ~n1517 & n1694;
  assign n1696 = n1516 & ~n1695;
  assign n1697 = n1518 & n1694;
  assign n1698 = ~n1696 & ~n1697;
  assign n1699 = ~n1693 & n1698;
  assign n1700 = ~n1691 & ~n1699;
  assign n1701 = po53  & ~n1700;
  assign n1702 = ~po53  & n1700;
  assign n1703 = ~n1520 & ~n1522;
  assign n1704 = po46  & n1703;
  assign n1705 = n1527 & n1704;
  assign n1706 = ~n1527 & ~n1704;
  assign n1707 = ~n1705 & ~n1706;
  assign n1708 = ~n1702 & n1707;
  assign n1709 = ~n1701 & ~n1708;
  assign n1710 = po54  & ~n1709;
  assign n1711 = ~po54  & ~n1701;
  assign n1712 = ~n1708 & n1711;
  assign n1713 = ~n1530 & po46 ;
  assign n1714 = ~n1536 & n1713;
  assign n1715 = n1535 & ~n1714;
  assign n1716 = n1537 & n1713;
  assign n1717 = ~n1715 & ~n1716;
  assign n1718 = ~n1712 & n1717;
  assign n1719 = ~n1710 & ~n1718;
  assign n1720 = po55  & ~n1719;
  assign n1721 = ~po55  & n1719;
  assign n1722 = ~n1539 & ~n1541;
  assign n1723 = po46  & n1722;
  assign n1724 = ~n1546 & ~n1723;
  assign n1725 = n1546 & n1723;
  assign n1726 = ~n1724 & ~n1725;
  assign n1727 = ~n1721 & n1726;
  assign n1728 = ~n1720 & ~n1727;
  assign n1729 = po56  & ~n1728;
  assign n1730 = ~po56  & ~n1720;
  assign n1731 = ~n1727 & n1730;
  assign n1732 = ~n1549 & po46 ;
  assign n1733 = ~n1555 & n1732;
  assign n1734 = n1554 & ~n1733;
  assign n1735 = n1556 & n1732;
  assign n1736 = ~n1734 & ~n1735;
  assign n1737 = ~n1731 & n1736;
  assign n1738 = ~n1729 & ~n1737;
  assign n1739 = po57  & ~n1738;
  assign n1740 = ~n1558 & ~n1560;
  assign n1741 = po46  & n1740;
  assign n1742 = n1565 & ~n1741;
  assign n1743 = ~n1565 & n1741;
  assign n1744 = ~n1742 & ~n1743;
  assign n1745 = ~po57  & n1738;
  assign n1746 = ~n1744 & ~n1745;
  assign n1747 = ~n1739 & ~n1746;
  assign n1748 = po58  & ~n1747;
  assign n1749 = ~po58  & ~n1739;
  assign n1750 = ~n1746 & n1749;
  assign n1751 = ~n1568 & po46 ;
  assign n1752 = ~n1574 & n1751;
  assign n1753 = n1573 & ~n1752;
  assign n1754 = n1575 & n1751;
  assign n1755 = ~n1753 & ~n1754;
  assign n1756 = ~n1750 & n1755;
  assign n1757 = ~n1748 & ~n1756;
  assign n1758 = po59  & ~n1757;
  assign n1759 = ~po59  & n1757;
  assign n1760 = ~n1577 & po46 ;
  assign n1761 = ~n1584 & n1760;
  assign n1762 = n1582 & ~n1761;
  assign n1763 = n1585 & n1760;
  assign n1764 = ~n1762 & ~n1763;
  assign n1765 = ~n1759 & n1764;
  assign n1766 = ~n1758 & ~n1765;
  assign n1767 = po60  & ~n1766;
  assign n1768 = ~po60  & ~n1758;
  assign n1769 = ~n1765 & n1768;
  assign n1770 = ~n1587 & po46 ;
  assign n1771 = ~n1593 & n1770;
  assign n1772 = n1592 & ~n1771;
  assign n1773 = n1594 & n1770;
  assign n1774 = ~n1772 & ~n1773;
  assign n1775 = ~n1769 & n1774;
  assign n1776 = ~n1767 & ~n1775;
  assign n1777 = po61  & ~n1776;
  assign n1778 = ~n1596 & ~n1598;
  assign n1779 = po46  & n1778;
  assign n1780 = n1603 & ~n1779;
  assign n1781 = ~n1603 & n1779;
  assign n1782 = ~n1780 & ~n1781;
  assign n1783 = ~po61  & n1776;
  assign n1784 = ~n1782 & ~n1783;
  assign n1785 = ~n1777 & ~n1784;
  assign n1786 = po62  & ~n1785;
  assign n1787 = ~po62  & ~n1777;
  assign n1788 = ~n1784 & n1787;
  assign n1789 = ~n1606 & po46 ;
  assign n1790 = ~n1612 & n1789;
  assign n1791 = n1611 & ~n1790;
  assign n1792 = n1613 & n1789;
  assign n1793 = ~n1791 & ~n1792;
  assign n1794 = ~n1788 & n1793;
  assign n1795 = ~n1786 & ~n1794;
  assign n1796 = n1624 & po46 ;
  assign n1797 = ~n1629 & ~n1796;
  assign n1798 = ~n1637 & ~n1797;
  assign n1799 = po46  & ~n1798;
  assign n1800 = ~n1615 & po46 ;
  assign n1801 = ~n1622 & n1800;
  assign n1802 = n1620 & ~n1801;
  assign n1803 = n1623 & n1800;
  assign n1804 = ~n1802 & ~n1803;
  assign n1805 = ~n1799 & n1804;
  assign n1806 = ~n1795 & n1805;
  assign n1807 = ~po63  & ~n1806;
  assign n1808 = n1795 & ~n1804;
  assign n1809 = po63  & n1798;
  assign n1810 = ~n1808 & ~n1809;
  assign po45  = n1807 | ~n1810;
  assign n1812 = pi90  & po45 ;
  assign n1813 = ~pi88  & ~pi89 ;
  assign n1814 = ~pi90  & n1813;
  assign n1815 = ~n1812 & ~n1814;
  assign n1816 = po46  & ~n1815;
  assign n1817 = ~po46  & n1815;
  assign n1818 = ~pi90  & po45 ;
  assign n1819 = pi91  & ~n1818;
  assign n1820 = ~pi91  & n1818;
  assign n1821 = ~n1819 & ~n1820;
  assign n1822 = ~n1817 & n1821;
  assign n1823 = ~n1816 & ~n1822;
  assign n1824 = po47  & ~n1823;
  assign n1825 = po46  & ~po45 ;
  assign n1826 = ~n1820 & ~n1825;
  assign n1827 = pi92  & ~n1826;
  assign n1828 = ~pi92  & n1826;
  assign n1829 = ~n1827 & ~n1828;
  assign n1830 = ~po47  & n1823;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = ~n1824 & ~n1831;
  assign n1833 = po48  & ~n1832;
  assign n1834 = ~po48  & ~n1824;
  assign n1835 = ~n1831 & n1834;
  assign n1836 = ~n1645 & ~n1650;
  assign n1837 = po45  & n1836;
  assign n1838 = n1649 & ~n1837;
  assign n1839 = ~n1649 & n1837;
  assign n1840 = ~n1838 & ~n1839;
  assign n1841 = ~n1835 & ~n1840;
  assign n1842 = ~n1833 & ~n1841;
  assign n1843 = po49  & ~n1842;
  assign n1844 = ~n1653 & ~n1655;
  assign n1845 = po45  & n1844;
  assign n1846 = ~n1660 & ~n1845;
  assign n1847 = n1660 & n1845;
  assign n1848 = ~n1846 & ~n1847;
  assign n1849 = ~po49  & n1842;
  assign n1850 = ~n1848 & ~n1849;
  assign n1851 = ~n1843 & ~n1850;
  assign n1852 = po50  & ~n1851;
  assign n1853 = ~po50  & ~n1843;
  assign n1854 = ~n1850 & n1853;
  assign n1855 = ~n1663 & ~n1664;
  assign n1856 = po45  & n1855;
  assign n1857 = n1669 & ~n1856;
  assign n1858 = ~n1669 & n1856;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = ~n1854 & n1859;
  assign n1861 = ~n1852 & ~n1860;
  assign n1862 = po51  & ~n1861;
  assign n1863 = ~n1672 & ~n1674;
  assign n1864 = po45  & n1863;
  assign n1865 = n1679 & ~n1864;
  assign n1866 = ~n1679 & n1864;
  assign n1867 = ~n1865 & ~n1866;
  assign n1868 = ~po51  & n1861;
  assign n1869 = ~n1867 & ~n1868;
  assign n1870 = ~n1862 & ~n1869;
  assign n1871 = po52  & ~n1870;
  assign n1872 = ~po52  & ~n1862;
  assign n1873 = ~n1869 & n1872;
  assign n1874 = ~n1682 & ~n1683;
  assign n1875 = po45  & n1874;
  assign n1876 = n1688 & n1875;
  assign n1877 = ~n1688 & ~n1875;
  assign n1878 = ~n1876 & ~n1877;
  assign n1879 = ~n1873 & n1878;
  assign n1880 = ~n1871 & ~n1879;
  assign n1881 = po53  & ~n1880;
  assign n1882 = ~n1691 & ~n1693;
  assign n1883 = po45  & n1882;
  assign n1884 = n1698 & ~n1883;
  assign n1885 = ~n1698 & n1883;
  assign n1886 = ~n1884 & ~n1885;
  assign n1887 = ~po53  & n1880;
  assign n1888 = ~n1886 & ~n1887;
  assign n1889 = ~n1881 & ~n1888;
  assign n1890 = po54  & ~n1889;
  assign n1891 = ~po54  & ~n1881;
  assign n1892 = ~n1888 & n1891;
  assign n1893 = ~n1701 & ~n1702;
  assign n1894 = po45  & n1893;
  assign n1895 = ~n1707 & ~n1894;
  assign n1896 = n1707 & n1894;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = ~n1892 & n1897;
  assign n1899 = ~n1890 & ~n1898;
  assign n1900 = po55  & ~n1899;
  assign n1901 = ~n1710 & ~n1712;
  assign n1902 = po45  & n1901;
  assign n1903 = n1717 & ~n1902;
  assign n1904 = ~n1717 & n1902;
  assign n1905 = ~n1903 & ~n1904;
  assign n1906 = ~po55  & n1899;
  assign n1907 = ~n1905 & ~n1906;
  assign n1908 = ~n1900 & ~n1907;
  assign n1909 = po56  & ~n1908;
  assign n1910 = ~n1720 & ~n1721;
  assign n1911 = po45  & n1910;
  assign n1912 = n1726 & ~n1911;
  assign n1913 = ~n1726 & n1911;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = ~po56  & ~n1900;
  assign n1916 = ~n1907 & n1915;
  assign n1917 = ~n1914 & ~n1916;
  assign n1918 = ~n1909 & ~n1917;
  assign n1919 = po57  & ~n1918;
  assign n1920 = ~n1729 & ~n1731;
  assign n1921 = po45  & n1920;
  assign n1922 = n1736 & ~n1921;
  assign n1923 = ~n1736 & n1921;
  assign n1924 = ~n1922 & ~n1923;
  assign n1925 = ~po57  & n1918;
  assign n1926 = ~n1924 & ~n1925;
  assign n1927 = ~n1919 & ~n1926;
  assign n1928 = po58  & ~n1927;
  assign n1929 = ~po58  & ~n1919;
  assign n1930 = ~n1926 & n1929;
  assign n1931 = ~n1739 & po45 ;
  assign n1932 = ~n1745 & n1931;
  assign n1933 = n1744 & ~n1932;
  assign n1934 = n1746 & n1931;
  assign n1935 = ~n1933 & ~n1934;
  assign n1936 = ~n1930 & n1935;
  assign n1937 = ~n1928 & ~n1936;
  assign n1938 = po59  & ~n1937;
  assign n1939 = ~n1748 & ~n1750;
  assign n1940 = po45  & n1939;
  assign n1941 = n1755 & ~n1940;
  assign n1942 = ~n1755 & n1940;
  assign n1943 = ~n1941 & ~n1942;
  assign n1944 = ~po59  & n1937;
  assign n1945 = ~n1943 & ~n1944;
  assign n1946 = ~n1938 & ~n1945;
  assign n1947 = po60  & ~n1946;
  assign n1948 = ~n1758 & ~n1759;
  assign n1949 = po45  & n1948;
  assign n1950 = n1764 & ~n1949;
  assign n1951 = ~n1764 & n1949;
  assign n1952 = ~n1950 & ~n1951;
  assign n1953 = ~po60  & ~n1938;
  assign n1954 = ~n1945 & n1953;
  assign n1955 = ~n1952 & ~n1954;
  assign n1956 = ~n1947 & ~n1955;
  assign n1957 = po61  & ~n1956;
  assign n1958 = ~n1767 & ~n1769;
  assign n1959 = po45  & n1958;
  assign n1960 = n1774 & ~n1959;
  assign n1961 = ~n1774 & n1959;
  assign n1962 = ~n1960 & ~n1961;
  assign n1963 = ~po61  & n1956;
  assign n1964 = ~n1962 & ~n1963;
  assign n1965 = ~n1957 & ~n1964;
  assign n1966 = po62  & ~n1965;
  assign n1967 = ~po62  & ~n1957;
  assign n1968 = ~n1964 & n1967;
  assign n1969 = ~n1777 & po45 ;
  assign n1970 = ~n1783 & n1969;
  assign n1971 = n1782 & ~n1970;
  assign n1972 = n1784 & n1969;
  assign n1973 = ~n1971 & ~n1972;
  assign n1974 = ~n1968 & n1973;
  assign n1975 = ~n1966 & ~n1974;
  assign n1976 = n1804 & po45 ;
  assign n1977 = ~n1795 & n1976;
  assign n1978 = ~n1786 & ~n1788;
  assign n1979 = po45  & n1978;
  assign n1980 = n1793 & ~n1979;
  assign n1981 = ~n1793 & n1979;
  assign n1982 = ~n1980 & ~n1981;
  assign n1983 = ~n1808 & ~n1977;
  assign n1984 = ~n1982 & n1983;
  assign n1985 = ~n1975 & n1984;
  assign n1986 = ~po63  & ~n1985;
  assign n1987 = n1975 & n1982;
  assign n1988 = n1795 & ~n1976;
  assign n1989 = ~n1795 & n1804;
  assign n1990 = po63  & ~n1989;
  assign n1991 = ~n1988 & n1990;
  assign n1992 = ~n1987 & ~n1991;
  assign po44  = n1986 | ~n1992;
  assign n1994 = pi88  & po44 ;
  assign n1995 = ~pi86  & ~pi87 ;
  assign n1996 = ~pi88  & n1995;
  assign n1997 = ~n1994 & ~n1996;
  assign n1998 = po45  & ~n1997;
  assign n1999 = ~pi88  & po44 ;
  assign n2000 = pi89  & ~n1999;
  assign n2001 = ~pi89  & n1999;
  assign n2002 = ~n2000 & ~n2001;
  assign n2003 = ~po45  & n1997;
  assign n2004 = n2002 & ~n2003;
  assign n2005 = ~n1998 & ~n2004;
  assign n2006 = po46  & ~n2005;
  assign n2007 = ~po46  & ~n1998;
  assign n2008 = ~n2004 & n2007;
  assign n2009 = po45  & ~po44 ;
  assign n2010 = ~n2001 & ~n2009;
  assign n2011 = pi90  & ~n2010;
  assign n2012 = ~pi90  & n2010;
  assign n2013 = ~n2011 & ~n2012;
  assign n2014 = ~n2008 & ~n2013;
  assign n2015 = ~n2006 & ~n2014;
  assign n2016 = po47  & ~n2015;
  assign n2017 = ~po47  & n2015;
  assign n2018 = ~n1816 & ~n1817;
  assign n2019 = po44  & n2018;
  assign n2020 = n1821 & ~n2019;
  assign n2021 = ~n1821 & n2019;
  assign n2022 = ~n2020 & ~n2021;
  assign n2023 = ~n2017 & ~n2022;
  assign n2024 = ~n2016 & ~n2023;
  assign n2025 = po48  & ~n2024;
  assign n2026 = ~po48  & ~n2016;
  assign n2027 = ~n2023 & n2026;
  assign n2028 = ~n1824 & po44 ;
  assign n2029 = ~n1830 & n2028;
  assign n2030 = n1829 & ~n2029;
  assign n2031 = n1831 & n2028;
  assign n2032 = ~n2030 & ~n2031;
  assign n2033 = ~n2027 & n2032;
  assign n2034 = ~n2025 & ~n2033;
  assign n2035 = po49  & ~n2034;
  assign n2036 = ~po49  & n2034;
  assign n2037 = ~n1833 & ~n1835;
  assign n2038 = po44  & n2037;
  assign n2039 = n1840 & ~n2038;
  assign n2040 = ~n1840 & n2038;
  assign n2041 = ~n2039 & ~n2040;
  assign n2042 = ~n2036 & n2041;
  assign n2043 = ~n2035 & ~n2042;
  assign n2044 = po50  & ~n2043;
  assign n2045 = ~po50  & ~n2035;
  assign n2046 = ~n2042 & n2045;
  assign n2047 = ~n1843 & po44 ;
  assign n2048 = ~n1849 & n2047;
  assign n2049 = n1848 & ~n2048;
  assign n2050 = n1850 & n2047;
  assign n2051 = ~n2049 & ~n2050;
  assign n2052 = ~n2046 & n2051;
  assign n2053 = ~n2044 & ~n2052;
  assign n2054 = po51  & ~n2053;
  assign n2055 = ~po51  & n2053;
  assign n2056 = ~n1852 & ~n1854;
  assign n2057 = po44  & n2056;
  assign n2058 = n1859 & n2057;
  assign n2059 = ~n1859 & ~n2057;
  assign n2060 = ~n2058 & ~n2059;
  assign n2061 = ~n2055 & n2060;
  assign n2062 = ~n2054 & ~n2061;
  assign n2063 = po52  & ~n2062;
  assign n2064 = ~po52  & ~n2054;
  assign n2065 = ~n2061 & n2064;
  assign n2066 = ~n1862 & po44 ;
  assign n2067 = ~n1868 & n2066;
  assign n2068 = n1867 & ~n2067;
  assign n2069 = n1869 & n2066;
  assign n2070 = ~n2068 & ~n2069;
  assign n2071 = ~n2065 & n2070;
  assign n2072 = ~n2063 & ~n2071;
  assign n2073 = po53  & ~n2072;
  assign n2074 = ~po53  & n2072;
  assign n2075 = ~n1871 & ~n1873;
  assign n2076 = po44  & n2075;
  assign n2077 = n1878 & n2076;
  assign n2078 = ~n1878 & ~n2076;
  assign n2079 = ~n2077 & ~n2078;
  assign n2080 = ~n2074 & n2079;
  assign n2081 = ~n2073 & ~n2080;
  assign n2082 = po54  & ~n2081;
  assign n2083 = ~po54  & ~n2073;
  assign n2084 = ~n2080 & n2083;
  assign n2085 = ~n1881 & po44 ;
  assign n2086 = ~n1887 & n2085;
  assign n2087 = n1886 & ~n2086;
  assign n2088 = n1888 & n2085;
  assign n2089 = ~n2087 & ~n2088;
  assign n2090 = ~n2084 & n2089;
  assign n2091 = ~n2082 & ~n2090;
  assign n2092 = po55  & ~n2091;
  assign n2093 = ~n1890 & ~n1892;
  assign n2094 = po44  & n2093;
  assign n2095 = n1897 & ~n2094;
  assign n2096 = ~n1897 & n2094;
  assign n2097 = ~n2095 & ~n2096;
  assign n2098 = ~po55  & n2091;
  assign n2099 = ~n2097 & ~n2098;
  assign n2100 = ~n2092 & ~n2099;
  assign n2101 = po56  & ~n2100;
  assign n2102 = ~po56  & ~n2092;
  assign n2103 = ~n2099 & n2102;
  assign n2104 = ~n1900 & po44 ;
  assign n2105 = ~n1906 & n2104;
  assign n2106 = n1905 & ~n2105;
  assign n2107 = n1907 & n2104;
  assign n2108 = ~n2106 & ~n2107;
  assign n2109 = ~n2103 & n2108;
  assign n2110 = ~n2101 & ~n2109;
  assign n2111 = po57  & ~n2110;
  assign n2112 = ~po57  & n2110;
  assign n2113 = ~n1909 & po44 ;
  assign n2114 = ~n1916 & n2113;
  assign n2115 = n1914 & ~n2114;
  assign n2116 = n1917 & n2113;
  assign n2117 = ~n2115 & ~n2116;
  assign n2118 = ~n2112 & n2117;
  assign n2119 = ~n2111 & ~n2118;
  assign n2120 = po58  & ~n2119;
  assign n2121 = ~po58  & ~n2111;
  assign n2122 = ~n2118 & n2121;
  assign n2123 = ~n1919 & po44 ;
  assign n2124 = ~n1925 & n2123;
  assign n2125 = n1924 & ~n2124;
  assign n2126 = n1926 & n2123;
  assign n2127 = ~n2125 & ~n2126;
  assign n2128 = ~n2122 & n2127;
  assign n2129 = ~n2120 & ~n2128;
  assign n2130 = po59  & ~n2129;
  assign n2131 = ~n1928 & ~n1930;
  assign n2132 = po44  & n2131;
  assign n2133 = n1935 & ~n2132;
  assign n2134 = ~n1935 & n2132;
  assign n2135 = ~n2133 & ~n2134;
  assign n2136 = ~po59  & n2129;
  assign n2137 = ~n2135 & ~n2136;
  assign n2138 = ~n2130 & ~n2137;
  assign n2139 = po60  & ~n2138;
  assign n2140 = ~po60  & ~n2130;
  assign n2141 = ~n2137 & n2140;
  assign n2142 = ~n1938 & po44 ;
  assign n2143 = ~n1944 & n2142;
  assign n2144 = n1943 & ~n2143;
  assign n2145 = n1945 & n2142;
  assign n2146 = ~n2144 & ~n2145;
  assign n2147 = ~n2141 & n2146;
  assign n2148 = ~n2139 & ~n2147;
  assign n2149 = po61  & ~n2148;
  assign n2150 = ~po61  & n2148;
  assign n2151 = ~n1947 & po44 ;
  assign n2152 = ~n1954 & n2151;
  assign n2153 = n1952 & ~n2152;
  assign n2154 = n1955 & n2151;
  assign n2155 = ~n2153 & ~n2154;
  assign n2156 = ~n2150 & n2155;
  assign n2157 = ~n2149 & ~n2156;
  assign n2158 = po62  & ~n2157;
  assign n2159 = ~po62  & ~n2149;
  assign n2160 = ~n2156 & n2159;
  assign n2161 = ~n1957 & po44 ;
  assign n2162 = ~n1963 & n2161;
  assign n2163 = n1962 & ~n2162;
  assign n2164 = n1964 & n2161;
  assign n2165 = ~n2163 & ~n2164;
  assign n2166 = ~n2160 & n2165;
  assign n2167 = ~n2158 & ~n2166;
  assign n2168 = ~n1966 & ~n1968;
  assign n2169 = po44  & n2168;
  assign n2170 = n1973 & ~n2169;
  assign n2171 = ~n1973 & n2169;
  assign n2172 = ~n2170 & ~n2171;
  assign n2173 = n1975 & po44 ;
  assign n2174 = ~n1982 & ~n2173;
  assign n2175 = ~n1987 & ~n2174;
  assign n2176 = po44  & ~n2175;
  assign n2177 = ~n2172 & ~n2176;
  assign n2178 = ~n2167 & n2177;
  assign n2179 = ~po63  & ~n2178;
  assign n2180 = n2167 & n2172;
  assign n2181 = po63  & n2175;
  assign n2182 = ~n2180 & ~n2181;
  assign po43  = n2179 | ~n2182;
  assign n2184 = pi86  & po43 ;
  assign n2185 = ~pi84  & ~pi85 ;
  assign n2186 = ~pi86  & n2185;
  assign n2187 = ~n2184 & ~n2186;
  assign n2188 = po44  & ~n2187;
  assign n2189 = ~po44  & n2187;
  assign n2190 = ~pi86  & po43 ;
  assign n2191 = pi87  & ~n2190;
  assign n2192 = ~pi87  & n2190;
  assign n2193 = ~n2191 & ~n2192;
  assign n2194 = ~n2189 & n2193;
  assign n2195 = ~n2188 & ~n2194;
  assign n2196 = po45  & ~n2195;
  assign n2197 = po44  & ~po43 ;
  assign n2198 = ~n2192 & ~n2197;
  assign n2199 = pi88  & ~n2198;
  assign n2200 = ~pi88  & n2198;
  assign n2201 = ~n2199 & ~n2200;
  assign n2202 = ~po45  & n2195;
  assign n2203 = ~n2201 & ~n2202;
  assign n2204 = ~n2196 & ~n2203;
  assign n2205 = po46  & ~n2204;
  assign n2206 = ~po46  & ~n2196;
  assign n2207 = ~n2203 & n2206;
  assign n2208 = ~n1998 & ~n2003;
  assign n2209 = po43  & n2208;
  assign n2210 = n2002 & ~n2209;
  assign n2211 = ~n2002 & n2209;
  assign n2212 = ~n2210 & ~n2211;
  assign n2213 = ~n2207 & ~n2212;
  assign n2214 = ~n2205 & ~n2213;
  assign n2215 = po47  & ~n2214;
  assign n2216 = ~n2006 & ~n2008;
  assign n2217 = po43  & n2216;
  assign n2218 = ~n2013 & ~n2217;
  assign n2219 = n2013 & n2217;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = ~po47  & n2214;
  assign n2222 = ~n2220 & ~n2221;
  assign n2223 = ~n2215 & ~n2222;
  assign n2224 = po48  & ~n2223;
  assign n2225 = ~po48  & ~n2215;
  assign n2226 = ~n2222 & n2225;
  assign n2227 = ~n2016 & ~n2017;
  assign n2228 = po43  & n2227;
  assign n2229 = n2022 & ~n2228;
  assign n2230 = ~n2022 & n2228;
  assign n2231 = ~n2229 & ~n2230;
  assign n2232 = ~n2226 & n2231;
  assign n2233 = ~n2224 & ~n2232;
  assign n2234 = po49  & ~n2233;
  assign n2235 = ~n2025 & ~n2027;
  assign n2236 = po43  & n2235;
  assign n2237 = n2032 & ~n2236;
  assign n2238 = ~n2032 & n2236;
  assign n2239 = ~n2237 & ~n2238;
  assign n2240 = ~po49  & n2233;
  assign n2241 = ~n2239 & ~n2240;
  assign n2242 = ~n2234 & ~n2241;
  assign n2243 = po50  & ~n2242;
  assign n2244 = ~po50  & ~n2234;
  assign n2245 = ~n2241 & n2244;
  assign n2246 = ~n2035 & ~n2036;
  assign n2247 = po43  & n2246;
  assign n2248 = n2041 & n2247;
  assign n2249 = ~n2041 & ~n2247;
  assign n2250 = ~n2248 & ~n2249;
  assign n2251 = ~n2245 & n2250;
  assign n2252 = ~n2243 & ~n2251;
  assign n2253 = po51  & ~n2252;
  assign n2254 = ~n2044 & ~n2046;
  assign n2255 = po43  & n2254;
  assign n2256 = n2051 & ~n2255;
  assign n2257 = ~n2051 & n2255;
  assign n2258 = ~n2256 & ~n2257;
  assign n2259 = ~po51  & n2252;
  assign n2260 = ~n2258 & ~n2259;
  assign n2261 = ~n2253 & ~n2260;
  assign n2262 = po52  & ~n2261;
  assign n2263 = ~po52  & ~n2253;
  assign n2264 = ~n2260 & n2263;
  assign n2265 = ~n2054 & ~n2055;
  assign n2266 = po43  & n2265;
  assign n2267 = ~n2060 & ~n2266;
  assign n2268 = n2060 & n2266;
  assign n2269 = ~n2267 & ~n2268;
  assign n2270 = ~n2264 & n2269;
  assign n2271 = ~n2262 & ~n2270;
  assign n2272 = po53  & ~n2271;
  assign n2273 = ~n2063 & ~n2065;
  assign n2274 = po43  & n2273;
  assign n2275 = n2070 & ~n2274;
  assign n2276 = ~n2070 & n2274;
  assign n2277 = ~n2275 & ~n2276;
  assign n2278 = ~po53  & n2271;
  assign n2279 = ~n2277 & ~n2278;
  assign n2280 = ~n2272 & ~n2279;
  assign n2281 = po54  & ~n2280;
  assign n2282 = ~po54  & ~n2272;
  assign n2283 = ~n2279 & n2282;
  assign n2284 = ~n2073 & ~n2074;
  assign n2285 = po43  & n2284;
  assign n2286 = ~n2079 & ~n2285;
  assign n2287 = n2079 & n2285;
  assign n2288 = ~n2286 & ~n2287;
  assign n2289 = ~n2283 & n2288;
  assign n2290 = ~n2281 & ~n2289;
  assign n2291 = po55  & ~n2290;
  assign n2292 = ~n2082 & ~n2084;
  assign n2293 = po43  & n2292;
  assign n2294 = n2089 & ~n2293;
  assign n2295 = ~n2089 & n2293;
  assign n2296 = ~n2294 & ~n2295;
  assign n2297 = ~po55  & n2290;
  assign n2298 = ~n2296 & ~n2297;
  assign n2299 = ~n2291 & ~n2298;
  assign n2300 = po56  & ~n2299;
  assign n2301 = ~po56  & ~n2291;
  assign n2302 = ~n2298 & n2301;
  assign n2303 = ~n2092 & po43 ;
  assign n2304 = ~n2098 & n2303;
  assign n2305 = n2097 & ~n2304;
  assign n2306 = n2099 & n2303;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = ~n2302 & n2307;
  assign n2309 = ~n2300 & ~n2308;
  assign n2310 = po57  & ~n2309;
  assign n2311 = ~n2101 & ~n2103;
  assign n2312 = po43  & n2311;
  assign n2313 = n2108 & ~n2312;
  assign n2314 = ~n2108 & n2312;
  assign n2315 = ~n2313 & ~n2314;
  assign n2316 = ~po57  & n2309;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = ~n2310 & ~n2317;
  assign n2319 = po58  & ~n2318;
  assign n2320 = ~n2111 & ~n2112;
  assign n2321 = po43  & n2320;
  assign n2322 = n2117 & ~n2321;
  assign n2323 = ~n2117 & n2321;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = ~po58  & ~n2310;
  assign n2326 = ~n2317 & n2325;
  assign n2327 = ~n2324 & ~n2326;
  assign n2328 = ~n2319 & ~n2327;
  assign n2329 = po59  & ~n2328;
  assign n2330 = ~n2120 & ~n2122;
  assign n2331 = po43  & n2330;
  assign n2332 = n2127 & ~n2331;
  assign n2333 = ~n2127 & n2331;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = ~po59  & n2328;
  assign n2336 = ~n2334 & ~n2335;
  assign n2337 = ~n2329 & ~n2336;
  assign n2338 = po60  & ~n2337;
  assign n2339 = ~po60  & ~n2329;
  assign n2340 = ~n2336 & n2339;
  assign n2341 = ~n2130 & po43 ;
  assign n2342 = ~n2136 & n2341;
  assign n2343 = n2135 & ~n2342;
  assign n2344 = n2137 & n2341;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = ~n2340 & n2345;
  assign n2347 = ~n2338 & ~n2346;
  assign n2348 = po61  & ~n2347;
  assign n2349 = ~n2139 & ~n2141;
  assign n2350 = po43  & n2349;
  assign n2351 = n2146 & ~n2350;
  assign n2352 = ~n2146 & n2350;
  assign n2353 = ~n2351 & ~n2352;
  assign n2354 = ~po61  & n2347;
  assign n2355 = ~n2353 & ~n2354;
  assign n2356 = ~n2348 & ~n2355;
  assign n2357 = po62  & ~n2356;
  assign n2358 = ~n2149 & ~n2150;
  assign n2359 = po43  & n2358;
  assign n2360 = n2155 & ~n2359;
  assign n2361 = ~n2155 & n2359;
  assign n2362 = ~n2360 & ~n2361;
  assign n2363 = ~po62  & ~n2348;
  assign n2364 = ~n2355 & n2363;
  assign n2365 = ~n2362 & ~n2364;
  assign n2366 = ~n2357 & ~n2365;
  assign n2367 = ~n2158 & ~n2160;
  assign n2368 = po43  & n2367;
  assign n2369 = n2165 & ~n2368;
  assign n2370 = ~n2165 & n2368;
  assign n2371 = ~n2369 & ~n2370;
  assign n2372 = n2167 & po43 ;
  assign n2373 = ~n2172 & ~n2372;
  assign n2374 = ~n2180 & ~n2373;
  assign n2375 = po43  & ~n2374;
  assign n2376 = ~n2371 & ~n2375;
  assign n2377 = ~n2366 & n2376;
  assign n2378 = ~po63  & ~n2377;
  assign n2379 = n2366 & n2371;
  assign n2380 = po63  & n2374;
  assign n2381 = ~n2379 & ~n2380;
  assign po42  = n2378 | ~n2381;
  assign n2383 = pi84  & po42 ;
  assign n2384 = ~pi82  & ~pi83 ;
  assign n2385 = ~pi84  & n2384;
  assign n2386 = ~n2383 & ~n2385;
  assign n2387 = po43  & ~n2386;
  assign n2388 = ~pi84  & po42 ;
  assign n2389 = pi85  & ~n2388;
  assign n2390 = ~pi85  & n2388;
  assign n2391 = ~n2389 & ~n2390;
  assign n2392 = ~po43  & n2386;
  assign n2393 = n2391 & ~n2392;
  assign n2394 = ~n2387 & ~n2393;
  assign n2395 = po44  & ~n2394;
  assign n2396 = ~po44  & ~n2387;
  assign n2397 = ~n2393 & n2396;
  assign n2398 = po43  & ~po42 ;
  assign n2399 = ~n2390 & ~n2398;
  assign n2400 = pi86  & ~n2399;
  assign n2401 = ~pi86  & n2399;
  assign n2402 = ~n2400 & ~n2401;
  assign n2403 = ~n2397 & ~n2402;
  assign n2404 = ~n2395 & ~n2403;
  assign n2405 = po45  & ~n2404;
  assign n2406 = ~po45  & n2404;
  assign n2407 = ~n2188 & ~n2189;
  assign n2408 = po42  & n2407;
  assign n2409 = n2193 & ~n2408;
  assign n2410 = ~n2193 & n2408;
  assign n2411 = ~n2409 & ~n2410;
  assign n2412 = ~n2406 & ~n2411;
  assign n2413 = ~n2405 & ~n2412;
  assign n2414 = po46  & ~n2413;
  assign n2415 = ~po46  & ~n2405;
  assign n2416 = ~n2412 & n2415;
  assign n2417 = ~n2196 & po42 ;
  assign n2418 = ~n2202 & n2417;
  assign n2419 = n2201 & ~n2418;
  assign n2420 = n2203 & n2417;
  assign n2421 = ~n2419 & ~n2420;
  assign n2422 = ~n2416 & n2421;
  assign n2423 = ~n2414 & ~n2422;
  assign n2424 = po47  & ~n2423;
  assign n2425 = ~po47  & n2423;
  assign n2426 = ~n2205 & ~n2207;
  assign n2427 = po42  & n2426;
  assign n2428 = n2212 & ~n2427;
  assign n2429 = ~n2212 & n2427;
  assign n2430 = ~n2428 & ~n2429;
  assign n2431 = ~n2425 & n2430;
  assign n2432 = ~n2424 & ~n2431;
  assign n2433 = po48  & ~n2432;
  assign n2434 = ~po48  & ~n2424;
  assign n2435 = ~n2431 & n2434;
  assign n2436 = ~n2215 & po42 ;
  assign n2437 = ~n2221 & n2436;
  assign n2438 = n2220 & ~n2437;
  assign n2439 = n2222 & n2436;
  assign n2440 = ~n2438 & ~n2439;
  assign n2441 = ~n2435 & n2440;
  assign n2442 = ~n2433 & ~n2441;
  assign n2443 = po49  & ~n2442;
  assign n2444 = ~po49  & n2442;
  assign n2445 = ~n2224 & ~n2226;
  assign n2446 = po42  & n2445;
  assign n2447 = n2231 & n2446;
  assign n2448 = ~n2231 & ~n2446;
  assign n2449 = ~n2447 & ~n2448;
  assign n2450 = ~n2444 & n2449;
  assign n2451 = ~n2443 & ~n2450;
  assign n2452 = po50  & ~n2451;
  assign n2453 = ~po50  & ~n2443;
  assign n2454 = ~n2450 & n2453;
  assign n2455 = ~n2234 & po42 ;
  assign n2456 = ~n2240 & n2455;
  assign n2457 = n2239 & ~n2456;
  assign n2458 = n2241 & n2455;
  assign n2459 = ~n2457 & ~n2458;
  assign n2460 = ~n2454 & n2459;
  assign n2461 = ~n2452 & ~n2460;
  assign n2462 = po51  & ~n2461;
  assign n2463 = ~po51  & n2461;
  assign n2464 = ~n2243 & ~n2245;
  assign n2465 = po42  & n2464;
  assign n2466 = ~n2250 & ~n2465;
  assign n2467 = n2250 & n2465;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = ~n2463 & n2468;
  assign n2470 = ~n2462 & ~n2469;
  assign n2471 = po52  & ~n2470;
  assign n2472 = ~po52  & ~n2462;
  assign n2473 = ~n2469 & n2472;
  assign n2474 = ~n2253 & po42 ;
  assign n2475 = ~n2259 & n2474;
  assign n2476 = n2258 & ~n2475;
  assign n2477 = n2260 & n2474;
  assign n2478 = ~n2476 & ~n2477;
  assign n2479 = ~n2473 & n2478;
  assign n2480 = ~n2471 & ~n2479;
  assign n2481 = po53  & ~n2480;
  assign n2482 = ~n2262 & ~n2264;
  assign n2483 = po42  & n2482;
  assign n2484 = n2269 & ~n2483;
  assign n2485 = ~n2269 & n2483;
  assign n2486 = ~n2484 & ~n2485;
  assign n2487 = ~po53  & n2480;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = ~n2481 & ~n2488;
  assign n2490 = po54  & ~n2489;
  assign n2491 = ~po54  & ~n2481;
  assign n2492 = ~n2488 & n2491;
  assign n2493 = ~n2272 & po42 ;
  assign n2494 = ~n2278 & n2493;
  assign n2495 = n2277 & ~n2494;
  assign n2496 = n2279 & n2493;
  assign n2497 = ~n2495 & ~n2496;
  assign n2498 = ~n2492 & n2497;
  assign n2499 = ~n2490 & ~n2498;
  assign n2500 = po55  & ~n2499;
  assign n2501 = ~n2281 & ~n2283;
  assign n2502 = po42  & n2501;
  assign n2503 = n2288 & ~n2502;
  assign n2504 = ~n2288 & n2502;
  assign n2505 = ~n2503 & ~n2504;
  assign n2506 = ~po55  & n2499;
  assign n2507 = ~n2505 & ~n2506;
  assign n2508 = ~n2500 & ~n2507;
  assign n2509 = po56  & ~n2508;
  assign n2510 = ~po56  & ~n2500;
  assign n2511 = ~n2507 & n2510;
  assign n2512 = ~n2291 & po42 ;
  assign n2513 = ~n2297 & n2512;
  assign n2514 = n2296 & ~n2513;
  assign n2515 = n2298 & n2512;
  assign n2516 = ~n2514 & ~n2515;
  assign n2517 = ~n2511 & n2516;
  assign n2518 = ~n2509 & ~n2517;
  assign n2519 = po57  & ~n2518;
  assign n2520 = ~n2300 & ~n2302;
  assign n2521 = po42  & n2520;
  assign n2522 = n2307 & ~n2521;
  assign n2523 = ~n2307 & n2521;
  assign n2524 = ~n2522 & ~n2523;
  assign n2525 = ~po57  & n2518;
  assign n2526 = ~n2524 & ~n2525;
  assign n2527 = ~n2519 & ~n2526;
  assign n2528 = po58  & ~n2527;
  assign n2529 = ~po58  & ~n2519;
  assign n2530 = ~n2526 & n2529;
  assign n2531 = ~n2310 & po42 ;
  assign n2532 = ~n2316 & n2531;
  assign n2533 = n2315 & ~n2532;
  assign n2534 = n2317 & n2531;
  assign n2535 = ~n2533 & ~n2534;
  assign n2536 = ~n2530 & n2535;
  assign n2537 = ~n2528 & ~n2536;
  assign n2538 = po59  & ~n2537;
  assign n2539 = ~po59  & n2537;
  assign n2540 = ~n2319 & po42 ;
  assign n2541 = ~n2326 & n2540;
  assign n2542 = n2324 & ~n2541;
  assign n2543 = n2327 & n2540;
  assign n2544 = ~n2542 & ~n2543;
  assign n2545 = ~n2539 & n2544;
  assign n2546 = ~n2538 & ~n2545;
  assign n2547 = po60  & ~n2546;
  assign n2548 = ~po60  & ~n2538;
  assign n2549 = ~n2545 & n2548;
  assign n2550 = ~n2329 & po42 ;
  assign n2551 = ~n2335 & n2550;
  assign n2552 = n2334 & ~n2551;
  assign n2553 = n2336 & n2550;
  assign n2554 = ~n2552 & ~n2553;
  assign n2555 = ~n2549 & n2554;
  assign n2556 = ~n2547 & ~n2555;
  assign n2557 = po61  & ~n2556;
  assign n2558 = ~n2338 & ~n2340;
  assign n2559 = po42  & n2558;
  assign n2560 = n2345 & ~n2559;
  assign n2561 = ~n2345 & n2559;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = ~po61  & n2556;
  assign n2564 = ~n2562 & ~n2563;
  assign n2565 = ~n2557 & ~n2564;
  assign n2566 = po62  & ~n2565;
  assign n2567 = ~po62  & ~n2557;
  assign n2568 = ~n2564 & n2567;
  assign n2569 = ~n2348 & po42 ;
  assign n2570 = ~n2354 & n2569;
  assign n2571 = n2353 & ~n2570;
  assign n2572 = n2355 & n2569;
  assign n2573 = ~n2571 & ~n2572;
  assign n2574 = ~n2568 & n2573;
  assign n2575 = ~n2566 & ~n2574;
  assign n2576 = n2366 & po42 ;
  assign n2577 = ~n2371 & ~n2576;
  assign n2578 = ~n2379 & ~n2577;
  assign n2579 = po42  & ~n2578;
  assign n2580 = ~n2357 & po42 ;
  assign n2581 = ~n2364 & n2580;
  assign n2582 = n2362 & ~n2581;
  assign n2583 = n2365 & n2580;
  assign n2584 = ~n2582 & ~n2583;
  assign n2585 = ~n2579 & n2584;
  assign n2586 = ~n2575 & n2585;
  assign n2587 = ~po63  & ~n2586;
  assign n2588 = n2575 & ~n2584;
  assign n2589 = po63  & n2578;
  assign n2590 = ~n2588 & ~n2589;
  assign po41  = n2587 | ~n2590;
  assign n2592 = pi82  & po41 ;
  assign n2593 = ~pi80  & ~pi81 ;
  assign n2594 = ~pi82  & n2593;
  assign n2595 = ~n2592 & ~n2594;
  assign n2596 = po42  & ~n2595;
  assign n2597 = ~po42  & n2595;
  assign n2598 = ~pi82  & po41 ;
  assign n2599 = pi83  & ~n2598;
  assign n2600 = ~pi83  & n2598;
  assign n2601 = ~n2599 & ~n2600;
  assign n2602 = ~n2597 & n2601;
  assign n2603 = ~n2596 & ~n2602;
  assign n2604 = po43  & ~n2603;
  assign n2605 = po42  & ~po41 ;
  assign n2606 = ~n2600 & ~n2605;
  assign n2607 = pi84  & ~n2606;
  assign n2608 = ~pi84  & n2606;
  assign n2609 = ~n2607 & ~n2608;
  assign n2610 = ~po43  & n2603;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = ~n2604 & ~n2611;
  assign n2613 = po44  & ~n2612;
  assign n2614 = ~po44  & ~n2604;
  assign n2615 = ~n2611 & n2614;
  assign n2616 = ~n2387 & ~n2392;
  assign n2617 = po41  & n2616;
  assign n2618 = n2391 & ~n2617;
  assign n2619 = ~n2391 & n2617;
  assign n2620 = ~n2618 & ~n2619;
  assign n2621 = ~n2615 & ~n2620;
  assign n2622 = ~n2613 & ~n2621;
  assign n2623 = po45  & ~n2622;
  assign n2624 = ~n2395 & ~n2397;
  assign n2625 = po41  & n2624;
  assign n2626 = ~n2402 & ~n2625;
  assign n2627 = n2402 & n2625;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = ~po45  & n2622;
  assign n2630 = ~n2628 & ~n2629;
  assign n2631 = ~n2623 & ~n2630;
  assign n2632 = po46  & ~n2631;
  assign n2633 = ~po46  & ~n2623;
  assign n2634 = ~n2630 & n2633;
  assign n2635 = ~n2405 & ~n2406;
  assign n2636 = po41  & n2635;
  assign n2637 = n2411 & ~n2636;
  assign n2638 = ~n2411 & n2636;
  assign n2639 = ~n2637 & ~n2638;
  assign n2640 = ~n2634 & n2639;
  assign n2641 = ~n2632 & ~n2640;
  assign n2642 = po47  & ~n2641;
  assign n2643 = ~n2414 & ~n2416;
  assign n2644 = po41  & n2643;
  assign n2645 = n2421 & ~n2644;
  assign n2646 = ~n2421 & n2644;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = ~po47  & n2641;
  assign n2649 = ~n2647 & ~n2648;
  assign n2650 = ~n2642 & ~n2649;
  assign n2651 = po48  & ~n2650;
  assign n2652 = ~po48  & ~n2642;
  assign n2653 = ~n2649 & n2652;
  assign n2654 = ~n2424 & ~n2425;
  assign n2655 = po41  & n2654;
  assign n2656 = n2430 & n2655;
  assign n2657 = ~n2430 & ~n2655;
  assign n2658 = ~n2656 & ~n2657;
  assign n2659 = ~n2653 & n2658;
  assign n2660 = ~n2651 & ~n2659;
  assign n2661 = po49  & ~n2660;
  assign n2662 = ~n2433 & ~n2435;
  assign n2663 = po41  & n2662;
  assign n2664 = n2440 & ~n2663;
  assign n2665 = ~n2440 & n2663;
  assign n2666 = ~n2664 & ~n2665;
  assign n2667 = ~po49  & n2660;
  assign n2668 = ~n2666 & ~n2667;
  assign n2669 = ~n2661 & ~n2668;
  assign n2670 = po50  & ~n2669;
  assign n2671 = ~po50  & ~n2661;
  assign n2672 = ~n2668 & n2671;
  assign n2673 = ~n2443 & ~n2444;
  assign n2674 = po41  & n2673;
  assign n2675 = ~n2449 & ~n2674;
  assign n2676 = n2449 & n2674;
  assign n2677 = ~n2675 & ~n2676;
  assign n2678 = ~n2672 & n2677;
  assign n2679 = ~n2670 & ~n2678;
  assign n2680 = po51  & ~n2679;
  assign n2681 = ~n2452 & ~n2454;
  assign n2682 = po41  & n2681;
  assign n2683 = n2459 & ~n2682;
  assign n2684 = ~n2459 & n2682;
  assign n2685 = ~n2683 & ~n2684;
  assign n2686 = ~po51  & n2679;
  assign n2687 = ~n2685 & ~n2686;
  assign n2688 = ~n2680 & ~n2687;
  assign n2689 = po52  & ~n2688;
  assign n2690 = ~n2462 & ~n2463;
  assign n2691 = po41  & n2690;
  assign n2692 = n2468 & ~n2691;
  assign n2693 = ~n2468 & n2691;
  assign n2694 = ~n2692 & ~n2693;
  assign n2695 = ~po52  & ~n2680;
  assign n2696 = ~n2687 & n2695;
  assign n2697 = ~n2694 & ~n2696;
  assign n2698 = ~n2689 & ~n2697;
  assign n2699 = po53  & ~n2698;
  assign n2700 = ~n2471 & ~n2473;
  assign n2701 = po41  & n2700;
  assign n2702 = n2478 & ~n2701;
  assign n2703 = ~n2478 & n2701;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = ~po53  & n2698;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = ~n2699 & ~n2706;
  assign n2708 = po54  & ~n2707;
  assign n2709 = ~po54  & ~n2699;
  assign n2710 = ~n2706 & n2709;
  assign n2711 = ~n2481 & po41 ;
  assign n2712 = ~n2487 & n2711;
  assign n2713 = n2486 & ~n2712;
  assign n2714 = n2488 & n2711;
  assign n2715 = ~n2713 & ~n2714;
  assign n2716 = ~n2710 & n2715;
  assign n2717 = ~n2708 & ~n2716;
  assign n2718 = po55  & ~n2717;
  assign n2719 = ~n2490 & ~n2492;
  assign n2720 = po41  & n2719;
  assign n2721 = n2497 & ~n2720;
  assign n2722 = ~n2497 & n2720;
  assign n2723 = ~n2721 & ~n2722;
  assign n2724 = ~po55  & n2717;
  assign n2725 = ~n2723 & ~n2724;
  assign n2726 = ~n2718 & ~n2725;
  assign n2727 = po56  & ~n2726;
  assign n2728 = ~po56  & ~n2718;
  assign n2729 = ~n2725 & n2728;
  assign n2730 = ~n2500 & po41 ;
  assign n2731 = ~n2506 & n2730;
  assign n2732 = n2505 & ~n2731;
  assign n2733 = n2507 & n2730;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = ~n2729 & n2734;
  assign n2736 = ~n2727 & ~n2735;
  assign n2737 = po57  & ~n2736;
  assign n2738 = ~n2509 & ~n2511;
  assign n2739 = po41  & n2738;
  assign n2740 = n2516 & ~n2739;
  assign n2741 = ~n2516 & n2739;
  assign n2742 = ~n2740 & ~n2741;
  assign n2743 = ~po57  & n2736;
  assign n2744 = ~n2742 & ~n2743;
  assign n2745 = ~n2737 & ~n2744;
  assign n2746 = po58  & ~n2745;
  assign n2747 = ~po58  & ~n2737;
  assign n2748 = ~n2744 & n2747;
  assign n2749 = ~n2519 & po41 ;
  assign n2750 = ~n2525 & n2749;
  assign n2751 = n2524 & ~n2750;
  assign n2752 = n2526 & n2749;
  assign n2753 = ~n2751 & ~n2752;
  assign n2754 = ~n2748 & n2753;
  assign n2755 = ~n2746 & ~n2754;
  assign n2756 = po59  & ~n2755;
  assign n2757 = ~n2528 & ~n2530;
  assign n2758 = po41  & n2757;
  assign n2759 = n2535 & ~n2758;
  assign n2760 = ~n2535 & n2758;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = ~po59  & n2755;
  assign n2763 = ~n2761 & ~n2762;
  assign n2764 = ~n2756 & ~n2763;
  assign n2765 = po60  & ~n2764;
  assign n2766 = ~n2538 & ~n2539;
  assign n2767 = po41  & n2766;
  assign n2768 = n2544 & ~n2767;
  assign n2769 = ~n2544 & n2767;
  assign n2770 = ~n2768 & ~n2769;
  assign n2771 = ~po60  & ~n2756;
  assign n2772 = ~n2763 & n2771;
  assign n2773 = ~n2770 & ~n2772;
  assign n2774 = ~n2765 & ~n2773;
  assign n2775 = po61  & ~n2774;
  assign n2776 = ~n2547 & ~n2549;
  assign n2777 = po41  & n2776;
  assign n2778 = n2554 & ~n2777;
  assign n2779 = ~n2554 & n2777;
  assign n2780 = ~n2778 & ~n2779;
  assign n2781 = ~po61  & n2774;
  assign n2782 = ~n2780 & ~n2781;
  assign n2783 = ~n2775 & ~n2782;
  assign n2784 = po62  & ~n2783;
  assign n2785 = ~po62  & ~n2775;
  assign n2786 = ~n2782 & n2785;
  assign n2787 = ~n2557 & po41 ;
  assign n2788 = ~n2563 & n2787;
  assign n2789 = n2562 & ~n2788;
  assign n2790 = n2564 & n2787;
  assign n2791 = ~n2789 & ~n2790;
  assign n2792 = ~n2786 & n2791;
  assign n2793 = ~n2784 & ~n2792;
  assign n2794 = n2584 & po41 ;
  assign n2795 = ~n2575 & n2794;
  assign n2796 = ~n2566 & ~n2568;
  assign n2797 = po41  & n2796;
  assign n2798 = n2573 & ~n2797;
  assign n2799 = ~n2573 & n2797;
  assign n2800 = ~n2798 & ~n2799;
  assign n2801 = ~n2588 & ~n2795;
  assign n2802 = ~n2800 & n2801;
  assign n2803 = ~n2793 & n2802;
  assign n2804 = ~po63  & ~n2803;
  assign n2805 = n2793 & n2800;
  assign n2806 = n2575 & ~n2794;
  assign n2807 = ~n2575 & n2584;
  assign n2808 = po63  & ~n2807;
  assign n2809 = ~n2806 & n2808;
  assign n2810 = ~n2805 & ~n2809;
  assign po40  = n2804 | ~n2810;
  assign n2812 = pi80  & po40 ;
  assign n2813 = ~pi78  & ~pi79 ;
  assign n2814 = ~pi80  & n2813;
  assign n2815 = ~n2812 & ~n2814;
  assign n2816 = po41  & ~n2815;
  assign n2817 = ~pi80  & po40 ;
  assign n2818 = pi81  & ~n2817;
  assign n2819 = ~pi81  & n2817;
  assign n2820 = ~n2818 & ~n2819;
  assign n2821 = ~po41  & n2815;
  assign n2822 = n2820 & ~n2821;
  assign n2823 = ~n2816 & ~n2822;
  assign n2824 = po42  & ~n2823;
  assign n2825 = ~po42  & ~n2816;
  assign n2826 = ~n2822 & n2825;
  assign n2827 = po41  & ~po40 ;
  assign n2828 = ~n2819 & ~n2827;
  assign n2829 = pi82  & ~n2828;
  assign n2830 = ~pi82  & n2828;
  assign n2831 = ~n2829 & ~n2830;
  assign n2832 = ~n2826 & ~n2831;
  assign n2833 = ~n2824 & ~n2832;
  assign n2834 = po43  & ~n2833;
  assign n2835 = ~po43  & n2833;
  assign n2836 = ~n2596 & ~n2597;
  assign n2837 = po40  & n2836;
  assign n2838 = n2601 & ~n2837;
  assign n2839 = ~n2601 & n2837;
  assign n2840 = ~n2838 & ~n2839;
  assign n2841 = ~n2835 & ~n2840;
  assign n2842 = ~n2834 & ~n2841;
  assign n2843 = po44  & ~n2842;
  assign n2844 = ~po44  & ~n2834;
  assign n2845 = ~n2841 & n2844;
  assign n2846 = ~n2604 & po40 ;
  assign n2847 = ~n2610 & n2846;
  assign n2848 = n2609 & ~n2847;
  assign n2849 = n2611 & n2846;
  assign n2850 = ~n2848 & ~n2849;
  assign n2851 = ~n2845 & n2850;
  assign n2852 = ~n2843 & ~n2851;
  assign n2853 = po45  & ~n2852;
  assign n2854 = ~po45  & n2852;
  assign n2855 = ~n2613 & ~n2615;
  assign n2856 = po40  & n2855;
  assign n2857 = n2620 & ~n2856;
  assign n2858 = ~n2620 & n2856;
  assign n2859 = ~n2857 & ~n2858;
  assign n2860 = ~n2854 & n2859;
  assign n2861 = ~n2853 & ~n2860;
  assign n2862 = po46  & ~n2861;
  assign n2863 = ~po46  & ~n2853;
  assign n2864 = ~n2860 & n2863;
  assign n2865 = ~n2623 & po40 ;
  assign n2866 = ~n2629 & n2865;
  assign n2867 = n2628 & ~n2866;
  assign n2868 = n2630 & n2865;
  assign n2869 = ~n2867 & ~n2868;
  assign n2870 = ~n2864 & n2869;
  assign n2871 = ~n2862 & ~n2870;
  assign n2872 = po47  & ~n2871;
  assign n2873 = ~po47  & n2871;
  assign n2874 = ~n2632 & ~n2634;
  assign n2875 = po40  & n2874;
  assign n2876 = n2639 & n2875;
  assign n2877 = ~n2639 & ~n2875;
  assign n2878 = ~n2876 & ~n2877;
  assign n2879 = ~n2873 & n2878;
  assign n2880 = ~n2872 & ~n2879;
  assign n2881 = po48  & ~n2880;
  assign n2882 = ~po48  & ~n2872;
  assign n2883 = ~n2879 & n2882;
  assign n2884 = ~n2642 & po40 ;
  assign n2885 = ~n2648 & n2884;
  assign n2886 = n2647 & ~n2885;
  assign n2887 = n2649 & n2884;
  assign n2888 = ~n2886 & ~n2887;
  assign n2889 = ~n2883 & n2888;
  assign n2890 = ~n2881 & ~n2889;
  assign n2891 = po49  & ~n2890;
  assign n2892 = ~po49  & n2890;
  assign n2893 = ~n2651 & ~n2653;
  assign n2894 = po40  & n2893;
  assign n2895 = ~n2658 & ~n2894;
  assign n2896 = n2658 & n2894;
  assign n2897 = ~n2895 & ~n2896;
  assign n2898 = ~n2892 & n2897;
  assign n2899 = ~n2891 & ~n2898;
  assign n2900 = po50  & ~n2899;
  assign n2901 = ~po50  & ~n2891;
  assign n2902 = ~n2898 & n2901;
  assign n2903 = ~n2661 & po40 ;
  assign n2904 = ~n2667 & n2903;
  assign n2905 = n2666 & ~n2904;
  assign n2906 = n2668 & n2903;
  assign n2907 = ~n2905 & ~n2906;
  assign n2908 = ~n2902 & n2907;
  assign n2909 = ~n2900 & ~n2908;
  assign n2910 = po51  & ~n2909;
  assign n2911 = ~n2670 & ~n2672;
  assign n2912 = po40  & n2911;
  assign n2913 = n2677 & ~n2912;
  assign n2914 = ~n2677 & n2912;
  assign n2915 = ~n2913 & ~n2914;
  assign n2916 = ~po51  & n2909;
  assign n2917 = ~n2915 & ~n2916;
  assign n2918 = ~n2910 & ~n2917;
  assign n2919 = po52  & ~n2918;
  assign n2920 = ~po52  & ~n2910;
  assign n2921 = ~n2917 & n2920;
  assign n2922 = ~n2680 & po40 ;
  assign n2923 = ~n2686 & n2922;
  assign n2924 = n2685 & ~n2923;
  assign n2925 = n2687 & n2922;
  assign n2926 = ~n2924 & ~n2925;
  assign n2927 = ~n2921 & n2926;
  assign n2928 = ~n2919 & ~n2927;
  assign n2929 = po53  & ~n2928;
  assign n2930 = ~po53  & n2928;
  assign n2931 = ~n2689 & po40 ;
  assign n2932 = ~n2696 & n2931;
  assign n2933 = n2694 & ~n2932;
  assign n2934 = n2697 & n2931;
  assign n2935 = ~n2933 & ~n2934;
  assign n2936 = ~n2930 & n2935;
  assign n2937 = ~n2929 & ~n2936;
  assign n2938 = po54  & ~n2937;
  assign n2939 = ~po54  & ~n2929;
  assign n2940 = ~n2936 & n2939;
  assign n2941 = ~n2699 & po40 ;
  assign n2942 = ~n2705 & n2941;
  assign n2943 = n2704 & ~n2942;
  assign n2944 = n2706 & n2941;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = ~n2940 & n2945;
  assign n2947 = ~n2938 & ~n2946;
  assign n2948 = po55  & ~n2947;
  assign n2949 = ~n2708 & ~n2710;
  assign n2950 = po40  & n2949;
  assign n2951 = n2715 & ~n2950;
  assign n2952 = ~n2715 & n2950;
  assign n2953 = ~n2951 & ~n2952;
  assign n2954 = ~po55  & n2947;
  assign n2955 = ~n2953 & ~n2954;
  assign n2956 = ~n2948 & ~n2955;
  assign n2957 = po56  & ~n2956;
  assign n2958 = ~po56  & ~n2948;
  assign n2959 = ~n2955 & n2958;
  assign n2960 = ~n2718 & po40 ;
  assign n2961 = ~n2724 & n2960;
  assign n2962 = n2723 & ~n2961;
  assign n2963 = n2725 & n2960;
  assign n2964 = ~n2962 & ~n2963;
  assign n2965 = ~n2959 & n2964;
  assign n2966 = ~n2957 & ~n2965;
  assign n2967 = po57  & ~n2966;
  assign n2968 = ~n2727 & ~n2729;
  assign n2969 = po40  & n2968;
  assign n2970 = n2734 & ~n2969;
  assign n2971 = ~n2734 & n2969;
  assign n2972 = ~n2970 & ~n2971;
  assign n2973 = ~po57  & n2966;
  assign n2974 = ~n2972 & ~n2973;
  assign n2975 = ~n2967 & ~n2974;
  assign n2976 = po58  & ~n2975;
  assign n2977 = ~po58  & ~n2967;
  assign n2978 = ~n2974 & n2977;
  assign n2979 = ~n2737 & po40 ;
  assign n2980 = ~n2743 & n2979;
  assign n2981 = n2742 & ~n2980;
  assign n2982 = n2744 & n2979;
  assign n2983 = ~n2981 & ~n2982;
  assign n2984 = ~n2978 & n2983;
  assign n2985 = ~n2976 & ~n2984;
  assign n2986 = po59  & ~n2985;
  assign n2987 = ~n2746 & ~n2748;
  assign n2988 = po40  & n2987;
  assign n2989 = n2753 & ~n2988;
  assign n2990 = ~n2753 & n2988;
  assign n2991 = ~n2989 & ~n2990;
  assign n2992 = ~po59  & n2985;
  assign n2993 = ~n2991 & ~n2992;
  assign n2994 = ~n2986 & ~n2993;
  assign n2995 = po60  & ~n2994;
  assign n2996 = ~po60  & ~n2986;
  assign n2997 = ~n2993 & n2996;
  assign n2998 = ~n2756 & po40 ;
  assign n2999 = ~n2762 & n2998;
  assign n3000 = n2761 & ~n2999;
  assign n3001 = n2763 & n2998;
  assign n3002 = ~n3000 & ~n3001;
  assign n3003 = ~n2997 & n3002;
  assign n3004 = ~n2995 & ~n3003;
  assign n3005 = po61  & ~n3004;
  assign n3006 = ~po61  & n3004;
  assign n3007 = ~n2765 & po40 ;
  assign n3008 = ~n2772 & n3007;
  assign n3009 = n2770 & ~n3008;
  assign n3010 = n2773 & n3007;
  assign n3011 = ~n3009 & ~n3010;
  assign n3012 = ~n3006 & n3011;
  assign n3013 = ~n3005 & ~n3012;
  assign n3014 = po62  & ~n3013;
  assign n3015 = ~po62  & ~n3005;
  assign n3016 = ~n3012 & n3015;
  assign n3017 = ~n2775 & po40 ;
  assign n3018 = ~n2781 & n3017;
  assign n3019 = n2780 & ~n3018;
  assign n3020 = n2782 & n3017;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = ~n3016 & n3021;
  assign n3023 = ~n3014 & ~n3022;
  assign n3024 = ~n2784 & ~n2786;
  assign n3025 = po40  & n3024;
  assign n3026 = n2791 & ~n3025;
  assign n3027 = ~n2791 & n3025;
  assign n3028 = ~n3026 & ~n3027;
  assign n3029 = n2793 & po40 ;
  assign n3030 = ~n2800 & ~n3029;
  assign n3031 = ~n2805 & ~n3030;
  assign n3032 = po40  & ~n3031;
  assign n3033 = ~n3028 & ~n3032;
  assign n3034 = ~n3023 & n3033;
  assign n3035 = ~po63  & ~n3034;
  assign n3036 = n3023 & n3028;
  assign n3037 = po63  & n3031;
  assign n3038 = ~n3036 & ~n3037;
  assign po39  = n3035 | ~n3038;
  assign n3040 = pi78  & po39 ;
  assign n3041 = ~pi76  & ~pi77 ;
  assign n3042 = ~pi78  & n3041;
  assign n3043 = ~n3040 & ~n3042;
  assign n3044 = po40  & ~n3043;
  assign n3045 = ~po40  & n3043;
  assign n3046 = ~pi78  & po39 ;
  assign n3047 = pi79  & ~n3046;
  assign n3048 = ~pi79  & n3046;
  assign n3049 = ~n3047 & ~n3048;
  assign n3050 = ~n3045 & n3049;
  assign n3051 = ~n3044 & ~n3050;
  assign n3052 = po41  & ~n3051;
  assign n3053 = po40  & ~po39 ;
  assign n3054 = ~n3048 & ~n3053;
  assign n3055 = pi80  & ~n3054;
  assign n3056 = ~pi80  & n3054;
  assign n3057 = ~n3055 & ~n3056;
  assign n3058 = ~po41  & n3051;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = ~n3052 & ~n3059;
  assign n3061 = po42  & ~n3060;
  assign n3062 = ~po42  & ~n3052;
  assign n3063 = ~n3059 & n3062;
  assign n3064 = ~n2816 & ~n2821;
  assign n3065 = po39  & n3064;
  assign n3066 = n2820 & ~n3065;
  assign n3067 = ~n2820 & n3065;
  assign n3068 = ~n3066 & ~n3067;
  assign n3069 = ~n3063 & ~n3068;
  assign n3070 = ~n3061 & ~n3069;
  assign n3071 = po43  & ~n3070;
  assign n3072 = ~n2824 & ~n2826;
  assign n3073 = po39  & n3072;
  assign n3074 = ~n2831 & ~n3073;
  assign n3075 = n2831 & n3073;
  assign n3076 = ~n3074 & ~n3075;
  assign n3077 = ~po43  & n3070;
  assign n3078 = ~n3076 & ~n3077;
  assign n3079 = ~n3071 & ~n3078;
  assign n3080 = po44  & ~n3079;
  assign n3081 = ~po44  & ~n3071;
  assign n3082 = ~n3078 & n3081;
  assign n3083 = ~n2834 & ~n2835;
  assign n3084 = po39  & n3083;
  assign n3085 = n2840 & ~n3084;
  assign n3086 = ~n2840 & n3084;
  assign n3087 = ~n3085 & ~n3086;
  assign n3088 = ~n3082 & n3087;
  assign n3089 = ~n3080 & ~n3088;
  assign n3090 = po45  & ~n3089;
  assign n3091 = ~n2843 & ~n2845;
  assign n3092 = po39  & n3091;
  assign n3093 = n2850 & ~n3092;
  assign n3094 = ~n2850 & n3092;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = ~po45  & n3089;
  assign n3097 = ~n3095 & ~n3096;
  assign n3098 = ~n3090 & ~n3097;
  assign n3099 = po46  & ~n3098;
  assign n3100 = ~po46  & ~n3090;
  assign n3101 = ~n3097 & n3100;
  assign n3102 = ~n2853 & ~n2854;
  assign n3103 = po39  & n3102;
  assign n3104 = n2859 & n3103;
  assign n3105 = ~n2859 & ~n3103;
  assign n3106 = ~n3104 & ~n3105;
  assign n3107 = ~n3101 & n3106;
  assign n3108 = ~n3099 & ~n3107;
  assign n3109 = po47  & ~n3108;
  assign n3110 = ~n2862 & ~n2864;
  assign n3111 = po39  & n3110;
  assign n3112 = n2869 & ~n3111;
  assign n3113 = ~n2869 & n3111;
  assign n3114 = ~n3112 & ~n3113;
  assign n3115 = ~po47  & n3108;
  assign n3116 = ~n3114 & ~n3115;
  assign n3117 = ~n3109 & ~n3116;
  assign n3118 = po48  & ~n3117;
  assign n3119 = ~po48  & ~n3109;
  assign n3120 = ~n3116 & n3119;
  assign n3121 = ~n2872 & ~n2873;
  assign n3122 = po39  & n3121;
  assign n3123 = ~n2878 & ~n3122;
  assign n3124 = n2878 & n3122;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = ~n3120 & n3125;
  assign n3127 = ~n3118 & ~n3126;
  assign n3128 = po49  & ~n3127;
  assign n3129 = ~n2881 & ~n2883;
  assign n3130 = po39  & n3129;
  assign n3131 = n2888 & ~n3130;
  assign n3132 = ~n2888 & n3130;
  assign n3133 = ~n3131 & ~n3132;
  assign n3134 = ~po49  & n3127;
  assign n3135 = ~n3133 & ~n3134;
  assign n3136 = ~n3128 & ~n3135;
  assign n3137 = po50  & ~n3136;
  assign n3138 = ~n2891 & ~n2892;
  assign n3139 = po39  & n3138;
  assign n3140 = n2897 & ~n3139;
  assign n3141 = ~n2897 & n3139;
  assign n3142 = ~n3140 & ~n3141;
  assign n3143 = ~po50  & ~n3128;
  assign n3144 = ~n3135 & n3143;
  assign n3145 = ~n3142 & ~n3144;
  assign n3146 = ~n3137 & ~n3145;
  assign n3147 = po51  & ~n3146;
  assign n3148 = ~n2900 & ~n2902;
  assign n3149 = po39  & n3148;
  assign n3150 = n2907 & ~n3149;
  assign n3151 = ~n2907 & n3149;
  assign n3152 = ~n3150 & ~n3151;
  assign n3153 = ~po51  & n3146;
  assign n3154 = ~n3152 & ~n3153;
  assign n3155 = ~n3147 & ~n3154;
  assign n3156 = po52  & ~n3155;
  assign n3157 = ~po52  & ~n3147;
  assign n3158 = ~n3154 & n3157;
  assign n3159 = ~n2910 & po39 ;
  assign n3160 = ~n2916 & n3159;
  assign n3161 = n2915 & ~n3160;
  assign n3162 = n2917 & n3159;
  assign n3163 = ~n3161 & ~n3162;
  assign n3164 = ~n3158 & n3163;
  assign n3165 = ~n3156 & ~n3164;
  assign n3166 = po53  & ~n3165;
  assign n3167 = ~n2919 & ~n2921;
  assign n3168 = po39  & n3167;
  assign n3169 = n2926 & ~n3168;
  assign n3170 = ~n2926 & n3168;
  assign n3171 = ~n3169 & ~n3170;
  assign n3172 = ~po53  & n3165;
  assign n3173 = ~n3171 & ~n3172;
  assign n3174 = ~n3166 & ~n3173;
  assign n3175 = po54  & ~n3174;
  assign n3176 = ~n2929 & ~n2930;
  assign n3177 = po39  & n3176;
  assign n3178 = n2935 & ~n3177;
  assign n3179 = ~n2935 & n3177;
  assign n3180 = ~n3178 & ~n3179;
  assign n3181 = ~po54  & ~n3166;
  assign n3182 = ~n3173 & n3181;
  assign n3183 = ~n3180 & ~n3182;
  assign n3184 = ~n3175 & ~n3183;
  assign n3185 = po55  & ~n3184;
  assign n3186 = ~n2938 & ~n2940;
  assign n3187 = po39  & n3186;
  assign n3188 = n2945 & ~n3187;
  assign n3189 = ~n2945 & n3187;
  assign n3190 = ~n3188 & ~n3189;
  assign n3191 = ~po55  & n3184;
  assign n3192 = ~n3190 & ~n3191;
  assign n3193 = ~n3185 & ~n3192;
  assign n3194 = po56  & ~n3193;
  assign n3195 = ~po56  & ~n3185;
  assign n3196 = ~n3192 & n3195;
  assign n3197 = ~n2948 & po39 ;
  assign n3198 = ~n2954 & n3197;
  assign n3199 = n2953 & ~n3198;
  assign n3200 = n2955 & n3197;
  assign n3201 = ~n3199 & ~n3200;
  assign n3202 = ~n3196 & n3201;
  assign n3203 = ~n3194 & ~n3202;
  assign n3204 = po57  & ~n3203;
  assign n3205 = ~n2957 & ~n2959;
  assign n3206 = po39  & n3205;
  assign n3207 = n2964 & ~n3206;
  assign n3208 = ~n2964 & n3206;
  assign n3209 = ~n3207 & ~n3208;
  assign n3210 = ~po57  & n3203;
  assign n3211 = ~n3209 & ~n3210;
  assign n3212 = ~n3204 & ~n3211;
  assign n3213 = po58  & ~n3212;
  assign n3214 = ~po58  & ~n3204;
  assign n3215 = ~n3211 & n3214;
  assign n3216 = ~n2967 & po39 ;
  assign n3217 = ~n2973 & n3216;
  assign n3218 = n2972 & ~n3217;
  assign n3219 = n2974 & n3216;
  assign n3220 = ~n3218 & ~n3219;
  assign n3221 = ~n3215 & n3220;
  assign n3222 = ~n3213 & ~n3221;
  assign n3223 = po59  & ~n3222;
  assign n3224 = ~n2976 & ~n2978;
  assign n3225 = po39  & n3224;
  assign n3226 = n2983 & ~n3225;
  assign n3227 = ~n2983 & n3225;
  assign n3228 = ~n3226 & ~n3227;
  assign n3229 = ~po59  & n3222;
  assign n3230 = ~n3228 & ~n3229;
  assign n3231 = ~n3223 & ~n3230;
  assign n3232 = po60  & ~n3231;
  assign n3233 = ~po60  & ~n3223;
  assign n3234 = ~n3230 & n3233;
  assign n3235 = ~n2986 & po39 ;
  assign n3236 = ~n2992 & n3235;
  assign n3237 = n2991 & ~n3236;
  assign n3238 = n2993 & n3235;
  assign n3239 = ~n3237 & ~n3238;
  assign n3240 = ~n3234 & n3239;
  assign n3241 = ~n3232 & ~n3240;
  assign n3242 = po61  & ~n3241;
  assign n3243 = ~n2995 & ~n2997;
  assign n3244 = po39  & n3243;
  assign n3245 = n3002 & ~n3244;
  assign n3246 = ~n3002 & n3244;
  assign n3247 = ~n3245 & ~n3246;
  assign n3248 = ~po61  & n3241;
  assign n3249 = ~n3247 & ~n3248;
  assign n3250 = ~n3242 & ~n3249;
  assign n3251 = po62  & ~n3250;
  assign n3252 = ~n3005 & ~n3006;
  assign n3253 = po39  & n3252;
  assign n3254 = n3011 & ~n3253;
  assign n3255 = ~n3011 & n3253;
  assign n3256 = ~n3254 & ~n3255;
  assign n3257 = ~po62  & ~n3242;
  assign n3258 = ~n3249 & n3257;
  assign n3259 = ~n3256 & ~n3258;
  assign n3260 = ~n3251 & ~n3259;
  assign n3261 = ~n3014 & ~n3016;
  assign n3262 = po39  & n3261;
  assign n3263 = n3021 & ~n3262;
  assign n3264 = ~n3021 & n3262;
  assign n3265 = ~n3263 & ~n3264;
  assign n3266 = n3023 & po39 ;
  assign n3267 = ~n3028 & ~n3266;
  assign n3268 = ~n3036 & ~n3267;
  assign n3269 = po39  & ~n3268;
  assign n3270 = ~n3265 & ~n3269;
  assign n3271 = ~n3260 & n3270;
  assign n3272 = ~po63  & ~n3271;
  assign n3273 = n3260 & n3265;
  assign n3274 = po63  & n3268;
  assign n3275 = ~n3273 & ~n3274;
  assign po38  = n3272 | ~n3275;
  assign n3277 = pi76  & po38 ;
  assign n3278 = ~pi74  & ~pi75 ;
  assign n3279 = ~pi76  & n3278;
  assign n3280 = ~n3277 & ~n3279;
  assign n3281 = po39  & ~n3280;
  assign n3282 = ~pi76  & po38 ;
  assign n3283 = pi77  & ~n3282;
  assign n3284 = ~pi77  & n3282;
  assign n3285 = ~n3283 & ~n3284;
  assign n3286 = ~po39  & n3280;
  assign n3287 = n3285 & ~n3286;
  assign n3288 = ~n3281 & ~n3287;
  assign n3289 = po40  & ~n3288;
  assign n3290 = ~po40  & ~n3281;
  assign n3291 = ~n3287 & n3290;
  assign n3292 = po39  & ~po38 ;
  assign n3293 = ~n3284 & ~n3292;
  assign n3294 = pi78  & ~n3293;
  assign n3295 = ~pi78  & n3293;
  assign n3296 = ~n3294 & ~n3295;
  assign n3297 = ~n3291 & ~n3296;
  assign n3298 = ~n3289 & ~n3297;
  assign n3299 = po41  & ~n3298;
  assign n3300 = ~po41  & n3298;
  assign n3301 = ~n3044 & ~n3045;
  assign n3302 = po38  & n3301;
  assign n3303 = n3049 & ~n3302;
  assign n3304 = ~n3049 & n3302;
  assign n3305 = ~n3303 & ~n3304;
  assign n3306 = ~n3300 & ~n3305;
  assign n3307 = ~n3299 & ~n3306;
  assign n3308 = po42  & ~n3307;
  assign n3309 = ~po42  & ~n3299;
  assign n3310 = ~n3306 & n3309;
  assign n3311 = ~n3052 & po38 ;
  assign n3312 = ~n3058 & n3311;
  assign n3313 = n3057 & ~n3312;
  assign n3314 = n3059 & n3311;
  assign n3315 = ~n3313 & ~n3314;
  assign n3316 = ~n3310 & n3315;
  assign n3317 = ~n3308 & ~n3316;
  assign n3318 = po43  & ~n3317;
  assign n3319 = ~po43  & n3317;
  assign n3320 = ~n3061 & ~n3063;
  assign n3321 = po38  & n3320;
  assign n3322 = n3068 & ~n3321;
  assign n3323 = ~n3068 & n3321;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = ~n3319 & n3324;
  assign n3326 = ~n3318 & ~n3325;
  assign n3327 = po44  & ~n3326;
  assign n3328 = ~po44  & ~n3318;
  assign n3329 = ~n3325 & n3328;
  assign n3330 = ~n3071 & po38 ;
  assign n3331 = ~n3077 & n3330;
  assign n3332 = n3076 & ~n3331;
  assign n3333 = n3078 & n3330;
  assign n3334 = ~n3332 & ~n3333;
  assign n3335 = ~n3329 & n3334;
  assign n3336 = ~n3327 & ~n3335;
  assign n3337 = po45  & ~n3336;
  assign n3338 = ~po45  & n3336;
  assign n3339 = ~n3080 & ~n3082;
  assign n3340 = po38  & n3339;
  assign n3341 = n3087 & n3340;
  assign n3342 = ~n3087 & ~n3340;
  assign n3343 = ~n3341 & ~n3342;
  assign n3344 = ~n3338 & n3343;
  assign n3345 = ~n3337 & ~n3344;
  assign n3346 = po46  & ~n3345;
  assign n3347 = ~po46  & ~n3337;
  assign n3348 = ~n3344 & n3347;
  assign n3349 = ~n3090 & po38 ;
  assign n3350 = ~n3096 & n3349;
  assign n3351 = n3095 & ~n3350;
  assign n3352 = n3097 & n3349;
  assign n3353 = ~n3351 & ~n3352;
  assign n3354 = ~n3348 & n3353;
  assign n3355 = ~n3346 & ~n3354;
  assign n3356 = po47  & ~n3355;
  assign n3357 = ~po47  & n3355;
  assign n3358 = ~n3099 & ~n3101;
  assign n3359 = po38  & n3358;
  assign n3360 = ~n3106 & ~n3359;
  assign n3361 = n3106 & n3359;
  assign n3362 = ~n3360 & ~n3361;
  assign n3363 = ~n3357 & n3362;
  assign n3364 = ~n3356 & ~n3363;
  assign n3365 = po48  & ~n3364;
  assign n3366 = ~po48  & ~n3356;
  assign n3367 = ~n3363 & n3366;
  assign n3368 = ~n3109 & po38 ;
  assign n3369 = ~n3115 & n3368;
  assign n3370 = n3114 & ~n3369;
  assign n3371 = n3116 & n3368;
  assign n3372 = ~n3370 & ~n3371;
  assign n3373 = ~n3367 & n3372;
  assign n3374 = ~n3365 & ~n3373;
  assign n3375 = po49  & ~n3374;
  assign n3376 = ~n3118 & ~n3120;
  assign n3377 = po38  & n3376;
  assign n3378 = n3125 & ~n3377;
  assign n3379 = ~n3125 & n3377;
  assign n3380 = ~n3378 & ~n3379;
  assign n3381 = ~po49  & n3374;
  assign n3382 = ~n3380 & ~n3381;
  assign n3383 = ~n3375 & ~n3382;
  assign n3384 = po50  & ~n3383;
  assign n3385 = ~po50  & ~n3375;
  assign n3386 = ~n3382 & n3385;
  assign n3387 = ~n3128 & po38 ;
  assign n3388 = ~n3134 & n3387;
  assign n3389 = n3133 & ~n3388;
  assign n3390 = n3135 & n3387;
  assign n3391 = ~n3389 & ~n3390;
  assign n3392 = ~n3386 & n3391;
  assign n3393 = ~n3384 & ~n3392;
  assign n3394 = po51  & ~n3393;
  assign n3395 = ~po51  & n3393;
  assign n3396 = ~n3137 & po38 ;
  assign n3397 = ~n3144 & n3396;
  assign n3398 = n3142 & ~n3397;
  assign n3399 = n3145 & n3396;
  assign n3400 = ~n3398 & ~n3399;
  assign n3401 = ~n3395 & n3400;
  assign n3402 = ~n3394 & ~n3401;
  assign n3403 = po52  & ~n3402;
  assign n3404 = ~po52  & ~n3394;
  assign n3405 = ~n3401 & n3404;
  assign n3406 = ~n3147 & po38 ;
  assign n3407 = ~n3153 & n3406;
  assign n3408 = n3152 & ~n3407;
  assign n3409 = n3154 & n3406;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = ~n3405 & n3410;
  assign n3412 = ~n3403 & ~n3411;
  assign n3413 = po53  & ~n3412;
  assign n3414 = ~n3156 & ~n3158;
  assign n3415 = po38  & n3414;
  assign n3416 = n3163 & ~n3415;
  assign n3417 = ~n3163 & n3415;
  assign n3418 = ~n3416 & ~n3417;
  assign n3419 = ~po53  & n3412;
  assign n3420 = ~n3418 & ~n3419;
  assign n3421 = ~n3413 & ~n3420;
  assign n3422 = po54  & ~n3421;
  assign n3423 = ~po54  & ~n3413;
  assign n3424 = ~n3420 & n3423;
  assign n3425 = ~n3166 & po38 ;
  assign n3426 = ~n3172 & n3425;
  assign n3427 = n3171 & ~n3426;
  assign n3428 = n3173 & n3425;
  assign n3429 = ~n3427 & ~n3428;
  assign n3430 = ~n3424 & n3429;
  assign n3431 = ~n3422 & ~n3430;
  assign n3432 = po55  & ~n3431;
  assign n3433 = ~po55  & n3431;
  assign n3434 = ~n3175 & po38 ;
  assign n3435 = ~n3182 & n3434;
  assign n3436 = n3180 & ~n3435;
  assign n3437 = n3183 & n3434;
  assign n3438 = ~n3436 & ~n3437;
  assign n3439 = ~n3433 & n3438;
  assign n3440 = ~n3432 & ~n3439;
  assign n3441 = po56  & ~n3440;
  assign n3442 = ~po56  & ~n3432;
  assign n3443 = ~n3439 & n3442;
  assign n3444 = ~n3185 & po38 ;
  assign n3445 = ~n3191 & n3444;
  assign n3446 = n3190 & ~n3445;
  assign n3447 = n3192 & n3444;
  assign n3448 = ~n3446 & ~n3447;
  assign n3449 = ~n3443 & n3448;
  assign n3450 = ~n3441 & ~n3449;
  assign n3451 = po57  & ~n3450;
  assign n3452 = ~n3194 & ~n3196;
  assign n3453 = po38  & n3452;
  assign n3454 = n3201 & ~n3453;
  assign n3455 = ~n3201 & n3453;
  assign n3456 = ~n3454 & ~n3455;
  assign n3457 = ~po57  & n3450;
  assign n3458 = ~n3456 & ~n3457;
  assign n3459 = ~n3451 & ~n3458;
  assign n3460 = po58  & ~n3459;
  assign n3461 = ~po58  & ~n3451;
  assign n3462 = ~n3458 & n3461;
  assign n3463 = ~n3204 & po38 ;
  assign n3464 = ~n3210 & n3463;
  assign n3465 = n3209 & ~n3464;
  assign n3466 = n3211 & n3463;
  assign n3467 = ~n3465 & ~n3466;
  assign n3468 = ~n3462 & n3467;
  assign n3469 = ~n3460 & ~n3468;
  assign n3470 = po59  & ~n3469;
  assign n3471 = ~n3213 & ~n3215;
  assign n3472 = po38  & n3471;
  assign n3473 = n3220 & ~n3472;
  assign n3474 = ~n3220 & n3472;
  assign n3475 = ~n3473 & ~n3474;
  assign n3476 = ~po59  & n3469;
  assign n3477 = ~n3475 & ~n3476;
  assign n3478 = ~n3470 & ~n3477;
  assign n3479 = po60  & ~n3478;
  assign n3480 = ~po60  & ~n3470;
  assign n3481 = ~n3477 & n3480;
  assign n3482 = ~n3223 & po38 ;
  assign n3483 = ~n3229 & n3482;
  assign n3484 = n3228 & ~n3483;
  assign n3485 = n3230 & n3482;
  assign n3486 = ~n3484 & ~n3485;
  assign n3487 = ~n3481 & n3486;
  assign n3488 = ~n3479 & ~n3487;
  assign n3489 = po61  & ~n3488;
  assign n3490 = ~n3232 & ~n3234;
  assign n3491 = po38  & n3490;
  assign n3492 = n3239 & ~n3491;
  assign n3493 = ~n3239 & n3491;
  assign n3494 = ~n3492 & ~n3493;
  assign n3495 = ~po61  & n3488;
  assign n3496 = ~n3494 & ~n3495;
  assign n3497 = ~n3489 & ~n3496;
  assign n3498 = po62  & ~n3497;
  assign n3499 = ~po62  & ~n3489;
  assign n3500 = ~n3496 & n3499;
  assign n3501 = ~n3242 & po38 ;
  assign n3502 = ~n3248 & n3501;
  assign n3503 = n3247 & ~n3502;
  assign n3504 = n3249 & n3501;
  assign n3505 = ~n3503 & ~n3504;
  assign n3506 = ~n3500 & n3505;
  assign n3507 = ~n3498 & ~n3506;
  assign n3508 = n3260 & po38 ;
  assign n3509 = ~n3265 & ~n3508;
  assign n3510 = ~n3273 & ~n3509;
  assign n3511 = po38  & ~n3510;
  assign n3512 = ~n3251 & po38 ;
  assign n3513 = ~n3258 & n3512;
  assign n3514 = n3256 & ~n3513;
  assign n3515 = n3259 & n3512;
  assign n3516 = ~n3514 & ~n3515;
  assign n3517 = ~n3511 & n3516;
  assign n3518 = ~n3507 & n3517;
  assign n3519 = ~po63  & ~n3518;
  assign n3520 = n3507 & ~n3516;
  assign n3521 = po63  & n3510;
  assign n3522 = ~n3520 & ~n3521;
  assign po37  = n3519 | ~n3522;
  assign n3524 = pi74  & po37 ;
  assign n3525 = ~pi72  & ~pi73 ;
  assign n3526 = ~pi74  & n3525;
  assign n3527 = ~n3524 & ~n3526;
  assign n3528 = po38  & ~n3527;
  assign n3529 = ~po38  & n3527;
  assign n3530 = ~pi74  & po37 ;
  assign n3531 = pi75  & ~n3530;
  assign n3532 = ~pi75  & n3530;
  assign n3533 = ~n3531 & ~n3532;
  assign n3534 = ~n3529 & n3533;
  assign n3535 = ~n3528 & ~n3534;
  assign n3536 = po39  & ~n3535;
  assign n3537 = po38  & ~po37 ;
  assign n3538 = ~n3532 & ~n3537;
  assign n3539 = pi76  & ~n3538;
  assign n3540 = ~pi76  & n3538;
  assign n3541 = ~n3539 & ~n3540;
  assign n3542 = ~po39  & n3535;
  assign n3543 = ~n3541 & ~n3542;
  assign n3544 = ~n3536 & ~n3543;
  assign n3545 = po40  & ~n3544;
  assign n3546 = ~po40  & ~n3536;
  assign n3547 = ~n3543 & n3546;
  assign n3548 = ~n3281 & ~n3286;
  assign n3549 = po37  & n3548;
  assign n3550 = n3285 & ~n3549;
  assign n3551 = ~n3285 & n3549;
  assign n3552 = ~n3550 & ~n3551;
  assign n3553 = ~n3547 & ~n3552;
  assign n3554 = ~n3545 & ~n3553;
  assign n3555 = po41  & ~n3554;
  assign n3556 = ~n3289 & ~n3291;
  assign n3557 = po37  & n3556;
  assign n3558 = ~n3296 & ~n3557;
  assign n3559 = n3296 & n3557;
  assign n3560 = ~n3558 & ~n3559;
  assign n3561 = ~po41  & n3554;
  assign n3562 = ~n3560 & ~n3561;
  assign n3563 = ~n3555 & ~n3562;
  assign n3564 = po42  & ~n3563;
  assign n3565 = ~po42  & ~n3555;
  assign n3566 = ~n3562 & n3565;
  assign n3567 = ~n3299 & ~n3300;
  assign n3568 = po37  & n3567;
  assign n3569 = n3305 & ~n3568;
  assign n3570 = ~n3305 & n3568;
  assign n3571 = ~n3569 & ~n3570;
  assign n3572 = ~n3566 & n3571;
  assign n3573 = ~n3564 & ~n3572;
  assign n3574 = po43  & ~n3573;
  assign n3575 = ~n3308 & ~n3310;
  assign n3576 = po37  & n3575;
  assign n3577 = n3315 & ~n3576;
  assign n3578 = ~n3315 & n3576;
  assign n3579 = ~n3577 & ~n3578;
  assign n3580 = ~po43  & n3573;
  assign n3581 = ~n3579 & ~n3580;
  assign n3582 = ~n3574 & ~n3581;
  assign n3583 = po44  & ~n3582;
  assign n3584 = ~po44  & ~n3574;
  assign n3585 = ~n3581 & n3584;
  assign n3586 = ~n3318 & ~n3319;
  assign n3587 = po37  & n3586;
  assign n3588 = n3324 & n3587;
  assign n3589 = ~n3324 & ~n3587;
  assign n3590 = ~n3588 & ~n3589;
  assign n3591 = ~n3585 & n3590;
  assign n3592 = ~n3583 & ~n3591;
  assign n3593 = po45  & ~n3592;
  assign n3594 = ~n3327 & ~n3329;
  assign n3595 = po37  & n3594;
  assign n3596 = n3334 & ~n3595;
  assign n3597 = ~n3334 & n3595;
  assign n3598 = ~n3596 & ~n3597;
  assign n3599 = ~po45  & n3592;
  assign n3600 = ~n3598 & ~n3599;
  assign n3601 = ~n3593 & ~n3600;
  assign n3602 = po46  & ~n3601;
  assign n3603 = ~po46  & ~n3593;
  assign n3604 = ~n3600 & n3603;
  assign n3605 = ~n3337 & ~n3338;
  assign n3606 = po37  & n3605;
  assign n3607 = ~n3343 & ~n3606;
  assign n3608 = n3343 & n3606;
  assign n3609 = ~n3607 & ~n3608;
  assign n3610 = ~n3604 & n3609;
  assign n3611 = ~n3602 & ~n3610;
  assign n3612 = po47  & ~n3611;
  assign n3613 = ~n3346 & ~n3348;
  assign n3614 = po37  & n3613;
  assign n3615 = n3353 & ~n3614;
  assign n3616 = ~n3353 & n3614;
  assign n3617 = ~n3615 & ~n3616;
  assign n3618 = ~po47  & n3611;
  assign n3619 = ~n3617 & ~n3618;
  assign n3620 = ~n3612 & ~n3619;
  assign n3621 = po48  & ~n3620;
  assign n3622 = ~n3356 & ~n3357;
  assign n3623 = po37  & n3622;
  assign n3624 = n3362 & ~n3623;
  assign n3625 = ~n3362 & n3623;
  assign n3626 = ~n3624 & ~n3625;
  assign n3627 = ~po48  & ~n3612;
  assign n3628 = ~n3619 & n3627;
  assign n3629 = ~n3626 & ~n3628;
  assign n3630 = ~n3621 & ~n3629;
  assign n3631 = po49  & ~n3630;
  assign n3632 = ~n3365 & ~n3367;
  assign n3633 = po37  & n3632;
  assign n3634 = n3372 & ~n3633;
  assign n3635 = ~n3372 & n3633;
  assign n3636 = ~n3634 & ~n3635;
  assign n3637 = ~po49  & n3630;
  assign n3638 = ~n3636 & ~n3637;
  assign n3639 = ~n3631 & ~n3638;
  assign n3640 = po50  & ~n3639;
  assign n3641 = ~po50  & ~n3631;
  assign n3642 = ~n3638 & n3641;
  assign n3643 = ~n3375 & po37 ;
  assign n3644 = ~n3381 & n3643;
  assign n3645 = n3380 & ~n3644;
  assign n3646 = n3382 & n3643;
  assign n3647 = ~n3645 & ~n3646;
  assign n3648 = ~n3642 & n3647;
  assign n3649 = ~n3640 & ~n3648;
  assign n3650 = po51  & ~n3649;
  assign n3651 = ~n3384 & ~n3386;
  assign n3652 = po37  & n3651;
  assign n3653 = n3391 & ~n3652;
  assign n3654 = ~n3391 & n3652;
  assign n3655 = ~n3653 & ~n3654;
  assign n3656 = ~po51  & n3649;
  assign n3657 = ~n3655 & ~n3656;
  assign n3658 = ~n3650 & ~n3657;
  assign n3659 = po52  & ~n3658;
  assign n3660 = ~n3394 & ~n3395;
  assign n3661 = po37  & n3660;
  assign n3662 = n3400 & ~n3661;
  assign n3663 = ~n3400 & n3661;
  assign n3664 = ~n3662 & ~n3663;
  assign n3665 = ~po52  & ~n3650;
  assign n3666 = ~n3657 & n3665;
  assign n3667 = ~n3664 & ~n3666;
  assign n3668 = ~n3659 & ~n3667;
  assign n3669 = po53  & ~n3668;
  assign n3670 = ~n3403 & ~n3405;
  assign n3671 = po37  & n3670;
  assign n3672 = n3410 & ~n3671;
  assign n3673 = ~n3410 & n3671;
  assign n3674 = ~n3672 & ~n3673;
  assign n3675 = ~po53  & n3668;
  assign n3676 = ~n3674 & ~n3675;
  assign n3677 = ~n3669 & ~n3676;
  assign n3678 = po54  & ~n3677;
  assign n3679 = ~po54  & ~n3669;
  assign n3680 = ~n3676 & n3679;
  assign n3681 = ~n3413 & po37 ;
  assign n3682 = ~n3419 & n3681;
  assign n3683 = n3418 & ~n3682;
  assign n3684 = n3420 & n3681;
  assign n3685 = ~n3683 & ~n3684;
  assign n3686 = ~n3680 & n3685;
  assign n3687 = ~n3678 & ~n3686;
  assign n3688 = po55  & ~n3687;
  assign n3689 = ~n3422 & ~n3424;
  assign n3690 = po37  & n3689;
  assign n3691 = n3429 & ~n3690;
  assign n3692 = ~n3429 & n3690;
  assign n3693 = ~n3691 & ~n3692;
  assign n3694 = ~po55  & n3687;
  assign n3695 = ~n3693 & ~n3694;
  assign n3696 = ~n3688 & ~n3695;
  assign n3697 = po56  & ~n3696;
  assign n3698 = ~n3432 & ~n3433;
  assign n3699 = po37  & n3698;
  assign n3700 = n3438 & ~n3699;
  assign n3701 = ~n3438 & n3699;
  assign n3702 = ~n3700 & ~n3701;
  assign n3703 = ~po56  & ~n3688;
  assign n3704 = ~n3695 & n3703;
  assign n3705 = ~n3702 & ~n3704;
  assign n3706 = ~n3697 & ~n3705;
  assign n3707 = po57  & ~n3706;
  assign n3708 = ~n3441 & ~n3443;
  assign n3709 = po37  & n3708;
  assign n3710 = n3448 & ~n3709;
  assign n3711 = ~n3448 & n3709;
  assign n3712 = ~n3710 & ~n3711;
  assign n3713 = ~po57  & n3706;
  assign n3714 = ~n3712 & ~n3713;
  assign n3715 = ~n3707 & ~n3714;
  assign n3716 = po58  & ~n3715;
  assign n3717 = ~po58  & ~n3707;
  assign n3718 = ~n3714 & n3717;
  assign n3719 = ~n3451 & po37 ;
  assign n3720 = ~n3457 & n3719;
  assign n3721 = n3456 & ~n3720;
  assign n3722 = n3458 & n3719;
  assign n3723 = ~n3721 & ~n3722;
  assign n3724 = ~n3718 & n3723;
  assign n3725 = ~n3716 & ~n3724;
  assign n3726 = po59  & ~n3725;
  assign n3727 = ~n3460 & ~n3462;
  assign n3728 = po37  & n3727;
  assign n3729 = n3467 & ~n3728;
  assign n3730 = ~n3467 & n3728;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = ~po59  & n3725;
  assign n3733 = ~n3731 & ~n3732;
  assign n3734 = ~n3726 & ~n3733;
  assign n3735 = po60  & ~n3734;
  assign n3736 = ~po60  & ~n3726;
  assign n3737 = ~n3733 & n3736;
  assign n3738 = ~n3470 & po37 ;
  assign n3739 = ~n3476 & n3738;
  assign n3740 = n3475 & ~n3739;
  assign n3741 = n3477 & n3738;
  assign n3742 = ~n3740 & ~n3741;
  assign n3743 = ~n3737 & n3742;
  assign n3744 = ~n3735 & ~n3743;
  assign n3745 = po61  & ~n3744;
  assign n3746 = ~n3479 & ~n3481;
  assign n3747 = po37  & n3746;
  assign n3748 = n3486 & ~n3747;
  assign n3749 = ~n3486 & n3747;
  assign n3750 = ~n3748 & ~n3749;
  assign n3751 = ~po61  & n3744;
  assign n3752 = ~n3750 & ~n3751;
  assign n3753 = ~n3745 & ~n3752;
  assign n3754 = po62  & ~n3753;
  assign n3755 = ~po62  & ~n3745;
  assign n3756 = ~n3752 & n3755;
  assign n3757 = ~n3489 & po37 ;
  assign n3758 = ~n3495 & n3757;
  assign n3759 = n3494 & ~n3758;
  assign n3760 = n3496 & n3757;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = ~n3756 & n3761;
  assign n3763 = ~n3754 & ~n3762;
  assign n3764 = n3516 & po37 ;
  assign n3765 = ~n3507 & n3764;
  assign n3766 = ~n3498 & ~n3500;
  assign n3767 = po37  & n3766;
  assign n3768 = n3505 & ~n3767;
  assign n3769 = ~n3505 & n3767;
  assign n3770 = ~n3768 & ~n3769;
  assign n3771 = ~n3520 & ~n3765;
  assign n3772 = ~n3770 & n3771;
  assign n3773 = ~n3763 & n3772;
  assign n3774 = ~po63  & ~n3773;
  assign n3775 = n3763 & n3770;
  assign n3776 = n3507 & ~n3764;
  assign n3777 = ~n3507 & n3516;
  assign n3778 = po63  & ~n3777;
  assign n3779 = ~n3776 & n3778;
  assign n3780 = ~n3775 & ~n3779;
  assign po36  = n3774 | ~n3780;
  assign n3782 = pi72  & po36 ;
  assign n3783 = ~pi70  & ~pi71 ;
  assign n3784 = ~pi72  & n3783;
  assign n3785 = ~n3782 & ~n3784;
  assign n3786 = po37  & ~n3785;
  assign n3787 = ~pi72  & po36 ;
  assign n3788 = pi73  & ~n3787;
  assign n3789 = ~pi73  & n3787;
  assign n3790 = ~n3788 & ~n3789;
  assign n3791 = ~po37  & n3785;
  assign n3792 = n3790 & ~n3791;
  assign n3793 = ~n3786 & ~n3792;
  assign n3794 = po38  & ~n3793;
  assign n3795 = ~po38  & ~n3786;
  assign n3796 = ~n3792 & n3795;
  assign n3797 = po37  & ~po36 ;
  assign n3798 = ~n3789 & ~n3797;
  assign n3799 = pi74  & ~n3798;
  assign n3800 = ~pi74  & n3798;
  assign n3801 = ~n3799 & ~n3800;
  assign n3802 = ~n3796 & ~n3801;
  assign n3803 = ~n3794 & ~n3802;
  assign n3804 = po39  & ~n3803;
  assign n3805 = ~po39  & n3803;
  assign n3806 = ~n3528 & ~n3529;
  assign n3807 = po36  & n3806;
  assign n3808 = n3533 & ~n3807;
  assign n3809 = ~n3533 & n3807;
  assign n3810 = ~n3808 & ~n3809;
  assign n3811 = ~n3805 & ~n3810;
  assign n3812 = ~n3804 & ~n3811;
  assign n3813 = po40  & ~n3812;
  assign n3814 = ~po40  & ~n3804;
  assign n3815 = ~n3811 & n3814;
  assign n3816 = ~n3536 & po36 ;
  assign n3817 = ~n3542 & n3816;
  assign n3818 = n3541 & ~n3817;
  assign n3819 = n3543 & n3816;
  assign n3820 = ~n3818 & ~n3819;
  assign n3821 = ~n3815 & n3820;
  assign n3822 = ~n3813 & ~n3821;
  assign n3823 = po41  & ~n3822;
  assign n3824 = ~po41  & n3822;
  assign n3825 = ~n3545 & ~n3547;
  assign n3826 = po36  & n3825;
  assign n3827 = n3552 & ~n3826;
  assign n3828 = ~n3552 & n3826;
  assign n3829 = ~n3827 & ~n3828;
  assign n3830 = ~n3824 & n3829;
  assign n3831 = ~n3823 & ~n3830;
  assign n3832 = po42  & ~n3831;
  assign n3833 = ~po42  & ~n3823;
  assign n3834 = ~n3830 & n3833;
  assign n3835 = ~n3555 & po36 ;
  assign n3836 = ~n3561 & n3835;
  assign n3837 = n3560 & ~n3836;
  assign n3838 = n3562 & n3835;
  assign n3839 = ~n3837 & ~n3838;
  assign n3840 = ~n3834 & n3839;
  assign n3841 = ~n3832 & ~n3840;
  assign n3842 = po43  & ~n3841;
  assign n3843 = ~po43  & n3841;
  assign n3844 = ~n3564 & ~n3566;
  assign n3845 = po36  & n3844;
  assign n3846 = n3571 & n3845;
  assign n3847 = ~n3571 & ~n3845;
  assign n3848 = ~n3846 & ~n3847;
  assign n3849 = ~n3843 & n3848;
  assign n3850 = ~n3842 & ~n3849;
  assign n3851 = po44  & ~n3850;
  assign n3852 = ~po44  & ~n3842;
  assign n3853 = ~n3849 & n3852;
  assign n3854 = ~n3574 & po36 ;
  assign n3855 = ~n3580 & n3854;
  assign n3856 = n3579 & ~n3855;
  assign n3857 = n3581 & n3854;
  assign n3858 = ~n3856 & ~n3857;
  assign n3859 = ~n3853 & n3858;
  assign n3860 = ~n3851 & ~n3859;
  assign n3861 = po45  & ~n3860;
  assign n3862 = ~po45  & n3860;
  assign n3863 = ~n3583 & ~n3585;
  assign n3864 = po36  & n3863;
  assign n3865 = ~n3590 & ~n3864;
  assign n3866 = n3590 & n3864;
  assign n3867 = ~n3865 & ~n3866;
  assign n3868 = ~n3862 & n3867;
  assign n3869 = ~n3861 & ~n3868;
  assign n3870 = po46  & ~n3869;
  assign n3871 = ~po46  & ~n3861;
  assign n3872 = ~n3868 & n3871;
  assign n3873 = ~n3593 & po36 ;
  assign n3874 = ~n3599 & n3873;
  assign n3875 = n3598 & ~n3874;
  assign n3876 = n3600 & n3873;
  assign n3877 = ~n3875 & ~n3876;
  assign n3878 = ~n3872 & n3877;
  assign n3879 = ~n3870 & ~n3878;
  assign n3880 = po47  & ~n3879;
  assign n3881 = ~n3602 & ~n3604;
  assign n3882 = po36  & n3881;
  assign n3883 = n3609 & ~n3882;
  assign n3884 = ~n3609 & n3882;
  assign n3885 = ~n3883 & ~n3884;
  assign n3886 = ~po47  & n3879;
  assign n3887 = ~n3885 & ~n3886;
  assign n3888 = ~n3880 & ~n3887;
  assign n3889 = po48  & ~n3888;
  assign n3890 = ~po48  & ~n3880;
  assign n3891 = ~n3887 & n3890;
  assign n3892 = ~n3612 & po36 ;
  assign n3893 = ~n3618 & n3892;
  assign n3894 = n3617 & ~n3893;
  assign n3895 = n3619 & n3892;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = ~n3891 & n3896;
  assign n3898 = ~n3889 & ~n3897;
  assign n3899 = po49  & ~n3898;
  assign n3900 = ~po49  & n3898;
  assign n3901 = ~n3621 & po36 ;
  assign n3902 = ~n3628 & n3901;
  assign n3903 = n3626 & ~n3902;
  assign n3904 = n3629 & n3901;
  assign n3905 = ~n3903 & ~n3904;
  assign n3906 = ~n3900 & n3905;
  assign n3907 = ~n3899 & ~n3906;
  assign n3908 = po50  & ~n3907;
  assign n3909 = ~po50  & ~n3899;
  assign n3910 = ~n3906 & n3909;
  assign n3911 = ~n3631 & po36 ;
  assign n3912 = ~n3637 & n3911;
  assign n3913 = n3636 & ~n3912;
  assign n3914 = n3638 & n3911;
  assign n3915 = ~n3913 & ~n3914;
  assign n3916 = ~n3910 & n3915;
  assign n3917 = ~n3908 & ~n3916;
  assign n3918 = po51  & ~n3917;
  assign n3919 = ~n3640 & ~n3642;
  assign n3920 = po36  & n3919;
  assign n3921 = n3647 & ~n3920;
  assign n3922 = ~n3647 & n3920;
  assign n3923 = ~n3921 & ~n3922;
  assign n3924 = ~po51  & n3917;
  assign n3925 = ~n3923 & ~n3924;
  assign n3926 = ~n3918 & ~n3925;
  assign n3927 = po52  & ~n3926;
  assign n3928 = ~po52  & ~n3918;
  assign n3929 = ~n3925 & n3928;
  assign n3930 = ~n3650 & po36 ;
  assign n3931 = ~n3656 & n3930;
  assign n3932 = n3655 & ~n3931;
  assign n3933 = n3657 & n3930;
  assign n3934 = ~n3932 & ~n3933;
  assign n3935 = ~n3929 & n3934;
  assign n3936 = ~n3927 & ~n3935;
  assign n3937 = po53  & ~n3936;
  assign n3938 = ~po53  & n3936;
  assign n3939 = ~n3659 & po36 ;
  assign n3940 = ~n3666 & n3939;
  assign n3941 = n3664 & ~n3940;
  assign n3942 = n3667 & n3939;
  assign n3943 = ~n3941 & ~n3942;
  assign n3944 = ~n3938 & n3943;
  assign n3945 = ~n3937 & ~n3944;
  assign n3946 = po54  & ~n3945;
  assign n3947 = ~po54  & ~n3937;
  assign n3948 = ~n3944 & n3947;
  assign n3949 = ~n3669 & po36 ;
  assign n3950 = ~n3675 & n3949;
  assign n3951 = n3674 & ~n3950;
  assign n3952 = n3676 & n3949;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = ~n3948 & n3953;
  assign n3955 = ~n3946 & ~n3954;
  assign n3956 = po55  & ~n3955;
  assign n3957 = ~n3678 & ~n3680;
  assign n3958 = po36  & n3957;
  assign n3959 = n3685 & ~n3958;
  assign n3960 = ~n3685 & n3958;
  assign n3961 = ~n3959 & ~n3960;
  assign n3962 = ~po55  & n3955;
  assign n3963 = ~n3961 & ~n3962;
  assign n3964 = ~n3956 & ~n3963;
  assign n3965 = po56  & ~n3964;
  assign n3966 = ~po56  & ~n3956;
  assign n3967 = ~n3963 & n3966;
  assign n3968 = ~n3688 & po36 ;
  assign n3969 = ~n3694 & n3968;
  assign n3970 = n3693 & ~n3969;
  assign n3971 = n3695 & n3968;
  assign n3972 = ~n3970 & ~n3971;
  assign n3973 = ~n3967 & n3972;
  assign n3974 = ~n3965 & ~n3973;
  assign n3975 = po57  & ~n3974;
  assign n3976 = ~po57  & n3974;
  assign n3977 = ~n3697 & po36 ;
  assign n3978 = ~n3704 & n3977;
  assign n3979 = n3702 & ~n3978;
  assign n3980 = n3705 & n3977;
  assign n3981 = ~n3979 & ~n3980;
  assign n3982 = ~n3976 & n3981;
  assign n3983 = ~n3975 & ~n3982;
  assign n3984 = po58  & ~n3983;
  assign n3985 = ~po58  & ~n3975;
  assign n3986 = ~n3982 & n3985;
  assign n3987 = ~n3707 & po36 ;
  assign n3988 = ~n3713 & n3987;
  assign n3989 = n3712 & ~n3988;
  assign n3990 = n3714 & n3987;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992 = ~n3986 & n3991;
  assign n3993 = ~n3984 & ~n3992;
  assign n3994 = po59  & ~n3993;
  assign n3995 = ~n3716 & ~n3718;
  assign n3996 = po36  & n3995;
  assign n3997 = n3723 & ~n3996;
  assign n3998 = ~n3723 & n3996;
  assign n3999 = ~n3997 & ~n3998;
  assign n4000 = ~po59  & n3993;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = ~n3994 & ~n4001;
  assign n4003 = po60  & ~n4002;
  assign n4004 = ~po60  & ~n3994;
  assign n4005 = ~n4001 & n4004;
  assign n4006 = ~n3726 & po36 ;
  assign n4007 = ~n3732 & n4006;
  assign n4008 = n3731 & ~n4007;
  assign n4009 = n3733 & n4006;
  assign n4010 = ~n4008 & ~n4009;
  assign n4011 = ~n4005 & n4010;
  assign n4012 = ~n4003 & ~n4011;
  assign n4013 = po61  & ~n4012;
  assign n4014 = ~n3735 & ~n3737;
  assign n4015 = po36  & n4014;
  assign n4016 = n3742 & ~n4015;
  assign n4017 = ~n3742 & n4015;
  assign n4018 = ~n4016 & ~n4017;
  assign n4019 = ~po61  & n4012;
  assign n4020 = ~n4018 & ~n4019;
  assign n4021 = ~n4013 & ~n4020;
  assign n4022 = po62  & ~n4021;
  assign n4023 = ~po62  & ~n4013;
  assign n4024 = ~n4020 & n4023;
  assign n4025 = ~n3745 & po36 ;
  assign n4026 = ~n3751 & n4025;
  assign n4027 = n3750 & ~n4026;
  assign n4028 = n3752 & n4025;
  assign n4029 = ~n4027 & ~n4028;
  assign n4030 = ~n4024 & n4029;
  assign n4031 = ~n4022 & ~n4030;
  assign n4032 = ~n3754 & ~n3756;
  assign n4033 = po36  & n4032;
  assign n4034 = n3761 & ~n4033;
  assign n4035 = ~n3761 & n4033;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = n3763 & po36 ;
  assign n4038 = ~n3770 & ~n4037;
  assign n4039 = ~n3775 & ~n4038;
  assign n4040 = po36  & ~n4039;
  assign n4041 = ~n4036 & ~n4040;
  assign n4042 = ~n4031 & n4041;
  assign n4043 = ~po63  & ~n4042;
  assign n4044 = n4031 & n4036;
  assign n4045 = po63  & n4039;
  assign n4046 = ~n4044 & ~n4045;
  assign po35  = n4043 | ~n4046;
  assign n4048 = pi70  & po35 ;
  assign n4049 = ~pi68  & ~pi69 ;
  assign n4050 = ~pi70  & n4049;
  assign n4051 = ~n4048 & ~n4050;
  assign n4052 = po36  & ~n4051;
  assign n4053 = ~po36  & n4051;
  assign n4054 = ~pi70  & po35 ;
  assign n4055 = pi71  & ~n4054;
  assign n4056 = ~pi71  & n4054;
  assign n4057 = ~n4055 & ~n4056;
  assign n4058 = ~n4053 & n4057;
  assign n4059 = ~n4052 & ~n4058;
  assign n4060 = po37  & ~n4059;
  assign n4061 = po36  & ~po35 ;
  assign n4062 = ~n4056 & ~n4061;
  assign n4063 = pi72  & ~n4062;
  assign n4064 = ~pi72  & n4062;
  assign n4065 = ~n4063 & ~n4064;
  assign n4066 = ~po37  & n4059;
  assign n4067 = ~n4065 & ~n4066;
  assign n4068 = ~n4060 & ~n4067;
  assign n4069 = po38  & ~n4068;
  assign n4070 = ~po38  & ~n4060;
  assign n4071 = ~n4067 & n4070;
  assign n4072 = ~n3786 & ~n3791;
  assign n4073 = po35  & n4072;
  assign n4074 = n3790 & ~n4073;
  assign n4075 = ~n3790 & n4073;
  assign n4076 = ~n4074 & ~n4075;
  assign n4077 = ~n4071 & ~n4076;
  assign n4078 = ~n4069 & ~n4077;
  assign n4079 = po39  & ~n4078;
  assign n4080 = ~n3794 & ~n3796;
  assign n4081 = po35  & n4080;
  assign n4082 = ~n3801 & ~n4081;
  assign n4083 = n3801 & n4081;
  assign n4084 = ~n4082 & ~n4083;
  assign n4085 = ~po39  & n4078;
  assign n4086 = ~n4084 & ~n4085;
  assign n4087 = ~n4079 & ~n4086;
  assign n4088 = po40  & ~n4087;
  assign n4089 = ~po40  & ~n4079;
  assign n4090 = ~n4086 & n4089;
  assign n4091 = ~n3804 & ~n3805;
  assign n4092 = po35  & n4091;
  assign n4093 = n3810 & ~n4092;
  assign n4094 = ~n3810 & n4092;
  assign n4095 = ~n4093 & ~n4094;
  assign n4096 = ~n4090 & n4095;
  assign n4097 = ~n4088 & ~n4096;
  assign n4098 = po41  & ~n4097;
  assign n4099 = ~n3813 & ~n3815;
  assign n4100 = po35  & n4099;
  assign n4101 = n3820 & ~n4100;
  assign n4102 = ~n3820 & n4100;
  assign n4103 = ~n4101 & ~n4102;
  assign n4104 = ~po41  & n4097;
  assign n4105 = ~n4103 & ~n4104;
  assign n4106 = ~n4098 & ~n4105;
  assign n4107 = po42  & ~n4106;
  assign n4108 = ~po42  & ~n4098;
  assign n4109 = ~n4105 & n4108;
  assign n4110 = ~n3823 & ~n3824;
  assign n4111 = po35  & n4110;
  assign n4112 = n3829 & n4111;
  assign n4113 = ~n3829 & ~n4111;
  assign n4114 = ~n4112 & ~n4113;
  assign n4115 = ~n4109 & n4114;
  assign n4116 = ~n4107 & ~n4115;
  assign n4117 = po43  & ~n4116;
  assign n4118 = ~n3832 & ~n3834;
  assign n4119 = po35  & n4118;
  assign n4120 = n3839 & ~n4119;
  assign n4121 = ~n3839 & n4119;
  assign n4122 = ~n4120 & ~n4121;
  assign n4123 = ~po43  & n4116;
  assign n4124 = ~n4122 & ~n4123;
  assign n4125 = ~n4117 & ~n4124;
  assign n4126 = po44  & ~n4125;
  assign n4127 = ~po44  & ~n4117;
  assign n4128 = ~n4124 & n4127;
  assign n4129 = ~n3842 & ~n3843;
  assign n4130 = po35  & n4129;
  assign n4131 = ~n3848 & ~n4130;
  assign n4132 = n3848 & n4130;
  assign n4133 = ~n4131 & ~n4132;
  assign n4134 = ~n4128 & n4133;
  assign n4135 = ~n4126 & ~n4134;
  assign n4136 = po45  & ~n4135;
  assign n4137 = ~n3851 & ~n3853;
  assign n4138 = po35  & n4137;
  assign n4139 = n3858 & ~n4138;
  assign n4140 = ~n3858 & n4138;
  assign n4141 = ~n4139 & ~n4140;
  assign n4142 = ~po45  & n4135;
  assign n4143 = ~n4141 & ~n4142;
  assign n4144 = ~n4136 & ~n4143;
  assign n4145 = po46  & ~n4144;
  assign n4146 = ~n3861 & ~n3862;
  assign n4147 = po35  & n4146;
  assign n4148 = n3867 & ~n4147;
  assign n4149 = ~n3867 & n4147;
  assign n4150 = ~n4148 & ~n4149;
  assign n4151 = ~po46  & ~n4136;
  assign n4152 = ~n4143 & n4151;
  assign n4153 = ~n4150 & ~n4152;
  assign n4154 = ~n4145 & ~n4153;
  assign n4155 = po47  & ~n4154;
  assign n4156 = ~n3870 & ~n3872;
  assign n4157 = po35  & n4156;
  assign n4158 = n3877 & ~n4157;
  assign n4159 = ~n3877 & n4157;
  assign n4160 = ~n4158 & ~n4159;
  assign n4161 = ~po47  & n4154;
  assign n4162 = ~n4160 & ~n4161;
  assign n4163 = ~n4155 & ~n4162;
  assign n4164 = po48  & ~n4163;
  assign n4165 = ~po48  & ~n4155;
  assign n4166 = ~n4162 & n4165;
  assign n4167 = ~n3880 & po35 ;
  assign n4168 = ~n3886 & n4167;
  assign n4169 = n3885 & ~n4168;
  assign n4170 = n3887 & n4167;
  assign n4171 = ~n4169 & ~n4170;
  assign n4172 = ~n4166 & n4171;
  assign n4173 = ~n4164 & ~n4172;
  assign n4174 = po49  & ~n4173;
  assign n4175 = ~n3889 & ~n3891;
  assign n4176 = po35  & n4175;
  assign n4177 = n3896 & ~n4176;
  assign n4178 = ~n3896 & n4176;
  assign n4179 = ~n4177 & ~n4178;
  assign n4180 = ~po49  & n4173;
  assign n4181 = ~n4179 & ~n4180;
  assign n4182 = ~n4174 & ~n4181;
  assign n4183 = po50  & ~n4182;
  assign n4184 = ~n3899 & ~n3900;
  assign n4185 = po35  & n4184;
  assign n4186 = n3905 & ~n4185;
  assign n4187 = ~n3905 & n4185;
  assign n4188 = ~n4186 & ~n4187;
  assign n4189 = ~po50  & ~n4174;
  assign n4190 = ~n4181 & n4189;
  assign n4191 = ~n4188 & ~n4190;
  assign n4192 = ~n4183 & ~n4191;
  assign n4193 = po51  & ~n4192;
  assign n4194 = ~n3908 & ~n3910;
  assign n4195 = po35  & n4194;
  assign n4196 = n3915 & ~n4195;
  assign n4197 = ~n3915 & n4195;
  assign n4198 = ~n4196 & ~n4197;
  assign n4199 = ~po51  & n4192;
  assign n4200 = ~n4198 & ~n4199;
  assign n4201 = ~n4193 & ~n4200;
  assign n4202 = po52  & ~n4201;
  assign n4203 = ~po52  & ~n4193;
  assign n4204 = ~n4200 & n4203;
  assign n4205 = ~n3918 & po35 ;
  assign n4206 = ~n3924 & n4205;
  assign n4207 = n3923 & ~n4206;
  assign n4208 = n3925 & n4205;
  assign n4209 = ~n4207 & ~n4208;
  assign n4210 = ~n4204 & n4209;
  assign n4211 = ~n4202 & ~n4210;
  assign n4212 = po53  & ~n4211;
  assign n4213 = ~n3927 & ~n3929;
  assign n4214 = po35  & n4213;
  assign n4215 = n3934 & ~n4214;
  assign n4216 = ~n3934 & n4214;
  assign n4217 = ~n4215 & ~n4216;
  assign n4218 = ~po53  & n4211;
  assign n4219 = ~n4217 & ~n4218;
  assign n4220 = ~n4212 & ~n4219;
  assign n4221 = po54  & ~n4220;
  assign n4222 = ~n3937 & ~n3938;
  assign n4223 = po35  & n4222;
  assign n4224 = n3943 & ~n4223;
  assign n4225 = ~n3943 & n4223;
  assign n4226 = ~n4224 & ~n4225;
  assign n4227 = ~po54  & ~n4212;
  assign n4228 = ~n4219 & n4227;
  assign n4229 = ~n4226 & ~n4228;
  assign n4230 = ~n4221 & ~n4229;
  assign n4231 = po55  & ~n4230;
  assign n4232 = ~n3946 & ~n3948;
  assign n4233 = po35  & n4232;
  assign n4234 = n3953 & ~n4233;
  assign n4235 = ~n3953 & n4233;
  assign n4236 = ~n4234 & ~n4235;
  assign n4237 = ~po55  & n4230;
  assign n4238 = ~n4236 & ~n4237;
  assign n4239 = ~n4231 & ~n4238;
  assign n4240 = po56  & ~n4239;
  assign n4241 = ~po56  & ~n4231;
  assign n4242 = ~n4238 & n4241;
  assign n4243 = ~n3956 & po35 ;
  assign n4244 = ~n3962 & n4243;
  assign n4245 = n3961 & ~n4244;
  assign n4246 = n3963 & n4243;
  assign n4247 = ~n4245 & ~n4246;
  assign n4248 = ~n4242 & n4247;
  assign n4249 = ~n4240 & ~n4248;
  assign n4250 = po57  & ~n4249;
  assign n4251 = ~n3965 & ~n3967;
  assign n4252 = po35  & n4251;
  assign n4253 = n3972 & ~n4252;
  assign n4254 = ~n3972 & n4252;
  assign n4255 = ~n4253 & ~n4254;
  assign n4256 = ~po57  & n4249;
  assign n4257 = ~n4255 & ~n4256;
  assign n4258 = ~n4250 & ~n4257;
  assign n4259 = po58  & ~n4258;
  assign n4260 = ~n3975 & ~n3976;
  assign n4261 = po35  & n4260;
  assign n4262 = n3981 & ~n4261;
  assign n4263 = ~n3981 & n4261;
  assign n4264 = ~n4262 & ~n4263;
  assign n4265 = ~po58  & ~n4250;
  assign n4266 = ~n4257 & n4265;
  assign n4267 = ~n4264 & ~n4266;
  assign n4268 = ~n4259 & ~n4267;
  assign n4269 = po59  & ~n4268;
  assign n4270 = ~n3984 & ~n3986;
  assign n4271 = po35  & n4270;
  assign n4272 = n3991 & ~n4271;
  assign n4273 = ~n3991 & n4271;
  assign n4274 = ~n4272 & ~n4273;
  assign n4275 = ~po59  & n4268;
  assign n4276 = ~n4274 & ~n4275;
  assign n4277 = ~n4269 & ~n4276;
  assign n4278 = po60  & ~n4277;
  assign n4279 = ~po60  & ~n4269;
  assign n4280 = ~n4276 & n4279;
  assign n4281 = ~n3994 & po35 ;
  assign n4282 = ~n4000 & n4281;
  assign n4283 = n3999 & ~n4282;
  assign n4284 = n4001 & n4281;
  assign n4285 = ~n4283 & ~n4284;
  assign n4286 = ~n4280 & n4285;
  assign n4287 = ~n4278 & ~n4286;
  assign n4288 = po61  & ~n4287;
  assign n4289 = ~n4003 & ~n4005;
  assign n4290 = po35  & n4289;
  assign n4291 = n4010 & ~n4290;
  assign n4292 = ~n4010 & n4290;
  assign n4293 = ~n4291 & ~n4292;
  assign n4294 = ~po61  & n4287;
  assign n4295 = ~n4293 & ~n4294;
  assign n4296 = ~n4288 & ~n4295;
  assign n4297 = po62  & ~n4296;
  assign n4298 = ~po62  & ~n4288;
  assign n4299 = ~n4295 & n4298;
  assign n4300 = ~n4013 & po35 ;
  assign n4301 = ~n4019 & n4300;
  assign n4302 = n4018 & ~n4301;
  assign n4303 = n4020 & n4300;
  assign n4304 = ~n4302 & ~n4303;
  assign n4305 = ~n4299 & n4304;
  assign n4306 = ~n4297 & ~n4305;
  assign n4307 = ~n4022 & ~n4024;
  assign n4308 = po35  & n4307;
  assign n4309 = n4029 & ~n4308;
  assign n4310 = ~n4029 & n4308;
  assign n4311 = ~n4309 & ~n4310;
  assign n4312 = n4031 & po35 ;
  assign n4313 = ~n4036 & ~n4312;
  assign n4314 = ~n4044 & ~n4313;
  assign n4315 = po35  & ~n4314;
  assign n4316 = ~n4311 & ~n4315;
  assign n4317 = ~n4306 & n4316;
  assign n4318 = ~po63  & ~n4317;
  assign n4319 = n4306 & n4311;
  assign n4320 = po63  & n4314;
  assign n4321 = ~n4319 & ~n4320;
  assign po34  = n4318 | ~n4321;
  assign n4323 = pi68  & po34 ;
  assign n4324 = ~pi66  & ~pi67 ;
  assign n4325 = ~pi68  & n4324;
  assign n4326 = ~n4323 & ~n4325;
  assign n4327 = po35  & ~n4326;
  assign n4328 = ~pi68  & po34 ;
  assign n4329 = pi69  & ~n4328;
  assign n4330 = ~pi69  & n4328;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = ~po35  & n4326;
  assign n4333 = n4331 & ~n4332;
  assign n4334 = ~n4327 & ~n4333;
  assign n4335 = po36  & ~n4334;
  assign n4336 = ~po36  & ~n4327;
  assign n4337 = ~n4333 & n4336;
  assign n4338 = po35  & ~po34 ;
  assign n4339 = ~n4330 & ~n4338;
  assign n4340 = pi70  & ~n4339;
  assign n4341 = ~pi70  & n4339;
  assign n4342 = ~n4340 & ~n4341;
  assign n4343 = ~n4337 & ~n4342;
  assign n4344 = ~n4335 & ~n4343;
  assign n4345 = po37  & ~n4344;
  assign n4346 = ~po37  & n4344;
  assign n4347 = ~n4052 & ~n4053;
  assign n4348 = po34  & n4347;
  assign n4349 = n4057 & ~n4348;
  assign n4350 = ~n4057 & n4348;
  assign n4351 = ~n4349 & ~n4350;
  assign n4352 = ~n4346 & ~n4351;
  assign n4353 = ~n4345 & ~n4352;
  assign n4354 = po38  & ~n4353;
  assign n4355 = ~po38  & ~n4345;
  assign n4356 = ~n4352 & n4355;
  assign n4357 = ~n4060 & po34 ;
  assign n4358 = ~n4066 & n4357;
  assign n4359 = n4065 & ~n4358;
  assign n4360 = n4067 & n4357;
  assign n4361 = ~n4359 & ~n4360;
  assign n4362 = ~n4356 & n4361;
  assign n4363 = ~n4354 & ~n4362;
  assign n4364 = po39  & ~n4363;
  assign n4365 = ~po39  & n4363;
  assign n4366 = ~n4069 & ~n4071;
  assign n4367 = po34  & n4366;
  assign n4368 = n4076 & ~n4367;
  assign n4369 = ~n4076 & n4367;
  assign n4370 = ~n4368 & ~n4369;
  assign n4371 = ~n4365 & n4370;
  assign n4372 = ~n4364 & ~n4371;
  assign n4373 = po40  & ~n4372;
  assign n4374 = ~po40  & ~n4364;
  assign n4375 = ~n4371 & n4374;
  assign n4376 = ~n4079 & po34 ;
  assign n4377 = ~n4085 & n4376;
  assign n4378 = n4084 & ~n4377;
  assign n4379 = n4086 & n4376;
  assign n4380 = ~n4378 & ~n4379;
  assign n4381 = ~n4375 & n4380;
  assign n4382 = ~n4373 & ~n4381;
  assign n4383 = po41  & ~n4382;
  assign n4384 = ~po41  & n4382;
  assign n4385 = ~n4088 & ~n4090;
  assign n4386 = po34  & n4385;
  assign n4387 = n4095 & n4386;
  assign n4388 = ~n4095 & ~n4386;
  assign n4389 = ~n4387 & ~n4388;
  assign n4390 = ~n4384 & n4389;
  assign n4391 = ~n4383 & ~n4390;
  assign n4392 = po42  & ~n4391;
  assign n4393 = ~po42  & ~n4383;
  assign n4394 = ~n4390 & n4393;
  assign n4395 = ~n4098 & po34 ;
  assign n4396 = ~n4104 & n4395;
  assign n4397 = n4103 & ~n4396;
  assign n4398 = n4105 & n4395;
  assign n4399 = ~n4397 & ~n4398;
  assign n4400 = ~n4394 & n4399;
  assign n4401 = ~n4392 & ~n4400;
  assign n4402 = po43  & ~n4401;
  assign n4403 = ~po43  & n4401;
  assign n4404 = ~n4107 & ~n4109;
  assign n4405 = po34  & n4404;
  assign n4406 = ~n4114 & ~n4405;
  assign n4407 = n4114 & n4405;
  assign n4408 = ~n4406 & ~n4407;
  assign n4409 = ~n4403 & n4408;
  assign n4410 = ~n4402 & ~n4409;
  assign n4411 = po44  & ~n4410;
  assign n4412 = ~po44  & ~n4402;
  assign n4413 = ~n4409 & n4412;
  assign n4414 = ~n4117 & po34 ;
  assign n4415 = ~n4123 & n4414;
  assign n4416 = n4122 & ~n4415;
  assign n4417 = n4124 & n4414;
  assign n4418 = ~n4416 & ~n4417;
  assign n4419 = ~n4413 & n4418;
  assign n4420 = ~n4411 & ~n4419;
  assign n4421 = po45  & ~n4420;
  assign n4422 = ~n4126 & ~n4128;
  assign n4423 = po34  & n4422;
  assign n4424 = n4133 & ~n4423;
  assign n4425 = ~n4133 & n4423;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = ~po45  & n4420;
  assign n4428 = ~n4426 & ~n4427;
  assign n4429 = ~n4421 & ~n4428;
  assign n4430 = po46  & ~n4429;
  assign n4431 = ~po46  & ~n4421;
  assign n4432 = ~n4428 & n4431;
  assign n4433 = ~n4136 & po34 ;
  assign n4434 = ~n4142 & n4433;
  assign n4435 = n4141 & ~n4434;
  assign n4436 = n4143 & n4433;
  assign n4437 = ~n4435 & ~n4436;
  assign n4438 = ~n4432 & n4437;
  assign n4439 = ~n4430 & ~n4438;
  assign n4440 = po47  & ~n4439;
  assign n4441 = ~po47  & n4439;
  assign n4442 = ~n4145 & po34 ;
  assign n4443 = ~n4152 & n4442;
  assign n4444 = n4150 & ~n4443;
  assign n4445 = n4153 & n4442;
  assign n4446 = ~n4444 & ~n4445;
  assign n4447 = ~n4441 & n4446;
  assign n4448 = ~n4440 & ~n4447;
  assign n4449 = po48  & ~n4448;
  assign n4450 = ~po48  & ~n4440;
  assign n4451 = ~n4447 & n4450;
  assign n4452 = ~n4155 & po34 ;
  assign n4453 = ~n4161 & n4452;
  assign n4454 = n4160 & ~n4453;
  assign n4455 = n4162 & n4452;
  assign n4456 = ~n4454 & ~n4455;
  assign n4457 = ~n4451 & n4456;
  assign n4458 = ~n4449 & ~n4457;
  assign n4459 = po49  & ~n4458;
  assign n4460 = ~n4164 & ~n4166;
  assign n4461 = po34  & n4460;
  assign n4462 = n4171 & ~n4461;
  assign n4463 = ~n4171 & n4461;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = ~po49  & n4458;
  assign n4466 = ~n4464 & ~n4465;
  assign n4467 = ~n4459 & ~n4466;
  assign n4468 = po50  & ~n4467;
  assign n4469 = ~po50  & ~n4459;
  assign n4470 = ~n4466 & n4469;
  assign n4471 = ~n4174 & po34 ;
  assign n4472 = ~n4180 & n4471;
  assign n4473 = n4179 & ~n4472;
  assign n4474 = n4181 & n4471;
  assign n4475 = ~n4473 & ~n4474;
  assign n4476 = ~n4470 & n4475;
  assign n4477 = ~n4468 & ~n4476;
  assign n4478 = po51  & ~n4477;
  assign n4479 = ~po51  & n4477;
  assign n4480 = ~n4183 & po34 ;
  assign n4481 = ~n4190 & n4480;
  assign n4482 = n4188 & ~n4481;
  assign n4483 = n4191 & n4480;
  assign n4484 = ~n4482 & ~n4483;
  assign n4485 = ~n4479 & n4484;
  assign n4486 = ~n4478 & ~n4485;
  assign n4487 = po52  & ~n4486;
  assign n4488 = ~po52  & ~n4478;
  assign n4489 = ~n4485 & n4488;
  assign n4490 = ~n4193 & po34 ;
  assign n4491 = ~n4199 & n4490;
  assign n4492 = n4198 & ~n4491;
  assign n4493 = n4200 & n4490;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495 = ~n4489 & n4494;
  assign n4496 = ~n4487 & ~n4495;
  assign n4497 = po53  & ~n4496;
  assign n4498 = ~n4202 & ~n4204;
  assign n4499 = po34  & n4498;
  assign n4500 = n4209 & ~n4499;
  assign n4501 = ~n4209 & n4499;
  assign n4502 = ~n4500 & ~n4501;
  assign n4503 = ~po53  & n4496;
  assign n4504 = ~n4502 & ~n4503;
  assign n4505 = ~n4497 & ~n4504;
  assign n4506 = po54  & ~n4505;
  assign n4507 = ~po54  & ~n4497;
  assign n4508 = ~n4504 & n4507;
  assign n4509 = ~n4212 & po34 ;
  assign n4510 = ~n4218 & n4509;
  assign n4511 = n4217 & ~n4510;
  assign n4512 = n4219 & n4509;
  assign n4513 = ~n4511 & ~n4512;
  assign n4514 = ~n4508 & n4513;
  assign n4515 = ~n4506 & ~n4514;
  assign n4516 = po55  & ~n4515;
  assign n4517 = ~po55  & n4515;
  assign n4518 = ~n4221 & po34 ;
  assign n4519 = ~n4228 & n4518;
  assign n4520 = n4226 & ~n4519;
  assign n4521 = n4229 & n4518;
  assign n4522 = ~n4520 & ~n4521;
  assign n4523 = ~n4517 & n4522;
  assign n4524 = ~n4516 & ~n4523;
  assign n4525 = po56  & ~n4524;
  assign n4526 = ~po56  & ~n4516;
  assign n4527 = ~n4523 & n4526;
  assign n4528 = ~n4231 & po34 ;
  assign n4529 = ~n4237 & n4528;
  assign n4530 = n4236 & ~n4529;
  assign n4531 = n4238 & n4528;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = ~n4527 & n4532;
  assign n4534 = ~n4525 & ~n4533;
  assign n4535 = po57  & ~n4534;
  assign n4536 = ~n4240 & ~n4242;
  assign n4537 = po34  & n4536;
  assign n4538 = n4247 & ~n4537;
  assign n4539 = ~n4247 & n4537;
  assign n4540 = ~n4538 & ~n4539;
  assign n4541 = ~po57  & n4534;
  assign n4542 = ~n4540 & ~n4541;
  assign n4543 = ~n4535 & ~n4542;
  assign n4544 = po58  & ~n4543;
  assign n4545 = ~po58  & ~n4535;
  assign n4546 = ~n4542 & n4545;
  assign n4547 = ~n4250 & po34 ;
  assign n4548 = ~n4256 & n4547;
  assign n4549 = n4255 & ~n4548;
  assign n4550 = n4257 & n4547;
  assign n4551 = ~n4549 & ~n4550;
  assign n4552 = ~n4546 & n4551;
  assign n4553 = ~n4544 & ~n4552;
  assign n4554 = po59  & ~n4553;
  assign n4555 = ~po59  & n4553;
  assign n4556 = ~n4259 & po34 ;
  assign n4557 = ~n4266 & n4556;
  assign n4558 = n4264 & ~n4557;
  assign n4559 = n4267 & n4556;
  assign n4560 = ~n4558 & ~n4559;
  assign n4561 = ~n4555 & n4560;
  assign n4562 = ~n4554 & ~n4561;
  assign n4563 = po60  & ~n4562;
  assign n4564 = ~po60  & ~n4554;
  assign n4565 = ~n4561 & n4564;
  assign n4566 = ~n4269 & po34 ;
  assign n4567 = ~n4275 & n4566;
  assign n4568 = n4274 & ~n4567;
  assign n4569 = n4276 & n4566;
  assign n4570 = ~n4568 & ~n4569;
  assign n4571 = ~n4565 & n4570;
  assign n4572 = ~n4563 & ~n4571;
  assign n4573 = po61  & ~n4572;
  assign n4574 = ~n4278 & ~n4280;
  assign n4575 = po34  & n4574;
  assign n4576 = n4285 & ~n4575;
  assign n4577 = ~n4285 & n4575;
  assign n4578 = ~n4576 & ~n4577;
  assign n4579 = ~po61  & n4572;
  assign n4580 = ~n4578 & ~n4579;
  assign n4581 = ~n4573 & ~n4580;
  assign n4582 = po62  & ~n4581;
  assign n4583 = ~po62  & ~n4573;
  assign n4584 = ~n4580 & n4583;
  assign n4585 = ~n4288 & po34 ;
  assign n4586 = ~n4294 & n4585;
  assign n4587 = n4293 & ~n4586;
  assign n4588 = n4295 & n4585;
  assign n4589 = ~n4587 & ~n4588;
  assign n4590 = ~n4584 & n4589;
  assign n4591 = ~n4582 & ~n4590;
  assign n4592 = ~n4297 & ~n4299;
  assign n4593 = po34  & n4592;
  assign n4594 = n4304 & ~n4593;
  assign n4595 = ~n4304 & n4593;
  assign n4596 = ~n4594 & ~n4595;
  assign n4597 = n4306 & po34 ;
  assign n4598 = ~n4311 & ~n4597;
  assign n4599 = ~n4319 & ~n4598;
  assign n4600 = po34  & ~n4599;
  assign n4601 = ~n4596 & ~n4600;
  assign n4602 = ~n4591 & n4601;
  assign n4603 = ~po63  & ~n4602;
  assign n4604 = n4591 & n4596;
  assign n4605 = po63  & n4599;
  assign n4606 = ~n4604 & ~n4605;
  assign po33  = n4603 | ~n4606;
  assign n4608 = pi66  & po33 ;
  assign n4609 = ~pi64  & ~pi65 ;
  assign n4610 = ~pi66  & n4609;
  assign n4611 = ~n4608 & ~n4610;
  assign n4612 = po34  & ~n4611;
  assign n4613 = ~po34  & n4611;
  assign n4614 = ~pi66  & po33 ;
  assign n4615 = pi67  & ~n4614;
  assign n4616 = ~pi67  & n4614;
  assign n4617 = ~n4615 & ~n4616;
  assign n4618 = ~n4613 & n4617;
  assign n4619 = ~n4612 & ~n4618;
  assign n4620 = po35  & ~n4619;
  assign n4621 = po34  & ~po33 ;
  assign n4622 = ~n4616 & ~n4621;
  assign n4623 = pi68  & ~n4622;
  assign n4624 = ~pi68  & n4622;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = ~po35  & n4619;
  assign n4627 = ~n4625 & ~n4626;
  assign n4628 = ~n4620 & ~n4627;
  assign n4629 = po36  & ~n4628;
  assign n4630 = ~po36  & ~n4620;
  assign n4631 = ~n4627 & n4630;
  assign n4632 = ~n4327 & ~n4332;
  assign n4633 = po33  & n4632;
  assign n4634 = n4331 & ~n4633;
  assign n4635 = ~n4331 & n4633;
  assign n4636 = ~n4634 & ~n4635;
  assign n4637 = ~n4631 & ~n4636;
  assign n4638 = ~n4629 & ~n4637;
  assign n4639 = po37  & ~n4638;
  assign n4640 = ~n4335 & ~n4337;
  assign n4641 = po33  & n4640;
  assign n4642 = ~n4342 & ~n4641;
  assign n4643 = n4342 & n4641;
  assign n4644 = ~n4642 & ~n4643;
  assign n4645 = ~po37  & n4638;
  assign n4646 = ~n4644 & ~n4645;
  assign n4647 = ~n4639 & ~n4646;
  assign n4648 = po38  & ~n4647;
  assign n4649 = ~po38  & ~n4639;
  assign n4650 = ~n4646 & n4649;
  assign n4651 = ~n4345 & ~n4346;
  assign n4652 = po33  & n4651;
  assign n4653 = n4351 & ~n4652;
  assign n4654 = ~n4351 & n4652;
  assign n4655 = ~n4653 & ~n4654;
  assign n4656 = ~n4650 & n4655;
  assign n4657 = ~n4648 & ~n4656;
  assign n4658 = po39  & ~n4657;
  assign n4659 = ~n4354 & ~n4356;
  assign n4660 = po33  & n4659;
  assign n4661 = n4361 & ~n4660;
  assign n4662 = ~n4361 & n4660;
  assign n4663 = ~n4661 & ~n4662;
  assign n4664 = ~po39  & n4657;
  assign n4665 = ~n4663 & ~n4664;
  assign n4666 = ~n4658 & ~n4665;
  assign n4667 = po40  & ~n4666;
  assign n4668 = ~po40  & ~n4658;
  assign n4669 = ~n4665 & n4668;
  assign n4670 = ~n4364 & ~n4365;
  assign n4671 = po33  & n4670;
  assign n4672 = n4370 & n4671;
  assign n4673 = ~n4370 & ~n4671;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = ~n4669 & n4674;
  assign n4676 = ~n4667 & ~n4675;
  assign n4677 = po41  & ~n4676;
  assign n4678 = ~n4373 & ~n4375;
  assign n4679 = po33  & n4678;
  assign n4680 = n4380 & ~n4679;
  assign n4681 = ~n4380 & n4679;
  assign n4682 = ~n4680 & ~n4681;
  assign n4683 = ~po41  & n4676;
  assign n4684 = ~n4682 & ~n4683;
  assign n4685 = ~n4677 & ~n4684;
  assign n4686 = po42  & ~n4685;
  assign n4687 = ~po42  & ~n4677;
  assign n4688 = ~n4684 & n4687;
  assign n4689 = ~n4383 & ~n4384;
  assign n4690 = po33  & n4689;
  assign n4691 = ~n4389 & ~n4690;
  assign n4692 = n4389 & n4690;
  assign n4693 = ~n4691 & ~n4692;
  assign n4694 = ~n4688 & n4693;
  assign n4695 = ~n4686 & ~n4694;
  assign n4696 = po43  & ~n4695;
  assign n4697 = ~n4392 & ~n4394;
  assign n4698 = po33  & n4697;
  assign n4699 = n4399 & ~n4698;
  assign n4700 = ~n4399 & n4698;
  assign n4701 = ~n4699 & ~n4700;
  assign n4702 = ~po43  & n4695;
  assign n4703 = ~n4701 & ~n4702;
  assign n4704 = ~n4696 & ~n4703;
  assign n4705 = po44  & ~n4704;
  assign n4706 = ~n4402 & ~n4403;
  assign n4707 = po33  & n4706;
  assign n4708 = n4408 & ~n4707;
  assign n4709 = ~n4408 & n4707;
  assign n4710 = ~n4708 & ~n4709;
  assign n4711 = ~po44  & ~n4696;
  assign n4712 = ~n4703 & n4711;
  assign n4713 = ~n4710 & ~n4712;
  assign n4714 = ~n4705 & ~n4713;
  assign n4715 = po45  & ~n4714;
  assign n4716 = ~n4411 & ~n4413;
  assign n4717 = po33  & n4716;
  assign n4718 = n4418 & ~n4717;
  assign n4719 = ~n4418 & n4717;
  assign n4720 = ~n4718 & ~n4719;
  assign n4721 = ~po45  & n4714;
  assign n4722 = ~n4720 & ~n4721;
  assign n4723 = ~n4715 & ~n4722;
  assign n4724 = po46  & ~n4723;
  assign n4725 = ~po46  & ~n4715;
  assign n4726 = ~n4722 & n4725;
  assign n4727 = ~n4421 & po33 ;
  assign n4728 = ~n4427 & n4727;
  assign n4729 = n4426 & ~n4728;
  assign n4730 = n4428 & n4727;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = ~n4726 & n4731;
  assign n4733 = ~n4724 & ~n4732;
  assign n4734 = po47  & ~n4733;
  assign n4735 = ~n4430 & ~n4432;
  assign n4736 = po33  & n4735;
  assign n4737 = n4437 & ~n4736;
  assign n4738 = ~n4437 & n4736;
  assign n4739 = ~n4737 & ~n4738;
  assign n4740 = ~po47  & n4733;
  assign n4741 = ~n4739 & ~n4740;
  assign n4742 = ~n4734 & ~n4741;
  assign n4743 = po48  & ~n4742;
  assign n4744 = ~n4440 & ~n4441;
  assign n4745 = po33  & n4744;
  assign n4746 = n4446 & ~n4745;
  assign n4747 = ~n4446 & n4745;
  assign n4748 = ~n4746 & ~n4747;
  assign n4749 = ~po48  & ~n4734;
  assign n4750 = ~n4741 & n4749;
  assign n4751 = ~n4748 & ~n4750;
  assign n4752 = ~n4743 & ~n4751;
  assign n4753 = po49  & ~n4752;
  assign n4754 = ~n4449 & ~n4451;
  assign n4755 = po33  & n4754;
  assign n4756 = n4456 & ~n4755;
  assign n4757 = ~n4456 & n4755;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = ~po49  & n4752;
  assign n4760 = ~n4758 & ~n4759;
  assign n4761 = ~n4753 & ~n4760;
  assign n4762 = po50  & ~n4761;
  assign n4763 = ~po50  & ~n4753;
  assign n4764 = ~n4760 & n4763;
  assign n4765 = ~n4459 & po33 ;
  assign n4766 = ~n4465 & n4765;
  assign n4767 = n4464 & ~n4766;
  assign n4768 = n4466 & n4765;
  assign n4769 = ~n4767 & ~n4768;
  assign n4770 = ~n4764 & n4769;
  assign n4771 = ~n4762 & ~n4770;
  assign n4772 = po51  & ~n4771;
  assign n4773 = ~n4468 & ~n4470;
  assign n4774 = po33  & n4773;
  assign n4775 = n4475 & ~n4774;
  assign n4776 = ~n4475 & n4774;
  assign n4777 = ~n4775 & ~n4776;
  assign n4778 = ~po51  & n4771;
  assign n4779 = ~n4777 & ~n4778;
  assign n4780 = ~n4772 & ~n4779;
  assign n4781 = po52  & ~n4780;
  assign n4782 = ~n4478 & ~n4479;
  assign n4783 = po33  & n4782;
  assign n4784 = n4484 & ~n4783;
  assign n4785 = ~n4484 & n4783;
  assign n4786 = ~n4784 & ~n4785;
  assign n4787 = ~po52  & ~n4772;
  assign n4788 = ~n4779 & n4787;
  assign n4789 = ~n4786 & ~n4788;
  assign n4790 = ~n4781 & ~n4789;
  assign n4791 = po53  & ~n4790;
  assign n4792 = ~n4487 & ~n4489;
  assign n4793 = po33  & n4792;
  assign n4794 = n4494 & ~n4793;
  assign n4795 = ~n4494 & n4793;
  assign n4796 = ~n4794 & ~n4795;
  assign n4797 = ~po53  & n4790;
  assign n4798 = ~n4796 & ~n4797;
  assign n4799 = ~n4791 & ~n4798;
  assign n4800 = po54  & ~n4799;
  assign n4801 = ~po54  & ~n4791;
  assign n4802 = ~n4798 & n4801;
  assign n4803 = ~n4497 & po33 ;
  assign n4804 = ~n4503 & n4803;
  assign n4805 = n4502 & ~n4804;
  assign n4806 = n4504 & n4803;
  assign n4807 = ~n4805 & ~n4806;
  assign n4808 = ~n4802 & n4807;
  assign n4809 = ~n4800 & ~n4808;
  assign n4810 = po55  & ~n4809;
  assign n4811 = ~n4506 & ~n4508;
  assign n4812 = po33  & n4811;
  assign n4813 = n4513 & ~n4812;
  assign n4814 = ~n4513 & n4812;
  assign n4815 = ~n4813 & ~n4814;
  assign n4816 = ~po55  & n4809;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = ~n4810 & ~n4817;
  assign n4819 = po56  & ~n4818;
  assign n4820 = ~n4516 & ~n4517;
  assign n4821 = po33  & n4820;
  assign n4822 = n4522 & ~n4821;
  assign n4823 = ~n4522 & n4821;
  assign n4824 = ~n4822 & ~n4823;
  assign n4825 = ~po56  & ~n4810;
  assign n4826 = ~n4817 & n4825;
  assign n4827 = ~n4824 & ~n4826;
  assign n4828 = ~n4819 & ~n4827;
  assign n4829 = po57  & ~n4828;
  assign n4830 = ~n4525 & ~n4527;
  assign n4831 = po33  & n4830;
  assign n4832 = n4532 & ~n4831;
  assign n4833 = ~n4532 & n4831;
  assign n4834 = ~n4832 & ~n4833;
  assign n4835 = ~po57  & n4828;
  assign n4836 = ~n4834 & ~n4835;
  assign n4837 = ~n4829 & ~n4836;
  assign n4838 = po58  & ~n4837;
  assign n4839 = ~po58  & ~n4829;
  assign n4840 = ~n4836 & n4839;
  assign n4841 = ~n4535 & po33 ;
  assign n4842 = ~n4541 & n4841;
  assign n4843 = n4540 & ~n4842;
  assign n4844 = n4542 & n4841;
  assign n4845 = ~n4843 & ~n4844;
  assign n4846 = ~n4840 & n4845;
  assign n4847 = ~n4838 & ~n4846;
  assign n4848 = po59  & ~n4847;
  assign n4849 = ~n4544 & ~n4546;
  assign n4850 = po33  & n4849;
  assign n4851 = n4551 & ~n4850;
  assign n4852 = ~n4551 & n4850;
  assign n4853 = ~n4851 & ~n4852;
  assign n4854 = ~po59  & n4847;
  assign n4855 = ~n4853 & ~n4854;
  assign n4856 = ~n4848 & ~n4855;
  assign n4857 = po60  & ~n4856;
  assign n4858 = ~n4554 & ~n4555;
  assign n4859 = po33  & n4858;
  assign n4860 = n4560 & ~n4859;
  assign n4861 = ~n4560 & n4859;
  assign n4862 = ~n4860 & ~n4861;
  assign n4863 = ~po60  & ~n4848;
  assign n4864 = ~n4855 & n4863;
  assign n4865 = ~n4862 & ~n4864;
  assign n4866 = ~n4857 & ~n4865;
  assign n4867 = po61  & ~n4866;
  assign n4868 = ~n4563 & ~n4565;
  assign n4869 = po33  & n4868;
  assign n4870 = n4570 & ~n4869;
  assign n4871 = ~n4570 & n4869;
  assign n4872 = ~n4870 & ~n4871;
  assign n4873 = ~po61  & n4866;
  assign n4874 = ~n4872 & ~n4873;
  assign n4875 = ~n4867 & ~n4874;
  assign n4876 = po62  & ~n4875;
  assign n4877 = ~po62  & ~n4867;
  assign n4878 = ~n4874 & n4877;
  assign n4879 = ~n4573 & po33 ;
  assign n4880 = ~n4579 & n4879;
  assign n4881 = n4578 & ~n4880;
  assign n4882 = n4580 & n4879;
  assign n4883 = ~n4881 & ~n4882;
  assign n4884 = ~n4878 & n4883;
  assign n4885 = ~n4876 & ~n4884;
  assign n4886 = ~n4582 & ~n4584;
  assign n4887 = po33  & n4886;
  assign n4888 = n4589 & ~n4887;
  assign n4889 = ~n4589 & n4887;
  assign n4890 = ~n4888 & ~n4889;
  assign n4891 = n4591 & po33 ;
  assign n4892 = ~n4596 & ~n4891;
  assign n4893 = ~n4604 & ~n4892;
  assign n4894 = po33  & ~n4893;
  assign n4895 = ~n4890 & ~n4894;
  assign n4896 = ~n4885 & n4895;
  assign n4897 = ~po63  & ~n4896;
  assign n4898 = n4885 & n4890;
  assign n4899 = po63  & n4893;
  assign n4900 = ~n4898 & ~n4899;
  assign po32  = n4897 | ~n4900;
  assign n4902 = pi64  & po32 ;
  assign n4903 = ~pi62  & ~pi63 ;
  assign n4904 = ~pi64  & n4903;
  assign n4905 = ~n4902 & ~n4904;
  assign n4906 = po33  & ~n4905;
  assign n4907 = ~pi64  & po32 ;
  assign n4908 = pi65  & ~n4907;
  assign n4909 = ~pi65  & n4907;
  assign n4910 = ~n4908 & ~n4909;
  assign n4911 = ~po33  & n4905;
  assign n4912 = n4910 & ~n4911;
  assign n4913 = ~n4906 & ~n4912;
  assign n4914 = po34  & ~n4913;
  assign n4915 = ~po34  & ~n4906;
  assign n4916 = ~n4912 & n4915;
  assign n4917 = po33  & ~po32 ;
  assign n4918 = ~n4909 & ~n4917;
  assign n4919 = pi66  & ~n4918;
  assign n4920 = ~pi66  & n4918;
  assign n4921 = ~n4919 & ~n4920;
  assign n4922 = ~n4916 & ~n4921;
  assign n4923 = ~n4914 & ~n4922;
  assign n4924 = po35  & ~n4923;
  assign n4925 = ~po35  & n4923;
  assign n4926 = ~n4612 & ~n4613;
  assign n4927 = po32  & n4926;
  assign n4928 = n4617 & ~n4927;
  assign n4929 = ~n4617 & n4927;
  assign n4930 = ~n4928 & ~n4929;
  assign n4931 = ~n4925 & ~n4930;
  assign n4932 = ~n4924 & ~n4931;
  assign n4933 = po36  & ~n4932;
  assign n4934 = ~po36  & ~n4924;
  assign n4935 = ~n4931 & n4934;
  assign n4936 = ~n4620 & po32 ;
  assign n4937 = ~n4626 & n4936;
  assign n4938 = n4625 & ~n4937;
  assign n4939 = n4627 & n4936;
  assign n4940 = ~n4938 & ~n4939;
  assign n4941 = ~n4935 & n4940;
  assign n4942 = ~n4933 & ~n4941;
  assign n4943 = po37  & ~n4942;
  assign n4944 = ~po37  & n4942;
  assign n4945 = ~n4629 & ~n4631;
  assign n4946 = po32  & n4945;
  assign n4947 = n4636 & ~n4946;
  assign n4948 = ~n4636 & n4946;
  assign n4949 = ~n4947 & ~n4948;
  assign n4950 = ~n4944 & n4949;
  assign n4951 = ~n4943 & ~n4950;
  assign n4952 = po38  & ~n4951;
  assign n4953 = ~po38  & ~n4943;
  assign n4954 = ~n4950 & n4953;
  assign n4955 = ~n4639 & po32 ;
  assign n4956 = ~n4645 & n4955;
  assign n4957 = n4644 & ~n4956;
  assign n4958 = n4646 & n4955;
  assign n4959 = ~n4957 & ~n4958;
  assign n4960 = ~n4954 & n4959;
  assign n4961 = ~n4952 & ~n4960;
  assign n4962 = po39  & ~n4961;
  assign n4963 = ~po39  & n4961;
  assign n4964 = ~n4648 & ~n4650;
  assign n4965 = po32  & n4964;
  assign n4966 = n4655 & n4965;
  assign n4967 = ~n4655 & ~n4965;
  assign n4968 = ~n4966 & ~n4967;
  assign n4969 = ~n4963 & n4968;
  assign n4970 = ~n4962 & ~n4969;
  assign n4971 = po40  & ~n4970;
  assign n4972 = ~po40  & ~n4962;
  assign n4973 = ~n4969 & n4972;
  assign n4974 = ~n4658 & po32 ;
  assign n4975 = ~n4664 & n4974;
  assign n4976 = n4663 & ~n4975;
  assign n4977 = n4665 & n4974;
  assign n4978 = ~n4976 & ~n4977;
  assign n4979 = ~n4973 & n4978;
  assign n4980 = ~n4971 & ~n4979;
  assign n4981 = po41  & ~n4980;
  assign n4982 = ~po41  & n4980;
  assign n4983 = ~n4667 & ~n4669;
  assign n4984 = po32  & n4983;
  assign n4985 = ~n4674 & ~n4984;
  assign n4986 = n4674 & n4984;
  assign n4987 = ~n4985 & ~n4986;
  assign n4988 = ~n4982 & n4987;
  assign n4989 = ~n4981 & ~n4988;
  assign n4990 = po42  & ~n4989;
  assign n4991 = ~po42  & ~n4981;
  assign n4992 = ~n4988 & n4991;
  assign n4993 = ~n4677 & po32 ;
  assign n4994 = ~n4683 & n4993;
  assign n4995 = n4682 & ~n4994;
  assign n4996 = n4684 & n4993;
  assign n4997 = ~n4995 & ~n4996;
  assign n4998 = ~n4992 & n4997;
  assign n4999 = ~n4990 & ~n4998;
  assign n5000 = po43  & ~n4999;
  assign n5001 = ~n4686 & ~n4688;
  assign n5002 = po32  & n5001;
  assign n5003 = n4693 & ~n5002;
  assign n5004 = ~n4693 & n5002;
  assign n5005 = ~n5003 & ~n5004;
  assign n5006 = ~po43  & n4999;
  assign n5007 = ~n5005 & ~n5006;
  assign n5008 = ~n5000 & ~n5007;
  assign n5009 = po44  & ~n5008;
  assign n5010 = ~po44  & ~n5000;
  assign n5011 = ~n5007 & n5010;
  assign n5012 = ~n4696 & po32 ;
  assign n5013 = ~n4702 & n5012;
  assign n5014 = n4701 & ~n5013;
  assign n5015 = n4703 & n5012;
  assign n5016 = ~n5014 & ~n5015;
  assign n5017 = ~n5011 & n5016;
  assign n5018 = ~n5009 & ~n5017;
  assign n5019 = po45  & ~n5018;
  assign n5020 = ~po45  & n5018;
  assign n5021 = ~n4705 & po32 ;
  assign n5022 = ~n4712 & n5021;
  assign n5023 = n4710 & ~n5022;
  assign n5024 = n4713 & n5021;
  assign n5025 = ~n5023 & ~n5024;
  assign n5026 = ~n5020 & n5025;
  assign n5027 = ~n5019 & ~n5026;
  assign n5028 = po46  & ~n5027;
  assign n5029 = ~po46  & ~n5019;
  assign n5030 = ~n5026 & n5029;
  assign n5031 = ~n4715 & po32 ;
  assign n5032 = ~n4721 & n5031;
  assign n5033 = n4720 & ~n5032;
  assign n5034 = n4722 & n5031;
  assign n5035 = ~n5033 & ~n5034;
  assign n5036 = ~n5030 & n5035;
  assign n5037 = ~n5028 & ~n5036;
  assign n5038 = po47  & ~n5037;
  assign n5039 = ~n4724 & ~n4726;
  assign n5040 = po32  & n5039;
  assign n5041 = n4731 & ~n5040;
  assign n5042 = ~n4731 & n5040;
  assign n5043 = ~n5041 & ~n5042;
  assign n5044 = ~po47  & n5037;
  assign n5045 = ~n5043 & ~n5044;
  assign n5046 = ~n5038 & ~n5045;
  assign n5047 = po48  & ~n5046;
  assign n5048 = ~po48  & ~n5038;
  assign n5049 = ~n5045 & n5048;
  assign n5050 = ~n4734 & po32 ;
  assign n5051 = ~n4740 & n5050;
  assign n5052 = n4739 & ~n5051;
  assign n5053 = n4741 & n5050;
  assign n5054 = ~n5052 & ~n5053;
  assign n5055 = ~n5049 & n5054;
  assign n5056 = ~n5047 & ~n5055;
  assign n5057 = po49  & ~n5056;
  assign n5058 = ~po49  & n5056;
  assign n5059 = ~n4743 & po32 ;
  assign n5060 = ~n4750 & n5059;
  assign n5061 = n4748 & ~n5060;
  assign n5062 = n4751 & n5059;
  assign n5063 = ~n5061 & ~n5062;
  assign n5064 = ~n5058 & n5063;
  assign n5065 = ~n5057 & ~n5064;
  assign n5066 = po50  & ~n5065;
  assign n5067 = ~po50  & ~n5057;
  assign n5068 = ~n5064 & n5067;
  assign n5069 = ~n4753 & po32 ;
  assign n5070 = ~n4759 & n5069;
  assign n5071 = n4758 & ~n5070;
  assign n5072 = n4760 & n5069;
  assign n5073 = ~n5071 & ~n5072;
  assign n5074 = ~n5068 & n5073;
  assign n5075 = ~n5066 & ~n5074;
  assign n5076 = po51  & ~n5075;
  assign n5077 = ~n4762 & ~n4764;
  assign n5078 = po32  & n5077;
  assign n5079 = n4769 & ~n5078;
  assign n5080 = ~n4769 & n5078;
  assign n5081 = ~n5079 & ~n5080;
  assign n5082 = ~po51  & n5075;
  assign n5083 = ~n5081 & ~n5082;
  assign n5084 = ~n5076 & ~n5083;
  assign n5085 = po52  & ~n5084;
  assign n5086 = ~po52  & ~n5076;
  assign n5087 = ~n5083 & n5086;
  assign n5088 = ~n4772 & po32 ;
  assign n5089 = ~n4778 & n5088;
  assign n5090 = n4777 & ~n5089;
  assign n5091 = n4779 & n5088;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = ~n5087 & n5092;
  assign n5094 = ~n5085 & ~n5093;
  assign n5095 = po53  & ~n5094;
  assign n5096 = ~po53  & n5094;
  assign n5097 = ~n4781 & po32 ;
  assign n5098 = ~n4788 & n5097;
  assign n5099 = n4786 & ~n5098;
  assign n5100 = n4789 & n5097;
  assign n5101 = ~n5099 & ~n5100;
  assign n5102 = ~n5096 & n5101;
  assign n5103 = ~n5095 & ~n5102;
  assign n5104 = po54  & ~n5103;
  assign n5105 = ~po54  & ~n5095;
  assign n5106 = ~n5102 & n5105;
  assign n5107 = ~n4791 & po32 ;
  assign n5108 = ~n4797 & n5107;
  assign n5109 = n4796 & ~n5108;
  assign n5110 = n4798 & n5107;
  assign n5111 = ~n5109 & ~n5110;
  assign n5112 = ~n5106 & n5111;
  assign n5113 = ~n5104 & ~n5112;
  assign n5114 = po55  & ~n5113;
  assign n5115 = ~n4800 & ~n4802;
  assign n5116 = po32  & n5115;
  assign n5117 = n4807 & ~n5116;
  assign n5118 = ~n4807 & n5116;
  assign n5119 = ~n5117 & ~n5118;
  assign n5120 = ~po55  & n5113;
  assign n5121 = ~n5119 & ~n5120;
  assign n5122 = ~n5114 & ~n5121;
  assign n5123 = po56  & ~n5122;
  assign n5124 = ~po56  & ~n5114;
  assign n5125 = ~n5121 & n5124;
  assign n5126 = ~n4810 & po32 ;
  assign n5127 = ~n4816 & n5126;
  assign n5128 = n4815 & ~n5127;
  assign n5129 = n4817 & n5126;
  assign n5130 = ~n5128 & ~n5129;
  assign n5131 = ~n5125 & n5130;
  assign n5132 = ~n5123 & ~n5131;
  assign n5133 = po57  & ~n5132;
  assign n5134 = ~po57  & n5132;
  assign n5135 = ~n4819 & po32 ;
  assign n5136 = ~n4826 & n5135;
  assign n5137 = n4824 & ~n5136;
  assign n5138 = n4827 & n5135;
  assign n5139 = ~n5137 & ~n5138;
  assign n5140 = ~n5134 & n5139;
  assign n5141 = ~n5133 & ~n5140;
  assign n5142 = po58  & ~n5141;
  assign n5143 = ~po58  & ~n5133;
  assign n5144 = ~n5140 & n5143;
  assign n5145 = ~n4829 & po32 ;
  assign n5146 = ~n4835 & n5145;
  assign n5147 = n4834 & ~n5146;
  assign n5148 = n4836 & n5145;
  assign n5149 = ~n5147 & ~n5148;
  assign n5150 = ~n5144 & n5149;
  assign n5151 = ~n5142 & ~n5150;
  assign n5152 = po59  & ~n5151;
  assign n5153 = ~n4838 & ~n4840;
  assign n5154 = po32  & n5153;
  assign n5155 = n4845 & ~n5154;
  assign n5156 = ~n4845 & n5154;
  assign n5157 = ~n5155 & ~n5156;
  assign n5158 = ~po59  & n5151;
  assign n5159 = ~n5157 & ~n5158;
  assign n5160 = ~n5152 & ~n5159;
  assign n5161 = po60  & ~n5160;
  assign n5162 = ~po60  & ~n5152;
  assign n5163 = ~n5159 & n5162;
  assign n5164 = ~n4848 & po32 ;
  assign n5165 = ~n4854 & n5164;
  assign n5166 = n4853 & ~n5165;
  assign n5167 = n4855 & n5164;
  assign n5168 = ~n5166 & ~n5167;
  assign n5169 = ~n5163 & n5168;
  assign n5170 = ~n5161 & ~n5169;
  assign n5171 = po61  & ~n5170;
  assign n5172 = ~po61  & n5170;
  assign n5173 = ~n4857 & po32 ;
  assign n5174 = ~n4864 & n5173;
  assign n5175 = n4862 & ~n5174;
  assign n5176 = n4865 & n5173;
  assign n5177 = ~n5175 & ~n5176;
  assign n5178 = ~n5172 & n5177;
  assign n5179 = ~n5171 & ~n5178;
  assign n5180 = po62  & ~n5179;
  assign n5181 = ~po62  & ~n5171;
  assign n5182 = ~n5178 & n5181;
  assign n5183 = ~n4867 & po32 ;
  assign n5184 = ~n4873 & n5183;
  assign n5185 = n4872 & ~n5184;
  assign n5186 = n4874 & n5183;
  assign n5187 = ~n5185 & ~n5186;
  assign n5188 = ~n5182 & n5187;
  assign n5189 = ~n5180 & ~n5188;
  assign n5190 = ~n4876 & ~n4878;
  assign n5191 = po32  & n5190;
  assign n5192 = n4883 & ~n5191;
  assign n5193 = ~n4883 & n5191;
  assign n5194 = ~n5192 & ~n5193;
  assign n5195 = n4885 & po32 ;
  assign n5196 = ~n4890 & ~n5195;
  assign n5197 = ~n4898 & ~n5196;
  assign n5198 = po32  & ~n5197;
  assign n5199 = ~n5194 & ~n5198;
  assign n5200 = ~n5189 & n5199;
  assign n5201 = ~po63  & ~n5200;
  assign n5202 = n5189 & n5194;
  assign n5203 = po63  & n5197;
  assign n5204 = ~n5202 & ~n5203;
  assign po31  = n5201 | ~n5204;
  assign n5206 = ~pi62  & po31 ;
  assign n5207 = ~pi63  & n5206;
  assign n5208 = po32  & ~po31 ;
  assign n5209 = ~n5207 & ~n5208;
  assign n5210 = pi64  & ~n5209;
  assign n5211 = ~pi64  & n5209;
  assign n5212 = ~n5210 & ~n5211;
  assign n5213 = pi62  & po31 ;
  assign n5214 = ~pi60  & ~pi61 ;
  assign n5215 = ~pi62  & n5214;
  assign n5216 = ~n5213 & ~n5215;
  assign n5217 = po32  & ~n5216;
  assign n5218 = pi63  & ~n5206;
  assign n5219 = ~n5207 & ~n5218;
  assign n5220 = ~po32  & n5216;
  assign n5221 = n5219 & ~n5220;
  assign n5222 = ~n5217 & ~n5221;
  assign n5223 = ~po33  & n5222;
  assign n5224 = po33  & ~n5222;
  assign n5225 = ~n5212 & ~n5223;
  assign n5226 = ~n5224 & ~n5225;
  assign n5227 = po34  & ~n5226;
  assign n5228 = ~po34  & ~n5224;
  assign n5229 = ~n5225 & n5228;
  assign n5230 = ~n4906 & ~n4911;
  assign n5231 = po31  & n5230;
  assign n5232 = n4910 & ~n5231;
  assign n5233 = ~n4910 & n5231;
  assign n5234 = ~n5232 & ~n5233;
  assign n5235 = ~n5229 & ~n5234;
  assign n5236 = ~n5227 & ~n5235;
  assign n5237 = po35  & ~n5236;
  assign n5238 = ~n4914 & ~n4916;
  assign n5239 = po31  & n5238;
  assign n5240 = ~n4921 & ~n5239;
  assign n5241 = n4921 & n5239;
  assign n5242 = ~n5240 & ~n5241;
  assign n5243 = ~po35  & n5236;
  assign n5244 = ~n5242 & ~n5243;
  assign n5245 = ~n5237 & ~n5244;
  assign n5246 = po36  & ~n5245;
  assign n5247 = ~po36  & ~n5237;
  assign n5248 = ~n5244 & n5247;
  assign n5249 = ~n4924 & ~n4925;
  assign n5250 = po31  & n5249;
  assign n5251 = n4930 & ~n5250;
  assign n5252 = ~n4930 & n5250;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = ~n5248 & n5253;
  assign n5255 = ~n5246 & ~n5254;
  assign n5256 = po37  & ~n5255;
  assign n5257 = ~n4933 & ~n4935;
  assign n5258 = po31  & n5257;
  assign n5259 = n4940 & ~n5258;
  assign n5260 = ~n4940 & n5258;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = ~po37  & n5255;
  assign n5263 = ~n5261 & ~n5262;
  assign n5264 = ~n5256 & ~n5263;
  assign n5265 = po38  & ~n5264;
  assign n5266 = ~po38  & ~n5256;
  assign n5267 = ~n5263 & n5266;
  assign n5268 = ~n4943 & ~n4944;
  assign n5269 = po31  & n5268;
  assign n5270 = n4949 & n5269;
  assign n5271 = ~n4949 & ~n5269;
  assign n5272 = ~n5270 & ~n5271;
  assign n5273 = ~n5267 & n5272;
  assign n5274 = ~n5265 & ~n5273;
  assign n5275 = po39  & ~n5274;
  assign n5276 = ~n4952 & ~n4954;
  assign n5277 = po31  & n5276;
  assign n5278 = n4959 & ~n5277;
  assign n5279 = ~n4959 & n5277;
  assign n5280 = ~n5278 & ~n5279;
  assign n5281 = ~po39  & n5274;
  assign n5282 = ~n5280 & ~n5281;
  assign n5283 = ~n5275 & ~n5282;
  assign n5284 = po40  & ~n5283;
  assign n5285 = ~po40  & ~n5275;
  assign n5286 = ~n5282 & n5285;
  assign n5287 = ~n4962 & ~n4963;
  assign n5288 = po31  & n5287;
  assign n5289 = ~n4968 & ~n5288;
  assign n5290 = n4968 & n5288;
  assign n5291 = ~n5289 & ~n5290;
  assign n5292 = ~n5286 & n5291;
  assign n5293 = ~n5284 & ~n5292;
  assign n5294 = po41  & ~n5293;
  assign n5295 = ~n4971 & ~n4973;
  assign n5296 = po31  & n5295;
  assign n5297 = n4978 & ~n5296;
  assign n5298 = ~n4978 & n5296;
  assign n5299 = ~n5297 & ~n5298;
  assign n5300 = ~po41  & n5293;
  assign n5301 = ~n5299 & ~n5300;
  assign n5302 = ~n5294 & ~n5301;
  assign n5303 = po42  & ~n5302;
  assign n5304 = ~n4981 & ~n4982;
  assign n5305 = po31  & n5304;
  assign n5306 = n4987 & ~n5305;
  assign n5307 = ~n4987 & n5305;
  assign n5308 = ~n5306 & ~n5307;
  assign n5309 = ~po42  & ~n5294;
  assign n5310 = ~n5301 & n5309;
  assign n5311 = ~n5308 & ~n5310;
  assign n5312 = ~n5303 & ~n5311;
  assign n5313 = po43  & ~n5312;
  assign n5314 = ~n4990 & ~n4992;
  assign n5315 = po31  & n5314;
  assign n5316 = n4997 & ~n5315;
  assign n5317 = ~n4997 & n5315;
  assign n5318 = ~n5316 & ~n5317;
  assign n5319 = ~po43  & n5312;
  assign n5320 = ~n5318 & ~n5319;
  assign n5321 = ~n5313 & ~n5320;
  assign n5322 = po44  & ~n5321;
  assign n5323 = ~po44  & ~n5313;
  assign n5324 = ~n5320 & n5323;
  assign n5325 = ~n5000 & po31 ;
  assign n5326 = ~n5006 & n5325;
  assign n5327 = n5005 & ~n5326;
  assign n5328 = n5007 & n5325;
  assign n5329 = ~n5327 & ~n5328;
  assign n5330 = ~n5324 & n5329;
  assign n5331 = ~n5322 & ~n5330;
  assign n5332 = po45  & ~n5331;
  assign n5333 = ~n5009 & ~n5011;
  assign n5334 = po31  & n5333;
  assign n5335 = n5016 & ~n5334;
  assign n5336 = ~n5016 & n5334;
  assign n5337 = ~n5335 & ~n5336;
  assign n5338 = ~po45  & n5331;
  assign n5339 = ~n5337 & ~n5338;
  assign n5340 = ~n5332 & ~n5339;
  assign n5341 = po46  & ~n5340;
  assign n5342 = ~n5019 & ~n5020;
  assign n5343 = po31  & n5342;
  assign n5344 = n5025 & ~n5343;
  assign n5345 = ~n5025 & n5343;
  assign n5346 = ~n5344 & ~n5345;
  assign n5347 = ~po46  & ~n5332;
  assign n5348 = ~n5339 & n5347;
  assign n5349 = ~n5346 & ~n5348;
  assign n5350 = ~n5341 & ~n5349;
  assign n5351 = po47  & ~n5350;
  assign n5352 = ~n5028 & ~n5030;
  assign n5353 = po31  & n5352;
  assign n5354 = n5035 & ~n5353;
  assign n5355 = ~n5035 & n5353;
  assign n5356 = ~n5354 & ~n5355;
  assign n5357 = ~po47  & n5350;
  assign n5358 = ~n5356 & ~n5357;
  assign n5359 = ~n5351 & ~n5358;
  assign n5360 = po48  & ~n5359;
  assign n5361 = ~po48  & ~n5351;
  assign n5362 = ~n5358 & n5361;
  assign n5363 = ~n5038 & po31 ;
  assign n5364 = ~n5044 & n5363;
  assign n5365 = n5043 & ~n5364;
  assign n5366 = n5045 & n5363;
  assign n5367 = ~n5365 & ~n5366;
  assign n5368 = ~n5362 & n5367;
  assign n5369 = ~n5360 & ~n5368;
  assign n5370 = po49  & ~n5369;
  assign n5371 = ~n5047 & ~n5049;
  assign n5372 = po31  & n5371;
  assign n5373 = n5054 & ~n5372;
  assign n5374 = ~n5054 & n5372;
  assign n5375 = ~n5373 & ~n5374;
  assign n5376 = ~po49  & n5369;
  assign n5377 = ~n5375 & ~n5376;
  assign n5378 = ~n5370 & ~n5377;
  assign n5379 = po50  & ~n5378;
  assign n5380 = ~n5057 & ~n5058;
  assign n5381 = po31  & n5380;
  assign n5382 = n5063 & ~n5381;
  assign n5383 = ~n5063 & n5381;
  assign n5384 = ~n5382 & ~n5383;
  assign n5385 = ~po50  & ~n5370;
  assign n5386 = ~n5377 & n5385;
  assign n5387 = ~n5384 & ~n5386;
  assign n5388 = ~n5379 & ~n5387;
  assign n5389 = po51  & ~n5388;
  assign n5390 = ~n5066 & ~n5068;
  assign n5391 = po31  & n5390;
  assign n5392 = n5073 & ~n5391;
  assign n5393 = ~n5073 & n5391;
  assign n5394 = ~n5392 & ~n5393;
  assign n5395 = ~po51  & n5388;
  assign n5396 = ~n5394 & ~n5395;
  assign n5397 = ~n5389 & ~n5396;
  assign n5398 = po52  & ~n5397;
  assign n5399 = ~po52  & ~n5389;
  assign n5400 = ~n5396 & n5399;
  assign n5401 = ~n5076 & po31 ;
  assign n5402 = ~n5082 & n5401;
  assign n5403 = n5081 & ~n5402;
  assign n5404 = n5083 & n5401;
  assign n5405 = ~n5403 & ~n5404;
  assign n5406 = ~n5400 & n5405;
  assign n5407 = ~n5398 & ~n5406;
  assign n5408 = po53  & ~n5407;
  assign n5409 = ~n5085 & ~n5087;
  assign n5410 = po31  & n5409;
  assign n5411 = n5092 & ~n5410;
  assign n5412 = ~n5092 & n5410;
  assign n5413 = ~n5411 & ~n5412;
  assign n5414 = ~po53  & n5407;
  assign n5415 = ~n5413 & ~n5414;
  assign n5416 = ~n5408 & ~n5415;
  assign n5417 = po54  & ~n5416;
  assign n5418 = ~n5095 & ~n5096;
  assign n5419 = po31  & n5418;
  assign n5420 = n5101 & ~n5419;
  assign n5421 = ~n5101 & n5419;
  assign n5422 = ~n5420 & ~n5421;
  assign n5423 = ~po54  & ~n5408;
  assign n5424 = ~n5415 & n5423;
  assign n5425 = ~n5422 & ~n5424;
  assign n5426 = ~n5417 & ~n5425;
  assign n5427 = po55  & ~n5426;
  assign n5428 = ~n5104 & ~n5106;
  assign n5429 = po31  & n5428;
  assign n5430 = n5111 & ~n5429;
  assign n5431 = ~n5111 & n5429;
  assign n5432 = ~n5430 & ~n5431;
  assign n5433 = ~po55  & n5426;
  assign n5434 = ~n5432 & ~n5433;
  assign n5435 = ~n5427 & ~n5434;
  assign n5436 = po56  & ~n5435;
  assign n5437 = ~po56  & ~n5427;
  assign n5438 = ~n5434 & n5437;
  assign n5439 = ~n5114 & po31 ;
  assign n5440 = ~n5120 & n5439;
  assign n5441 = n5119 & ~n5440;
  assign n5442 = n5121 & n5439;
  assign n5443 = ~n5441 & ~n5442;
  assign n5444 = ~n5438 & n5443;
  assign n5445 = ~n5436 & ~n5444;
  assign n5446 = po57  & ~n5445;
  assign n5447 = ~n5123 & ~n5125;
  assign n5448 = po31  & n5447;
  assign n5449 = n5130 & ~n5448;
  assign n5450 = ~n5130 & n5448;
  assign n5451 = ~n5449 & ~n5450;
  assign n5452 = ~po57  & n5445;
  assign n5453 = ~n5451 & ~n5452;
  assign n5454 = ~n5446 & ~n5453;
  assign n5455 = po58  & ~n5454;
  assign n5456 = ~n5133 & ~n5134;
  assign n5457 = po31  & n5456;
  assign n5458 = n5139 & ~n5457;
  assign n5459 = ~n5139 & n5457;
  assign n5460 = ~n5458 & ~n5459;
  assign n5461 = ~po58  & ~n5446;
  assign n5462 = ~n5453 & n5461;
  assign n5463 = ~n5460 & ~n5462;
  assign n5464 = ~n5455 & ~n5463;
  assign n5465 = po59  & ~n5464;
  assign n5466 = ~n5142 & ~n5144;
  assign n5467 = po31  & n5466;
  assign n5468 = n5149 & ~n5467;
  assign n5469 = ~n5149 & n5467;
  assign n5470 = ~n5468 & ~n5469;
  assign n5471 = ~po59  & n5464;
  assign n5472 = ~n5470 & ~n5471;
  assign n5473 = ~n5465 & ~n5472;
  assign n5474 = po60  & ~n5473;
  assign n5475 = ~po60  & ~n5465;
  assign n5476 = ~n5472 & n5475;
  assign n5477 = ~n5152 & po31 ;
  assign n5478 = ~n5158 & n5477;
  assign n5479 = n5157 & ~n5478;
  assign n5480 = n5159 & n5477;
  assign n5481 = ~n5479 & ~n5480;
  assign n5482 = ~n5476 & n5481;
  assign n5483 = ~n5474 & ~n5482;
  assign n5484 = po61  & ~n5483;
  assign n5485 = ~n5161 & ~n5163;
  assign n5486 = po31  & n5485;
  assign n5487 = n5168 & ~n5486;
  assign n5488 = ~n5168 & n5486;
  assign n5489 = ~n5487 & ~n5488;
  assign n5490 = ~po61  & n5483;
  assign n5491 = ~n5489 & ~n5490;
  assign n5492 = ~n5484 & ~n5491;
  assign n5493 = po62  & ~n5492;
  assign n5494 = ~n5171 & ~n5172;
  assign n5495 = po31  & n5494;
  assign n5496 = n5177 & ~n5495;
  assign n5497 = ~n5177 & n5495;
  assign n5498 = ~n5496 & ~n5497;
  assign n5499 = ~po62  & ~n5484;
  assign n5500 = ~n5491 & n5499;
  assign n5501 = ~n5498 & ~n5500;
  assign n5502 = ~n5493 & ~n5501;
  assign n5503 = ~n5180 & ~n5182;
  assign n5504 = po31  & n5503;
  assign n5505 = n5187 & ~n5504;
  assign n5506 = ~n5187 & n5504;
  assign n5507 = ~n5505 & ~n5506;
  assign n5508 = n5189 & po31 ;
  assign n5509 = ~n5194 & ~n5508;
  assign n5510 = ~n5202 & ~n5509;
  assign n5511 = po31  & ~n5510;
  assign n5512 = ~n5507 & ~n5511;
  assign n5513 = ~n5502 & n5512;
  assign n5514 = ~po63  & ~n5513;
  assign n5515 = n5502 & n5507;
  assign n5516 = po63  & n5510;
  assign n5517 = ~n5515 & ~n5516;
  assign po30  = n5514 | ~n5517;
  assign n5519 = ~n5224 & po30 ;
  assign n5520 = ~n5223 & n5519;
  assign n5521 = n5212 & ~n5520;
  assign n5522 = n5225 & n5519;
  assign n5523 = ~n5521 & ~n5522;
  assign n5524 = pi60  & po30 ;
  assign n5525 = ~pi58  & ~pi59 ;
  assign n5526 = ~pi60  & n5525;
  assign n5527 = ~n5524 & ~n5526;
  assign n5528 = po31  & ~n5527;
  assign n5529 = ~pi60  & po30 ;
  assign n5530 = pi61  & ~n5529;
  assign n5531 = ~pi61  & n5529;
  assign n5532 = ~n5530 & ~n5531;
  assign n5533 = ~po31  & n5527;
  assign n5534 = n5532 & ~n5533;
  assign n5535 = ~n5528 & ~n5534;
  assign n5536 = po32  & ~n5535;
  assign n5537 = po31  & ~po30 ;
  assign n5538 = ~n5531 & ~n5537;
  assign n5539 = pi62  & ~n5538;
  assign n5540 = ~pi62  & n5538;
  assign n5541 = ~n5539 & ~n5540;
  assign n5542 = ~po32  & ~n5528;
  assign n5543 = ~n5534 & n5542;
  assign n5544 = ~n5541 & ~n5543;
  assign n5545 = ~n5536 & ~n5544;
  assign n5546 = ~po33  & n5545;
  assign n5547 = ~n5217 & ~n5220;
  assign n5548 = po30  & n5547;
  assign n5549 = n5219 & ~n5548;
  assign n5550 = ~n5219 & n5548;
  assign n5551 = ~n5549 & ~n5550;
  assign n5552 = ~n5546 & ~n5551;
  assign n5553 = po33  & ~n5545;
  assign n5554 = ~po34  & ~n5553;
  assign n5555 = ~n5552 & n5554;
  assign n5556 = ~n5552 & ~n5553;
  assign n5557 = po34  & ~n5556;
  assign n5558 = n5523 & ~n5555;
  assign n5559 = ~n5557 & ~n5558;
  assign n5560 = po35  & ~n5559;
  assign n5561 = ~po35  & n5559;
  assign n5562 = ~n5227 & ~n5229;
  assign n5563 = po30  & n5562;
  assign n5564 = n5234 & ~n5563;
  assign n5565 = ~n5234 & n5563;
  assign n5566 = ~n5564 & ~n5565;
  assign n5567 = ~n5561 & n5566;
  assign n5568 = ~n5560 & ~n5567;
  assign n5569 = po36  & ~n5568;
  assign n5570 = ~po36  & ~n5560;
  assign n5571 = ~n5567 & n5570;
  assign n5572 = ~n5237 & po30 ;
  assign n5573 = ~n5243 & n5572;
  assign n5574 = n5242 & ~n5573;
  assign n5575 = n5244 & n5572;
  assign n5576 = ~n5574 & ~n5575;
  assign n5577 = ~n5571 & n5576;
  assign n5578 = ~n5569 & ~n5577;
  assign n5579 = po37  & ~n5578;
  assign n5580 = ~po37  & n5578;
  assign n5581 = ~n5246 & ~n5248;
  assign n5582 = po30  & n5581;
  assign n5583 = n5253 & n5582;
  assign n5584 = ~n5253 & ~n5582;
  assign n5585 = ~n5583 & ~n5584;
  assign n5586 = ~n5580 & n5585;
  assign n5587 = ~n5579 & ~n5586;
  assign n5588 = po38  & ~n5587;
  assign n5589 = ~po38  & ~n5579;
  assign n5590 = ~n5586 & n5589;
  assign n5591 = ~n5256 & po30 ;
  assign n5592 = ~n5262 & n5591;
  assign n5593 = n5261 & ~n5592;
  assign n5594 = n5263 & n5591;
  assign n5595 = ~n5593 & ~n5594;
  assign n5596 = ~n5590 & n5595;
  assign n5597 = ~n5588 & ~n5596;
  assign n5598 = po39  & ~n5597;
  assign n5599 = ~po39  & n5597;
  assign n5600 = ~n5265 & ~n5267;
  assign n5601 = po30  & n5600;
  assign n5602 = ~n5272 & ~n5601;
  assign n5603 = n5272 & n5601;
  assign n5604 = ~n5602 & ~n5603;
  assign n5605 = ~n5599 & n5604;
  assign n5606 = ~n5598 & ~n5605;
  assign n5607 = po40  & ~n5606;
  assign n5608 = ~po40  & ~n5598;
  assign n5609 = ~n5605 & n5608;
  assign n5610 = ~n5275 & po30 ;
  assign n5611 = ~n5281 & n5610;
  assign n5612 = n5280 & ~n5611;
  assign n5613 = n5282 & n5610;
  assign n5614 = ~n5612 & ~n5613;
  assign n5615 = ~n5609 & n5614;
  assign n5616 = ~n5607 & ~n5615;
  assign n5617 = po41  & ~n5616;
  assign n5618 = ~n5284 & ~n5286;
  assign n5619 = po30  & n5618;
  assign n5620 = n5291 & ~n5619;
  assign n5621 = ~n5291 & n5619;
  assign n5622 = ~n5620 & ~n5621;
  assign n5623 = ~po41  & n5616;
  assign n5624 = ~n5622 & ~n5623;
  assign n5625 = ~n5617 & ~n5624;
  assign n5626 = po42  & ~n5625;
  assign n5627 = ~po42  & ~n5617;
  assign n5628 = ~n5624 & n5627;
  assign n5629 = ~n5294 & po30 ;
  assign n5630 = ~n5300 & n5629;
  assign n5631 = n5299 & ~n5630;
  assign n5632 = n5301 & n5629;
  assign n5633 = ~n5631 & ~n5632;
  assign n5634 = ~n5628 & n5633;
  assign n5635 = ~n5626 & ~n5634;
  assign n5636 = po43  & ~n5635;
  assign n5637 = ~po43  & n5635;
  assign n5638 = ~n5303 & po30 ;
  assign n5639 = ~n5310 & n5638;
  assign n5640 = n5308 & ~n5639;
  assign n5641 = n5311 & n5638;
  assign n5642 = ~n5640 & ~n5641;
  assign n5643 = ~n5637 & n5642;
  assign n5644 = ~n5636 & ~n5643;
  assign n5645 = po44  & ~n5644;
  assign n5646 = ~po44  & ~n5636;
  assign n5647 = ~n5643 & n5646;
  assign n5648 = ~n5313 & po30 ;
  assign n5649 = ~n5319 & n5648;
  assign n5650 = n5318 & ~n5649;
  assign n5651 = n5320 & n5648;
  assign n5652 = ~n5650 & ~n5651;
  assign n5653 = ~n5647 & n5652;
  assign n5654 = ~n5645 & ~n5653;
  assign n5655 = po45  & ~n5654;
  assign n5656 = ~n5322 & ~n5324;
  assign n5657 = po30  & n5656;
  assign n5658 = n5329 & ~n5657;
  assign n5659 = ~n5329 & n5657;
  assign n5660 = ~n5658 & ~n5659;
  assign n5661 = ~po45  & n5654;
  assign n5662 = ~n5660 & ~n5661;
  assign n5663 = ~n5655 & ~n5662;
  assign n5664 = po46  & ~n5663;
  assign n5665 = ~po46  & ~n5655;
  assign n5666 = ~n5662 & n5665;
  assign n5667 = ~n5332 & po30 ;
  assign n5668 = ~n5338 & n5667;
  assign n5669 = n5337 & ~n5668;
  assign n5670 = n5339 & n5667;
  assign n5671 = ~n5669 & ~n5670;
  assign n5672 = ~n5666 & n5671;
  assign n5673 = ~n5664 & ~n5672;
  assign n5674 = po47  & ~n5673;
  assign n5675 = ~po47  & n5673;
  assign n5676 = ~n5341 & po30 ;
  assign n5677 = ~n5348 & n5676;
  assign n5678 = n5346 & ~n5677;
  assign n5679 = n5349 & n5676;
  assign n5680 = ~n5678 & ~n5679;
  assign n5681 = ~n5675 & n5680;
  assign n5682 = ~n5674 & ~n5681;
  assign n5683 = po48  & ~n5682;
  assign n5684 = ~po48  & ~n5674;
  assign n5685 = ~n5681 & n5684;
  assign n5686 = ~n5351 & po30 ;
  assign n5687 = ~n5357 & n5686;
  assign n5688 = n5356 & ~n5687;
  assign n5689 = n5358 & n5686;
  assign n5690 = ~n5688 & ~n5689;
  assign n5691 = ~n5685 & n5690;
  assign n5692 = ~n5683 & ~n5691;
  assign n5693 = po49  & ~n5692;
  assign n5694 = ~n5360 & ~n5362;
  assign n5695 = po30  & n5694;
  assign n5696 = n5367 & ~n5695;
  assign n5697 = ~n5367 & n5695;
  assign n5698 = ~n5696 & ~n5697;
  assign n5699 = ~po49  & n5692;
  assign n5700 = ~n5698 & ~n5699;
  assign n5701 = ~n5693 & ~n5700;
  assign n5702 = po50  & ~n5701;
  assign n5703 = ~po50  & ~n5693;
  assign n5704 = ~n5700 & n5703;
  assign n5705 = ~n5370 & po30 ;
  assign n5706 = ~n5376 & n5705;
  assign n5707 = n5375 & ~n5706;
  assign n5708 = n5377 & n5705;
  assign n5709 = ~n5707 & ~n5708;
  assign n5710 = ~n5704 & n5709;
  assign n5711 = ~n5702 & ~n5710;
  assign n5712 = po51  & ~n5711;
  assign n5713 = ~po51  & n5711;
  assign n5714 = ~n5379 & po30 ;
  assign n5715 = ~n5386 & n5714;
  assign n5716 = n5384 & ~n5715;
  assign n5717 = n5387 & n5714;
  assign n5718 = ~n5716 & ~n5717;
  assign n5719 = ~n5713 & n5718;
  assign n5720 = ~n5712 & ~n5719;
  assign n5721 = po52  & ~n5720;
  assign n5722 = ~po52  & ~n5712;
  assign n5723 = ~n5719 & n5722;
  assign n5724 = ~n5389 & po30 ;
  assign n5725 = ~n5395 & n5724;
  assign n5726 = n5394 & ~n5725;
  assign n5727 = n5396 & n5724;
  assign n5728 = ~n5726 & ~n5727;
  assign n5729 = ~n5723 & n5728;
  assign n5730 = ~n5721 & ~n5729;
  assign n5731 = po53  & ~n5730;
  assign n5732 = ~n5398 & ~n5400;
  assign n5733 = po30  & n5732;
  assign n5734 = n5405 & ~n5733;
  assign n5735 = ~n5405 & n5733;
  assign n5736 = ~n5734 & ~n5735;
  assign n5737 = ~po53  & n5730;
  assign n5738 = ~n5736 & ~n5737;
  assign n5739 = ~n5731 & ~n5738;
  assign n5740 = po54  & ~n5739;
  assign n5741 = ~po54  & ~n5731;
  assign n5742 = ~n5738 & n5741;
  assign n5743 = ~n5408 & po30 ;
  assign n5744 = ~n5414 & n5743;
  assign n5745 = n5413 & ~n5744;
  assign n5746 = n5415 & n5743;
  assign n5747 = ~n5745 & ~n5746;
  assign n5748 = ~n5742 & n5747;
  assign n5749 = ~n5740 & ~n5748;
  assign n5750 = po55  & ~n5749;
  assign n5751 = ~po55  & n5749;
  assign n5752 = ~n5417 & po30 ;
  assign n5753 = ~n5424 & n5752;
  assign n5754 = n5422 & ~n5753;
  assign n5755 = n5425 & n5752;
  assign n5756 = ~n5754 & ~n5755;
  assign n5757 = ~n5751 & n5756;
  assign n5758 = ~n5750 & ~n5757;
  assign n5759 = po56  & ~n5758;
  assign n5760 = ~po56  & ~n5750;
  assign n5761 = ~n5757 & n5760;
  assign n5762 = ~n5427 & po30 ;
  assign n5763 = ~n5433 & n5762;
  assign n5764 = n5432 & ~n5763;
  assign n5765 = n5434 & n5762;
  assign n5766 = ~n5764 & ~n5765;
  assign n5767 = ~n5761 & n5766;
  assign n5768 = ~n5759 & ~n5767;
  assign n5769 = po57  & ~n5768;
  assign n5770 = ~n5436 & ~n5438;
  assign n5771 = po30  & n5770;
  assign n5772 = n5443 & ~n5771;
  assign n5773 = ~n5443 & n5771;
  assign n5774 = ~n5772 & ~n5773;
  assign n5775 = ~po57  & n5768;
  assign n5776 = ~n5774 & ~n5775;
  assign n5777 = ~n5769 & ~n5776;
  assign n5778 = po58  & ~n5777;
  assign n5779 = ~po58  & ~n5769;
  assign n5780 = ~n5776 & n5779;
  assign n5781 = ~n5446 & po30 ;
  assign n5782 = ~n5452 & n5781;
  assign n5783 = n5451 & ~n5782;
  assign n5784 = n5453 & n5781;
  assign n5785 = ~n5783 & ~n5784;
  assign n5786 = ~n5780 & n5785;
  assign n5787 = ~n5778 & ~n5786;
  assign n5788 = po59  & ~n5787;
  assign n5789 = ~po59  & n5787;
  assign n5790 = ~n5455 & po30 ;
  assign n5791 = ~n5462 & n5790;
  assign n5792 = n5460 & ~n5791;
  assign n5793 = n5463 & n5790;
  assign n5794 = ~n5792 & ~n5793;
  assign n5795 = ~n5789 & n5794;
  assign n5796 = ~n5788 & ~n5795;
  assign n5797 = po60  & ~n5796;
  assign n5798 = ~po60  & ~n5788;
  assign n5799 = ~n5795 & n5798;
  assign n5800 = ~n5465 & po30 ;
  assign n5801 = ~n5471 & n5800;
  assign n5802 = n5470 & ~n5801;
  assign n5803 = n5472 & n5800;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = ~n5799 & n5804;
  assign n5806 = ~n5797 & ~n5805;
  assign n5807 = po61  & ~n5806;
  assign n5808 = ~n5474 & ~n5476;
  assign n5809 = po30  & n5808;
  assign n5810 = n5481 & ~n5809;
  assign n5811 = ~n5481 & n5809;
  assign n5812 = ~n5810 & ~n5811;
  assign n5813 = ~po61  & n5806;
  assign n5814 = ~n5812 & ~n5813;
  assign n5815 = ~n5807 & ~n5814;
  assign n5816 = po62  & ~n5815;
  assign n5817 = ~po62  & ~n5807;
  assign n5818 = ~n5814 & n5817;
  assign n5819 = ~n5484 & po30 ;
  assign n5820 = ~n5490 & n5819;
  assign n5821 = n5489 & ~n5820;
  assign n5822 = n5491 & n5819;
  assign n5823 = ~n5821 & ~n5822;
  assign n5824 = ~n5818 & n5823;
  assign n5825 = ~n5816 & ~n5824;
  assign n5826 = n5502 & po30 ;
  assign n5827 = ~n5507 & ~n5826;
  assign n5828 = ~n5515 & ~n5827;
  assign n5829 = po30  & ~n5828;
  assign n5830 = ~n5493 & po30 ;
  assign n5831 = ~n5500 & n5830;
  assign n5832 = n5498 & ~n5831;
  assign n5833 = n5501 & n5830;
  assign n5834 = ~n5832 & ~n5833;
  assign n5835 = ~n5829 & n5834;
  assign n5836 = ~n5825 & n5835;
  assign n5837 = ~po63  & ~n5836;
  assign n5838 = n5825 & ~n5834;
  assign n5839 = po63  & n5828;
  assign n5840 = ~n5838 & ~n5839;
  assign po29  = n5837 | ~n5840;
  assign n5842 = ~n5555 & ~n5557;
  assign n5843 = po29  & n5842;
  assign n5844 = n5523 & ~n5843;
  assign n5845 = ~n5523 & n5843;
  assign n5846 = ~n5844 & ~n5845;
  assign n5847 = pi58  & po29 ;
  assign n5848 = ~pi56  & ~pi57 ;
  assign n5849 = ~pi58  & n5848;
  assign n5850 = ~n5847 & ~n5849;
  assign n5851 = po30  & ~n5850;
  assign n5852 = ~po30  & n5850;
  assign n5853 = ~pi58  & po29 ;
  assign n5854 = pi59  & ~n5853;
  assign n5855 = ~pi59  & n5853;
  assign n5856 = ~n5854 & ~n5855;
  assign n5857 = ~n5852 & n5856;
  assign n5858 = ~n5851 & ~n5857;
  assign n5859 = po31  & ~n5858;
  assign n5860 = po30  & ~po29 ;
  assign n5861 = ~n5855 & ~n5860;
  assign n5862 = pi60  & ~n5861;
  assign n5863 = ~pi60  & n5861;
  assign n5864 = ~n5862 & ~n5863;
  assign n5865 = ~po31  & n5858;
  assign n5866 = ~n5864 & ~n5865;
  assign n5867 = ~n5859 & ~n5866;
  assign n5868 = po32  & ~n5867;
  assign n5869 = ~po32  & ~n5859;
  assign n5870 = ~n5866 & n5869;
  assign n5871 = ~n5528 & ~n5533;
  assign n5872 = po29  & n5871;
  assign n5873 = n5532 & ~n5872;
  assign n5874 = ~n5532 & n5872;
  assign n5875 = ~n5873 & ~n5874;
  assign n5876 = ~n5870 & ~n5875;
  assign n5877 = ~n5868 & ~n5876;
  assign n5878 = ~po33  & n5877;
  assign n5879 = ~n5536 & po29 ;
  assign n5880 = ~n5543 & n5879;
  assign n5881 = n5541 & ~n5880;
  assign n5882 = n5544 & n5879;
  assign n5883 = ~n5881 & ~n5882;
  assign n5884 = ~n5878 & n5883;
  assign n5885 = po33  & ~n5877;
  assign n5886 = ~n5884 & ~n5885;
  assign n5887 = po34  & ~n5886;
  assign n5888 = ~po34  & ~n5885;
  assign n5889 = ~n5884 & n5888;
  assign n5890 = ~n5546 & ~n5553;
  assign n5891 = po29  & n5890;
  assign n5892 = n5551 & ~n5891;
  assign n5893 = ~n5551 & n5891;
  assign n5894 = ~n5892 & ~n5893;
  assign n5895 = ~n5889 & n5894;
  assign n5896 = ~n5887 & ~n5895;
  assign n5897 = ~po35  & n5896;
  assign n5898 = po35  & ~n5896;
  assign n5899 = ~n5846 & ~n5897;
  assign n5900 = ~n5898 & ~n5899;
  assign n5901 = po36  & ~n5900;
  assign n5902 = ~po36  & ~n5898;
  assign n5903 = ~n5899 & n5902;
  assign n5904 = ~n5560 & ~n5561;
  assign n5905 = po29  & n5904;
  assign n5906 = n5566 & n5905;
  assign n5907 = ~n5566 & ~n5905;
  assign n5908 = ~n5906 & ~n5907;
  assign n5909 = ~n5903 & n5908;
  assign n5910 = ~n5901 & ~n5909;
  assign n5911 = po37  & ~n5910;
  assign n5912 = ~n5569 & ~n5571;
  assign n5913 = po29  & n5912;
  assign n5914 = n5576 & ~n5913;
  assign n5915 = ~n5576 & n5913;
  assign n5916 = ~n5914 & ~n5915;
  assign n5917 = ~po37  & n5910;
  assign n5918 = ~n5916 & ~n5917;
  assign n5919 = ~n5911 & ~n5918;
  assign n5920 = po38  & ~n5919;
  assign n5921 = ~po38  & ~n5911;
  assign n5922 = ~n5918 & n5921;
  assign n5923 = ~n5579 & ~n5580;
  assign n5924 = po29  & n5923;
  assign n5925 = ~n5585 & ~n5924;
  assign n5926 = n5585 & n5924;
  assign n5927 = ~n5925 & ~n5926;
  assign n5928 = ~n5922 & n5927;
  assign n5929 = ~n5920 & ~n5928;
  assign n5930 = po39  & ~n5929;
  assign n5931 = ~n5588 & ~n5590;
  assign n5932 = po29  & n5931;
  assign n5933 = n5595 & ~n5932;
  assign n5934 = ~n5595 & n5932;
  assign n5935 = ~n5933 & ~n5934;
  assign n5936 = ~po39  & n5929;
  assign n5937 = ~n5935 & ~n5936;
  assign n5938 = ~n5930 & ~n5937;
  assign n5939 = po40  & ~n5938;
  assign n5940 = ~n5598 & ~n5599;
  assign n5941 = po29  & n5940;
  assign n5942 = n5604 & ~n5941;
  assign n5943 = ~n5604 & n5941;
  assign n5944 = ~n5942 & ~n5943;
  assign n5945 = ~po40  & ~n5930;
  assign n5946 = ~n5937 & n5945;
  assign n5947 = ~n5944 & ~n5946;
  assign n5948 = ~n5939 & ~n5947;
  assign n5949 = po41  & ~n5948;
  assign n5950 = ~n5607 & ~n5609;
  assign n5951 = po29  & n5950;
  assign n5952 = n5614 & ~n5951;
  assign n5953 = ~n5614 & n5951;
  assign n5954 = ~n5952 & ~n5953;
  assign n5955 = ~po41  & n5948;
  assign n5956 = ~n5954 & ~n5955;
  assign n5957 = ~n5949 & ~n5956;
  assign n5958 = po42  & ~n5957;
  assign n5959 = ~po42  & ~n5949;
  assign n5960 = ~n5956 & n5959;
  assign n5961 = ~n5617 & po29 ;
  assign n5962 = ~n5623 & n5961;
  assign n5963 = n5622 & ~n5962;
  assign n5964 = n5624 & n5961;
  assign n5965 = ~n5963 & ~n5964;
  assign n5966 = ~n5960 & n5965;
  assign n5967 = ~n5958 & ~n5966;
  assign n5968 = po43  & ~n5967;
  assign n5969 = ~n5626 & ~n5628;
  assign n5970 = po29  & n5969;
  assign n5971 = n5633 & ~n5970;
  assign n5972 = ~n5633 & n5970;
  assign n5973 = ~n5971 & ~n5972;
  assign n5974 = ~po43  & n5967;
  assign n5975 = ~n5973 & ~n5974;
  assign n5976 = ~n5968 & ~n5975;
  assign n5977 = po44  & ~n5976;
  assign n5978 = ~n5636 & ~n5637;
  assign n5979 = po29  & n5978;
  assign n5980 = n5642 & ~n5979;
  assign n5981 = ~n5642 & n5979;
  assign n5982 = ~n5980 & ~n5981;
  assign n5983 = ~po44  & ~n5968;
  assign n5984 = ~n5975 & n5983;
  assign n5985 = ~n5982 & ~n5984;
  assign n5986 = ~n5977 & ~n5985;
  assign n5987 = po45  & ~n5986;
  assign n5988 = ~n5645 & ~n5647;
  assign n5989 = po29  & n5988;
  assign n5990 = n5652 & ~n5989;
  assign n5991 = ~n5652 & n5989;
  assign n5992 = ~n5990 & ~n5991;
  assign n5993 = ~po45  & n5986;
  assign n5994 = ~n5992 & ~n5993;
  assign n5995 = ~n5987 & ~n5994;
  assign n5996 = po46  & ~n5995;
  assign n5997 = ~po46  & ~n5987;
  assign n5998 = ~n5994 & n5997;
  assign n5999 = ~n5655 & po29 ;
  assign n6000 = ~n5661 & n5999;
  assign n6001 = n5660 & ~n6000;
  assign n6002 = n5662 & n5999;
  assign n6003 = ~n6001 & ~n6002;
  assign n6004 = ~n5998 & n6003;
  assign n6005 = ~n5996 & ~n6004;
  assign n6006 = po47  & ~n6005;
  assign n6007 = ~n5664 & ~n5666;
  assign n6008 = po29  & n6007;
  assign n6009 = n5671 & ~n6008;
  assign n6010 = ~n5671 & n6008;
  assign n6011 = ~n6009 & ~n6010;
  assign n6012 = ~po47  & n6005;
  assign n6013 = ~n6011 & ~n6012;
  assign n6014 = ~n6006 & ~n6013;
  assign n6015 = po48  & ~n6014;
  assign n6016 = ~n5674 & ~n5675;
  assign n6017 = po29  & n6016;
  assign n6018 = n5680 & ~n6017;
  assign n6019 = ~n5680 & n6017;
  assign n6020 = ~n6018 & ~n6019;
  assign n6021 = ~po48  & ~n6006;
  assign n6022 = ~n6013 & n6021;
  assign n6023 = ~n6020 & ~n6022;
  assign n6024 = ~n6015 & ~n6023;
  assign n6025 = po49  & ~n6024;
  assign n6026 = ~n5683 & ~n5685;
  assign n6027 = po29  & n6026;
  assign n6028 = n5690 & ~n6027;
  assign n6029 = ~n5690 & n6027;
  assign n6030 = ~n6028 & ~n6029;
  assign n6031 = ~po49  & n6024;
  assign n6032 = ~n6030 & ~n6031;
  assign n6033 = ~n6025 & ~n6032;
  assign n6034 = po50  & ~n6033;
  assign n6035 = ~po50  & ~n6025;
  assign n6036 = ~n6032 & n6035;
  assign n6037 = ~n5693 & po29 ;
  assign n6038 = ~n5699 & n6037;
  assign n6039 = n5698 & ~n6038;
  assign n6040 = n5700 & n6037;
  assign n6041 = ~n6039 & ~n6040;
  assign n6042 = ~n6036 & n6041;
  assign n6043 = ~n6034 & ~n6042;
  assign n6044 = po51  & ~n6043;
  assign n6045 = ~n5702 & ~n5704;
  assign n6046 = po29  & n6045;
  assign n6047 = n5709 & ~n6046;
  assign n6048 = ~n5709 & n6046;
  assign n6049 = ~n6047 & ~n6048;
  assign n6050 = ~po51  & n6043;
  assign n6051 = ~n6049 & ~n6050;
  assign n6052 = ~n6044 & ~n6051;
  assign n6053 = po52  & ~n6052;
  assign n6054 = ~n5712 & ~n5713;
  assign n6055 = po29  & n6054;
  assign n6056 = n5718 & ~n6055;
  assign n6057 = ~n5718 & n6055;
  assign n6058 = ~n6056 & ~n6057;
  assign n6059 = ~po52  & ~n6044;
  assign n6060 = ~n6051 & n6059;
  assign n6061 = ~n6058 & ~n6060;
  assign n6062 = ~n6053 & ~n6061;
  assign n6063 = po53  & ~n6062;
  assign n6064 = ~n5721 & ~n5723;
  assign n6065 = po29  & n6064;
  assign n6066 = n5728 & ~n6065;
  assign n6067 = ~n5728 & n6065;
  assign n6068 = ~n6066 & ~n6067;
  assign n6069 = ~po53  & n6062;
  assign n6070 = ~n6068 & ~n6069;
  assign n6071 = ~n6063 & ~n6070;
  assign n6072 = po54  & ~n6071;
  assign n6073 = ~po54  & ~n6063;
  assign n6074 = ~n6070 & n6073;
  assign n6075 = ~n5731 & po29 ;
  assign n6076 = ~n5737 & n6075;
  assign n6077 = n5736 & ~n6076;
  assign n6078 = n5738 & n6075;
  assign n6079 = ~n6077 & ~n6078;
  assign n6080 = ~n6074 & n6079;
  assign n6081 = ~n6072 & ~n6080;
  assign n6082 = po55  & ~n6081;
  assign n6083 = ~n5740 & ~n5742;
  assign n6084 = po29  & n6083;
  assign n6085 = n5747 & ~n6084;
  assign n6086 = ~n5747 & n6084;
  assign n6087 = ~n6085 & ~n6086;
  assign n6088 = ~po55  & n6081;
  assign n6089 = ~n6087 & ~n6088;
  assign n6090 = ~n6082 & ~n6089;
  assign n6091 = po56  & ~n6090;
  assign n6092 = ~n5750 & ~n5751;
  assign n6093 = po29  & n6092;
  assign n6094 = n5756 & ~n6093;
  assign n6095 = ~n5756 & n6093;
  assign n6096 = ~n6094 & ~n6095;
  assign n6097 = ~po56  & ~n6082;
  assign n6098 = ~n6089 & n6097;
  assign n6099 = ~n6096 & ~n6098;
  assign n6100 = ~n6091 & ~n6099;
  assign n6101 = po57  & ~n6100;
  assign n6102 = ~n5759 & ~n5761;
  assign n6103 = po29  & n6102;
  assign n6104 = n5766 & ~n6103;
  assign n6105 = ~n5766 & n6103;
  assign n6106 = ~n6104 & ~n6105;
  assign n6107 = ~po57  & n6100;
  assign n6108 = ~n6106 & ~n6107;
  assign n6109 = ~n6101 & ~n6108;
  assign n6110 = po58  & ~n6109;
  assign n6111 = ~po58  & ~n6101;
  assign n6112 = ~n6108 & n6111;
  assign n6113 = ~n5769 & po29 ;
  assign n6114 = ~n5775 & n6113;
  assign n6115 = n5774 & ~n6114;
  assign n6116 = n5776 & n6113;
  assign n6117 = ~n6115 & ~n6116;
  assign n6118 = ~n6112 & n6117;
  assign n6119 = ~n6110 & ~n6118;
  assign n6120 = po59  & ~n6119;
  assign n6121 = ~n5778 & ~n5780;
  assign n6122 = po29  & n6121;
  assign n6123 = n5785 & ~n6122;
  assign n6124 = ~n5785 & n6122;
  assign n6125 = ~n6123 & ~n6124;
  assign n6126 = ~po59  & n6119;
  assign n6127 = ~n6125 & ~n6126;
  assign n6128 = ~n6120 & ~n6127;
  assign n6129 = po60  & ~n6128;
  assign n6130 = ~n5788 & ~n5789;
  assign n6131 = po29  & n6130;
  assign n6132 = n5794 & ~n6131;
  assign n6133 = ~n5794 & n6131;
  assign n6134 = ~n6132 & ~n6133;
  assign n6135 = ~po60  & ~n6120;
  assign n6136 = ~n6127 & n6135;
  assign n6137 = ~n6134 & ~n6136;
  assign n6138 = ~n6129 & ~n6137;
  assign n6139 = po61  & ~n6138;
  assign n6140 = ~n5797 & ~n5799;
  assign n6141 = po29  & n6140;
  assign n6142 = n5804 & ~n6141;
  assign n6143 = ~n5804 & n6141;
  assign n6144 = ~n6142 & ~n6143;
  assign n6145 = ~po61  & n6138;
  assign n6146 = ~n6144 & ~n6145;
  assign n6147 = ~n6139 & ~n6146;
  assign n6148 = po62  & ~n6147;
  assign n6149 = ~po62  & ~n6139;
  assign n6150 = ~n6146 & n6149;
  assign n6151 = ~n5807 & po29 ;
  assign n6152 = ~n5813 & n6151;
  assign n6153 = n5812 & ~n6152;
  assign n6154 = n5814 & n6151;
  assign n6155 = ~n6153 & ~n6154;
  assign n6156 = ~n6150 & n6155;
  assign n6157 = ~n6148 & ~n6156;
  assign n6158 = n5834 & po29 ;
  assign n6159 = ~n5825 & n6158;
  assign n6160 = ~n5816 & ~n5818;
  assign n6161 = po29  & n6160;
  assign n6162 = n5823 & ~n6161;
  assign n6163 = ~n5823 & n6161;
  assign n6164 = ~n6162 & ~n6163;
  assign n6165 = ~n5838 & ~n6159;
  assign n6166 = ~n6164 & n6165;
  assign n6167 = ~n6157 & n6166;
  assign n6168 = ~po63  & ~n6167;
  assign n6169 = n6157 & n6164;
  assign n6170 = n5825 & ~n6158;
  assign n6171 = ~n5825 & n5834;
  assign n6172 = po63  & ~n6171;
  assign n6173 = ~n6170 & n6172;
  assign n6174 = ~n6169 & ~n6173;
  assign po28  = n6168 | ~n6174;
  assign n6176 = ~n5898 & po28 ;
  assign n6177 = ~n5897 & n6176;
  assign n6178 = n5846 & ~n6177;
  assign n6179 = n5899 & n6176;
  assign n6180 = ~n6178 & ~n6179;
  assign n6181 = pi56  & po28 ;
  assign n6182 = ~pi54  & ~pi55 ;
  assign n6183 = ~pi56  & n6182;
  assign n6184 = ~n6181 & ~n6183;
  assign n6185 = po29  & ~n6184;
  assign n6186 = ~pi56  & po28 ;
  assign n6187 = pi57  & ~n6186;
  assign n6188 = ~pi57  & n6186;
  assign n6189 = ~n6187 & ~n6188;
  assign n6190 = ~po29  & n6184;
  assign n6191 = n6189 & ~n6190;
  assign n6192 = ~n6185 & ~n6191;
  assign n6193 = po30  & ~n6192;
  assign n6194 = ~po30  & ~n6185;
  assign n6195 = ~n6191 & n6194;
  assign n6196 = po29  & ~po28 ;
  assign n6197 = ~n6188 & ~n6196;
  assign n6198 = pi58  & ~n6197;
  assign n6199 = ~pi58  & n6197;
  assign n6200 = ~n6198 & ~n6199;
  assign n6201 = ~n6195 & ~n6200;
  assign n6202 = ~n6193 & ~n6201;
  assign n6203 = po31  & ~n6202;
  assign n6204 = ~po31  & n6202;
  assign n6205 = ~n5851 & ~n5852;
  assign n6206 = po28  & n6205;
  assign n6207 = n5856 & ~n6206;
  assign n6208 = ~n5856 & n6206;
  assign n6209 = ~n6207 & ~n6208;
  assign n6210 = ~n6204 & ~n6209;
  assign n6211 = ~n6203 & ~n6210;
  assign n6212 = po32  & ~n6211;
  assign n6213 = ~po32  & ~n6203;
  assign n6214 = ~n6210 & n6213;
  assign n6215 = ~n5859 & po28 ;
  assign n6216 = ~n5865 & n6215;
  assign n6217 = n5864 & ~n6216;
  assign n6218 = n5866 & n6215;
  assign n6219 = ~n6217 & ~n6218;
  assign n6220 = ~n6214 & n6219;
  assign n6221 = ~n6212 & ~n6220;
  assign n6222 = po33  & ~n6221;
  assign n6223 = ~po33  & n6221;
  assign n6224 = ~n5868 & ~n5870;
  assign n6225 = po28  & n6224;
  assign n6226 = n5875 & ~n6225;
  assign n6227 = ~n5875 & n6225;
  assign n6228 = ~n6226 & ~n6227;
  assign n6229 = ~n6223 & n6228;
  assign n6230 = ~n6222 & ~n6229;
  assign n6231 = po34  & ~n6230;
  assign n6232 = ~n5878 & ~n5885;
  assign n6233 = po28  & n6232;
  assign n6234 = n5883 & ~n6233;
  assign n6235 = ~n5883 & n6233;
  assign n6236 = ~n6234 & ~n6235;
  assign n6237 = ~po34  & ~n6222;
  assign n6238 = ~n6229 & n6237;
  assign n6239 = ~n6236 & ~n6238;
  assign n6240 = ~n6231 & ~n6239;
  assign n6241 = ~po35  & n6240;
  assign n6242 = ~n5887 & ~n5889;
  assign n6243 = po28  & n6242;
  assign n6244 = n5894 & n6243;
  assign n6245 = ~n5894 & ~n6243;
  assign n6246 = ~n6244 & ~n6245;
  assign n6247 = ~n6241 & n6246;
  assign n6248 = po35  & ~n6240;
  assign n6249 = ~po36  & ~n6248;
  assign n6250 = ~n6247 & n6249;
  assign n6251 = ~n6247 & ~n6248;
  assign n6252 = po36  & ~n6251;
  assign n6253 = n6180 & ~n6250;
  assign n6254 = ~n6252 & ~n6253;
  assign n6255 = po37  & ~n6254;
  assign n6256 = ~po37  & n6254;
  assign n6257 = ~n5901 & ~n5903;
  assign n6258 = po28  & n6257;
  assign n6259 = n5908 & n6258;
  assign n6260 = ~n5908 & ~n6258;
  assign n6261 = ~n6259 & ~n6260;
  assign n6262 = ~n6256 & n6261;
  assign n6263 = ~n6255 & ~n6262;
  assign n6264 = po38  & ~n6263;
  assign n6265 = ~po38  & ~n6255;
  assign n6266 = ~n6262 & n6265;
  assign n6267 = ~n5911 & po28 ;
  assign n6268 = ~n5917 & n6267;
  assign n6269 = n5916 & ~n6268;
  assign n6270 = n5918 & n6267;
  assign n6271 = ~n6269 & ~n6270;
  assign n6272 = ~n6266 & n6271;
  assign n6273 = ~n6264 & ~n6272;
  assign n6274 = po39  & ~n6273;
  assign n6275 = ~n5920 & ~n5922;
  assign n6276 = po28  & n6275;
  assign n6277 = n5927 & ~n6276;
  assign n6278 = ~n5927 & n6276;
  assign n6279 = ~n6277 & ~n6278;
  assign n6280 = ~po39  & n6273;
  assign n6281 = ~n6279 & ~n6280;
  assign n6282 = ~n6274 & ~n6281;
  assign n6283 = po40  & ~n6282;
  assign n6284 = ~po40  & ~n6274;
  assign n6285 = ~n6281 & n6284;
  assign n6286 = ~n5930 & po28 ;
  assign n6287 = ~n5936 & n6286;
  assign n6288 = n5935 & ~n6287;
  assign n6289 = n5937 & n6286;
  assign n6290 = ~n6288 & ~n6289;
  assign n6291 = ~n6285 & n6290;
  assign n6292 = ~n6283 & ~n6291;
  assign n6293 = po41  & ~n6292;
  assign n6294 = ~po41  & n6292;
  assign n6295 = ~n5939 & po28 ;
  assign n6296 = ~n5946 & n6295;
  assign n6297 = n5944 & ~n6296;
  assign n6298 = n5947 & n6295;
  assign n6299 = ~n6297 & ~n6298;
  assign n6300 = ~n6294 & n6299;
  assign n6301 = ~n6293 & ~n6300;
  assign n6302 = po42  & ~n6301;
  assign n6303 = ~po42  & ~n6293;
  assign n6304 = ~n6300 & n6303;
  assign n6305 = ~n5949 & po28 ;
  assign n6306 = ~n5955 & n6305;
  assign n6307 = n5954 & ~n6306;
  assign n6308 = n5956 & n6305;
  assign n6309 = ~n6307 & ~n6308;
  assign n6310 = ~n6304 & n6309;
  assign n6311 = ~n6302 & ~n6310;
  assign n6312 = po43  & ~n6311;
  assign n6313 = ~n5958 & ~n5960;
  assign n6314 = po28  & n6313;
  assign n6315 = n5965 & ~n6314;
  assign n6316 = ~n5965 & n6314;
  assign n6317 = ~n6315 & ~n6316;
  assign n6318 = ~po43  & n6311;
  assign n6319 = ~n6317 & ~n6318;
  assign n6320 = ~n6312 & ~n6319;
  assign n6321 = po44  & ~n6320;
  assign n6322 = ~po44  & ~n6312;
  assign n6323 = ~n6319 & n6322;
  assign n6324 = ~n5968 & po28 ;
  assign n6325 = ~n5974 & n6324;
  assign n6326 = n5973 & ~n6325;
  assign n6327 = n5975 & n6324;
  assign n6328 = ~n6326 & ~n6327;
  assign n6329 = ~n6323 & n6328;
  assign n6330 = ~n6321 & ~n6329;
  assign n6331 = po45  & ~n6330;
  assign n6332 = ~po45  & n6330;
  assign n6333 = ~n5977 & po28 ;
  assign n6334 = ~n5984 & n6333;
  assign n6335 = n5982 & ~n6334;
  assign n6336 = n5985 & n6333;
  assign n6337 = ~n6335 & ~n6336;
  assign n6338 = ~n6332 & n6337;
  assign n6339 = ~n6331 & ~n6338;
  assign n6340 = po46  & ~n6339;
  assign n6341 = ~po46  & ~n6331;
  assign n6342 = ~n6338 & n6341;
  assign n6343 = ~n5987 & po28 ;
  assign n6344 = ~n5993 & n6343;
  assign n6345 = n5992 & ~n6344;
  assign n6346 = n5994 & n6343;
  assign n6347 = ~n6345 & ~n6346;
  assign n6348 = ~n6342 & n6347;
  assign n6349 = ~n6340 & ~n6348;
  assign n6350 = po47  & ~n6349;
  assign n6351 = ~n5996 & ~n5998;
  assign n6352 = po28  & n6351;
  assign n6353 = n6003 & ~n6352;
  assign n6354 = ~n6003 & n6352;
  assign n6355 = ~n6353 & ~n6354;
  assign n6356 = ~po47  & n6349;
  assign n6357 = ~n6355 & ~n6356;
  assign n6358 = ~n6350 & ~n6357;
  assign n6359 = po48  & ~n6358;
  assign n6360 = ~po48  & ~n6350;
  assign n6361 = ~n6357 & n6360;
  assign n6362 = ~n6006 & po28 ;
  assign n6363 = ~n6012 & n6362;
  assign n6364 = n6011 & ~n6363;
  assign n6365 = n6013 & n6362;
  assign n6366 = ~n6364 & ~n6365;
  assign n6367 = ~n6361 & n6366;
  assign n6368 = ~n6359 & ~n6367;
  assign n6369 = po49  & ~n6368;
  assign n6370 = ~po49  & n6368;
  assign n6371 = ~n6015 & po28 ;
  assign n6372 = ~n6022 & n6371;
  assign n6373 = n6020 & ~n6372;
  assign n6374 = n6023 & n6371;
  assign n6375 = ~n6373 & ~n6374;
  assign n6376 = ~n6370 & n6375;
  assign n6377 = ~n6369 & ~n6376;
  assign n6378 = po50  & ~n6377;
  assign n6379 = ~po50  & ~n6369;
  assign n6380 = ~n6376 & n6379;
  assign n6381 = ~n6025 & po28 ;
  assign n6382 = ~n6031 & n6381;
  assign n6383 = n6030 & ~n6382;
  assign n6384 = n6032 & n6381;
  assign n6385 = ~n6383 & ~n6384;
  assign n6386 = ~n6380 & n6385;
  assign n6387 = ~n6378 & ~n6386;
  assign n6388 = po51  & ~n6387;
  assign n6389 = ~n6034 & ~n6036;
  assign n6390 = po28  & n6389;
  assign n6391 = n6041 & ~n6390;
  assign n6392 = ~n6041 & n6390;
  assign n6393 = ~n6391 & ~n6392;
  assign n6394 = ~po51  & n6387;
  assign n6395 = ~n6393 & ~n6394;
  assign n6396 = ~n6388 & ~n6395;
  assign n6397 = po52  & ~n6396;
  assign n6398 = ~po52  & ~n6388;
  assign n6399 = ~n6395 & n6398;
  assign n6400 = ~n6044 & po28 ;
  assign n6401 = ~n6050 & n6400;
  assign n6402 = n6049 & ~n6401;
  assign n6403 = n6051 & n6400;
  assign n6404 = ~n6402 & ~n6403;
  assign n6405 = ~n6399 & n6404;
  assign n6406 = ~n6397 & ~n6405;
  assign n6407 = po53  & ~n6406;
  assign n6408 = ~po53  & n6406;
  assign n6409 = ~n6053 & po28 ;
  assign n6410 = ~n6060 & n6409;
  assign n6411 = n6058 & ~n6410;
  assign n6412 = n6061 & n6409;
  assign n6413 = ~n6411 & ~n6412;
  assign n6414 = ~n6408 & n6413;
  assign n6415 = ~n6407 & ~n6414;
  assign n6416 = po54  & ~n6415;
  assign n6417 = ~po54  & ~n6407;
  assign n6418 = ~n6414 & n6417;
  assign n6419 = ~n6063 & po28 ;
  assign n6420 = ~n6069 & n6419;
  assign n6421 = n6068 & ~n6420;
  assign n6422 = n6070 & n6419;
  assign n6423 = ~n6421 & ~n6422;
  assign n6424 = ~n6418 & n6423;
  assign n6425 = ~n6416 & ~n6424;
  assign n6426 = po55  & ~n6425;
  assign n6427 = ~n6072 & ~n6074;
  assign n6428 = po28  & n6427;
  assign n6429 = n6079 & ~n6428;
  assign n6430 = ~n6079 & n6428;
  assign n6431 = ~n6429 & ~n6430;
  assign n6432 = ~po55  & n6425;
  assign n6433 = ~n6431 & ~n6432;
  assign n6434 = ~n6426 & ~n6433;
  assign n6435 = po56  & ~n6434;
  assign n6436 = ~po56  & ~n6426;
  assign n6437 = ~n6433 & n6436;
  assign n6438 = ~n6082 & po28 ;
  assign n6439 = ~n6088 & n6438;
  assign n6440 = n6087 & ~n6439;
  assign n6441 = n6089 & n6438;
  assign n6442 = ~n6440 & ~n6441;
  assign n6443 = ~n6437 & n6442;
  assign n6444 = ~n6435 & ~n6443;
  assign n6445 = po57  & ~n6444;
  assign n6446 = ~po57  & n6444;
  assign n6447 = ~n6091 & po28 ;
  assign n6448 = ~n6098 & n6447;
  assign n6449 = n6096 & ~n6448;
  assign n6450 = n6099 & n6447;
  assign n6451 = ~n6449 & ~n6450;
  assign n6452 = ~n6446 & n6451;
  assign n6453 = ~n6445 & ~n6452;
  assign n6454 = po58  & ~n6453;
  assign n6455 = ~po58  & ~n6445;
  assign n6456 = ~n6452 & n6455;
  assign n6457 = ~n6101 & po28 ;
  assign n6458 = ~n6107 & n6457;
  assign n6459 = n6106 & ~n6458;
  assign n6460 = n6108 & n6457;
  assign n6461 = ~n6459 & ~n6460;
  assign n6462 = ~n6456 & n6461;
  assign n6463 = ~n6454 & ~n6462;
  assign n6464 = po59  & ~n6463;
  assign n6465 = ~n6110 & ~n6112;
  assign n6466 = po28  & n6465;
  assign n6467 = n6117 & ~n6466;
  assign n6468 = ~n6117 & n6466;
  assign n6469 = ~n6467 & ~n6468;
  assign n6470 = ~po59  & n6463;
  assign n6471 = ~n6469 & ~n6470;
  assign n6472 = ~n6464 & ~n6471;
  assign n6473 = po60  & ~n6472;
  assign n6474 = ~po60  & ~n6464;
  assign n6475 = ~n6471 & n6474;
  assign n6476 = ~n6120 & po28 ;
  assign n6477 = ~n6126 & n6476;
  assign n6478 = n6125 & ~n6477;
  assign n6479 = n6127 & n6476;
  assign n6480 = ~n6478 & ~n6479;
  assign n6481 = ~n6475 & n6480;
  assign n6482 = ~n6473 & ~n6481;
  assign n6483 = po61  & ~n6482;
  assign n6484 = ~po61  & n6482;
  assign n6485 = ~n6129 & po28 ;
  assign n6486 = ~n6136 & n6485;
  assign n6487 = n6134 & ~n6486;
  assign n6488 = n6137 & n6485;
  assign n6489 = ~n6487 & ~n6488;
  assign n6490 = ~n6484 & n6489;
  assign n6491 = ~n6483 & ~n6490;
  assign n6492 = po62  & ~n6491;
  assign n6493 = ~po62  & ~n6483;
  assign n6494 = ~n6490 & n6493;
  assign n6495 = ~n6139 & po28 ;
  assign n6496 = ~n6145 & n6495;
  assign n6497 = n6144 & ~n6496;
  assign n6498 = n6146 & n6495;
  assign n6499 = ~n6497 & ~n6498;
  assign n6500 = ~n6494 & n6499;
  assign n6501 = ~n6492 & ~n6500;
  assign n6502 = ~n6148 & ~n6150;
  assign n6503 = po28  & n6502;
  assign n6504 = n6155 & ~n6503;
  assign n6505 = ~n6155 & n6503;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = n6157 & po28 ;
  assign n6508 = ~n6164 & ~n6507;
  assign n6509 = ~n6169 & ~n6508;
  assign n6510 = po28  & ~n6509;
  assign n6511 = ~n6506 & ~n6510;
  assign n6512 = ~n6501 & n6511;
  assign n6513 = ~po63  & ~n6512;
  assign n6514 = n6501 & n6506;
  assign n6515 = po63  & n6509;
  assign n6516 = ~n6514 & ~n6515;
  assign po27  = n6513 | ~n6516;
  assign n6518 = ~n6250 & ~n6252;
  assign n6519 = po27  & n6518;
  assign n6520 = n6180 & ~n6519;
  assign n6521 = ~n6180 & n6519;
  assign n6522 = ~n6520 & ~n6521;
  assign n6523 = pi54  & po27 ;
  assign n6524 = ~pi52  & ~pi53 ;
  assign n6525 = ~pi54  & n6524;
  assign n6526 = ~n6523 & ~n6525;
  assign n6527 = po28  & ~n6526;
  assign n6528 = ~po28  & n6526;
  assign n6529 = ~pi54  & po27 ;
  assign n6530 = pi55  & ~n6529;
  assign n6531 = ~pi55  & n6529;
  assign n6532 = ~n6530 & ~n6531;
  assign n6533 = ~n6528 & n6532;
  assign n6534 = ~n6527 & ~n6533;
  assign n6535 = po29  & ~n6534;
  assign n6536 = po28  & ~po27 ;
  assign n6537 = ~n6531 & ~n6536;
  assign n6538 = pi56  & ~n6537;
  assign n6539 = ~pi56  & n6537;
  assign n6540 = ~n6538 & ~n6539;
  assign n6541 = ~po29  & n6534;
  assign n6542 = ~n6540 & ~n6541;
  assign n6543 = ~n6535 & ~n6542;
  assign n6544 = po30  & ~n6543;
  assign n6545 = ~po30  & ~n6535;
  assign n6546 = ~n6542 & n6545;
  assign n6547 = ~n6185 & ~n6190;
  assign n6548 = po27  & n6547;
  assign n6549 = n6189 & ~n6548;
  assign n6550 = ~n6189 & n6548;
  assign n6551 = ~n6549 & ~n6550;
  assign n6552 = ~n6546 & ~n6551;
  assign n6553 = ~n6544 & ~n6552;
  assign n6554 = po31  & ~n6553;
  assign n6555 = ~n6193 & ~n6195;
  assign n6556 = po27  & n6555;
  assign n6557 = ~n6200 & ~n6556;
  assign n6558 = n6200 & n6556;
  assign n6559 = ~n6557 & ~n6558;
  assign n6560 = ~po31  & n6553;
  assign n6561 = ~n6559 & ~n6560;
  assign n6562 = ~n6554 & ~n6561;
  assign n6563 = po32  & ~n6562;
  assign n6564 = ~po32  & ~n6554;
  assign n6565 = ~n6561 & n6564;
  assign n6566 = ~n6203 & ~n6204;
  assign n6567 = po27  & n6566;
  assign n6568 = n6209 & ~n6567;
  assign n6569 = ~n6209 & n6567;
  assign n6570 = ~n6568 & ~n6569;
  assign n6571 = ~n6565 & n6570;
  assign n6572 = ~n6563 & ~n6571;
  assign n6573 = po33  & ~n6572;
  assign n6574 = ~n6212 & ~n6214;
  assign n6575 = po27  & n6574;
  assign n6576 = n6219 & ~n6575;
  assign n6577 = ~n6219 & n6575;
  assign n6578 = ~n6576 & ~n6577;
  assign n6579 = ~po33  & n6572;
  assign n6580 = ~n6578 & ~n6579;
  assign n6581 = ~n6573 & ~n6580;
  assign n6582 = po34  & ~n6581;
  assign n6583 = ~po34  & ~n6573;
  assign n6584 = ~n6580 & n6583;
  assign n6585 = ~n6222 & ~n6223;
  assign n6586 = po27  & n6585;
  assign n6587 = n6228 & n6586;
  assign n6588 = ~n6228 & ~n6586;
  assign n6589 = ~n6587 & ~n6588;
  assign n6590 = ~n6584 & n6589;
  assign n6591 = ~n6582 & ~n6590;
  assign n6592 = ~po35  & n6591;
  assign n6593 = ~n6231 & po27 ;
  assign n6594 = ~n6238 & n6593;
  assign n6595 = n6236 & ~n6594;
  assign n6596 = n6239 & n6593;
  assign n6597 = ~n6595 & ~n6596;
  assign n6598 = ~n6592 & n6597;
  assign n6599 = po35  & ~n6591;
  assign n6600 = ~n6598 & ~n6599;
  assign n6601 = po36  & ~n6600;
  assign n6602 = ~n6241 & ~n6248;
  assign n6603 = po27  & n6602;
  assign n6604 = ~n6246 & ~n6603;
  assign n6605 = n6246 & n6603;
  assign n6606 = ~n6604 & ~n6605;
  assign n6607 = ~po36  & ~n6599;
  assign n6608 = ~n6598 & n6607;
  assign n6609 = n6606 & ~n6608;
  assign n6610 = ~n6601 & ~n6609;
  assign n6611 = ~po37  & n6610;
  assign n6612 = po37  & ~n6610;
  assign n6613 = ~n6522 & ~n6611;
  assign n6614 = ~n6612 & ~n6613;
  assign n6615 = po38  & ~n6614;
  assign n6616 = ~po38  & ~n6612;
  assign n6617 = ~n6613 & n6616;
  assign n6618 = ~n6255 & ~n6256;
  assign n6619 = po27  & n6618;
  assign n6620 = ~n6261 & ~n6619;
  assign n6621 = n6261 & n6619;
  assign n6622 = ~n6620 & ~n6621;
  assign n6623 = ~n6617 & n6622;
  assign n6624 = ~n6615 & ~n6623;
  assign n6625 = po39  & ~n6624;
  assign n6626 = ~n6264 & ~n6266;
  assign n6627 = po27  & n6626;
  assign n6628 = n6271 & ~n6627;
  assign n6629 = ~n6271 & n6627;
  assign n6630 = ~n6628 & ~n6629;
  assign n6631 = ~po39  & n6624;
  assign n6632 = ~n6630 & ~n6631;
  assign n6633 = ~n6625 & ~n6632;
  assign n6634 = po40  & ~n6633;
  assign n6635 = ~po40  & ~n6625;
  assign n6636 = ~n6632 & n6635;
  assign n6637 = ~n6274 & po27 ;
  assign n6638 = ~n6280 & n6637;
  assign n6639 = n6279 & ~n6638;
  assign n6640 = n6281 & n6637;
  assign n6641 = ~n6639 & ~n6640;
  assign n6642 = ~n6636 & n6641;
  assign n6643 = ~n6634 & ~n6642;
  assign n6644 = po41  & ~n6643;
  assign n6645 = ~n6283 & ~n6285;
  assign n6646 = po27  & n6645;
  assign n6647 = n6290 & ~n6646;
  assign n6648 = ~n6290 & n6646;
  assign n6649 = ~n6647 & ~n6648;
  assign n6650 = ~po41  & n6643;
  assign n6651 = ~n6649 & ~n6650;
  assign n6652 = ~n6644 & ~n6651;
  assign n6653 = po42  & ~n6652;
  assign n6654 = ~n6293 & ~n6294;
  assign n6655 = po27  & n6654;
  assign n6656 = n6299 & ~n6655;
  assign n6657 = ~n6299 & n6655;
  assign n6658 = ~n6656 & ~n6657;
  assign n6659 = ~po42  & ~n6644;
  assign n6660 = ~n6651 & n6659;
  assign n6661 = ~n6658 & ~n6660;
  assign n6662 = ~n6653 & ~n6661;
  assign n6663 = po43  & ~n6662;
  assign n6664 = ~n6302 & ~n6304;
  assign n6665 = po27  & n6664;
  assign n6666 = n6309 & ~n6665;
  assign n6667 = ~n6309 & n6665;
  assign n6668 = ~n6666 & ~n6667;
  assign n6669 = ~po43  & n6662;
  assign n6670 = ~n6668 & ~n6669;
  assign n6671 = ~n6663 & ~n6670;
  assign n6672 = po44  & ~n6671;
  assign n6673 = ~po44  & ~n6663;
  assign n6674 = ~n6670 & n6673;
  assign n6675 = ~n6312 & po27 ;
  assign n6676 = ~n6318 & n6675;
  assign n6677 = n6317 & ~n6676;
  assign n6678 = n6319 & n6675;
  assign n6679 = ~n6677 & ~n6678;
  assign n6680 = ~n6674 & n6679;
  assign n6681 = ~n6672 & ~n6680;
  assign n6682 = po45  & ~n6681;
  assign n6683 = ~n6321 & ~n6323;
  assign n6684 = po27  & n6683;
  assign n6685 = n6328 & ~n6684;
  assign n6686 = ~n6328 & n6684;
  assign n6687 = ~n6685 & ~n6686;
  assign n6688 = ~po45  & n6681;
  assign n6689 = ~n6687 & ~n6688;
  assign n6690 = ~n6682 & ~n6689;
  assign n6691 = po46  & ~n6690;
  assign n6692 = ~n6331 & ~n6332;
  assign n6693 = po27  & n6692;
  assign n6694 = n6337 & ~n6693;
  assign n6695 = ~n6337 & n6693;
  assign n6696 = ~n6694 & ~n6695;
  assign n6697 = ~po46  & ~n6682;
  assign n6698 = ~n6689 & n6697;
  assign n6699 = ~n6696 & ~n6698;
  assign n6700 = ~n6691 & ~n6699;
  assign n6701 = po47  & ~n6700;
  assign n6702 = ~n6340 & ~n6342;
  assign n6703 = po27  & n6702;
  assign n6704 = n6347 & ~n6703;
  assign n6705 = ~n6347 & n6703;
  assign n6706 = ~n6704 & ~n6705;
  assign n6707 = ~po47  & n6700;
  assign n6708 = ~n6706 & ~n6707;
  assign n6709 = ~n6701 & ~n6708;
  assign n6710 = po48  & ~n6709;
  assign n6711 = ~po48  & ~n6701;
  assign n6712 = ~n6708 & n6711;
  assign n6713 = ~n6350 & po27 ;
  assign n6714 = ~n6356 & n6713;
  assign n6715 = n6355 & ~n6714;
  assign n6716 = n6357 & n6713;
  assign n6717 = ~n6715 & ~n6716;
  assign n6718 = ~n6712 & n6717;
  assign n6719 = ~n6710 & ~n6718;
  assign n6720 = po49  & ~n6719;
  assign n6721 = ~n6359 & ~n6361;
  assign n6722 = po27  & n6721;
  assign n6723 = n6366 & ~n6722;
  assign n6724 = ~n6366 & n6722;
  assign n6725 = ~n6723 & ~n6724;
  assign n6726 = ~po49  & n6719;
  assign n6727 = ~n6725 & ~n6726;
  assign n6728 = ~n6720 & ~n6727;
  assign n6729 = po50  & ~n6728;
  assign n6730 = ~n6369 & ~n6370;
  assign n6731 = po27  & n6730;
  assign n6732 = n6375 & ~n6731;
  assign n6733 = ~n6375 & n6731;
  assign n6734 = ~n6732 & ~n6733;
  assign n6735 = ~po50  & ~n6720;
  assign n6736 = ~n6727 & n6735;
  assign n6737 = ~n6734 & ~n6736;
  assign n6738 = ~n6729 & ~n6737;
  assign n6739 = po51  & ~n6738;
  assign n6740 = ~n6378 & ~n6380;
  assign n6741 = po27  & n6740;
  assign n6742 = n6385 & ~n6741;
  assign n6743 = ~n6385 & n6741;
  assign n6744 = ~n6742 & ~n6743;
  assign n6745 = ~po51  & n6738;
  assign n6746 = ~n6744 & ~n6745;
  assign n6747 = ~n6739 & ~n6746;
  assign n6748 = po52  & ~n6747;
  assign n6749 = ~po52  & ~n6739;
  assign n6750 = ~n6746 & n6749;
  assign n6751 = ~n6388 & po27 ;
  assign n6752 = ~n6394 & n6751;
  assign n6753 = n6393 & ~n6752;
  assign n6754 = n6395 & n6751;
  assign n6755 = ~n6753 & ~n6754;
  assign n6756 = ~n6750 & n6755;
  assign n6757 = ~n6748 & ~n6756;
  assign n6758 = po53  & ~n6757;
  assign n6759 = ~n6397 & ~n6399;
  assign n6760 = po27  & n6759;
  assign n6761 = n6404 & ~n6760;
  assign n6762 = ~n6404 & n6760;
  assign n6763 = ~n6761 & ~n6762;
  assign n6764 = ~po53  & n6757;
  assign n6765 = ~n6763 & ~n6764;
  assign n6766 = ~n6758 & ~n6765;
  assign n6767 = po54  & ~n6766;
  assign n6768 = ~n6407 & ~n6408;
  assign n6769 = po27  & n6768;
  assign n6770 = n6413 & ~n6769;
  assign n6771 = ~n6413 & n6769;
  assign n6772 = ~n6770 & ~n6771;
  assign n6773 = ~po54  & ~n6758;
  assign n6774 = ~n6765 & n6773;
  assign n6775 = ~n6772 & ~n6774;
  assign n6776 = ~n6767 & ~n6775;
  assign n6777 = po55  & ~n6776;
  assign n6778 = ~n6416 & ~n6418;
  assign n6779 = po27  & n6778;
  assign n6780 = n6423 & ~n6779;
  assign n6781 = ~n6423 & n6779;
  assign n6782 = ~n6780 & ~n6781;
  assign n6783 = ~po55  & n6776;
  assign n6784 = ~n6782 & ~n6783;
  assign n6785 = ~n6777 & ~n6784;
  assign n6786 = po56  & ~n6785;
  assign n6787 = ~po56  & ~n6777;
  assign n6788 = ~n6784 & n6787;
  assign n6789 = ~n6426 & po27 ;
  assign n6790 = ~n6432 & n6789;
  assign n6791 = n6431 & ~n6790;
  assign n6792 = n6433 & n6789;
  assign n6793 = ~n6791 & ~n6792;
  assign n6794 = ~n6788 & n6793;
  assign n6795 = ~n6786 & ~n6794;
  assign n6796 = po57  & ~n6795;
  assign n6797 = ~n6435 & ~n6437;
  assign n6798 = po27  & n6797;
  assign n6799 = n6442 & ~n6798;
  assign n6800 = ~n6442 & n6798;
  assign n6801 = ~n6799 & ~n6800;
  assign n6802 = ~po57  & n6795;
  assign n6803 = ~n6801 & ~n6802;
  assign n6804 = ~n6796 & ~n6803;
  assign n6805 = po58  & ~n6804;
  assign n6806 = ~n6445 & ~n6446;
  assign n6807 = po27  & n6806;
  assign n6808 = n6451 & ~n6807;
  assign n6809 = ~n6451 & n6807;
  assign n6810 = ~n6808 & ~n6809;
  assign n6811 = ~po58  & ~n6796;
  assign n6812 = ~n6803 & n6811;
  assign n6813 = ~n6810 & ~n6812;
  assign n6814 = ~n6805 & ~n6813;
  assign n6815 = po59  & ~n6814;
  assign n6816 = ~n6454 & ~n6456;
  assign n6817 = po27  & n6816;
  assign n6818 = n6461 & ~n6817;
  assign n6819 = ~n6461 & n6817;
  assign n6820 = ~n6818 & ~n6819;
  assign n6821 = ~po59  & n6814;
  assign n6822 = ~n6820 & ~n6821;
  assign n6823 = ~n6815 & ~n6822;
  assign n6824 = po60  & ~n6823;
  assign n6825 = ~po60  & ~n6815;
  assign n6826 = ~n6822 & n6825;
  assign n6827 = ~n6464 & po27 ;
  assign n6828 = ~n6470 & n6827;
  assign n6829 = n6469 & ~n6828;
  assign n6830 = n6471 & n6827;
  assign n6831 = ~n6829 & ~n6830;
  assign n6832 = ~n6826 & n6831;
  assign n6833 = ~n6824 & ~n6832;
  assign n6834 = po61  & ~n6833;
  assign n6835 = ~n6473 & ~n6475;
  assign n6836 = po27  & n6835;
  assign n6837 = n6480 & ~n6836;
  assign n6838 = ~n6480 & n6836;
  assign n6839 = ~n6837 & ~n6838;
  assign n6840 = ~po61  & n6833;
  assign n6841 = ~n6839 & ~n6840;
  assign n6842 = ~n6834 & ~n6841;
  assign n6843 = po62  & ~n6842;
  assign n6844 = ~n6483 & ~n6484;
  assign n6845 = po27  & n6844;
  assign n6846 = n6489 & ~n6845;
  assign n6847 = ~n6489 & n6845;
  assign n6848 = ~n6846 & ~n6847;
  assign n6849 = ~po62  & ~n6834;
  assign n6850 = ~n6841 & n6849;
  assign n6851 = ~n6848 & ~n6850;
  assign n6852 = ~n6843 & ~n6851;
  assign n6853 = ~n6492 & ~n6494;
  assign n6854 = po27  & n6853;
  assign n6855 = n6499 & ~n6854;
  assign n6856 = ~n6499 & n6854;
  assign n6857 = ~n6855 & ~n6856;
  assign n6858 = n6501 & po27 ;
  assign n6859 = ~n6506 & ~n6858;
  assign n6860 = ~n6514 & ~n6859;
  assign n6861 = po27  & ~n6860;
  assign n6862 = ~n6857 & ~n6861;
  assign n6863 = ~n6852 & n6862;
  assign n6864 = ~po63  & ~n6863;
  assign n6865 = n6852 & n6857;
  assign n6866 = po63  & n6860;
  assign n6867 = ~n6865 & ~n6866;
  assign po26  = n6864 | ~n6867;
  assign n6869 = ~n6612 & po26 ;
  assign n6870 = ~n6611 & n6869;
  assign n6871 = n6522 & ~n6870;
  assign n6872 = n6613 & n6869;
  assign n6873 = ~n6871 & ~n6872;
  assign n6874 = ~n6601 & ~n6608;
  assign n6875 = po26  & n6874;
  assign n6876 = n6606 & ~n6875;
  assign n6877 = ~n6606 & n6875;
  assign n6878 = ~n6876 & ~n6877;
  assign n6879 = pi52  & po26 ;
  assign n6880 = ~pi50  & ~pi51 ;
  assign n6881 = ~pi52  & n6880;
  assign n6882 = ~n6879 & ~n6881;
  assign n6883 = po27  & ~n6882;
  assign n6884 = ~pi52  & po26 ;
  assign n6885 = pi53  & ~n6884;
  assign n6886 = ~pi53  & n6884;
  assign n6887 = ~n6885 & ~n6886;
  assign n6888 = ~po27  & n6882;
  assign n6889 = n6887 & ~n6888;
  assign n6890 = ~n6883 & ~n6889;
  assign n6891 = po28  & ~n6890;
  assign n6892 = ~po28  & ~n6883;
  assign n6893 = ~n6889 & n6892;
  assign n6894 = po27  & ~po26 ;
  assign n6895 = ~n6886 & ~n6894;
  assign n6896 = pi54  & ~n6895;
  assign n6897 = ~pi54  & n6895;
  assign n6898 = ~n6896 & ~n6897;
  assign n6899 = ~n6893 & ~n6898;
  assign n6900 = ~n6891 & ~n6899;
  assign n6901 = po29  & ~n6900;
  assign n6902 = ~po29  & n6900;
  assign n6903 = ~n6527 & ~n6528;
  assign n6904 = po26  & n6903;
  assign n6905 = n6532 & ~n6904;
  assign n6906 = ~n6532 & n6904;
  assign n6907 = ~n6905 & ~n6906;
  assign n6908 = ~n6902 & ~n6907;
  assign n6909 = ~n6901 & ~n6908;
  assign n6910 = po30  & ~n6909;
  assign n6911 = ~po30  & ~n6901;
  assign n6912 = ~n6908 & n6911;
  assign n6913 = ~n6535 & po26 ;
  assign n6914 = ~n6541 & n6913;
  assign n6915 = n6540 & ~n6914;
  assign n6916 = n6542 & n6913;
  assign n6917 = ~n6915 & ~n6916;
  assign n6918 = ~n6912 & n6917;
  assign n6919 = ~n6910 & ~n6918;
  assign n6920 = po31  & ~n6919;
  assign n6921 = ~po31  & n6919;
  assign n6922 = ~n6544 & ~n6546;
  assign n6923 = po26  & n6922;
  assign n6924 = n6551 & ~n6923;
  assign n6925 = ~n6551 & n6923;
  assign n6926 = ~n6924 & ~n6925;
  assign n6927 = ~n6921 & n6926;
  assign n6928 = ~n6920 & ~n6927;
  assign n6929 = po32  & ~n6928;
  assign n6930 = ~po32  & ~n6920;
  assign n6931 = ~n6927 & n6930;
  assign n6932 = ~n6554 & po26 ;
  assign n6933 = ~n6560 & n6932;
  assign n6934 = n6559 & ~n6933;
  assign n6935 = n6561 & n6932;
  assign n6936 = ~n6934 & ~n6935;
  assign n6937 = ~n6931 & n6936;
  assign n6938 = ~n6929 & ~n6937;
  assign n6939 = po33  & ~n6938;
  assign n6940 = ~po33  & n6938;
  assign n6941 = ~n6563 & ~n6565;
  assign n6942 = po26  & n6941;
  assign n6943 = n6570 & n6942;
  assign n6944 = ~n6570 & ~n6942;
  assign n6945 = ~n6943 & ~n6944;
  assign n6946 = ~n6940 & n6945;
  assign n6947 = ~n6939 & ~n6946;
  assign n6948 = po34  & ~n6947;
  assign n6949 = ~po34  & ~n6939;
  assign n6950 = ~n6946 & n6949;
  assign n6951 = ~n6573 & po26 ;
  assign n6952 = ~n6579 & n6951;
  assign n6953 = n6578 & ~n6952;
  assign n6954 = n6580 & n6951;
  assign n6955 = ~n6953 & ~n6954;
  assign n6956 = ~n6950 & n6955;
  assign n6957 = ~n6948 & ~n6956;
  assign n6958 = po35  & ~n6957;
  assign n6959 = ~po35  & n6957;
  assign n6960 = ~n6582 & ~n6584;
  assign n6961 = po26  & n6960;
  assign n6962 = ~n6589 & ~n6961;
  assign n6963 = n6589 & n6961;
  assign n6964 = ~n6962 & ~n6963;
  assign n6965 = ~n6959 & n6964;
  assign n6966 = ~n6958 & ~n6965;
  assign n6967 = po36  & ~n6966;
  assign n6968 = ~n6592 & ~n6599;
  assign n6969 = po26  & n6968;
  assign n6970 = n6597 & ~n6969;
  assign n6971 = ~n6597 & n6969;
  assign n6972 = ~n6970 & ~n6971;
  assign n6973 = ~po36  & ~n6958;
  assign n6974 = ~n6965 & n6973;
  assign n6975 = ~n6972 & ~n6974;
  assign n6976 = ~n6967 & ~n6975;
  assign n6977 = ~po37  & n6976;
  assign n6978 = ~n6878 & ~n6977;
  assign n6979 = po37  & ~n6976;
  assign n6980 = ~po38  & ~n6979;
  assign n6981 = ~n6978 & n6980;
  assign n6982 = ~n6978 & ~n6979;
  assign n6983 = po38  & ~n6982;
  assign n6984 = n6873 & ~n6981;
  assign n6985 = ~n6983 & ~n6984;
  assign n6986 = po39  & ~n6985;
  assign n6987 = ~n6615 & ~n6617;
  assign n6988 = po26  & n6987;
  assign n6989 = n6622 & ~n6988;
  assign n6990 = ~n6622 & n6988;
  assign n6991 = ~n6989 & ~n6990;
  assign n6992 = ~po39  & n6985;
  assign n6993 = ~n6991 & ~n6992;
  assign n6994 = ~n6986 & ~n6993;
  assign n6995 = po40  & ~n6994;
  assign n6996 = ~po40  & ~n6986;
  assign n6997 = ~n6993 & n6996;
  assign n6998 = ~n6625 & po26 ;
  assign n6999 = ~n6631 & n6998;
  assign n7000 = n6630 & ~n6999;
  assign n7001 = n6632 & n6998;
  assign n7002 = ~n7000 & ~n7001;
  assign n7003 = ~n6997 & n7002;
  assign n7004 = ~n6995 & ~n7003;
  assign n7005 = po41  & ~n7004;
  assign n7006 = ~n6634 & ~n6636;
  assign n7007 = po26  & n7006;
  assign n7008 = n6641 & ~n7007;
  assign n7009 = ~n6641 & n7007;
  assign n7010 = ~n7008 & ~n7009;
  assign n7011 = ~po41  & n7004;
  assign n7012 = ~n7010 & ~n7011;
  assign n7013 = ~n7005 & ~n7012;
  assign n7014 = po42  & ~n7013;
  assign n7015 = ~po42  & ~n7005;
  assign n7016 = ~n7012 & n7015;
  assign n7017 = ~n6644 & po26 ;
  assign n7018 = ~n6650 & n7017;
  assign n7019 = n6649 & ~n7018;
  assign n7020 = n6651 & n7017;
  assign n7021 = ~n7019 & ~n7020;
  assign n7022 = ~n7016 & n7021;
  assign n7023 = ~n7014 & ~n7022;
  assign n7024 = po43  & ~n7023;
  assign n7025 = ~po43  & n7023;
  assign n7026 = ~n6653 & po26 ;
  assign n7027 = ~n6660 & n7026;
  assign n7028 = n6658 & ~n7027;
  assign n7029 = n6661 & n7026;
  assign n7030 = ~n7028 & ~n7029;
  assign n7031 = ~n7025 & n7030;
  assign n7032 = ~n7024 & ~n7031;
  assign n7033 = po44  & ~n7032;
  assign n7034 = ~po44  & ~n7024;
  assign n7035 = ~n7031 & n7034;
  assign n7036 = ~n6663 & po26 ;
  assign n7037 = ~n6669 & n7036;
  assign n7038 = n6668 & ~n7037;
  assign n7039 = n6670 & n7036;
  assign n7040 = ~n7038 & ~n7039;
  assign n7041 = ~n7035 & n7040;
  assign n7042 = ~n7033 & ~n7041;
  assign n7043 = po45  & ~n7042;
  assign n7044 = ~n6672 & ~n6674;
  assign n7045 = po26  & n7044;
  assign n7046 = n6679 & ~n7045;
  assign n7047 = ~n6679 & n7045;
  assign n7048 = ~n7046 & ~n7047;
  assign n7049 = ~po45  & n7042;
  assign n7050 = ~n7048 & ~n7049;
  assign n7051 = ~n7043 & ~n7050;
  assign n7052 = po46  & ~n7051;
  assign n7053 = ~po46  & ~n7043;
  assign n7054 = ~n7050 & n7053;
  assign n7055 = ~n6682 & po26 ;
  assign n7056 = ~n6688 & n7055;
  assign n7057 = n6687 & ~n7056;
  assign n7058 = n6689 & n7055;
  assign n7059 = ~n7057 & ~n7058;
  assign n7060 = ~n7054 & n7059;
  assign n7061 = ~n7052 & ~n7060;
  assign n7062 = po47  & ~n7061;
  assign n7063 = ~po47  & n7061;
  assign n7064 = ~n6691 & po26 ;
  assign n7065 = ~n6698 & n7064;
  assign n7066 = n6696 & ~n7065;
  assign n7067 = n6699 & n7064;
  assign n7068 = ~n7066 & ~n7067;
  assign n7069 = ~n7063 & n7068;
  assign n7070 = ~n7062 & ~n7069;
  assign n7071 = po48  & ~n7070;
  assign n7072 = ~po48  & ~n7062;
  assign n7073 = ~n7069 & n7072;
  assign n7074 = ~n6701 & po26 ;
  assign n7075 = ~n6707 & n7074;
  assign n7076 = n6706 & ~n7075;
  assign n7077 = n6708 & n7074;
  assign n7078 = ~n7076 & ~n7077;
  assign n7079 = ~n7073 & n7078;
  assign n7080 = ~n7071 & ~n7079;
  assign n7081 = po49  & ~n7080;
  assign n7082 = ~n6710 & ~n6712;
  assign n7083 = po26  & n7082;
  assign n7084 = n6717 & ~n7083;
  assign n7085 = ~n6717 & n7083;
  assign n7086 = ~n7084 & ~n7085;
  assign n7087 = ~po49  & n7080;
  assign n7088 = ~n7086 & ~n7087;
  assign n7089 = ~n7081 & ~n7088;
  assign n7090 = po50  & ~n7089;
  assign n7091 = ~po50  & ~n7081;
  assign n7092 = ~n7088 & n7091;
  assign n7093 = ~n6720 & po26 ;
  assign n7094 = ~n6726 & n7093;
  assign n7095 = n6725 & ~n7094;
  assign n7096 = n6727 & n7093;
  assign n7097 = ~n7095 & ~n7096;
  assign n7098 = ~n7092 & n7097;
  assign n7099 = ~n7090 & ~n7098;
  assign n7100 = po51  & ~n7099;
  assign n7101 = ~po51  & n7099;
  assign n7102 = ~n6729 & po26 ;
  assign n7103 = ~n6736 & n7102;
  assign n7104 = n6734 & ~n7103;
  assign n7105 = n6737 & n7102;
  assign n7106 = ~n7104 & ~n7105;
  assign n7107 = ~n7101 & n7106;
  assign n7108 = ~n7100 & ~n7107;
  assign n7109 = po52  & ~n7108;
  assign n7110 = ~po52  & ~n7100;
  assign n7111 = ~n7107 & n7110;
  assign n7112 = ~n6739 & po26 ;
  assign n7113 = ~n6745 & n7112;
  assign n7114 = n6744 & ~n7113;
  assign n7115 = n6746 & n7112;
  assign n7116 = ~n7114 & ~n7115;
  assign n7117 = ~n7111 & n7116;
  assign n7118 = ~n7109 & ~n7117;
  assign n7119 = po53  & ~n7118;
  assign n7120 = ~n6748 & ~n6750;
  assign n7121 = po26  & n7120;
  assign n7122 = n6755 & ~n7121;
  assign n7123 = ~n6755 & n7121;
  assign n7124 = ~n7122 & ~n7123;
  assign n7125 = ~po53  & n7118;
  assign n7126 = ~n7124 & ~n7125;
  assign n7127 = ~n7119 & ~n7126;
  assign n7128 = po54  & ~n7127;
  assign n7129 = ~po54  & ~n7119;
  assign n7130 = ~n7126 & n7129;
  assign n7131 = ~n6758 & po26 ;
  assign n7132 = ~n6764 & n7131;
  assign n7133 = n6763 & ~n7132;
  assign n7134 = n6765 & n7131;
  assign n7135 = ~n7133 & ~n7134;
  assign n7136 = ~n7130 & n7135;
  assign n7137 = ~n7128 & ~n7136;
  assign n7138 = po55  & ~n7137;
  assign n7139 = ~po55  & n7137;
  assign n7140 = ~n6767 & po26 ;
  assign n7141 = ~n6774 & n7140;
  assign n7142 = n6772 & ~n7141;
  assign n7143 = n6775 & n7140;
  assign n7144 = ~n7142 & ~n7143;
  assign n7145 = ~n7139 & n7144;
  assign n7146 = ~n7138 & ~n7145;
  assign n7147 = po56  & ~n7146;
  assign n7148 = ~po56  & ~n7138;
  assign n7149 = ~n7145 & n7148;
  assign n7150 = ~n6777 & po26 ;
  assign n7151 = ~n6783 & n7150;
  assign n7152 = n6782 & ~n7151;
  assign n7153 = n6784 & n7150;
  assign n7154 = ~n7152 & ~n7153;
  assign n7155 = ~n7149 & n7154;
  assign n7156 = ~n7147 & ~n7155;
  assign n7157 = po57  & ~n7156;
  assign n7158 = ~n6786 & ~n6788;
  assign n7159 = po26  & n7158;
  assign n7160 = n6793 & ~n7159;
  assign n7161 = ~n6793 & n7159;
  assign n7162 = ~n7160 & ~n7161;
  assign n7163 = ~po57  & n7156;
  assign n7164 = ~n7162 & ~n7163;
  assign n7165 = ~n7157 & ~n7164;
  assign n7166 = po58  & ~n7165;
  assign n7167 = ~po58  & ~n7157;
  assign n7168 = ~n7164 & n7167;
  assign n7169 = ~n6796 & po26 ;
  assign n7170 = ~n6802 & n7169;
  assign n7171 = n6801 & ~n7170;
  assign n7172 = n6803 & n7169;
  assign n7173 = ~n7171 & ~n7172;
  assign n7174 = ~n7168 & n7173;
  assign n7175 = ~n7166 & ~n7174;
  assign n7176 = po59  & ~n7175;
  assign n7177 = ~po59  & n7175;
  assign n7178 = ~n6805 & po26 ;
  assign n7179 = ~n6812 & n7178;
  assign n7180 = n6810 & ~n7179;
  assign n7181 = n6813 & n7178;
  assign n7182 = ~n7180 & ~n7181;
  assign n7183 = ~n7177 & n7182;
  assign n7184 = ~n7176 & ~n7183;
  assign n7185 = po60  & ~n7184;
  assign n7186 = ~po60  & ~n7176;
  assign n7187 = ~n7183 & n7186;
  assign n7188 = ~n6815 & po26 ;
  assign n7189 = ~n6821 & n7188;
  assign n7190 = n6820 & ~n7189;
  assign n7191 = n6822 & n7188;
  assign n7192 = ~n7190 & ~n7191;
  assign n7193 = ~n7187 & n7192;
  assign n7194 = ~n7185 & ~n7193;
  assign n7195 = po61  & ~n7194;
  assign n7196 = ~n6824 & ~n6826;
  assign n7197 = po26  & n7196;
  assign n7198 = n6831 & ~n7197;
  assign n7199 = ~n6831 & n7197;
  assign n7200 = ~n7198 & ~n7199;
  assign n7201 = ~po61  & n7194;
  assign n7202 = ~n7200 & ~n7201;
  assign n7203 = ~n7195 & ~n7202;
  assign n7204 = po62  & ~n7203;
  assign n7205 = ~po62  & ~n7195;
  assign n7206 = ~n7202 & n7205;
  assign n7207 = ~n6834 & po26 ;
  assign n7208 = ~n6840 & n7207;
  assign n7209 = n6839 & ~n7208;
  assign n7210 = n6841 & n7207;
  assign n7211 = ~n7209 & ~n7210;
  assign n7212 = ~n7206 & n7211;
  assign n7213 = ~n7204 & ~n7212;
  assign n7214 = n6852 & po26 ;
  assign n7215 = ~n6857 & ~n7214;
  assign n7216 = ~n6865 & ~n7215;
  assign n7217 = po26  & ~n7216;
  assign n7218 = ~n6843 & po26 ;
  assign n7219 = ~n6850 & n7218;
  assign n7220 = n6848 & ~n7219;
  assign n7221 = n6851 & n7218;
  assign n7222 = ~n7220 & ~n7221;
  assign n7223 = ~n7217 & n7222;
  assign n7224 = ~n7213 & n7223;
  assign n7225 = ~po63  & ~n7224;
  assign n7226 = n7213 & ~n7222;
  assign n7227 = po63  & n7216;
  assign n7228 = ~n7226 & ~n7227;
  assign po25  = n7225 | ~n7228;
  assign n7230 = ~n6981 & ~n6983;
  assign n7231 = po25  & n7230;
  assign n7232 = n6873 & ~n7231;
  assign n7233 = ~n6873 & n7231;
  assign n7234 = ~n7232 & ~n7233;
  assign n7235 = pi50  & po25 ;
  assign n7236 = ~pi48  & ~pi49 ;
  assign n7237 = ~pi50  & n7236;
  assign n7238 = ~n7235 & ~n7237;
  assign n7239 = po26  & ~n7238;
  assign n7240 = ~po26  & n7238;
  assign n7241 = ~pi50  & po25 ;
  assign n7242 = pi51  & ~n7241;
  assign n7243 = ~pi51  & n7241;
  assign n7244 = ~n7242 & ~n7243;
  assign n7245 = ~n7240 & n7244;
  assign n7246 = ~n7239 & ~n7245;
  assign n7247 = po27  & ~n7246;
  assign n7248 = po26  & ~po25 ;
  assign n7249 = ~n7243 & ~n7248;
  assign n7250 = pi52  & ~n7249;
  assign n7251 = ~pi52  & n7249;
  assign n7252 = ~n7250 & ~n7251;
  assign n7253 = ~po27  & n7246;
  assign n7254 = ~n7252 & ~n7253;
  assign n7255 = ~n7247 & ~n7254;
  assign n7256 = po28  & ~n7255;
  assign n7257 = ~po28  & ~n7247;
  assign n7258 = ~n7254 & n7257;
  assign n7259 = ~n6883 & ~n6888;
  assign n7260 = po25  & n7259;
  assign n7261 = n6887 & ~n7260;
  assign n7262 = ~n6887 & n7260;
  assign n7263 = ~n7261 & ~n7262;
  assign n7264 = ~n7258 & ~n7263;
  assign n7265 = ~n7256 & ~n7264;
  assign n7266 = po29  & ~n7265;
  assign n7267 = ~n6891 & ~n6893;
  assign n7268 = po25  & n7267;
  assign n7269 = ~n6898 & ~n7268;
  assign n7270 = n6898 & n7268;
  assign n7271 = ~n7269 & ~n7270;
  assign n7272 = ~po29  & n7265;
  assign n7273 = ~n7271 & ~n7272;
  assign n7274 = ~n7266 & ~n7273;
  assign n7275 = po30  & ~n7274;
  assign n7276 = ~po30  & ~n7266;
  assign n7277 = ~n7273 & n7276;
  assign n7278 = ~n6901 & ~n6902;
  assign n7279 = po25  & n7278;
  assign n7280 = n6907 & ~n7279;
  assign n7281 = ~n6907 & n7279;
  assign n7282 = ~n7280 & ~n7281;
  assign n7283 = ~n7277 & n7282;
  assign n7284 = ~n7275 & ~n7283;
  assign n7285 = po31  & ~n7284;
  assign n7286 = ~n6910 & ~n6912;
  assign n7287 = po25  & n7286;
  assign n7288 = n6917 & ~n7287;
  assign n7289 = ~n6917 & n7287;
  assign n7290 = ~n7288 & ~n7289;
  assign n7291 = ~po31  & n7284;
  assign n7292 = ~n7290 & ~n7291;
  assign n7293 = ~n7285 & ~n7292;
  assign n7294 = po32  & ~n7293;
  assign n7295 = ~po32  & ~n7285;
  assign n7296 = ~n7292 & n7295;
  assign n7297 = ~n6920 & ~n6921;
  assign n7298 = po25  & n7297;
  assign n7299 = n6926 & n7298;
  assign n7300 = ~n6926 & ~n7298;
  assign n7301 = ~n7299 & ~n7300;
  assign n7302 = ~n7296 & n7301;
  assign n7303 = ~n7294 & ~n7302;
  assign n7304 = po33  & ~n7303;
  assign n7305 = ~n6929 & ~n6931;
  assign n7306 = po25  & n7305;
  assign n7307 = n6936 & ~n7306;
  assign n7308 = ~n6936 & n7306;
  assign n7309 = ~n7307 & ~n7308;
  assign n7310 = ~po33  & n7303;
  assign n7311 = ~n7309 & ~n7310;
  assign n7312 = ~n7304 & ~n7311;
  assign n7313 = po34  & ~n7312;
  assign n7314 = ~po34  & ~n7304;
  assign n7315 = ~n7311 & n7314;
  assign n7316 = ~n6939 & ~n6940;
  assign n7317 = po25  & n7316;
  assign n7318 = ~n6945 & ~n7317;
  assign n7319 = n6945 & n7317;
  assign n7320 = ~n7318 & ~n7319;
  assign n7321 = ~n7315 & n7320;
  assign n7322 = ~n7313 & ~n7321;
  assign n7323 = po35  & ~n7322;
  assign n7324 = ~n6948 & ~n6950;
  assign n7325 = po25  & n7324;
  assign n7326 = n6955 & ~n7325;
  assign n7327 = ~n6955 & n7325;
  assign n7328 = ~n7326 & ~n7327;
  assign n7329 = ~po35  & n7322;
  assign n7330 = ~n7328 & ~n7329;
  assign n7331 = ~n7323 & ~n7330;
  assign n7332 = po36  & ~n7331;
  assign n7333 = ~n6958 & ~n6959;
  assign n7334 = po25  & n7333;
  assign n7335 = n6964 & ~n7334;
  assign n7336 = ~n6964 & n7334;
  assign n7337 = ~n7335 & ~n7336;
  assign n7338 = ~po36  & ~n7323;
  assign n7339 = ~n7330 & n7338;
  assign n7340 = ~n7337 & ~n7339;
  assign n7341 = ~n7332 & ~n7340;
  assign n7342 = ~po37  & n7341;
  assign n7343 = ~n6967 & po25 ;
  assign n7344 = ~n6974 & n7343;
  assign n7345 = n6972 & ~n7344;
  assign n7346 = n6975 & n7343;
  assign n7347 = ~n7345 & ~n7346;
  assign n7348 = ~n7342 & n7347;
  assign n7349 = po37  & ~n7341;
  assign n7350 = ~n7348 & ~n7349;
  assign n7351 = po38  & ~n7350;
  assign n7352 = ~po38  & ~n7349;
  assign n7353 = ~n7348 & n7352;
  assign n7354 = ~n6977 & ~n6979;
  assign n7355 = po25  & n7354;
  assign n7356 = n6878 & n7355;
  assign n7357 = ~n6878 & ~n7355;
  assign n7358 = ~n7356 & ~n7357;
  assign n7359 = ~n7353 & ~n7358;
  assign n7360 = ~n7351 & ~n7359;
  assign n7361 = ~po39  & n7360;
  assign n7362 = po39  & ~n7360;
  assign n7363 = ~n7234 & ~n7361;
  assign n7364 = ~n7362 & ~n7363;
  assign n7365 = po40  & ~n7364;
  assign n7366 = ~po40  & ~n7362;
  assign n7367 = ~n7363 & n7366;
  assign n7368 = ~n6986 & po25 ;
  assign n7369 = ~n6992 & n7368;
  assign n7370 = n6991 & ~n7369;
  assign n7371 = n6993 & n7368;
  assign n7372 = ~n7370 & ~n7371;
  assign n7373 = ~n7367 & n7372;
  assign n7374 = ~n7365 & ~n7373;
  assign n7375 = po41  & ~n7374;
  assign n7376 = ~n6995 & ~n6997;
  assign n7377 = po25  & n7376;
  assign n7378 = n7002 & ~n7377;
  assign n7379 = ~n7002 & n7377;
  assign n7380 = ~n7378 & ~n7379;
  assign n7381 = ~po41  & n7374;
  assign n7382 = ~n7380 & ~n7381;
  assign n7383 = ~n7375 & ~n7382;
  assign n7384 = po42  & ~n7383;
  assign n7385 = ~po42  & ~n7375;
  assign n7386 = ~n7382 & n7385;
  assign n7387 = ~n7005 & po25 ;
  assign n7388 = ~n7011 & n7387;
  assign n7389 = n7010 & ~n7388;
  assign n7390 = n7012 & n7387;
  assign n7391 = ~n7389 & ~n7390;
  assign n7392 = ~n7386 & n7391;
  assign n7393 = ~n7384 & ~n7392;
  assign n7394 = po43  & ~n7393;
  assign n7395 = ~n7014 & ~n7016;
  assign n7396 = po25  & n7395;
  assign n7397 = n7021 & ~n7396;
  assign n7398 = ~n7021 & n7396;
  assign n7399 = ~n7397 & ~n7398;
  assign n7400 = ~po43  & n7393;
  assign n7401 = ~n7399 & ~n7400;
  assign n7402 = ~n7394 & ~n7401;
  assign n7403 = po44  & ~n7402;
  assign n7404 = ~n7024 & ~n7025;
  assign n7405 = po25  & n7404;
  assign n7406 = n7030 & ~n7405;
  assign n7407 = ~n7030 & n7405;
  assign n7408 = ~n7406 & ~n7407;
  assign n7409 = ~po44  & ~n7394;
  assign n7410 = ~n7401 & n7409;
  assign n7411 = ~n7408 & ~n7410;
  assign n7412 = ~n7403 & ~n7411;
  assign n7413 = po45  & ~n7412;
  assign n7414 = ~n7033 & ~n7035;
  assign n7415 = po25  & n7414;
  assign n7416 = n7040 & ~n7415;
  assign n7417 = ~n7040 & n7415;
  assign n7418 = ~n7416 & ~n7417;
  assign n7419 = ~po45  & n7412;
  assign n7420 = ~n7418 & ~n7419;
  assign n7421 = ~n7413 & ~n7420;
  assign n7422 = po46  & ~n7421;
  assign n7423 = ~po46  & ~n7413;
  assign n7424 = ~n7420 & n7423;
  assign n7425 = ~n7043 & po25 ;
  assign n7426 = ~n7049 & n7425;
  assign n7427 = n7048 & ~n7426;
  assign n7428 = n7050 & n7425;
  assign n7429 = ~n7427 & ~n7428;
  assign n7430 = ~n7424 & n7429;
  assign n7431 = ~n7422 & ~n7430;
  assign n7432 = po47  & ~n7431;
  assign n7433 = ~n7052 & ~n7054;
  assign n7434 = po25  & n7433;
  assign n7435 = n7059 & ~n7434;
  assign n7436 = ~n7059 & n7434;
  assign n7437 = ~n7435 & ~n7436;
  assign n7438 = ~po47  & n7431;
  assign n7439 = ~n7437 & ~n7438;
  assign n7440 = ~n7432 & ~n7439;
  assign n7441 = po48  & ~n7440;
  assign n7442 = ~n7062 & ~n7063;
  assign n7443 = po25  & n7442;
  assign n7444 = n7068 & ~n7443;
  assign n7445 = ~n7068 & n7443;
  assign n7446 = ~n7444 & ~n7445;
  assign n7447 = ~po48  & ~n7432;
  assign n7448 = ~n7439 & n7447;
  assign n7449 = ~n7446 & ~n7448;
  assign n7450 = ~n7441 & ~n7449;
  assign n7451 = po49  & ~n7450;
  assign n7452 = ~n7071 & ~n7073;
  assign n7453 = po25  & n7452;
  assign n7454 = n7078 & ~n7453;
  assign n7455 = ~n7078 & n7453;
  assign n7456 = ~n7454 & ~n7455;
  assign n7457 = ~po49  & n7450;
  assign n7458 = ~n7456 & ~n7457;
  assign n7459 = ~n7451 & ~n7458;
  assign n7460 = po50  & ~n7459;
  assign n7461 = ~po50  & ~n7451;
  assign n7462 = ~n7458 & n7461;
  assign n7463 = ~n7081 & po25 ;
  assign n7464 = ~n7087 & n7463;
  assign n7465 = n7086 & ~n7464;
  assign n7466 = n7088 & n7463;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = ~n7462 & n7467;
  assign n7469 = ~n7460 & ~n7468;
  assign n7470 = po51  & ~n7469;
  assign n7471 = ~n7090 & ~n7092;
  assign n7472 = po25  & n7471;
  assign n7473 = n7097 & ~n7472;
  assign n7474 = ~n7097 & n7472;
  assign n7475 = ~n7473 & ~n7474;
  assign n7476 = ~po51  & n7469;
  assign n7477 = ~n7475 & ~n7476;
  assign n7478 = ~n7470 & ~n7477;
  assign n7479 = po52  & ~n7478;
  assign n7480 = ~n7100 & ~n7101;
  assign n7481 = po25  & n7480;
  assign n7482 = n7106 & ~n7481;
  assign n7483 = ~n7106 & n7481;
  assign n7484 = ~n7482 & ~n7483;
  assign n7485 = ~po52  & ~n7470;
  assign n7486 = ~n7477 & n7485;
  assign n7487 = ~n7484 & ~n7486;
  assign n7488 = ~n7479 & ~n7487;
  assign n7489 = po53  & ~n7488;
  assign n7490 = ~n7109 & ~n7111;
  assign n7491 = po25  & n7490;
  assign n7492 = n7116 & ~n7491;
  assign n7493 = ~n7116 & n7491;
  assign n7494 = ~n7492 & ~n7493;
  assign n7495 = ~po53  & n7488;
  assign n7496 = ~n7494 & ~n7495;
  assign n7497 = ~n7489 & ~n7496;
  assign n7498 = po54  & ~n7497;
  assign n7499 = ~po54  & ~n7489;
  assign n7500 = ~n7496 & n7499;
  assign n7501 = ~n7119 & po25 ;
  assign n7502 = ~n7125 & n7501;
  assign n7503 = n7124 & ~n7502;
  assign n7504 = n7126 & n7501;
  assign n7505 = ~n7503 & ~n7504;
  assign n7506 = ~n7500 & n7505;
  assign n7507 = ~n7498 & ~n7506;
  assign n7508 = po55  & ~n7507;
  assign n7509 = ~n7128 & ~n7130;
  assign n7510 = po25  & n7509;
  assign n7511 = n7135 & ~n7510;
  assign n7512 = ~n7135 & n7510;
  assign n7513 = ~n7511 & ~n7512;
  assign n7514 = ~po55  & n7507;
  assign n7515 = ~n7513 & ~n7514;
  assign n7516 = ~n7508 & ~n7515;
  assign n7517 = po56  & ~n7516;
  assign n7518 = ~n7138 & ~n7139;
  assign n7519 = po25  & n7518;
  assign n7520 = n7144 & ~n7519;
  assign n7521 = ~n7144 & n7519;
  assign n7522 = ~n7520 & ~n7521;
  assign n7523 = ~po56  & ~n7508;
  assign n7524 = ~n7515 & n7523;
  assign n7525 = ~n7522 & ~n7524;
  assign n7526 = ~n7517 & ~n7525;
  assign n7527 = po57  & ~n7526;
  assign n7528 = ~n7147 & ~n7149;
  assign n7529 = po25  & n7528;
  assign n7530 = n7154 & ~n7529;
  assign n7531 = ~n7154 & n7529;
  assign n7532 = ~n7530 & ~n7531;
  assign n7533 = ~po57  & n7526;
  assign n7534 = ~n7532 & ~n7533;
  assign n7535 = ~n7527 & ~n7534;
  assign n7536 = po58  & ~n7535;
  assign n7537 = ~po58  & ~n7527;
  assign n7538 = ~n7534 & n7537;
  assign n7539 = ~n7157 & po25 ;
  assign n7540 = ~n7163 & n7539;
  assign n7541 = n7162 & ~n7540;
  assign n7542 = n7164 & n7539;
  assign n7543 = ~n7541 & ~n7542;
  assign n7544 = ~n7538 & n7543;
  assign n7545 = ~n7536 & ~n7544;
  assign n7546 = po59  & ~n7545;
  assign n7547 = ~n7166 & ~n7168;
  assign n7548 = po25  & n7547;
  assign n7549 = n7173 & ~n7548;
  assign n7550 = ~n7173 & n7548;
  assign n7551 = ~n7549 & ~n7550;
  assign n7552 = ~po59  & n7545;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = ~n7546 & ~n7553;
  assign n7555 = po60  & ~n7554;
  assign n7556 = ~n7176 & ~n7177;
  assign n7557 = po25  & n7556;
  assign n7558 = n7182 & ~n7557;
  assign n7559 = ~n7182 & n7557;
  assign n7560 = ~n7558 & ~n7559;
  assign n7561 = ~po60  & ~n7546;
  assign n7562 = ~n7553 & n7561;
  assign n7563 = ~n7560 & ~n7562;
  assign n7564 = ~n7555 & ~n7563;
  assign n7565 = po61  & ~n7564;
  assign n7566 = ~n7185 & ~n7187;
  assign n7567 = po25  & n7566;
  assign n7568 = n7192 & ~n7567;
  assign n7569 = ~n7192 & n7567;
  assign n7570 = ~n7568 & ~n7569;
  assign n7571 = ~po61  & n7564;
  assign n7572 = ~n7570 & ~n7571;
  assign n7573 = ~n7565 & ~n7572;
  assign n7574 = po62  & ~n7573;
  assign n7575 = ~po62  & ~n7565;
  assign n7576 = ~n7572 & n7575;
  assign n7577 = ~n7195 & po25 ;
  assign n7578 = ~n7201 & n7577;
  assign n7579 = n7200 & ~n7578;
  assign n7580 = n7202 & n7577;
  assign n7581 = ~n7579 & ~n7580;
  assign n7582 = ~n7576 & n7581;
  assign n7583 = ~n7574 & ~n7582;
  assign n7584 = n7222 & po25 ;
  assign n7585 = ~n7213 & n7584;
  assign n7586 = ~n7204 & ~n7206;
  assign n7587 = po25  & n7586;
  assign n7588 = n7211 & ~n7587;
  assign n7589 = ~n7211 & n7587;
  assign n7590 = ~n7588 & ~n7589;
  assign n7591 = ~n7226 & ~n7585;
  assign n7592 = ~n7590 & n7591;
  assign n7593 = ~n7583 & n7592;
  assign n7594 = ~po63  & ~n7593;
  assign n7595 = n7583 & n7590;
  assign n7596 = n7213 & ~n7584;
  assign n7597 = ~n7213 & n7222;
  assign n7598 = po63  & ~n7597;
  assign n7599 = ~n7596 & n7598;
  assign n7600 = ~n7595 & ~n7599;
  assign po24  = n7594 | ~n7600;
  assign n7602 = ~n7362 & po24 ;
  assign n7603 = ~n7361 & n7602;
  assign n7604 = n7234 & ~n7603;
  assign n7605 = n7363 & n7602;
  assign n7606 = ~n7604 & ~n7605;
  assign n7607 = ~n7351 & ~n7353;
  assign n7608 = po24  & n7607;
  assign n7609 = ~n7358 & ~n7608;
  assign n7610 = n7358 & n7608;
  assign n7611 = ~n7609 & ~n7610;
  assign n7612 = pi48  & po24 ;
  assign n7613 = ~pi46  & ~pi47 ;
  assign n7614 = ~pi48  & n7613;
  assign n7615 = ~n7612 & ~n7614;
  assign n7616 = po25  & ~n7615;
  assign n7617 = ~pi48  & po24 ;
  assign n7618 = pi49  & ~n7617;
  assign n7619 = ~pi49  & n7617;
  assign n7620 = ~n7618 & ~n7619;
  assign n7621 = ~po25  & n7615;
  assign n7622 = n7620 & ~n7621;
  assign n7623 = ~n7616 & ~n7622;
  assign n7624 = po26  & ~n7623;
  assign n7625 = ~po26  & ~n7616;
  assign n7626 = ~n7622 & n7625;
  assign n7627 = po25  & ~po24 ;
  assign n7628 = ~n7619 & ~n7627;
  assign n7629 = pi50  & ~n7628;
  assign n7630 = ~pi50  & n7628;
  assign n7631 = ~n7629 & ~n7630;
  assign n7632 = ~n7626 & ~n7631;
  assign n7633 = ~n7624 & ~n7632;
  assign n7634 = po27  & ~n7633;
  assign n7635 = ~po27  & n7633;
  assign n7636 = ~n7239 & ~n7240;
  assign n7637 = po24  & n7636;
  assign n7638 = n7244 & ~n7637;
  assign n7639 = ~n7244 & n7637;
  assign n7640 = ~n7638 & ~n7639;
  assign n7641 = ~n7635 & ~n7640;
  assign n7642 = ~n7634 & ~n7641;
  assign n7643 = po28  & ~n7642;
  assign n7644 = ~po28  & ~n7634;
  assign n7645 = ~n7641 & n7644;
  assign n7646 = ~n7247 & po24 ;
  assign n7647 = ~n7253 & n7646;
  assign n7648 = n7252 & ~n7647;
  assign n7649 = n7254 & n7646;
  assign n7650 = ~n7648 & ~n7649;
  assign n7651 = ~n7645 & n7650;
  assign n7652 = ~n7643 & ~n7651;
  assign n7653 = po29  & ~n7652;
  assign n7654 = ~po29  & n7652;
  assign n7655 = ~n7256 & ~n7258;
  assign n7656 = po24  & n7655;
  assign n7657 = n7263 & ~n7656;
  assign n7658 = ~n7263 & n7656;
  assign n7659 = ~n7657 & ~n7658;
  assign n7660 = ~n7654 & n7659;
  assign n7661 = ~n7653 & ~n7660;
  assign n7662 = po30  & ~n7661;
  assign n7663 = ~po30  & ~n7653;
  assign n7664 = ~n7660 & n7663;
  assign n7665 = ~n7266 & po24 ;
  assign n7666 = ~n7272 & n7665;
  assign n7667 = n7271 & ~n7666;
  assign n7668 = n7273 & n7665;
  assign n7669 = ~n7667 & ~n7668;
  assign n7670 = ~n7664 & n7669;
  assign n7671 = ~n7662 & ~n7670;
  assign n7672 = po31  & ~n7671;
  assign n7673 = ~po31  & n7671;
  assign n7674 = ~n7275 & ~n7277;
  assign n7675 = po24  & n7674;
  assign n7676 = n7282 & n7675;
  assign n7677 = ~n7282 & ~n7675;
  assign n7678 = ~n7676 & ~n7677;
  assign n7679 = ~n7673 & n7678;
  assign n7680 = ~n7672 & ~n7679;
  assign n7681 = po32  & ~n7680;
  assign n7682 = ~po32  & ~n7672;
  assign n7683 = ~n7679 & n7682;
  assign n7684 = ~n7285 & po24 ;
  assign n7685 = ~n7291 & n7684;
  assign n7686 = n7290 & ~n7685;
  assign n7687 = n7292 & n7684;
  assign n7688 = ~n7686 & ~n7687;
  assign n7689 = ~n7683 & n7688;
  assign n7690 = ~n7681 & ~n7689;
  assign n7691 = po33  & ~n7690;
  assign n7692 = ~po33  & n7690;
  assign n7693 = ~n7294 & ~n7296;
  assign n7694 = po24  & n7693;
  assign n7695 = ~n7301 & ~n7694;
  assign n7696 = n7301 & n7694;
  assign n7697 = ~n7695 & ~n7696;
  assign n7698 = ~n7692 & n7697;
  assign n7699 = ~n7691 & ~n7698;
  assign n7700 = po34  & ~n7699;
  assign n7701 = ~po34  & ~n7691;
  assign n7702 = ~n7698 & n7701;
  assign n7703 = ~n7304 & po24 ;
  assign n7704 = ~n7310 & n7703;
  assign n7705 = n7309 & ~n7704;
  assign n7706 = n7311 & n7703;
  assign n7707 = ~n7705 & ~n7706;
  assign n7708 = ~n7702 & n7707;
  assign n7709 = ~n7700 & ~n7708;
  assign n7710 = po35  & ~n7709;
  assign n7711 = ~n7313 & ~n7315;
  assign n7712 = po24  & n7711;
  assign n7713 = n7320 & ~n7712;
  assign n7714 = ~n7320 & n7712;
  assign n7715 = ~n7713 & ~n7714;
  assign n7716 = ~po35  & n7709;
  assign n7717 = ~n7715 & ~n7716;
  assign n7718 = ~n7710 & ~n7717;
  assign n7719 = po36  & ~n7718;
  assign n7720 = ~po36  & ~n7710;
  assign n7721 = ~n7717 & n7720;
  assign n7722 = ~n7323 & po24 ;
  assign n7723 = ~n7329 & n7722;
  assign n7724 = n7328 & ~n7723;
  assign n7725 = n7330 & n7722;
  assign n7726 = ~n7724 & ~n7725;
  assign n7727 = ~n7721 & n7726;
  assign n7728 = ~n7719 & ~n7727;
  assign n7729 = po37  & ~n7728;
  assign n7730 = ~po37  & n7728;
  assign n7731 = ~n7332 & po24 ;
  assign n7732 = ~n7339 & n7731;
  assign n7733 = n7337 & ~n7732;
  assign n7734 = n7340 & n7731;
  assign n7735 = ~n7733 & ~n7734;
  assign n7736 = ~n7730 & n7735;
  assign n7737 = ~n7729 & ~n7736;
  assign n7738 = po38  & ~n7737;
  assign n7739 = ~n7342 & ~n7349;
  assign n7740 = po24  & n7739;
  assign n7741 = n7347 & ~n7740;
  assign n7742 = ~n7347 & n7740;
  assign n7743 = ~n7741 & ~n7742;
  assign n7744 = ~po38  & ~n7729;
  assign n7745 = ~n7736 & n7744;
  assign n7746 = ~n7743 & ~n7745;
  assign n7747 = ~n7738 & ~n7746;
  assign n7748 = ~po39  & n7747;
  assign n7749 = ~n7611 & ~n7748;
  assign n7750 = po39  & ~n7747;
  assign n7751 = ~po40  & ~n7750;
  assign n7752 = ~n7749 & n7751;
  assign n7753 = ~n7749 & ~n7750;
  assign n7754 = po40  & ~n7753;
  assign n7755 = n7606 & ~n7752;
  assign n7756 = ~n7754 & ~n7755;
  assign n7757 = po41  & ~n7756;
  assign n7758 = ~n7365 & ~n7367;
  assign n7759 = po24  & n7758;
  assign n7760 = n7372 & ~n7759;
  assign n7761 = ~n7372 & n7759;
  assign n7762 = ~n7760 & ~n7761;
  assign n7763 = ~po41  & n7756;
  assign n7764 = ~n7762 & ~n7763;
  assign n7765 = ~n7757 & ~n7764;
  assign n7766 = po42  & ~n7765;
  assign n7767 = ~po42  & ~n7757;
  assign n7768 = ~n7764 & n7767;
  assign n7769 = ~n7375 & po24 ;
  assign n7770 = ~n7381 & n7769;
  assign n7771 = n7380 & ~n7770;
  assign n7772 = n7382 & n7769;
  assign n7773 = ~n7771 & ~n7772;
  assign n7774 = ~n7768 & n7773;
  assign n7775 = ~n7766 & ~n7774;
  assign n7776 = po43  & ~n7775;
  assign n7777 = ~n7384 & ~n7386;
  assign n7778 = po24  & n7777;
  assign n7779 = n7391 & ~n7778;
  assign n7780 = ~n7391 & n7778;
  assign n7781 = ~n7779 & ~n7780;
  assign n7782 = ~po43  & n7775;
  assign n7783 = ~n7781 & ~n7782;
  assign n7784 = ~n7776 & ~n7783;
  assign n7785 = po44  & ~n7784;
  assign n7786 = ~po44  & ~n7776;
  assign n7787 = ~n7783 & n7786;
  assign n7788 = ~n7394 & po24 ;
  assign n7789 = ~n7400 & n7788;
  assign n7790 = n7399 & ~n7789;
  assign n7791 = n7401 & n7788;
  assign n7792 = ~n7790 & ~n7791;
  assign n7793 = ~n7787 & n7792;
  assign n7794 = ~n7785 & ~n7793;
  assign n7795 = po45  & ~n7794;
  assign n7796 = ~po45  & n7794;
  assign n7797 = ~n7403 & po24 ;
  assign n7798 = ~n7410 & n7797;
  assign n7799 = n7408 & ~n7798;
  assign n7800 = n7411 & n7797;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = ~n7796 & n7801;
  assign n7803 = ~n7795 & ~n7802;
  assign n7804 = po46  & ~n7803;
  assign n7805 = ~po46  & ~n7795;
  assign n7806 = ~n7802 & n7805;
  assign n7807 = ~n7413 & po24 ;
  assign n7808 = ~n7419 & n7807;
  assign n7809 = n7418 & ~n7808;
  assign n7810 = n7420 & n7807;
  assign n7811 = ~n7809 & ~n7810;
  assign n7812 = ~n7806 & n7811;
  assign n7813 = ~n7804 & ~n7812;
  assign n7814 = po47  & ~n7813;
  assign n7815 = ~n7422 & ~n7424;
  assign n7816 = po24  & n7815;
  assign n7817 = n7429 & ~n7816;
  assign n7818 = ~n7429 & n7816;
  assign n7819 = ~n7817 & ~n7818;
  assign n7820 = ~po47  & n7813;
  assign n7821 = ~n7819 & ~n7820;
  assign n7822 = ~n7814 & ~n7821;
  assign n7823 = po48  & ~n7822;
  assign n7824 = ~po48  & ~n7814;
  assign n7825 = ~n7821 & n7824;
  assign n7826 = ~n7432 & po24 ;
  assign n7827 = ~n7438 & n7826;
  assign n7828 = n7437 & ~n7827;
  assign n7829 = n7439 & n7826;
  assign n7830 = ~n7828 & ~n7829;
  assign n7831 = ~n7825 & n7830;
  assign n7832 = ~n7823 & ~n7831;
  assign n7833 = po49  & ~n7832;
  assign n7834 = ~po49  & n7832;
  assign n7835 = ~n7441 & po24 ;
  assign n7836 = ~n7448 & n7835;
  assign n7837 = n7446 & ~n7836;
  assign n7838 = n7449 & n7835;
  assign n7839 = ~n7837 & ~n7838;
  assign n7840 = ~n7834 & n7839;
  assign n7841 = ~n7833 & ~n7840;
  assign n7842 = po50  & ~n7841;
  assign n7843 = ~po50  & ~n7833;
  assign n7844 = ~n7840 & n7843;
  assign n7845 = ~n7451 & po24 ;
  assign n7846 = ~n7457 & n7845;
  assign n7847 = n7456 & ~n7846;
  assign n7848 = n7458 & n7845;
  assign n7849 = ~n7847 & ~n7848;
  assign n7850 = ~n7844 & n7849;
  assign n7851 = ~n7842 & ~n7850;
  assign n7852 = po51  & ~n7851;
  assign n7853 = ~n7460 & ~n7462;
  assign n7854 = po24  & n7853;
  assign n7855 = n7467 & ~n7854;
  assign n7856 = ~n7467 & n7854;
  assign n7857 = ~n7855 & ~n7856;
  assign n7858 = ~po51  & n7851;
  assign n7859 = ~n7857 & ~n7858;
  assign n7860 = ~n7852 & ~n7859;
  assign n7861 = po52  & ~n7860;
  assign n7862 = ~po52  & ~n7852;
  assign n7863 = ~n7859 & n7862;
  assign n7864 = ~n7470 & po24 ;
  assign n7865 = ~n7476 & n7864;
  assign n7866 = n7475 & ~n7865;
  assign n7867 = n7477 & n7864;
  assign n7868 = ~n7866 & ~n7867;
  assign n7869 = ~n7863 & n7868;
  assign n7870 = ~n7861 & ~n7869;
  assign n7871 = po53  & ~n7870;
  assign n7872 = ~po53  & n7870;
  assign n7873 = ~n7479 & po24 ;
  assign n7874 = ~n7486 & n7873;
  assign n7875 = n7484 & ~n7874;
  assign n7876 = n7487 & n7873;
  assign n7877 = ~n7875 & ~n7876;
  assign n7878 = ~n7872 & n7877;
  assign n7879 = ~n7871 & ~n7878;
  assign n7880 = po54  & ~n7879;
  assign n7881 = ~po54  & ~n7871;
  assign n7882 = ~n7878 & n7881;
  assign n7883 = ~n7489 & po24 ;
  assign n7884 = ~n7495 & n7883;
  assign n7885 = n7494 & ~n7884;
  assign n7886 = n7496 & n7883;
  assign n7887 = ~n7885 & ~n7886;
  assign n7888 = ~n7882 & n7887;
  assign n7889 = ~n7880 & ~n7888;
  assign n7890 = po55  & ~n7889;
  assign n7891 = ~n7498 & ~n7500;
  assign n7892 = po24  & n7891;
  assign n7893 = n7505 & ~n7892;
  assign n7894 = ~n7505 & n7892;
  assign n7895 = ~n7893 & ~n7894;
  assign n7896 = ~po55  & n7889;
  assign n7897 = ~n7895 & ~n7896;
  assign n7898 = ~n7890 & ~n7897;
  assign n7899 = po56  & ~n7898;
  assign n7900 = ~po56  & ~n7890;
  assign n7901 = ~n7897 & n7900;
  assign n7902 = ~n7508 & po24 ;
  assign n7903 = ~n7514 & n7902;
  assign n7904 = n7513 & ~n7903;
  assign n7905 = n7515 & n7902;
  assign n7906 = ~n7904 & ~n7905;
  assign n7907 = ~n7901 & n7906;
  assign n7908 = ~n7899 & ~n7907;
  assign n7909 = po57  & ~n7908;
  assign n7910 = ~po57  & n7908;
  assign n7911 = ~n7517 & po24 ;
  assign n7912 = ~n7524 & n7911;
  assign n7913 = n7522 & ~n7912;
  assign n7914 = n7525 & n7911;
  assign n7915 = ~n7913 & ~n7914;
  assign n7916 = ~n7910 & n7915;
  assign n7917 = ~n7909 & ~n7916;
  assign n7918 = po58  & ~n7917;
  assign n7919 = ~po58  & ~n7909;
  assign n7920 = ~n7916 & n7919;
  assign n7921 = ~n7527 & po24 ;
  assign n7922 = ~n7533 & n7921;
  assign n7923 = n7532 & ~n7922;
  assign n7924 = n7534 & n7921;
  assign n7925 = ~n7923 & ~n7924;
  assign n7926 = ~n7920 & n7925;
  assign n7927 = ~n7918 & ~n7926;
  assign n7928 = po59  & ~n7927;
  assign n7929 = ~n7536 & ~n7538;
  assign n7930 = po24  & n7929;
  assign n7931 = n7543 & ~n7930;
  assign n7932 = ~n7543 & n7930;
  assign n7933 = ~n7931 & ~n7932;
  assign n7934 = ~po59  & n7927;
  assign n7935 = ~n7933 & ~n7934;
  assign n7936 = ~n7928 & ~n7935;
  assign n7937 = po60  & ~n7936;
  assign n7938 = ~po60  & ~n7928;
  assign n7939 = ~n7935 & n7938;
  assign n7940 = ~n7546 & po24 ;
  assign n7941 = ~n7552 & n7940;
  assign n7942 = n7551 & ~n7941;
  assign n7943 = n7553 & n7940;
  assign n7944 = ~n7942 & ~n7943;
  assign n7945 = ~n7939 & n7944;
  assign n7946 = ~n7937 & ~n7945;
  assign n7947 = po61  & ~n7946;
  assign n7948 = ~po61  & n7946;
  assign n7949 = ~n7555 & po24 ;
  assign n7950 = ~n7562 & n7949;
  assign n7951 = n7560 & ~n7950;
  assign n7952 = n7563 & n7949;
  assign n7953 = ~n7951 & ~n7952;
  assign n7954 = ~n7948 & n7953;
  assign n7955 = ~n7947 & ~n7954;
  assign n7956 = po62  & ~n7955;
  assign n7957 = ~po62  & ~n7947;
  assign n7958 = ~n7954 & n7957;
  assign n7959 = ~n7565 & po24 ;
  assign n7960 = ~n7571 & n7959;
  assign n7961 = n7570 & ~n7960;
  assign n7962 = n7572 & n7959;
  assign n7963 = ~n7961 & ~n7962;
  assign n7964 = ~n7958 & n7963;
  assign n7965 = ~n7956 & ~n7964;
  assign n7966 = ~n7574 & ~n7576;
  assign n7967 = po24  & n7966;
  assign n7968 = n7581 & ~n7967;
  assign n7969 = ~n7581 & n7967;
  assign n7970 = ~n7968 & ~n7969;
  assign n7971 = n7583 & po24 ;
  assign n7972 = ~n7590 & ~n7971;
  assign n7973 = ~n7595 & ~n7972;
  assign n7974 = po24  & ~n7973;
  assign n7975 = ~n7970 & ~n7974;
  assign n7976 = ~n7965 & n7975;
  assign n7977 = ~po63  & ~n7976;
  assign n7978 = n7965 & n7970;
  assign n7979 = po63  & n7973;
  assign n7980 = ~n7978 & ~n7979;
  assign po23  = n7977 | ~n7980;
  assign n7982 = ~n7752 & ~n7754;
  assign n7983 = po23  & n7982;
  assign n7984 = n7606 & ~n7983;
  assign n7985 = ~n7606 & n7983;
  assign n7986 = ~n7984 & ~n7985;
  assign n7987 = pi46  & po23 ;
  assign n7988 = ~pi44  & ~pi45 ;
  assign n7989 = ~pi46  & n7988;
  assign n7990 = ~n7987 & ~n7989;
  assign n7991 = po24  & ~n7990;
  assign n7992 = ~po24  & n7990;
  assign n7993 = ~pi46  & po23 ;
  assign n7994 = pi47  & ~n7993;
  assign n7995 = ~pi47  & n7993;
  assign n7996 = ~n7994 & ~n7995;
  assign n7997 = ~n7992 & n7996;
  assign n7998 = ~n7991 & ~n7997;
  assign n7999 = po25  & ~n7998;
  assign n8000 = po24  & ~po23 ;
  assign n8001 = ~n7995 & ~n8000;
  assign n8002 = pi48  & ~n8001;
  assign n8003 = ~pi48  & n8001;
  assign n8004 = ~n8002 & ~n8003;
  assign n8005 = ~po25  & n7998;
  assign n8006 = ~n8004 & ~n8005;
  assign n8007 = ~n7999 & ~n8006;
  assign n8008 = po26  & ~n8007;
  assign n8009 = ~po26  & ~n7999;
  assign n8010 = ~n8006 & n8009;
  assign n8011 = ~n7616 & ~n7621;
  assign n8012 = po23  & n8011;
  assign n8013 = n7620 & ~n8012;
  assign n8014 = ~n7620 & n8012;
  assign n8015 = ~n8013 & ~n8014;
  assign n8016 = ~n8010 & ~n8015;
  assign n8017 = ~n8008 & ~n8016;
  assign n8018 = po27  & ~n8017;
  assign n8019 = ~n7624 & ~n7626;
  assign n8020 = po23  & n8019;
  assign n8021 = ~n7631 & ~n8020;
  assign n8022 = n7631 & n8020;
  assign n8023 = ~n8021 & ~n8022;
  assign n8024 = ~po27  & n8017;
  assign n8025 = ~n8023 & ~n8024;
  assign n8026 = ~n8018 & ~n8025;
  assign n8027 = po28  & ~n8026;
  assign n8028 = ~po28  & ~n8018;
  assign n8029 = ~n8025 & n8028;
  assign n8030 = ~n7634 & ~n7635;
  assign n8031 = po23  & n8030;
  assign n8032 = n7640 & ~n8031;
  assign n8033 = ~n7640 & n8031;
  assign n8034 = ~n8032 & ~n8033;
  assign n8035 = ~n8029 & n8034;
  assign n8036 = ~n8027 & ~n8035;
  assign n8037 = po29  & ~n8036;
  assign n8038 = ~n7643 & ~n7645;
  assign n8039 = po23  & n8038;
  assign n8040 = n7650 & ~n8039;
  assign n8041 = ~n7650 & n8039;
  assign n8042 = ~n8040 & ~n8041;
  assign n8043 = ~po29  & n8036;
  assign n8044 = ~n8042 & ~n8043;
  assign n8045 = ~n8037 & ~n8044;
  assign n8046 = po30  & ~n8045;
  assign n8047 = ~po30  & ~n8037;
  assign n8048 = ~n8044 & n8047;
  assign n8049 = ~n7653 & ~n7654;
  assign n8050 = po23  & n8049;
  assign n8051 = n7659 & n8050;
  assign n8052 = ~n7659 & ~n8050;
  assign n8053 = ~n8051 & ~n8052;
  assign n8054 = ~n8048 & n8053;
  assign n8055 = ~n8046 & ~n8054;
  assign n8056 = po31  & ~n8055;
  assign n8057 = ~n7662 & ~n7664;
  assign n8058 = po23  & n8057;
  assign n8059 = n7669 & ~n8058;
  assign n8060 = ~n7669 & n8058;
  assign n8061 = ~n8059 & ~n8060;
  assign n8062 = ~po31  & n8055;
  assign n8063 = ~n8061 & ~n8062;
  assign n8064 = ~n8056 & ~n8063;
  assign n8065 = po32  & ~n8064;
  assign n8066 = ~po32  & ~n8056;
  assign n8067 = ~n8063 & n8066;
  assign n8068 = ~n7672 & ~n7673;
  assign n8069 = po23  & n8068;
  assign n8070 = ~n7678 & ~n8069;
  assign n8071 = n7678 & n8069;
  assign n8072 = ~n8070 & ~n8071;
  assign n8073 = ~n8067 & n8072;
  assign n8074 = ~n8065 & ~n8073;
  assign n8075 = po33  & ~n8074;
  assign n8076 = ~n7681 & ~n7683;
  assign n8077 = po23  & n8076;
  assign n8078 = n7688 & ~n8077;
  assign n8079 = ~n7688 & n8077;
  assign n8080 = ~n8078 & ~n8079;
  assign n8081 = ~po33  & n8074;
  assign n8082 = ~n8080 & ~n8081;
  assign n8083 = ~n8075 & ~n8082;
  assign n8084 = po34  & ~n8083;
  assign n8085 = ~n7691 & ~n7692;
  assign n8086 = po23  & n8085;
  assign n8087 = n7697 & ~n8086;
  assign n8088 = ~n7697 & n8086;
  assign n8089 = ~n8087 & ~n8088;
  assign n8090 = ~po34  & ~n8075;
  assign n8091 = ~n8082 & n8090;
  assign n8092 = ~n8089 & ~n8091;
  assign n8093 = ~n8084 & ~n8092;
  assign n8094 = po35  & ~n8093;
  assign n8095 = ~n7700 & ~n7702;
  assign n8096 = po23  & n8095;
  assign n8097 = n7707 & ~n8096;
  assign n8098 = ~n7707 & n8096;
  assign n8099 = ~n8097 & ~n8098;
  assign n8100 = ~po35  & n8093;
  assign n8101 = ~n8099 & ~n8100;
  assign n8102 = ~n8094 & ~n8101;
  assign n8103 = po36  & ~n8102;
  assign n8104 = ~po36  & ~n8094;
  assign n8105 = ~n8101 & n8104;
  assign n8106 = ~n7710 & po23 ;
  assign n8107 = ~n7716 & n8106;
  assign n8108 = n7715 & ~n8107;
  assign n8109 = n7717 & n8106;
  assign n8110 = ~n8108 & ~n8109;
  assign n8111 = ~n8105 & n8110;
  assign n8112 = ~n8103 & ~n8111;
  assign n8113 = po37  & ~n8112;
  assign n8114 = ~n7719 & ~n7721;
  assign n8115 = po23  & n8114;
  assign n8116 = n7726 & ~n8115;
  assign n8117 = ~n7726 & n8115;
  assign n8118 = ~n8116 & ~n8117;
  assign n8119 = ~po37  & n8112;
  assign n8120 = ~n8118 & ~n8119;
  assign n8121 = ~n8113 & ~n8120;
  assign n8122 = po38  & ~n8121;
  assign n8123 = ~n7729 & ~n7730;
  assign n8124 = po23  & n8123;
  assign n8125 = n7735 & ~n8124;
  assign n8126 = ~n7735 & n8124;
  assign n8127 = ~n8125 & ~n8126;
  assign n8128 = ~po38  & ~n8113;
  assign n8129 = ~n8120 & n8128;
  assign n8130 = ~n8127 & ~n8129;
  assign n8131 = ~n8122 & ~n8130;
  assign n8132 = ~po39  & n8131;
  assign n8133 = ~n7738 & po23 ;
  assign n8134 = ~n7745 & n8133;
  assign n8135 = n7743 & ~n8134;
  assign n8136 = n7746 & n8133;
  assign n8137 = ~n8135 & ~n8136;
  assign n8138 = ~n8132 & n8137;
  assign n8139 = po39  & ~n8131;
  assign n8140 = ~n8138 & ~n8139;
  assign n8141 = po40  & ~n8140;
  assign n8142 = ~n7748 & ~n7750;
  assign n8143 = po23  & n8142;
  assign n8144 = n7611 & ~n8143;
  assign n8145 = ~n7611 & n8143;
  assign n8146 = ~n8144 & ~n8145;
  assign n8147 = ~po40  & ~n8139;
  assign n8148 = ~n8138 & n8147;
  assign n8149 = n8146 & ~n8148;
  assign n8150 = ~n8141 & ~n8149;
  assign n8151 = ~po41  & n8150;
  assign n8152 = po41  & ~n8150;
  assign n8153 = ~n7986 & ~n8151;
  assign n8154 = ~n8152 & ~n8153;
  assign n8155 = po42  & ~n8154;
  assign n8156 = ~po42  & ~n8152;
  assign n8157 = ~n8153 & n8156;
  assign n8158 = ~n7757 & po23 ;
  assign n8159 = ~n7763 & n8158;
  assign n8160 = n7762 & ~n8159;
  assign n8161 = n7764 & n8158;
  assign n8162 = ~n8160 & ~n8161;
  assign n8163 = ~n8157 & n8162;
  assign n8164 = ~n8155 & ~n8163;
  assign n8165 = po43  & ~n8164;
  assign n8166 = ~n7766 & ~n7768;
  assign n8167 = po23  & n8166;
  assign n8168 = n7773 & ~n8167;
  assign n8169 = ~n7773 & n8167;
  assign n8170 = ~n8168 & ~n8169;
  assign n8171 = ~po43  & n8164;
  assign n8172 = ~n8170 & ~n8171;
  assign n8173 = ~n8165 & ~n8172;
  assign n8174 = po44  & ~n8173;
  assign n8175 = ~po44  & ~n8165;
  assign n8176 = ~n8172 & n8175;
  assign n8177 = ~n7776 & po23 ;
  assign n8178 = ~n7782 & n8177;
  assign n8179 = n7781 & ~n8178;
  assign n8180 = n7783 & n8177;
  assign n8181 = ~n8179 & ~n8180;
  assign n8182 = ~n8176 & n8181;
  assign n8183 = ~n8174 & ~n8182;
  assign n8184 = po45  & ~n8183;
  assign n8185 = ~n7785 & ~n7787;
  assign n8186 = po23  & n8185;
  assign n8187 = n7792 & ~n8186;
  assign n8188 = ~n7792 & n8186;
  assign n8189 = ~n8187 & ~n8188;
  assign n8190 = ~po45  & n8183;
  assign n8191 = ~n8189 & ~n8190;
  assign n8192 = ~n8184 & ~n8191;
  assign n8193 = po46  & ~n8192;
  assign n8194 = ~n7795 & ~n7796;
  assign n8195 = po23  & n8194;
  assign n8196 = n7801 & ~n8195;
  assign n8197 = ~n7801 & n8195;
  assign n8198 = ~n8196 & ~n8197;
  assign n8199 = ~po46  & ~n8184;
  assign n8200 = ~n8191 & n8199;
  assign n8201 = ~n8198 & ~n8200;
  assign n8202 = ~n8193 & ~n8201;
  assign n8203 = po47  & ~n8202;
  assign n8204 = ~n7804 & ~n7806;
  assign n8205 = po23  & n8204;
  assign n8206 = n7811 & ~n8205;
  assign n8207 = ~n7811 & n8205;
  assign n8208 = ~n8206 & ~n8207;
  assign n8209 = ~po47  & n8202;
  assign n8210 = ~n8208 & ~n8209;
  assign n8211 = ~n8203 & ~n8210;
  assign n8212 = po48  & ~n8211;
  assign n8213 = ~po48  & ~n8203;
  assign n8214 = ~n8210 & n8213;
  assign n8215 = ~n7814 & po23 ;
  assign n8216 = ~n7820 & n8215;
  assign n8217 = n7819 & ~n8216;
  assign n8218 = n7821 & n8215;
  assign n8219 = ~n8217 & ~n8218;
  assign n8220 = ~n8214 & n8219;
  assign n8221 = ~n8212 & ~n8220;
  assign n8222 = po49  & ~n8221;
  assign n8223 = ~n7823 & ~n7825;
  assign n8224 = po23  & n8223;
  assign n8225 = n7830 & ~n8224;
  assign n8226 = ~n7830 & n8224;
  assign n8227 = ~n8225 & ~n8226;
  assign n8228 = ~po49  & n8221;
  assign n8229 = ~n8227 & ~n8228;
  assign n8230 = ~n8222 & ~n8229;
  assign n8231 = po50  & ~n8230;
  assign n8232 = ~n7833 & ~n7834;
  assign n8233 = po23  & n8232;
  assign n8234 = n7839 & ~n8233;
  assign n8235 = ~n7839 & n8233;
  assign n8236 = ~n8234 & ~n8235;
  assign n8237 = ~po50  & ~n8222;
  assign n8238 = ~n8229 & n8237;
  assign n8239 = ~n8236 & ~n8238;
  assign n8240 = ~n8231 & ~n8239;
  assign n8241 = po51  & ~n8240;
  assign n8242 = ~n7842 & ~n7844;
  assign n8243 = po23  & n8242;
  assign n8244 = n7849 & ~n8243;
  assign n8245 = ~n7849 & n8243;
  assign n8246 = ~n8244 & ~n8245;
  assign n8247 = ~po51  & n8240;
  assign n8248 = ~n8246 & ~n8247;
  assign n8249 = ~n8241 & ~n8248;
  assign n8250 = po52  & ~n8249;
  assign n8251 = ~po52  & ~n8241;
  assign n8252 = ~n8248 & n8251;
  assign n8253 = ~n7852 & po23 ;
  assign n8254 = ~n7858 & n8253;
  assign n8255 = n7857 & ~n8254;
  assign n8256 = n7859 & n8253;
  assign n8257 = ~n8255 & ~n8256;
  assign n8258 = ~n8252 & n8257;
  assign n8259 = ~n8250 & ~n8258;
  assign n8260 = po53  & ~n8259;
  assign n8261 = ~n7861 & ~n7863;
  assign n8262 = po23  & n8261;
  assign n8263 = n7868 & ~n8262;
  assign n8264 = ~n7868 & n8262;
  assign n8265 = ~n8263 & ~n8264;
  assign n8266 = ~po53  & n8259;
  assign n8267 = ~n8265 & ~n8266;
  assign n8268 = ~n8260 & ~n8267;
  assign n8269 = po54  & ~n8268;
  assign n8270 = ~n7871 & ~n7872;
  assign n8271 = po23  & n8270;
  assign n8272 = n7877 & ~n8271;
  assign n8273 = ~n7877 & n8271;
  assign n8274 = ~n8272 & ~n8273;
  assign n8275 = ~po54  & ~n8260;
  assign n8276 = ~n8267 & n8275;
  assign n8277 = ~n8274 & ~n8276;
  assign n8278 = ~n8269 & ~n8277;
  assign n8279 = po55  & ~n8278;
  assign n8280 = ~n7880 & ~n7882;
  assign n8281 = po23  & n8280;
  assign n8282 = n7887 & ~n8281;
  assign n8283 = ~n7887 & n8281;
  assign n8284 = ~n8282 & ~n8283;
  assign n8285 = ~po55  & n8278;
  assign n8286 = ~n8284 & ~n8285;
  assign n8287 = ~n8279 & ~n8286;
  assign n8288 = po56  & ~n8287;
  assign n8289 = ~po56  & ~n8279;
  assign n8290 = ~n8286 & n8289;
  assign n8291 = ~n7890 & po23 ;
  assign n8292 = ~n7896 & n8291;
  assign n8293 = n7895 & ~n8292;
  assign n8294 = n7897 & n8291;
  assign n8295 = ~n8293 & ~n8294;
  assign n8296 = ~n8290 & n8295;
  assign n8297 = ~n8288 & ~n8296;
  assign n8298 = po57  & ~n8297;
  assign n8299 = ~n7899 & ~n7901;
  assign n8300 = po23  & n8299;
  assign n8301 = n7906 & ~n8300;
  assign n8302 = ~n7906 & n8300;
  assign n8303 = ~n8301 & ~n8302;
  assign n8304 = ~po57  & n8297;
  assign n8305 = ~n8303 & ~n8304;
  assign n8306 = ~n8298 & ~n8305;
  assign n8307 = po58  & ~n8306;
  assign n8308 = ~n7909 & ~n7910;
  assign n8309 = po23  & n8308;
  assign n8310 = n7915 & ~n8309;
  assign n8311 = ~n7915 & n8309;
  assign n8312 = ~n8310 & ~n8311;
  assign n8313 = ~po58  & ~n8298;
  assign n8314 = ~n8305 & n8313;
  assign n8315 = ~n8312 & ~n8314;
  assign n8316 = ~n8307 & ~n8315;
  assign n8317 = po59  & ~n8316;
  assign n8318 = ~n7918 & ~n7920;
  assign n8319 = po23  & n8318;
  assign n8320 = n7925 & ~n8319;
  assign n8321 = ~n7925 & n8319;
  assign n8322 = ~n8320 & ~n8321;
  assign n8323 = ~po59  & n8316;
  assign n8324 = ~n8322 & ~n8323;
  assign n8325 = ~n8317 & ~n8324;
  assign n8326 = po60  & ~n8325;
  assign n8327 = ~po60  & ~n8317;
  assign n8328 = ~n8324 & n8327;
  assign n8329 = ~n7928 & po23 ;
  assign n8330 = ~n7934 & n8329;
  assign n8331 = n7933 & ~n8330;
  assign n8332 = n7935 & n8329;
  assign n8333 = ~n8331 & ~n8332;
  assign n8334 = ~n8328 & n8333;
  assign n8335 = ~n8326 & ~n8334;
  assign n8336 = po61  & ~n8335;
  assign n8337 = ~n7937 & ~n7939;
  assign n8338 = po23  & n8337;
  assign n8339 = n7944 & ~n8338;
  assign n8340 = ~n7944 & n8338;
  assign n8341 = ~n8339 & ~n8340;
  assign n8342 = ~po61  & n8335;
  assign n8343 = ~n8341 & ~n8342;
  assign n8344 = ~n8336 & ~n8343;
  assign n8345 = po62  & ~n8344;
  assign n8346 = ~n7947 & ~n7948;
  assign n8347 = po23  & n8346;
  assign n8348 = n7953 & ~n8347;
  assign n8349 = ~n7953 & n8347;
  assign n8350 = ~n8348 & ~n8349;
  assign n8351 = ~po62  & ~n8336;
  assign n8352 = ~n8343 & n8351;
  assign n8353 = ~n8350 & ~n8352;
  assign n8354 = ~n8345 & ~n8353;
  assign n8355 = ~n7956 & ~n7958;
  assign n8356 = po23  & n8355;
  assign n8357 = n7963 & ~n8356;
  assign n8358 = ~n7963 & n8356;
  assign n8359 = ~n8357 & ~n8358;
  assign n8360 = n7965 & po23 ;
  assign n8361 = ~n7970 & ~n8360;
  assign n8362 = ~n7978 & ~n8361;
  assign n8363 = po23  & ~n8362;
  assign n8364 = ~n8359 & ~n8363;
  assign n8365 = ~n8354 & n8364;
  assign n8366 = ~po63  & ~n8365;
  assign n8367 = n8354 & n8359;
  assign n8368 = po63  & n8362;
  assign n8369 = ~n8367 & ~n8368;
  assign po22  = n8366 | ~n8369;
  assign n8371 = ~n8152 & po22 ;
  assign n8372 = ~n8151 & n8371;
  assign n8373 = n7986 & ~n8372;
  assign n8374 = n8153 & n8371;
  assign n8375 = ~n8373 & ~n8374;
  assign n8376 = pi44  & po22 ;
  assign n8377 = ~pi42  & ~pi43 ;
  assign n8378 = ~pi44  & n8377;
  assign n8379 = ~n8376 & ~n8378;
  assign n8380 = po23  & ~n8379;
  assign n8381 = ~pi44  & po22 ;
  assign n8382 = pi45  & ~n8381;
  assign n8383 = ~pi45  & n8381;
  assign n8384 = ~n8382 & ~n8383;
  assign n8385 = ~po23  & n8379;
  assign n8386 = n8384 & ~n8385;
  assign n8387 = ~n8380 & ~n8386;
  assign n8388 = po24  & ~n8387;
  assign n8389 = ~po24  & ~n8380;
  assign n8390 = ~n8386 & n8389;
  assign n8391 = po23  & ~po22 ;
  assign n8392 = ~n8383 & ~n8391;
  assign n8393 = pi46  & ~n8392;
  assign n8394 = ~pi46  & n8392;
  assign n8395 = ~n8393 & ~n8394;
  assign n8396 = ~n8390 & ~n8395;
  assign n8397 = ~n8388 & ~n8396;
  assign n8398 = po25  & ~n8397;
  assign n8399 = ~po25  & n8397;
  assign n8400 = ~n7991 & ~n7992;
  assign n8401 = po22  & n8400;
  assign n8402 = n7996 & ~n8401;
  assign n8403 = ~n7996 & n8401;
  assign n8404 = ~n8402 & ~n8403;
  assign n8405 = ~n8399 & ~n8404;
  assign n8406 = ~n8398 & ~n8405;
  assign n8407 = po26  & ~n8406;
  assign n8408 = ~po26  & ~n8398;
  assign n8409 = ~n8405 & n8408;
  assign n8410 = ~n7999 & po22 ;
  assign n8411 = ~n8005 & n8410;
  assign n8412 = n8004 & ~n8411;
  assign n8413 = n8006 & n8410;
  assign n8414 = ~n8412 & ~n8413;
  assign n8415 = ~n8409 & n8414;
  assign n8416 = ~n8407 & ~n8415;
  assign n8417 = po27  & ~n8416;
  assign n8418 = ~po27  & n8416;
  assign n8419 = ~n8008 & ~n8010;
  assign n8420 = po22  & n8419;
  assign n8421 = n8015 & ~n8420;
  assign n8422 = ~n8015 & n8420;
  assign n8423 = ~n8421 & ~n8422;
  assign n8424 = ~n8418 & n8423;
  assign n8425 = ~n8417 & ~n8424;
  assign n8426 = po28  & ~n8425;
  assign n8427 = ~po28  & ~n8417;
  assign n8428 = ~n8424 & n8427;
  assign n8429 = ~n8018 & po22 ;
  assign n8430 = ~n8024 & n8429;
  assign n8431 = n8023 & ~n8430;
  assign n8432 = n8025 & n8429;
  assign n8433 = ~n8431 & ~n8432;
  assign n8434 = ~n8428 & n8433;
  assign n8435 = ~n8426 & ~n8434;
  assign n8436 = po29  & ~n8435;
  assign n8437 = ~po29  & n8435;
  assign n8438 = ~n8027 & ~n8029;
  assign n8439 = po22  & n8438;
  assign n8440 = n8034 & n8439;
  assign n8441 = ~n8034 & ~n8439;
  assign n8442 = ~n8440 & ~n8441;
  assign n8443 = ~n8437 & n8442;
  assign n8444 = ~n8436 & ~n8443;
  assign n8445 = po30  & ~n8444;
  assign n8446 = ~po30  & ~n8436;
  assign n8447 = ~n8443 & n8446;
  assign n8448 = ~n8037 & po22 ;
  assign n8449 = ~n8043 & n8448;
  assign n8450 = n8042 & ~n8449;
  assign n8451 = n8044 & n8448;
  assign n8452 = ~n8450 & ~n8451;
  assign n8453 = ~n8447 & n8452;
  assign n8454 = ~n8445 & ~n8453;
  assign n8455 = po31  & ~n8454;
  assign n8456 = ~po31  & n8454;
  assign n8457 = ~n8046 & ~n8048;
  assign n8458 = po22  & n8457;
  assign n8459 = ~n8053 & ~n8458;
  assign n8460 = n8053 & n8458;
  assign n8461 = ~n8459 & ~n8460;
  assign n8462 = ~n8456 & n8461;
  assign n8463 = ~n8455 & ~n8462;
  assign n8464 = po32  & ~n8463;
  assign n8465 = ~po32  & ~n8455;
  assign n8466 = ~n8462 & n8465;
  assign n8467 = ~n8056 & po22 ;
  assign n8468 = ~n8062 & n8467;
  assign n8469 = n8061 & ~n8468;
  assign n8470 = n8063 & n8467;
  assign n8471 = ~n8469 & ~n8470;
  assign n8472 = ~n8466 & n8471;
  assign n8473 = ~n8464 & ~n8472;
  assign n8474 = po33  & ~n8473;
  assign n8475 = ~n8065 & ~n8067;
  assign n8476 = po22  & n8475;
  assign n8477 = n8072 & ~n8476;
  assign n8478 = ~n8072 & n8476;
  assign n8479 = ~n8477 & ~n8478;
  assign n8480 = ~po33  & n8473;
  assign n8481 = ~n8479 & ~n8480;
  assign n8482 = ~n8474 & ~n8481;
  assign n8483 = po34  & ~n8482;
  assign n8484 = ~po34  & ~n8474;
  assign n8485 = ~n8481 & n8484;
  assign n8486 = ~n8075 & po22 ;
  assign n8487 = ~n8081 & n8486;
  assign n8488 = n8080 & ~n8487;
  assign n8489 = n8082 & n8486;
  assign n8490 = ~n8488 & ~n8489;
  assign n8491 = ~n8485 & n8490;
  assign n8492 = ~n8483 & ~n8491;
  assign n8493 = po35  & ~n8492;
  assign n8494 = ~po35  & n8492;
  assign n8495 = ~n8084 & po22 ;
  assign n8496 = ~n8091 & n8495;
  assign n8497 = n8089 & ~n8496;
  assign n8498 = n8092 & n8495;
  assign n8499 = ~n8497 & ~n8498;
  assign n8500 = ~n8494 & n8499;
  assign n8501 = ~n8493 & ~n8500;
  assign n8502 = po36  & ~n8501;
  assign n8503 = ~po36  & ~n8493;
  assign n8504 = ~n8500 & n8503;
  assign n8505 = ~n8094 & po22 ;
  assign n8506 = ~n8100 & n8505;
  assign n8507 = n8099 & ~n8506;
  assign n8508 = n8101 & n8505;
  assign n8509 = ~n8507 & ~n8508;
  assign n8510 = ~n8504 & n8509;
  assign n8511 = ~n8502 & ~n8510;
  assign n8512 = po37  & ~n8511;
  assign n8513 = ~n8103 & ~n8105;
  assign n8514 = po22  & n8513;
  assign n8515 = n8110 & ~n8514;
  assign n8516 = ~n8110 & n8514;
  assign n8517 = ~n8515 & ~n8516;
  assign n8518 = ~po37  & n8511;
  assign n8519 = ~n8517 & ~n8518;
  assign n8520 = ~n8512 & ~n8519;
  assign n8521 = po38  & ~n8520;
  assign n8522 = ~po38  & ~n8512;
  assign n8523 = ~n8519 & n8522;
  assign n8524 = ~n8113 & po22 ;
  assign n8525 = ~n8119 & n8524;
  assign n8526 = n8118 & ~n8525;
  assign n8527 = n8120 & n8524;
  assign n8528 = ~n8526 & ~n8527;
  assign n8529 = ~n8523 & n8528;
  assign n8530 = ~n8521 & ~n8529;
  assign n8531 = po39  & ~n8530;
  assign n8532 = ~po39  & n8530;
  assign n8533 = ~n8122 & po22 ;
  assign n8534 = ~n8129 & n8533;
  assign n8535 = n8127 & ~n8534;
  assign n8536 = n8130 & n8533;
  assign n8537 = ~n8535 & ~n8536;
  assign n8538 = ~n8532 & n8537;
  assign n8539 = ~n8531 & ~n8538;
  assign n8540 = po40  & ~n8539;
  assign n8541 = ~n8132 & ~n8139;
  assign n8542 = po22  & n8541;
  assign n8543 = n8137 & ~n8542;
  assign n8544 = ~n8137 & n8542;
  assign n8545 = ~n8543 & ~n8544;
  assign n8546 = ~po40  & ~n8531;
  assign n8547 = ~n8538 & n8546;
  assign n8548 = ~n8545 & ~n8547;
  assign n8549 = ~n8540 & ~n8548;
  assign n8550 = ~po41  & n8549;
  assign n8551 = ~n8141 & ~n8148;
  assign n8552 = po22  & n8551;
  assign n8553 = n8146 & n8552;
  assign n8554 = ~n8146 & ~n8552;
  assign n8555 = ~n8553 & ~n8554;
  assign n8556 = ~n8550 & n8555;
  assign n8557 = po41  & ~n8549;
  assign n8558 = ~po42  & ~n8557;
  assign n8559 = ~n8556 & n8558;
  assign n8560 = ~n8556 & ~n8557;
  assign n8561 = po42  & ~n8560;
  assign n8562 = n8375 & ~n8559;
  assign n8563 = ~n8561 & ~n8562;
  assign n8564 = po43  & ~n8563;
  assign n8565 = ~n8155 & ~n8157;
  assign n8566 = po22  & n8565;
  assign n8567 = n8162 & ~n8566;
  assign n8568 = ~n8162 & n8566;
  assign n8569 = ~n8567 & ~n8568;
  assign n8570 = ~po43  & n8563;
  assign n8571 = ~n8569 & ~n8570;
  assign n8572 = ~n8564 & ~n8571;
  assign n8573 = po44  & ~n8572;
  assign n8574 = ~po44  & ~n8564;
  assign n8575 = ~n8571 & n8574;
  assign n8576 = ~n8165 & po22 ;
  assign n8577 = ~n8171 & n8576;
  assign n8578 = n8170 & ~n8577;
  assign n8579 = n8172 & n8576;
  assign n8580 = ~n8578 & ~n8579;
  assign n8581 = ~n8575 & n8580;
  assign n8582 = ~n8573 & ~n8581;
  assign n8583 = po45  & ~n8582;
  assign n8584 = ~n8174 & ~n8176;
  assign n8585 = po22  & n8584;
  assign n8586 = n8181 & ~n8585;
  assign n8587 = ~n8181 & n8585;
  assign n8588 = ~n8586 & ~n8587;
  assign n8589 = ~po45  & n8582;
  assign n8590 = ~n8588 & ~n8589;
  assign n8591 = ~n8583 & ~n8590;
  assign n8592 = po46  & ~n8591;
  assign n8593 = ~po46  & ~n8583;
  assign n8594 = ~n8590 & n8593;
  assign n8595 = ~n8184 & po22 ;
  assign n8596 = ~n8190 & n8595;
  assign n8597 = n8189 & ~n8596;
  assign n8598 = n8191 & n8595;
  assign n8599 = ~n8597 & ~n8598;
  assign n8600 = ~n8594 & n8599;
  assign n8601 = ~n8592 & ~n8600;
  assign n8602 = po47  & ~n8601;
  assign n8603 = ~po47  & n8601;
  assign n8604 = ~n8193 & po22 ;
  assign n8605 = ~n8200 & n8604;
  assign n8606 = n8198 & ~n8605;
  assign n8607 = n8201 & n8604;
  assign n8608 = ~n8606 & ~n8607;
  assign n8609 = ~n8603 & n8608;
  assign n8610 = ~n8602 & ~n8609;
  assign n8611 = po48  & ~n8610;
  assign n8612 = ~po48  & ~n8602;
  assign n8613 = ~n8609 & n8612;
  assign n8614 = ~n8203 & po22 ;
  assign n8615 = ~n8209 & n8614;
  assign n8616 = n8208 & ~n8615;
  assign n8617 = n8210 & n8614;
  assign n8618 = ~n8616 & ~n8617;
  assign n8619 = ~n8613 & n8618;
  assign n8620 = ~n8611 & ~n8619;
  assign n8621 = po49  & ~n8620;
  assign n8622 = ~n8212 & ~n8214;
  assign n8623 = po22  & n8622;
  assign n8624 = n8219 & ~n8623;
  assign n8625 = ~n8219 & n8623;
  assign n8626 = ~n8624 & ~n8625;
  assign n8627 = ~po49  & n8620;
  assign n8628 = ~n8626 & ~n8627;
  assign n8629 = ~n8621 & ~n8628;
  assign n8630 = po50  & ~n8629;
  assign n8631 = ~po50  & ~n8621;
  assign n8632 = ~n8628 & n8631;
  assign n8633 = ~n8222 & po22 ;
  assign n8634 = ~n8228 & n8633;
  assign n8635 = n8227 & ~n8634;
  assign n8636 = n8229 & n8633;
  assign n8637 = ~n8635 & ~n8636;
  assign n8638 = ~n8632 & n8637;
  assign n8639 = ~n8630 & ~n8638;
  assign n8640 = po51  & ~n8639;
  assign n8641 = ~po51  & n8639;
  assign n8642 = ~n8231 & po22 ;
  assign n8643 = ~n8238 & n8642;
  assign n8644 = n8236 & ~n8643;
  assign n8645 = n8239 & n8642;
  assign n8646 = ~n8644 & ~n8645;
  assign n8647 = ~n8641 & n8646;
  assign n8648 = ~n8640 & ~n8647;
  assign n8649 = po52  & ~n8648;
  assign n8650 = ~po52  & ~n8640;
  assign n8651 = ~n8647 & n8650;
  assign n8652 = ~n8241 & po22 ;
  assign n8653 = ~n8247 & n8652;
  assign n8654 = n8246 & ~n8653;
  assign n8655 = n8248 & n8652;
  assign n8656 = ~n8654 & ~n8655;
  assign n8657 = ~n8651 & n8656;
  assign n8658 = ~n8649 & ~n8657;
  assign n8659 = po53  & ~n8658;
  assign n8660 = ~n8250 & ~n8252;
  assign n8661 = po22  & n8660;
  assign n8662 = n8257 & ~n8661;
  assign n8663 = ~n8257 & n8661;
  assign n8664 = ~n8662 & ~n8663;
  assign n8665 = ~po53  & n8658;
  assign n8666 = ~n8664 & ~n8665;
  assign n8667 = ~n8659 & ~n8666;
  assign n8668 = po54  & ~n8667;
  assign n8669 = ~po54  & ~n8659;
  assign n8670 = ~n8666 & n8669;
  assign n8671 = ~n8260 & po22 ;
  assign n8672 = ~n8266 & n8671;
  assign n8673 = n8265 & ~n8672;
  assign n8674 = n8267 & n8671;
  assign n8675 = ~n8673 & ~n8674;
  assign n8676 = ~n8670 & n8675;
  assign n8677 = ~n8668 & ~n8676;
  assign n8678 = po55  & ~n8677;
  assign n8679 = ~po55  & n8677;
  assign n8680 = ~n8269 & po22 ;
  assign n8681 = ~n8276 & n8680;
  assign n8682 = n8274 & ~n8681;
  assign n8683 = n8277 & n8680;
  assign n8684 = ~n8682 & ~n8683;
  assign n8685 = ~n8679 & n8684;
  assign n8686 = ~n8678 & ~n8685;
  assign n8687 = po56  & ~n8686;
  assign n8688 = ~po56  & ~n8678;
  assign n8689 = ~n8685 & n8688;
  assign n8690 = ~n8279 & po22 ;
  assign n8691 = ~n8285 & n8690;
  assign n8692 = n8284 & ~n8691;
  assign n8693 = n8286 & n8690;
  assign n8694 = ~n8692 & ~n8693;
  assign n8695 = ~n8689 & n8694;
  assign n8696 = ~n8687 & ~n8695;
  assign n8697 = po57  & ~n8696;
  assign n8698 = ~n8288 & ~n8290;
  assign n8699 = po22  & n8698;
  assign n8700 = n8295 & ~n8699;
  assign n8701 = ~n8295 & n8699;
  assign n8702 = ~n8700 & ~n8701;
  assign n8703 = ~po57  & n8696;
  assign n8704 = ~n8702 & ~n8703;
  assign n8705 = ~n8697 & ~n8704;
  assign n8706 = po58  & ~n8705;
  assign n8707 = ~po58  & ~n8697;
  assign n8708 = ~n8704 & n8707;
  assign n8709 = ~n8298 & po22 ;
  assign n8710 = ~n8304 & n8709;
  assign n8711 = n8303 & ~n8710;
  assign n8712 = n8305 & n8709;
  assign n8713 = ~n8711 & ~n8712;
  assign n8714 = ~n8708 & n8713;
  assign n8715 = ~n8706 & ~n8714;
  assign n8716 = po59  & ~n8715;
  assign n8717 = ~po59  & n8715;
  assign n8718 = ~n8307 & po22 ;
  assign n8719 = ~n8314 & n8718;
  assign n8720 = n8312 & ~n8719;
  assign n8721 = n8315 & n8718;
  assign n8722 = ~n8720 & ~n8721;
  assign n8723 = ~n8717 & n8722;
  assign n8724 = ~n8716 & ~n8723;
  assign n8725 = po60  & ~n8724;
  assign n8726 = ~po60  & ~n8716;
  assign n8727 = ~n8723 & n8726;
  assign n8728 = ~n8317 & po22 ;
  assign n8729 = ~n8323 & n8728;
  assign n8730 = n8322 & ~n8729;
  assign n8731 = n8324 & n8728;
  assign n8732 = ~n8730 & ~n8731;
  assign n8733 = ~n8727 & n8732;
  assign n8734 = ~n8725 & ~n8733;
  assign n8735 = po61  & ~n8734;
  assign n8736 = ~n8326 & ~n8328;
  assign n8737 = po22  & n8736;
  assign n8738 = n8333 & ~n8737;
  assign n8739 = ~n8333 & n8737;
  assign n8740 = ~n8738 & ~n8739;
  assign n8741 = ~po61  & n8734;
  assign n8742 = ~n8740 & ~n8741;
  assign n8743 = ~n8735 & ~n8742;
  assign n8744 = po62  & ~n8743;
  assign n8745 = ~po62  & ~n8735;
  assign n8746 = ~n8742 & n8745;
  assign n8747 = ~n8336 & po22 ;
  assign n8748 = ~n8342 & n8747;
  assign n8749 = n8341 & ~n8748;
  assign n8750 = n8343 & n8747;
  assign n8751 = ~n8749 & ~n8750;
  assign n8752 = ~n8746 & n8751;
  assign n8753 = ~n8744 & ~n8752;
  assign n8754 = n8354 & po22 ;
  assign n8755 = ~n8359 & ~n8754;
  assign n8756 = ~n8367 & ~n8755;
  assign n8757 = po22  & ~n8756;
  assign n8758 = ~n8345 & po22 ;
  assign n8759 = ~n8352 & n8758;
  assign n8760 = n8350 & ~n8759;
  assign n8761 = n8353 & n8758;
  assign n8762 = ~n8760 & ~n8761;
  assign n8763 = ~n8757 & n8762;
  assign n8764 = ~n8753 & n8763;
  assign n8765 = ~po63  & ~n8764;
  assign n8766 = n8753 & ~n8762;
  assign n8767 = po63  & n8756;
  assign n8768 = ~n8766 & ~n8767;
  assign po21  = n8765 | ~n8768;
  assign n8770 = ~n8559 & ~n8561;
  assign n8771 = po21  & n8770;
  assign n8772 = n8375 & ~n8771;
  assign n8773 = ~n8375 & n8771;
  assign n8774 = ~n8772 & ~n8773;
  assign n8775 = pi42  & po21 ;
  assign n8776 = ~pi40  & ~pi41 ;
  assign n8777 = ~pi42  & n8776;
  assign n8778 = ~n8775 & ~n8777;
  assign n8779 = po22  & ~n8778;
  assign n8780 = ~po22  & n8778;
  assign n8781 = ~pi42  & po21 ;
  assign n8782 = pi43  & ~n8781;
  assign n8783 = ~pi43  & n8781;
  assign n8784 = ~n8782 & ~n8783;
  assign n8785 = ~n8780 & n8784;
  assign n8786 = ~n8779 & ~n8785;
  assign n8787 = po23  & ~n8786;
  assign n8788 = po22  & ~po21 ;
  assign n8789 = ~n8783 & ~n8788;
  assign n8790 = pi44  & ~n8789;
  assign n8791 = ~pi44  & n8789;
  assign n8792 = ~n8790 & ~n8791;
  assign n8793 = ~po23  & n8786;
  assign n8794 = ~n8792 & ~n8793;
  assign n8795 = ~n8787 & ~n8794;
  assign n8796 = po24  & ~n8795;
  assign n8797 = ~po24  & ~n8787;
  assign n8798 = ~n8794 & n8797;
  assign n8799 = ~n8380 & ~n8385;
  assign n8800 = po21  & n8799;
  assign n8801 = n8384 & ~n8800;
  assign n8802 = ~n8384 & n8800;
  assign n8803 = ~n8801 & ~n8802;
  assign n8804 = ~n8798 & ~n8803;
  assign n8805 = ~n8796 & ~n8804;
  assign n8806 = po25  & ~n8805;
  assign n8807 = ~n8388 & ~n8390;
  assign n8808 = po21  & n8807;
  assign n8809 = ~n8395 & ~n8808;
  assign n8810 = n8395 & n8808;
  assign n8811 = ~n8809 & ~n8810;
  assign n8812 = ~po25  & n8805;
  assign n8813 = ~n8811 & ~n8812;
  assign n8814 = ~n8806 & ~n8813;
  assign n8815 = po26  & ~n8814;
  assign n8816 = ~po26  & ~n8806;
  assign n8817 = ~n8813 & n8816;
  assign n8818 = ~n8398 & ~n8399;
  assign n8819 = po21  & n8818;
  assign n8820 = n8404 & ~n8819;
  assign n8821 = ~n8404 & n8819;
  assign n8822 = ~n8820 & ~n8821;
  assign n8823 = ~n8817 & n8822;
  assign n8824 = ~n8815 & ~n8823;
  assign n8825 = po27  & ~n8824;
  assign n8826 = ~n8407 & ~n8409;
  assign n8827 = po21  & n8826;
  assign n8828 = n8414 & ~n8827;
  assign n8829 = ~n8414 & n8827;
  assign n8830 = ~n8828 & ~n8829;
  assign n8831 = ~po27  & n8824;
  assign n8832 = ~n8830 & ~n8831;
  assign n8833 = ~n8825 & ~n8832;
  assign n8834 = po28  & ~n8833;
  assign n8835 = ~po28  & ~n8825;
  assign n8836 = ~n8832 & n8835;
  assign n8837 = ~n8417 & ~n8418;
  assign n8838 = po21  & n8837;
  assign n8839 = n8423 & n8838;
  assign n8840 = ~n8423 & ~n8838;
  assign n8841 = ~n8839 & ~n8840;
  assign n8842 = ~n8836 & n8841;
  assign n8843 = ~n8834 & ~n8842;
  assign n8844 = po29  & ~n8843;
  assign n8845 = ~n8426 & ~n8428;
  assign n8846 = po21  & n8845;
  assign n8847 = n8433 & ~n8846;
  assign n8848 = ~n8433 & n8846;
  assign n8849 = ~n8847 & ~n8848;
  assign n8850 = ~po29  & n8843;
  assign n8851 = ~n8849 & ~n8850;
  assign n8852 = ~n8844 & ~n8851;
  assign n8853 = po30  & ~n8852;
  assign n8854 = ~po30  & ~n8844;
  assign n8855 = ~n8851 & n8854;
  assign n8856 = ~n8436 & ~n8437;
  assign n8857 = po21  & n8856;
  assign n8858 = ~n8442 & ~n8857;
  assign n8859 = n8442 & n8857;
  assign n8860 = ~n8858 & ~n8859;
  assign n8861 = ~n8855 & n8860;
  assign n8862 = ~n8853 & ~n8861;
  assign n8863 = po31  & ~n8862;
  assign n8864 = ~n8445 & ~n8447;
  assign n8865 = po21  & n8864;
  assign n8866 = n8452 & ~n8865;
  assign n8867 = ~n8452 & n8865;
  assign n8868 = ~n8866 & ~n8867;
  assign n8869 = ~po31  & n8862;
  assign n8870 = ~n8868 & ~n8869;
  assign n8871 = ~n8863 & ~n8870;
  assign n8872 = po32  & ~n8871;
  assign n8873 = ~n8455 & ~n8456;
  assign n8874 = po21  & n8873;
  assign n8875 = n8461 & ~n8874;
  assign n8876 = ~n8461 & n8874;
  assign n8877 = ~n8875 & ~n8876;
  assign n8878 = ~po32  & ~n8863;
  assign n8879 = ~n8870 & n8878;
  assign n8880 = ~n8877 & ~n8879;
  assign n8881 = ~n8872 & ~n8880;
  assign n8882 = po33  & ~n8881;
  assign n8883 = ~n8464 & ~n8466;
  assign n8884 = po21  & n8883;
  assign n8885 = n8471 & ~n8884;
  assign n8886 = ~n8471 & n8884;
  assign n8887 = ~n8885 & ~n8886;
  assign n8888 = ~po33  & n8881;
  assign n8889 = ~n8887 & ~n8888;
  assign n8890 = ~n8882 & ~n8889;
  assign n8891 = po34  & ~n8890;
  assign n8892 = ~po34  & ~n8882;
  assign n8893 = ~n8889 & n8892;
  assign n8894 = ~n8474 & po21 ;
  assign n8895 = ~n8480 & n8894;
  assign n8896 = n8479 & ~n8895;
  assign n8897 = n8481 & n8894;
  assign n8898 = ~n8896 & ~n8897;
  assign n8899 = ~n8893 & n8898;
  assign n8900 = ~n8891 & ~n8899;
  assign n8901 = po35  & ~n8900;
  assign n8902 = ~n8483 & ~n8485;
  assign n8903 = po21  & n8902;
  assign n8904 = n8490 & ~n8903;
  assign n8905 = ~n8490 & n8903;
  assign n8906 = ~n8904 & ~n8905;
  assign n8907 = ~po35  & n8900;
  assign n8908 = ~n8906 & ~n8907;
  assign n8909 = ~n8901 & ~n8908;
  assign n8910 = po36  & ~n8909;
  assign n8911 = ~n8493 & ~n8494;
  assign n8912 = po21  & n8911;
  assign n8913 = n8499 & ~n8912;
  assign n8914 = ~n8499 & n8912;
  assign n8915 = ~n8913 & ~n8914;
  assign n8916 = ~po36  & ~n8901;
  assign n8917 = ~n8908 & n8916;
  assign n8918 = ~n8915 & ~n8917;
  assign n8919 = ~n8910 & ~n8918;
  assign n8920 = po37  & ~n8919;
  assign n8921 = ~n8502 & ~n8504;
  assign n8922 = po21  & n8921;
  assign n8923 = n8509 & ~n8922;
  assign n8924 = ~n8509 & n8922;
  assign n8925 = ~n8923 & ~n8924;
  assign n8926 = ~po37  & n8919;
  assign n8927 = ~n8925 & ~n8926;
  assign n8928 = ~n8920 & ~n8927;
  assign n8929 = po38  & ~n8928;
  assign n8930 = ~po38  & ~n8920;
  assign n8931 = ~n8927 & n8930;
  assign n8932 = ~n8512 & po21 ;
  assign n8933 = ~n8518 & n8932;
  assign n8934 = n8517 & ~n8933;
  assign n8935 = n8519 & n8932;
  assign n8936 = ~n8934 & ~n8935;
  assign n8937 = ~n8931 & n8936;
  assign n8938 = ~n8929 & ~n8937;
  assign n8939 = po39  & ~n8938;
  assign n8940 = ~n8521 & ~n8523;
  assign n8941 = po21  & n8940;
  assign n8942 = n8528 & ~n8941;
  assign n8943 = ~n8528 & n8941;
  assign n8944 = ~n8942 & ~n8943;
  assign n8945 = ~po39  & n8938;
  assign n8946 = ~n8944 & ~n8945;
  assign n8947 = ~n8939 & ~n8946;
  assign n8948 = po40  & ~n8947;
  assign n8949 = ~n8531 & ~n8532;
  assign n8950 = po21  & n8949;
  assign n8951 = n8537 & ~n8950;
  assign n8952 = ~n8537 & n8950;
  assign n8953 = ~n8951 & ~n8952;
  assign n8954 = ~po40  & ~n8939;
  assign n8955 = ~n8946 & n8954;
  assign n8956 = ~n8953 & ~n8955;
  assign n8957 = ~n8948 & ~n8956;
  assign n8958 = ~po41  & n8957;
  assign n8959 = ~n8540 & po21 ;
  assign n8960 = ~n8547 & n8959;
  assign n8961 = n8545 & ~n8960;
  assign n8962 = n8548 & n8959;
  assign n8963 = ~n8961 & ~n8962;
  assign n8964 = ~n8958 & n8963;
  assign n8965 = po41  & ~n8957;
  assign n8966 = ~n8964 & ~n8965;
  assign n8967 = po42  & ~n8966;
  assign n8968 = ~n8550 & ~n8557;
  assign n8969 = po21  & n8968;
  assign n8970 = ~n8555 & ~n8969;
  assign n8971 = n8555 & n8969;
  assign n8972 = ~n8970 & ~n8971;
  assign n8973 = ~po42  & ~n8965;
  assign n8974 = ~n8964 & n8973;
  assign n8975 = n8972 & ~n8974;
  assign n8976 = ~n8967 & ~n8975;
  assign n8977 = ~po43  & n8976;
  assign n8978 = po43  & ~n8976;
  assign n8979 = ~n8774 & ~n8977;
  assign n8980 = ~n8978 & ~n8979;
  assign n8981 = po44  & ~n8980;
  assign n8982 = ~po44  & ~n8978;
  assign n8983 = ~n8979 & n8982;
  assign n8984 = ~n8564 & po21 ;
  assign n8985 = ~n8570 & n8984;
  assign n8986 = n8569 & ~n8985;
  assign n8987 = n8571 & n8984;
  assign n8988 = ~n8986 & ~n8987;
  assign n8989 = ~n8983 & n8988;
  assign n8990 = ~n8981 & ~n8989;
  assign n8991 = po45  & ~n8990;
  assign n8992 = ~n8573 & ~n8575;
  assign n8993 = po21  & n8992;
  assign n8994 = n8580 & ~n8993;
  assign n8995 = ~n8580 & n8993;
  assign n8996 = ~n8994 & ~n8995;
  assign n8997 = ~po45  & n8990;
  assign n8998 = ~n8996 & ~n8997;
  assign n8999 = ~n8991 & ~n8998;
  assign n9000 = po46  & ~n8999;
  assign n9001 = ~po46  & ~n8991;
  assign n9002 = ~n8998 & n9001;
  assign n9003 = ~n8583 & po21 ;
  assign n9004 = ~n8589 & n9003;
  assign n9005 = n8588 & ~n9004;
  assign n9006 = n8590 & n9003;
  assign n9007 = ~n9005 & ~n9006;
  assign n9008 = ~n9002 & n9007;
  assign n9009 = ~n9000 & ~n9008;
  assign n9010 = po47  & ~n9009;
  assign n9011 = ~n8592 & ~n8594;
  assign n9012 = po21  & n9011;
  assign n9013 = n8599 & ~n9012;
  assign n9014 = ~n8599 & n9012;
  assign n9015 = ~n9013 & ~n9014;
  assign n9016 = ~po47  & n9009;
  assign n9017 = ~n9015 & ~n9016;
  assign n9018 = ~n9010 & ~n9017;
  assign n9019 = po48  & ~n9018;
  assign n9020 = ~n8602 & ~n8603;
  assign n9021 = po21  & n9020;
  assign n9022 = n8608 & ~n9021;
  assign n9023 = ~n8608 & n9021;
  assign n9024 = ~n9022 & ~n9023;
  assign n9025 = ~po48  & ~n9010;
  assign n9026 = ~n9017 & n9025;
  assign n9027 = ~n9024 & ~n9026;
  assign n9028 = ~n9019 & ~n9027;
  assign n9029 = po49  & ~n9028;
  assign n9030 = ~n8611 & ~n8613;
  assign n9031 = po21  & n9030;
  assign n9032 = n8618 & ~n9031;
  assign n9033 = ~n8618 & n9031;
  assign n9034 = ~n9032 & ~n9033;
  assign n9035 = ~po49  & n9028;
  assign n9036 = ~n9034 & ~n9035;
  assign n9037 = ~n9029 & ~n9036;
  assign n9038 = po50  & ~n9037;
  assign n9039 = ~po50  & ~n9029;
  assign n9040 = ~n9036 & n9039;
  assign n9041 = ~n8621 & po21 ;
  assign n9042 = ~n8627 & n9041;
  assign n9043 = n8626 & ~n9042;
  assign n9044 = n8628 & n9041;
  assign n9045 = ~n9043 & ~n9044;
  assign n9046 = ~n9040 & n9045;
  assign n9047 = ~n9038 & ~n9046;
  assign n9048 = po51  & ~n9047;
  assign n9049 = ~n8630 & ~n8632;
  assign n9050 = po21  & n9049;
  assign n9051 = n8637 & ~n9050;
  assign n9052 = ~n8637 & n9050;
  assign n9053 = ~n9051 & ~n9052;
  assign n9054 = ~po51  & n9047;
  assign n9055 = ~n9053 & ~n9054;
  assign n9056 = ~n9048 & ~n9055;
  assign n9057 = po52  & ~n9056;
  assign n9058 = ~n8640 & ~n8641;
  assign n9059 = po21  & n9058;
  assign n9060 = n8646 & ~n9059;
  assign n9061 = ~n8646 & n9059;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = ~po52  & ~n9048;
  assign n9064 = ~n9055 & n9063;
  assign n9065 = ~n9062 & ~n9064;
  assign n9066 = ~n9057 & ~n9065;
  assign n9067 = po53  & ~n9066;
  assign n9068 = ~n8649 & ~n8651;
  assign n9069 = po21  & n9068;
  assign n9070 = n8656 & ~n9069;
  assign n9071 = ~n8656 & n9069;
  assign n9072 = ~n9070 & ~n9071;
  assign n9073 = ~po53  & n9066;
  assign n9074 = ~n9072 & ~n9073;
  assign n9075 = ~n9067 & ~n9074;
  assign n9076 = po54  & ~n9075;
  assign n9077 = ~po54  & ~n9067;
  assign n9078 = ~n9074 & n9077;
  assign n9079 = ~n8659 & po21 ;
  assign n9080 = ~n8665 & n9079;
  assign n9081 = n8664 & ~n9080;
  assign n9082 = n8666 & n9079;
  assign n9083 = ~n9081 & ~n9082;
  assign n9084 = ~n9078 & n9083;
  assign n9085 = ~n9076 & ~n9084;
  assign n9086 = po55  & ~n9085;
  assign n9087 = ~n8668 & ~n8670;
  assign n9088 = po21  & n9087;
  assign n9089 = n8675 & ~n9088;
  assign n9090 = ~n8675 & n9088;
  assign n9091 = ~n9089 & ~n9090;
  assign n9092 = ~po55  & n9085;
  assign n9093 = ~n9091 & ~n9092;
  assign n9094 = ~n9086 & ~n9093;
  assign n9095 = po56  & ~n9094;
  assign n9096 = ~n8678 & ~n8679;
  assign n9097 = po21  & n9096;
  assign n9098 = n8684 & ~n9097;
  assign n9099 = ~n8684 & n9097;
  assign n9100 = ~n9098 & ~n9099;
  assign n9101 = ~po56  & ~n9086;
  assign n9102 = ~n9093 & n9101;
  assign n9103 = ~n9100 & ~n9102;
  assign n9104 = ~n9095 & ~n9103;
  assign n9105 = po57  & ~n9104;
  assign n9106 = ~n8687 & ~n8689;
  assign n9107 = po21  & n9106;
  assign n9108 = n8694 & ~n9107;
  assign n9109 = ~n8694 & n9107;
  assign n9110 = ~n9108 & ~n9109;
  assign n9111 = ~po57  & n9104;
  assign n9112 = ~n9110 & ~n9111;
  assign n9113 = ~n9105 & ~n9112;
  assign n9114 = po58  & ~n9113;
  assign n9115 = ~po58  & ~n9105;
  assign n9116 = ~n9112 & n9115;
  assign n9117 = ~n8697 & po21 ;
  assign n9118 = ~n8703 & n9117;
  assign n9119 = n8702 & ~n9118;
  assign n9120 = n8704 & n9117;
  assign n9121 = ~n9119 & ~n9120;
  assign n9122 = ~n9116 & n9121;
  assign n9123 = ~n9114 & ~n9122;
  assign n9124 = po59  & ~n9123;
  assign n9125 = ~n8706 & ~n8708;
  assign n9126 = po21  & n9125;
  assign n9127 = n8713 & ~n9126;
  assign n9128 = ~n8713 & n9126;
  assign n9129 = ~n9127 & ~n9128;
  assign n9130 = ~po59  & n9123;
  assign n9131 = ~n9129 & ~n9130;
  assign n9132 = ~n9124 & ~n9131;
  assign n9133 = po60  & ~n9132;
  assign n9134 = ~n8716 & ~n8717;
  assign n9135 = po21  & n9134;
  assign n9136 = n8722 & ~n9135;
  assign n9137 = ~n8722 & n9135;
  assign n9138 = ~n9136 & ~n9137;
  assign n9139 = ~po60  & ~n9124;
  assign n9140 = ~n9131 & n9139;
  assign n9141 = ~n9138 & ~n9140;
  assign n9142 = ~n9133 & ~n9141;
  assign n9143 = po61  & ~n9142;
  assign n9144 = ~n8725 & ~n8727;
  assign n9145 = po21  & n9144;
  assign n9146 = n8732 & ~n9145;
  assign n9147 = ~n8732 & n9145;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = ~po61  & n9142;
  assign n9150 = ~n9148 & ~n9149;
  assign n9151 = ~n9143 & ~n9150;
  assign n9152 = po62  & ~n9151;
  assign n9153 = ~po62  & ~n9143;
  assign n9154 = ~n9150 & n9153;
  assign n9155 = ~n8735 & po21 ;
  assign n9156 = ~n8741 & n9155;
  assign n9157 = n8740 & ~n9156;
  assign n9158 = n8742 & n9155;
  assign n9159 = ~n9157 & ~n9158;
  assign n9160 = ~n9154 & n9159;
  assign n9161 = ~n9152 & ~n9160;
  assign n9162 = n8762 & po21 ;
  assign n9163 = ~n8753 & n9162;
  assign n9164 = ~n8744 & ~n8746;
  assign n9165 = po21  & n9164;
  assign n9166 = n8751 & ~n9165;
  assign n9167 = ~n8751 & n9165;
  assign n9168 = ~n9166 & ~n9167;
  assign n9169 = ~n8766 & ~n9163;
  assign n9170 = ~n9168 & n9169;
  assign n9171 = ~n9161 & n9170;
  assign n9172 = ~po63  & ~n9171;
  assign n9173 = n9161 & n9168;
  assign n9174 = n8753 & ~n9162;
  assign n9175 = ~n8753 & n8762;
  assign n9176 = po63  & ~n9175;
  assign n9177 = ~n9174 & n9176;
  assign n9178 = ~n9173 & ~n9177;
  assign po20  = n9172 | ~n9178;
  assign n9180 = ~n8978 & po20 ;
  assign n9181 = ~n8977 & n9180;
  assign n9182 = n8774 & ~n9181;
  assign n9183 = n8979 & n9180;
  assign n9184 = ~n9182 & ~n9183;
  assign n9185 = ~n8967 & ~n8974;
  assign n9186 = po20  & n9185;
  assign n9187 = n8972 & ~n9186;
  assign n9188 = ~n8972 & n9186;
  assign n9189 = ~n9187 & ~n9188;
  assign n9190 = pi40  & po20 ;
  assign n9191 = ~pi38  & ~pi39 ;
  assign n9192 = ~pi40  & n9191;
  assign n9193 = ~n9190 & ~n9192;
  assign n9194 = po21  & ~n9193;
  assign n9195 = ~pi40  & po20 ;
  assign n9196 = pi41  & ~n9195;
  assign n9197 = ~pi41  & n9195;
  assign n9198 = ~n9196 & ~n9197;
  assign n9199 = ~po21  & n9193;
  assign n9200 = n9198 & ~n9199;
  assign n9201 = ~n9194 & ~n9200;
  assign n9202 = po22  & ~n9201;
  assign n9203 = ~po22  & ~n9194;
  assign n9204 = ~n9200 & n9203;
  assign n9205 = po21  & ~po20 ;
  assign n9206 = ~n9197 & ~n9205;
  assign n9207 = pi42  & ~n9206;
  assign n9208 = ~pi42  & n9206;
  assign n9209 = ~n9207 & ~n9208;
  assign n9210 = ~n9204 & ~n9209;
  assign n9211 = ~n9202 & ~n9210;
  assign n9212 = po23  & ~n9211;
  assign n9213 = ~po23  & n9211;
  assign n9214 = ~n8779 & ~n8780;
  assign n9215 = po20  & n9214;
  assign n9216 = n8784 & ~n9215;
  assign n9217 = ~n8784 & n9215;
  assign n9218 = ~n9216 & ~n9217;
  assign n9219 = ~n9213 & ~n9218;
  assign n9220 = ~n9212 & ~n9219;
  assign n9221 = po24  & ~n9220;
  assign n9222 = ~po24  & ~n9212;
  assign n9223 = ~n9219 & n9222;
  assign n9224 = ~n8787 & po20 ;
  assign n9225 = ~n8793 & n9224;
  assign n9226 = n8792 & ~n9225;
  assign n9227 = n8794 & n9224;
  assign n9228 = ~n9226 & ~n9227;
  assign n9229 = ~n9223 & n9228;
  assign n9230 = ~n9221 & ~n9229;
  assign n9231 = po25  & ~n9230;
  assign n9232 = ~po25  & n9230;
  assign n9233 = ~n8796 & ~n8798;
  assign n9234 = po20  & n9233;
  assign n9235 = n8803 & ~n9234;
  assign n9236 = ~n8803 & n9234;
  assign n9237 = ~n9235 & ~n9236;
  assign n9238 = ~n9232 & n9237;
  assign n9239 = ~n9231 & ~n9238;
  assign n9240 = po26  & ~n9239;
  assign n9241 = ~po26  & ~n9231;
  assign n9242 = ~n9238 & n9241;
  assign n9243 = ~n8806 & po20 ;
  assign n9244 = ~n8812 & n9243;
  assign n9245 = n8811 & ~n9244;
  assign n9246 = n8813 & n9243;
  assign n9247 = ~n9245 & ~n9246;
  assign n9248 = ~n9242 & n9247;
  assign n9249 = ~n9240 & ~n9248;
  assign n9250 = po27  & ~n9249;
  assign n9251 = ~po27  & n9249;
  assign n9252 = ~n8815 & ~n8817;
  assign n9253 = po20  & n9252;
  assign n9254 = n8822 & n9253;
  assign n9255 = ~n8822 & ~n9253;
  assign n9256 = ~n9254 & ~n9255;
  assign n9257 = ~n9251 & n9256;
  assign n9258 = ~n9250 & ~n9257;
  assign n9259 = po28  & ~n9258;
  assign n9260 = ~po28  & ~n9250;
  assign n9261 = ~n9257 & n9260;
  assign n9262 = ~n8825 & po20 ;
  assign n9263 = ~n8831 & n9262;
  assign n9264 = n8830 & ~n9263;
  assign n9265 = n8832 & n9262;
  assign n9266 = ~n9264 & ~n9265;
  assign n9267 = ~n9261 & n9266;
  assign n9268 = ~n9259 & ~n9267;
  assign n9269 = po29  & ~n9268;
  assign n9270 = ~po29  & n9268;
  assign n9271 = ~n8834 & ~n8836;
  assign n9272 = po20  & n9271;
  assign n9273 = ~n8841 & ~n9272;
  assign n9274 = n8841 & n9272;
  assign n9275 = ~n9273 & ~n9274;
  assign n9276 = ~n9270 & n9275;
  assign n9277 = ~n9269 & ~n9276;
  assign n9278 = po30  & ~n9277;
  assign n9279 = ~po30  & ~n9269;
  assign n9280 = ~n9276 & n9279;
  assign n9281 = ~n8844 & po20 ;
  assign n9282 = ~n8850 & n9281;
  assign n9283 = n8849 & ~n9282;
  assign n9284 = n8851 & n9281;
  assign n9285 = ~n9283 & ~n9284;
  assign n9286 = ~n9280 & n9285;
  assign n9287 = ~n9278 & ~n9286;
  assign n9288 = po31  & ~n9287;
  assign n9289 = ~n8853 & ~n8855;
  assign n9290 = po20  & n9289;
  assign n9291 = n8860 & ~n9290;
  assign n9292 = ~n8860 & n9290;
  assign n9293 = ~n9291 & ~n9292;
  assign n9294 = ~po31  & n9287;
  assign n9295 = ~n9293 & ~n9294;
  assign n9296 = ~n9288 & ~n9295;
  assign n9297 = po32  & ~n9296;
  assign n9298 = ~po32  & ~n9288;
  assign n9299 = ~n9295 & n9298;
  assign n9300 = ~n8863 & po20 ;
  assign n9301 = ~n8869 & n9300;
  assign n9302 = n8868 & ~n9301;
  assign n9303 = n8870 & n9300;
  assign n9304 = ~n9302 & ~n9303;
  assign n9305 = ~n9299 & n9304;
  assign n9306 = ~n9297 & ~n9305;
  assign n9307 = po33  & ~n9306;
  assign n9308 = ~po33  & n9306;
  assign n9309 = ~n8872 & po20 ;
  assign n9310 = ~n8879 & n9309;
  assign n9311 = n8877 & ~n9310;
  assign n9312 = n8880 & n9309;
  assign n9313 = ~n9311 & ~n9312;
  assign n9314 = ~n9308 & n9313;
  assign n9315 = ~n9307 & ~n9314;
  assign n9316 = po34  & ~n9315;
  assign n9317 = ~po34  & ~n9307;
  assign n9318 = ~n9314 & n9317;
  assign n9319 = ~n8882 & po20 ;
  assign n9320 = ~n8888 & n9319;
  assign n9321 = n8887 & ~n9320;
  assign n9322 = n8889 & n9319;
  assign n9323 = ~n9321 & ~n9322;
  assign n9324 = ~n9318 & n9323;
  assign n9325 = ~n9316 & ~n9324;
  assign n9326 = po35  & ~n9325;
  assign n9327 = ~n8891 & ~n8893;
  assign n9328 = po20  & n9327;
  assign n9329 = n8898 & ~n9328;
  assign n9330 = ~n8898 & n9328;
  assign n9331 = ~n9329 & ~n9330;
  assign n9332 = ~po35  & n9325;
  assign n9333 = ~n9331 & ~n9332;
  assign n9334 = ~n9326 & ~n9333;
  assign n9335 = po36  & ~n9334;
  assign n9336 = ~po36  & ~n9326;
  assign n9337 = ~n9333 & n9336;
  assign n9338 = ~n8901 & po20 ;
  assign n9339 = ~n8907 & n9338;
  assign n9340 = n8906 & ~n9339;
  assign n9341 = n8908 & n9338;
  assign n9342 = ~n9340 & ~n9341;
  assign n9343 = ~n9337 & n9342;
  assign n9344 = ~n9335 & ~n9343;
  assign n9345 = po37  & ~n9344;
  assign n9346 = ~po37  & n9344;
  assign n9347 = ~n8910 & po20 ;
  assign n9348 = ~n8917 & n9347;
  assign n9349 = n8915 & ~n9348;
  assign n9350 = n8918 & n9347;
  assign n9351 = ~n9349 & ~n9350;
  assign n9352 = ~n9346 & n9351;
  assign n9353 = ~n9345 & ~n9352;
  assign n9354 = po38  & ~n9353;
  assign n9355 = ~po38  & ~n9345;
  assign n9356 = ~n9352 & n9355;
  assign n9357 = ~n8920 & po20 ;
  assign n9358 = ~n8926 & n9357;
  assign n9359 = n8925 & ~n9358;
  assign n9360 = n8927 & n9357;
  assign n9361 = ~n9359 & ~n9360;
  assign n9362 = ~n9356 & n9361;
  assign n9363 = ~n9354 & ~n9362;
  assign n9364 = po39  & ~n9363;
  assign n9365 = ~n8929 & ~n8931;
  assign n9366 = po20  & n9365;
  assign n9367 = n8936 & ~n9366;
  assign n9368 = ~n8936 & n9366;
  assign n9369 = ~n9367 & ~n9368;
  assign n9370 = ~po39  & n9363;
  assign n9371 = ~n9369 & ~n9370;
  assign n9372 = ~n9364 & ~n9371;
  assign n9373 = po40  & ~n9372;
  assign n9374 = ~po40  & ~n9364;
  assign n9375 = ~n9371 & n9374;
  assign n9376 = ~n8939 & po20 ;
  assign n9377 = ~n8945 & n9376;
  assign n9378 = n8944 & ~n9377;
  assign n9379 = n8946 & n9376;
  assign n9380 = ~n9378 & ~n9379;
  assign n9381 = ~n9375 & n9380;
  assign n9382 = ~n9373 & ~n9381;
  assign n9383 = po41  & ~n9382;
  assign n9384 = ~po41  & n9382;
  assign n9385 = ~n8948 & po20 ;
  assign n9386 = ~n8955 & n9385;
  assign n9387 = n8953 & ~n9386;
  assign n9388 = n8956 & n9385;
  assign n9389 = ~n9387 & ~n9388;
  assign n9390 = ~n9384 & n9389;
  assign n9391 = ~n9383 & ~n9390;
  assign n9392 = po42  & ~n9391;
  assign n9393 = ~n8958 & ~n8965;
  assign n9394 = po20  & n9393;
  assign n9395 = n8963 & ~n9394;
  assign n9396 = ~n8963 & n9394;
  assign n9397 = ~n9395 & ~n9396;
  assign n9398 = ~po42  & ~n9383;
  assign n9399 = ~n9390 & n9398;
  assign n9400 = ~n9397 & ~n9399;
  assign n9401 = ~n9392 & ~n9400;
  assign n9402 = ~po43  & n9401;
  assign n9403 = ~n9189 & ~n9402;
  assign n9404 = po43  & ~n9401;
  assign n9405 = ~po44  & ~n9404;
  assign n9406 = ~n9403 & n9405;
  assign n9407 = ~n9403 & ~n9404;
  assign n9408 = po44  & ~n9407;
  assign n9409 = n9184 & ~n9406;
  assign n9410 = ~n9408 & ~n9409;
  assign n9411 = po45  & ~n9410;
  assign n9412 = ~n8981 & ~n8983;
  assign n9413 = po20  & n9412;
  assign n9414 = n8988 & ~n9413;
  assign n9415 = ~n8988 & n9413;
  assign n9416 = ~n9414 & ~n9415;
  assign n9417 = ~po45  & n9410;
  assign n9418 = ~n9416 & ~n9417;
  assign n9419 = ~n9411 & ~n9418;
  assign n9420 = po46  & ~n9419;
  assign n9421 = ~po46  & ~n9411;
  assign n9422 = ~n9418 & n9421;
  assign n9423 = ~n8991 & po20 ;
  assign n9424 = ~n8997 & n9423;
  assign n9425 = n8996 & ~n9424;
  assign n9426 = n8998 & n9423;
  assign n9427 = ~n9425 & ~n9426;
  assign n9428 = ~n9422 & n9427;
  assign n9429 = ~n9420 & ~n9428;
  assign n9430 = po47  & ~n9429;
  assign n9431 = ~n9000 & ~n9002;
  assign n9432 = po20  & n9431;
  assign n9433 = n9007 & ~n9432;
  assign n9434 = ~n9007 & n9432;
  assign n9435 = ~n9433 & ~n9434;
  assign n9436 = ~po47  & n9429;
  assign n9437 = ~n9435 & ~n9436;
  assign n9438 = ~n9430 & ~n9437;
  assign n9439 = po48  & ~n9438;
  assign n9440 = ~po48  & ~n9430;
  assign n9441 = ~n9437 & n9440;
  assign n9442 = ~n9010 & po20 ;
  assign n9443 = ~n9016 & n9442;
  assign n9444 = n9015 & ~n9443;
  assign n9445 = n9017 & n9442;
  assign n9446 = ~n9444 & ~n9445;
  assign n9447 = ~n9441 & n9446;
  assign n9448 = ~n9439 & ~n9447;
  assign n9449 = po49  & ~n9448;
  assign n9450 = ~po49  & n9448;
  assign n9451 = ~n9019 & po20 ;
  assign n9452 = ~n9026 & n9451;
  assign n9453 = n9024 & ~n9452;
  assign n9454 = n9027 & n9451;
  assign n9455 = ~n9453 & ~n9454;
  assign n9456 = ~n9450 & n9455;
  assign n9457 = ~n9449 & ~n9456;
  assign n9458 = po50  & ~n9457;
  assign n9459 = ~po50  & ~n9449;
  assign n9460 = ~n9456 & n9459;
  assign n9461 = ~n9029 & po20 ;
  assign n9462 = ~n9035 & n9461;
  assign n9463 = n9034 & ~n9462;
  assign n9464 = n9036 & n9461;
  assign n9465 = ~n9463 & ~n9464;
  assign n9466 = ~n9460 & n9465;
  assign n9467 = ~n9458 & ~n9466;
  assign n9468 = po51  & ~n9467;
  assign n9469 = ~n9038 & ~n9040;
  assign n9470 = po20  & n9469;
  assign n9471 = n9045 & ~n9470;
  assign n9472 = ~n9045 & n9470;
  assign n9473 = ~n9471 & ~n9472;
  assign n9474 = ~po51  & n9467;
  assign n9475 = ~n9473 & ~n9474;
  assign n9476 = ~n9468 & ~n9475;
  assign n9477 = po52  & ~n9476;
  assign n9478 = ~po52  & ~n9468;
  assign n9479 = ~n9475 & n9478;
  assign n9480 = ~n9048 & po20 ;
  assign n9481 = ~n9054 & n9480;
  assign n9482 = n9053 & ~n9481;
  assign n9483 = n9055 & n9480;
  assign n9484 = ~n9482 & ~n9483;
  assign n9485 = ~n9479 & n9484;
  assign n9486 = ~n9477 & ~n9485;
  assign n9487 = po53  & ~n9486;
  assign n9488 = ~po53  & n9486;
  assign n9489 = ~n9057 & po20 ;
  assign n9490 = ~n9064 & n9489;
  assign n9491 = n9062 & ~n9490;
  assign n9492 = n9065 & n9489;
  assign n9493 = ~n9491 & ~n9492;
  assign n9494 = ~n9488 & n9493;
  assign n9495 = ~n9487 & ~n9494;
  assign n9496 = po54  & ~n9495;
  assign n9497 = ~po54  & ~n9487;
  assign n9498 = ~n9494 & n9497;
  assign n9499 = ~n9067 & po20 ;
  assign n9500 = ~n9073 & n9499;
  assign n9501 = n9072 & ~n9500;
  assign n9502 = n9074 & n9499;
  assign n9503 = ~n9501 & ~n9502;
  assign n9504 = ~n9498 & n9503;
  assign n9505 = ~n9496 & ~n9504;
  assign n9506 = po55  & ~n9505;
  assign n9507 = ~n9076 & ~n9078;
  assign n9508 = po20  & n9507;
  assign n9509 = n9083 & ~n9508;
  assign n9510 = ~n9083 & n9508;
  assign n9511 = ~n9509 & ~n9510;
  assign n9512 = ~po55  & n9505;
  assign n9513 = ~n9511 & ~n9512;
  assign n9514 = ~n9506 & ~n9513;
  assign n9515 = po56  & ~n9514;
  assign n9516 = ~po56  & ~n9506;
  assign n9517 = ~n9513 & n9516;
  assign n9518 = ~n9086 & po20 ;
  assign n9519 = ~n9092 & n9518;
  assign n9520 = n9091 & ~n9519;
  assign n9521 = n9093 & n9518;
  assign n9522 = ~n9520 & ~n9521;
  assign n9523 = ~n9517 & n9522;
  assign n9524 = ~n9515 & ~n9523;
  assign n9525 = po57  & ~n9524;
  assign n9526 = ~po57  & n9524;
  assign n9527 = ~n9095 & po20 ;
  assign n9528 = ~n9102 & n9527;
  assign n9529 = n9100 & ~n9528;
  assign n9530 = n9103 & n9527;
  assign n9531 = ~n9529 & ~n9530;
  assign n9532 = ~n9526 & n9531;
  assign n9533 = ~n9525 & ~n9532;
  assign n9534 = po58  & ~n9533;
  assign n9535 = ~po58  & ~n9525;
  assign n9536 = ~n9532 & n9535;
  assign n9537 = ~n9105 & po20 ;
  assign n9538 = ~n9111 & n9537;
  assign n9539 = n9110 & ~n9538;
  assign n9540 = n9112 & n9537;
  assign n9541 = ~n9539 & ~n9540;
  assign n9542 = ~n9536 & n9541;
  assign n9543 = ~n9534 & ~n9542;
  assign n9544 = po59  & ~n9543;
  assign n9545 = ~n9114 & ~n9116;
  assign n9546 = po20  & n9545;
  assign n9547 = n9121 & ~n9546;
  assign n9548 = ~n9121 & n9546;
  assign n9549 = ~n9547 & ~n9548;
  assign n9550 = ~po59  & n9543;
  assign n9551 = ~n9549 & ~n9550;
  assign n9552 = ~n9544 & ~n9551;
  assign n9553 = po60  & ~n9552;
  assign n9554 = ~po60  & ~n9544;
  assign n9555 = ~n9551 & n9554;
  assign n9556 = ~n9124 & po20 ;
  assign n9557 = ~n9130 & n9556;
  assign n9558 = n9129 & ~n9557;
  assign n9559 = n9131 & n9556;
  assign n9560 = ~n9558 & ~n9559;
  assign n9561 = ~n9555 & n9560;
  assign n9562 = ~n9553 & ~n9561;
  assign n9563 = po61  & ~n9562;
  assign n9564 = ~po61  & n9562;
  assign n9565 = ~n9133 & po20 ;
  assign n9566 = ~n9140 & n9565;
  assign n9567 = n9138 & ~n9566;
  assign n9568 = n9141 & n9565;
  assign n9569 = ~n9567 & ~n9568;
  assign n9570 = ~n9564 & n9569;
  assign n9571 = ~n9563 & ~n9570;
  assign n9572 = po62  & ~n9571;
  assign n9573 = ~po62  & ~n9563;
  assign n9574 = ~n9570 & n9573;
  assign n9575 = ~n9143 & po20 ;
  assign n9576 = ~n9149 & n9575;
  assign n9577 = n9148 & ~n9576;
  assign n9578 = n9150 & n9575;
  assign n9579 = ~n9577 & ~n9578;
  assign n9580 = ~n9574 & n9579;
  assign n9581 = ~n9572 & ~n9580;
  assign n9582 = ~n9152 & ~n9154;
  assign n9583 = po20  & n9582;
  assign n9584 = n9159 & ~n9583;
  assign n9585 = ~n9159 & n9583;
  assign n9586 = ~n9584 & ~n9585;
  assign n9587 = n9161 & po20 ;
  assign n9588 = ~n9168 & ~n9587;
  assign n9589 = ~n9173 & ~n9588;
  assign n9590 = po20  & ~n9589;
  assign n9591 = ~n9586 & ~n9590;
  assign n9592 = ~n9581 & n9591;
  assign n9593 = ~po63  & ~n9592;
  assign n9594 = n9581 & n9586;
  assign n9595 = po63  & n9589;
  assign n9596 = ~n9594 & ~n9595;
  assign po19  = n9593 | ~n9596;
  assign n9598 = ~n9406 & ~n9408;
  assign n9599 = po19  & n9598;
  assign n9600 = n9184 & ~n9599;
  assign n9601 = ~n9184 & n9599;
  assign n9602 = ~n9600 & ~n9601;
  assign n9603 = pi38  & po19 ;
  assign n9604 = ~pi36  & ~pi37 ;
  assign n9605 = ~pi38  & n9604;
  assign n9606 = ~n9603 & ~n9605;
  assign n9607 = po20  & ~n9606;
  assign n9608 = ~po20  & n9606;
  assign n9609 = ~pi38  & po19 ;
  assign n9610 = pi39  & ~n9609;
  assign n9611 = ~pi39  & n9609;
  assign n9612 = ~n9610 & ~n9611;
  assign n9613 = ~n9608 & n9612;
  assign n9614 = ~n9607 & ~n9613;
  assign n9615 = po21  & ~n9614;
  assign n9616 = po20  & ~po19 ;
  assign n9617 = ~n9611 & ~n9616;
  assign n9618 = pi40  & ~n9617;
  assign n9619 = ~pi40  & n9617;
  assign n9620 = ~n9618 & ~n9619;
  assign n9621 = ~po21  & n9614;
  assign n9622 = ~n9620 & ~n9621;
  assign n9623 = ~n9615 & ~n9622;
  assign n9624 = po22  & ~n9623;
  assign n9625 = ~po22  & ~n9615;
  assign n9626 = ~n9622 & n9625;
  assign n9627 = ~n9194 & ~n9199;
  assign n9628 = po19  & n9627;
  assign n9629 = n9198 & ~n9628;
  assign n9630 = ~n9198 & n9628;
  assign n9631 = ~n9629 & ~n9630;
  assign n9632 = ~n9626 & ~n9631;
  assign n9633 = ~n9624 & ~n9632;
  assign n9634 = po23  & ~n9633;
  assign n9635 = ~n9202 & ~n9204;
  assign n9636 = po19  & n9635;
  assign n9637 = ~n9209 & ~n9636;
  assign n9638 = n9209 & n9636;
  assign n9639 = ~n9637 & ~n9638;
  assign n9640 = ~po23  & n9633;
  assign n9641 = ~n9639 & ~n9640;
  assign n9642 = ~n9634 & ~n9641;
  assign n9643 = po24  & ~n9642;
  assign n9644 = ~po24  & ~n9634;
  assign n9645 = ~n9641 & n9644;
  assign n9646 = ~n9212 & ~n9213;
  assign n9647 = po19  & n9646;
  assign n9648 = n9218 & ~n9647;
  assign n9649 = ~n9218 & n9647;
  assign n9650 = ~n9648 & ~n9649;
  assign n9651 = ~n9645 & n9650;
  assign n9652 = ~n9643 & ~n9651;
  assign n9653 = po25  & ~n9652;
  assign n9654 = ~n9221 & ~n9223;
  assign n9655 = po19  & n9654;
  assign n9656 = n9228 & ~n9655;
  assign n9657 = ~n9228 & n9655;
  assign n9658 = ~n9656 & ~n9657;
  assign n9659 = ~po25  & n9652;
  assign n9660 = ~n9658 & ~n9659;
  assign n9661 = ~n9653 & ~n9660;
  assign n9662 = po26  & ~n9661;
  assign n9663 = ~po26  & ~n9653;
  assign n9664 = ~n9660 & n9663;
  assign n9665 = ~n9231 & ~n9232;
  assign n9666 = po19  & n9665;
  assign n9667 = n9237 & n9666;
  assign n9668 = ~n9237 & ~n9666;
  assign n9669 = ~n9667 & ~n9668;
  assign n9670 = ~n9664 & n9669;
  assign n9671 = ~n9662 & ~n9670;
  assign n9672 = po27  & ~n9671;
  assign n9673 = ~n9240 & ~n9242;
  assign n9674 = po19  & n9673;
  assign n9675 = n9247 & ~n9674;
  assign n9676 = ~n9247 & n9674;
  assign n9677 = ~n9675 & ~n9676;
  assign n9678 = ~po27  & n9671;
  assign n9679 = ~n9677 & ~n9678;
  assign n9680 = ~n9672 & ~n9679;
  assign n9681 = po28  & ~n9680;
  assign n9682 = ~po28  & ~n9672;
  assign n9683 = ~n9679 & n9682;
  assign n9684 = ~n9250 & ~n9251;
  assign n9685 = po19  & n9684;
  assign n9686 = ~n9256 & ~n9685;
  assign n9687 = n9256 & n9685;
  assign n9688 = ~n9686 & ~n9687;
  assign n9689 = ~n9683 & n9688;
  assign n9690 = ~n9681 & ~n9689;
  assign n9691 = po29  & ~n9690;
  assign n9692 = ~n9259 & ~n9261;
  assign n9693 = po19  & n9692;
  assign n9694 = n9266 & ~n9693;
  assign n9695 = ~n9266 & n9693;
  assign n9696 = ~n9694 & ~n9695;
  assign n9697 = ~po29  & n9690;
  assign n9698 = ~n9696 & ~n9697;
  assign n9699 = ~n9691 & ~n9698;
  assign n9700 = po30  & ~n9699;
  assign n9701 = ~n9269 & ~n9270;
  assign n9702 = po19  & n9701;
  assign n9703 = n9275 & ~n9702;
  assign n9704 = ~n9275 & n9702;
  assign n9705 = ~n9703 & ~n9704;
  assign n9706 = ~po30  & ~n9691;
  assign n9707 = ~n9698 & n9706;
  assign n9708 = ~n9705 & ~n9707;
  assign n9709 = ~n9700 & ~n9708;
  assign n9710 = po31  & ~n9709;
  assign n9711 = ~n9278 & ~n9280;
  assign n9712 = po19  & n9711;
  assign n9713 = n9285 & ~n9712;
  assign n9714 = ~n9285 & n9712;
  assign n9715 = ~n9713 & ~n9714;
  assign n9716 = ~po31  & n9709;
  assign n9717 = ~n9715 & ~n9716;
  assign n9718 = ~n9710 & ~n9717;
  assign n9719 = po32  & ~n9718;
  assign n9720 = ~po32  & ~n9710;
  assign n9721 = ~n9717 & n9720;
  assign n9722 = ~n9288 & po19 ;
  assign n9723 = ~n9294 & n9722;
  assign n9724 = n9293 & ~n9723;
  assign n9725 = n9295 & n9722;
  assign n9726 = ~n9724 & ~n9725;
  assign n9727 = ~n9721 & n9726;
  assign n9728 = ~n9719 & ~n9727;
  assign n9729 = po33  & ~n9728;
  assign n9730 = ~n9297 & ~n9299;
  assign n9731 = po19  & n9730;
  assign n9732 = n9304 & ~n9731;
  assign n9733 = ~n9304 & n9731;
  assign n9734 = ~n9732 & ~n9733;
  assign n9735 = ~po33  & n9728;
  assign n9736 = ~n9734 & ~n9735;
  assign n9737 = ~n9729 & ~n9736;
  assign n9738 = po34  & ~n9737;
  assign n9739 = ~n9307 & ~n9308;
  assign n9740 = po19  & n9739;
  assign n9741 = n9313 & ~n9740;
  assign n9742 = ~n9313 & n9740;
  assign n9743 = ~n9741 & ~n9742;
  assign n9744 = ~po34  & ~n9729;
  assign n9745 = ~n9736 & n9744;
  assign n9746 = ~n9743 & ~n9745;
  assign n9747 = ~n9738 & ~n9746;
  assign n9748 = po35  & ~n9747;
  assign n9749 = ~n9316 & ~n9318;
  assign n9750 = po19  & n9749;
  assign n9751 = n9323 & ~n9750;
  assign n9752 = ~n9323 & n9750;
  assign n9753 = ~n9751 & ~n9752;
  assign n9754 = ~po35  & n9747;
  assign n9755 = ~n9753 & ~n9754;
  assign n9756 = ~n9748 & ~n9755;
  assign n9757 = po36  & ~n9756;
  assign n9758 = ~po36  & ~n9748;
  assign n9759 = ~n9755 & n9758;
  assign n9760 = ~n9326 & po19 ;
  assign n9761 = ~n9332 & n9760;
  assign n9762 = n9331 & ~n9761;
  assign n9763 = n9333 & n9760;
  assign n9764 = ~n9762 & ~n9763;
  assign n9765 = ~n9759 & n9764;
  assign n9766 = ~n9757 & ~n9765;
  assign n9767 = po37  & ~n9766;
  assign n9768 = ~n9335 & ~n9337;
  assign n9769 = po19  & n9768;
  assign n9770 = n9342 & ~n9769;
  assign n9771 = ~n9342 & n9769;
  assign n9772 = ~n9770 & ~n9771;
  assign n9773 = ~po37  & n9766;
  assign n9774 = ~n9772 & ~n9773;
  assign n9775 = ~n9767 & ~n9774;
  assign n9776 = po38  & ~n9775;
  assign n9777 = ~n9345 & ~n9346;
  assign n9778 = po19  & n9777;
  assign n9779 = n9351 & ~n9778;
  assign n9780 = ~n9351 & n9778;
  assign n9781 = ~n9779 & ~n9780;
  assign n9782 = ~po38  & ~n9767;
  assign n9783 = ~n9774 & n9782;
  assign n9784 = ~n9781 & ~n9783;
  assign n9785 = ~n9776 & ~n9784;
  assign n9786 = po39  & ~n9785;
  assign n9787 = ~n9354 & ~n9356;
  assign n9788 = po19  & n9787;
  assign n9789 = n9361 & ~n9788;
  assign n9790 = ~n9361 & n9788;
  assign n9791 = ~n9789 & ~n9790;
  assign n9792 = ~po39  & n9785;
  assign n9793 = ~n9791 & ~n9792;
  assign n9794 = ~n9786 & ~n9793;
  assign n9795 = po40  & ~n9794;
  assign n9796 = ~po40  & ~n9786;
  assign n9797 = ~n9793 & n9796;
  assign n9798 = ~n9364 & po19 ;
  assign n9799 = ~n9370 & n9798;
  assign n9800 = n9369 & ~n9799;
  assign n9801 = n9371 & n9798;
  assign n9802 = ~n9800 & ~n9801;
  assign n9803 = ~n9797 & n9802;
  assign n9804 = ~n9795 & ~n9803;
  assign n9805 = po41  & ~n9804;
  assign n9806 = ~n9373 & ~n9375;
  assign n9807 = po19  & n9806;
  assign n9808 = n9380 & ~n9807;
  assign n9809 = ~n9380 & n9807;
  assign n9810 = ~n9808 & ~n9809;
  assign n9811 = ~po41  & n9804;
  assign n9812 = ~n9810 & ~n9811;
  assign n9813 = ~n9805 & ~n9812;
  assign n9814 = po42  & ~n9813;
  assign n9815 = ~n9383 & ~n9384;
  assign n9816 = po19  & n9815;
  assign n9817 = n9389 & ~n9816;
  assign n9818 = ~n9389 & n9816;
  assign n9819 = ~n9817 & ~n9818;
  assign n9820 = ~po42  & ~n9805;
  assign n9821 = ~n9812 & n9820;
  assign n9822 = ~n9819 & ~n9821;
  assign n9823 = ~n9814 & ~n9822;
  assign n9824 = ~po43  & n9823;
  assign n9825 = ~n9392 & po19 ;
  assign n9826 = ~n9399 & n9825;
  assign n9827 = n9397 & ~n9826;
  assign n9828 = n9400 & n9825;
  assign n9829 = ~n9827 & ~n9828;
  assign n9830 = ~n9824 & n9829;
  assign n9831 = po43  & ~n9823;
  assign n9832 = ~n9830 & ~n9831;
  assign n9833 = po44  & ~n9832;
  assign n9834 = ~po44  & ~n9831;
  assign n9835 = ~n9830 & n9834;
  assign n9836 = ~n9402 & ~n9404;
  assign n9837 = po19  & n9836;
  assign n9838 = n9189 & n9837;
  assign n9839 = ~n9189 & ~n9837;
  assign n9840 = ~n9838 & ~n9839;
  assign n9841 = ~n9835 & ~n9840;
  assign n9842 = ~n9833 & ~n9841;
  assign n9843 = ~po45  & n9842;
  assign n9844 = po45  & ~n9842;
  assign n9845 = ~n9602 & ~n9843;
  assign n9846 = ~n9844 & ~n9845;
  assign n9847 = po46  & ~n9846;
  assign n9848 = ~po46  & ~n9844;
  assign n9849 = ~n9845 & n9848;
  assign n9850 = ~n9411 & po19 ;
  assign n9851 = ~n9417 & n9850;
  assign n9852 = n9416 & ~n9851;
  assign n9853 = n9418 & n9850;
  assign n9854 = ~n9852 & ~n9853;
  assign n9855 = ~n9849 & n9854;
  assign n9856 = ~n9847 & ~n9855;
  assign n9857 = po47  & ~n9856;
  assign n9858 = ~n9420 & ~n9422;
  assign n9859 = po19  & n9858;
  assign n9860 = n9427 & ~n9859;
  assign n9861 = ~n9427 & n9859;
  assign n9862 = ~n9860 & ~n9861;
  assign n9863 = ~po47  & n9856;
  assign n9864 = ~n9862 & ~n9863;
  assign n9865 = ~n9857 & ~n9864;
  assign n9866 = po48  & ~n9865;
  assign n9867 = ~po48  & ~n9857;
  assign n9868 = ~n9864 & n9867;
  assign n9869 = ~n9430 & po19 ;
  assign n9870 = ~n9436 & n9869;
  assign n9871 = n9435 & ~n9870;
  assign n9872 = n9437 & n9869;
  assign n9873 = ~n9871 & ~n9872;
  assign n9874 = ~n9868 & n9873;
  assign n9875 = ~n9866 & ~n9874;
  assign n9876 = po49  & ~n9875;
  assign n9877 = ~n9439 & ~n9441;
  assign n9878 = po19  & n9877;
  assign n9879 = n9446 & ~n9878;
  assign n9880 = ~n9446 & n9878;
  assign n9881 = ~n9879 & ~n9880;
  assign n9882 = ~po49  & n9875;
  assign n9883 = ~n9881 & ~n9882;
  assign n9884 = ~n9876 & ~n9883;
  assign n9885 = po50  & ~n9884;
  assign n9886 = ~n9449 & ~n9450;
  assign n9887 = po19  & n9886;
  assign n9888 = n9455 & ~n9887;
  assign n9889 = ~n9455 & n9887;
  assign n9890 = ~n9888 & ~n9889;
  assign n9891 = ~po50  & ~n9876;
  assign n9892 = ~n9883 & n9891;
  assign n9893 = ~n9890 & ~n9892;
  assign n9894 = ~n9885 & ~n9893;
  assign n9895 = po51  & ~n9894;
  assign n9896 = ~n9458 & ~n9460;
  assign n9897 = po19  & n9896;
  assign n9898 = n9465 & ~n9897;
  assign n9899 = ~n9465 & n9897;
  assign n9900 = ~n9898 & ~n9899;
  assign n9901 = ~po51  & n9894;
  assign n9902 = ~n9900 & ~n9901;
  assign n9903 = ~n9895 & ~n9902;
  assign n9904 = po52  & ~n9903;
  assign n9905 = ~po52  & ~n9895;
  assign n9906 = ~n9902 & n9905;
  assign n9907 = ~n9468 & po19 ;
  assign n9908 = ~n9474 & n9907;
  assign n9909 = n9473 & ~n9908;
  assign n9910 = n9475 & n9907;
  assign n9911 = ~n9909 & ~n9910;
  assign n9912 = ~n9906 & n9911;
  assign n9913 = ~n9904 & ~n9912;
  assign n9914 = po53  & ~n9913;
  assign n9915 = ~n9477 & ~n9479;
  assign n9916 = po19  & n9915;
  assign n9917 = n9484 & ~n9916;
  assign n9918 = ~n9484 & n9916;
  assign n9919 = ~n9917 & ~n9918;
  assign n9920 = ~po53  & n9913;
  assign n9921 = ~n9919 & ~n9920;
  assign n9922 = ~n9914 & ~n9921;
  assign n9923 = po54  & ~n9922;
  assign n9924 = ~n9487 & ~n9488;
  assign n9925 = po19  & n9924;
  assign n9926 = n9493 & ~n9925;
  assign n9927 = ~n9493 & n9925;
  assign n9928 = ~n9926 & ~n9927;
  assign n9929 = ~po54  & ~n9914;
  assign n9930 = ~n9921 & n9929;
  assign n9931 = ~n9928 & ~n9930;
  assign n9932 = ~n9923 & ~n9931;
  assign n9933 = po55  & ~n9932;
  assign n9934 = ~n9496 & ~n9498;
  assign n9935 = po19  & n9934;
  assign n9936 = n9503 & ~n9935;
  assign n9937 = ~n9503 & n9935;
  assign n9938 = ~n9936 & ~n9937;
  assign n9939 = ~po55  & n9932;
  assign n9940 = ~n9938 & ~n9939;
  assign n9941 = ~n9933 & ~n9940;
  assign n9942 = po56  & ~n9941;
  assign n9943 = ~po56  & ~n9933;
  assign n9944 = ~n9940 & n9943;
  assign n9945 = ~n9506 & po19 ;
  assign n9946 = ~n9512 & n9945;
  assign n9947 = n9511 & ~n9946;
  assign n9948 = n9513 & n9945;
  assign n9949 = ~n9947 & ~n9948;
  assign n9950 = ~n9944 & n9949;
  assign n9951 = ~n9942 & ~n9950;
  assign n9952 = po57  & ~n9951;
  assign n9953 = ~n9515 & ~n9517;
  assign n9954 = po19  & n9953;
  assign n9955 = n9522 & ~n9954;
  assign n9956 = ~n9522 & n9954;
  assign n9957 = ~n9955 & ~n9956;
  assign n9958 = ~po57  & n9951;
  assign n9959 = ~n9957 & ~n9958;
  assign n9960 = ~n9952 & ~n9959;
  assign n9961 = po58  & ~n9960;
  assign n9962 = ~n9525 & ~n9526;
  assign n9963 = po19  & n9962;
  assign n9964 = n9531 & ~n9963;
  assign n9965 = ~n9531 & n9963;
  assign n9966 = ~n9964 & ~n9965;
  assign n9967 = ~po58  & ~n9952;
  assign n9968 = ~n9959 & n9967;
  assign n9969 = ~n9966 & ~n9968;
  assign n9970 = ~n9961 & ~n9969;
  assign n9971 = po59  & ~n9970;
  assign n9972 = ~n9534 & ~n9536;
  assign n9973 = po19  & n9972;
  assign n9974 = n9541 & ~n9973;
  assign n9975 = ~n9541 & n9973;
  assign n9976 = ~n9974 & ~n9975;
  assign n9977 = ~po59  & n9970;
  assign n9978 = ~n9976 & ~n9977;
  assign n9979 = ~n9971 & ~n9978;
  assign n9980 = po60  & ~n9979;
  assign n9981 = ~po60  & ~n9971;
  assign n9982 = ~n9978 & n9981;
  assign n9983 = ~n9544 & po19 ;
  assign n9984 = ~n9550 & n9983;
  assign n9985 = n9549 & ~n9984;
  assign n9986 = n9551 & n9983;
  assign n9987 = ~n9985 & ~n9986;
  assign n9988 = ~n9982 & n9987;
  assign n9989 = ~n9980 & ~n9988;
  assign n9990 = po61  & ~n9989;
  assign n9991 = ~n9553 & ~n9555;
  assign n9992 = po19  & n9991;
  assign n9993 = n9560 & ~n9992;
  assign n9994 = ~n9560 & n9992;
  assign n9995 = ~n9993 & ~n9994;
  assign n9996 = ~po61  & n9989;
  assign n9997 = ~n9995 & ~n9996;
  assign n9998 = ~n9990 & ~n9997;
  assign n9999 = po62  & ~n9998;
  assign n10000 = ~n9563 & ~n9564;
  assign n10001 = po19  & n10000;
  assign n10002 = n9569 & ~n10001;
  assign n10003 = ~n9569 & n10001;
  assign n10004 = ~n10002 & ~n10003;
  assign n10005 = ~po62  & ~n9990;
  assign n10006 = ~n9997 & n10005;
  assign n10007 = ~n10004 & ~n10006;
  assign n10008 = ~n9999 & ~n10007;
  assign n10009 = ~n9572 & ~n9574;
  assign n10010 = po19  & n10009;
  assign n10011 = n9579 & ~n10010;
  assign n10012 = ~n9579 & n10010;
  assign n10013 = ~n10011 & ~n10012;
  assign n10014 = n9581 & po19 ;
  assign n10015 = ~n9586 & ~n10014;
  assign n10016 = ~n9594 & ~n10015;
  assign n10017 = po19  & ~n10016;
  assign n10018 = ~n10013 & ~n10017;
  assign n10019 = ~n10008 & n10018;
  assign n10020 = ~po63  & ~n10019;
  assign n10021 = n10008 & n10013;
  assign n10022 = po63  & n10016;
  assign n10023 = ~n10021 & ~n10022;
  assign po18  = n10020 | ~n10023;
  assign n10025 = ~n9844 & po18 ;
  assign n10026 = ~n9843 & n10025;
  assign n10027 = n9602 & ~n10026;
  assign n10028 = n9845 & n10025;
  assign n10029 = ~n10027 & ~n10028;
  assign n10030 = ~n9833 & ~n9835;
  assign n10031 = po18  & n10030;
  assign n10032 = ~n9840 & ~n10031;
  assign n10033 = n9840 & n10031;
  assign n10034 = ~n10032 & ~n10033;
  assign n10035 = pi36  & po18 ;
  assign n10036 = ~pi34  & ~pi35 ;
  assign n10037 = ~pi36  & n10036;
  assign n10038 = ~n10035 & ~n10037;
  assign n10039 = po19  & ~n10038;
  assign n10040 = ~pi36  & po18 ;
  assign n10041 = pi37  & ~n10040;
  assign n10042 = ~pi37  & n10040;
  assign n10043 = ~n10041 & ~n10042;
  assign n10044 = ~po19  & n10038;
  assign n10045 = n10043 & ~n10044;
  assign n10046 = ~n10039 & ~n10045;
  assign n10047 = po20  & ~n10046;
  assign n10048 = ~po20  & ~n10039;
  assign n10049 = ~n10045 & n10048;
  assign n10050 = po19  & ~po18 ;
  assign n10051 = ~n10042 & ~n10050;
  assign n10052 = pi38  & ~n10051;
  assign n10053 = ~pi38  & n10051;
  assign n10054 = ~n10052 & ~n10053;
  assign n10055 = ~n10049 & ~n10054;
  assign n10056 = ~n10047 & ~n10055;
  assign n10057 = po21  & ~n10056;
  assign n10058 = ~po21  & n10056;
  assign n10059 = ~n9607 & ~n9608;
  assign n10060 = po18  & n10059;
  assign n10061 = n9612 & ~n10060;
  assign n10062 = ~n9612 & n10060;
  assign n10063 = ~n10061 & ~n10062;
  assign n10064 = ~n10058 & ~n10063;
  assign n10065 = ~n10057 & ~n10064;
  assign n10066 = po22  & ~n10065;
  assign n10067 = ~po22  & ~n10057;
  assign n10068 = ~n10064 & n10067;
  assign n10069 = ~n9615 & po18 ;
  assign n10070 = ~n9621 & n10069;
  assign n10071 = n9620 & ~n10070;
  assign n10072 = n9622 & n10069;
  assign n10073 = ~n10071 & ~n10072;
  assign n10074 = ~n10068 & n10073;
  assign n10075 = ~n10066 & ~n10074;
  assign n10076 = po23  & ~n10075;
  assign n10077 = ~po23  & n10075;
  assign n10078 = ~n9624 & ~n9626;
  assign n10079 = po18  & n10078;
  assign n10080 = n9631 & ~n10079;
  assign n10081 = ~n9631 & n10079;
  assign n10082 = ~n10080 & ~n10081;
  assign n10083 = ~n10077 & n10082;
  assign n10084 = ~n10076 & ~n10083;
  assign n10085 = po24  & ~n10084;
  assign n10086 = ~po24  & ~n10076;
  assign n10087 = ~n10083 & n10086;
  assign n10088 = ~n9634 & po18 ;
  assign n10089 = ~n9640 & n10088;
  assign n10090 = n9639 & ~n10089;
  assign n10091 = n9641 & n10088;
  assign n10092 = ~n10090 & ~n10091;
  assign n10093 = ~n10087 & n10092;
  assign n10094 = ~n10085 & ~n10093;
  assign n10095 = po25  & ~n10094;
  assign n10096 = ~po25  & n10094;
  assign n10097 = ~n9643 & ~n9645;
  assign n10098 = po18  & n10097;
  assign n10099 = n9650 & n10098;
  assign n10100 = ~n9650 & ~n10098;
  assign n10101 = ~n10099 & ~n10100;
  assign n10102 = ~n10096 & n10101;
  assign n10103 = ~n10095 & ~n10102;
  assign n10104 = po26  & ~n10103;
  assign n10105 = ~po26  & ~n10095;
  assign n10106 = ~n10102 & n10105;
  assign n10107 = ~n9653 & po18 ;
  assign n10108 = ~n9659 & n10107;
  assign n10109 = n9658 & ~n10108;
  assign n10110 = n9660 & n10107;
  assign n10111 = ~n10109 & ~n10110;
  assign n10112 = ~n10106 & n10111;
  assign n10113 = ~n10104 & ~n10112;
  assign n10114 = po27  & ~n10113;
  assign n10115 = ~po27  & n10113;
  assign n10116 = ~n9662 & ~n9664;
  assign n10117 = po18  & n10116;
  assign n10118 = ~n9669 & ~n10117;
  assign n10119 = n9669 & n10117;
  assign n10120 = ~n10118 & ~n10119;
  assign n10121 = ~n10115 & n10120;
  assign n10122 = ~n10114 & ~n10121;
  assign n10123 = po28  & ~n10122;
  assign n10124 = ~po28  & ~n10114;
  assign n10125 = ~n10121 & n10124;
  assign n10126 = ~n9672 & po18 ;
  assign n10127 = ~n9678 & n10126;
  assign n10128 = n9677 & ~n10127;
  assign n10129 = n9679 & n10126;
  assign n10130 = ~n10128 & ~n10129;
  assign n10131 = ~n10125 & n10130;
  assign n10132 = ~n10123 & ~n10131;
  assign n10133 = po29  & ~n10132;
  assign n10134 = ~n9681 & ~n9683;
  assign n10135 = po18  & n10134;
  assign n10136 = n9688 & ~n10135;
  assign n10137 = ~n9688 & n10135;
  assign n10138 = ~n10136 & ~n10137;
  assign n10139 = ~po29  & n10132;
  assign n10140 = ~n10138 & ~n10139;
  assign n10141 = ~n10133 & ~n10140;
  assign n10142 = po30  & ~n10141;
  assign n10143 = ~po30  & ~n10133;
  assign n10144 = ~n10140 & n10143;
  assign n10145 = ~n9691 & po18 ;
  assign n10146 = ~n9697 & n10145;
  assign n10147 = n9696 & ~n10146;
  assign n10148 = n9698 & n10145;
  assign n10149 = ~n10147 & ~n10148;
  assign n10150 = ~n10144 & n10149;
  assign n10151 = ~n10142 & ~n10150;
  assign n10152 = po31  & ~n10151;
  assign n10153 = ~po31  & n10151;
  assign n10154 = ~n9700 & po18 ;
  assign n10155 = ~n9707 & n10154;
  assign n10156 = n9705 & ~n10155;
  assign n10157 = n9708 & n10154;
  assign n10158 = ~n10156 & ~n10157;
  assign n10159 = ~n10153 & n10158;
  assign n10160 = ~n10152 & ~n10159;
  assign n10161 = po32  & ~n10160;
  assign n10162 = ~po32  & ~n10152;
  assign n10163 = ~n10159 & n10162;
  assign n10164 = ~n9710 & po18 ;
  assign n10165 = ~n9716 & n10164;
  assign n10166 = n9715 & ~n10165;
  assign n10167 = n9717 & n10164;
  assign n10168 = ~n10166 & ~n10167;
  assign n10169 = ~n10163 & n10168;
  assign n10170 = ~n10161 & ~n10169;
  assign n10171 = po33  & ~n10170;
  assign n10172 = ~n9719 & ~n9721;
  assign n10173 = po18  & n10172;
  assign n10174 = n9726 & ~n10173;
  assign n10175 = ~n9726 & n10173;
  assign n10176 = ~n10174 & ~n10175;
  assign n10177 = ~po33  & n10170;
  assign n10178 = ~n10176 & ~n10177;
  assign n10179 = ~n10171 & ~n10178;
  assign n10180 = po34  & ~n10179;
  assign n10181 = ~po34  & ~n10171;
  assign n10182 = ~n10178 & n10181;
  assign n10183 = ~n9729 & po18 ;
  assign n10184 = ~n9735 & n10183;
  assign n10185 = n9734 & ~n10184;
  assign n10186 = n9736 & n10183;
  assign n10187 = ~n10185 & ~n10186;
  assign n10188 = ~n10182 & n10187;
  assign n10189 = ~n10180 & ~n10188;
  assign n10190 = po35  & ~n10189;
  assign n10191 = ~po35  & n10189;
  assign n10192 = ~n9738 & po18 ;
  assign n10193 = ~n9745 & n10192;
  assign n10194 = n9743 & ~n10193;
  assign n10195 = n9746 & n10192;
  assign n10196 = ~n10194 & ~n10195;
  assign n10197 = ~n10191 & n10196;
  assign n10198 = ~n10190 & ~n10197;
  assign n10199 = po36  & ~n10198;
  assign n10200 = ~po36  & ~n10190;
  assign n10201 = ~n10197 & n10200;
  assign n10202 = ~n9748 & po18 ;
  assign n10203 = ~n9754 & n10202;
  assign n10204 = n9753 & ~n10203;
  assign n10205 = n9755 & n10202;
  assign n10206 = ~n10204 & ~n10205;
  assign n10207 = ~n10201 & n10206;
  assign n10208 = ~n10199 & ~n10207;
  assign n10209 = po37  & ~n10208;
  assign n10210 = ~n9757 & ~n9759;
  assign n10211 = po18  & n10210;
  assign n10212 = n9764 & ~n10211;
  assign n10213 = ~n9764 & n10211;
  assign n10214 = ~n10212 & ~n10213;
  assign n10215 = ~po37  & n10208;
  assign n10216 = ~n10214 & ~n10215;
  assign n10217 = ~n10209 & ~n10216;
  assign n10218 = po38  & ~n10217;
  assign n10219 = ~po38  & ~n10209;
  assign n10220 = ~n10216 & n10219;
  assign n10221 = ~n9767 & po18 ;
  assign n10222 = ~n9773 & n10221;
  assign n10223 = n9772 & ~n10222;
  assign n10224 = n9774 & n10221;
  assign n10225 = ~n10223 & ~n10224;
  assign n10226 = ~n10220 & n10225;
  assign n10227 = ~n10218 & ~n10226;
  assign n10228 = po39  & ~n10227;
  assign n10229 = ~po39  & n10227;
  assign n10230 = ~n9776 & po18 ;
  assign n10231 = ~n9783 & n10230;
  assign n10232 = n9781 & ~n10231;
  assign n10233 = n9784 & n10230;
  assign n10234 = ~n10232 & ~n10233;
  assign n10235 = ~n10229 & n10234;
  assign n10236 = ~n10228 & ~n10235;
  assign n10237 = po40  & ~n10236;
  assign n10238 = ~po40  & ~n10228;
  assign n10239 = ~n10235 & n10238;
  assign n10240 = ~n9786 & po18 ;
  assign n10241 = ~n9792 & n10240;
  assign n10242 = n9791 & ~n10241;
  assign n10243 = n9793 & n10240;
  assign n10244 = ~n10242 & ~n10243;
  assign n10245 = ~n10239 & n10244;
  assign n10246 = ~n10237 & ~n10245;
  assign n10247 = po41  & ~n10246;
  assign n10248 = ~n9795 & ~n9797;
  assign n10249 = po18  & n10248;
  assign n10250 = n9802 & ~n10249;
  assign n10251 = ~n9802 & n10249;
  assign n10252 = ~n10250 & ~n10251;
  assign n10253 = ~po41  & n10246;
  assign n10254 = ~n10252 & ~n10253;
  assign n10255 = ~n10247 & ~n10254;
  assign n10256 = po42  & ~n10255;
  assign n10257 = ~po42  & ~n10247;
  assign n10258 = ~n10254 & n10257;
  assign n10259 = ~n9805 & po18 ;
  assign n10260 = ~n9811 & n10259;
  assign n10261 = n9810 & ~n10260;
  assign n10262 = n9812 & n10259;
  assign n10263 = ~n10261 & ~n10262;
  assign n10264 = ~n10258 & n10263;
  assign n10265 = ~n10256 & ~n10264;
  assign n10266 = po43  & ~n10265;
  assign n10267 = ~po43  & n10265;
  assign n10268 = ~n9814 & po18 ;
  assign n10269 = ~n9821 & n10268;
  assign n10270 = n9819 & ~n10269;
  assign n10271 = n9822 & n10268;
  assign n10272 = ~n10270 & ~n10271;
  assign n10273 = ~n10267 & n10272;
  assign n10274 = ~n10266 & ~n10273;
  assign n10275 = po44  & ~n10274;
  assign n10276 = ~n9824 & ~n9831;
  assign n10277 = po18  & n10276;
  assign n10278 = n9829 & ~n10277;
  assign n10279 = ~n9829 & n10277;
  assign n10280 = ~n10278 & ~n10279;
  assign n10281 = ~po44  & ~n10266;
  assign n10282 = ~n10273 & n10281;
  assign n10283 = ~n10280 & ~n10282;
  assign n10284 = ~n10275 & ~n10283;
  assign n10285 = ~po45  & n10284;
  assign n10286 = ~n10034 & ~n10285;
  assign n10287 = po45  & ~n10284;
  assign n10288 = ~po46  & ~n10287;
  assign n10289 = ~n10286 & n10288;
  assign n10290 = ~n10286 & ~n10287;
  assign n10291 = po46  & ~n10290;
  assign n10292 = n10029 & ~n10289;
  assign n10293 = ~n10291 & ~n10292;
  assign n10294 = po47  & ~n10293;
  assign n10295 = ~n9847 & ~n9849;
  assign n10296 = po18  & n10295;
  assign n10297 = n9854 & ~n10296;
  assign n10298 = ~n9854 & n10296;
  assign n10299 = ~n10297 & ~n10298;
  assign n10300 = ~po47  & n10293;
  assign n10301 = ~n10299 & ~n10300;
  assign n10302 = ~n10294 & ~n10301;
  assign n10303 = po48  & ~n10302;
  assign n10304 = ~po48  & ~n10294;
  assign n10305 = ~n10301 & n10304;
  assign n10306 = ~n9857 & po18 ;
  assign n10307 = ~n9863 & n10306;
  assign n10308 = n9862 & ~n10307;
  assign n10309 = n9864 & n10306;
  assign n10310 = ~n10308 & ~n10309;
  assign n10311 = ~n10305 & n10310;
  assign n10312 = ~n10303 & ~n10311;
  assign n10313 = po49  & ~n10312;
  assign n10314 = ~n9866 & ~n9868;
  assign n10315 = po18  & n10314;
  assign n10316 = n9873 & ~n10315;
  assign n10317 = ~n9873 & n10315;
  assign n10318 = ~n10316 & ~n10317;
  assign n10319 = ~po49  & n10312;
  assign n10320 = ~n10318 & ~n10319;
  assign n10321 = ~n10313 & ~n10320;
  assign n10322 = po50  & ~n10321;
  assign n10323 = ~po50  & ~n10313;
  assign n10324 = ~n10320 & n10323;
  assign n10325 = ~n9876 & po18 ;
  assign n10326 = ~n9882 & n10325;
  assign n10327 = n9881 & ~n10326;
  assign n10328 = n9883 & n10325;
  assign n10329 = ~n10327 & ~n10328;
  assign n10330 = ~n10324 & n10329;
  assign n10331 = ~n10322 & ~n10330;
  assign n10332 = po51  & ~n10331;
  assign n10333 = ~po51  & n10331;
  assign n10334 = ~n9885 & po18 ;
  assign n10335 = ~n9892 & n10334;
  assign n10336 = n9890 & ~n10335;
  assign n10337 = n9893 & n10334;
  assign n10338 = ~n10336 & ~n10337;
  assign n10339 = ~n10333 & n10338;
  assign n10340 = ~n10332 & ~n10339;
  assign n10341 = po52  & ~n10340;
  assign n10342 = ~po52  & ~n10332;
  assign n10343 = ~n10339 & n10342;
  assign n10344 = ~n9895 & po18 ;
  assign n10345 = ~n9901 & n10344;
  assign n10346 = n9900 & ~n10345;
  assign n10347 = n9902 & n10344;
  assign n10348 = ~n10346 & ~n10347;
  assign n10349 = ~n10343 & n10348;
  assign n10350 = ~n10341 & ~n10349;
  assign n10351 = po53  & ~n10350;
  assign n10352 = ~n9904 & ~n9906;
  assign n10353 = po18  & n10352;
  assign n10354 = n9911 & ~n10353;
  assign n10355 = ~n9911 & n10353;
  assign n10356 = ~n10354 & ~n10355;
  assign n10357 = ~po53  & n10350;
  assign n10358 = ~n10356 & ~n10357;
  assign n10359 = ~n10351 & ~n10358;
  assign n10360 = po54  & ~n10359;
  assign n10361 = ~po54  & ~n10351;
  assign n10362 = ~n10358 & n10361;
  assign n10363 = ~n9914 & po18 ;
  assign n10364 = ~n9920 & n10363;
  assign n10365 = n9919 & ~n10364;
  assign n10366 = n9921 & n10363;
  assign n10367 = ~n10365 & ~n10366;
  assign n10368 = ~n10362 & n10367;
  assign n10369 = ~n10360 & ~n10368;
  assign n10370 = po55  & ~n10369;
  assign n10371 = ~po55  & n10369;
  assign n10372 = ~n9923 & po18 ;
  assign n10373 = ~n9930 & n10372;
  assign n10374 = n9928 & ~n10373;
  assign n10375 = n9931 & n10372;
  assign n10376 = ~n10374 & ~n10375;
  assign n10377 = ~n10371 & n10376;
  assign n10378 = ~n10370 & ~n10377;
  assign n10379 = po56  & ~n10378;
  assign n10380 = ~po56  & ~n10370;
  assign n10381 = ~n10377 & n10380;
  assign n10382 = ~n9933 & po18 ;
  assign n10383 = ~n9939 & n10382;
  assign n10384 = n9938 & ~n10383;
  assign n10385 = n9940 & n10382;
  assign n10386 = ~n10384 & ~n10385;
  assign n10387 = ~n10381 & n10386;
  assign n10388 = ~n10379 & ~n10387;
  assign n10389 = po57  & ~n10388;
  assign n10390 = ~n9942 & ~n9944;
  assign n10391 = po18  & n10390;
  assign n10392 = n9949 & ~n10391;
  assign n10393 = ~n9949 & n10391;
  assign n10394 = ~n10392 & ~n10393;
  assign n10395 = ~po57  & n10388;
  assign n10396 = ~n10394 & ~n10395;
  assign n10397 = ~n10389 & ~n10396;
  assign n10398 = po58  & ~n10397;
  assign n10399 = ~po58  & ~n10389;
  assign n10400 = ~n10396 & n10399;
  assign n10401 = ~n9952 & po18 ;
  assign n10402 = ~n9958 & n10401;
  assign n10403 = n9957 & ~n10402;
  assign n10404 = n9959 & n10401;
  assign n10405 = ~n10403 & ~n10404;
  assign n10406 = ~n10400 & n10405;
  assign n10407 = ~n10398 & ~n10406;
  assign n10408 = po59  & ~n10407;
  assign n10409 = ~po59  & n10407;
  assign n10410 = ~n9961 & po18 ;
  assign n10411 = ~n9968 & n10410;
  assign n10412 = n9966 & ~n10411;
  assign n10413 = n9969 & n10410;
  assign n10414 = ~n10412 & ~n10413;
  assign n10415 = ~n10409 & n10414;
  assign n10416 = ~n10408 & ~n10415;
  assign n10417 = po60  & ~n10416;
  assign n10418 = ~po60  & ~n10408;
  assign n10419 = ~n10415 & n10418;
  assign n10420 = ~n9971 & po18 ;
  assign n10421 = ~n9977 & n10420;
  assign n10422 = n9976 & ~n10421;
  assign n10423 = n9978 & n10420;
  assign n10424 = ~n10422 & ~n10423;
  assign n10425 = ~n10419 & n10424;
  assign n10426 = ~n10417 & ~n10425;
  assign n10427 = po61  & ~n10426;
  assign n10428 = ~n9980 & ~n9982;
  assign n10429 = po18  & n10428;
  assign n10430 = n9987 & ~n10429;
  assign n10431 = ~n9987 & n10429;
  assign n10432 = ~n10430 & ~n10431;
  assign n10433 = ~po61  & n10426;
  assign n10434 = ~n10432 & ~n10433;
  assign n10435 = ~n10427 & ~n10434;
  assign n10436 = po62  & ~n10435;
  assign n10437 = ~po62  & ~n10427;
  assign n10438 = ~n10434 & n10437;
  assign n10439 = ~n9990 & po18 ;
  assign n10440 = ~n9996 & n10439;
  assign n10441 = n9995 & ~n10440;
  assign n10442 = n9997 & n10439;
  assign n10443 = ~n10441 & ~n10442;
  assign n10444 = ~n10438 & n10443;
  assign n10445 = ~n10436 & ~n10444;
  assign n10446 = n10008 & po18 ;
  assign n10447 = ~n10013 & ~n10446;
  assign n10448 = ~n10021 & ~n10447;
  assign n10449 = po18  & ~n10448;
  assign n10450 = ~n9999 & po18 ;
  assign n10451 = ~n10006 & n10450;
  assign n10452 = n10004 & ~n10451;
  assign n10453 = n10007 & n10450;
  assign n10454 = ~n10452 & ~n10453;
  assign n10455 = ~n10449 & n10454;
  assign n10456 = ~n10445 & n10455;
  assign n10457 = ~po63  & ~n10456;
  assign n10458 = n10445 & ~n10454;
  assign n10459 = po63  & n10448;
  assign n10460 = ~n10458 & ~n10459;
  assign po17  = n10457 | ~n10460;
  assign n10462 = ~n10289 & ~n10291;
  assign n10463 = po17  & n10462;
  assign n10464 = n10029 & ~n10463;
  assign n10465 = ~n10029 & n10463;
  assign n10466 = ~n10464 & ~n10465;
  assign n10467 = pi34  & po17 ;
  assign n10468 = ~pi32  & ~pi33 ;
  assign n10469 = ~pi34  & n10468;
  assign n10470 = ~n10467 & ~n10469;
  assign n10471 = po18  & ~n10470;
  assign n10472 = ~po18  & n10470;
  assign n10473 = ~pi34  & po17 ;
  assign n10474 = pi35  & ~n10473;
  assign n10475 = ~pi35  & n10473;
  assign n10476 = ~n10474 & ~n10475;
  assign n10477 = ~n10472 & n10476;
  assign n10478 = ~n10471 & ~n10477;
  assign n10479 = po19  & ~n10478;
  assign n10480 = po18  & ~po17 ;
  assign n10481 = ~n10475 & ~n10480;
  assign n10482 = pi36  & ~n10481;
  assign n10483 = ~pi36  & n10481;
  assign n10484 = ~n10482 & ~n10483;
  assign n10485 = ~po19  & n10478;
  assign n10486 = ~n10484 & ~n10485;
  assign n10487 = ~n10479 & ~n10486;
  assign n10488 = po20  & ~n10487;
  assign n10489 = ~po20  & ~n10479;
  assign n10490 = ~n10486 & n10489;
  assign n10491 = ~n10039 & ~n10044;
  assign n10492 = po17  & n10491;
  assign n10493 = n10043 & ~n10492;
  assign n10494 = ~n10043 & n10492;
  assign n10495 = ~n10493 & ~n10494;
  assign n10496 = ~n10490 & ~n10495;
  assign n10497 = ~n10488 & ~n10496;
  assign n10498 = po21  & ~n10497;
  assign n10499 = ~n10047 & ~n10049;
  assign n10500 = po17  & n10499;
  assign n10501 = ~n10054 & ~n10500;
  assign n10502 = n10054 & n10500;
  assign n10503 = ~n10501 & ~n10502;
  assign n10504 = ~po21  & n10497;
  assign n10505 = ~n10503 & ~n10504;
  assign n10506 = ~n10498 & ~n10505;
  assign n10507 = po22  & ~n10506;
  assign n10508 = ~po22  & ~n10498;
  assign n10509 = ~n10505 & n10508;
  assign n10510 = ~n10057 & ~n10058;
  assign n10511 = po17  & n10510;
  assign n10512 = n10063 & ~n10511;
  assign n10513 = ~n10063 & n10511;
  assign n10514 = ~n10512 & ~n10513;
  assign n10515 = ~n10509 & n10514;
  assign n10516 = ~n10507 & ~n10515;
  assign n10517 = po23  & ~n10516;
  assign n10518 = ~n10066 & ~n10068;
  assign n10519 = po17  & n10518;
  assign n10520 = n10073 & ~n10519;
  assign n10521 = ~n10073 & n10519;
  assign n10522 = ~n10520 & ~n10521;
  assign n10523 = ~po23  & n10516;
  assign n10524 = ~n10522 & ~n10523;
  assign n10525 = ~n10517 & ~n10524;
  assign n10526 = po24  & ~n10525;
  assign n10527 = ~po24  & ~n10517;
  assign n10528 = ~n10524 & n10527;
  assign n10529 = ~n10076 & ~n10077;
  assign n10530 = po17  & n10529;
  assign n10531 = n10082 & n10530;
  assign n10532 = ~n10082 & ~n10530;
  assign n10533 = ~n10531 & ~n10532;
  assign n10534 = ~n10528 & n10533;
  assign n10535 = ~n10526 & ~n10534;
  assign n10536 = po25  & ~n10535;
  assign n10537 = ~n10085 & ~n10087;
  assign n10538 = po17  & n10537;
  assign n10539 = n10092 & ~n10538;
  assign n10540 = ~n10092 & n10538;
  assign n10541 = ~n10539 & ~n10540;
  assign n10542 = ~po25  & n10535;
  assign n10543 = ~n10541 & ~n10542;
  assign n10544 = ~n10536 & ~n10543;
  assign n10545 = po26  & ~n10544;
  assign n10546 = ~po26  & ~n10536;
  assign n10547 = ~n10543 & n10546;
  assign n10548 = ~n10095 & ~n10096;
  assign n10549 = po17  & n10548;
  assign n10550 = ~n10101 & ~n10549;
  assign n10551 = n10101 & n10549;
  assign n10552 = ~n10550 & ~n10551;
  assign n10553 = ~n10547 & n10552;
  assign n10554 = ~n10545 & ~n10553;
  assign n10555 = po27  & ~n10554;
  assign n10556 = ~n10104 & ~n10106;
  assign n10557 = po17  & n10556;
  assign n10558 = n10111 & ~n10557;
  assign n10559 = ~n10111 & n10557;
  assign n10560 = ~n10558 & ~n10559;
  assign n10561 = ~po27  & n10554;
  assign n10562 = ~n10560 & ~n10561;
  assign n10563 = ~n10555 & ~n10562;
  assign n10564 = po28  & ~n10563;
  assign n10565 = ~n10114 & ~n10115;
  assign n10566 = po17  & n10565;
  assign n10567 = n10120 & ~n10566;
  assign n10568 = ~n10120 & n10566;
  assign n10569 = ~n10567 & ~n10568;
  assign n10570 = ~po28  & ~n10555;
  assign n10571 = ~n10562 & n10570;
  assign n10572 = ~n10569 & ~n10571;
  assign n10573 = ~n10564 & ~n10572;
  assign n10574 = po29  & ~n10573;
  assign n10575 = ~n10123 & ~n10125;
  assign n10576 = po17  & n10575;
  assign n10577 = n10130 & ~n10576;
  assign n10578 = ~n10130 & n10576;
  assign n10579 = ~n10577 & ~n10578;
  assign n10580 = ~po29  & n10573;
  assign n10581 = ~n10579 & ~n10580;
  assign n10582 = ~n10574 & ~n10581;
  assign n10583 = po30  & ~n10582;
  assign n10584 = ~po30  & ~n10574;
  assign n10585 = ~n10581 & n10584;
  assign n10586 = ~n10133 & po17 ;
  assign n10587 = ~n10139 & n10586;
  assign n10588 = n10138 & ~n10587;
  assign n10589 = n10140 & n10586;
  assign n10590 = ~n10588 & ~n10589;
  assign n10591 = ~n10585 & n10590;
  assign n10592 = ~n10583 & ~n10591;
  assign n10593 = po31  & ~n10592;
  assign n10594 = ~n10142 & ~n10144;
  assign n10595 = po17  & n10594;
  assign n10596 = n10149 & ~n10595;
  assign n10597 = ~n10149 & n10595;
  assign n10598 = ~n10596 & ~n10597;
  assign n10599 = ~po31  & n10592;
  assign n10600 = ~n10598 & ~n10599;
  assign n10601 = ~n10593 & ~n10600;
  assign n10602 = po32  & ~n10601;
  assign n10603 = ~n10152 & ~n10153;
  assign n10604 = po17  & n10603;
  assign n10605 = n10158 & ~n10604;
  assign n10606 = ~n10158 & n10604;
  assign n10607 = ~n10605 & ~n10606;
  assign n10608 = ~po32  & ~n10593;
  assign n10609 = ~n10600 & n10608;
  assign n10610 = ~n10607 & ~n10609;
  assign n10611 = ~n10602 & ~n10610;
  assign n10612 = po33  & ~n10611;
  assign n10613 = ~n10161 & ~n10163;
  assign n10614 = po17  & n10613;
  assign n10615 = n10168 & ~n10614;
  assign n10616 = ~n10168 & n10614;
  assign n10617 = ~n10615 & ~n10616;
  assign n10618 = ~po33  & n10611;
  assign n10619 = ~n10617 & ~n10618;
  assign n10620 = ~n10612 & ~n10619;
  assign n10621 = po34  & ~n10620;
  assign n10622 = ~po34  & ~n10612;
  assign n10623 = ~n10619 & n10622;
  assign n10624 = ~n10171 & po17 ;
  assign n10625 = ~n10177 & n10624;
  assign n10626 = n10176 & ~n10625;
  assign n10627 = n10178 & n10624;
  assign n10628 = ~n10626 & ~n10627;
  assign n10629 = ~n10623 & n10628;
  assign n10630 = ~n10621 & ~n10629;
  assign n10631 = po35  & ~n10630;
  assign n10632 = ~n10180 & ~n10182;
  assign n10633 = po17  & n10632;
  assign n10634 = n10187 & ~n10633;
  assign n10635 = ~n10187 & n10633;
  assign n10636 = ~n10634 & ~n10635;
  assign n10637 = ~po35  & n10630;
  assign n10638 = ~n10636 & ~n10637;
  assign n10639 = ~n10631 & ~n10638;
  assign n10640 = po36  & ~n10639;
  assign n10641 = ~n10190 & ~n10191;
  assign n10642 = po17  & n10641;
  assign n10643 = n10196 & ~n10642;
  assign n10644 = ~n10196 & n10642;
  assign n10645 = ~n10643 & ~n10644;
  assign n10646 = ~po36  & ~n10631;
  assign n10647 = ~n10638 & n10646;
  assign n10648 = ~n10645 & ~n10647;
  assign n10649 = ~n10640 & ~n10648;
  assign n10650 = po37  & ~n10649;
  assign n10651 = ~n10199 & ~n10201;
  assign n10652 = po17  & n10651;
  assign n10653 = n10206 & ~n10652;
  assign n10654 = ~n10206 & n10652;
  assign n10655 = ~n10653 & ~n10654;
  assign n10656 = ~po37  & n10649;
  assign n10657 = ~n10655 & ~n10656;
  assign n10658 = ~n10650 & ~n10657;
  assign n10659 = po38  & ~n10658;
  assign n10660 = ~po38  & ~n10650;
  assign n10661 = ~n10657 & n10660;
  assign n10662 = ~n10209 & po17 ;
  assign n10663 = ~n10215 & n10662;
  assign n10664 = n10214 & ~n10663;
  assign n10665 = n10216 & n10662;
  assign n10666 = ~n10664 & ~n10665;
  assign n10667 = ~n10661 & n10666;
  assign n10668 = ~n10659 & ~n10667;
  assign n10669 = po39  & ~n10668;
  assign n10670 = ~n10218 & ~n10220;
  assign n10671 = po17  & n10670;
  assign n10672 = n10225 & ~n10671;
  assign n10673 = ~n10225 & n10671;
  assign n10674 = ~n10672 & ~n10673;
  assign n10675 = ~po39  & n10668;
  assign n10676 = ~n10674 & ~n10675;
  assign n10677 = ~n10669 & ~n10676;
  assign n10678 = po40  & ~n10677;
  assign n10679 = ~n10228 & ~n10229;
  assign n10680 = po17  & n10679;
  assign n10681 = n10234 & ~n10680;
  assign n10682 = ~n10234 & n10680;
  assign n10683 = ~n10681 & ~n10682;
  assign n10684 = ~po40  & ~n10669;
  assign n10685 = ~n10676 & n10684;
  assign n10686 = ~n10683 & ~n10685;
  assign n10687 = ~n10678 & ~n10686;
  assign n10688 = po41  & ~n10687;
  assign n10689 = ~n10237 & ~n10239;
  assign n10690 = po17  & n10689;
  assign n10691 = n10244 & ~n10690;
  assign n10692 = ~n10244 & n10690;
  assign n10693 = ~n10691 & ~n10692;
  assign n10694 = ~po41  & n10687;
  assign n10695 = ~n10693 & ~n10694;
  assign n10696 = ~n10688 & ~n10695;
  assign n10697 = po42  & ~n10696;
  assign n10698 = ~po42  & ~n10688;
  assign n10699 = ~n10695 & n10698;
  assign n10700 = ~n10247 & po17 ;
  assign n10701 = ~n10253 & n10700;
  assign n10702 = n10252 & ~n10701;
  assign n10703 = n10254 & n10700;
  assign n10704 = ~n10702 & ~n10703;
  assign n10705 = ~n10699 & n10704;
  assign n10706 = ~n10697 & ~n10705;
  assign n10707 = po43  & ~n10706;
  assign n10708 = ~n10256 & ~n10258;
  assign n10709 = po17  & n10708;
  assign n10710 = n10263 & ~n10709;
  assign n10711 = ~n10263 & n10709;
  assign n10712 = ~n10710 & ~n10711;
  assign n10713 = ~po43  & n10706;
  assign n10714 = ~n10712 & ~n10713;
  assign n10715 = ~n10707 & ~n10714;
  assign n10716 = po44  & ~n10715;
  assign n10717 = ~n10266 & ~n10267;
  assign n10718 = po17  & n10717;
  assign n10719 = n10272 & ~n10718;
  assign n10720 = ~n10272 & n10718;
  assign n10721 = ~n10719 & ~n10720;
  assign n10722 = ~po44  & ~n10707;
  assign n10723 = ~n10714 & n10722;
  assign n10724 = ~n10721 & ~n10723;
  assign n10725 = ~n10716 & ~n10724;
  assign n10726 = ~po45  & n10725;
  assign n10727 = ~n10275 & po17 ;
  assign n10728 = ~n10282 & n10727;
  assign n10729 = n10280 & ~n10728;
  assign n10730 = n10283 & n10727;
  assign n10731 = ~n10729 & ~n10730;
  assign n10732 = ~n10726 & n10731;
  assign n10733 = po45  & ~n10725;
  assign n10734 = ~n10732 & ~n10733;
  assign n10735 = po46  & ~n10734;
  assign n10736 = ~n10285 & ~n10287;
  assign n10737 = po17  & n10736;
  assign n10738 = n10034 & ~n10737;
  assign n10739 = ~n10034 & n10737;
  assign n10740 = ~n10738 & ~n10739;
  assign n10741 = ~po46  & ~n10733;
  assign n10742 = ~n10732 & n10741;
  assign n10743 = n10740 & ~n10742;
  assign n10744 = ~n10735 & ~n10743;
  assign n10745 = ~po47  & n10744;
  assign n10746 = po47  & ~n10744;
  assign n10747 = ~n10466 & ~n10745;
  assign n10748 = ~n10746 & ~n10747;
  assign n10749 = po48  & ~n10748;
  assign n10750 = ~po48  & ~n10746;
  assign n10751 = ~n10747 & n10750;
  assign n10752 = ~n10294 & po17 ;
  assign n10753 = ~n10300 & n10752;
  assign n10754 = n10299 & ~n10753;
  assign n10755 = n10301 & n10752;
  assign n10756 = ~n10754 & ~n10755;
  assign n10757 = ~n10751 & n10756;
  assign n10758 = ~n10749 & ~n10757;
  assign n10759 = po49  & ~n10758;
  assign n10760 = ~n10303 & ~n10305;
  assign n10761 = po17  & n10760;
  assign n10762 = n10310 & ~n10761;
  assign n10763 = ~n10310 & n10761;
  assign n10764 = ~n10762 & ~n10763;
  assign n10765 = ~po49  & n10758;
  assign n10766 = ~n10764 & ~n10765;
  assign n10767 = ~n10759 & ~n10766;
  assign n10768 = po50  & ~n10767;
  assign n10769 = ~po50  & ~n10759;
  assign n10770 = ~n10766 & n10769;
  assign n10771 = ~n10313 & po17 ;
  assign n10772 = ~n10319 & n10771;
  assign n10773 = n10318 & ~n10772;
  assign n10774 = n10320 & n10771;
  assign n10775 = ~n10773 & ~n10774;
  assign n10776 = ~n10770 & n10775;
  assign n10777 = ~n10768 & ~n10776;
  assign n10778 = po51  & ~n10777;
  assign n10779 = ~n10322 & ~n10324;
  assign n10780 = po17  & n10779;
  assign n10781 = n10329 & ~n10780;
  assign n10782 = ~n10329 & n10780;
  assign n10783 = ~n10781 & ~n10782;
  assign n10784 = ~po51  & n10777;
  assign n10785 = ~n10783 & ~n10784;
  assign n10786 = ~n10778 & ~n10785;
  assign n10787 = po52  & ~n10786;
  assign n10788 = ~n10332 & ~n10333;
  assign n10789 = po17  & n10788;
  assign n10790 = n10338 & ~n10789;
  assign n10791 = ~n10338 & n10789;
  assign n10792 = ~n10790 & ~n10791;
  assign n10793 = ~po52  & ~n10778;
  assign n10794 = ~n10785 & n10793;
  assign n10795 = ~n10792 & ~n10794;
  assign n10796 = ~n10787 & ~n10795;
  assign n10797 = po53  & ~n10796;
  assign n10798 = ~n10341 & ~n10343;
  assign n10799 = po17  & n10798;
  assign n10800 = n10348 & ~n10799;
  assign n10801 = ~n10348 & n10799;
  assign n10802 = ~n10800 & ~n10801;
  assign n10803 = ~po53  & n10796;
  assign n10804 = ~n10802 & ~n10803;
  assign n10805 = ~n10797 & ~n10804;
  assign n10806 = po54  & ~n10805;
  assign n10807 = ~po54  & ~n10797;
  assign n10808 = ~n10804 & n10807;
  assign n10809 = ~n10351 & po17 ;
  assign n10810 = ~n10357 & n10809;
  assign n10811 = n10356 & ~n10810;
  assign n10812 = n10358 & n10809;
  assign n10813 = ~n10811 & ~n10812;
  assign n10814 = ~n10808 & n10813;
  assign n10815 = ~n10806 & ~n10814;
  assign n10816 = po55  & ~n10815;
  assign n10817 = ~n10360 & ~n10362;
  assign n10818 = po17  & n10817;
  assign n10819 = n10367 & ~n10818;
  assign n10820 = ~n10367 & n10818;
  assign n10821 = ~n10819 & ~n10820;
  assign n10822 = ~po55  & n10815;
  assign n10823 = ~n10821 & ~n10822;
  assign n10824 = ~n10816 & ~n10823;
  assign n10825 = po56  & ~n10824;
  assign n10826 = ~n10370 & ~n10371;
  assign n10827 = po17  & n10826;
  assign n10828 = n10376 & ~n10827;
  assign n10829 = ~n10376 & n10827;
  assign n10830 = ~n10828 & ~n10829;
  assign n10831 = ~po56  & ~n10816;
  assign n10832 = ~n10823 & n10831;
  assign n10833 = ~n10830 & ~n10832;
  assign n10834 = ~n10825 & ~n10833;
  assign n10835 = po57  & ~n10834;
  assign n10836 = ~n10379 & ~n10381;
  assign n10837 = po17  & n10836;
  assign n10838 = n10386 & ~n10837;
  assign n10839 = ~n10386 & n10837;
  assign n10840 = ~n10838 & ~n10839;
  assign n10841 = ~po57  & n10834;
  assign n10842 = ~n10840 & ~n10841;
  assign n10843 = ~n10835 & ~n10842;
  assign n10844 = po58  & ~n10843;
  assign n10845 = ~po58  & ~n10835;
  assign n10846 = ~n10842 & n10845;
  assign n10847 = ~n10389 & po17 ;
  assign n10848 = ~n10395 & n10847;
  assign n10849 = n10394 & ~n10848;
  assign n10850 = n10396 & n10847;
  assign n10851 = ~n10849 & ~n10850;
  assign n10852 = ~n10846 & n10851;
  assign n10853 = ~n10844 & ~n10852;
  assign n10854 = po59  & ~n10853;
  assign n10855 = ~n10398 & ~n10400;
  assign n10856 = po17  & n10855;
  assign n10857 = n10405 & ~n10856;
  assign n10858 = ~n10405 & n10856;
  assign n10859 = ~n10857 & ~n10858;
  assign n10860 = ~po59  & n10853;
  assign n10861 = ~n10859 & ~n10860;
  assign n10862 = ~n10854 & ~n10861;
  assign n10863 = po60  & ~n10862;
  assign n10864 = ~n10408 & ~n10409;
  assign n10865 = po17  & n10864;
  assign n10866 = n10414 & ~n10865;
  assign n10867 = ~n10414 & n10865;
  assign n10868 = ~n10866 & ~n10867;
  assign n10869 = ~po60  & ~n10854;
  assign n10870 = ~n10861 & n10869;
  assign n10871 = ~n10868 & ~n10870;
  assign n10872 = ~n10863 & ~n10871;
  assign n10873 = po61  & ~n10872;
  assign n10874 = ~n10417 & ~n10419;
  assign n10875 = po17  & n10874;
  assign n10876 = n10424 & ~n10875;
  assign n10877 = ~n10424 & n10875;
  assign n10878 = ~n10876 & ~n10877;
  assign n10879 = ~po61  & n10872;
  assign n10880 = ~n10878 & ~n10879;
  assign n10881 = ~n10873 & ~n10880;
  assign n10882 = po62  & ~n10881;
  assign n10883 = ~po62  & ~n10873;
  assign n10884 = ~n10880 & n10883;
  assign n10885 = ~n10427 & po17 ;
  assign n10886 = ~n10433 & n10885;
  assign n10887 = n10432 & ~n10886;
  assign n10888 = n10434 & n10885;
  assign n10889 = ~n10887 & ~n10888;
  assign n10890 = ~n10884 & n10889;
  assign n10891 = ~n10882 & ~n10890;
  assign n10892 = n10454 & po17 ;
  assign n10893 = ~n10445 & n10892;
  assign n10894 = ~n10436 & ~n10438;
  assign n10895 = po17  & n10894;
  assign n10896 = n10443 & ~n10895;
  assign n10897 = ~n10443 & n10895;
  assign n10898 = ~n10896 & ~n10897;
  assign n10899 = ~n10458 & ~n10893;
  assign n10900 = ~n10898 & n10899;
  assign n10901 = ~n10891 & n10900;
  assign n10902 = ~po63  & ~n10901;
  assign n10903 = n10891 & n10898;
  assign n10904 = n10445 & ~n10892;
  assign n10905 = ~n10445 & n10454;
  assign n10906 = po63  & ~n10905;
  assign n10907 = ~n10904 & n10906;
  assign n10908 = ~n10903 & ~n10907;
  assign po16  = n10902 | ~n10908;
  assign n10910 = ~n10746 & po16 ;
  assign n10911 = ~n10745 & n10910;
  assign n10912 = n10466 & ~n10911;
  assign n10913 = n10747 & n10910;
  assign n10914 = ~n10912 & ~n10913;
  assign n10915 = pi32  & po16 ;
  assign n10916 = ~pi30  & ~pi31 ;
  assign n10917 = ~pi32  & n10916;
  assign n10918 = ~n10915 & ~n10917;
  assign n10919 = po17  & ~n10918;
  assign n10920 = ~pi32  & po16 ;
  assign n10921 = pi33  & ~n10920;
  assign n10922 = ~pi33  & n10920;
  assign n10923 = ~n10921 & ~n10922;
  assign n10924 = ~po17  & n10918;
  assign n10925 = n10923 & ~n10924;
  assign n10926 = ~n10919 & ~n10925;
  assign n10927 = po18  & ~n10926;
  assign n10928 = ~po18  & ~n10919;
  assign n10929 = ~n10925 & n10928;
  assign n10930 = po17  & ~po16 ;
  assign n10931 = ~n10922 & ~n10930;
  assign n10932 = pi34  & ~n10931;
  assign n10933 = ~pi34  & n10931;
  assign n10934 = ~n10932 & ~n10933;
  assign n10935 = ~n10929 & ~n10934;
  assign n10936 = ~n10927 & ~n10935;
  assign n10937 = po19  & ~n10936;
  assign n10938 = ~po19  & n10936;
  assign n10939 = ~n10471 & ~n10472;
  assign n10940 = po16  & n10939;
  assign n10941 = n10476 & ~n10940;
  assign n10942 = ~n10476 & n10940;
  assign n10943 = ~n10941 & ~n10942;
  assign n10944 = ~n10938 & ~n10943;
  assign n10945 = ~n10937 & ~n10944;
  assign n10946 = po20  & ~n10945;
  assign n10947 = ~po20  & ~n10937;
  assign n10948 = ~n10944 & n10947;
  assign n10949 = ~n10479 & po16 ;
  assign n10950 = ~n10485 & n10949;
  assign n10951 = n10484 & ~n10950;
  assign n10952 = n10486 & n10949;
  assign n10953 = ~n10951 & ~n10952;
  assign n10954 = ~n10948 & n10953;
  assign n10955 = ~n10946 & ~n10954;
  assign n10956 = po21  & ~n10955;
  assign n10957 = ~po21  & n10955;
  assign n10958 = ~n10488 & ~n10490;
  assign n10959 = po16  & n10958;
  assign n10960 = n10495 & ~n10959;
  assign n10961 = ~n10495 & n10959;
  assign n10962 = ~n10960 & ~n10961;
  assign n10963 = ~n10957 & n10962;
  assign n10964 = ~n10956 & ~n10963;
  assign n10965 = po22  & ~n10964;
  assign n10966 = ~po22  & ~n10956;
  assign n10967 = ~n10963 & n10966;
  assign n10968 = ~n10498 & po16 ;
  assign n10969 = ~n10504 & n10968;
  assign n10970 = n10503 & ~n10969;
  assign n10971 = n10505 & n10968;
  assign n10972 = ~n10970 & ~n10971;
  assign n10973 = ~n10967 & n10972;
  assign n10974 = ~n10965 & ~n10973;
  assign n10975 = po23  & ~n10974;
  assign n10976 = ~po23  & n10974;
  assign n10977 = ~n10507 & ~n10509;
  assign n10978 = po16  & n10977;
  assign n10979 = n10514 & n10978;
  assign n10980 = ~n10514 & ~n10978;
  assign n10981 = ~n10979 & ~n10980;
  assign n10982 = ~n10976 & n10981;
  assign n10983 = ~n10975 & ~n10982;
  assign n10984 = po24  & ~n10983;
  assign n10985 = ~po24  & ~n10975;
  assign n10986 = ~n10982 & n10985;
  assign n10987 = ~n10517 & po16 ;
  assign n10988 = ~n10523 & n10987;
  assign n10989 = n10522 & ~n10988;
  assign n10990 = n10524 & n10987;
  assign n10991 = ~n10989 & ~n10990;
  assign n10992 = ~n10986 & n10991;
  assign n10993 = ~n10984 & ~n10992;
  assign n10994 = po25  & ~n10993;
  assign n10995 = ~po25  & n10993;
  assign n10996 = ~n10526 & ~n10528;
  assign n10997 = po16  & n10996;
  assign n10998 = ~n10533 & ~n10997;
  assign n10999 = n10533 & n10997;
  assign n11000 = ~n10998 & ~n10999;
  assign n11001 = ~n10995 & n11000;
  assign n11002 = ~n10994 & ~n11001;
  assign n11003 = po26  & ~n11002;
  assign n11004 = ~po26  & ~n10994;
  assign n11005 = ~n11001 & n11004;
  assign n11006 = ~n10536 & po16 ;
  assign n11007 = ~n10542 & n11006;
  assign n11008 = n10541 & ~n11007;
  assign n11009 = n10543 & n11006;
  assign n11010 = ~n11008 & ~n11009;
  assign n11011 = ~n11005 & n11010;
  assign n11012 = ~n11003 & ~n11011;
  assign n11013 = po27  & ~n11012;
  assign n11014 = ~n10545 & ~n10547;
  assign n11015 = po16  & n11014;
  assign n11016 = n10552 & ~n11015;
  assign n11017 = ~n10552 & n11015;
  assign n11018 = ~n11016 & ~n11017;
  assign n11019 = ~po27  & n11012;
  assign n11020 = ~n11018 & ~n11019;
  assign n11021 = ~n11013 & ~n11020;
  assign n11022 = po28  & ~n11021;
  assign n11023 = ~po28  & ~n11013;
  assign n11024 = ~n11020 & n11023;
  assign n11025 = ~n10555 & po16 ;
  assign n11026 = ~n10561 & n11025;
  assign n11027 = n10560 & ~n11026;
  assign n11028 = n10562 & n11025;
  assign n11029 = ~n11027 & ~n11028;
  assign n11030 = ~n11024 & n11029;
  assign n11031 = ~n11022 & ~n11030;
  assign n11032 = po29  & ~n11031;
  assign n11033 = ~po29  & n11031;
  assign n11034 = ~n10564 & po16 ;
  assign n11035 = ~n10571 & n11034;
  assign n11036 = n10569 & ~n11035;
  assign n11037 = n10572 & n11034;
  assign n11038 = ~n11036 & ~n11037;
  assign n11039 = ~n11033 & n11038;
  assign n11040 = ~n11032 & ~n11039;
  assign n11041 = po30  & ~n11040;
  assign n11042 = ~po30  & ~n11032;
  assign n11043 = ~n11039 & n11042;
  assign n11044 = ~n10574 & po16 ;
  assign n11045 = ~n10580 & n11044;
  assign n11046 = n10579 & ~n11045;
  assign n11047 = n10581 & n11044;
  assign n11048 = ~n11046 & ~n11047;
  assign n11049 = ~n11043 & n11048;
  assign n11050 = ~n11041 & ~n11049;
  assign n11051 = po31  & ~n11050;
  assign n11052 = ~n10583 & ~n10585;
  assign n11053 = po16  & n11052;
  assign n11054 = n10590 & ~n11053;
  assign n11055 = ~n10590 & n11053;
  assign n11056 = ~n11054 & ~n11055;
  assign n11057 = ~po31  & n11050;
  assign n11058 = ~n11056 & ~n11057;
  assign n11059 = ~n11051 & ~n11058;
  assign n11060 = po32  & ~n11059;
  assign n11061 = ~po32  & ~n11051;
  assign n11062 = ~n11058 & n11061;
  assign n11063 = ~n10593 & po16 ;
  assign n11064 = ~n10599 & n11063;
  assign n11065 = n10598 & ~n11064;
  assign n11066 = n10600 & n11063;
  assign n11067 = ~n11065 & ~n11066;
  assign n11068 = ~n11062 & n11067;
  assign n11069 = ~n11060 & ~n11068;
  assign n11070 = po33  & ~n11069;
  assign n11071 = ~po33  & n11069;
  assign n11072 = ~n10602 & po16 ;
  assign n11073 = ~n10609 & n11072;
  assign n11074 = n10607 & ~n11073;
  assign n11075 = n10610 & n11072;
  assign n11076 = ~n11074 & ~n11075;
  assign n11077 = ~n11071 & n11076;
  assign n11078 = ~n11070 & ~n11077;
  assign n11079 = po34  & ~n11078;
  assign n11080 = ~po34  & ~n11070;
  assign n11081 = ~n11077 & n11080;
  assign n11082 = ~n10612 & po16 ;
  assign n11083 = ~n10618 & n11082;
  assign n11084 = n10617 & ~n11083;
  assign n11085 = n10619 & n11082;
  assign n11086 = ~n11084 & ~n11085;
  assign n11087 = ~n11081 & n11086;
  assign n11088 = ~n11079 & ~n11087;
  assign n11089 = po35  & ~n11088;
  assign n11090 = ~n10621 & ~n10623;
  assign n11091 = po16  & n11090;
  assign n11092 = n10628 & ~n11091;
  assign n11093 = ~n10628 & n11091;
  assign n11094 = ~n11092 & ~n11093;
  assign n11095 = ~po35  & n11088;
  assign n11096 = ~n11094 & ~n11095;
  assign n11097 = ~n11089 & ~n11096;
  assign n11098 = po36  & ~n11097;
  assign n11099 = ~po36  & ~n11089;
  assign n11100 = ~n11096 & n11099;
  assign n11101 = ~n10631 & po16 ;
  assign n11102 = ~n10637 & n11101;
  assign n11103 = n10636 & ~n11102;
  assign n11104 = n10638 & n11101;
  assign n11105 = ~n11103 & ~n11104;
  assign n11106 = ~n11100 & n11105;
  assign n11107 = ~n11098 & ~n11106;
  assign n11108 = po37  & ~n11107;
  assign n11109 = ~po37  & n11107;
  assign n11110 = ~n10640 & po16 ;
  assign n11111 = ~n10647 & n11110;
  assign n11112 = n10645 & ~n11111;
  assign n11113 = n10648 & n11110;
  assign n11114 = ~n11112 & ~n11113;
  assign n11115 = ~n11109 & n11114;
  assign n11116 = ~n11108 & ~n11115;
  assign n11117 = po38  & ~n11116;
  assign n11118 = ~po38  & ~n11108;
  assign n11119 = ~n11115 & n11118;
  assign n11120 = ~n10650 & po16 ;
  assign n11121 = ~n10656 & n11120;
  assign n11122 = n10655 & ~n11121;
  assign n11123 = n10657 & n11120;
  assign n11124 = ~n11122 & ~n11123;
  assign n11125 = ~n11119 & n11124;
  assign n11126 = ~n11117 & ~n11125;
  assign n11127 = po39  & ~n11126;
  assign n11128 = ~n10659 & ~n10661;
  assign n11129 = po16  & n11128;
  assign n11130 = n10666 & ~n11129;
  assign n11131 = ~n10666 & n11129;
  assign n11132 = ~n11130 & ~n11131;
  assign n11133 = ~po39  & n11126;
  assign n11134 = ~n11132 & ~n11133;
  assign n11135 = ~n11127 & ~n11134;
  assign n11136 = po40  & ~n11135;
  assign n11137 = ~po40  & ~n11127;
  assign n11138 = ~n11134 & n11137;
  assign n11139 = ~n10669 & po16 ;
  assign n11140 = ~n10675 & n11139;
  assign n11141 = n10674 & ~n11140;
  assign n11142 = n10676 & n11139;
  assign n11143 = ~n11141 & ~n11142;
  assign n11144 = ~n11138 & n11143;
  assign n11145 = ~n11136 & ~n11144;
  assign n11146 = po41  & ~n11145;
  assign n11147 = ~po41  & n11145;
  assign n11148 = ~n10678 & po16 ;
  assign n11149 = ~n10685 & n11148;
  assign n11150 = n10683 & ~n11149;
  assign n11151 = n10686 & n11148;
  assign n11152 = ~n11150 & ~n11151;
  assign n11153 = ~n11147 & n11152;
  assign n11154 = ~n11146 & ~n11153;
  assign n11155 = po42  & ~n11154;
  assign n11156 = ~po42  & ~n11146;
  assign n11157 = ~n11153 & n11156;
  assign n11158 = ~n10688 & po16 ;
  assign n11159 = ~n10694 & n11158;
  assign n11160 = n10693 & ~n11159;
  assign n11161 = n10695 & n11158;
  assign n11162 = ~n11160 & ~n11161;
  assign n11163 = ~n11157 & n11162;
  assign n11164 = ~n11155 & ~n11163;
  assign n11165 = po43  & ~n11164;
  assign n11166 = ~n10697 & ~n10699;
  assign n11167 = po16  & n11166;
  assign n11168 = n10704 & ~n11167;
  assign n11169 = ~n10704 & n11167;
  assign n11170 = ~n11168 & ~n11169;
  assign n11171 = ~po43  & n11164;
  assign n11172 = ~n11170 & ~n11171;
  assign n11173 = ~n11165 & ~n11172;
  assign n11174 = po44  & ~n11173;
  assign n11175 = ~po44  & ~n11165;
  assign n11176 = ~n11172 & n11175;
  assign n11177 = ~n10707 & po16 ;
  assign n11178 = ~n10713 & n11177;
  assign n11179 = n10712 & ~n11178;
  assign n11180 = n10714 & n11177;
  assign n11181 = ~n11179 & ~n11180;
  assign n11182 = ~n11176 & n11181;
  assign n11183 = ~n11174 & ~n11182;
  assign n11184 = po45  & ~n11183;
  assign n11185 = ~po45  & n11183;
  assign n11186 = ~n10716 & po16 ;
  assign n11187 = ~n10723 & n11186;
  assign n11188 = n10721 & ~n11187;
  assign n11189 = n10724 & n11186;
  assign n11190 = ~n11188 & ~n11189;
  assign n11191 = ~n11185 & n11190;
  assign n11192 = ~n11184 & ~n11191;
  assign n11193 = po46  & ~n11192;
  assign n11194 = ~n10726 & ~n10733;
  assign n11195 = po16  & n11194;
  assign n11196 = n10731 & ~n11195;
  assign n11197 = ~n10731 & n11195;
  assign n11198 = ~n11196 & ~n11197;
  assign n11199 = ~po46  & ~n11184;
  assign n11200 = ~n11191 & n11199;
  assign n11201 = ~n11198 & ~n11200;
  assign n11202 = ~n11193 & ~n11201;
  assign n11203 = ~po47  & n11202;
  assign n11204 = ~n10735 & ~n10742;
  assign n11205 = po16  & n11204;
  assign n11206 = n10740 & n11205;
  assign n11207 = ~n10740 & ~n11205;
  assign n11208 = ~n11206 & ~n11207;
  assign n11209 = ~n11203 & n11208;
  assign n11210 = po47  & ~n11202;
  assign n11211 = ~po48  & ~n11210;
  assign n11212 = ~n11209 & n11211;
  assign n11213 = ~n11209 & ~n11210;
  assign n11214 = po48  & ~n11213;
  assign n11215 = n10914 & ~n11212;
  assign n11216 = ~n11214 & ~n11215;
  assign n11217 = po49  & ~n11216;
  assign n11218 = ~n10749 & ~n10751;
  assign n11219 = po16  & n11218;
  assign n11220 = n10756 & ~n11219;
  assign n11221 = ~n10756 & n11219;
  assign n11222 = ~n11220 & ~n11221;
  assign n11223 = ~po49  & n11216;
  assign n11224 = ~n11222 & ~n11223;
  assign n11225 = ~n11217 & ~n11224;
  assign n11226 = po50  & ~n11225;
  assign n11227 = ~po50  & ~n11217;
  assign n11228 = ~n11224 & n11227;
  assign n11229 = ~n10759 & po16 ;
  assign n11230 = ~n10765 & n11229;
  assign n11231 = n10764 & ~n11230;
  assign n11232 = n10766 & n11229;
  assign n11233 = ~n11231 & ~n11232;
  assign n11234 = ~n11228 & n11233;
  assign n11235 = ~n11226 & ~n11234;
  assign n11236 = po51  & ~n11235;
  assign n11237 = ~n10768 & ~n10770;
  assign n11238 = po16  & n11237;
  assign n11239 = n10775 & ~n11238;
  assign n11240 = ~n10775 & n11238;
  assign n11241 = ~n11239 & ~n11240;
  assign n11242 = ~po51  & n11235;
  assign n11243 = ~n11241 & ~n11242;
  assign n11244 = ~n11236 & ~n11243;
  assign n11245 = po52  & ~n11244;
  assign n11246 = ~po52  & ~n11236;
  assign n11247 = ~n11243 & n11246;
  assign n11248 = ~n10778 & po16 ;
  assign n11249 = ~n10784 & n11248;
  assign n11250 = n10783 & ~n11249;
  assign n11251 = n10785 & n11248;
  assign n11252 = ~n11250 & ~n11251;
  assign n11253 = ~n11247 & n11252;
  assign n11254 = ~n11245 & ~n11253;
  assign n11255 = po53  & ~n11254;
  assign n11256 = ~po53  & n11254;
  assign n11257 = ~n10787 & po16 ;
  assign n11258 = ~n10794 & n11257;
  assign n11259 = n10792 & ~n11258;
  assign n11260 = n10795 & n11257;
  assign n11261 = ~n11259 & ~n11260;
  assign n11262 = ~n11256 & n11261;
  assign n11263 = ~n11255 & ~n11262;
  assign n11264 = po54  & ~n11263;
  assign n11265 = ~po54  & ~n11255;
  assign n11266 = ~n11262 & n11265;
  assign n11267 = ~n10797 & po16 ;
  assign n11268 = ~n10803 & n11267;
  assign n11269 = n10802 & ~n11268;
  assign n11270 = n10804 & n11267;
  assign n11271 = ~n11269 & ~n11270;
  assign n11272 = ~n11266 & n11271;
  assign n11273 = ~n11264 & ~n11272;
  assign n11274 = po55  & ~n11273;
  assign n11275 = ~n10806 & ~n10808;
  assign n11276 = po16  & n11275;
  assign n11277 = n10813 & ~n11276;
  assign n11278 = ~n10813 & n11276;
  assign n11279 = ~n11277 & ~n11278;
  assign n11280 = ~po55  & n11273;
  assign n11281 = ~n11279 & ~n11280;
  assign n11282 = ~n11274 & ~n11281;
  assign n11283 = po56  & ~n11282;
  assign n11284 = ~po56  & ~n11274;
  assign n11285 = ~n11281 & n11284;
  assign n11286 = ~n10816 & po16 ;
  assign n11287 = ~n10822 & n11286;
  assign n11288 = n10821 & ~n11287;
  assign n11289 = n10823 & n11286;
  assign n11290 = ~n11288 & ~n11289;
  assign n11291 = ~n11285 & n11290;
  assign n11292 = ~n11283 & ~n11291;
  assign n11293 = po57  & ~n11292;
  assign n11294 = ~po57  & n11292;
  assign n11295 = ~n10825 & po16 ;
  assign n11296 = ~n10832 & n11295;
  assign n11297 = n10830 & ~n11296;
  assign n11298 = n10833 & n11295;
  assign n11299 = ~n11297 & ~n11298;
  assign n11300 = ~n11294 & n11299;
  assign n11301 = ~n11293 & ~n11300;
  assign n11302 = po58  & ~n11301;
  assign n11303 = ~po58  & ~n11293;
  assign n11304 = ~n11300 & n11303;
  assign n11305 = ~n10835 & po16 ;
  assign n11306 = ~n10841 & n11305;
  assign n11307 = n10840 & ~n11306;
  assign n11308 = n10842 & n11305;
  assign n11309 = ~n11307 & ~n11308;
  assign n11310 = ~n11304 & n11309;
  assign n11311 = ~n11302 & ~n11310;
  assign n11312 = po59  & ~n11311;
  assign n11313 = ~n10844 & ~n10846;
  assign n11314 = po16  & n11313;
  assign n11315 = n10851 & ~n11314;
  assign n11316 = ~n10851 & n11314;
  assign n11317 = ~n11315 & ~n11316;
  assign n11318 = ~po59  & n11311;
  assign n11319 = ~n11317 & ~n11318;
  assign n11320 = ~n11312 & ~n11319;
  assign n11321 = po60  & ~n11320;
  assign n11322 = ~po60  & ~n11312;
  assign n11323 = ~n11319 & n11322;
  assign n11324 = ~n10854 & po16 ;
  assign n11325 = ~n10860 & n11324;
  assign n11326 = n10859 & ~n11325;
  assign n11327 = n10861 & n11324;
  assign n11328 = ~n11326 & ~n11327;
  assign n11329 = ~n11323 & n11328;
  assign n11330 = ~n11321 & ~n11329;
  assign n11331 = po61  & ~n11330;
  assign n11332 = ~po61  & n11330;
  assign n11333 = ~n10863 & po16 ;
  assign n11334 = ~n10870 & n11333;
  assign n11335 = n10868 & ~n11334;
  assign n11336 = n10871 & n11333;
  assign n11337 = ~n11335 & ~n11336;
  assign n11338 = ~n11332 & n11337;
  assign n11339 = ~n11331 & ~n11338;
  assign n11340 = po62  & ~n11339;
  assign n11341 = ~po62  & ~n11331;
  assign n11342 = ~n11338 & n11341;
  assign n11343 = ~n10873 & po16 ;
  assign n11344 = ~n10879 & n11343;
  assign n11345 = n10878 & ~n11344;
  assign n11346 = n10880 & n11343;
  assign n11347 = ~n11345 & ~n11346;
  assign n11348 = ~n11342 & n11347;
  assign n11349 = ~n11340 & ~n11348;
  assign n11350 = ~n10882 & ~n10884;
  assign n11351 = po16  & n11350;
  assign n11352 = n10889 & ~n11351;
  assign n11353 = ~n10889 & n11351;
  assign n11354 = ~n11352 & ~n11353;
  assign n11355 = n10891 & po16 ;
  assign n11356 = ~n10898 & ~n11355;
  assign n11357 = ~n10903 & ~n11356;
  assign n11358 = po16  & ~n11357;
  assign n11359 = ~n11354 & ~n11358;
  assign n11360 = ~n11349 & n11359;
  assign n11361 = ~po63  & ~n11360;
  assign n11362 = n11349 & n11354;
  assign n11363 = po63  & n11357;
  assign n11364 = ~n11362 & ~n11363;
  assign po15  = n11361 | ~n11364;
  assign n11366 = ~n11212 & ~n11214;
  assign n11367 = po15  & n11366;
  assign n11368 = n10914 & ~n11367;
  assign n11369 = ~n10914 & n11367;
  assign n11370 = ~n11368 & ~n11369;
  assign n11371 = pi30  & po15 ;
  assign n11372 = ~pi28  & ~pi29 ;
  assign n11373 = ~pi30  & n11372;
  assign n11374 = ~n11371 & ~n11373;
  assign n11375 = po16  & ~n11374;
  assign n11376 = ~po16  & n11374;
  assign n11377 = ~pi30  & po15 ;
  assign n11378 = pi31  & ~n11377;
  assign n11379 = ~pi31  & n11377;
  assign n11380 = ~n11378 & ~n11379;
  assign n11381 = ~n11376 & n11380;
  assign n11382 = ~n11375 & ~n11381;
  assign n11383 = po17  & ~n11382;
  assign n11384 = po16  & ~po15 ;
  assign n11385 = ~n11379 & ~n11384;
  assign n11386 = pi32  & ~n11385;
  assign n11387 = ~pi32  & n11385;
  assign n11388 = ~n11386 & ~n11387;
  assign n11389 = ~po17  & n11382;
  assign n11390 = ~n11388 & ~n11389;
  assign n11391 = ~n11383 & ~n11390;
  assign n11392 = po18  & ~n11391;
  assign n11393 = ~po18  & ~n11383;
  assign n11394 = ~n11390 & n11393;
  assign n11395 = ~n10919 & ~n10924;
  assign n11396 = po15  & n11395;
  assign n11397 = n10923 & ~n11396;
  assign n11398 = ~n10923 & n11396;
  assign n11399 = ~n11397 & ~n11398;
  assign n11400 = ~n11394 & ~n11399;
  assign n11401 = ~n11392 & ~n11400;
  assign n11402 = po19  & ~n11401;
  assign n11403 = ~n10927 & ~n10929;
  assign n11404 = po15  & n11403;
  assign n11405 = ~n10934 & ~n11404;
  assign n11406 = n10934 & n11404;
  assign n11407 = ~n11405 & ~n11406;
  assign n11408 = ~po19  & n11401;
  assign n11409 = ~n11407 & ~n11408;
  assign n11410 = ~n11402 & ~n11409;
  assign n11411 = po20  & ~n11410;
  assign n11412 = ~po20  & ~n11402;
  assign n11413 = ~n11409 & n11412;
  assign n11414 = ~n10937 & ~n10938;
  assign n11415 = po15  & n11414;
  assign n11416 = n10943 & ~n11415;
  assign n11417 = ~n10943 & n11415;
  assign n11418 = ~n11416 & ~n11417;
  assign n11419 = ~n11413 & n11418;
  assign n11420 = ~n11411 & ~n11419;
  assign n11421 = po21  & ~n11420;
  assign n11422 = ~n10946 & ~n10948;
  assign n11423 = po15  & n11422;
  assign n11424 = n10953 & ~n11423;
  assign n11425 = ~n10953 & n11423;
  assign n11426 = ~n11424 & ~n11425;
  assign n11427 = ~po21  & n11420;
  assign n11428 = ~n11426 & ~n11427;
  assign n11429 = ~n11421 & ~n11428;
  assign n11430 = po22  & ~n11429;
  assign n11431 = ~po22  & ~n11421;
  assign n11432 = ~n11428 & n11431;
  assign n11433 = ~n10956 & ~n10957;
  assign n11434 = po15  & n11433;
  assign n11435 = n10962 & n11434;
  assign n11436 = ~n10962 & ~n11434;
  assign n11437 = ~n11435 & ~n11436;
  assign n11438 = ~n11432 & n11437;
  assign n11439 = ~n11430 & ~n11438;
  assign n11440 = po23  & ~n11439;
  assign n11441 = ~n10965 & ~n10967;
  assign n11442 = po15  & n11441;
  assign n11443 = n10972 & ~n11442;
  assign n11444 = ~n10972 & n11442;
  assign n11445 = ~n11443 & ~n11444;
  assign n11446 = ~po23  & n11439;
  assign n11447 = ~n11445 & ~n11446;
  assign n11448 = ~n11440 & ~n11447;
  assign n11449 = po24  & ~n11448;
  assign n11450 = ~po24  & ~n11440;
  assign n11451 = ~n11447 & n11450;
  assign n11452 = ~n10975 & ~n10976;
  assign n11453 = po15  & n11452;
  assign n11454 = ~n10981 & ~n11453;
  assign n11455 = n10981 & n11453;
  assign n11456 = ~n11454 & ~n11455;
  assign n11457 = ~n11451 & n11456;
  assign n11458 = ~n11449 & ~n11457;
  assign n11459 = po25  & ~n11458;
  assign n11460 = ~n10984 & ~n10986;
  assign n11461 = po15  & n11460;
  assign n11462 = n10991 & ~n11461;
  assign n11463 = ~n10991 & n11461;
  assign n11464 = ~n11462 & ~n11463;
  assign n11465 = ~po25  & n11458;
  assign n11466 = ~n11464 & ~n11465;
  assign n11467 = ~n11459 & ~n11466;
  assign n11468 = po26  & ~n11467;
  assign n11469 = ~n10994 & ~n10995;
  assign n11470 = po15  & n11469;
  assign n11471 = n11000 & ~n11470;
  assign n11472 = ~n11000 & n11470;
  assign n11473 = ~n11471 & ~n11472;
  assign n11474 = ~po26  & ~n11459;
  assign n11475 = ~n11466 & n11474;
  assign n11476 = ~n11473 & ~n11475;
  assign n11477 = ~n11468 & ~n11476;
  assign n11478 = po27  & ~n11477;
  assign n11479 = ~n11003 & ~n11005;
  assign n11480 = po15  & n11479;
  assign n11481 = n11010 & ~n11480;
  assign n11482 = ~n11010 & n11480;
  assign n11483 = ~n11481 & ~n11482;
  assign n11484 = ~po27  & n11477;
  assign n11485 = ~n11483 & ~n11484;
  assign n11486 = ~n11478 & ~n11485;
  assign n11487 = po28  & ~n11486;
  assign n11488 = ~po28  & ~n11478;
  assign n11489 = ~n11485 & n11488;
  assign n11490 = ~n11013 & po15 ;
  assign n11491 = ~n11019 & n11490;
  assign n11492 = n11018 & ~n11491;
  assign n11493 = n11020 & n11490;
  assign n11494 = ~n11492 & ~n11493;
  assign n11495 = ~n11489 & n11494;
  assign n11496 = ~n11487 & ~n11495;
  assign n11497 = po29  & ~n11496;
  assign n11498 = ~n11022 & ~n11024;
  assign n11499 = po15  & n11498;
  assign n11500 = n11029 & ~n11499;
  assign n11501 = ~n11029 & n11499;
  assign n11502 = ~n11500 & ~n11501;
  assign n11503 = ~po29  & n11496;
  assign n11504 = ~n11502 & ~n11503;
  assign n11505 = ~n11497 & ~n11504;
  assign n11506 = po30  & ~n11505;
  assign n11507 = ~n11032 & ~n11033;
  assign n11508 = po15  & n11507;
  assign n11509 = n11038 & ~n11508;
  assign n11510 = ~n11038 & n11508;
  assign n11511 = ~n11509 & ~n11510;
  assign n11512 = ~po30  & ~n11497;
  assign n11513 = ~n11504 & n11512;
  assign n11514 = ~n11511 & ~n11513;
  assign n11515 = ~n11506 & ~n11514;
  assign n11516 = po31  & ~n11515;
  assign n11517 = ~n11041 & ~n11043;
  assign n11518 = po15  & n11517;
  assign n11519 = n11048 & ~n11518;
  assign n11520 = ~n11048 & n11518;
  assign n11521 = ~n11519 & ~n11520;
  assign n11522 = ~po31  & n11515;
  assign n11523 = ~n11521 & ~n11522;
  assign n11524 = ~n11516 & ~n11523;
  assign n11525 = po32  & ~n11524;
  assign n11526 = ~po32  & ~n11516;
  assign n11527 = ~n11523 & n11526;
  assign n11528 = ~n11051 & po15 ;
  assign n11529 = ~n11057 & n11528;
  assign n11530 = n11056 & ~n11529;
  assign n11531 = n11058 & n11528;
  assign n11532 = ~n11530 & ~n11531;
  assign n11533 = ~n11527 & n11532;
  assign n11534 = ~n11525 & ~n11533;
  assign n11535 = po33  & ~n11534;
  assign n11536 = ~n11060 & ~n11062;
  assign n11537 = po15  & n11536;
  assign n11538 = n11067 & ~n11537;
  assign n11539 = ~n11067 & n11537;
  assign n11540 = ~n11538 & ~n11539;
  assign n11541 = ~po33  & n11534;
  assign n11542 = ~n11540 & ~n11541;
  assign n11543 = ~n11535 & ~n11542;
  assign n11544 = po34  & ~n11543;
  assign n11545 = ~n11070 & ~n11071;
  assign n11546 = po15  & n11545;
  assign n11547 = n11076 & ~n11546;
  assign n11548 = ~n11076 & n11546;
  assign n11549 = ~n11547 & ~n11548;
  assign n11550 = ~po34  & ~n11535;
  assign n11551 = ~n11542 & n11550;
  assign n11552 = ~n11549 & ~n11551;
  assign n11553 = ~n11544 & ~n11552;
  assign n11554 = po35  & ~n11553;
  assign n11555 = ~n11079 & ~n11081;
  assign n11556 = po15  & n11555;
  assign n11557 = n11086 & ~n11556;
  assign n11558 = ~n11086 & n11556;
  assign n11559 = ~n11557 & ~n11558;
  assign n11560 = ~po35  & n11553;
  assign n11561 = ~n11559 & ~n11560;
  assign n11562 = ~n11554 & ~n11561;
  assign n11563 = po36  & ~n11562;
  assign n11564 = ~po36  & ~n11554;
  assign n11565 = ~n11561 & n11564;
  assign n11566 = ~n11089 & po15 ;
  assign n11567 = ~n11095 & n11566;
  assign n11568 = n11094 & ~n11567;
  assign n11569 = n11096 & n11566;
  assign n11570 = ~n11568 & ~n11569;
  assign n11571 = ~n11565 & n11570;
  assign n11572 = ~n11563 & ~n11571;
  assign n11573 = po37  & ~n11572;
  assign n11574 = ~n11098 & ~n11100;
  assign n11575 = po15  & n11574;
  assign n11576 = n11105 & ~n11575;
  assign n11577 = ~n11105 & n11575;
  assign n11578 = ~n11576 & ~n11577;
  assign n11579 = ~po37  & n11572;
  assign n11580 = ~n11578 & ~n11579;
  assign n11581 = ~n11573 & ~n11580;
  assign n11582 = po38  & ~n11581;
  assign n11583 = ~n11108 & ~n11109;
  assign n11584 = po15  & n11583;
  assign n11585 = n11114 & ~n11584;
  assign n11586 = ~n11114 & n11584;
  assign n11587 = ~n11585 & ~n11586;
  assign n11588 = ~po38  & ~n11573;
  assign n11589 = ~n11580 & n11588;
  assign n11590 = ~n11587 & ~n11589;
  assign n11591 = ~n11582 & ~n11590;
  assign n11592 = po39  & ~n11591;
  assign n11593 = ~n11117 & ~n11119;
  assign n11594 = po15  & n11593;
  assign n11595 = n11124 & ~n11594;
  assign n11596 = ~n11124 & n11594;
  assign n11597 = ~n11595 & ~n11596;
  assign n11598 = ~po39  & n11591;
  assign n11599 = ~n11597 & ~n11598;
  assign n11600 = ~n11592 & ~n11599;
  assign n11601 = po40  & ~n11600;
  assign n11602 = ~po40  & ~n11592;
  assign n11603 = ~n11599 & n11602;
  assign n11604 = ~n11127 & po15 ;
  assign n11605 = ~n11133 & n11604;
  assign n11606 = n11132 & ~n11605;
  assign n11607 = n11134 & n11604;
  assign n11608 = ~n11606 & ~n11607;
  assign n11609 = ~n11603 & n11608;
  assign n11610 = ~n11601 & ~n11609;
  assign n11611 = po41  & ~n11610;
  assign n11612 = ~n11136 & ~n11138;
  assign n11613 = po15  & n11612;
  assign n11614 = n11143 & ~n11613;
  assign n11615 = ~n11143 & n11613;
  assign n11616 = ~n11614 & ~n11615;
  assign n11617 = ~po41  & n11610;
  assign n11618 = ~n11616 & ~n11617;
  assign n11619 = ~n11611 & ~n11618;
  assign n11620 = po42  & ~n11619;
  assign n11621 = ~n11146 & ~n11147;
  assign n11622 = po15  & n11621;
  assign n11623 = n11152 & ~n11622;
  assign n11624 = ~n11152 & n11622;
  assign n11625 = ~n11623 & ~n11624;
  assign n11626 = ~po42  & ~n11611;
  assign n11627 = ~n11618 & n11626;
  assign n11628 = ~n11625 & ~n11627;
  assign n11629 = ~n11620 & ~n11628;
  assign n11630 = po43  & ~n11629;
  assign n11631 = ~n11155 & ~n11157;
  assign n11632 = po15  & n11631;
  assign n11633 = n11162 & ~n11632;
  assign n11634 = ~n11162 & n11632;
  assign n11635 = ~n11633 & ~n11634;
  assign n11636 = ~po43  & n11629;
  assign n11637 = ~n11635 & ~n11636;
  assign n11638 = ~n11630 & ~n11637;
  assign n11639 = po44  & ~n11638;
  assign n11640 = ~po44  & ~n11630;
  assign n11641 = ~n11637 & n11640;
  assign n11642 = ~n11165 & po15 ;
  assign n11643 = ~n11171 & n11642;
  assign n11644 = n11170 & ~n11643;
  assign n11645 = n11172 & n11642;
  assign n11646 = ~n11644 & ~n11645;
  assign n11647 = ~n11641 & n11646;
  assign n11648 = ~n11639 & ~n11647;
  assign n11649 = po45  & ~n11648;
  assign n11650 = ~n11174 & ~n11176;
  assign n11651 = po15  & n11650;
  assign n11652 = n11181 & ~n11651;
  assign n11653 = ~n11181 & n11651;
  assign n11654 = ~n11652 & ~n11653;
  assign n11655 = ~po45  & n11648;
  assign n11656 = ~n11654 & ~n11655;
  assign n11657 = ~n11649 & ~n11656;
  assign n11658 = po46  & ~n11657;
  assign n11659 = ~n11184 & ~n11185;
  assign n11660 = po15  & n11659;
  assign n11661 = n11190 & ~n11660;
  assign n11662 = ~n11190 & n11660;
  assign n11663 = ~n11661 & ~n11662;
  assign n11664 = ~po46  & ~n11649;
  assign n11665 = ~n11656 & n11664;
  assign n11666 = ~n11663 & ~n11665;
  assign n11667 = ~n11658 & ~n11666;
  assign n11668 = ~po47  & n11667;
  assign n11669 = ~n11193 & po15 ;
  assign n11670 = ~n11200 & n11669;
  assign n11671 = n11198 & ~n11670;
  assign n11672 = n11201 & n11669;
  assign n11673 = ~n11671 & ~n11672;
  assign n11674 = ~n11668 & n11673;
  assign n11675 = po47  & ~n11667;
  assign n11676 = ~n11674 & ~n11675;
  assign n11677 = po48  & ~n11676;
  assign n11678 = ~n11203 & ~n11210;
  assign n11679 = po15  & n11678;
  assign n11680 = ~n11208 & ~n11679;
  assign n11681 = n11208 & n11679;
  assign n11682 = ~n11680 & ~n11681;
  assign n11683 = ~po48  & ~n11675;
  assign n11684 = ~n11674 & n11683;
  assign n11685 = n11682 & ~n11684;
  assign n11686 = ~n11677 & ~n11685;
  assign n11687 = ~po49  & n11686;
  assign n11688 = po49  & ~n11686;
  assign n11689 = ~n11370 & ~n11687;
  assign n11690 = ~n11688 & ~n11689;
  assign n11691 = po50  & ~n11690;
  assign n11692 = ~po50  & ~n11688;
  assign n11693 = ~n11689 & n11692;
  assign n11694 = ~n11217 & po15 ;
  assign n11695 = ~n11223 & n11694;
  assign n11696 = n11222 & ~n11695;
  assign n11697 = n11224 & n11694;
  assign n11698 = ~n11696 & ~n11697;
  assign n11699 = ~n11693 & n11698;
  assign n11700 = ~n11691 & ~n11699;
  assign n11701 = po51  & ~n11700;
  assign n11702 = ~n11226 & ~n11228;
  assign n11703 = po15  & n11702;
  assign n11704 = n11233 & ~n11703;
  assign n11705 = ~n11233 & n11703;
  assign n11706 = ~n11704 & ~n11705;
  assign n11707 = ~po51  & n11700;
  assign n11708 = ~n11706 & ~n11707;
  assign n11709 = ~n11701 & ~n11708;
  assign n11710 = po52  & ~n11709;
  assign n11711 = ~po52  & ~n11701;
  assign n11712 = ~n11708 & n11711;
  assign n11713 = ~n11236 & po15 ;
  assign n11714 = ~n11242 & n11713;
  assign n11715 = n11241 & ~n11714;
  assign n11716 = n11243 & n11713;
  assign n11717 = ~n11715 & ~n11716;
  assign n11718 = ~n11712 & n11717;
  assign n11719 = ~n11710 & ~n11718;
  assign n11720 = po53  & ~n11719;
  assign n11721 = ~n11245 & ~n11247;
  assign n11722 = po15  & n11721;
  assign n11723 = n11252 & ~n11722;
  assign n11724 = ~n11252 & n11722;
  assign n11725 = ~n11723 & ~n11724;
  assign n11726 = ~po53  & n11719;
  assign n11727 = ~n11725 & ~n11726;
  assign n11728 = ~n11720 & ~n11727;
  assign n11729 = po54  & ~n11728;
  assign n11730 = ~n11255 & ~n11256;
  assign n11731 = po15  & n11730;
  assign n11732 = n11261 & ~n11731;
  assign n11733 = ~n11261 & n11731;
  assign n11734 = ~n11732 & ~n11733;
  assign n11735 = ~po54  & ~n11720;
  assign n11736 = ~n11727 & n11735;
  assign n11737 = ~n11734 & ~n11736;
  assign n11738 = ~n11729 & ~n11737;
  assign n11739 = po55  & ~n11738;
  assign n11740 = ~n11264 & ~n11266;
  assign n11741 = po15  & n11740;
  assign n11742 = n11271 & ~n11741;
  assign n11743 = ~n11271 & n11741;
  assign n11744 = ~n11742 & ~n11743;
  assign n11745 = ~po55  & n11738;
  assign n11746 = ~n11744 & ~n11745;
  assign n11747 = ~n11739 & ~n11746;
  assign n11748 = po56  & ~n11747;
  assign n11749 = ~po56  & ~n11739;
  assign n11750 = ~n11746 & n11749;
  assign n11751 = ~n11274 & po15 ;
  assign n11752 = ~n11280 & n11751;
  assign n11753 = n11279 & ~n11752;
  assign n11754 = n11281 & n11751;
  assign n11755 = ~n11753 & ~n11754;
  assign n11756 = ~n11750 & n11755;
  assign n11757 = ~n11748 & ~n11756;
  assign n11758 = po57  & ~n11757;
  assign n11759 = ~n11283 & ~n11285;
  assign n11760 = po15  & n11759;
  assign n11761 = n11290 & ~n11760;
  assign n11762 = ~n11290 & n11760;
  assign n11763 = ~n11761 & ~n11762;
  assign n11764 = ~po57  & n11757;
  assign n11765 = ~n11763 & ~n11764;
  assign n11766 = ~n11758 & ~n11765;
  assign n11767 = po58  & ~n11766;
  assign n11768 = ~n11293 & ~n11294;
  assign n11769 = po15  & n11768;
  assign n11770 = n11299 & ~n11769;
  assign n11771 = ~n11299 & n11769;
  assign n11772 = ~n11770 & ~n11771;
  assign n11773 = ~po58  & ~n11758;
  assign n11774 = ~n11765 & n11773;
  assign n11775 = ~n11772 & ~n11774;
  assign n11776 = ~n11767 & ~n11775;
  assign n11777 = po59  & ~n11776;
  assign n11778 = ~n11302 & ~n11304;
  assign n11779 = po15  & n11778;
  assign n11780 = n11309 & ~n11779;
  assign n11781 = ~n11309 & n11779;
  assign n11782 = ~n11780 & ~n11781;
  assign n11783 = ~po59  & n11776;
  assign n11784 = ~n11782 & ~n11783;
  assign n11785 = ~n11777 & ~n11784;
  assign n11786 = po60  & ~n11785;
  assign n11787 = ~po60  & ~n11777;
  assign n11788 = ~n11784 & n11787;
  assign n11789 = ~n11312 & po15 ;
  assign n11790 = ~n11318 & n11789;
  assign n11791 = n11317 & ~n11790;
  assign n11792 = n11319 & n11789;
  assign n11793 = ~n11791 & ~n11792;
  assign n11794 = ~n11788 & n11793;
  assign n11795 = ~n11786 & ~n11794;
  assign n11796 = po61  & ~n11795;
  assign n11797 = ~n11321 & ~n11323;
  assign n11798 = po15  & n11797;
  assign n11799 = n11328 & ~n11798;
  assign n11800 = ~n11328 & n11798;
  assign n11801 = ~n11799 & ~n11800;
  assign n11802 = ~po61  & n11795;
  assign n11803 = ~n11801 & ~n11802;
  assign n11804 = ~n11796 & ~n11803;
  assign n11805 = po62  & ~n11804;
  assign n11806 = ~n11331 & ~n11332;
  assign n11807 = po15  & n11806;
  assign n11808 = n11337 & ~n11807;
  assign n11809 = ~n11337 & n11807;
  assign n11810 = ~n11808 & ~n11809;
  assign n11811 = ~po62  & ~n11796;
  assign n11812 = ~n11803 & n11811;
  assign n11813 = ~n11810 & ~n11812;
  assign n11814 = ~n11805 & ~n11813;
  assign n11815 = ~n11340 & ~n11342;
  assign n11816 = po15  & n11815;
  assign n11817 = n11347 & ~n11816;
  assign n11818 = ~n11347 & n11816;
  assign n11819 = ~n11817 & ~n11818;
  assign n11820 = n11349 & po15 ;
  assign n11821 = ~n11354 & ~n11820;
  assign n11822 = ~n11362 & ~n11821;
  assign n11823 = po15  & ~n11822;
  assign n11824 = ~n11819 & ~n11823;
  assign n11825 = ~n11814 & n11824;
  assign n11826 = ~po63  & ~n11825;
  assign n11827 = n11814 & n11819;
  assign n11828 = po63  & n11822;
  assign n11829 = ~n11827 & ~n11828;
  assign po14  = n11826 | ~n11829;
  assign n11831 = ~n11688 & po14 ;
  assign n11832 = ~n11687 & n11831;
  assign n11833 = n11370 & ~n11832;
  assign n11834 = n11689 & n11831;
  assign n11835 = ~n11833 & ~n11834;
  assign n11836 = ~n11677 & ~n11684;
  assign n11837 = po14  & n11836;
  assign n11838 = n11682 & ~n11837;
  assign n11839 = ~n11682 & n11837;
  assign n11840 = ~n11838 & ~n11839;
  assign n11841 = pi28  & po14 ;
  assign n11842 = ~pi26  & ~pi27 ;
  assign n11843 = ~pi28  & n11842;
  assign n11844 = ~n11841 & ~n11843;
  assign n11845 = po15  & ~n11844;
  assign n11846 = ~pi28  & po14 ;
  assign n11847 = pi29  & ~n11846;
  assign n11848 = ~pi29  & n11846;
  assign n11849 = ~n11847 & ~n11848;
  assign n11850 = ~po15  & n11844;
  assign n11851 = n11849 & ~n11850;
  assign n11852 = ~n11845 & ~n11851;
  assign n11853 = po16  & ~n11852;
  assign n11854 = ~po16  & ~n11845;
  assign n11855 = ~n11851 & n11854;
  assign n11856 = po15  & ~po14 ;
  assign n11857 = ~n11848 & ~n11856;
  assign n11858 = pi30  & ~n11857;
  assign n11859 = ~pi30  & n11857;
  assign n11860 = ~n11858 & ~n11859;
  assign n11861 = ~n11855 & ~n11860;
  assign n11862 = ~n11853 & ~n11861;
  assign n11863 = po17  & ~n11862;
  assign n11864 = ~po17  & n11862;
  assign n11865 = ~n11375 & ~n11376;
  assign n11866 = po14  & n11865;
  assign n11867 = n11380 & ~n11866;
  assign n11868 = ~n11380 & n11866;
  assign n11869 = ~n11867 & ~n11868;
  assign n11870 = ~n11864 & ~n11869;
  assign n11871 = ~n11863 & ~n11870;
  assign n11872 = po18  & ~n11871;
  assign n11873 = ~po18  & ~n11863;
  assign n11874 = ~n11870 & n11873;
  assign n11875 = ~n11383 & po14 ;
  assign n11876 = ~n11389 & n11875;
  assign n11877 = n11388 & ~n11876;
  assign n11878 = n11390 & n11875;
  assign n11879 = ~n11877 & ~n11878;
  assign n11880 = ~n11874 & n11879;
  assign n11881 = ~n11872 & ~n11880;
  assign n11882 = po19  & ~n11881;
  assign n11883 = ~po19  & n11881;
  assign n11884 = ~n11392 & ~n11394;
  assign n11885 = po14  & n11884;
  assign n11886 = n11399 & ~n11885;
  assign n11887 = ~n11399 & n11885;
  assign n11888 = ~n11886 & ~n11887;
  assign n11889 = ~n11883 & n11888;
  assign n11890 = ~n11882 & ~n11889;
  assign n11891 = po20  & ~n11890;
  assign n11892 = ~po20  & ~n11882;
  assign n11893 = ~n11889 & n11892;
  assign n11894 = ~n11402 & po14 ;
  assign n11895 = ~n11408 & n11894;
  assign n11896 = n11407 & ~n11895;
  assign n11897 = n11409 & n11894;
  assign n11898 = ~n11896 & ~n11897;
  assign n11899 = ~n11893 & n11898;
  assign n11900 = ~n11891 & ~n11899;
  assign n11901 = po21  & ~n11900;
  assign n11902 = ~po21  & n11900;
  assign n11903 = ~n11411 & ~n11413;
  assign n11904 = po14  & n11903;
  assign n11905 = n11418 & n11904;
  assign n11906 = ~n11418 & ~n11904;
  assign n11907 = ~n11905 & ~n11906;
  assign n11908 = ~n11902 & n11907;
  assign n11909 = ~n11901 & ~n11908;
  assign n11910 = po22  & ~n11909;
  assign n11911 = ~po22  & ~n11901;
  assign n11912 = ~n11908 & n11911;
  assign n11913 = ~n11421 & po14 ;
  assign n11914 = ~n11427 & n11913;
  assign n11915 = n11426 & ~n11914;
  assign n11916 = n11428 & n11913;
  assign n11917 = ~n11915 & ~n11916;
  assign n11918 = ~n11912 & n11917;
  assign n11919 = ~n11910 & ~n11918;
  assign n11920 = po23  & ~n11919;
  assign n11921 = ~po23  & n11919;
  assign n11922 = ~n11430 & ~n11432;
  assign n11923 = po14  & n11922;
  assign n11924 = ~n11437 & ~n11923;
  assign n11925 = n11437 & n11923;
  assign n11926 = ~n11924 & ~n11925;
  assign n11927 = ~n11921 & n11926;
  assign n11928 = ~n11920 & ~n11927;
  assign n11929 = po24  & ~n11928;
  assign n11930 = ~po24  & ~n11920;
  assign n11931 = ~n11927 & n11930;
  assign n11932 = ~n11440 & po14 ;
  assign n11933 = ~n11446 & n11932;
  assign n11934 = n11445 & ~n11933;
  assign n11935 = n11447 & n11932;
  assign n11936 = ~n11934 & ~n11935;
  assign n11937 = ~n11931 & n11936;
  assign n11938 = ~n11929 & ~n11937;
  assign n11939 = po25  & ~n11938;
  assign n11940 = ~n11449 & ~n11451;
  assign n11941 = po14  & n11940;
  assign n11942 = n11456 & ~n11941;
  assign n11943 = ~n11456 & n11941;
  assign n11944 = ~n11942 & ~n11943;
  assign n11945 = ~po25  & n11938;
  assign n11946 = ~n11944 & ~n11945;
  assign n11947 = ~n11939 & ~n11946;
  assign n11948 = po26  & ~n11947;
  assign n11949 = ~po26  & ~n11939;
  assign n11950 = ~n11946 & n11949;
  assign n11951 = ~n11459 & po14 ;
  assign n11952 = ~n11465 & n11951;
  assign n11953 = n11464 & ~n11952;
  assign n11954 = n11466 & n11951;
  assign n11955 = ~n11953 & ~n11954;
  assign n11956 = ~n11950 & n11955;
  assign n11957 = ~n11948 & ~n11956;
  assign n11958 = po27  & ~n11957;
  assign n11959 = ~po27  & n11957;
  assign n11960 = ~n11468 & po14 ;
  assign n11961 = ~n11475 & n11960;
  assign n11962 = n11473 & ~n11961;
  assign n11963 = n11476 & n11960;
  assign n11964 = ~n11962 & ~n11963;
  assign n11965 = ~n11959 & n11964;
  assign n11966 = ~n11958 & ~n11965;
  assign n11967 = po28  & ~n11966;
  assign n11968 = ~po28  & ~n11958;
  assign n11969 = ~n11965 & n11968;
  assign n11970 = ~n11478 & po14 ;
  assign n11971 = ~n11484 & n11970;
  assign n11972 = n11483 & ~n11971;
  assign n11973 = n11485 & n11970;
  assign n11974 = ~n11972 & ~n11973;
  assign n11975 = ~n11969 & n11974;
  assign n11976 = ~n11967 & ~n11975;
  assign n11977 = po29  & ~n11976;
  assign n11978 = ~n11487 & ~n11489;
  assign n11979 = po14  & n11978;
  assign n11980 = n11494 & ~n11979;
  assign n11981 = ~n11494 & n11979;
  assign n11982 = ~n11980 & ~n11981;
  assign n11983 = ~po29  & n11976;
  assign n11984 = ~n11982 & ~n11983;
  assign n11985 = ~n11977 & ~n11984;
  assign n11986 = po30  & ~n11985;
  assign n11987 = ~po30  & ~n11977;
  assign n11988 = ~n11984 & n11987;
  assign n11989 = ~n11497 & po14 ;
  assign n11990 = ~n11503 & n11989;
  assign n11991 = n11502 & ~n11990;
  assign n11992 = n11504 & n11989;
  assign n11993 = ~n11991 & ~n11992;
  assign n11994 = ~n11988 & n11993;
  assign n11995 = ~n11986 & ~n11994;
  assign n11996 = po31  & ~n11995;
  assign n11997 = ~po31  & n11995;
  assign n11998 = ~n11506 & po14 ;
  assign n11999 = ~n11513 & n11998;
  assign n12000 = n11511 & ~n11999;
  assign n12001 = n11514 & n11998;
  assign n12002 = ~n12000 & ~n12001;
  assign n12003 = ~n11997 & n12002;
  assign n12004 = ~n11996 & ~n12003;
  assign n12005 = po32  & ~n12004;
  assign n12006 = ~po32  & ~n11996;
  assign n12007 = ~n12003 & n12006;
  assign n12008 = ~n11516 & po14 ;
  assign n12009 = ~n11522 & n12008;
  assign n12010 = n11521 & ~n12009;
  assign n12011 = n11523 & n12008;
  assign n12012 = ~n12010 & ~n12011;
  assign n12013 = ~n12007 & n12012;
  assign n12014 = ~n12005 & ~n12013;
  assign n12015 = po33  & ~n12014;
  assign n12016 = ~n11525 & ~n11527;
  assign n12017 = po14  & n12016;
  assign n12018 = n11532 & ~n12017;
  assign n12019 = ~n11532 & n12017;
  assign n12020 = ~n12018 & ~n12019;
  assign n12021 = ~po33  & n12014;
  assign n12022 = ~n12020 & ~n12021;
  assign n12023 = ~n12015 & ~n12022;
  assign n12024 = po34  & ~n12023;
  assign n12025 = ~po34  & ~n12015;
  assign n12026 = ~n12022 & n12025;
  assign n12027 = ~n11535 & po14 ;
  assign n12028 = ~n11541 & n12027;
  assign n12029 = n11540 & ~n12028;
  assign n12030 = n11542 & n12027;
  assign n12031 = ~n12029 & ~n12030;
  assign n12032 = ~n12026 & n12031;
  assign n12033 = ~n12024 & ~n12032;
  assign n12034 = po35  & ~n12033;
  assign n12035 = ~po35  & n12033;
  assign n12036 = ~n11544 & po14 ;
  assign n12037 = ~n11551 & n12036;
  assign n12038 = n11549 & ~n12037;
  assign n12039 = n11552 & n12036;
  assign n12040 = ~n12038 & ~n12039;
  assign n12041 = ~n12035 & n12040;
  assign n12042 = ~n12034 & ~n12041;
  assign n12043 = po36  & ~n12042;
  assign n12044 = ~po36  & ~n12034;
  assign n12045 = ~n12041 & n12044;
  assign n12046 = ~n11554 & po14 ;
  assign n12047 = ~n11560 & n12046;
  assign n12048 = n11559 & ~n12047;
  assign n12049 = n11561 & n12046;
  assign n12050 = ~n12048 & ~n12049;
  assign n12051 = ~n12045 & n12050;
  assign n12052 = ~n12043 & ~n12051;
  assign n12053 = po37  & ~n12052;
  assign n12054 = ~n11563 & ~n11565;
  assign n12055 = po14  & n12054;
  assign n12056 = n11570 & ~n12055;
  assign n12057 = ~n11570 & n12055;
  assign n12058 = ~n12056 & ~n12057;
  assign n12059 = ~po37  & n12052;
  assign n12060 = ~n12058 & ~n12059;
  assign n12061 = ~n12053 & ~n12060;
  assign n12062 = po38  & ~n12061;
  assign n12063 = ~po38  & ~n12053;
  assign n12064 = ~n12060 & n12063;
  assign n12065 = ~n11573 & po14 ;
  assign n12066 = ~n11579 & n12065;
  assign n12067 = n11578 & ~n12066;
  assign n12068 = n11580 & n12065;
  assign n12069 = ~n12067 & ~n12068;
  assign n12070 = ~n12064 & n12069;
  assign n12071 = ~n12062 & ~n12070;
  assign n12072 = po39  & ~n12071;
  assign n12073 = ~po39  & n12071;
  assign n12074 = ~n11582 & po14 ;
  assign n12075 = ~n11589 & n12074;
  assign n12076 = n11587 & ~n12075;
  assign n12077 = n11590 & n12074;
  assign n12078 = ~n12076 & ~n12077;
  assign n12079 = ~n12073 & n12078;
  assign n12080 = ~n12072 & ~n12079;
  assign n12081 = po40  & ~n12080;
  assign n12082 = ~po40  & ~n12072;
  assign n12083 = ~n12079 & n12082;
  assign n12084 = ~n11592 & po14 ;
  assign n12085 = ~n11598 & n12084;
  assign n12086 = n11597 & ~n12085;
  assign n12087 = n11599 & n12084;
  assign n12088 = ~n12086 & ~n12087;
  assign n12089 = ~n12083 & n12088;
  assign n12090 = ~n12081 & ~n12089;
  assign n12091 = po41  & ~n12090;
  assign n12092 = ~n11601 & ~n11603;
  assign n12093 = po14  & n12092;
  assign n12094 = n11608 & ~n12093;
  assign n12095 = ~n11608 & n12093;
  assign n12096 = ~n12094 & ~n12095;
  assign n12097 = ~po41  & n12090;
  assign n12098 = ~n12096 & ~n12097;
  assign n12099 = ~n12091 & ~n12098;
  assign n12100 = po42  & ~n12099;
  assign n12101 = ~po42  & ~n12091;
  assign n12102 = ~n12098 & n12101;
  assign n12103 = ~n11611 & po14 ;
  assign n12104 = ~n11617 & n12103;
  assign n12105 = n11616 & ~n12104;
  assign n12106 = n11618 & n12103;
  assign n12107 = ~n12105 & ~n12106;
  assign n12108 = ~n12102 & n12107;
  assign n12109 = ~n12100 & ~n12108;
  assign n12110 = po43  & ~n12109;
  assign n12111 = ~po43  & n12109;
  assign n12112 = ~n11620 & po14 ;
  assign n12113 = ~n11627 & n12112;
  assign n12114 = n11625 & ~n12113;
  assign n12115 = n11628 & n12112;
  assign n12116 = ~n12114 & ~n12115;
  assign n12117 = ~n12111 & n12116;
  assign n12118 = ~n12110 & ~n12117;
  assign n12119 = po44  & ~n12118;
  assign n12120 = ~po44  & ~n12110;
  assign n12121 = ~n12117 & n12120;
  assign n12122 = ~n11630 & po14 ;
  assign n12123 = ~n11636 & n12122;
  assign n12124 = n11635 & ~n12123;
  assign n12125 = n11637 & n12122;
  assign n12126 = ~n12124 & ~n12125;
  assign n12127 = ~n12121 & n12126;
  assign n12128 = ~n12119 & ~n12127;
  assign n12129 = po45  & ~n12128;
  assign n12130 = ~n11639 & ~n11641;
  assign n12131 = po14  & n12130;
  assign n12132 = n11646 & ~n12131;
  assign n12133 = ~n11646 & n12131;
  assign n12134 = ~n12132 & ~n12133;
  assign n12135 = ~po45  & n12128;
  assign n12136 = ~n12134 & ~n12135;
  assign n12137 = ~n12129 & ~n12136;
  assign n12138 = po46  & ~n12137;
  assign n12139 = ~po46  & ~n12129;
  assign n12140 = ~n12136 & n12139;
  assign n12141 = ~n11649 & po14 ;
  assign n12142 = ~n11655 & n12141;
  assign n12143 = n11654 & ~n12142;
  assign n12144 = n11656 & n12141;
  assign n12145 = ~n12143 & ~n12144;
  assign n12146 = ~n12140 & n12145;
  assign n12147 = ~n12138 & ~n12146;
  assign n12148 = po47  & ~n12147;
  assign n12149 = ~po47  & n12147;
  assign n12150 = ~n11658 & po14 ;
  assign n12151 = ~n11665 & n12150;
  assign n12152 = n11663 & ~n12151;
  assign n12153 = n11666 & n12150;
  assign n12154 = ~n12152 & ~n12153;
  assign n12155 = ~n12149 & n12154;
  assign n12156 = ~n12148 & ~n12155;
  assign n12157 = po48  & ~n12156;
  assign n12158 = ~n11668 & ~n11675;
  assign n12159 = po14  & n12158;
  assign n12160 = n11673 & ~n12159;
  assign n12161 = ~n11673 & n12159;
  assign n12162 = ~n12160 & ~n12161;
  assign n12163 = ~po48  & ~n12148;
  assign n12164 = ~n12155 & n12163;
  assign n12165 = ~n12162 & ~n12164;
  assign n12166 = ~n12157 & ~n12165;
  assign n12167 = ~po49  & n12166;
  assign n12168 = ~n11840 & ~n12167;
  assign n12169 = po49  & ~n12166;
  assign n12170 = ~po50  & ~n12169;
  assign n12171 = ~n12168 & n12170;
  assign n12172 = ~n12168 & ~n12169;
  assign n12173 = po50  & ~n12172;
  assign n12174 = n11835 & ~n12171;
  assign n12175 = ~n12173 & ~n12174;
  assign n12176 = po51  & ~n12175;
  assign n12177 = ~n11691 & ~n11693;
  assign n12178 = po14  & n12177;
  assign n12179 = n11698 & ~n12178;
  assign n12180 = ~n11698 & n12178;
  assign n12181 = ~n12179 & ~n12180;
  assign n12182 = ~po51  & n12175;
  assign n12183 = ~n12181 & ~n12182;
  assign n12184 = ~n12176 & ~n12183;
  assign n12185 = po52  & ~n12184;
  assign n12186 = ~po52  & ~n12176;
  assign n12187 = ~n12183 & n12186;
  assign n12188 = ~n11701 & po14 ;
  assign n12189 = ~n11707 & n12188;
  assign n12190 = n11706 & ~n12189;
  assign n12191 = n11708 & n12188;
  assign n12192 = ~n12190 & ~n12191;
  assign n12193 = ~n12187 & n12192;
  assign n12194 = ~n12185 & ~n12193;
  assign n12195 = po53  & ~n12194;
  assign n12196 = ~n11710 & ~n11712;
  assign n12197 = po14  & n12196;
  assign n12198 = n11717 & ~n12197;
  assign n12199 = ~n11717 & n12197;
  assign n12200 = ~n12198 & ~n12199;
  assign n12201 = ~po53  & n12194;
  assign n12202 = ~n12200 & ~n12201;
  assign n12203 = ~n12195 & ~n12202;
  assign n12204 = po54  & ~n12203;
  assign n12205 = ~po54  & ~n12195;
  assign n12206 = ~n12202 & n12205;
  assign n12207 = ~n11720 & po14 ;
  assign n12208 = ~n11726 & n12207;
  assign n12209 = n11725 & ~n12208;
  assign n12210 = n11727 & n12207;
  assign n12211 = ~n12209 & ~n12210;
  assign n12212 = ~n12206 & n12211;
  assign n12213 = ~n12204 & ~n12212;
  assign n12214 = po55  & ~n12213;
  assign n12215 = ~po55  & n12213;
  assign n12216 = ~n11729 & po14 ;
  assign n12217 = ~n11736 & n12216;
  assign n12218 = n11734 & ~n12217;
  assign n12219 = n11737 & n12216;
  assign n12220 = ~n12218 & ~n12219;
  assign n12221 = ~n12215 & n12220;
  assign n12222 = ~n12214 & ~n12221;
  assign n12223 = po56  & ~n12222;
  assign n12224 = ~po56  & ~n12214;
  assign n12225 = ~n12221 & n12224;
  assign n12226 = ~n11739 & po14 ;
  assign n12227 = ~n11745 & n12226;
  assign n12228 = n11744 & ~n12227;
  assign n12229 = n11746 & n12226;
  assign n12230 = ~n12228 & ~n12229;
  assign n12231 = ~n12225 & n12230;
  assign n12232 = ~n12223 & ~n12231;
  assign n12233 = po57  & ~n12232;
  assign n12234 = ~n11748 & ~n11750;
  assign n12235 = po14  & n12234;
  assign n12236 = n11755 & ~n12235;
  assign n12237 = ~n11755 & n12235;
  assign n12238 = ~n12236 & ~n12237;
  assign n12239 = ~po57  & n12232;
  assign n12240 = ~n12238 & ~n12239;
  assign n12241 = ~n12233 & ~n12240;
  assign n12242 = po58  & ~n12241;
  assign n12243 = ~po58  & ~n12233;
  assign n12244 = ~n12240 & n12243;
  assign n12245 = ~n11758 & po14 ;
  assign n12246 = ~n11764 & n12245;
  assign n12247 = n11763 & ~n12246;
  assign n12248 = n11765 & n12245;
  assign n12249 = ~n12247 & ~n12248;
  assign n12250 = ~n12244 & n12249;
  assign n12251 = ~n12242 & ~n12250;
  assign n12252 = po59  & ~n12251;
  assign n12253 = ~po59  & n12251;
  assign n12254 = ~n11767 & po14 ;
  assign n12255 = ~n11774 & n12254;
  assign n12256 = n11772 & ~n12255;
  assign n12257 = n11775 & n12254;
  assign n12258 = ~n12256 & ~n12257;
  assign n12259 = ~n12253 & n12258;
  assign n12260 = ~n12252 & ~n12259;
  assign n12261 = po60  & ~n12260;
  assign n12262 = ~po60  & ~n12252;
  assign n12263 = ~n12259 & n12262;
  assign n12264 = ~n11777 & po14 ;
  assign n12265 = ~n11783 & n12264;
  assign n12266 = n11782 & ~n12265;
  assign n12267 = n11784 & n12264;
  assign n12268 = ~n12266 & ~n12267;
  assign n12269 = ~n12263 & n12268;
  assign n12270 = ~n12261 & ~n12269;
  assign n12271 = po61  & ~n12270;
  assign n12272 = ~n11786 & ~n11788;
  assign n12273 = po14  & n12272;
  assign n12274 = n11793 & ~n12273;
  assign n12275 = ~n11793 & n12273;
  assign n12276 = ~n12274 & ~n12275;
  assign n12277 = ~po61  & n12270;
  assign n12278 = ~n12276 & ~n12277;
  assign n12279 = ~n12271 & ~n12278;
  assign n12280 = po62  & ~n12279;
  assign n12281 = ~po62  & ~n12271;
  assign n12282 = ~n12278 & n12281;
  assign n12283 = ~n11796 & po14 ;
  assign n12284 = ~n11802 & n12283;
  assign n12285 = n11801 & ~n12284;
  assign n12286 = n11803 & n12283;
  assign n12287 = ~n12285 & ~n12286;
  assign n12288 = ~n12282 & n12287;
  assign n12289 = ~n12280 & ~n12288;
  assign n12290 = n11814 & po14 ;
  assign n12291 = ~n11819 & ~n12290;
  assign n12292 = ~n11827 & ~n12291;
  assign n12293 = po14  & ~n12292;
  assign n12294 = ~n11805 & po14 ;
  assign n12295 = ~n11812 & n12294;
  assign n12296 = n11810 & ~n12295;
  assign n12297 = n11813 & n12294;
  assign n12298 = ~n12296 & ~n12297;
  assign n12299 = ~n12293 & n12298;
  assign n12300 = ~n12289 & n12299;
  assign n12301 = ~po63  & ~n12300;
  assign n12302 = n12289 & ~n12298;
  assign n12303 = po63  & n12292;
  assign n12304 = ~n12302 & ~n12303;
  assign po13  = n12301 | ~n12304;
  assign n12306 = ~n12171 & ~n12173;
  assign n12307 = po13  & n12306;
  assign n12308 = n11835 & ~n12307;
  assign n12309 = ~n11835 & n12307;
  assign n12310 = ~n12308 & ~n12309;
  assign n12311 = pi26  & po13 ;
  assign n12312 = ~pi24  & ~pi25 ;
  assign n12313 = ~pi26  & n12312;
  assign n12314 = ~n12311 & ~n12313;
  assign n12315 = po14  & ~n12314;
  assign n12316 = ~po14  & n12314;
  assign n12317 = ~pi26  & po13 ;
  assign n12318 = pi27  & ~n12317;
  assign n12319 = ~pi27  & n12317;
  assign n12320 = ~n12318 & ~n12319;
  assign n12321 = ~n12316 & n12320;
  assign n12322 = ~n12315 & ~n12321;
  assign n12323 = po15  & ~n12322;
  assign n12324 = po14  & ~po13 ;
  assign n12325 = ~n12319 & ~n12324;
  assign n12326 = pi28  & ~n12325;
  assign n12327 = ~pi28  & n12325;
  assign n12328 = ~n12326 & ~n12327;
  assign n12329 = ~po15  & n12322;
  assign n12330 = ~n12328 & ~n12329;
  assign n12331 = ~n12323 & ~n12330;
  assign n12332 = po16  & ~n12331;
  assign n12333 = ~po16  & ~n12323;
  assign n12334 = ~n12330 & n12333;
  assign n12335 = ~n11845 & ~n11850;
  assign n12336 = po13  & n12335;
  assign n12337 = n11849 & ~n12336;
  assign n12338 = ~n11849 & n12336;
  assign n12339 = ~n12337 & ~n12338;
  assign n12340 = ~n12334 & ~n12339;
  assign n12341 = ~n12332 & ~n12340;
  assign n12342 = po17  & ~n12341;
  assign n12343 = ~n11853 & ~n11855;
  assign n12344 = po13  & n12343;
  assign n12345 = ~n11860 & ~n12344;
  assign n12346 = n11860 & n12344;
  assign n12347 = ~n12345 & ~n12346;
  assign n12348 = ~po17  & n12341;
  assign n12349 = ~n12347 & ~n12348;
  assign n12350 = ~n12342 & ~n12349;
  assign n12351 = po18  & ~n12350;
  assign n12352 = ~po18  & ~n12342;
  assign n12353 = ~n12349 & n12352;
  assign n12354 = ~n11863 & ~n11864;
  assign n12355 = po13  & n12354;
  assign n12356 = n11869 & ~n12355;
  assign n12357 = ~n11869 & n12355;
  assign n12358 = ~n12356 & ~n12357;
  assign n12359 = ~n12353 & n12358;
  assign n12360 = ~n12351 & ~n12359;
  assign n12361 = po19  & ~n12360;
  assign n12362 = ~n11872 & ~n11874;
  assign n12363 = po13  & n12362;
  assign n12364 = n11879 & ~n12363;
  assign n12365 = ~n11879 & n12363;
  assign n12366 = ~n12364 & ~n12365;
  assign n12367 = ~po19  & n12360;
  assign n12368 = ~n12366 & ~n12367;
  assign n12369 = ~n12361 & ~n12368;
  assign n12370 = po20  & ~n12369;
  assign n12371 = ~po20  & ~n12361;
  assign n12372 = ~n12368 & n12371;
  assign n12373 = ~n11882 & ~n11883;
  assign n12374 = po13  & n12373;
  assign n12375 = n11888 & n12374;
  assign n12376 = ~n11888 & ~n12374;
  assign n12377 = ~n12375 & ~n12376;
  assign n12378 = ~n12372 & n12377;
  assign n12379 = ~n12370 & ~n12378;
  assign n12380 = po21  & ~n12379;
  assign n12381 = ~n11891 & ~n11893;
  assign n12382 = po13  & n12381;
  assign n12383 = n11898 & ~n12382;
  assign n12384 = ~n11898 & n12382;
  assign n12385 = ~n12383 & ~n12384;
  assign n12386 = ~po21  & n12379;
  assign n12387 = ~n12385 & ~n12386;
  assign n12388 = ~n12380 & ~n12387;
  assign n12389 = po22  & ~n12388;
  assign n12390 = ~po22  & ~n12380;
  assign n12391 = ~n12387 & n12390;
  assign n12392 = ~n11901 & ~n11902;
  assign n12393 = po13  & n12392;
  assign n12394 = ~n11907 & ~n12393;
  assign n12395 = n11907 & n12393;
  assign n12396 = ~n12394 & ~n12395;
  assign n12397 = ~n12391 & n12396;
  assign n12398 = ~n12389 & ~n12397;
  assign n12399 = po23  & ~n12398;
  assign n12400 = ~n11910 & ~n11912;
  assign n12401 = po13  & n12400;
  assign n12402 = n11917 & ~n12401;
  assign n12403 = ~n11917 & n12401;
  assign n12404 = ~n12402 & ~n12403;
  assign n12405 = ~po23  & n12398;
  assign n12406 = ~n12404 & ~n12405;
  assign n12407 = ~n12399 & ~n12406;
  assign n12408 = po24  & ~n12407;
  assign n12409 = ~n11920 & ~n11921;
  assign n12410 = po13  & n12409;
  assign n12411 = n11926 & ~n12410;
  assign n12412 = ~n11926 & n12410;
  assign n12413 = ~n12411 & ~n12412;
  assign n12414 = ~po24  & ~n12399;
  assign n12415 = ~n12406 & n12414;
  assign n12416 = ~n12413 & ~n12415;
  assign n12417 = ~n12408 & ~n12416;
  assign n12418 = po25  & ~n12417;
  assign n12419 = ~n11929 & ~n11931;
  assign n12420 = po13  & n12419;
  assign n12421 = n11936 & ~n12420;
  assign n12422 = ~n11936 & n12420;
  assign n12423 = ~n12421 & ~n12422;
  assign n12424 = ~po25  & n12417;
  assign n12425 = ~n12423 & ~n12424;
  assign n12426 = ~n12418 & ~n12425;
  assign n12427 = po26  & ~n12426;
  assign n12428 = ~po26  & ~n12418;
  assign n12429 = ~n12425 & n12428;
  assign n12430 = ~n11939 & po13 ;
  assign n12431 = ~n11945 & n12430;
  assign n12432 = n11944 & ~n12431;
  assign n12433 = n11946 & n12430;
  assign n12434 = ~n12432 & ~n12433;
  assign n12435 = ~n12429 & n12434;
  assign n12436 = ~n12427 & ~n12435;
  assign n12437 = po27  & ~n12436;
  assign n12438 = ~n11948 & ~n11950;
  assign n12439 = po13  & n12438;
  assign n12440 = n11955 & ~n12439;
  assign n12441 = ~n11955 & n12439;
  assign n12442 = ~n12440 & ~n12441;
  assign n12443 = ~po27  & n12436;
  assign n12444 = ~n12442 & ~n12443;
  assign n12445 = ~n12437 & ~n12444;
  assign n12446 = po28  & ~n12445;
  assign n12447 = ~n11958 & ~n11959;
  assign n12448 = po13  & n12447;
  assign n12449 = n11964 & ~n12448;
  assign n12450 = ~n11964 & n12448;
  assign n12451 = ~n12449 & ~n12450;
  assign n12452 = ~po28  & ~n12437;
  assign n12453 = ~n12444 & n12452;
  assign n12454 = ~n12451 & ~n12453;
  assign n12455 = ~n12446 & ~n12454;
  assign n12456 = po29  & ~n12455;
  assign n12457 = ~n11967 & ~n11969;
  assign n12458 = po13  & n12457;
  assign n12459 = n11974 & ~n12458;
  assign n12460 = ~n11974 & n12458;
  assign n12461 = ~n12459 & ~n12460;
  assign n12462 = ~po29  & n12455;
  assign n12463 = ~n12461 & ~n12462;
  assign n12464 = ~n12456 & ~n12463;
  assign n12465 = po30  & ~n12464;
  assign n12466 = ~po30  & ~n12456;
  assign n12467 = ~n12463 & n12466;
  assign n12468 = ~n11977 & po13 ;
  assign n12469 = ~n11983 & n12468;
  assign n12470 = n11982 & ~n12469;
  assign n12471 = n11984 & n12468;
  assign n12472 = ~n12470 & ~n12471;
  assign n12473 = ~n12467 & n12472;
  assign n12474 = ~n12465 & ~n12473;
  assign n12475 = po31  & ~n12474;
  assign n12476 = ~n11986 & ~n11988;
  assign n12477 = po13  & n12476;
  assign n12478 = n11993 & ~n12477;
  assign n12479 = ~n11993 & n12477;
  assign n12480 = ~n12478 & ~n12479;
  assign n12481 = ~po31  & n12474;
  assign n12482 = ~n12480 & ~n12481;
  assign n12483 = ~n12475 & ~n12482;
  assign n12484 = po32  & ~n12483;
  assign n12485 = ~n11996 & ~n11997;
  assign n12486 = po13  & n12485;
  assign n12487 = n12002 & ~n12486;
  assign n12488 = ~n12002 & n12486;
  assign n12489 = ~n12487 & ~n12488;
  assign n12490 = ~po32  & ~n12475;
  assign n12491 = ~n12482 & n12490;
  assign n12492 = ~n12489 & ~n12491;
  assign n12493 = ~n12484 & ~n12492;
  assign n12494 = po33  & ~n12493;
  assign n12495 = ~n12005 & ~n12007;
  assign n12496 = po13  & n12495;
  assign n12497 = n12012 & ~n12496;
  assign n12498 = ~n12012 & n12496;
  assign n12499 = ~n12497 & ~n12498;
  assign n12500 = ~po33  & n12493;
  assign n12501 = ~n12499 & ~n12500;
  assign n12502 = ~n12494 & ~n12501;
  assign n12503 = po34  & ~n12502;
  assign n12504 = ~po34  & ~n12494;
  assign n12505 = ~n12501 & n12504;
  assign n12506 = ~n12015 & po13 ;
  assign n12507 = ~n12021 & n12506;
  assign n12508 = n12020 & ~n12507;
  assign n12509 = n12022 & n12506;
  assign n12510 = ~n12508 & ~n12509;
  assign n12511 = ~n12505 & n12510;
  assign n12512 = ~n12503 & ~n12511;
  assign n12513 = po35  & ~n12512;
  assign n12514 = ~n12024 & ~n12026;
  assign n12515 = po13  & n12514;
  assign n12516 = n12031 & ~n12515;
  assign n12517 = ~n12031 & n12515;
  assign n12518 = ~n12516 & ~n12517;
  assign n12519 = ~po35  & n12512;
  assign n12520 = ~n12518 & ~n12519;
  assign n12521 = ~n12513 & ~n12520;
  assign n12522 = po36  & ~n12521;
  assign n12523 = ~n12034 & ~n12035;
  assign n12524 = po13  & n12523;
  assign n12525 = n12040 & ~n12524;
  assign n12526 = ~n12040 & n12524;
  assign n12527 = ~n12525 & ~n12526;
  assign n12528 = ~po36  & ~n12513;
  assign n12529 = ~n12520 & n12528;
  assign n12530 = ~n12527 & ~n12529;
  assign n12531 = ~n12522 & ~n12530;
  assign n12532 = po37  & ~n12531;
  assign n12533 = ~n12043 & ~n12045;
  assign n12534 = po13  & n12533;
  assign n12535 = n12050 & ~n12534;
  assign n12536 = ~n12050 & n12534;
  assign n12537 = ~n12535 & ~n12536;
  assign n12538 = ~po37  & n12531;
  assign n12539 = ~n12537 & ~n12538;
  assign n12540 = ~n12532 & ~n12539;
  assign n12541 = po38  & ~n12540;
  assign n12542 = ~po38  & ~n12532;
  assign n12543 = ~n12539 & n12542;
  assign n12544 = ~n12053 & po13 ;
  assign n12545 = ~n12059 & n12544;
  assign n12546 = n12058 & ~n12545;
  assign n12547 = n12060 & n12544;
  assign n12548 = ~n12546 & ~n12547;
  assign n12549 = ~n12543 & n12548;
  assign n12550 = ~n12541 & ~n12549;
  assign n12551 = po39  & ~n12550;
  assign n12552 = ~n12062 & ~n12064;
  assign n12553 = po13  & n12552;
  assign n12554 = n12069 & ~n12553;
  assign n12555 = ~n12069 & n12553;
  assign n12556 = ~n12554 & ~n12555;
  assign n12557 = ~po39  & n12550;
  assign n12558 = ~n12556 & ~n12557;
  assign n12559 = ~n12551 & ~n12558;
  assign n12560 = po40  & ~n12559;
  assign n12561 = ~n12072 & ~n12073;
  assign n12562 = po13  & n12561;
  assign n12563 = n12078 & ~n12562;
  assign n12564 = ~n12078 & n12562;
  assign n12565 = ~n12563 & ~n12564;
  assign n12566 = ~po40  & ~n12551;
  assign n12567 = ~n12558 & n12566;
  assign n12568 = ~n12565 & ~n12567;
  assign n12569 = ~n12560 & ~n12568;
  assign n12570 = po41  & ~n12569;
  assign n12571 = ~n12081 & ~n12083;
  assign n12572 = po13  & n12571;
  assign n12573 = n12088 & ~n12572;
  assign n12574 = ~n12088 & n12572;
  assign n12575 = ~n12573 & ~n12574;
  assign n12576 = ~po41  & n12569;
  assign n12577 = ~n12575 & ~n12576;
  assign n12578 = ~n12570 & ~n12577;
  assign n12579 = po42  & ~n12578;
  assign n12580 = ~po42  & ~n12570;
  assign n12581 = ~n12577 & n12580;
  assign n12582 = ~n12091 & po13 ;
  assign n12583 = ~n12097 & n12582;
  assign n12584 = n12096 & ~n12583;
  assign n12585 = n12098 & n12582;
  assign n12586 = ~n12584 & ~n12585;
  assign n12587 = ~n12581 & n12586;
  assign n12588 = ~n12579 & ~n12587;
  assign n12589 = po43  & ~n12588;
  assign n12590 = ~n12100 & ~n12102;
  assign n12591 = po13  & n12590;
  assign n12592 = n12107 & ~n12591;
  assign n12593 = ~n12107 & n12591;
  assign n12594 = ~n12592 & ~n12593;
  assign n12595 = ~po43  & n12588;
  assign n12596 = ~n12594 & ~n12595;
  assign n12597 = ~n12589 & ~n12596;
  assign n12598 = po44  & ~n12597;
  assign n12599 = ~n12110 & ~n12111;
  assign n12600 = po13  & n12599;
  assign n12601 = n12116 & ~n12600;
  assign n12602 = ~n12116 & n12600;
  assign n12603 = ~n12601 & ~n12602;
  assign n12604 = ~po44  & ~n12589;
  assign n12605 = ~n12596 & n12604;
  assign n12606 = ~n12603 & ~n12605;
  assign n12607 = ~n12598 & ~n12606;
  assign n12608 = po45  & ~n12607;
  assign n12609 = ~n12119 & ~n12121;
  assign n12610 = po13  & n12609;
  assign n12611 = n12126 & ~n12610;
  assign n12612 = ~n12126 & n12610;
  assign n12613 = ~n12611 & ~n12612;
  assign n12614 = ~po45  & n12607;
  assign n12615 = ~n12613 & ~n12614;
  assign n12616 = ~n12608 & ~n12615;
  assign n12617 = po46  & ~n12616;
  assign n12618 = ~po46  & ~n12608;
  assign n12619 = ~n12615 & n12618;
  assign n12620 = ~n12129 & po13 ;
  assign n12621 = ~n12135 & n12620;
  assign n12622 = n12134 & ~n12621;
  assign n12623 = n12136 & n12620;
  assign n12624 = ~n12622 & ~n12623;
  assign n12625 = ~n12619 & n12624;
  assign n12626 = ~n12617 & ~n12625;
  assign n12627 = po47  & ~n12626;
  assign n12628 = ~n12138 & ~n12140;
  assign n12629 = po13  & n12628;
  assign n12630 = n12145 & ~n12629;
  assign n12631 = ~n12145 & n12629;
  assign n12632 = ~n12630 & ~n12631;
  assign n12633 = ~po47  & n12626;
  assign n12634 = ~n12632 & ~n12633;
  assign n12635 = ~n12627 & ~n12634;
  assign n12636 = po48  & ~n12635;
  assign n12637 = ~n12148 & ~n12149;
  assign n12638 = po13  & n12637;
  assign n12639 = n12154 & ~n12638;
  assign n12640 = ~n12154 & n12638;
  assign n12641 = ~n12639 & ~n12640;
  assign n12642 = ~po48  & ~n12627;
  assign n12643 = ~n12634 & n12642;
  assign n12644 = ~n12641 & ~n12643;
  assign n12645 = ~n12636 & ~n12644;
  assign n12646 = ~po49  & n12645;
  assign n12647 = ~n12157 & po13 ;
  assign n12648 = ~n12164 & n12647;
  assign n12649 = n12162 & ~n12648;
  assign n12650 = n12165 & n12647;
  assign n12651 = ~n12649 & ~n12650;
  assign n12652 = ~n12646 & n12651;
  assign n12653 = po49  & ~n12645;
  assign n12654 = ~n12652 & ~n12653;
  assign n12655 = po50  & ~n12654;
  assign n12656 = ~po50  & ~n12653;
  assign n12657 = ~n12652 & n12656;
  assign n12658 = ~n12167 & ~n12169;
  assign n12659 = po13  & n12658;
  assign n12660 = n11840 & n12659;
  assign n12661 = ~n11840 & ~n12659;
  assign n12662 = ~n12660 & ~n12661;
  assign n12663 = ~n12657 & ~n12662;
  assign n12664 = ~n12655 & ~n12663;
  assign n12665 = ~po51  & n12664;
  assign n12666 = po51  & ~n12664;
  assign n12667 = ~n12310 & ~n12665;
  assign n12668 = ~n12666 & ~n12667;
  assign n12669 = po52  & ~n12668;
  assign n12670 = ~po52  & ~n12666;
  assign n12671 = ~n12667 & n12670;
  assign n12672 = ~n12176 & po13 ;
  assign n12673 = ~n12182 & n12672;
  assign n12674 = n12181 & ~n12673;
  assign n12675 = n12183 & n12672;
  assign n12676 = ~n12674 & ~n12675;
  assign n12677 = ~n12671 & n12676;
  assign n12678 = ~n12669 & ~n12677;
  assign n12679 = po53  & ~n12678;
  assign n12680 = ~n12185 & ~n12187;
  assign n12681 = po13  & n12680;
  assign n12682 = n12192 & ~n12681;
  assign n12683 = ~n12192 & n12681;
  assign n12684 = ~n12682 & ~n12683;
  assign n12685 = ~po53  & n12678;
  assign n12686 = ~n12684 & ~n12685;
  assign n12687 = ~n12679 & ~n12686;
  assign n12688 = po54  & ~n12687;
  assign n12689 = ~po54  & ~n12679;
  assign n12690 = ~n12686 & n12689;
  assign n12691 = ~n12195 & po13 ;
  assign n12692 = ~n12201 & n12691;
  assign n12693 = n12200 & ~n12692;
  assign n12694 = n12202 & n12691;
  assign n12695 = ~n12693 & ~n12694;
  assign n12696 = ~n12690 & n12695;
  assign n12697 = ~n12688 & ~n12696;
  assign n12698 = po55  & ~n12697;
  assign n12699 = ~n12204 & ~n12206;
  assign n12700 = po13  & n12699;
  assign n12701 = n12211 & ~n12700;
  assign n12702 = ~n12211 & n12700;
  assign n12703 = ~n12701 & ~n12702;
  assign n12704 = ~po55  & n12697;
  assign n12705 = ~n12703 & ~n12704;
  assign n12706 = ~n12698 & ~n12705;
  assign n12707 = po56  & ~n12706;
  assign n12708 = ~n12214 & ~n12215;
  assign n12709 = po13  & n12708;
  assign n12710 = n12220 & ~n12709;
  assign n12711 = ~n12220 & n12709;
  assign n12712 = ~n12710 & ~n12711;
  assign n12713 = ~po56  & ~n12698;
  assign n12714 = ~n12705 & n12713;
  assign n12715 = ~n12712 & ~n12714;
  assign n12716 = ~n12707 & ~n12715;
  assign n12717 = po57  & ~n12716;
  assign n12718 = ~n12223 & ~n12225;
  assign n12719 = po13  & n12718;
  assign n12720 = n12230 & ~n12719;
  assign n12721 = ~n12230 & n12719;
  assign n12722 = ~n12720 & ~n12721;
  assign n12723 = ~po57  & n12716;
  assign n12724 = ~n12722 & ~n12723;
  assign n12725 = ~n12717 & ~n12724;
  assign n12726 = po58  & ~n12725;
  assign n12727 = ~po58  & ~n12717;
  assign n12728 = ~n12724 & n12727;
  assign n12729 = ~n12233 & po13 ;
  assign n12730 = ~n12239 & n12729;
  assign n12731 = n12238 & ~n12730;
  assign n12732 = n12240 & n12729;
  assign n12733 = ~n12731 & ~n12732;
  assign n12734 = ~n12728 & n12733;
  assign n12735 = ~n12726 & ~n12734;
  assign n12736 = po59  & ~n12735;
  assign n12737 = ~n12242 & ~n12244;
  assign n12738 = po13  & n12737;
  assign n12739 = n12249 & ~n12738;
  assign n12740 = ~n12249 & n12738;
  assign n12741 = ~n12739 & ~n12740;
  assign n12742 = ~po59  & n12735;
  assign n12743 = ~n12741 & ~n12742;
  assign n12744 = ~n12736 & ~n12743;
  assign n12745 = po60  & ~n12744;
  assign n12746 = ~n12252 & ~n12253;
  assign n12747 = po13  & n12746;
  assign n12748 = n12258 & ~n12747;
  assign n12749 = ~n12258 & n12747;
  assign n12750 = ~n12748 & ~n12749;
  assign n12751 = ~po60  & ~n12736;
  assign n12752 = ~n12743 & n12751;
  assign n12753 = ~n12750 & ~n12752;
  assign n12754 = ~n12745 & ~n12753;
  assign n12755 = po61  & ~n12754;
  assign n12756 = ~n12261 & ~n12263;
  assign n12757 = po13  & n12756;
  assign n12758 = n12268 & ~n12757;
  assign n12759 = ~n12268 & n12757;
  assign n12760 = ~n12758 & ~n12759;
  assign n12761 = ~po61  & n12754;
  assign n12762 = ~n12760 & ~n12761;
  assign n12763 = ~n12755 & ~n12762;
  assign n12764 = po62  & ~n12763;
  assign n12765 = ~po62  & ~n12755;
  assign n12766 = ~n12762 & n12765;
  assign n12767 = ~n12271 & po13 ;
  assign n12768 = ~n12277 & n12767;
  assign n12769 = n12276 & ~n12768;
  assign n12770 = n12278 & n12767;
  assign n12771 = ~n12769 & ~n12770;
  assign n12772 = ~n12766 & n12771;
  assign n12773 = ~n12764 & ~n12772;
  assign n12774 = n12298 & po13 ;
  assign n12775 = ~n12289 & n12774;
  assign n12776 = ~n12280 & ~n12282;
  assign n12777 = po13  & n12776;
  assign n12778 = n12287 & ~n12777;
  assign n12779 = ~n12287 & n12777;
  assign n12780 = ~n12778 & ~n12779;
  assign n12781 = ~n12302 & ~n12775;
  assign n12782 = ~n12780 & n12781;
  assign n12783 = ~n12773 & n12782;
  assign n12784 = ~po63  & ~n12783;
  assign n12785 = n12773 & n12780;
  assign n12786 = n12289 & ~n12774;
  assign n12787 = ~n12289 & n12298;
  assign n12788 = po63  & ~n12787;
  assign n12789 = ~n12786 & n12788;
  assign n12790 = ~n12785 & ~n12789;
  assign po12  = n12784 | ~n12790;
  assign n12792 = ~n12666 & po12 ;
  assign n12793 = ~n12665 & n12792;
  assign n12794 = n12310 & ~n12793;
  assign n12795 = n12667 & n12792;
  assign n12796 = ~n12794 & ~n12795;
  assign n12797 = ~n12655 & ~n12657;
  assign n12798 = po12  & n12797;
  assign n12799 = ~n12662 & ~n12798;
  assign n12800 = n12662 & n12798;
  assign n12801 = ~n12799 & ~n12800;
  assign n12802 = pi24  & po12 ;
  assign n12803 = ~pi22  & ~pi23 ;
  assign n12804 = ~pi24  & n12803;
  assign n12805 = ~n12802 & ~n12804;
  assign n12806 = po13  & ~n12805;
  assign n12807 = ~pi24  & po12 ;
  assign n12808 = pi25  & ~n12807;
  assign n12809 = ~pi25  & n12807;
  assign n12810 = ~n12808 & ~n12809;
  assign n12811 = ~po13  & n12805;
  assign n12812 = n12810 & ~n12811;
  assign n12813 = ~n12806 & ~n12812;
  assign n12814 = po14  & ~n12813;
  assign n12815 = ~po14  & ~n12806;
  assign n12816 = ~n12812 & n12815;
  assign n12817 = po13  & ~po12 ;
  assign n12818 = ~n12809 & ~n12817;
  assign n12819 = pi26  & ~n12818;
  assign n12820 = ~pi26  & n12818;
  assign n12821 = ~n12819 & ~n12820;
  assign n12822 = ~n12816 & ~n12821;
  assign n12823 = ~n12814 & ~n12822;
  assign n12824 = po15  & ~n12823;
  assign n12825 = ~po15  & n12823;
  assign n12826 = ~n12315 & ~n12316;
  assign n12827 = po12  & n12826;
  assign n12828 = n12320 & ~n12827;
  assign n12829 = ~n12320 & n12827;
  assign n12830 = ~n12828 & ~n12829;
  assign n12831 = ~n12825 & ~n12830;
  assign n12832 = ~n12824 & ~n12831;
  assign n12833 = po16  & ~n12832;
  assign n12834 = ~po16  & ~n12824;
  assign n12835 = ~n12831 & n12834;
  assign n12836 = ~n12323 & po12 ;
  assign n12837 = ~n12329 & n12836;
  assign n12838 = n12328 & ~n12837;
  assign n12839 = n12330 & n12836;
  assign n12840 = ~n12838 & ~n12839;
  assign n12841 = ~n12835 & n12840;
  assign n12842 = ~n12833 & ~n12841;
  assign n12843 = po17  & ~n12842;
  assign n12844 = ~po17  & n12842;
  assign n12845 = ~n12332 & ~n12334;
  assign n12846 = po12  & n12845;
  assign n12847 = n12339 & ~n12846;
  assign n12848 = ~n12339 & n12846;
  assign n12849 = ~n12847 & ~n12848;
  assign n12850 = ~n12844 & n12849;
  assign n12851 = ~n12843 & ~n12850;
  assign n12852 = po18  & ~n12851;
  assign n12853 = ~po18  & ~n12843;
  assign n12854 = ~n12850 & n12853;
  assign n12855 = ~n12342 & po12 ;
  assign n12856 = ~n12348 & n12855;
  assign n12857 = n12347 & ~n12856;
  assign n12858 = n12349 & n12855;
  assign n12859 = ~n12857 & ~n12858;
  assign n12860 = ~n12854 & n12859;
  assign n12861 = ~n12852 & ~n12860;
  assign n12862 = po19  & ~n12861;
  assign n12863 = ~po19  & n12861;
  assign n12864 = ~n12351 & ~n12353;
  assign n12865 = po12  & n12864;
  assign n12866 = n12358 & n12865;
  assign n12867 = ~n12358 & ~n12865;
  assign n12868 = ~n12866 & ~n12867;
  assign n12869 = ~n12863 & n12868;
  assign n12870 = ~n12862 & ~n12869;
  assign n12871 = po20  & ~n12870;
  assign n12872 = ~po20  & ~n12862;
  assign n12873 = ~n12869 & n12872;
  assign n12874 = ~n12361 & po12 ;
  assign n12875 = ~n12367 & n12874;
  assign n12876 = n12366 & ~n12875;
  assign n12877 = n12368 & n12874;
  assign n12878 = ~n12876 & ~n12877;
  assign n12879 = ~n12873 & n12878;
  assign n12880 = ~n12871 & ~n12879;
  assign n12881 = po21  & ~n12880;
  assign n12882 = ~po21  & n12880;
  assign n12883 = ~n12370 & ~n12372;
  assign n12884 = po12  & n12883;
  assign n12885 = ~n12377 & ~n12884;
  assign n12886 = n12377 & n12884;
  assign n12887 = ~n12885 & ~n12886;
  assign n12888 = ~n12882 & n12887;
  assign n12889 = ~n12881 & ~n12888;
  assign n12890 = po22  & ~n12889;
  assign n12891 = ~po22  & ~n12881;
  assign n12892 = ~n12888 & n12891;
  assign n12893 = ~n12380 & po12 ;
  assign n12894 = ~n12386 & n12893;
  assign n12895 = n12385 & ~n12894;
  assign n12896 = n12387 & n12893;
  assign n12897 = ~n12895 & ~n12896;
  assign n12898 = ~n12892 & n12897;
  assign n12899 = ~n12890 & ~n12898;
  assign n12900 = po23  & ~n12899;
  assign n12901 = ~n12389 & ~n12391;
  assign n12902 = po12  & n12901;
  assign n12903 = n12396 & ~n12902;
  assign n12904 = ~n12396 & n12902;
  assign n12905 = ~n12903 & ~n12904;
  assign n12906 = ~po23  & n12899;
  assign n12907 = ~n12905 & ~n12906;
  assign n12908 = ~n12900 & ~n12907;
  assign n12909 = po24  & ~n12908;
  assign n12910 = ~po24  & ~n12900;
  assign n12911 = ~n12907 & n12910;
  assign n12912 = ~n12399 & po12 ;
  assign n12913 = ~n12405 & n12912;
  assign n12914 = n12404 & ~n12913;
  assign n12915 = n12406 & n12912;
  assign n12916 = ~n12914 & ~n12915;
  assign n12917 = ~n12911 & n12916;
  assign n12918 = ~n12909 & ~n12917;
  assign n12919 = po25  & ~n12918;
  assign n12920 = ~po25  & n12918;
  assign n12921 = ~n12408 & po12 ;
  assign n12922 = ~n12415 & n12921;
  assign n12923 = n12413 & ~n12922;
  assign n12924 = n12416 & n12921;
  assign n12925 = ~n12923 & ~n12924;
  assign n12926 = ~n12920 & n12925;
  assign n12927 = ~n12919 & ~n12926;
  assign n12928 = po26  & ~n12927;
  assign n12929 = ~po26  & ~n12919;
  assign n12930 = ~n12926 & n12929;
  assign n12931 = ~n12418 & po12 ;
  assign n12932 = ~n12424 & n12931;
  assign n12933 = n12423 & ~n12932;
  assign n12934 = n12425 & n12931;
  assign n12935 = ~n12933 & ~n12934;
  assign n12936 = ~n12930 & n12935;
  assign n12937 = ~n12928 & ~n12936;
  assign n12938 = po27  & ~n12937;
  assign n12939 = ~n12427 & ~n12429;
  assign n12940 = po12  & n12939;
  assign n12941 = n12434 & ~n12940;
  assign n12942 = ~n12434 & n12940;
  assign n12943 = ~n12941 & ~n12942;
  assign n12944 = ~po27  & n12937;
  assign n12945 = ~n12943 & ~n12944;
  assign n12946 = ~n12938 & ~n12945;
  assign n12947 = po28  & ~n12946;
  assign n12948 = ~po28  & ~n12938;
  assign n12949 = ~n12945 & n12948;
  assign n12950 = ~n12437 & po12 ;
  assign n12951 = ~n12443 & n12950;
  assign n12952 = n12442 & ~n12951;
  assign n12953 = n12444 & n12950;
  assign n12954 = ~n12952 & ~n12953;
  assign n12955 = ~n12949 & n12954;
  assign n12956 = ~n12947 & ~n12955;
  assign n12957 = po29  & ~n12956;
  assign n12958 = ~po29  & n12956;
  assign n12959 = ~n12446 & po12 ;
  assign n12960 = ~n12453 & n12959;
  assign n12961 = n12451 & ~n12960;
  assign n12962 = n12454 & n12959;
  assign n12963 = ~n12961 & ~n12962;
  assign n12964 = ~n12958 & n12963;
  assign n12965 = ~n12957 & ~n12964;
  assign n12966 = po30  & ~n12965;
  assign n12967 = ~po30  & ~n12957;
  assign n12968 = ~n12964 & n12967;
  assign n12969 = ~n12456 & po12 ;
  assign n12970 = ~n12462 & n12969;
  assign n12971 = n12461 & ~n12970;
  assign n12972 = n12463 & n12969;
  assign n12973 = ~n12971 & ~n12972;
  assign n12974 = ~n12968 & n12973;
  assign n12975 = ~n12966 & ~n12974;
  assign n12976 = po31  & ~n12975;
  assign n12977 = ~n12465 & ~n12467;
  assign n12978 = po12  & n12977;
  assign n12979 = n12472 & ~n12978;
  assign n12980 = ~n12472 & n12978;
  assign n12981 = ~n12979 & ~n12980;
  assign n12982 = ~po31  & n12975;
  assign n12983 = ~n12981 & ~n12982;
  assign n12984 = ~n12976 & ~n12983;
  assign n12985 = po32  & ~n12984;
  assign n12986 = ~po32  & ~n12976;
  assign n12987 = ~n12983 & n12986;
  assign n12988 = ~n12475 & po12 ;
  assign n12989 = ~n12481 & n12988;
  assign n12990 = n12480 & ~n12989;
  assign n12991 = n12482 & n12988;
  assign n12992 = ~n12990 & ~n12991;
  assign n12993 = ~n12987 & n12992;
  assign n12994 = ~n12985 & ~n12993;
  assign n12995 = po33  & ~n12994;
  assign n12996 = ~po33  & n12994;
  assign n12997 = ~n12484 & po12 ;
  assign n12998 = ~n12491 & n12997;
  assign n12999 = n12489 & ~n12998;
  assign n13000 = n12492 & n12997;
  assign n13001 = ~n12999 & ~n13000;
  assign n13002 = ~n12996 & n13001;
  assign n13003 = ~n12995 & ~n13002;
  assign n13004 = po34  & ~n13003;
  assign n13005 = ~po34  & ~n12995;
  assign n13006 = ~n13002 & n13005;
  assign n13007 = ~n12494 & po12 ;
  assign n13008 = ~n12500 & n13007;
  assign n13009 = n12499 & ~n13008;
  assign n13010 = n12501 & n13007;
  assign n13011 = ~n13009 & ~n13010;
  assign n13012 = ~n13006 & n13011;
  assign n13013 = ~n13004 & ~n13012;
  assign n13014 = po35  & ~n13013;
  assign n13015 = ~n12503 & ~n12505;
  assign n13016 = po12  & n13015;
  assign n13017 = n12510 & ~n13016;
  assign n13018 = ~n12510 & n13016;
  assign n13019 = ~n13017 & ~n13018;
  assign n13020 = ~po35  & n13013;
  assign n13021 = ~n13019 & ~n13020;
  assign n13022 = ~n13014 & ~n13021;
  assign n13023 = po36  & ~n13022;
  assign n13024 = ~po36  & ~n13014;
  assign n13025 = ~n13021 & n13024;
  assign n13026 = ~n12513 & po12 ;
  assign n13027 = ~n12519 & n13026;
  assign n13028 = n12518 & ~n13027;
  assign n13029 = n12520 & n13026;
  assign n13030 = ~n13028 & ~n13029;
  assign n13031 = ~n13025 & n13030;
  assign n13032 = ~n13023 & ~n13031;
  assign n13033 = po37  & ~n13032;
  assign n13034 = ~po37  & n13032;
  assign n13035 = ~n12522 & po12 ;
  assign n13036 = ~n12529 & n13035;
  assign n13037 = n12527 & ~n13036;
  assign n13038 = n12530 & n13035;
  assign n13039 = ~n13037 & ~n13038;
  assign n13040 = ~n13034 & n13039;
  assign n13041 = ~n13033 & ~n13040;
  assign n13042 = po38  & ~n13041;
  assign n13043 = ~po38  & ~n13033;
  assign n13044 = ~n13040 & n13043;
  assign n13045 = ~n12532 & po12 ;
  assign n13046 = ~n12538 & n13045;
  assign n13047 = n12537 & ~n13046;
  assign n13048 = n12539 & n13045;
  assign n13049 = ~n13047 & ~n13048;
  assign n13050 = ~n13044 & n13049;
  assign n13051 = ~n13042 & ~n13050;
  assign n13052 = po39  & ~n13051;
  assign n13053 = ~n12541 & ~n12543;
  assign n13054 = po12  & n13053;
  assign n13055 = n12548 & ~n13054;
  assign n13056 = ~n12548 & n13054;
  assign n13057 = ~n13055 & ~n13056;
  assign n13058 = ~po39  & n13051;
  assign n13059 = ~n13057 & ~n13058;
  assign n13060 = ~n13052 & ~n13059;
  assign n13061 = po40  & ~n13060;
  assign n13062 = ~po40  & ~n13052;
  assign n13063 = ~n13059 & n13062;
  assign n13064 = ~n12551 & po12 ;
  assign n13065 = ~n12557 & n13064;
  assign n13066 = n12556 & ~n13065;
  assign n13067 = n12558 & n13064;
  assign n13068 = ~n13066 & ~n13067;
  assign n13069 = ~n13063 & n13068;
  assign n13070 = ~n13061 & ~n13069;
  assign n13071 = po41  & ~n13070;
  assign n13072 = ~po41  & n13070;
  assign n13073 = ~n12560 & po12 ;
  assign n13074 = ~n12567 & n13073;
  assign n13075 = n12565 & ~n13074;
  assign n13076 = n12568 & n13073;
  assign n13077 = ~n13075 & ~n13076;
  assign n13078 = ~n13072 & n13077;
  assign n13079 = ~n13071 & ~n13078;
  assign n13080 = po42  & ~n13079;
  assign n13081 = ~po42  & ~n13071;
  assign n13082 = ~n13078 & n13081;
  assign n13083 = ~n12570 & po12 ;
  assign n13084 = ~n12576 & n13083;
  assign n13085 = n12575 & ~n13084;
  assign n13086 = n12577 & n13083;
  assign n13087 = ~n13085 & ~n13086;
  assign n13088 = ~n13082 & n13087;
  assign n13089 = ~n13080 & ~n13088;
  assign n13090 = po43  & ~n13089;
  assign n13091 = ~n12579 & ~n12581;
  assign n13092 = po12  & n13091;
  assign n13093 = n12586 & ~n13092;
  assign n13094 = ~n12586 & n13092;
  assign n13095 = ~n13093 & ~n13094;
  assign n13096 = ~po43  & n13089;
  assign n13097 = ~n13095 & ~n13096;
  assign n13098 = ~n13090 & ~n13097;
  assign n13099 = po44  & ~n13098;
  assign n13100 = ~po44  & ~n13090;
  assign n13101 = ~n13097 & n13100;
  assign n13102 = ~n12589 & po12 ;
  assign n13103 = ~n12595 & n13102;
  assign n13104 = n12594 & ~n13103;
  assign n13105 = n12596 & n13102;
  assign n13106 = ~n13104 & ~n13105;
  assign n13107 = ~n13101 & n13106;
  assign n13108 = ~n13099 & ~n13107;
  assign n13109 = po45  & ~n13108;
  assign n13110 = ~po45  & n13108;
  assign n13111 = ~n12598 & po12 ;
  assign n13112 = ~n12605 & n13111;
  assign n13113 = n12603 & ~n13112;
  assign n13114 = n12606 & n13111;
  assign n13115 = ~n13113 & ~n13114;
  assign n13116 = ~n13110 & n13115;
  assign n13117 = ~n13109 & ~n13116;
  assign n13118 = po46  & ~n13117;
  assign n13119 = ~po46  & ~n13109;
  assign n13120 = ~n13116 & n13119;
  assign n13121 = ~n12608 & po12 ;
  assign n13122 = ~n12614 & n13121;
  assign n13123 = n12613 & ~n13122;
  assign n13124 = n12615 & n13121;
  assign n13125 = ~n13123 & ~n13124;
  assign n13126 = ~n13120 & n13125;
  assign n13127 = ~n13118 & ~n13126;
  assign n13128 = po47  & ~n13127;
  assign n13129 = ~n12617 & ~n12619;
  assign n13130 = po12  & n13129;
  assign n13131 = n12624 & ~n13130;
  assign n13132 = ~n12624 & n13130;
  assign n13133 = ~n13131 & ~n13132;
  assign n13134 = ~po47  & n13127;
  assign n13135 = ~n13133 & ~n13134;
  assign n13136 = ~n13128 & ~n13135;
  assign n13137 = po48  & ~n13136;
  assign n13138 = ~po48  & ~n13128;
  assign n13139 = ~n13135 & n13138;
  assign n13140 = ~n12627 & po12 ;
  assign n13141 = ~n12633 & n13140;
  assign n13142 = n12632 & ~n13141;
  assign n13143 = n12634 & n13140;
  assign n13144 = ~n13142 & ~n13143;
  assign n13145 = ~n13139 & n13144;
  assign n13146 = ~n13137 & ~n13145;
  assign n13147 = po49  & ~n13146;
  assign n13148 = ~po49  & n13146;
  assign n13149 = ~n12636 & po12 ;
  assign n13150 = ~n12643 & n13149;
  assign n13151 = n12641 & ~n13150;
  assign n13152 = n12644 & n13149;
  assign n13153 = ~n13151 & ~n13152;
  assign n13154 = ~n13148 & n13153;
  assign n13155 = ~n13147 & ~n13154;
  assign n13156 = po50  & ~n13155;
  assign n13157 = ~n12646 & ~n12653;
  assign n13158 = po12  & n13157;
  assign n13159 = n12651 & ~n13158;
  assign n13160 = ~n12651 & n13158;
  assign n13161 = ~n13159 & ~n13160;
  assign n13162 = ~po50  & ~n13147;
  assign n13163 = ~n13154 & n13162;
  assign n13164 = ~n13161 & ~n13163;
  assign n13165 = ~n13156 & ~n13164;
  assign n13166 = ~po51  & n13165;
  assign n13167 = ~n12801 & ~n13166;
  assign n13168 = po51  & ~n13165;
  assign n13169 = ~po52  & ~n13168;
  assign n13170 = ~n13167 & n13169;
  assign n13171 = ~n13167 & ~n13168;
  assign n13172 = po52  & ~n13171;
  assign n13173 = n12796 & ~n13170;
  assign n13174 = ~n13172 & ~n13173;
  assign n13175 = po53  & ~n13174;
  assign n13176 = ~n12669 & ~n12671;
  assign n13177 = po12  & n13176;
  assign n13178 = n12676 & ~n13177;
  assign n13179 = ~n12676 & n13177;
  assign n13180 = ~n13178 & ~n13179;
  assign n13181 = ~po53  & n13174;
  assign n13182 = ~n13180 & ~n13181;
  assign n13183 = ~n13175 & ~n13182;
  assign n13184 = po54  & ~n13183;
  assign n13185 = ~po54  & ~n13175;
  assign n13186 = ~n13182 & n13185;
  assign n13187 = ~n12679 & po12 ;
  assign n13188 = ~n12685 & n13187;
  assign n13189 = n12684 & ~n13188;
  assign n13190 = n12686 & n13187;
  assign n13191 = ~n13189 & ~n13190;
  assign n13192 = ~n13186 & n13191;
  assign n13193 = ~n13184 & ~n13192;
  assign n13194 = po55  & ~n13193;
  assign n13195 = ~n12688 & ~n12690;
  assign n13196 = po12  & n13195;
  assign n13197 = n12695 & ~n13196;
  assign n13198 = ~n12695 & n13196;
  assign n13199 = ~n13197 & ~n13198;
  assign n13200 = ~po55  & n13193;
  assign n13201 = ~n13199 & ~n13200;
  assign n13202 = ~n13194 & ~n13201;
  assign n13203 = po56  & ~n13202;
  assign n13204 = ~po56  & ~n13194;
  assign n13205 = ~n13201 & n13204;
  assign n13206 = ~n12698 & po12 ;
  assign n13207 = ~n12704 & n13206;
  assign n13208 = n12703 & ~n13207;
  assign n13209 = n12705 & n13206;
  assign n13210 = ~n13208 & ~n13209;
  assign n13211 = ~n13205 & n13210;
  assign n13212 = ~n13203 & ~n13211;
  assign n13213 = po57  & ~n13212;
  assign n13214 = ~po57  & n13212;
  assign n13215 = ~n12707 & po12 ;
  assign n13216 = ~n12714 & n13215;
  assign n13217 = n12712 & ~n13216;
  assign n13218 = n12715 & n13215;
  assign n13219 = ~n13217 & ~n13218;
  assign n13220 = ~n13214 & n13219;
  assign n13221 = ~n13213 & ~n13220;
  assign n13222 = po58  & ~n13221;
  assign n13223 = ~po58  & ~n13213;
  assign n13224 = ~n13220 & n13223;
  assign n13225 = ~n12717 & po12 ;
  assign n13226 = ~n12723 & n13225;
  assign n13227 = n12722 & ~n13226;
  assign n13228 = n12724 & n13225;
  assign n13229 = ~n13227 & ~n13228;
  assign n13230 = ~n13224 & n13229;
  assign n13231 = ~n13222 & ~n13230;
  assign n13232 = po59  & ~n13231;
  assign n13233 = ~n12726 & ~n12728;
  assign n13234 = po12  & n13233;
  assign n13235 = n12733 & ~n13234;
  assign n13236 = ~n12733 & n13234;
  assign n13237 = ~n13235 & ~n13236;
  assign n13238 = ~po59  & n13231;
  assign n13239 = ~n13237 & ~n13238;
  assign n13240 = ~n13232 & ~n13239;
  assign n13241 = po60  & ~n13240;
  assign n13242 = ~po60  & ~n13232;
  assign n13243 = ~n13239 & n13242;
  assign n13244 = ~n12736 & po12 ;
  assign n13245 = ~n12742 & n13244;
  assign n13246 = n12741 & ~n13245;
  assign n13247 = n12743 & n13244;
  assign n13248 = ~n13246 & ~n13247;
  assign n13249 = ~n13243 & n13248;
  assign n13250 = ~n13241 & ~n13249;
  assign n13251 = po61  & ~n13250;
  assign n13252 = ~po61  & n13250;
  assign n13253 = ~n12745 & po12 ;
  assign n13254 = ~n12752 & n13253;
  assign n13255 = n12750 & ~n13254;
  assign n13256 = n12753 & n13253;
  assign n13257 = ~n13255 & ~n13256;
  assign n13258 = ~n13252 & n13257;
  assign n13259 = ~n13251 & ~n13258;
  assign n13260 = po62  & ~n13259;
  assign n13261 = ~po62  & ~n13251;
  assign n13262 = ~n13258 & n13261;
  assign n13263 = ~n12755 & po12 ;
  assign n13264 = ~n12761 & n13263;
  assign n13265 = n12760 & ~n13264;
  assign n13266 = n12762 & n13263;
  assign n13267 = ~n13265 & ~n13266;
  assign n13268 = ~n13262 & n13267;
  assign n13269 = ~n13260 & ~n13268;
  assign n13270 = ~n12764 & ~n12766;
  assign n13271 = po12  & n13270;
  assign n13272 = n12771 & ~n13271;
  assign n13273 = ~n12771 & n13271;
  assign n13274 = ~n13272 & ~n13273;
  assign n13275 = n12773 & po12 ;
  assign n13276 = ~n12780 & ~n13275;
  assign n13277 = ~n12785 & ~n13276;
  assign n13278 = po12  & ~n13277;
  assign n13279 = ~n13274 & ~n13278;
  assign n13280 = ~n13269 & n13279;
  assign n13281 = ~po63  & ~n13280;
  assign n13282 = n13269 & n13274;
  assign n13283 = po63  & n13277;
  assign n13284 = ~n13282 & ~n13283;
  assign po11  = n13281 | ~n13284;
  assign n13286 = ~n13170 & ~n13172;
  assign n13287 = po11  & n13286;
  assign n13288 = n12796 & ~n13287;
  assign n13289 = ~n12796 & n13287;
  assign n13290 = ~n13288 & ~n13289;
  assign n13291 = pi22  & po11 ;
  assign n13292 = ~pi20  & ~pi21 ;
  assign n13293 = ~pi22  & n13292;
  assign n13294 = ~n13291 & ~n13293;
  assign n13295 = po12  & ~n13294;
  assign n13296 = ~po12  & n13294;
  assign n13297 = ~pi22  & po11 ;
  assign n13298 = pi23  & ~n13297;
  assign n13299 = ~pi23  & n13297;
  assign n13300 = ~n13298 & ~n13299;
  assign n13301 = ~n13296 & n13300;
  assign n13302 = ~n13295 & ~n13301;
  assign n13303 = po13  & ~n13302;
  assign n13304 = po12  & ~po11 ;
  assign n13305 = ~n13299 & ~n13304;
  assign n13306 = pi24  & ~n13305;
  assign n13307 = ~pi24  & n13305;
  assign n13308 = ~n13306 & ~n13307;
  assign n13309 = ~po13  & n13302;
  assign n13310 = ~n13308 & ~n13309;
  assign n13311 = ~n13303 & ~n13310;
  assign n13312 = po14  & ~n13311;
  assign n13313 = ~po14  & ~n13303;
  assign n13314 = ~n13310 & n13313;
  assign n13315 = ~n12806 & ~n12811;
  assign n13316 = po11  & n13315;
  assign n13317 = n12810 & ~n13316;
  assign n13318 = ~n12810 & n13316;
  assign n13319 = ~n13317 & ~n13318;
  assign n13320 = ~n13314 & ~n13319;
  assign n13321 = ~n13312 & ~n13320;
  assign n13322 = po15  & ~n13321;
  assign n13323 = ~n12814 & ~n12816;
  assign n13324 = po11  & n13323;
  assign n13325 = ~n12821 & ~n13324;
  assign n13326 = n12821 & n13324;
  assign n13327 = ~n13325 & ~n13326;
  assign n13328 = ~po15  & n13321;
  assign n13329 = ~n13327 & ~n13328;
  assign n13330 = ~n13322 & ~n13329;
  assign n13331 = po16  & ~n13330;
  assign n13332 = ~po16  & ~n13322;
  assign n13333 = ~n13329 & n13332;
  assign n13334 = ~n12824 & ~n12825;
  assign n13335 = po11  & n13334;
  assign n13336 = n12830 & ~n13335;
  assign n13337 = ~n12830 & n13335;
  assign n13338 = ~n13336 & ~n13337;
  assign n13339 = ~n13333 & n13338;
  assign n13340 = ~n13331 & ~n13339;
  assign n13341 = po17  & ~n13340;
  assign n13342 = ~n12833 & ~n12835;
  assign n13343 = po11  & n13342;
  assign n13344 = n12840 & ~n13343;
  assign n13345 = ~n12840 & n13343;
  assign n13346 = ~n13344 & ~n13345;
  assign n13347 = ~po17  & n13340;
  assign n13348 = ~n13346 & ~n13347;
  assign n13349 = ~n13341 & ~n13348;
  assign n13350 = po18  & ~n13349;
  assign n13351 = ~po18  & ~n13341;
  assign n13352 = ~n13348 & n13351;
  assign n13353 = ~n12843 & ~n12844;
  assign n13354 = po11  & n13353;
  assign n13355 = n12849 & n13354;
  assign n13356 = ~n12849 & ~n13354;
  assign n13357 = ~n13355 & ~n13356;
  assign n13358 = ~n13352 & n13357;
  assign n13359 = ~n13350 & ~n13358;
  assign n13360 = po19  & ~n13359;
  assign n13361 = ~n12852 & ~n12854;
  assign n13362 = po11  & n13361;
  assign n13363 = n12859 & ~n13362;
  assign n13364 = ~n12859 & n13362;
  assign n13365 = ~n13363 & ~n13364;
  assign n13366 = ~po19  & n13359;
  assign n13367 = ~n13365 & ~n13366;
  assign n13368 = ~n13360 & ~n13367;
  assign n13369 = po20  & ~n13368;
  assign n13370 = ~po20  & ~n13360;
  assign n13371 = ~n13367 & n13370;
  assign n13372 = ~n12862 & ~n12863;
  assign n13373 = po11  & n13372;
  assign n13374 = ~n12868 & ~n13373;
  assign n13375 = n12868 & n13373;
  assign n13376 = ~n13374 & ~n13375;
  assign n13377 = ~n13371 & n13376;
  assign n13378 = ~n13369 & ~n13377;
  assign n13379 = po21  & ~n13378;
  assign n13380 = ~n12871 & ~n12873;
  assign n13381 = po11  & n13380;
  assign n13382 = n12878 & ~n13381;
  assign n13383 = ~n12878 & n13381;
  assign n13384 = ~n13382 & ~n13383;
  assign n13385 = ~po21  & n13378;
  assign n13386 = ~n13384 & ~n13385;
  assign n13387 = ~n13379 & ~n13386;
  assign n13388 = po22  & ~n13387;
  assign n13389 = ~n12881 & ~n12882;
  assign n13390 = po11  & n13389;
  assign n13391 = n12887 & ~n13390;
  assign n13392 = ~n12887 & n13390;
  assign n13393 = ~n13391 & ~n13392;
  assign n13394 = ~po22  & ~n13379;
  assign n13395 = ~n13386 & n13394;
  assign n13396 = ~n13393 & ~n13395;
  assign n13397 = ~n13388 & ~n13396;
  assign n13398 = po23  & ~n13397;
  assign n13399 = ~n12890 & ~n12892;
  assign n13400 = po11  & n13399;
  assign n13401 = n12897 & ~n13400;
  assign n13402 = ~n12897 & n13400;
  assign n13403 = ~n13401 & ~n13402;
  assign n13404 = ~po23  & n13397;
  assign n13405 = ~n13403 & ~n13404;
  assign n13406 = ~n13398 & ~n13405;
  assign n13407 = po24  & ~n13406;
  assign n13408 = ~po24  & ~n13398;
  assign n13409 = ~n13405 & n13408;
  assign n13410 = ~n12900 & po11 ;
  assign n13411 = ~n12906 & n13410;
  assign n13412 = n12905 & ~n13411;
  assign n13413 = n12907 & n13410;
  assign n13414 = ~n13412 & ~n13413;
  assign n13415 = ~n13409 & n13414;
  assign n13416 = ~n13407 & ~n13415;
  assign n13417 = po25  & ~n13416;
  assign n13418 = ~n12909 & ~n12911;
  assign n13419 = po11  & n13418;
  assign n13420 = n12916 & ~n13419;
  assign n13421 = ~n12916 & n13419;
  assign n13422 = ~n13420 & ~n13421;
  assign n13423 = ~po25  & n13416;
  assign n13424 = ~n13422 & ~n13423;
  assign n13425 = ~n13417 & ~n13424;
  assign n13426 = po26  & ~n13425;
  assign n13427 = ~n12919 & ~n12920;
  assign n13428 = po11  & n13427;
  assign n13429 = n12925 & ~n13428;
  assign n13430 = ~n12925 & n13428;
  assign n13431 = ~n13429 & ~n13430;
  assign n13432 = ~po26  & ~n13417;
  assign n13433 = ~n13424 & n13432;
  assign n13434 = ~n13431 & ~n13433;
  assign n13435 = ~n13426 & ~n13434;
  assign n13436 = po27  & ~n13435;
  assign n13437 = ~n12928 & ~n12930;
  assign n13438 = po11  & n13437;
  assign n13439 = n12935 & ~n13438;
  assign n13440 = ~n12935 & n13438;
  assign n13441 = ~n13439 & ~n13440;
  assign n13442 = ~po27  & n13435;
  assign n13443 = ~n13441 & ~n13442;
  assign n13444 = ~n13436 & ~n13443;
  assign n13445 = po28  & ~n13444;
  assign n13446 = ~po28  & ~n13436;
  assign n13447 = ~n13443 & n13446;
  assign n13448 = ~n12938 & po11 ;
  assign n13449 = ~n12944 & n13448;
  assign n13450 = n12943 & ~n13449;
  assign n13451 = n12945 & n13448;
  assign n13452 = ~n13450 & ~n13451;
  assign n13453 = ~n13447 & n13452;
  assign n13454 = ~n13445 & ~n13453;
  assign n13455 = po29  & ~n13454;
  assign n13456 = ~n12947 & ~n12949;
  assign n13457 = po11  & n13456;
  assign n13458 = n12954 & ~n13457;
  assign n13459 = ~n12954 & n13457;
  assign n13460 = ~n13458 & ~n13459;
  assign n13461 = ~po29  & n13454;
  assign n13462 = ~n13460 & ~n13461;
  assign n13463 = ~n13455 & ~n13462;
  assign n13464 = po30  & ~n13463;
  assign n13465 = ~n12957 & ~n12958;
  assign n13466 = po11  & n13465;
  assign n13467 = n12963 & ~n13466;
  assign n13468 = ~n12963 & n13466;
  assign n13469 = ~n13467 & ~n13468;
  assign n13470 = ~po30  & ~n13455;
  assign n13471 = ~n13462 & n13470;
  assign n13472 = ~n13469 & ~n13471;
  assign n13473 = ~n13464 & ~n13472;
  assign n13474 = po31  & ~n13473;
  assign n13475 = ~n12966 & ~n12968;
  assign n13476 = po11  & n13475;
  assign n13477 = n12973 & ~n13476;
  assign n13478 = ~n12973 & n13476;
  assign n13479 = ~n13477 & ~n13478;
  assign n13480 = ~po31  & n13473;
  assign n13481 = ~n13479 & ~n13480;
  assign n13482 = ~n13474 & ~n13481;
  assign n13483 = po32  & ~n13482;
  assign n13484 = ~po32  & ~n13474;
  assign n13485 = ~n13481 & n13484;
  assign n13486 = ~n12976 & po11 ;
  assign n13487 = ~n12982 & n13486;
  assign n13488 = n12981 & ~n13487;
  assign n13489 = n12983 & n13486;
  assign n13490 = ~n13488 & ~n13489;
  assign n13491 = ~n13485 & n13490;
  assign n13492 = ~n13483 & ~n13491;
  assign n13493 = po33  & ~n13492;
  assign n13494 = ~n12985 & ~n12987;
  assign n13495 = po11  & n13494;
  assign n13496 = n12992 & ~n13495;
  assign n13497 = ~n12992 & n13495;
  assign n13498 = ~n13496 & ~n13497;
  assign n13499 = ~po33  & n13492;
  assign n13500 = ~n13498 & ~n13499;
  assign n13501 = ~n13493 & ~n13500;
  assign n13502 = po34  & ~n13501;
  assign n13503 = ~n12995 & ~n12996;
  assign n13504 = po11  & n13503;
  assign n13505 = n13001 & ~n13504;
  assign n13506 = ~n13001 & n13504;
  assign n13507 = ~n13505 & ~n13506;
  assign n13508 = ~po34  & ~n13493;
  assign n13509 = ~n13500 & n13508;
  assign n13510 = ~n13507 & ~n13509;
  assign n13511 = ~n13502 & ~n13510;
  assign n13512 = po35  & ~n13511;
  assign n13513 = ~n13004 & ~n13006;
  assign n13514 = po11  & n13513;
  assign n13515 = n13011 & ~n13514;
  assign n13516 = ~n13011 & n13514;
  assign n13517 = ~n13515 & ~n13516;
  assign n13518 = ~po35  & n13511;
  assign n13519 = ~n13517 & ~n13518;
  assign n13520 = ~n13512 & ~n13519;
  assign n13521 = po36  & ~n13520;
  assign n13522 = ~po36  & ~n13512;
  assign n13523 = ~n13519 & n13522;
  assign n13524 = ~n13014 & po11 ;
  assign n13525 = ~n13020 & n13524;
  assign n13526 = n13019 & ~n13525;
  assign n13527 = n13021 & n13524;
  assign n13528 = ~n13526 & ~n13527;
  assign n13529 = ~n13523 & n13528;
  assign n13530 = ~n13521 & ~n13529;
  assign n13531 = po37  & ~n13530;
  assign n13532 = ~n13023 & ~n13025;
  assign n13533 = po11  & n13532;
  assign n13534 = n13030 & ~n13533;
  assign n13535 = ~n13030 & n13533;
  assign n13536 = ~n13534 & ~n13535;
  assign n13537 = ~po37  & n13530;
  assign n13538 = ~n13536 & ~n13537;
  assign n13539 = ~n13531 & ~n13538;
  assign n13540 = po38  & ~n13539;
  assign n13541 = ~n13033 & ~n13034;
  assign n13542 = po11  & n13541;
  assign n13543 = n13039 & ~n13542;
  assign n13544 = ~n13039 & n13542;
  assign n13545 = ~n13543 & ~n13544;
  assign n13546 = ~po38  & ~n13531;
  assign n13547 = ~n13538 & n13546;
  assign n13548 = ~n13545 & ~n13547;
  assign n13549 = ~n13540 & ~n13548;
  assign n13550 = po39  & ~n13549;
  assign n13551 = ~n13042 & ~n13044;
  assign n13552 = po11  & n13551;
  assign n13553 = n13049 & ~n13552;
  assign n13554 = ~n13049 & n13552;
  assign n13555 = ~n13553 & ~n13554;
  assign n13556 = ~po39  & n13549;
  assign n13557 = ~n13555 & ~n13556;
  assign n13558 = ~n13550 & ~n13557;
  assign n13559 = po40  & ~n13558;
  assign n13560 = ~po40  & ~n13550;
  assign n13561 = ~n13557 & n13560;
  assign n13562 = ~n13052 & po11 ;
  assign n13563 = ~n13058 & n13562;
  assign n13564 = n13057 & ~n13563;
  assign n13565 = n13059 & n13562;
  assign n13566 = ~n13564 & ~n13565;
  assign n13567 = ~n13561 & n13566;
  assign n13568 = ~n13559 & ~n13567;
  assign n13569 = po41  & ~n13568;
  assign n13570 = ~n13061 & ~n13063;
  assign n13571 = po11  & n13570;
  assign n13572 = n13068 & ~n13571;
  assign n13573 = ~n13068 & n13571;
  assign n13574 = ~n13572 & ~n13573;
  assign n13575 = ~po41  & n13568;
  assign n13576 = ~n13574 & ~n13575;
  assign n13577 = ~n13569 & ~n13576;
  assign n13578 = po42  & ~n13577;
  assign n13579 = ~n13071 & ~n13072;
  assign n13580 = po11  & n13579;
  assign n13581 = n13077 & ~n13580;
  assign n13582 = ~n13077 & n13580;
  assign n13583 = ~n13581 & ~n13582;
  assign n13584 = ~po42  & ~n13569;
  assign n13585 = ~n13576 & n13584;
  assign n13586 = ~n13583 & ~n13585;
  assign n13587 = ~n13578 & ~n13586;
  assign n13588 = po43  & ~n13587;
  assign n13589 = ~n13080 & ~n13082;
  assign n13590 = po11  & n13589;
  assign n13591 = n13087 & ~n13590;
  assign n13592 = ~n13087 & n13590;
  assign n13593 = ~n13591 & ~n13592;
  assign n13594 = ~po43  & n13587;
  assign n13595 = ~n13593 & ~n13594;
  assign n13596 = ~n13588 & ~n13595;
  assign n13597 = po44  & ~n13596;
  assign n13598 = ~po44  & ~n13588;
  assign n13599 = ~n13595 & n13598;
  assign n13600 = ~n13090 & po11 ;
  assign n13601 = ~n13096 & n13600;
  assign n13602 = n13095 & ~n13601;
  assign n13603 = n13097 & n13600;
  assign n13604 = ~n13602 & ~n13603;
  assign n13605 = ~n13599 & n13604;
  assign n13606 = ~n13597 & ~n13605;
  assign n13607 = po45  & ~n13606;
  assign n13608 = ~n13099 & ~n13101;
  assign n13609 = po11  & n13608;
  assign n13610 = n13106 & ~n13609;
  assign n13611 = ~n13106 & n13609;
  assign n13612 = ~n13610 & ~n13611;
  assign n13613 = ~po45  & n13606;
  assign n13614 = ~n13612 & ~n13613;
  assign n13615 = ~n13607 & ~n13614;
  assign n13616 = po46  & ~n13615;
  assign n13617 = ~n13109 & ~n13110;
  assign n13618 = po11  & n13617;
  assign n13619 = n13115 & ~n13618;
  assign n13620 = ~n13115 & n13618;
  assign n13621 = ~n13619 & ~n13620;
  assign n13622 = ~po46  & ~n13607;
  assign n13623 = ~n13614 & n13622;
  assign n13624 = ~n13621 & ~n13623;
  assign n13625 = ~n13616 & ~n13624;
  assign n13626 = po47  & ~n13625;
  assign n13627 = ~n13118 & ~n13120;
  assign n13628 = po11  & n13627;
  assign n13629 = n13125 & ~n13628;
  assign n13630 = ~n13125 & n13628;
  assign n13631 = ~n13629 & ~n13630;
  assign n13632 = ~po47  & n13625;
  assign n13633 = ~n13631 & ~n13632;
  assign n13634 = ~n13626 & ~n13633;
  assign n13635 = po48  & ~n13634;
  assign n13636 = ~po48  & ~n13626;
  assign n13637 = ~n13633 & n13636;
  assign n13638 = ~n13128 & po11 ;
  assign n13639 = ~n13134 & n13638;
  assign n13640 = n13133 & ~n13639;
  assign n13641 = n13135 & n13638;
  assign n13642 = ~n13640 & ~n13641;
  assign n13643 = ~n13637 & n13642;
  assign n13644 = ~n13635 & ~n13643;
  assign n13645 = po49  & ~n13644;
  assign n13646 = ~n13137 & ~n13139;
  assign n13647 = po11  & n13646;
  assign n13648 = n13144 & ~n13647;
  assign n13649 = ~n13144 & n13647;
  assign n13650 = ~n13648 & ~n13649;
  assign n13651 = ~po49  & n13644;
  assign n13652 = ~n13650 & ~n13651;
  assign n13653 = ~n13645 & ~n13652;
  assign n13654 = po50  & ~n13653;
  assign n13655 = ~n13147 & ~n13148;
  assign n13656 = po11  & n13655;
  assign n13657 = n13153 & ~n13656;
  assign n13658 = ~n13153 & n13656;
  assign n13659 = ~n13657 & ~n13658;
  assign n13660 = ~po50  & ~n13645;
  assign n13661 = ~n13652 & n13660;
  assign n13662 = ~n13659 & ~n13661;
  assign n13663 = ~n13654 & ~n13662;
  assign n13664 = ~po51  & n13663;
  assign n13665 = ~n13156 & po11 ;
  assign n13666 = ~n13163 & n13665;
  assign n13667 = n13161 & ~n13666;
  assign n13668 = n13164 & n13665;
  assign n13669 = ~n13667 & ~n13668;
  assign n13670 = ~n13664 & n13669;
  assign n13671 = po51  & ~n13663;
  assign n13672 = ~n13670 & ~n13671;
  assign n13673 = po52  & ~n13672;
  assign n13674 = ~n13166 & ~n13168;
  assign n13675 = po11  & n13674;
  assign n13676 = n12801 & ~n13675;
  assign n13677 = ~n12801 & n13675;
  assign n13678 = ~n13676 & ~n13677;
  assign n13679 = ~po52  & ~n13671;
  assign n13680 = ~n13670 & n13679;
  assign n13681 = n13678 & ~n13680;
  assign n13682 = ~n13673 & ~n13681;
  assign n13683 = ~po53  & n13682;
  assign n13684 = po53  & ~n13682;
  assign n13685 = ~n13290 & ~n13683;
  assign n13686 = ~n13684 & ~n13685;
  assign n13687 = po54  & ~n13686;
  assign n13688 = ~po54  & ~n13684;
  assign n13689 = ~n13685 & n13688;
  assign n13690 = ~n13175 & po11 ;
  assign n13691 = ~n13181 & n13690;
  assign n13692 = n13180 & ~n13691;
  assign n13693 = n13182 & n13690;
  assign n13694 = ~n13692 & ~n13693;
  assign n13695 = ~n13689 & n13694;
  assign n13696 = ~n13687 & ~n13695;
  assign n13697 = po55  & ~n13696;
  assign n13698 = ~n13184 & ~n13186;
  assign n13699 = po11  & n13698;
  assign n13700 = n13191 & ~n13699;
  assign n13701 = ~n13191 & n13699;
  assign n13702 = ~n13700 & ~n13701;
  assign n13703 = ~po55  & n13696;
  assign n13704 = ~n13702 & ~n13703;
  assign n13705 = ~n13697 & ~n13704;
  assign n13706 = po56  & ~n13705;
  assign n13707 = ~po56  & ~n13697;
  assign n13708 = ~n13704 & n13707;
  assign n13709 = ~n13194 & po11 ;
  assign n13710 = ~n13200 & n13709;
  assign n13711 = n13199 & ~n13710;
  assign n13712 = n13201 & n13709;
  assign n13713 = ~n13711 & ~n13712;
  assign n13714 = ~n13708 & n13713;
  assign n13715 = ~n13706 & ~n13714;
  assign n13716 = po57  & ~n13715;
  assign n13717 = ~n13203 & ~n13205;
  assign n13718 = po11  & n13717;
  assign n13719 = n13210 & ~n13718;
  assign n13720 = ~n13210 & n13718;
  assign n13721 = ~n13719 & ~n13720;
  assign n13722 = ~po57  & n13715;
  assign n13723 = ~n13721 & ~n13722;
  assign n13724 = ~n13716 & ~n13723;
  assign n13725 = po58  & ~n13724;
  assign n13726 = ~n13213 & ~n13214;
  assign n13727 = po11  & n13726;
  assign n13728 = n13219 & ~n13727;
  assign n13729 = ~n13219 & n13727;
  assign n13730 = ~n13728 & ~n13729;
  assign n13731 = ~po58  & ~n13716;
  assign n13732 = ~n13723 & n13731;
  assign n13733 = ~n13730 & ~n13732;
  assign n13734 = ~n13725 & ~n13733;
  assign n13735 = po59  & ~n13734;
  assign n13736 = ~n13222 & ~n13224;
  assign n13737 = po11  & n13736;
  assign n13738 = n13229 & ~n13737;
  assign n13739 = ~n13229 & n13737;
  assign n13740 = ~n13738 & ~n13739;
  assign n13741 = ~po59  & n13734;
  assign n13742 = ~n13740 & ~n13741;
  assign n13743 = ~n13735 & ~n13742;
  assign n13744 = po60  & ~n13743;
  assign n13745 = ~po60  & ~n13735;
  assign n13746 = ~n13742 & n13745;
  assign n13747 = ~n13232 & po11 ;
  assign n13748 = ~n13238 & n13747;
  assign n13749 = n13237 & ~n13748;
  assign n13750 = n13239 & n13747;
  assign n13751 = ~n13749 & ~n13750;
  assign n13752 = ~n13746 & n13751;
  assign n13753 = ~n13744 & ~n13752;
  assign n13754 = po61  & ~n13753;
  assign n13755 = ~n13241 & ~n13243;
  assign n13756 = po11  & n13755;
  assign n13757 = n13248 & ~n13756;
  assign n13758 = ~n13248 & n13756;
  assign n13759 = ~n13757 & ~n13758;
  assign n13760 = ~po61  & n13753;
  assign n13761 = ~n13759 & ~n13760;
  assign n13762 = ~n13754 & ~n13761;
  assign n13763 = po62  & ~n13762;
  assign n13764 = ~n13251 & ~n13252;
  assign n13765 = po11  & n13764;
  assign n13766 = n13257 & ~n13765;
  assign n13767 = ~n13257 & n13765;
  assign n13768 = ~n13766 & ~n13767;
  assign n13769 = ~po62  & ~n13754;
  assign n13770 = ~n13761 & n13769;
  assign n13771 = ~n13768 & ~n13770;
  assign n13772 = ~n13763 & ~n13771;
  assign n13773 = ~n13260 & ~n13262;
  assign n13774 = po11  & n13773;
  assign n13775 = n13267 & ~n13774;
  assign n13776 = ~n13267 & n13774;
  assign n13777 = ~n13775 & ~n13776;
  assign n13778 = n13269 & po11 ;
  assign n13779 = ~n13274 & ~n13778;
  assign n13780 = ~n13282 & ~n13779;
  assign n13781 = po11  & ~n13780;
  assign n13782 = ~n13777 & ~n13781;
  assign n13783 = ~n13772 & n13782;
  assign n13784 = ~po63  & ~n13783;
  assign n13785 = n13772 & n13777;
  assign n13786 = po63  & n13780;
  assign n13787 = ~n13785 & ~n13786;
  assign po10  = n13784 | ~n13787;
  assign n13789 = ~n13684 & po10 ;
  assign n13790 = ~n13683 & n13789;
  assign n13791 = n13290 & ~n13790;
  assign n13792 = n13685 & n13789;
  assign n13793 = ~n13791 & ~n13792;
  assign n13794 = pi20  & po10 ;
  assign n13795 = ~pi18  & ~pi19 ;
  assign n13796 = ~pi20  & n13795;
  assign n13797 = ~n13794 & ~n13796;
  assign n13798 = po11  & ~n13797;
  assign n13799 = ~pi20  & po10 ;
  assign n13800 = pi21  & ~n13799;
  assign n13801 = ~pi21  & n13799;
  assign n13802 = ~n13800 & ~n13801;
  assign n13803 = ~po11  & n13797;
  assign n13804 = n13802 & ~n13803;
  assign n13805 = ~n13798 & ~n13804;
  assign n13806 = po12  & ~n13805;
  assign n13807 = ~po12  & ~n13798;
  assign n13808 = ~n13804 & n13807;
  assign n13809 = po11  & ~po10 ;
  assign n13810 = ~n13801 & ~n13809;
  assign n13811 = pi22  & ~n13810;
  assign n13812 = ~pi22  & n13810;
  assign n13813 = ~n13811 & ~n13812;
  assign n13814 = ~n13808 & ~n13813;
  assign n13815 = ~n13806 & ~n13814;
  assign n13816 = po13  & ~n13815;
  assign n13817 = ~po13  & n13815;
  assign n13818 = ~n13295 & ~n13296;
  assign n13819 = po10  & n13818;
  assign n13820 = n13300 & ~n13819;
  assign n13821 = ~n13300 & n13819;
  assign n13822 = ~n13820 & ~n13821;
  assign n13823 = ~n13817 & ~n13822;
  assign n13824 = ~n13816 & ~n13823;
  assign n13825 = po14  & ~n13824;
  assign n13826 = ~po14  & ~n13816;
  assign n13827 = ~n13823 & n13826;
  assign n13828 = ~n13303 & po10 ;
  assign n13829 = ~n13309 & n13828;
  assign n13830 = n13308 & ~n13829;
  assign n13831 = n13310 & n13828;
  assign n13832 = ~n13830 & ~n13831;
  assign n13833 = ~n13827 & n13832;
  assign n13834 = ~n13825 & ~n13833;
  assign n13835 = po15  & ~n13834;
  assign n13836 = ~po15  & n13834;
  assign n13837 = ~n13312 & ~n13314;
  assign n13838 = po10  & n13837;
  assign n13839 = n13319 & ~n13838;
  assign n13840 = ~n13319 & n13838;
  assign n13841 = ~n13839 & ~n13840;
  assign n13842 = ~n13836 & n13841;
  assign n13843 = ~n13835 & ~n13842;
  assign n13844 = po16  & ~n13843;
  assign n13845 = ~po16  & ~n13835;
  assign n13846 = ~n13842 & n13845;
  assign n13847 = ~n13322 & po10 ;
  assign n13848 = ~n13328 & n13847;
  assign n13849 = n13327 & ~n13848;
  assign n13850 = n13329 & n13847;
  assign n13851 = ~n13849 & ~n13850;
  assign n13852 = ~n13846 & n13851;
  assign n13853 = ~n13844 & ~n13852;
  assign n13854 = po17  & ~n13853;
  assign n13855 = ~po17  & n13853;
  assign n13856 = ~n13331 & ~n13333;
  assign n13857 = po10  & n13856;
  assign n13858 = n13338 & n13857;
  assign n13859 = ~n13338 & ~n13857;
  assign n13860 = ~n13858 & ~n13859;
  assign n13861 = ~n13855 & n13860;
  assign n13862 = ~n13854 & ~n13861;
  assign n13863 = po18  & ~n13862;
  assign n13864 = ~po18  & ~n13854;
  assign n13865 = ~n13861 & n13864;
  assign n13866 = ~n13341 & po10 ;
  assign n13867 = ~n13347 & n13866;
  assign n13868 = n13346 & ~n13867;
  assign n13869 = n13348 & n13866;
  assign n13870 = ~n13868 & ~n13869;
  assign n13871 = ~n13865 & n13870;
  assign n13872 = ~n13863 & ~n13871;
  assign n13873 = po19  & ~n13872;
  assign n13874 = ~po19  & n13872;
  assign n13875 = ~n13350 & ~n13352;
  assign n13876 = po10  & n13875;
  assign n13877 = ~n13357 & ~n13876;
  assign n13878 = n13357 & n13876;
  assign n13879 = ~n13877 & ~n13878;
  assign n13880 = ~n13874 & n13879;
  assign n13881 = ~n13873 & ~n13880;
  assign n13882 = po20  & ~n13881;
  assign n13883 = ~po20  & ~n13873;
  assign n13884 = ~n13880 & n13883;
  assign n13885 = ~n13360 & po10 ;
  assign n13886 = ~n13366 & n13885;
  assign n13887 = n13365 & ~n13886;
  assign n13888 = n13367 & n13885;
  assign n13889 = ~n13887 & ~n13888;
  assign n13890 = ~n13884 & n13889;
  assign n13891 = ~n13882 & ~n13890;
  assign n13892 = po21  & ~n13891;
  assign n13893 = ~n13369 & ~n13371;
  assign n13894 = po10  & n13893;
  assign n13895 = n13376 & ~n13894;
  assign n13896 = ~n13376 & n13894;
  assign n13897 = ~n13895 & ~n13896;
  assign n13898 = ~po21  & n13891;
  assign n13899 = ~n13897 & ~n13898;
  assign n13900 = ~n13892 & ~n13899;
  assign n13901 = po22  & ~n13900;
  assign n13902 = ~po22  & ~n13892;
  assign n13903 = ~n13899 & n13902;
  assign n13904 = ~n13379 & po10 ;
  assign n13905 = ~n13385 & n13904;
  assign n13906 = n13384 & ~n13905;
  assign n13907 = n13386 & n13904;
  assign n13908 = ~n13906 & ~n13907;
  assign n13909 = ~n13903 & n13908;
  assign n13910 = ~n13901 & ~n13909;
  assign n13911 = po23  & ~n13910;
  assign n13912 = ~po23  & n13910;
  assign n13913 = ~n13388 & po10 ;
  assign n13914 = ~n13395 & n13913;
  assign n13915 = n13393 & ~n13914;
  assign n13916 = n13396 & n13913;
  assign n13917 = ~n13915 & ~n13916;
  assign n13918 = ~n13912 & n13917;
  assign n13919 = ~n13911 & ~n13918;
  assign n13920 = po24  & ~n13919;
  assign n13921 = ~po24  & ~n13911;
  assign n13922 = ~n13918 & n13921;
  assign n13923 = ~n13398 & po10 ;
  assign n13924 = ~n13404 & n13923;
  assign n13925 = n13403 & ~n13924;
  assign n13926 = n13405 & n13923;
  assign n13927 = ~n13925 & ~n13926;
  assign n13928 = ~n13922 & n13927;
  assign n13929 = ~n13920 & ~n13928;
  assign n13930 = po25  & ~n13929;
  assign n13931 = ~n13407 & ~n13409;
  assign n13932 = po10  & n13931;
  assign n13933 = n13414 & ~n13932;
  assign n13934 = ~n13414 & n13932;
  assign n13935 = ~n13933 & ~n13934;
  assign n13936 = ~po25  & n13929;
  assign n13937 = ~n13935 & ~n13936;
  assign n13938 = ~n13930 & ~n13937;
  assign n13939 = po26  & ~n13938;
  assign n13940 = ~po26  & ~n13930;
  assign n13941 = ~n13937 & n13940;
  assign n13942 = ~n13417 & po10 ;
  assign n13943 = ~n13423 & n13942;
  assign n13944 = n13422 & ~n13943;
  assign n13945 = n13424 & n13942;
  assign n13946 = ~n13944 & ~n13945;
  assign n13947 = ~n13941 & n13946;
  assign n13948 = ~n13939 & ~n13947;
  assign n13949 = po27  & ~n13948;
  assign n13950 = ~po27  & n13948;
  assign n13951 = ~n13426 & po10 ;
  assign n13952 = ~n13433 & n13951;
  assign n13953 = n13431 & ~n13952;
  assign n13954 = n13434 & n13951;
  assign n13955 = ~n13953 & ~n13954;
  assign n13956 = ~n13950 & n13955;
  assign n13957 = ~n13949 & ~n13956;
  assign n13958 = po28  & ~n13957;
  assign n13959 = ~po28  & ~n13949;
  assign n13960 = ~n13956 & n13959;
  assign n13961 = ~n13436 & po10 ;
  assign n13962 = ~n13442 & n13961;
  assign n13963 = n13441 & ~n13962;
  assign n13964 = n13443 & n13961;
  assign n13965 = ~n13963 & ~n13964;
  assign n13966 = ~n13960 & n13965;
  assign n13967 = ~n13958 & ~n13966;
  assign n13968 = po29  & ~n13967;
  assign n13969 = ~n13445 & ~n13447;
  assign n13970 = po10  & n13969;
  assign n13971 = n13452 & ~n13970;
  assign n13972 = ~n13452 & n13970;
  assign n13973 = ~n13971 & ~n13972;
  assign n13974 = ~po29  & n13967;
  assign n13975 = ~n13973 & ~n13974;
  assign n13976 = ~n13968 & ~n13975;
  assign n13977 = po30  & ~n13976;
  assign n13978 = ~po30  & ~n13968;
  assign n13979 = ~n13975 & n13978;
  assign n13980 = ~n13455 & po10 ;
  assign n13981 = ~n13461 & n13980;
  assign n13982 = n13460 & ~n13981;
  assign n13983 = n13462 & n13980;
  assign n13984 = ~n13982 & ~n13983;
  assign n13985 = ~n13979 & n13984;
  assign n13986 = ~n13977 & ~n13985;
  assign n13987 = po31  & ~n13986;
  assign n13988 = ~po31  & n13986;
  assign n13989 = ~n13464 & po10 ;
  assign n13990 = ~n13471 & n13989;
  assign n13991 = n13469 & ~n13990;
  assign n13992 = n13472 & n13989;
  assign n13993 = ~n13991 & ~n13992;
  assign n13994 = ~n13988 & n13993;
  assign n13995 = ~n13987 & ~n13994;
  assign n13996 = po32  & ~n13995;
  assign n13997 = ~po32  & ~n13987;
  assign n13998 = ~n13994 & n13997;
  assign n13999 = ~n13474 & po10 ;
  assign n14000 = ~n13480 & n13999;
  assign n14001 = n13479 & ~n14000;
  assign n14002 = n13481 & n13999;
  assign n14003 = ~n14001 & ~n14002;
  assign n14004 = ~n13998 & n14003;
  assign n14005 = ~n13996 & ~n14004;
  assign n14006 = po33  & ~n14005;
  assign n14007 = ~n13483 & ~n13485;
  assign n14008 = po10  & n14007;
  assign n14009 = n13490 & ~n14008;
  assign n14010 = ~n13490 & n14008;
  assign n14011 = ~n14009 & ~n14010;
  assign n14012 = ~po33  & n14005;
  assign n14013 = ~n14011 & ~n14012;
  assign n14014 = ~n14006 & ~n14013;
  assign n14015 = po34  & ~n14014;
  assign n14016 = ~po34  & ~n14006;
  assign n14017 = ~n14013 & n14016;
  assign n14018 = ~n13493 & po10 ;
  assign n14019 = ~n13499 & n14018;
  assign n14020 = n13498 & ~n14019;
  assign n14021 = n13500 & n14018;
  assign n14022 = ~n14020 & ~n14021;
  assign n14023 = ~n14017 & n14022;
  assign n14024 = ~n14015 & ~n14023;
  assign n14025 = po35  & ~n14024;
  assign n14026 = ~po35  & n14024;
  assign n14027 = ~n13502 & po10 ;
  assign n14028 = ~n13509 & n14027;
  assign n14029 = n13507 & ~n14028;
  assign n14030 = n13510 & n14027;
  assign n14031 = ~n14029 & ~n14030;
  assign n14032 = ~n14026 & n14031;
  assign n14033 = ~n14025 & ~n14032;
  assign n14034 = po36  & ~n14033;
  assign n14035 = ~po36  & ~n14025;
  assign n14036 = ~n14032 & n14035;
  assign n14037 = ~n13512 & po10 ;
  assign n14038 = ~n13518 & n14037;
  assign n14039 = n13517 & ~n14038;
  assign n14040 = n13519 & n14037;
  assign n14041 = ~n14039 & ~n14040;
  assign n14042 = ~n14036 & n14041;
  assign n14043 = ~n14034 & ~n14042;
  assign n14044 = po37  & ~n14043;
  assign n14045 = ~n13521 & ~n13523;
  assign n14046 = po10  & n14045;
  assign n14047 = n13528 & ~n14046;
  assign n14048 = ~n13528 & n14046;
  assign n14049 = ~n14047 & ~n14048;
  assign n14050 = ~po37  & n14043;
  assign n14051 = ~n14049 & ~n14050;
  assign n14052 = ~n14044 & ~n14051;
  assign n14053 = po38  & ~n14052;
  assign n14054 = ~po38  & ~n14044;
  assign n14055 = ~n14051 & n14054;
  assign n14056 = ~n13531 & po10 ;
  assign n14057 = ~n13537 & n14056;
  assign n14058 = n13536 & ~n14057;
  assign n14059 = n13538 & n14056;
  assign n14060 = ~n14058 & ~n14059;
  assign n14061 = ~n14055 & n14060;
  assign n14062 = ~n14053 & ~n14061;
  assign n14063 = po39  & ~n14062;
  assign n14064 = ~po39  & n14062;
  assign n14065 = ~n13540 & po10 ;
  assign n14066 = ~n13547 & n14065;
  assign n14067 = n13545 & ~n14066;
  assign n14068 = n13548 & n14065;
  assign n14069 = ~n14067 & ~n14068;
  assign n14070 = ~n14064 & n14069;
  assign n14071 = ~n14063 & ~n14070;
  assign n14072 = po40  & ~n14071;
  assign n14073 = ~po40  & ~n14063;
  assign n14074 = ~n14070 & n14073;
  assign n14075 = ~n13550 & po10 ;
  assign n14076 = ~n13556 & n14075;
  assign n14077 = n13555 & ~n14076;
  assign n14078 = n13557 & n14075;
  assign n14079 = ~n14077 & ~n14078;
  assign n14080 = ~n14074 & n14079;
  assign n14081 = ~n14072 & ~n14080;
  assign n14082 = po41  & ~n14081;
  assign n14083 = ~n13559 & ~n13561;
  assign n14084 = po10  & n14083;
  assign n14085 = n13566 & ~n14084;
  assign n14086 = ~n13566 & n14084;
  assign n14087 = ~n14085 & ~n14086;
  assign n14088 = ~po41  & n14081;
  assign n14089 = ~n14087 & ~n14088;
  assign n14090 = ~n14082 & ~n14089;
  assign n14091 = po42  & ~n14090;
  assign n14092 = ~po42  & ~n14082;
  assign n14093 = ~n14089 & n14092;
  assign n14094 = ~n13569 & po10 ;
  assign n14095 = ~n13575 & n14094;
  assign n14096 = n13574 & ~n14095;
  assign n14097 = n13576 & n14094;
  assign n14098 = ~n14096 & ~n14097;
  assign n14099 = ~n14093 & n14098;
  assign n14100 = ~n14091 & ~n14099;
  assign n14101 = po43  & ~n14100;
  assign n14102 = ~po43  & n14100;
  assign n14103 = ~n13578 & po10 ;
  assign n14104 = ~n13585 & n14103;
  assign n14105 = n13583 & ~n14104;
  assign n14106 = n13586 & n14103;
  assign n14107 = ~n14105 & ~n14106;
  assign n14108 = ~n14102 & n14107;
  assign n14109 = ~n14101 & ~n14108;
  assign n14110 = po44  & ~n14109;
  assign n14111 = ~po44  & ~n14101;
  assign n14112 = ~n14108 & n14111;
  assign n14113 = ~n13588 & po10 ;
  assign n14114 = ~n13594 & n14113;
  assign n14115 = n13593 & ~n14114;
  assign n14116 = n13595 & n14113;
  assign n14117 = ~n14115 & ~n14116;
  assign n14118 = ~n14112 & n14117;
  assign n14119 = ~n14110 & ~n14118;
  assign n14120 = po45  & ~n14119;
  assign n14121 = ~n13597 & ~n13599;
  assign n14122 = po10  & n14121;
  assign n14123 = n13604 & ~n14122;
  assign n14124 = ~n13604 & n14122;
  assign n14125 = ~n14123 & ~n14124;
  assign n14126 = ~po45  & n14119;
  assign n14127 = ~n14125 & ~n14126;
  assign n14128 = ~n14120 & ~n14127;
  assign n14129 = po46  & ~n14128;
  assign n14130 = ~po46  & ~n14120;
  assign n14131 = ~n14127 & n14130;
  assign n14132 = ~n13607 & po10 ;
  assign n14133 = ~n13613 & n14132;
  assign n14134 = n13612 & ~n14133;
  assign n14135 = n13614 & n14132;
  assign n14136 = ~n14134 & ~n14135;
  assign n14137 = ~n14131 & n14136;
  assign n14138 = ~n14129 & ~n14137;
  assign n14139 = po47  & ~n14138;
  assign n14140 = ~po47  & n14138;
  assign n14141 = ~n13616 & po10 ;
  assign n14142 = ~n13623 & n14141;
  assign n14143 = n13621 & ~n14142;
  assign n14144 = n13624 & n14141;
  assign n14145 = ~n14143 & ~n14144;
  assign n14146 = ~n14140 & n14145;
  assign n14147 = ~n14139 & ~n14146;
  assign n14148 = po48  & ~n14147;
  assign n14149 = ~po48  & ~n14139;
  assign n14150 = ~n14146 & n14149;
  assign n14151 = ~n13626 & po10 ;
  assign n14152 = ~n13632 & n14151;
  assign n14153 = n13631 & ~n14152;
  assign n14154 = n13633 & n14151;
  assign n14155 = ~n14153 & ~n14154;
  assign n14156 = ~n14150 & n14155;
  assign n14157 = ~n14148 & ~n14156;
  assign n14158 = po49  & ~n14157;
  assign n14159 = ~n13635 & ~n13637;
  assign n14160 = po10  & n14159;
  assign n14161 = n13642 & ~n14160;
  assign n14162 = ~n13642 & n14160;
  assign n14163 = ~n14161 & ~n14162;
  assign n14164 = ~po49  & n14157;
  assign n14165 = ~n14163 & ~n14164;
  assign n14166 = ~n14158 & ~n14165;
  assign n14167 = po50  & ~n14166;
  assign n14168 = ~po50  & ~n14158;
  assign n14169 = ~n14165 & n14168;
  assign n14170 = ~n13645 & po10 ;
  assign n14171 = ~n13651 & n14170;
  assign n14172 = n13650 & ~n14171;
  assign n14173 = n13652 & n14170;
  assign n14174 = ~n14172 & ~n14173;
  assign n14175 = ~n14169 & n14174;
  assign n14176 = ~n14167 & ~n14175;
  assign n14177 = po51  & ~n14176;
  assign n14178 = ~po51  & n14176;
  assign n14179 = ~n13654 & po10 ;
  assign n14180 = ~n13661 & n14179;
  assign n14181 = n13659 & ~n14180;
  assign n14182 = n13662 & n14179;
  assign n14183 = ~n14181 & ~n14182;
  assign n14184 = ~n14178 & n14183;
  assign n14185 = ~n14177 & ~n14184;
  assign n14186 = po52  & ~n14185;
  assign n14187 = ~n13664 & ~n13671;
  assign n14188 = po10  & n14187;
  assign n14189 = n13669 & ~n14188;
  assign n14190 = ~n13669 & n14188;
  assign n14191 = ~n14189 & ~n14190;
  assign n14192 = ~po52  & ~n14177;
  assign n14193 = ~n14184 & n14192;
  assign n14194 = ~n14191 & ~n14193;
  assign n14195 = ~n14186 & ~n14194;
  assign n14196 = ~po53  & n14195;
  assign n14197 = ~n13673 & ~n13680;
  assign n14198 = po10  & n14197;
  assign n14199 = n13678 & n14198;
  assign n14200 = ~n13678 & ~n14198;
  assign n14201 = ~n14199 & ~n14200;
  assign n14202 = ~n14196 & n14201;
  assign n14203 = po53  & ~n14195;
  assign n14204 = ~po54  & ~n14203;
  assign n14205 = ~n14202 & n14204;
  assign n14206 = ~n14202 & ~n14203;
  assign n14207 = po54  & ~n14206;
  assign n14208 = n13793 & ~n14205;
  assign n14209 = ~n14207 & ~n14208;
  assign n14210 = po55  & ~n14209;
  assign n14211 = ~n13687 & ~n13689;
  assign n14212 = po10  & n14211;
  assign n14213 = n13694 & ~n14212;
  assign n14214 = ~n13694 & n14212;
  assign n14215 = ~n14213 & ~n14214;
  assign n14216 = ~po55  & n14209;
  assign n14217 = ~n14215 & ~n14216;
  assign n14218 = ~n14210 & ~n14217;
  assign n14219 = po56  & ~n14218;
  assign n14220 = ~po56  & ~n14210;
  assign n14221 = ~n14217 & n14220;
  assign n14222 = ~n13697 & po10 ;
  assign n14223 = ~n13703 & n14222;
  assign n14224 = n13702 & ~n14223;
  assign n14225 = n13704 & n14222;
  assign n14226 = ~n14224 & ~n14225;
  assign n14227 = ~n14221 & n14226;
  assign n14228 = ~n14219 & ~n14227;
  assign n14229 = po57  & ~n14228;
  assign n14230 = ~n13706 & ~n13708;
  assign n14231 = po10  & n14230;
  assign n14232 = n13713 & ~n14231;
  assign n14233 = ~n13713 & n14231;
  assign n14234 = ~n14232 & ~n14233;
  assign n14235 = ~po57  & n14228;
  assign n14236 = ~n14234 & ~n14235;
  assign n14237 = ~n14229 & ~n14236;
  assign n14238 = po58  & ~n14237;
  assign n14239 = ~po58  & ~n14229;
  assign n14240 = ~n14236 & n14239;
  assign n14241 = ~n13716 & po10 ;
  assign n14242 = ~n13722 & n14241;
  assign n14243 = n13721 & ~n14242;
  assign n14244 = n13723 & n14241;
  assign n14245 = ~n14243 & ~n14244;
  assign n14246 = ~n14240 & n14245;
  assign n14247 = ~n14238 & ~n14246;
  assign n14248 = po59  & ~n14247;
  assign n14249 = ~po59  & n14247;
  assign n14250 = ~n13725 & po10 ;
  assign n14251 = ~n13732 & n14250;
  assign n14252 = n13730 & ~n14251;
  assign n14253 = n13733 & n14250;
  assign n14254 = ~n14252 & ~n14253;
  assign n14255 = ~n14249 & n14254;
  assign n14256 = ~n14248 & ~n14255;
  assign n14257 = po60  & ~n14256;
  assign n14258 = ~po60  & ~n14248;
  assign n14259 = ~n14255 & n14258;
  assign n14260 = ~n13735 & po10 ;
  assign n14261 = ~n13741 & n14260;
  assign n14262 = n13740 & ~n14261;
  assign n14263 = n13742 & n14260;
  assign n14264 = ~n14262 & ~n14263;
  assign n14265 = ~n14259 & n14264;
  assign n14266 = ~n14257 & ~n14265;
  assign n14267 = po61  & ~n14266;
  assign n14268 = ~n13744 & ~n13746;
  assign n14269 = po10  & n14268;
  assign n14270 = n13751 & ~n14269;
  assign n14271 = ~n13751 & n14269;
  assign n14272 = ~n14270 & ~n14271;
  assign n14273 = ~po61  & n14266;
  assign n14274 = ~n14272 & ~n14273;
  assign n14275 = ~n14267 & ~n14274;
  assign n14276 = po62  & ~n14275;
  assign n14277 = ~po62  & ~n14267;
  assign n14278 = ~n14274 & n14277;
  assign n14279 = ~n13754 & po10 ;
  assign n14280 = ~n13760 & n14279;
  assign n14281 = n13759 & ~n14280;
  assign n14282 = n13761 & n14279;
  assign n14283 = ~n14281 & ~n14282;
  assign n14284 = ~n14278 & n14283;
  assign n14285 = ~n14276 & ~n14284;
  assign n14286 = n13772 & po10 ;
  assign n14287 = ~n13777 & ~n14286;
  assign n14288 = ~n13785 & ~n14287;
  assign n14289 = po10  & ~n14288;
  assign n14290 = ~n13763 & po10 ;
  assign n14291 = ~n13770 & n14290;
  assign n14292 = n13768 & ~n14291;
  assign n14293 = n13771 & n14290;
  assign n14294 = ~n14292 & ~n14293;
  assign n14295 = ~n14289 & n14294;
  assign n14296 = ~n14285 & n14295;
  assign n14297 = ~po63  & ~n14296;
  assign n14298 = n14285 & ~n14294;
  assign n14299 = po63  & n14288;
  assign n14300 = ~n14298 & ~n14299;
  assign po9  = n14297 | ~n14300;
  assign n14302 = ~n14205 & ~n14207;
  assign n14303 = po9  & n14302;
  assign n14304 = n13793 & ~n14303;
  assign n14305 = ~n13793 & n14303;
  assign n14306 = ~n14304 & ~n14305;
  assign n14307 = pi18  & po9 ;
  assign n14308 = ~pi16  & ~pi17 ;
  assign n14309 = ~pi18  & n14308;
  assign n14310 = ~n14307 & ~n14309;
  assign n14311 = po10  & ~n14310;
  assign n14312 = ~po10  & n14310;
  assign n14313 = ~pi18  & po9 ;
  assign n14314 = pi19  & ~n14313;
  assign n14315 = ~pi19  & n14313;
  assign n14316 = ~n14314 & ~n14315;
  assign n14317 = ~n14312 & n14316;
  assign n14318 = ~n14311 & ~n14317;
  assign n14319 = po11  & ~n14318;
  assign n14320 = po10  & ~po9 ;
  assign n14321 = ~n14315 & ~n14320;
  assign n14322 = pi20  & ~n14321;
  assign n14323 = ~pi20  & n14321;
  assign n14324 = ~n14322 & ~n14323;
  assign n14325 = ~po11  & n14318;
  assign n14326 = ~n14324 & ~n14325;
  assign n14327 = ~n14319 & ~n14326;
  assign n14328 = po12  & ~n14327;
  assign n14329 = ~po12  & ~n14319;
  assign n14330 = ~n14326 & n14329;
  assign n14331 = ~n13798 & ~n13803;
  assign n14332 = po9  & n14331;
  assign n14333 = n13802 & ~n14332;
  assign n14334 = ~n13802 & n14332;
  assign n14335 = ~n14333 & ~n14334;
  assign n14336 = ~n14330 & ~n14335;
  assign n14337 = ~n14328 & ~n14336;
  assign n14338 = po13  & ~n14337;
  assign n14339 = ~n13806 & ~n13808;
  assign n14340 = po9  & n14339;
  assign n14341 = ~n13813 & ~n14340;
  assign n14342 = n13813 & n14340;
  assign n14343 = ~n14341 & ~n14342;
  assign n14344 = ~po13  & n14337;
  assign n14345 = ~n14343 & ~n14344;
  assign n14346 = ~n14338 & ~n14345;
  assign n14347 = po14  & ~n14346;
  assign n14348 = ~po14  & ~n14338;
  assign n14349 = ~n14345 & n14348;
  assign n14350 = ~n13816 & ~n13817;
  assign n14351 = po9  & n14350;
  assign n14352 = n13822 & ~n14351;
  assign n14353 = ~n13822 & n14351;
  assign n14354 = ~n14352 & ~n14353;
  assign n14355 = ~n14349 & n14354;
  assign n14356 = ~n14347 & ~n14355;
  assign n14357 = po15  & ~n14356;
  assign n14358 = ~n13825 & ~n13827;
  assign n14359 = po9  & n14358;
  assign n14360 = n13832 & ~n14359;
  assign n14361 = ~n13832 & n14359;
  assign n14362 = ~n14360 & ~n14361;
  assign n14363 = ~po15  & n14356;
  assign n14364 = ~n14362 & ~n14363;
  assign n14365 = ~n14357 & ~n14364;
  assign n14366 = po16  & ~n14365;
  assign n14367 = ~po16  & ~n14357;
  assign n14368 = ~n14364 & n14367;
  assign n14369 = ~n13835 & ~n13836;
  assign n14370 = po9  & n14369;
  assign n14371 = n13841 & n14370;
  assign n14372 = ~n13841 & ~n14370;
  assign n14373 = ~n14371 & ~n14372;
  assign n14374 = ~n14368 & n14373;
  assign n14375 = ~n14366 & ~n14374;
  assign n14376 = po17  & ~n14375;
  assign n14377 = ~n13844 & ~n13846;
  assign n14378 = po9  & n14377;
  assign n14379 = n13851 & ~n14378;
  assign n14380 = ~n13851 & n14378;
  assign n14381 = ~n14379 & ~n14380;
  assign n14382 = ~po17  & n14375;
  assign n14383 = ~n14381 & ~n14382;
  assign n14384 = ~n14376 & ~n14383;
  assign n14385 = po18  & ~n14384;
  assign n14386 = ~po18  & ~n14376;
  assign n14387 = ~n14383 & n14386;
  assign n14388 = ~n13854 & ~n13855;
  assign n14389 = po9  & n14388;
  assign n14390 = ~n13860 & ~n14389;
  assign n14391 = n13860 & n14389;
  assign n14392 = ~n14390 & ~n14391;
  assign n14393 = ~n14387 & n14392;
  assign n14394 = ~n14385 & ~n14393;
  assign n14395 = po19  & ~n14394;
  assign n14396 = ~n13863 & ~n13865;
  assign n14397 = po9  & n14396;
  assign n14398 = n13870 & ~n14397;
  assign n14399 = ~n13870 & n14397;
  assign n14400 = ~n14398 & ~n14399;
  assign n14401 = ~po19  & n14394;
  assign n14402 = ~n14400 & ~n14401;
  assign n14403 = ~n14395 & ~n14402;
  assign n14404 = po20  & ~n14403;
  assign n14405 = ~n13873 & ~n13874;
  assign n14406 = po9  & n14405;
  assign n14407 = n13879 & ~n14406;
  assign n14408 = ~n13879 & n14406;
  assign n14409 = ~n14407 & ~n14408;
  assign n14410 = ~po20  & ~n14395;
  assign n14411 = ~n14402 & n14410;
  assign n14412 = ~n14409 & ~n14411;
  assign n14413 = ~n14404 & ~n14412;
  assign n14414 = po21  & ~n14413;
  assign n14415 = ~n13882 & ~n13884;
  assign n14416 = po9  & n14415;
  assign n14417 = n13889 & ~n14416;
  assign n14418 = ~n13889 & n14416;
  assign n14419 = ~n14417 & ~n14418;
  assign n14420 = ~po21  & n14413;
  assign n14421 = ~n14419 & ~n14420;
  assign n14422 = ~n14414 & ~n14421;
  assign n14423 = po22  & ~n14422;
  assign n14424 = ~po22  & ~n14414;
  assign n14425 = ~n14421 & n14424;
  assign n14426 = ~n13892 & po9 ;
  assign n14427 = ~n13898 & n14426;
  assign n14428 = n13897 & ~n14427;
  assign n14429 = n13899 & n14426;
  assign n14430 = ~n14428 & ~n14429;
  assign n14431 = ~n14425 & n14430;
  assign n14432 = ~n14423 & ~n14431;
  assign n14433 = po23  & ~n14432;
  assign n14434 = ~n13901 & ~n13903;
  assign n14435 = po9  & n14434;
  assign n14436 = n13908 & ~n14435;
  assign n14437 = ~n13908 & n14435;
  assign n14438 = ~n14436 & ~n14437;
  assign n14439 = ~po23  & n14432;
  assign n14440 = ~n14438 & ~n14439;
  assign n14441 = ~n14433 & ~n14440;
  assign n14442 = po24  & ~n14441;
  assign n14443 = ~n13911 & ~n13912;
  assign n14444 = po9  & n14443;
  assign n14445 = n13917 & ~n14444;
  assign n14446 = ~n13917 & n14444;
  assign n14447 = ~n14445 & ~n14446;
  assign n14448 = ~po24  & ~n14433;
  assign n14449 = ~n14440 & n14448;
  assign n14450 = ~n14447 & ~n14449;
  assign n14451 = ~n14442 & ~n14450;
  assign n14452 = po25  & ~n14451;
  assign n14453 = ~n13920 & ~n13922;
  assign n14454 = po9  & n14453;
  assign n14455 = n13927 & ~n14454;
  assign n14456 = ~n13927 & n14454;
  assign n14457 = ~n14455 & ~n14456;
  assign n14458 = ~po25  & n14451;
  assign n14459 = ~n14457 & ~n14458;
  assign n14460 = ~n14452 & ~n14459;
  assign n14461 = po26  & ~n14460;
  assign n14462 = ~po26  & ~n14452;
  assign n14463 = ~n14459 & n14462;
  assign n14464 = ~n13930 & po9 ;
  assign n14465 = ~n13936 & n14464;
  assign n14466 = n13935 & ~n14465;
  assign n14467 = n13937 & n14464;
  assign n14468 = ~n14466 & ~n14467;
  assign n14469 = ~n14463 & n14468;
  assign n14470 = ~n14461 & ~n14469;
  assign n14471 = po27  & ~n14470;
  assign n14472 = ~n13939 & ~n13941;
  assign n14473 = po9  & n14472;
  assign n14474 = n13946 & ~n14473;
  assign n14475 = ~n13946 & n14473;
  assign n14476 = ~n14474 & ~n14475;
  assign n14477 = ~po27  & n14470;
  assign n14478 = ~n14476 & ~n14477;
  assign n14479 = ~n14471 & ~n14478;
  assign n14480 = po28  & ~n14479;
  assign n14481 = ~n13949 & ~n13950;
  assign n14482 = po9  & n14481;
  assign n14483 = n13955 & ~n14482;
  assign n14484 = ~n13955 & n14482;
  assign n14485 = ~n14483 & ~n14484;
  assign n14486 = ~po28  & ~n14471;
  assign n14487 = ~n14478 & n14486;
  assign n14488 = ~n14485 & ~n14487;
  assign n14489 = ~n14480 & ~n14488;
  assign n14490 = po29  & ~n14489;
  assign n14491 = ~n13958 & ~n13960;
  assign n14492 = po9  & n14491;
  assign n14493 = n13965 & ~n14492;
  assign n14494 = ~n13965 & n14492;
  assign n14495 = ~n14493 & ~n14494;
  assign n14496 = ~po29  & n14489;
  assign n14497 = ~n14495 & ~n14496;
  assign n14498 = ~n14490 & ~n14497;
  assign n14499 = po30  & ~n14498;
  assign n14500 = ~po30  & ~n14490;
  assign n14501 = ~n14497 & n14500;
  assign n14502 = ~n13968 & po9 ;
  assign n14503 = ~n13974 & n14502;
  assign n14504 = n13973 & ~n14503;
  assign n14505 = n13975 & n14502;
  assign n14506 = ~n14504 & ~n14505;
  assign n14507 = ~n14501 & n14506;
  assign n14508 = ~n14499 & ~n14507;
  assign n14509 = po31  & ~n14508;
  assign n14510 = ~n13977 & ~n13979;
  assign n14511 = po9  & n14510;
  assign n14512 = n13984 & ~n14511;
  assign n14513 = ~n13984 & n14511;
  assign n14514 = ~n14512 & ~n14513;
  assign n14515 = ~po31  & n14508;
  assign n14516 = ~n14514 & ~n14515;
  assign n14517 = ~n14509 & ~n14516;
  assign n14518 = po32  & ~n14517;
  assign n14519 = ~n13987 & ~n13988;
  assign n14520 = po9  & n14519;
  assign n14521 = n13993 & ~n14520;
  assign n14522 = ~n13993 & n14520;
  assign n14523 = ~n14521 & ~n14522;
  assign n14524 = ~po32  & ~n14509;
  assign n14525 = ~n14516 & n14524;
  assign n14526 = ~n14523 & ~n14525;
  assign n14527 = ~n14518 & ~n14526;
  assign n14528 = po33  & ~n14527;
  assign n14529 = ~n13996 & ~n13998;
  assign n14530 = po9  & n14529;
  assign n14531 = n14003 & ~n14530;
  assign n14532 = ~n14003 & n14530;
  assign n14533 = ~n14531 & ~n14532;
  assign n14534 = ~po33  & n14527;
  assign n14535 = ~n14533 & ~n14534;
  assign n14536 = ~n14528 & ~n14535;
  assign n14537 = po34  & ~n14536;
  assign n14538 = ~po34  & ~n14528;
  assign n14539 = ~n14535 & n14538;
  assign n14540 = ~n14006 & po9 ;
  assign n14541 = ~n14012 & n14540;
  assign n14542 = n14011 & ~n14541;
  assign n14543 = n14013 & n14540;
  assign n14544 = ~n14542 & ~n14543;
  assign n14545 = ~n14539 & n14544;
  assign n14546 = ~n14537 & ~n14545;
  assign n14547 = po35  & ~n14546;
  assign n14548 = ~n14015 & ~n14017;
  assign n14549 = po9  & n14548;
  assign n14550 = n14022 & ~n14549;
  assign n14551 = ~n14022 & n14549;
  assign n14552 = ~n14550 & ~n14551;
  assign n14553 = ~po35  & n14546;
  assign n14554 = ~n14552 & ~n14553;
  assign n14555 = ~n14547 & ~n14554;
  assign n14556 = po36  & ~n14555;
  assign n14557 = ~n14025 & ~n14026;
  assign n14558 = po9  & n14557;
  assign n14559 = n14031 & ~n14558;
  assign n14560 = ~n14031 & n14558;
  assign n14561 = ~n14559 & ~n14560;
  assign n14562 = ~po36  & ~n14547;
  assign n14563 = ~n14554 & n14562;
  assign n14564 = ~n14561 & ~n14563;
  assign n14565 = ~n14556 & ~n14564;
  assign n14566 = po37  & ~n14565;
  assign n14567 = ~n14034 & ~n14036;
  assign n14568 = po9  & n14567;
  assign n14569 = n14041 & ~n14568;
  assign n14570 = ~n14041 & n14568;
  assign n14571 = ~n14569 & ~n14570;
  assign n14572 = ~po37  & n14565;
  assign n14573 = ~n14571 & ~n14572;
  assign n14574 = ~n14566 & ~n14573;
  assign n14575 = po38  & ~n14574;
  assign n14576 = ~po38  & ~n14566;
  assign n14577 = ~n14573 & n14576;
  assign n14578 = ~n14044 & po9 ;
  assign n14579 = ~n14050 & n14578;
  assign n14580 = n14049 & ~n14579;
  assign n14581 = n14051 & n14578;
  assign n14582 = ~n14580 & ~n14581;
  assign n14583 = ~n14577 & n14582;
  assign n14584 = ~n14575 & ~n14583;
  assign n14585 = po39  & ~n14584;
  assign n14586 = ~n14053 & ~n14055;
  assign n14587 = po9  & n14586;
  assign n14588 = n14060 & ~n14587;
  assign n14589 = ~n14060 & n14587;
  assign n14590 = ~n14588 & ~n14589;
  assign n14591 = ~po39  & n14584;
  assign n14592 = ~n14590 & ~n14591;
  assign n14593 = ~n14585 & ~n14592;
  assign n14594 = po40  & ~n14593;
  assign n14595 = ~n14063 & ~n14064;
  assign n14596 = po9  & n14595;
  assign n14597 = n14069 & ~n14596;
  assign n14598 = ~n14069 & n14596;
  assign n14599 = ~n14597 & ~n14598;
  assign n14600 = ~po40  & ~n14585;
  assign n14601 = ~n14592 & n14600;
  assign n14602 = ~n14599 & ~n14601;
  assign n14603 = ~n14594 & ~n14602;
  assign n14604 = po41  & ~n14603;
  assign n14605 = ~n14072 & ~n14074;
  assign n14606 = po9  & n14605;
  assign n14607 = n14079 & ~n14606;
  assign n14608 = ~n14079 & n14606;
  assign n14609 = ~n14607 & ~n14608;
  assign n14610 = ~po41  & n14603;
  assign n14611 = ~n14609 & ~n14610;
  assign n14612 = ~n14604 & ~n14611;
  assign n14613 = po42  & ~n14612;
  assign n14614 = ~po42  & ~n14604;
  assign n14615 = ~n14611 & n14614;
  assign n14616 = ~n14082 & po9 ;
  assign n14617 = ~n14088 & n14616;
  assign n14618 = n14087 & ~n14617;
  assign n14619 = n14089 & n14616;
  assign n14620 = ~n14618 & ~n14619;
  assign n14621 = ~n14615 & n14620;
  assign n14622 = ~n14613 & ~n14621;
  assign n14623 = po43  & ~n14622;
  assign n14624 = ~n14091 & ~n14093;
  assign n14625 = po9  & n14624;
  assign n14626 = n14098 & ~n14625;
  assign n14627 = ~n14098 & n14625;
  assign n14628 = ~n14626 & ~n14627;
  assign n14629 = ~po43  & n14622;
  assign n14630 = ~n14628 & ~n14629;
  assign n14631 = ~n14623 & ~n14630;
  assign n14632 = po44  & ~n14631;
  assign n14633 = ~n14101 & ~n14102;
  assign n14634 = po9  & n14633;
  assign n14635 = n14107 & ~n14634;
  assign n14636 = ~n14107 & n14634;
  assign n14637 = ~n14635 & ~n14636;
  assign n14638 = ~po44  & ~n14623;
  assign n14639 = ~n14630 & n14638;
  assign n14640 = ~n14637 & ~n14639;
  assign n14641 = ~n14632 & ~n14640;
  assign n14642 = po45  & ~n14641;
  assign n14643 = ~n14110 & ~n14112;
  assign n14644 = po9  & n14643;
  assign n14645 = n14117 & ~n14644;
  assign n14646 = ~n14117 & n14644;
  assign n14647 = ~n14645 & ~n14646;
  assign n14648 = ~po45  & n14641;
  assign n14649 = ~n14647 & ~n14648;
  assign n14650 = ~n14642 & ~n14649;
  assign n14651 = po46  & ~n14650;
  assign n14652 = ~po46  & ~n14642;
  assign n14653 = ~n14649 & n14652;
  assign n14654 = ~n14120 & po9 ;
  assign n14655 = ~n14126 & n14654;
  assign n14656 = n14125 & ~n14655;
  assign n14657 = n14127 & n14654;
  assign n14658 = ~n14656 & ~n14657;
  assign n14659 = ~n14653 & n14658;
  assign n14660 = ~n14651 & ~n14659;
  assign n14661 = po47  & ~n14660;
  assign n14662 = ~n14129 & ~n14131;
  assign n14663 = po9  & n14662;
  assign n14664 = n14136 & ~n14663;
  assign n14665 = ~n14136 & n14663;
  assign n14666 = ~n14664 & ~n14665;
  assign n14667 = ~po47  & n14660;
  assign n14668 = ~n14666 & ~n14667;
  assign n14669 = ~n14661 & ~n14668;
  assign n14670 = po48  & ~n14669;
  assign n14671 = ~n14139 & ~n14140;
  assign n14672 = po9  & n14671;
  assign n14673 = n14145 & ~n14672;
  assign n14674 = ~n14145 & n14672;
  assign n14675 = ~n14673 & ~n14674;
  assign n14676 = ~po48  & ~n14661;
  assign n14677 = ~n14668 & n14676;
  assign n14678 = ~n14675 & ~n14677;
  assign n14679 = ~n14670 & ~n14678;
  assign n14680 = po49  & ~n14679;
  assign n14681 = ~n14148 & ~n14150;
  assign n14682 = po9  & n14681;
  assign n14683 = n14155 & ~n14682;
  assign n14684 = ~n14155 & n14682;
  assign n14685 = ~n14683 & ~n14684;
  assign n14686 = ~po49  & n14679;
  assign n14687 = ~n14685 & ~n14686;
  assign n14688 = ~n14680 & ~n14687;
  assign n14689 = po50  & ~n14688;
  assign n14690 = ~po50  & ~n14680;
  assign n14691 = ~n14687 & n14690;
  assign n14692 = ~n14158 & po9 ;
  assign n14693 = ~n14164 & n14692;
  assign n14694 = n14163 & ~n14693;
  assign n14695 = n14165 & n14692;
  assign n14696 = ~n14694 & ~n14695;
  assign n14697 = ~n14691 & n14696;
  assign n14698 = ~n14689 & ~n14697;
  assign n14699 = po51  & ~n14698;
  assign n14700 = ~n14167 & ~n14169;
  assign n14701 = po9  & n14700;
  assign n14702 = n14174 & ~n14701;
  assign n14703 = ~n14174 & n14701;
  assign n14704 = ~n14702 & ~n14703;
  assign n14705 = ~po51  & n14698;
  assign n14706 = ~n14704 & ~n14705;
  assign n14707 = ~n14699 & ~n14706;
  assign n14708 = po52  & ~n14707;
  assign n14709 = ~n14177 & ~n14178;
  assign n14710 = po9  & n14709;
  assign n14711 = n14183 & ~n14710;
  assign n14712 = ~n14183 & n14710;
  assign n14713 = ~n14711 & ~n14712;
  assign n14714 = ~po52  & ~n14699;
  assign n14715 = ~n14706 & n14714;
  assign n14716 = ~n14713 & ~n14715;
  assign n14717 = ~n14708 & ~n14716;
  assign n14718 = ~po53  & n14717;
  assign n14719 = ~n14186 & po9 ;
  assign n14720 = ~n14193 & n14719;
  assign n14721 = n14191 & ~n14720;
  assign n14722 = n14194 & n14719;
  assign n14723 = ~n14721 & ~n14722;
  assign n14724 = ~n14718 & n14723;
  assign n14725 = po53  & ~n14717;
  assign n14726 = ~n14724 & ~n14725;
  assign n14727 = po54  & ~n14726;
  assign n14728 = ~n14196 & ~n14203;
  assign n14729 = po9  & n14728;
  assign n14730 = ~n14201 & ~n14729;
  assign n14731 = n14201 & n14729;
  assign n14732 = ~n14730 & ~n14731;
  assign n14733 = ~po54  & ~n14725;
  assign n14734 = ~n14724 & n14733;
  assign n14735 = n14732 & ~n14734;
  assign n14736 = ~n14727 & ~n14735;
  assign n14737 = ~po55  & n14736;
  assign n14738 = po55  & ~n14736;
  assign n14739 = ~n14306 & ~n14737;
  assign n14740 = ~n14738 & ~n14739;
  assign n14741 = po56  & ~n14740;
  assign n14742 = ~po56  & ~n14738;
  assign n14743 = ~n14739 & n14742;
  assign n14744 = ~n14210 & po9 ;
  assign n14745 = ~n14216 & n14744;
  assign n14746 = n14215 & ~n14745;
  assign n14747 = n14217 & n14744;
  assign n14748 = ~n14746 & ~n14747;
  assign n14749 = ~n14743 & n14748;
  assign n14750 = ~n14741 & ~n14749;
  assign n14751 = po57  & ~n14750;
  assign n14752 = ~n14219 & ~n14221;
  assign n14753 = po9  & n14752;
  assign n14754 = n14226 & ~n14753;
  assign n14755 = ~n14226 & n14753;
  assign n14756 = ~n14754 & ~n14755;
  assign n14757 = ~po57  & n14750;
  assign n14758 = ~n14756 & ~n14757;
  assign n14759 = ~n14751 & ~n14758;
  assign n14760 = po58  & ~n14759;
  assign n14761 = ~po58  & ~n14751;
  assign n14762 = ~n14758 & n14761;
  assign n14763 = ~n14229 & po9 ;
  assign n14764 = ~n14235 & n14763;
  assign n14765 = n14234 & ~n14764;
  assign n14766 = n14236 & n14763;
  assign n14767 = ~n14765 & ~n14766;
  assign n14768 = ~n14762 & n14767;
  assign n14769 = ~n14760 & ~n14768;
  assign n14770 = po59  & ~n14769;
  assign n14771 = ~n14238 & ~n14240;
  assign n14772 = po9  & n14771;
  assign n14773 = n14245 & ~n14772;
  assign n14774 = ~n14245 & n14772;
  assign n14775 = ~n14773 & ~n14774;
  assign n14776 = ~po59  & n14769;
  assign n14777 = ~n14775 & ~n14776;
  assign n14778 = ~n14770 & ~n14777;
  assign n14779 = po60  & ~n14778;
  assign n14780 = ~n14248 & ~n14249;
  assign n14781 = po9  & n14780;
  assign n14782 = n14254 & ~n14781;
  assign n14783 = ~n14254 & n14781;
  assign n14784 = ~n14782 & ~n14783;
  assign n14785 = ~po60  & ~n14770;
  assign n14786 = ~n14777 & n14785;
  assign n14787 = ~n14784 & ~n14786;
  assign n14788 = ~n14779 & ~n14787;
  assign n14789 = po61  & ~n14788;
  assign n14790 = ~n14257 & ~n14259;
  assign n14791 = po9  & n14790;
  assign n14792 = n14264 & ~n14791;
  assign n14793 = ~n14264 & n14791;
  assign n14794 = ~n14792 & ~n14793;
  assign n14795 = ~po61  & n14788;
  assign n14796 = ~n14794 & ~n14795;
  assign n14797 = ~n14789 & ~n14796;
  assign n14798 = po62  & ~n14797;
  assign n14799 = ~po62  & ~n14789;
  assign n14800 = ~n14796 & n14799;
  assign n14801 = ~n14267 & po9 ;
  assign n14802 = ~n14273 & n14801;
  assign n14803 = n14272 & ~n14802;
  assign n14804 = n14274 & n14801;
  assign n14805 = ~n14803 & ~n14804;
  assign n14806 = ~n14800 & n14805;
  assign n14807 = ~n14798 & ~n14806;
  assign n14808 = n14294 & po9 ;
  assign n14809 = ~n14285 & n14808;
  assign n14810 = ~n14276 & ~n14278;
  assign n14811 = po9  & n14810;
  assign n14812 = n14283 & ~n14811;
  assign n14813 = ~n14283 & n14811;
  assign n14814 = ~n14812 & ~n14813;
  assign n14815 = ~n14298 & ~n14809;
  assign n14816 = ~n14814 & n14815;
  assign n14817 = ~n14807 & n14816;
  assign n14818 = ~po63  & ~n14817;
  assign n14819 = n14807 & n14814;
  assign n14820 = n14285 & ~n14808;
  assign n14821 = ~n14285 & n14294;
  assign n14822 = po63  & ~n14821;
  assign n14823 = ~n14820 & n14822;
  assign n14824 = ~n14819 & ~n14823;
  assign po8  = n14818 | ~n14824;
  assign n14826 = ~n14738 & po8 ;
  assign n14827 = ~n14737 & n14826;
  assign n14828 = n14306 & ~n14827;
  assign n14829 = n14739 & n14826;
  assign n14830 = ~n14828 & ~n14829;
  assign n14831 = ~n14727 & ~n14734;
  assign n14832 = po8  & n14831;
  assign n14833 = n14732 & ~n14832;
  assign n14834 = ~n14732 & n14832;
  assign n14835 = ~n14833 & ~n14834;
  assign n14836 = pi16  & po8 ;
  assign n14837 = ~pi14  & ~pi15 ;
  assign n14838 = ~pi16  & n14837;
  assign n14839 = ~n14836 & ~n14838;
  assign n14840 = po9  & ~n14839;
  assign n14841 = ~pi16  & po8 ;
  assign n14842 = pi17  & ~n14841;
  assign n14843 = ~pi17  & n14841;
  assign n14844 = ~n14842 & ~n14843;
  assign n14845 = ~po9  & n14839;
  assign n14846 = n14844 & ~n14845;
  assign n14847 = ~n14840 & ~n14846;
  assign n14848 = po10  & ~n14847;
  assign n14849 = ~po10  & ~n14840;
  assign n14850 = ~n14846 & n14849;
  assign n14851 = po9  & ~po8 ;
  assign n14852 = ~n14843 & ~n14851;
  assign n14853 = pi18  & ~n14852;
  assign n14854 = ~pi18  & n14852;
  assign n14855 = ~n14853 & ~n14854;
  assign n14856 = ~n14850 & ~n14855;
  assign n14857 = ~n14848 & ~n14856;
  assign n14858 = po11  & ~n14857;
  assign n14859 = ~po11  & n14857;
  assign n14860 = ~n14311 & ~n14312;
  assign n14861 = po8  & n14860;
  assign n14862 = n14316 & ~n14861;
  assign n14863 = ~n14316 & n14861;
  assign n14864 = ~n14862 & ~n14863;
  assign n14865 = ~n14859 & ~n14864;
  assign n14866 = ~n14858 & ~n14865;
  assign n14867 = po12  & ~n14866;
  assign n14868 = ~po12  & ~n14858;
  assign n14869 = ~n14865 & n14868;
  assign n14870 = ~n14319 & po8 ;
  assign n14871 = ~n14325 & n14870;
  assign n14872 = n14324 & ~n14871;
  assign n14873 = n14326 & n14870;
  assign n14874 = ~n14872 & ~n14873;
  assign n14875 = ~n14869 & n14874;
  assign n14876 = ~n14867 & ~n14875;
  assign n14877 = po13  & ~n14876;
  assign n14878 = ~po13  & n14876;
  assign n14879 = ~n14328 & ~n14330;
  assign n14880 = po8  & n14879;
  assign n14881 = n14335 & ~n14880;
  assign n14882 = ~n14335 & n14880;
  assign n14883 = ~n14881 & ~n14882;
  assign n14884 = ~n14878 & n14883;
  assign n14885 = ~n14877 & ~n14884;
  assign n14886 = po14  & ~n14885;
  assign n14887 = ~po14  & ~n14877;
  assign n14888 = ~n14884 & n14887;
  assign n14889 = ~n14338 & po8 ;
  assign n14890 = ~n14344 & n14889;
  assign n14891 = n14343 & ~n14890;
  assign n14892 = n14345 & n14889;
  assign n14893 = ~n14891 & ~n14892;
  assign n14894 = ~n14888 & n14893;
  assign n14895 = ~n14886 & ~n14894;
  assign n14896 = po15  & ~n14895;
  assign n14897 = ~po15  & n14895;
  assign n14898 = ~n14347 & ~n14349;
  assign n14899 = po8  & n14898;
  assign n14900 = n14354 & n14899;
  assign n14901 = ~n14354 & ~n14899;
  assign n14902 = ~n14900 & ~n14901;
  assign n14903 = ~n14897 & n14902;
  assign n14904 = ~n14896 & ~n14903;
  assign n14905 = po16  & ~n14904;
  assign n14906 = ~po16  & ~n14896;
  assign n14907 = ~n14903 & n14906;
  assign n14908 = ~n14357 & po8 ;
  assign n14909 = ~n14363 & n14908;
  assign n14910 = n14362 & ~n14909;
  assign n14911 = n14364 & n14908;
  assign n14912 = ~n14910 & ~n14911;
  assign n14913 = ~n14907 & n14912;
  assign n14914 = ~n14905 & ~n14913;
  assign n14915 = po17  & ~n14914;
  assign n14916 = ~po17  & n14914;
  assign n14917 = ~n14366 & ~n14368;
  assign n14918 = po8  & n14917;
  assign n14919 = ~n14373 & ~n14918;
  assign n14920 = n14373 & n14918;
  assign n14921 = ~n14919 & ~n14920;
  assign n14922 = ~n14916 & n14921;
  assign n14923 = ~n14915 & ~n14922;
  assign n14924 = po18  & ~n14923;
  assign n14925 = ~po18  & ~n14915;
  assign n14926 = ~n14922 & n14925;
  assign n14927 = ~n14376 & po8 ;
  assign n14928 = ~n14382 & n14927;
  assign n14929 = n14381 & ~n14928;
  assign n14930 = n14383 & n14927;
  assign n14931 = ~n14929 & ~n14930;
  assign n14932 = ~n14926 & n14931;
  assign n14933 = ~n14924 & ~n14932;
  assign n14934 = po19  & ~n14933;
  assign n14935 = ~n14385 & ~n14387;
  assign n14936 = po8  & n14935;
  assign n14937 = n14392 & ~n14936;
  assign n14938 = ~n14392 & n14936;
  assign n14939 = ~n14937 & ~n14938;
  assign n14940 = ~po19  & n14933;
  assign n14941 = ~n14939 & ~n14940;
  assign n14942 = ~n14934 & ~n14941;
  assign n14943 = po20  & ~n14942;
  assign n14944 = ~po20  & ~n14934;
  assign n14945 = ~n14941 & n14944;
  assign n14946 = ~n14395 & po8 ;
  assign n14947 = ~n14401 & n14946;
  assign n14948 = n14400 & ~n14947;
  assign n14949 = n14402 & n14946;
  assign n14950 = ~n14948 & ~n14949;
  assign n14951 = ~n14945 & n14950;
  assign n14952 = ~n14943 & ~n14951;
  assign n14953 = po21  & ~n14952;
  assign n14954 = ~po21  & n14952;
  assign n14955 = ~n14404 & po8 ;
  assign n14956 = ~n14411 & n14955;
  assign n14957 = n14409 & ~n14956;
  assign n14958 = n14412 & n14955;
  assign n14959 = ~n14957 & ~n14958;
  assign n14960 = ~n14954 & n14959;
  assign n14961 = ~n14953 & ~n14960;
  assign n14962 = po22  & ~n14961;
  assign n14963 = ~po22  & ~n14953;
  assign n14964 = ~n14960 & n14963;
  assign n14965 = ~n14414 & po8 ;
  assign n14966 = ~n14420 & n14965;
  assign n14967 = n14419 & ~n14966;
  assign n14968 = n14421 & n14965;
  assign n14969 = ~n14967 & ~n14968;
  assign n14970 = ~n14964 & n14969;
  assign n14971 = ~n14962 & ~n14970;
  assign n14972 = po23  & ~n14971;
  assign n14973 = ~n14423 & ~n14425;
  assign n14974 = po8  & n14973;
  assign n14975 = n14430 & ~n14974;
  assign n14976 = ~n14430 & n14974;
  assign n14977 = ~n14975 & ~n14976;
  assign n14978 = ~po23  & n14971;
  assign n14979 = ~n14977 & ~n14978;
  assign n14980 = ~n14972 & ~n14979;
  assign n14981 = po24  & ~n14980;
  assign n14982 = ~po24  & ~n14972;
  assign n14983 = ~n14979 & n14982;
  assign n14984 = ~n14433 & po8 ;
  assign n14985 = ~n14439 & n14984;
  assign n14986 = n14438 & ~n14985;
  assign n14987 = n14440 & n14984;
  assign n14988 = ~n14986 & ~n14987;
  assign n14989 = ~n14983 & n14988;
  assign n14990 = ~n14981 & ~n14989;
  assign n14991 = po25  & ~n14990;
  assign n14992 = ~po25  & n14990;
  assign n14993 = ~n14442 & po8 ;
  assign n14994 = ~n14449 & n14993;
  assign n14995 = n14447 & ~n14994;
  assign n14996 = n14450 & n14993;
  assign n14997 = ~n14995 & ~n14996;
  assign n14998 = ~n14992 & n14997;
  assign n14999 = ~n14991 & ~n14998;
  assign n15000 = po26  & ~n14999;
  assign n15001 = ~po26  & ~n14991;
  assign n15002 = ~n14998 & n15001;
  assign n15003 = ~n14452 & po8 ;
  assign n15004 = ~n14458 & n15003;
  assign n15005 = n14457 & ~n15004;
  assign n15006 = n14459 & n15003;
  assign n15007 = ~n15005 & ~n15006;
  assign n15008 = ~n15002 & n15007;
  assign n15009 = ~n15000 & ~n15008;
  assign n15010 = po27  & ~n15009;
  assign n15011 = ~n14461 & ~n14463;
  assign n15012 = po8  & n15011;
  assign n15013 = n14468 & ~n15012;
  assign n15014 = ~n14468 & n15012;
  assign n15015 = ~n15013 & ~n15014;
  assign n15016 = ~po27  & n15009;
  assign n15017 = ~n15015 & ~n15016;
  assign n15018 = ~n15010 & ~n15017;
  assign n15019 = po28  & ~n15018;
  assign n15020 = ~po28  & ~n15010;
  assign n15021 = ~n15017 & n15020;
  assign n15022 = ~n14471 & po8 ;
  assign n15023 = ~n14477 & n15022;
  assign n15024 = n14476 & ~n15023;
  assign n15025 = n14478 & n15022;
  assign n15026 = ~n15024 & ~n15025;
  assign n15027 = ~n15021 & n15026;
  assign n15028 = ~n15019 & ~n15027;
  assign n15029 = po29  & ~n15028;
  assign n15030 = ~po29  & n15028;
  assign n15031 = ~n14480 & po8 ;
  assign n15032 = ~n14487 & n15031;
  assign n15033 = n14485 & ~n15032;
  assign n15034 = n14488 & n15031;
  assign n15035 = ~n15033 & ~n15034;
  assign n15036 = ~n15030 & n15035;
  assign n15037 = ~n15029 & ~n15036;
  assign n15038 = po30  & ~n15037;
  assign n15039 = ~po30  & ~n15029;
  assign n15040 = ~n15036 & n15039;
  assign n15041 = ~n14490 & po8 ;
  assign n15042 = ~n14496 & n15041;
  assign n15043 = n14495 & ~n15042;
  assign n15044 = n14497 & n15041;
  assign n15045 = ~n15043 & ~n15044;
  assign n15046 = ~n15040 & n15045;
  assign n15047 = ~n15038 & ~n15046;
  assign n15048 = po31  & ~n15047;
  assign n15049 = ~n14499 & ~n14501;
  assign n15050 = po8  & n15049;
  assign n15051 = n14506 & ~n15050;
  assign n15052 = ~n14506 & n15050;
  assign n15053 = ~n15051 & ~n15052;
  assign n15054 = ~po31  & n15047;
  assign n15055 = ~n15053 & ~n15054;
  assign n15056 = ~n15048 & ~n15055;
  assign n15057 = po32  & ~n15056;
  assign n15058 = ~po32  & ~n15048;
  assign n15059 = ~n15055 & n15058;
  assign n15060 = ~n14509 & po8 ;
  assign n15061 = ~n14515 & n15060;
  assign n15062 = n14514 & ~n15061;
  assign n15063 = n14516 & n15060;
  assign n15064 = ~n15062 & ~n15063;
  assign n15065 = ~n15059 & n15064;
  assign n15066 = ~n15057 & ~n15065;
  assign n15067 = po33  & ~n15066;
  assign n15068 = ~po33  & n15066;
  assign n15069 = ~n14518 & po8 ;
  assign n15070 = ~n14525 & n15069;
  assign n15071 = n14523 & ~n15070;
  assign n15072 = n14526 & n15069;
  assign n15073 = ~n15071 & ~n15072;
  assign n15074 = ~n15068 & n15073;
  assign n15075 = ~n15067 & ~n15074;
  assign n15076 = po34  & ~n15075;
  assign n15077 = ~po34  & ~n15067;
  assign n15078 = ~n15074 & n15077;
  assign n15079 = ~n14528 & po8 ;
  assign n15080 = ~n14534 & n15079;
  assign n15081 = n14533 & ~n15080;
  assign n15082 = n14535 & n15079;
  assign n15083 = ~n15081 & ~n15082;
  assign n15084 = ~n15078 & n15083;
  assign n15085 = ~n15076 & ~n15084;
  assign n15086 = po35  & ~n15085;
  assign n15087 = ~n14537 & ~n14539;
  assign n15088 = po8  & n15087;
  assign n15089 = n14544 & ~n15088;
  assign n15090 = ~n14544 & n15088;
  assign n15091 = ~n15089 & ~n15090;
  assign n15092 = ~po35  & n15085;
  assign n15093 = ~n15091 & ~n15092;
  assign n15094 = ~n15086 & ~n15093;
  assign n15095 = po36  & ~n15094;
  assign n15096 = ~po36  & ~n15086;
  assign n15097 = ~n15093 & n15096;
  assign n15098 = ~n14547 & po8 ;
  assign n15099 = ~n14553 & n15098;
  assign n15100 = n14552 & ~n15099;
  assign n15101 = n14554 & n15098;
  assign n15102 = ~n15100 & ~n15101;
  assign n15103 = ~n15097 & n15102;
  assign n15104 = ~n15095 & ~n15103;
  assign n15105 = po37  & ~n15104;
  assign n15106 = ~po37  & n15104;
  assign n15107 = ~n14556 & po8 ;
  assign n15108 = ~n14563 & n15107;
  assign n15109 = n14561 & ~n15108;
  assign n15110 = n14564 & n15107;
  assign n15111 = ~n15109 & ~n15110;
  assign n15112 = ~n15106 & n15111;
  assign n15113 = ~n15105 & ~n15112;
  assign n15114 = po38  & ~n15113;
  assign n15115 = ~po38  & ~n15105;
  assign n15116 = ~n15112 & n15115;
  assign n15117 = ~n14566 & po8 ;
  assign n15118 = ~n14572 & n15117;
  assign n15119 = n14571 & ~n15118;
  assign n15120 = n14573 & n15117;
  assign n15121 = ~n15119 & ~n15120;
  assign n15122 = ~n15116 & n15121;
  assign n15123 = ~n15114 & ~n15122;
  assign n15124 = po39  & ~n15123;
  assign n15125 = ~n14575 & ~n14577;
  assign n15126 = po8  & n15125;
  assign n15127 = n14582 & ~n15126;
  assign n15128 = ~n14582 & n15126;
  assign n15129 = ~n15127 & ~n15128;
  assign n15130 = ~po39  & n15123;
  assign n15131 = ~n15129 & ~n15130;
  assign n15132 = ~n15124 & ~n15131;
  assign n15133 = po40  & ~n15132;
  assign n15134 = ~po40  & ~n15124;
  assign n15135 = ~n15131 & n15134;
  assign n15136 = ~n14585 & po8 ;
  assign n15137 = ~n14591 & n15136;
  assign n15138 = n14590 & ~n15137;
  assign n15139 = n14592 & n15136;
  assign n15140 = ~n15138 & ~n15139;
  assign n15141 = ~n15135 & n15140;
  assign n15142 = ~n15133 & ~n15141;
  assign n15143 = po41  & ~n15142;
  assign n15144 = ~po41  & n15142;
  assign n15145 = ~n14594 & po8 ;
  assign n15146 = ~n14601 & n15145;
  assign n15147 = n14599 & ~n15146;
  assign n15148 = n14602 & n15145;
  assign n15149 = ~n15147 & ~n15148;
  assign n15150 = ~n15144 & n15149;
  assign n15151 = ~n15143 & ~n15150;
  assign n15152 = po42  & ~n15151;
  assign n15153 = ~po42  & ~n15143;
  assign n15154 = ~n15150 & n15153;
  assign n15155 = ~n14604 & po8 ;
  assign n15156 = ~n14610 & n15155;
  assign n15157 = n14609 & ~n15156;
  assign n15158 = n14611 & n15155;
  assign n15159 = ~n15157 & ~n15158;
  assign n15160 = ~n15154 & n15159;
  assign n15161 = ~n15152 & ~n15160;
  assign n15162 = po43  & ~n15161;
  assign n15163 = ~n14613 & ~n14615;
  assign n15164 = po8  & n15163;
  assign n15165 = n14620 & ~n15164;
  assign n15166 = ~n14620 & n15164;
  assign n15167 = ~n15165 & ~n15166;
  assign n15168 = ~po43  & n15161;
  assign n15169 = ~n15167 & ~n15168;
  assign n15170 = ~n15162 & ~n15169;
  assign n15171 = po44  & ~n15170;
  assign n15172 = ~po44  & ~n15162;
  assign n15173 = ~n15169 & n15172;
  assign n15174 = ~n14623 & po8 ;
  assign n15175 = ~n14629 & n15174;
  assign n15176 = n14628 & ~n15175;
  assign n15177 = n14630 & n15174;
  assign n15178 = ~n15176 & ~n15177;
  assign n15179 = ~n15173 & n15178;
  assign n15180 = ~n15171 & ~n15179;
  assign n15181 = po45  & ~n15180;
  assign n15182 = ~po45  & n15180;
  assign n15183 = ~n14632 & po8 ;
  assign n15184 = ~n14639 & n15183;
  assign n15185 = n14637 & ~n15184;
  assign n15186 = n14640 & n15183;
  assign n15187 = ~n15185 & ~n15186;
  assign n15188 = ~n15182 & n15187;
  assign n15189 = ~n15181 & ~n15188;
  assign n15190 = po46  & ~n15189;
  assign n15191 = ~po46  & ~n15181;
  assign n15192 = ~n15188 & n15191;
  assign n15193 = ~n14642 & po8 ;
  assign n15194 = ~n14648 & n15193;
  assign n15195 = n14647 & ~n15194;
  assign n15196 = n14649 & n15193;
  assign n15197 = ~n15195 & ~n15196;
  assign n15198 = ~n15192 & n15197;
  assign n15199 = ~n15190 & ~n15198;
  assign n15200 = po47  & ~n15199;
  assign n15201 = ~n14651 & ~n14653;
  assign n15202 = po8  & n15201;
  assign n15203 = n14658 & ~n15202;
  assign n15204 = ~n14658 & n15202;
  assign n15205 = ~n15203 & ~n15204;
  assign n15206 = ~po47  & n15199;
  assign n15207 = ~n15205 & ~n15206;
  assign n15208 = ~n15200 & ~n15207;
  assign n15209 = po48  & ~n15208;
  assign n15210 = ~po48  & ~n15200;
  assign n15211 = ~n15207 & n15210;
  assign n15212 = ~n14661 & po8 ;
  assign n15213 = ~n14667 & n15212;
  assign n15214 = n14666 & ~n15213;
  assign n15215 = n14668 & n15212;
  assign n15216 = ~n15214 & ~n15215;
  assign n15217 = ~n15211 & n15216;
  assign n15218 = ~n15209 & ~n15217;
  assign n15219 = po49  & ~n15218;
  assign n15220 = ~po49  & n15218;
  assign n15221 = ~n14670 & po8 ;
  assign n15222 = ~n14677 & n15221;
  assign n15223 = n14675 & ~n15222;
  assign n15224 = n14678 & n15221;
  assign n15225 = ~n15223 & ~n15224;
  assign n15226 = ~n15220 & n15225;
  assign n15227 = ~n15219 & ~n15226;
  assign n15228 = po50  & ~n15227;
  assign n15229 = ~po50  & ~n15219;
  assign n15230 = ~n15226 & n15229;
  assign n15231 = ~n14680 & po8 ;
  assign n15232 = ~n14686 & n15231;
  assign n15233 = n14685 & ~n15232;
  assign n15234 = n14687 & n15231;
  assign n15235 = ~n15233 & ~n15234;
  assign n15236 = ~n15230 & n15235;
  assign n15237 = ~n15228 & ~n15236;
  assign n15238 = po51  & ~n15237;
  assign n15239 = ~n14689 & ~n14691;
  assign n15240 = po8  & n15239;
  assign n15241 = n14696 & ~n15240;
  assign n15242 = ~n14696 & n15240;
  assign n15243 = ~n15241 & ~n15242;
  assign n15244 = ~po51  & n15237;
  assign n15245 = ~n15243 & ~n15244;
  assign n15246 = ~n15238 & ~n15245;
  assign n15247 = po52  & ~n15246;
  assign n15248 = ~po52  & ~n15238;
  assign n15249 = ~n15245 & n15248;
  assign n15250 = ~n14699 & po8 ;
  assign n15251 = ~n14705 & n15250;
  assign n15252 = n14704 & ~n15251;
  assign n15253 = n14706 & n15250;
  assign n15254 = ~n15252 & ~n15253;
  assign n15255 = ~n15249 & n15254;
  assign n15256 = ~n15247 & ~n15255;
  assign n15257 = po53  & ~n15256;
  assign n15258 = ~po53  & n15256;
  assign n15259 = ~n14708 & po8 ;
  assign n15260 = ~n14715 & n15259;
  assign n15261 = n14713 & ~n15260;
  assign n15262 = n14716 & n15259;
  assign n15263 = ~n15261 & ~n15262;
  assign n15264 = ~n15258 & n15263;
  assign n15265 = ~n15257 & ~n15264;
  assign n15266 = po54  & ~n15265;
  assign n15267 = ~n14718 & ~n14725;
  assign n15268 = po8  & n15267;
  assign n15269 = n14723 & ~n15268;
  assign n15270 = ~n14723 & n15268;
  assign n15271 = ~n15269 & ~n15270;
  assign n15272 = ~po54  & ~n15257;
  assign n15273 = ~n15264 & n15272;
  assign n15274 = ~n15271 & ~n15273;
  assign n15275 = ~n15266 & ~n15274;
  assign n15276 = ~po55  & n15275;
  assign n15277 = ~n14835 & ~n15276;
  assign n15278 = po55  & ~n15275;
  assign n15279 = ~po56  & ~n15278;
  assign n15280 = ~n15277 & n15279;
  assign n15281 = ~n15277 & ~n15278;
  assign n15282 = po56  & ~n15281;
  assign n15283 = n14830 & ~n15280;
  assign n15284 = ~n15282 & ~n15283;
  assign n15285 = po57  & ~n15284;
  assign n15286 = ~n14741 & ~n14743;
  assign n15287 = po8  & n15286;
  assign n15288 = n14748 & ~n15287;
  assign n15289 = ~n14748 & n15287;
  assign n15290 = ~n15288 & ~n15289;
  assign n15291 = ~po57  & n15284;
  assign n15292 = ~n15290 & ~n15291;
  assign n15293 = ~n15285 & ~n15292;
  assign n15294 = po58  & ~n15293;
  assign n15295 = ~po58  & ~n15285;
  assign n15296 = ~n15292 & n15295;
  assign n15297 = ~n14751 & po8 ;
  assign n15298 = ~n14757 & n15297;
  assign n15299 = n14756 & ~n15298;
  assign n15300 = n14758 & n15297;
  assign n15301 = ~n15299 & ~n15300;
  assign n15302 = ~n15296 & n15301;
  assign n15303 = ~n15294 & ~n15302;
  assign n15304 = po59  & ~n15303;
  assign n15305 = ~n14760 & ~n14762;
  assign n15306 = po8  & n15305;
  assign n15307 = n14767 & ~n15306;
  assign n15308 = ~n14767 & n15306;
  assign n15309 = ~n15307 & ~n15308;
  assign n15310 = ~po59  & n15303;
  assign n15311 = ~n15309 & ~n15310;
  assign n15312 = ~n15304 & ~n15311;
  assign n15313 = po60  & ~n15312;
  assign n15314 = ~po60  & ~n15304;
  assign n15315 = ~n15311 & n15314;
  assign n15316 = ~n14770 & po8 ;
  assign n15317 = ~n14776 & n15316;
  assign n15318 = n14775 & ~n15317;
  assign n15319 = n14777 & n15316;
  assign n15320 = ~n15318 & ~n15319;
  assign n15321 = ~n15315 & n15320;
  assign n15322 = ~n15313 & ~n15321;
  assign n15323 = po61  & ~n15322;
  assign n15324 = ~po61  & n15322;
  assign n15325 = ~n14779 & po8 ;
  assign n15326 = ~n14786 & n15325;
  assign n15327 = n14784 & ~n15326;
  assign n15328 = n14787 & n15325;
  assign n15329 = ~n15327 & ~n15328;
  assign n15330 = ~n15324 & n15329;
  assign n15331 = ~n15323 & ~n15330;
  assign n15332 = po62  & ~n15331;
  assign n15333 = ~po62  & ~n15323;
  assign n15334 = ~n15330 & n15333;
  assign n15335 = ~n14789 & po8 ;
  assign n15336 = ~n14795 & n15335;
  assign n15337 = n14794 & ~n15336;
  assign n15338 = n14796 & n15335;
  assign n15339 = ~n15337 & ~n15338;
  assign n15340 = ~n15334 & n15339;
  assign n15341 = ~n15332 & ~n15340;
  assign n15342 = ~n14798 & ~n14800;
  assign n15343 = po8  & n15342;
  assign n15344 = n14805 & ~n15343;
  assign n15345 = ~n14805 & n15343;
  assign n15346 = ~n15344 & ~n15345;
  assign n15347 = n14807 & po8 ;
  assign n15348 = ~n14814 & ~n15347;
  assign n15349 = ~n14819 & ~n15348;
  assign n15350 = po8  & ~n15349;
  assign n15351 = ~n15346 & ~n15350;
  assign n15352 = ~n15341 & n15351;
  assign n15353 = ~po63  & ~n15352;
  assign n15354 = n15341 & n15346;
  assign n15355 = po63  & n15349;
  assign n15356 = ~n15354 & ~n15355;
  assign po7  = n15353 | ~n15356;
  assign n15358 = ~n15280 & ~n15282;
  assign n15359 = po7  & n15358;
  assign n15360 = n14830 & ~n15359;
  assign n15361 = ~n14830 & n15359;
  assign n15362 = ~n15360 & ~n15361;
  assign n15363 = pi14  & po7 ;
  assign n15364 = ~pi12  & ~pi13 ;
  assign n15365 = ~pi14  & n15364;
  assign n15366 = ~n15363 & ~n15365;
  assign n15367 = po8  & ~n15366;
  assign n15368 = ~po8  & n15366;
  assign n15369 = ~pi14  & po7 ;
  assign n15370 = pi15  & ~n15369;
  assign n15371 = ~pi15  & n15369;
  assign n15372 = ~n15370 & ~n15371;
  assign n15373 = ~n15368 & n15372;
  assign n15374 = ~n15367 & ~n15373;
  assign n15375 = po9  & ~n15374;
  assign n15376 = po8  & ~po7 ;
  assign n15377 = ~n15371 & ~n15376;
  assign n15378 = pi16  & ~n15377;
  assign n15379 = ~pi16  & n15377;
  assign n15380 = ~n15378 & ~n15379;
  assign n15381 = ~po9  & n15374;
  assign n15382 = ~n15380 & ~n15381;
  assign n15383 = ~n15375 & ~n15382;
  assign n15384 = po10  & ~n15383;
  assign n15385 = ~po10  & ~n15375;
  assign n15386 = ~n15382 & n15385;
  assign n15387 = ~n14840 & ~n14845;
  assign n15388 = po7  & n15387;
  assign n15389 = n14844 & ~n15388;
  assign n15390 = ~n14844 & n15388;
  assign n15391 = ~n15389 & ~n15390;
  assign n15392 = ~n15386 & ~n15391;
  assign n15393 = ~n15384 & ~n15392;
  assign n15394 = po11  & ~n15393;
  assign n15395 = ~n14848 & ~n14850;
  assign n15396 = po7  & n15395;
  assign n15397 = ~n14855 & ~n15396;
  assign n15398 = n14855 & n15396;
  assign n15399 = ~n15397 & ~n15398;
  assign n15400 = ~po11  & n15393;
  assign n15401 = ~n15399 & ~n15400;
  assign n15402 = ~n15394 & ~n15401;
  assign n15403 = po12  & ~n15402;
  assign n15404 = ~po12  & ~n15394;
  assign n15405 = ~n15401 & n15404;
  assign n15406 = ~n14858 & ~n14859;
  assign n15407 = po7  & n15406;
  assign n15408 = n14864 & ~n15407;
  assign n15409 = ~n14864 & n15407;
  assign n15410 = ~n15408 & ~n15409;
  assign n15411 = ~n15405 & n15410;
  assign n15412 = ~n15403 & ~n15411;
  assign n15413 = po13  & ~n15412;
  assign n15414 = ~n14867 & ~n14869;
  assign n15415 = po7  & n15414;
  assign n15416 = n14874 & ~n15415;
  assign n15417 = ~n14874 & n15415;
  assign n15418 = ~n15416 & ~n15417;
  assign n15419 = ~po13  & n15412;
  assign n15420 = ~n15418 & ~n15419;
  assign n15421 = ~n15413 & ~n15420;
  assign n15422 = po14  & ~n15421;
  assign n15423 = ~po14  & ~n15413;
  assign n15424 = ~n15420 & n15423;
  assign n15425 = ~n14877 & ~n14878;
  assign n15426 = po7  & n15425;
  assign n15427 = n14883 & n15426;
  assign n15428 = ~n14883 & ~n15426;
  assign n15429 = ~n15427 & ~n15428;
  assign n15430 = ~n15424 & n15429;
  assign n15431 = ~n15422 & ~n15430;
  assign n15432 = po15  & ~n15431;
  assign n15433 = ~n14886 & ~n14888;
  assign n15434 = po7  & n15433;
  assign n15435 = n14893 & ~n15434;
  assign n15436 = ~n14893 & n15434;
  assign n15437 = ~n15435 & ~n15436;
  assign n15438 = ~po15  & n15431;
  assign n15439 = ~n15437 & ~n15438;
  assign n15440 = ~n15432 & ~n15439;
  assign n15441 = po16  & ~n15440;
  assign n15442 = ~po16  & ~n15432;
  assign n15443 = ~n15439 & n15442;
  assign n15444 = ~n14896 & ~n14897;
  assign n15445 = po7  & n15444;
  assign n15446 = ~n14902 & ~n15445;
  assign n15447 = n14902 & n15445;
  assign n15448 = ~n15446 & ~n15447;
  assign n15449 = ~n15443 & n15448;
  assign n15450 = ~n15441 & ~n15449;
  assign n15451 = po17  & ~n15450;
  assign n15452 = ~n14905 & ~n14907;
  assign n15453 = po7  & n15452;
  assign n15454 = n14912 & ~n15453;
  assign n15455 = ~n14912 & n15453;
  assign n15456 = ~n15454 & ~n15455;
  assign n15457 = ~po17  & n15450;
  assign n15458 = ~n15456 & ~n15457;
  assign n15459 = ~n15451 & ~n15458;
  assign n15460 = po18  & ~n15459;
  assign n15461 = ~n14915 & ~n14916;
  assign n15462 = po7  & n15461;
  assign n15463 = n14921 & ~n15462;
  assign n15464 = ~n14921 & n15462;
  assign n15465 = ~n15463 & ~n15464;
  assign n15466 = ~po18  & ~n15451;
  assign n15467 = ~n15458 & n15466;
  assign n15468 = ~n15465 & ~n15467;
  assign n15469 = ~n15460 & ~n15468;
  assign n15470 = po19  & ~n15469;
  assign n15471 = ~n14924 & ~n14926;
  assign n15472 = po7  & n15471;
  assign n15473 = n14931 & ~n15472;
  assign n15474 = ~n14931 & n15472;
  assign n15475 = ~n15473 & ~n15474;
  assign n15476 = ~po19  & n15469;
  assign n15477 = ~n15475 & ~n15476;
  assign n15478 = ~n15470 & ~n15477;
  assign n15479 = po20  & ~n15478;
  assign n15480 = ~po20  & ~n15470;
  assign n15481 = ~n15477 & n15480;
  assign n15482 = ~n14934 & po7 ;
  assign n15483 = ~n14940 & n15482;
  assign n15484 = n14939 & ~n15483;
  assign n15485 = n14941 & n15482;
  assign n15486 = ~n15484 & ~n15485;
  assign n15487 = ~n15481 & n15486;
  assign n15488 = ~n15479 & ~n15487;
  assign n15489 = po21  & ~n15488;
  assign n15490 = ~n14943 & ~n14945;
  assign n15491 = po7  & n15490;
  assign n15492 = n14950 & ~n15491;
  assign n15493 = ~n14950 & n15491;
  assign n15494 = ~n15492 & ~n15493;
  assign n15495 = ~po21  & n15488;
  assign n15496 = ~n15494 & ~n15495;
  assign n15497 = ~n15489 & ~n15496;
  assign n15498 = po22  & ~n15497;
  assign n15499 = ~n14953 & ~n14954;
  assign n15500 = po7  & n15499;
  assign n15501 = n14959 & ~n15500;
  assign n15502 = ~n14959 & n15500;
  assign n15503 = ~n15501 & ~n15502;
  assign n15504 = ~po22  & ~n15489;
  assign n15505 = ~n15496 & n15504;
  assign n15506 = ~n15503 & ~n15505;
  assign n15507 = ~n15498 & ~n15506;
  assign n15508 = po23  & ~n15507;
  assign n15509 = ~n14962 & ~n14964;
  assign n15510 = po7  & n15509;
  assign n15511 = n14969 & ~n15510;
  assign n15512 = ~n14969 & n15510;
  assign n15513 = ~n15511 & ~n15512;
  assign n15514 = ~po23  & n15507;
  assign n15515 = ~n15513 & ~n15514;
  assign n15516 = ~n15508 & ~n15515;
  assign n15517 = po24  & ~n15516;
  assign n15518 = ~po24  & ~n15508;
  assign n15519 = ~n15515 & n15518;
  assign n15520 = ~n14972 & po7 ;
  assign n15521 = ~n14978 & n15520;
  assign n15522 = n14977 & ~n15521;
  assign n15523 = n14979 & n15520;
  assign n15524 = ~n15522 & ~n15523;
  assign n15525 = ~n15519 & n15524;
  assign n15526 = ~n15517 & ~n15525;
  assign n15527 = po25  & ~n15526;
  assign n15528 = ~n14981 & ~n14983;
  assign n15529 = po7  & n15528;
  assign n15530 = n14988 & ~n15529;
  assign n15531 = ~n14988 & n15529;
  assign n15532 = ~n15530 & ~n15531;
  assign n15533 = ~po25  & n15526;
  assign n15534 = ~n15532 & ~n15533;
  assign n15535 = ~n15527 & ~n15534;
  assign n15536 = po26  & ~n15535;
  assign n15537 = ~n14991 & ~n14992;
  assign n15538 = po7  & n15537;
  assign n15539 = n14997 & ~n15538;
  assign n15540 = ~n14997 & n15538;
  assign n15541 = ~n15539 & ~n15540;
  assign n15542 = ~po26  & ~n15527;
  assign n15543 = ~n15534 & n15542;
  assign n15544 = ~n15541 & ~n15543;
  assign n15545 = ~n15536 & ~n15544;
  assign n15546 = po27  & ~n15545;
  assign n15547 = ~n15000 & ~n15002;
  assign n15548 = po7  & n15547;
  assign n15549 = n15007 & ~n15548;
  assign n15550 = ~n15007 & n15548;
  assign n15551 = ~n15549 & ~n15550;
  assign n15552 = ~po27  & n15545;
  assign n15553 = ~n15551 & ~n15552;
  assign n15554 = ~n15546 & ~n15553;
  assign n15555 = po28  & ~n15554;
  assign n15556 = ~po28  & ~n15546;
  assign n15557 = ~n15553 & n15556;
  assign n15558 = ~n15010 & po7 ;
  assign n15559 = ~n15016 & n15558;
  assign n15560 = n15015 & ~n15559;
  assign n15561 = n15017 & n15558;
  assign n15562 = ~n15560 & ~n15561;
  assign n15563 = ~n15557 & n15562;
  assign n15564 = ~n15555 & ~n15563;
  assign n15565 = po29  & ~n15564;
  assign n15566 = ~n15019 & ~n15021;
  assign n15567 = po7  & n15566;
  assign n15568 = n15026 & ~n15567;
  assign n15569 = ~n15026 & n15567;
  assign n15570 = ~n15568 & ~n15569;
  assign n15571 = ~po29  & n15564;
  assign n15572 = ~n15570 & ~n15571;
  assign n15573 = ~n15565 & ~n15572;
  assign n15574 = po30  & ~n15573;
  assign n15575 = ~n15029 & ~n15030;
  assign n15576 = po7  & n15575;
  assign n15577 = n15035 & ~n15576;
  assign n15578 = ~n15035 & n15576;
  assign n15579 = ~n15577 & ~n15578;
  assign n15580 = ~po30  & ~n15565;
  assign n15581 = ~n15572 & n15580;
  assign n15582 = ~n15579 & ~n15581;
  assign n15583 = ~n15574 & ~n15582;
  assign n15584 = po31  & ~n15583;
  assign n15585 = ~n15038 & ~n15040;
  assign n15586 = po7  & n15585;
  assign n15587 = n15045 & ~n15586;
  assign n15588 = ~n15045 & n15586;
  assign n15589 = ~n15587 & ~n15588;
  assign n15590 = ~po31  & n15583;
  assign n15591 = ~n15589 & ~n15590;
  assign n15592 = ~n15584 & ~n15591;
  assign n15593 = po32  & ~n15592;
  assign n15594 = ~po32  & ~n15584;
  assign n15595 = ~n15591 & n15594;
  assign n15596 = ~n15048 & po7 ;
  assign n15597 = ~n15054 & n15596;
  assign n15598 = n15053 & ~n15597;
  assign n15599 = n15055 & n15596;
  assign n15600 = ~n15598 & ~n15599;
  assign n15601 = ~n15595 & n15600;
  assign n15602 = ~n15593 & ~n15601;
  assign n15603 = po33  & ~n15602;
  assign n15604 = ~n15057 & ~n15059;
  assign n15605 = po7  & n15604;
  assign n15606 = n15064 & ~n15605;
  assign n15607 = ~n15064 & n15605;
  assign n15608 = ~n15606 & ~n15607;
  assign n15609 = ~po33  & n15602;
  assign n15610 = ~n15608 & ~n15609;
  assign n15611 = ~n15603 & ~n15610;
  assign n15612 = po34  & ~n15611;
  assign n15613 = ~n15067 & ~n15068;
  assign n15614 = po7  & n15613;
  assign n15615 = n15073 & ~n15614;
  assign n15616 = ~n15073 & n15614;
  assign n15617 = ~n15615 & ~n15616;
  assign n15618 = ~po34  & ~n15603;
  assign n15619 = ~n15610 & n15618;
  assign n15620 = ~n15617 & ~n15619;
  assign n15621 = ~n15612 & ~n15620;
  assign n15622 = po35  & ~n15621;
  assign n15623 = ~n15076 & ~n15078;
  assign n15624 = po7  & n15623;
  assign n15625 = n15083 & ~n15624;
  assign n15626 = ~n15083 & n15624;
  assign n15627 = ~n15625 & ~n15626;
  assign n15628 = ~po35  & n15621;
  assign n15629 = ~n15627 & ~n15628;
  assign n15630 = ~n15622 & ~n15629;
  assign n15631 = po36  & ~n15630;
  assign n15632 = ~po36  & ~n15622;
  assign n15633 = ~n15629 & n15632;
  assign n15634 = ~n15086 & po7 ;
  assign n15635 = ~n15092 & n15634;
  assign n15636 = n15091 & ~n15635;
  assign n15637 = n15093 & n15634;
  assign n15638 = ~n15636 & ~n15637;
  assign n15639 = ~n15633 & n15638;
  assign n15640 = ~n15631 & ~n15639;
  assign n15641 = po37  & ~n15640;
  assign n15642 = ~n15095 & ~n15097;
  assign n15643 = po7  & n15642;
  assign n15644 = n15102 & ~n15643;
  assign n15645 = ~n15102 & n15643;
  assign n15646 = ~n15644 & ~n15645;
  assign n15647 = ~po37  & n15640;
  assign n15648 = ~n15646 & ~n15647;
  assign n15649 = ~n15641 & ~n15648;
  assign n15650 = po38  & ~n15649;
  assign n15651 = ~n15105 & ~n15106;
  assign n15652 = po7  & n15651;
  assign n15653 = n15111 & ~n15652;
  assign n15654 = ~n15111 & n15652;
  assign n15655 = ~n15653 & ~n15654;
  assign n15656 = ~po38  & ~n15641;
  assign n15657 = ~n15648 & n15656;
  assign n15658 = ~n15655 & ~n15657;
  assign n15659 = ~n15650 & ~n15658;
  assign n15660 = po39  & ~n15659;
  assign n15661 = ~n15114 & ~n15116;
  assign n15662 = po7  & n15661;
  assign n15663 = n15121 & ~n15662;
  assign n15664 = ~n15121 & n15662;
  assign n15665 = ~n15663 & ~n15664;
  assign n15666 = ~po39  & n15659;
  assign n15667 = ~n15665 & ~n15666;
  assign n15668 = ~n15660 & ~n15667;
  assign n15669 = po40  & ~n15668;
  assign n15670 = ~po40  & ~n15660;
  assign n15671 = ~n15667 & n15670;
  assign n15672 = ~n15124 & po7 ;
  assign n15673 = ~n15130 & n15672;
  assign n15674 = n15129 & ~n15673;
  assign n15675 = n15131 & n15672;
  assign n15676 = ~n15674 & ~n15675;
  assign n15677 = ~n15671 & n15676;
  assign n15678 = ~n15669 & ~n15677;
  assign n15679 = po41  & ~n15678;
  assign n15680 = ~n15133 & ~n15135;
  assign n15681 = po7  & n15680;
  assign n15682 = n15140 & ~n15681;
  assign n15683 = ~n15140 & n15681;
  assign n15684 = ~n15682 & ~n15683;
  assign n15685 = ~po41  & n15678;
  assign n15686 = ~n15684 & ~n15685;
  assign n15687 = ~n15679 & ~n15686;
  assign n15688 = po42  & ~n15687;
  assign n15689 = ~n15143 & ~n15144;
  assign n15690 = po7  & n15689;
  assign n15691 = n15149 & ~n15690;
  assign n15692 = ~n15149 & n15690;
  assign n15693 = ~n15691 & ~n15692;
  assign n15694 = ~po42  & ~n15679;
  assign n15695 = ~n15686 & n15694;
  assign n15696 = ~n15693 & ~n15695;
  assign n15697 = ~n15688 & ~n15696;
  assign n15698 = po43  & ~n15697;
  assign n15699 = ~n15152 & ~n15154;
  assign n15700 = po7  & n15699;
  assign n15701 = n15159 & ~n15700;
  assign n15702 = ~n15159 & n15700;
  assign n15703 = ~n15701 & ~n15702;
  assign n15704 = ~po43  & n15697;
  assign n15705 = ~n15703 & ~n15704;
  assign n15706 = ~n15698 & ~n15705;
  assign n15707 = po44  & ~n15706;
  assign n15708 = ~po44  & ~n15698;
  assign n15709 = ~n15705 & n15708;
  assign n15710 = ~n15162 & po7 ;
  assign n15711 = ~n15168 & n15710;
  assign n15712 = n15167 & ~n15711;
  assign n15713 = n15169 & n15710;
  assign n15714 = ~n15712 & ~n15713;
  assign n15715 = ~n15709 & n15714;
  assign n15716 = ~n15707 & ~n15715;
  assign n15717 = po45  & ~n15716;
  assign n15718 = ~n15171 & ~n15173;
  assign n15719 = po7  & n15718;
  assign n15720 = n15178 & ~n15719;
  assign n15721 = ~n15178 & n15719;
  assign n15722 = ~n15720 & ~n15721;
  assign n15723 = ~po45  & n15716;
  assign n15724 = ~n15722 & ~n15723;
  assign n15725 = ~n15717 & ~n15724;
  assign n15726 = po46  & ~n15725;
  assign n15727 = ~n15181 & ~n15182;
  assign n15728 = po7  & n15727;
  assign n15729 = n15187 & ~n15728;
  assign n15730 = ~n15187 & n15728;
  assign n15731 = ~n15729 & ~n15730;
  assign n15732 = ~po46  & ~n15717;
  assign n15733 = ~n15724 & n15732;
  assign n15734 = ~n15731 & ~n15733;
  assign n15735 = ~n15726 & ~n15734;
  assign n15736 = po47  & ~n15735;
  assign n15737 = ~n15190 & ~n15192;
  assign n15738 = po7  & n15737;
  assign n15739 = n15197 & ~n15738;
  assign n15740 = ~n15197 & n15738;
  assign n15741 = ~n15739 & ~n15740;
  assign n15742 = ~po47  & n15735;
  assign n15743 = ~n15741 & ~n15742;
  assign n15744 = ~n15736 & ~n15743;
  assign n15745 = po48  & ~n15744;
  assign n15746 = ~po48  & ~n15736;
  assign n15747 = ~n15743 & n15746;
  assign n15748 = ~n15200 & po7 ;
  assign n15749 = ~n15206 & n15748;
  assign n15750 = n15205 & ~n15749;
  assign n15751 = n15207 & n15748;
  assign n15752 = ~n15750 & ~n15751;
  assign n15753 = ~n15747 & n15752;
  assign n15754 = ~n15745 & ~n15753;
  assign n15755 = po49  & ~n15754;
  assign n15756 = ~n15209 & ~n15211;
  assign n15757 = po7  & n15756;
  assign n15758 = n15216 & ~n15757;
  assign n15759 = ~n15216 & n15757;
  assign n15760 = ~n15758 & ~n15759;
  assign n15761 = ~po49  & n15754;
  assign n15762 = ~n15760 & ~n15761;
  assign n15763 = ~n15755 & ~n15762;
  assign n15764 = po50  & ~n15763;
  assign n15765 = ~n15219 & ~n15220;
  assign n15766 = po7  & n15765;
  assign n15767 = n15225 & ~n15766;
  assign n15768 = ~n15225 & n15766;
  assign n15769 = ~n15767 & ~n15768;
  assign n15770 = ~po50  & ~n15755;
  assign n15771 = ~n15762 & n15770;
  assign n15772 = ~n15769 & ~n15771;
  assign n15773 = ~n15764 & ~n15772;
  assign n15774 = po51  & ~n15773;
  assign n15775 = ~n15228 & ~n15230;
  assign n15776 = po7  & n15775;
  assign n15777 = n15235 & ~n15776;
  assign n15778 = ~n15235 & n15776;
  assign n15779 = ~n15777 & ~n15778;
  assign n15780 = ~po51  & n15773;
  assign n15781 = ~n15779 & ~n15780;
  assign n15782 = ~n15774 & ~n15781;
  assign n15783 = po52  & ~n15782;
  assign n15784 = ~po52  & ~n15774;
  assign n15785 = ~n15781 & n15784;
  assign n15786 = ~n15238 & po7 ;
  assign n15787 = ~n15244 & n15786;
  assign n15788 = n15243 & ~n15787;
  assign n15789 = n15245 & n15786;
  assign n15790 = ~n15788 & ~n15789;
  assign n15791 = ~n15785 & n15790;
  assign n15792 = ~n15783 & ~n15791;
  assign n15793 = po53  & ~n15792;
  assign n15794 = ~n15247 & ~n15249;
  assign n15795 = po7  & n15794;
  assign n15796 = n15254 & ~n15795;
  assign n15797 = ~n15254 & n15795;
  assign n15798 = ~n15796 & ~n15797;
  assign n15799 = ~po53  & n15792;
  assign n15800 = ~n15798 & ~n15799;
  assign n15801 = ~n15793 & ~n15800;
  assign n15802 = po54  & ~n15801;
  assign n15803 = ~n15257 & ~n15258;
  assign n15804 = po7  & n15803;
  assign n15805 = n15263 & ~n15804;
  assign n15806 = ~n15263 & n15804;
  assign n15807 = ~n15805 & ~n15806;
  assign n15808 = ~po54  & ~n15793;
  assign n15809 = ~n15800 & n15808;
  assign n15810 = ~n15807 & ~n15809;
  assign n15811 = ~n15802 & ~n15810;
  assign n15812 = ~po55  & n15811;
  assign n15813 = ~n15266 & po7 ;
  assign n15814 = ~n15273 & n15813;
  assign n15815 = n15271 & ~n15814;
  assign n15816 = n15274 & n15813;
  assign n15817 = ~n15815 & ~n15816;
  assign n15818 = ~n15812 & n15817;
  assign n15819 = po55  & ~n15811;
  assign n15820 = ~n15818 & ~n15819;
  assign n15821 = po56  & ~n15820;
  assign n15822 = ~po56  & ~n15819;
  assign n15823 = ~n15818 & n15822;
  assign n15824 = ~n15276 & ~n15278;
  assign n15825 = po7  & n15824;
  assign n15826 = n14835 & n15825;
  assign n15827 = ~n14835 & ~n15825;
  assign n15828 = ~n15826 & ~n15827;
  assign n15829 = ~n15823 & ~n15828;
  assign n15830 = ~n15821 & ~n15829;
  assign n15831 = ~po57  & n15830;
  assign n15832 = po57  & ~n15830;
  assign n15833 = ~n15362 & ~n15831;
  assign n15834 = ~n15832 & ~n15833;
  assign n15835 = po58  & ~n15834;
  assign n15836 = ~po58  & ~n15832;
  assign n15837 = ~n15833 & n15836;
  assign n15838 = ~n15285 & po7 ;
  assign n15839 = ~n15291 & n15838;
  assign n15840 = n15290 & ~n15839;
  assign n15841 = n15292 & n15838;
  assign n15842 = ~n15840 & ~n15841;
  assign n15843 = ~n15837 & n15842;
  assign n15844 = ~n15835 & ~n15843;
  assign n15845 = po59  & ~n15844;
  assign n15846 = ~n15294 & ~n15296;
  assign n15847 = po7  & n15846;
  assign n15848 = n15301 & ~n15847;
  assign n15849 = ~n15301 & n15847;
  assign n15850 = ~n15848 & ~n15849;
  assign n15851 = ~po59  & n15844;
  assign n15852 = ~n15850 & ~n15851;
  assign n15853 = ~n15845 & ~n15852;
  assign n15854 = po60  & ~n15853;
  assign n15855 = ~po60  & ~n15845;
  assign n15856 = ~n15852 & n15855;
  assign n15857 = ~n15304 & po7 ;
  assign n15858 = ~n15310 & n15857;
  assign n15859 = n15309 & ~n15858;
  assign n15860 = n15311 & n15857;
  assign n15861 = ~n15859 & ~n15860;
  assign n15862 = ~n15856 & n15861;
  assign n15863 = ~n15854 & ~n15862;
  assign n15864 = po61  & ~n15863;
  assign n15865 = ~n15313 & ~n15315;
  assign n15866 = po7  & n15865;
  assign n15867 = n15320 & ~n15866;
  assign n15868 = ~n15320 & n15866;
  assign n15869 = ~n15867 & ~n15868;
  assign n15870 = ~po61  & n15863;
  assign n15871 = ~n15869 & ~n15870;
  assign n15872 = ~n15864 & ~n15871;
  assign n15873 = po62  & ~n15872;
  assign n15874 = ~n15323 & ~n15324;
  assign n15875 = po7  & n15874;
  assign n15876 = n15329 & ~n15875;
  assign n15877 = ~n15329 & n15875;
  assign n15878 = ~n15876 & ~n15877;
  assign n15879 = ~po62  & ~n15864;
  assign n15880 = ~n15871 & n15879;
  assign n15881 = ~n15878 & ~n15880;
  assign n15882 = ~n15873 & ~n15881;
  assign n15883 = ~n15332 & ~n15334;
  assign n15884 = po7  & n15883;
  assign n15885 = n15339 & ~n15884;
  assign n15886 = ~n15339 & n15884;
  assign n15887 = ~n15885 & ~n15886;
  assign n15888 = n15341 & po7 ;
  assign n15889 = ~n15346 & ~n15888;
  assign n15890 = ~n15354 & ~n15889;
  assign n15891 = po7  & ~n15890;
  assign n15892 = ~n15887 & ~n15891;
  assign n15893 = ~n15882 & n15892;
  assign n15894 = ~po63  & ~n15893;
  assign n15895 = n15882 & n15887;
  assign n15896 = po63  & n15890;
  assign n15897 = ~n15895 & ~n15896;
  assign po6  = n15894 | ~n15897;
  assign n15899 = ~n15832 & po6 ;
  assign n15900 = ~n15831 & n15899;
  assign n15901 = n15362 & ~n15900;
  assign n15902 = n15833 & n15899;
  assign n15903 = ~n15901 & ~n15902;
  assign n15904 = ~n15821 & ~n15823;
  assign n15905 = po6  & n15904;
  assign n15906 = ~n15828 & ~n15905;
  assign n15907 = n15828 & n15905;
  assign n15908 = ~n15906 & ~n15907;
  assign n15909 = pi12  & po6 ;
  assign n15910 = ~pi10  & ~pi11 ;
  assign n15911 = ~pi12  & n15910;
  assign n15912 = ~n15909 & ~n15911;
  assign n15913 = po7  & ~n15912;
  assign n15914 = ~pi12  & po6 ;
  assign n15915 = pi13  & ~n15914;
  assign n15916 = ~pi13  & n15914;
  assign n15917 = ~n15915 & ~n15916;
  assign n15918 = ~po7  & n15912;
  assign n15919 = n15917 & ~n15918;
  assign n15920 = ~n15913 & ~n15919;
  assign n15921 = po8  & ~n15920;
  assign n15922 = ~po8  & ~n15913;
  assign n15923 = ~n15919 & n15922;
  assign n15924 = po7  & ~po6 ;
  assign n15925 = ~n15916 & ~n15924;
  assign n15926 = pi14  & ~n15925;
  assign n15927 = ~pi14  & n15925;
  assign n15928 = ~n15926 & ~n15927;
  assign n15929 = ~n15923 & ~n15928;
  assign n15930 = ~n15921 & ~n15929;
  assign n15931 = po9  & ~n15930;
  assign n15932 = ~po9  & n15930;
  assign n15933 = ~n15367 & ~n15368;
  assign n15934 = po6  & n15933;
  assign n15935 = n15372 & ~n15934;
  assign n15936 = ~n15372 & n15934;
  assign n15937 = ~n15935 & ~n15936;
  assign n15938 = ~n15932 & ~n15937;
  assign n15939 = ~n15931 & ~n15938;
  assign n15940 = po10  & ~n15939;
  assign n15941 = ~po10  & ~n15931;
  assign n15942 = ~n15938 & n15941;
  assign n15943 = ~n15375 & po6 ;
  assign n15944 = ~n15381 & n15943;
  assign n15945 = n15380 & ~n15944;
  assign n15946 = n15382 & n15943;
  assign n15947 = ~n15945 & ~n15946;
  assign n15948 = ~n15942 & n15947;
  assign n15949 = ~n15940 & ~n15948;
  assign n15950 = po11  & ~n15949;
  assign n15951 = ~po11  & n15949;
  assign n15952 = ~n15384 & ~n15386;
  assign n15953 = po6  & n15952;
  assign n15954 = n15391 & ~n15953;
  assign n15955 = ~n15391 & n15953;
  assign n15956 = ~n15954 & ~n15955;
  assign n15957 = ~n15951 & n15956;
  assign n15958 = ~n15950 & ~n15957;
  assign n15959 = po12  & ~n15958;
  assign n15960 = ~po12  & ~n15950;
  assign n15961 = ~n15957 & n15960;
  assign n15962 = ~n15394 & po6 ;
  assign n15963 = ~n15400 & n15962;
  assign n15964 = n15399 & ~n15963;
  assign n15965 = n15401 & n15962;
  assign n15966 = ~n15964 & ~n15965;
  assign n15967 = ~n15961 & n15966;
  assign n15968 = ~n15959 & ~n15967;
  assign n15969 = po13  & ~n15968;
  assign n15970 = ~po13  & n15968;
  assign n15971 = ~n15403 & ~n15405;
  assign n15972 = po6  & n15971;
  assign n15973 = n15410 & n15972;
  assign n15974 = ~n15410 & ~n15972;
  assign n15975 = ~n15973 & ~n15974;
  assign n15976 = ~n15970 & n15975;
  assign n15977 = ~n15969 & ~n15976;
  assign n15978 = po14  & ~n15977;
  assign n15979 = ~po14  & ~n15969;
  assign n15980 = ~n15976 & n15979;
  assign n15981 = ~n15413 & po6 ;
  assign n15982 = ~n15419 & n15981;
  assign n15983 = n15418 & ~n15982;
  assign n15984 = n15420 & n15981;
  assign n15985 = ~n15983 & ~n15984;
  assign n15986 = ~n15980 & n15985;
  assign n15987 = ~n15978 & ~n15986;
  assign n15988 = po15  & ~n15987;
  assign n15989 = ~po15  & n15987;
  assign n15990 = ~n15422 & ~n15424;
  assign n15991 = po6  & n15990;
  assign n15992 = ~n15429 & ~n15991;
  assign n15993 = n15429 & n15991;
  assign n15994 = ~n15992 & ~n15993;
  assign n15995 = ~n15989 & n15994;
  assign n15996 = ~n15988 & ~n15995;
  assign n15997 = po16  & ~n15996;
  assign n15998 = ~po16  & ~n15988;
  assign n15999 = ~n15995 & n15998;
  assign n16000 = ~n15432 & po6 ;
  assign n16001 = ~n15438 & n16000;
  assign n16002 = n15437 & ~n16001;
  assign n16003 = n15439 & n16000;
  assign n16004 = ~n16002 & ~n16003;
  assign n16005 = ~n15999 & n16004;
  assign n16006 = ~n15997 & ~n16005;
  assign n16007 = po17  & ~n16006;
  assign n16008 = ~n15441 & ~n15443;
  assign n16009 = po6  & n16008;
  assign n16010 = n15448 & ~n16009;
  assign n16011 = ~n15448 & n16009;
  assign n16012 = ~n16010 & ~n16011;
  assign n16013 = ~po17  & n16006;
  assign n16014 = ~n16012 & ~n16013;
  assign n16015 = ~n16007 & ~n16014;
  assign n16016 = po18  & ~n16015;
  assign n16017 = ~po18  & ~n16007;
  assign n16018 = ~n16014 & n16017;
  assign n16019 = ~n15451 & po6 ;
  assign n16020 = ~n15457 & n16019;
  assign n16021 = n15456 & ~n16020;
  assign n16022 = n15458 & n16019;
  assign n16023 = ~n16021 & ~n16022;
  assign n16024 = ~n16018 & n16023;
  assign n16025 = ~n16016 & ~n16024;
  assign n16026 = po19  & ~n16025;
  assign n16027 = ~po19  & n16025;
  assign n16028 = ~n15460 & po6 ;
  assign n16029 = ~n15467 & n16028;
  assign n16030 = n15465 & ~n16029;
  assign n16031 = n15468 & n16028;
  assign n16032 = ~n16030 & ~n16031;
  assign n16033 = ~n16027 & n16032;
  assign n16034 = ~n16026 & ~n16033;
  assign n16035 = po20  & ~n16034;
  assign n16036 = ~po20  & ~n16026;
  assign n16037 = ~n16033 & n16036;
  assign n16038 = ~n15470 & po6 ;
  assign n16039 = ~n15476 & n16038;
  assign n16040 = n15475 & ~n16039;
  assign n16041 = n15477 & n16038;
  assign n16042 = ~n16040 & ~n16041;
  assign n16043 = ~n16037 & n16042;
  assign n16044 = ~n16035 & ~n16043;
  assign n16045 = po21  & ~n16044;
  assign n16046 = ~n15479 & ~n15481;
  assign n16047 = po6  & n16046;
  assign n16048 = n15486 & ~n16047;
  assign n16049 = ~n15486 & n16047;
  assign n16050 = ~n16048 & ~n16049;
  assign n16051 = ~po21  & n16044;
  assign n16052 = ~n16050 & ~n16051;
  assign n16053 = ~n16045 & ~n16052;
  assign n16054 = po22  & ~n16053;
  assign n16055 = ~po22  & ~n16045;
  assign n16056 = ~n16052 & n16055;
  assign n16057 = ~n15489 & po6 ;
  assign n16058 = ~n15495 & n16057;
  assign n16059 = n15494 & ~n16058;
  assign n16060 = n15496 & n16057;
  assign n16061 = ~n16059 & ~n16060;
  assign n16062 = ~n16056 & n16061;
  assign n16063 = ~n16054 & ~n16062;
  assign n16064 = po23  & ~n16063;
  assign n16065 = ~po23  & n16063;
  assign n16066 = ~n15498 & po6 ;
  assign n16067 = ~n15505 & n16066;
  assign n16068 = n15503 & ~n16067;
  assign n16069 = n15506 & n16066;
  assign n16070 = ~n16068 & ~n16069;
  assign n16071 = ~n16065 & n16070;
  assign n16072 = ~n16064 & ~n16071;
  assign n16073 = po24  & ~n16072;
  assign n16074 = ~po24  & ~n16064;
  assign n16075 = ~n16071 & n16074;
  assign n16076 = ~n15508 & po6 ;
  assign n16077 = ~n15514 & n16076;
  assign n16078 = n15513 & ~n16077;
  assign n16079 = n15515 & n16076;
  assign n16080 = ~n16078 & ~n16079;
  assign n16081 = ~n16075 & n16080;
  assign n16082 = ~n16073 & ~n16081;
  assign n16083 = po25  & ~n16082;
  assign n16084 = ~n15517 & ~n15519;
  assign n16085 = po6  & n16084;
  assign n16086 = n15524 & ~n16085;
  assign n16087 = ~n15524 & n16085;
  assign n16088 = ~n16086 & ~n16087;
  assign n16089 = ~po25  & n16082;
  assign n16090 = ~n16088 & ~n16089;
  assign n16091 = ~n16083 & ~n16090;
  assign n16092 = po26  & ~n16091;
  assign n16093 = ~po26  & ~n16083;
  assign n16094 = ~n16090 & n16093;
  assign n16095 = ~n15527 & po6 ;
  assign n16096 = ~n15533 & n16095;
  assign n16097 = n15532 & ~n16096;
  assign n16098 = n15534 & n16095;
  assign n16099 = ~n16097 & ~n16098;
  assign n16100 = ~n16094 & n16099;
  assign n16101 = ~n16092 & ~n16100;
  assign n16102 = po27  & ~n16101;
  assign n16103 = ~po27  & n16101;
  assign n16104 = ~n15536 & po6 ;
  assign n16105 = ~n15543 & n16104;
  assign n16106 = n15541 & ~n16105;
  assign n16107 = n15544 & n16104;
  assign n16108 = ~n16106 & ~n16107;
  assign n16109 = ~n16103 & n16108;
  assign n16110 = ~n16102 & ~n16109;
  assign n16111 = po28  & ~n16110;
  assign n16112 = ~po28  & ~n16102;
  assign n16113 = ~n16109 & n16112;
  assign n16114 = ~n15546 & po6 ;
  assign n16115 = ~n15552 & n16114;
  assign n16116 = n15551 & ~n16115;
  assign n16117 = n15553 & n16114;
  assign n16118 = ~n16116 & ~n16117;
  assign n16119 = ~n16113 & n16118;
  assign n16120 = ~n16111 & ~n16119;
  assign n16121 = po29  & ~n16120;
  assign n16122 = ~n15555 & ~n15557;
  assign n16123 = po6  & n16122;
  assign n16124 = n15562 & ~n16123;
  assign n16125 = ~n15562 & n16123;
  assign n16126 = ~n16124 & ~n16125;
  assign n16127 = ~po29  & n16120;
  assign n16128 = ~n16126 & ~n16127;
  assign n16129 = ~n16121 & ~n16128;
  assign n16130 = po30  & ~n16129;
  assign n16131 = ~po30  & ~n16121;
  assign n16132 = ~n16128 & n16131;
  assign n16133 = ~n15565 & po6 ;
  assign n16134 = ~n15571 & n16133;
  assign n16135 = n15570 & ~n16134;
  assign n16136 = n15572 & n16133;
  assign n16137 = ~n16135 & ~n16136;
  assign n16138 = ~n16132 & n16137;
  assign n16139 = ~n16130 & ~n16138;
  assign n16140 = po31  & ~n16139;
  assign n16141 = ~po31  & n16139;
  assign n16142 = ~n15574 & po6 ;
  assign n16143 = ~n15581 & n16142;
  assign n16144 = n15579 & ~n16143;
  assign n16145 = n15582 & n16142;
  assign n16146 = ~n16144 & ~n16145;
  assign n16147 = ~n16141 & n16146;
  assign n16148 = ~n16140 & ~n16147;
  assign n16149 = po32  & ~n16148;
  assign n16150 = ~po32  & ~n16140;
  assign n16151 = ~n16147 & n16150;
  assign n16152 = ~n15584 & po6 ;
  assign n16153 = ~n15590 & n16152;
  assign n16154 = n15589 & ~n16153;
  assign n16155 = n15591 & n16152;
  assign n16156 = ~n16154 & ~n16155;
  assign n16157 = ~n16151 & n16156;
  assign n16158 = ~n16149 & ~n16157;
  assign n16159 = po33  & ~n16158;
  assign n16160 = ~n15593 & ~n15595;
  assign n16161 = po6  & n16160;
  assign n16162 = n15600 & ~n16161;
  assign n16163 = ~n15600 & n16161;
  assign n16164 = ~n16162 & ~n16163;
  assign n16165 = ~po33  & n16158;
  assign n16166 = ~n16164 & ~n16165;
  assign n16167 = ~n16159 & ~n16166;
  assign n16168 = po34  & ~n16167;
  assign n16169 = ~po34  & ~n16159;
  assign n16170 = ~n16166 & n16169;
  assign n16171 = ~n15603 & po6 ;
  assign n16172 = ~n15609 & n16171;
  assign n16173 = n15608 & ~n16172;
  assign n16174 = n15610 & n16171;
  assign n16175 = ~n16173 & ~n16174;
  assign n16176 = ~n16170 & n16175;
  assign n16177 = ~n16168 & ~n16176;
  assign n16178 = po35  & ~n16177;
  assign n16179 = ~po35  & n16177;
  assign n16180 = ~n15612 & po6 ;
  assign n16181 = ~n15619 & n16180;
  assign n16182 = n15617 & ~n16181;
  assign n16183 = n15620 & n16180;
  assign n16184 = ~n16182 & ~n16183;
  assign n16185 = ~n16179 & n16184;
  assign n16186 = ~n16178 & ~n16185;
  assign n16187 = po36  & ~n16186;
  assign n16188 = ~po36  & ~n16178;
  assign n16189 = ~n16185 & n16188;
  assign n16190 = ~n15622 & po6 ;
  assign n16191 = ~n15628 & n16190;
  assign n16192 = n15627 & ~n16191;
  assign n16193 = n15629 & n16190;
  assign n16194 = ~n16192 & ~n16193;
  assign n16195 = ~n16189 & n16194;
  assign n16196 = ~n16187 & ~n16195;
  assign n16197 = po37  & ~n16196;
  assign n16198 = ~n15631 & ~n15633;
  assign n16199 = po6  & n16198;
  assign n16200 = n15638 & ~n16199;
  assign n16201 = ~n15638 & n16199;
  assign n16202 = ~n16200 & ~n16201;
  assign n16203 = ~po37  & n16196;
  assign n16204 = ~n16202 & ~n16203;
  assign n16205 = ~n16197 & ~n16204;
  assign n16206 = po38  & ~n16205;
  assign n16207 = ~po38  & ~n16197;
  assign n16208 = ~n16204 & n16207;
  assign n16209 = ~n15641 & po6 ;
  assign n16210 = ~n15647 & n16209;
  assign n16211 = n15646 & ~n16210;
  assign n16212 = n15648 & n16209;
  assign n16213 = ~n16211 & ~n16212;
  assign n16214 = ~n16208 & n16213;
  assign n16215 = ~n16206 & ~n16214;
  assign n16216 = po39  & ~n16215;
  assign n16217 = ~po39  & n16215;
  assign n16218 = ~n15650 & po6 ;
  assign n16219 = ~n15657 & n16218;
  assign n16220 = n15655 & ~n16219;
  assign n16221 = n15658 & n16218;
  assign n16222 = ~n16220 & ~n16221;
  assign n16223 = ~n16217 & n16222;
  assign n16224 = ~n16216 & ~n16223;
  assign n16225 = po40  & ~n16224;
  assign n16226 = ~po40  & ~n16216;
  assign n16227 = ~n16223 & n16226;
  assign n16228 = ~n15660 & po6 ;
  assign n16229 = ~n15666 & n16228;
  assign n16230 = n15665 & ~n16229;
  assign n16231 = n15667 & n16228;
  assign n16232 = ~n16230 & ~n16231;
  assign n16233 = ~n16227 & n16232;
  assign n16234 = ~n16225 & ~n16233;
  assign n16235 = po41  & ~n16234;
  assign n16236 = ~n15669 & ~n15671;
  assign n16237 = po6  & n16236;
  assign n16238 = n15676 & ~n16237;
  assign n16239 = ~n15676 & n16237;
  assign n16240 = ~n16238 & ~n16239;
  assign n16241 = ~po41  & n16234;
  assign n16242 = ~n16240 & ~n16241;
  assign n16243 = ~n16235 & ~n16242;
  assign n16244 = po42  & ~n16243;
  assign n16245 = ~po42  & ~n16235;
  assign n16246 = ~n16242 & n16245;
  assign n16247 = ~n15679 & po6 ;
  assign n16248 = ~n15685 & n16247;
  assign n16249 = n15684 & ~n16248;
  assign n16250 = n15686 & n16247;
  assign n16251 = ~n16249 & ~n16250;
  assign n16252 = ~n16246 & n16251;
  assign n16253 = ~n16244 & ~n16252;
  assign n16254 = po43  & ~n16253;
  assign n16255 = ~po43  & n16253;
  assign n16256 = ~n15688 & po6 ;
  assign n16257 = ~n15695 & n16256;
  assign n16258 = n15693 & ~n16257;
  assign n16259 = n15696 & n16256;
  assign n16260 = ~n16258 & ~n16259;
  assign n16261 = ~n16255 & n16260;
  assign n16262 = ~n16254 & ~n16261;
  assign n16263 = po44  & ~n16262;
  assign n16264 = ~po44  & ~n16254;
  assign n16265 = ~n16261 & n16264;
  assign n16266 = ~n15698 & po6 ;
  assign n16267 = ~n15704 & n16266;
  assign n16268 = n15703 & ~n16267;
  assign n16269 = n15705 & n16266;
  assign n16270 = ~n16268 & ~n16269;
  assign n16271 = ~n16265 & n16270;
  assign n16272 = ~n16263 & ~n16271;
  assign n16273 = po45  & ~n16272;
  assign n16274 = ~n15707 & ~n15709;
  assign n16275 = po6  & n16274;
  assign n16276 = n15714 & ~n16275;
  assign n16277 = ~n15714 & n16275;
  assign n16278 = ~n16276 & ~n16277;
  assign n16279 = ~po45  & n16272;
  assign n16280 = ~n16278 & ~n16279;
  assign n16281 = ~n16273 & ~n16280;
  assign n16282 = po46  & ~n16281;
  assign n16283 = ~po46  & ~n16273;
  assign n16284 = ~n16280 & n16283;
  assign n16285 = ~n15717 & po6 ;
  assign n16286 = ~n15723 & n16285;
  assign n16287 = n15722 & ~n16286;
  assign n16288 = n15724 & n16285;
  assign n16289 = ~n16287 & ~n16288;
  assign n16290 = ~n16284 & n16289;
  assign n16291 = ~n16282 & ~n16290;
  assign n16292 = po47  & ~n16291;
  assign n16293 = ~po47  & n16291;
  assign n16294 = ~n15726 & po6 ;
  assign n16295 = ~n15733 & n16294;
  assign n16296 = n15731 & ~n16295;
  assign n16297 = n15734 & n16294;
  assign n16298 = ~n16296 & ~n16297;
  assign n16299 = ~n16293 & n16298;
  assign n16300 = ~n16292 & ~n16299;
  assign n16301 = po48  & ~n16300;
  assign n16302 = ~po48  & ~n16292;
  assign n16303 = ~n16299 & n16302;
  assign n16304 = ~n15736 & po6 ;
  assign n16305 = ~n15742 & n16304;
  assign n16306 = n15741 & ~n16305;
  assign n16307 = n15743 & n16304;
  assign n16308 = ~n16306 & ~n16307;
  assign n16309 = ~n16303 & n16308;
  assign n16310 = ~n16301 & ~n16309;
  assign n16311 = po49  & ~n16310;
  assign n16312 = ~n15745 & ~n15747;
  assign n16313 = po6  & n16312;
  assign n16314 = n15752 & ~n16313;
  assign n16315 = ~n15752 & n16313;
  assign n16316 = ~n16314 & ~n16315;
  assign n16317 = ~po49  & n16310;
  assign n16318 = ~n16316 & ~n16317;
  assign n16319 = ~n16311 & ~n16318;
  assign n16320 = po50  & ~n16319;
  assign n16321 = ~po50  & ~n16311;
  assign n16322 = ~n16318 & n16321;
  assign n16323 = ~n15755 & po6 ;
  assign n16324 = ~n15761 & n16323;
  assign n16325 = n15760 & ~n16324;
  assign n16326 = n15762 & n16323;
  assign n16327 = ~n16325 & ~n16326;
  assign n16328 = ~n16322 & n16327;
  assign n16329 = ~n16320 & ~n16328;
  assign n16330 = po51  & ~n16329;
  assign n16331 = ~po51  & n16329;
  assign n16332 = ~n15764 & po6 ;
  assign n16333 = ~n15771 & n16332;
  assign n16334 = n15769 & ~n16333;
  assign n16335 = n15772 & n16332;
  assign n16336 = ~n16334 & ~n16335;
  assign n16337 = ~n16331 & n16336;
  assign n16338 = ~n16330 & ~n16337;
  assign n16339 = po52  & ~n16338;
  assign n16340 = ~po52  & ~n16330;
  assign n16341 = ~n16337 & n16340;
  assign n16342 = ~n15774 & po6 ;
  assign n16343 = ~n15780 & n16342;
  assign n16344 = n15779 & ~n16343;
  assign n16345 = n15781 & n16342;
  assign n16346 = ~n16344 & ~n16345;
  assign n16347 = ~n16341 & n16346;
  assign n16348 = ~n16339 & ~n16347;
  assign n16349 = po53  & ~n16348;
  assign n16350 = ~n15783 & ~n15785;
  assign n16351 = po6  & n16350;
  assign n16352 = n15790 & ~n16351;
  assign n16353 = ~n15790 & n16351;
  assign n16354 = ~n16352 & ~n16353;
  assign n16355 = ~po53  & n16348;
  assign n16356 = ~n16354 & ~n16355;
  assign n16357 = ~n16349 & ~n16356;
  assign n16358 = po54  & ~n16357;
  assign n16359 = ~po54  & ~n16349;
  assign n16360 = ~n16356 & n16359;
  assign n16361 = ~n15793 & po6 ;
  assign n16362 = ~n15799 & n16361;
  assign n16363 = n15798 & ~n16362;
  assign n16364 = n15800 & n16361;
  assign n16365 = ~n16363 & ~n16364;
  assign n16366 = ~n16360 & n16365;
  assign n16367 = ~n16358 & ~n16366;
  assign n16368 = po55  & ~n16367;
  assign n16369 = ~po55  & n16367;
  assign n16370 = ~n15802 & po6 ;
  assign n16371 = ~n15809 & n16370;
  assign n16372 = n15807 & ~n16371;
  assign n16373 = n15810 & n16370;
  assign n16374 = ~n16372 & ~n16373;
  assign n16375 = ~n16369 & n16374;
  assign n16376 = ~n16368 & ~n16375;
  assign n16377 = po56  & ~n16376;
  assign n16378 = ~n15812 & ~n15819;
  assign n16379 = po6  & n16378;
  assign n16380 = n15817 & ~n16379;
  assign n16381 = ~n15817 & n16379;
  assign n16382 = ~n16380 & ~n16381;
  assign n16383 = ~po56  & ~n16368;
  assign n16384 = ~n16375 & n16383;
  assign n16385 = ~n16382 & ~n16384;
  assign n16386 = ~n16377 & ~n16385;
  assign n16387 = ~po57  & n16386;
  assign n16388 = ~n15908 & ~n16387;
  assign n16389 = po57  & ~n16386;
  assign n16390 = ~po58  & ~n16389;
  assign n16391 = ~n16388 & n16390;
  assign n16392 = ~n16388 & ~n16389;
  assign n16393 = po58  & ~n16392;
  assign n16394 = n15903 & ~n16391;
  assign n16395 = ~n16393 & ~n16394;
  assign n16396 = po59  & ~n16395;
  assign n16397 = ~n15835 & ~n15837;
  assign n16398 = po6  & n16397;
  assign n16399 = n15842 & ~n16398;
  assign n16400 = ~n15842 & n16398;
  assign n16401 = ~n16399 & ~n16400;
  assign n16402 = ~po59  & n16395;
  assign n16403 = ~n16401 & ~n16402;
  assign n16404 = ~n16396 & ~n16403;
  assign n16405 = po60  & ~n16404;
  assign n16406 = ~po60  & ~n16396;
  assign n16407 = ~n16403 & n16406;
  assign n16408 = ~n15845 & po6 ;
  assign n16409 = ~n15851 & n16408;
  assign n16410 = n15850 & ~n16409;
  assign n16411 = n15852 & n16408;
  assign n16412 = ~n16410 & ~n16411;
  assign n16413 = ~n16407 & n16412;
  assign n16414 = ~n16405 & ~n16413;
  assign n16415 = po61  & ~n16414;
  assign n16416 = ~n15854 & ~n15856;
  assign n16417 = po6  & n16416;
  assign n16418 = n15861 & ~n16417;
  assign n16419 = ~n15861 & n16417;
  assign n16420 = ~n16418 & ~n16419;
  assign n16421 = ~po61  & n16414;
  assign n16422 = ~n16420 & ~n16421;
  assign n16423 = ~n16415 & ~n16422;
  assign n16424 = po62  & ~n16423;
  assign n16425 = ~po62  & ~n16415;
  assign n16426 = ~n16422 & n16425;
  assign n16427 = ~n15864 & po6 ;
  assign n16428 = ~n15870 & n16427;
  assign n16429 = n15869 & ~n16428;
  assign n16430 = n15871 & n16427;
  assign n16431 = ~n16429 & ~n16430;
  assign n16432 = ~n16426 & n16431;
  assign n16433 = ~n16424 & ~n16432;
  assign n16434 = n15882 & po6 ;
  assign n16435 = ~n15887 & ~n16434;
  assign n16436 = ~n15895 & ~n16435;
  assign n16437 = po6  & ~n16436;
  assign n16438 = ~n15873 & po6 ;
  assign n16439 = ~n15880 & n16438;
  assign n16440 = n15878 & ~n16439;
  assign n16441 = n15881 & n16438;
  assign n16442 = ~n16440 & ~n16441;
  assign n16443 = ~n16437 & n16442;
  assign n16444 = ~n16433 & n16443;
  assign n16445 = ~po63  & ~n16444;
  assign n16446 = n16433 & ~n16442;
  assign n16447 = po63  & n16436;
  assign n16448 = ~n16446 & ~n16447;
  assign po5  = n16445 | ~n16448;
  assign n16450 = ~n16391 & ~n16393;
  assign n16451 = po5  & n16450;
  assign n16452 = n15903 & ~n16451;
  assign n16453 = ~n15903 & n16451;
  assign n16454 = ~n16452 & ~n16453;
  assign n16455 = pi10  & po5 ;
  assign n16456 = ~pi8  & ~pi9 ;
  assign n16457 = ~pi10  & n16456;
  assign n16458 = ~n16455 & ~n16457;
  assign n16459 = po6  & ~n16458;
  assign n16460 = ~po6  & n16458;
  assign n16461 = ~pi10  & po5 ;
  assign n16462 = pi11  & ~n16461;
  assign n16463 = ~pi11  & n16461;
  assign n16464 = ~n16462 & ~n16463;
  assign n16465 = ~n16460 & n16464;
  assign n16466 = ~n16459 & ~n16465;
  assign n16467 = po7  & ~n16466;
  assign n16468 = po6  & ~po5 ;
  assign n16469 = ~n16463 & ~n16468;
  assign n16470 = pi12  & ~n16469;
  assign n16471 = ~pi12  & n16469;
  assign n16472 = ~n16470 & ~n16471;
  assign n16473 = ~po7  & n16466;
  assign n16474 = ~n16472 & ~n16473;
  assign n16475 = ~n16467 & ~n16474;
  assign n16476 = po8  & ~n16475;
  assign n16477 = ~po8  & ~n16467;
  assign n16478 = ~n16474 & n16477;
  assign n16479 = ~n15913 & ~n15918;
  assign n16480 = po5  & n16479;
  assign n16481 = n15917 & ~n16480;
  assign n16482 = ~n15917 & n16480;
  assign n16483 = ~n16481 & ~n16482;
  assign n16484 = ~n16478 & ~n16483;
  assign n16485 = ~n16476 & ~n16484;
  assign n16486 = po9  & ~n16485;
  assign n16487 = ~n15921 & ~n15923;
  assign n16488 = po5  & n16487;
  assign n16489 = ~n15928 & ~n16488;
  assign n16490 = n15928 & n16488;
  assign n16491 = ~n16489 & ~n16490;
  assign n16492 = ~po9  & n16485;
  assign n16493 = ~n16491 & ~n16492;
  assign n16494 = ~n16486 & ~n16493;
  assign n16495 = po10  & ~n16494;
  assign n16496 = ~po10  & ~n16486;
  assign n16497 = ~n16493 & n16496;
  assign n16498 = ~n15931 & ~n15932;
  assign n16499 = po5  & n16498;
  assign n16500 = n15937 & ~n16499;
  assign n16501 = ~n15937 & n16499;
  assign n16502 = ~n16500 & ~n16501;
  assign n16503 = ~n16497 & n16502;
  assign n16504 = ~n16495 & ~n16503;
  assign n16505 = po11  & ~n16504;
  assign n16506 = ~n15940 & ~n15942;
  assign n16507 = po5  & n16506;
  assign n16508 = n15947 & ~n16507;
  assign n16509 = ~n15947 & n16507;
  assign n16510 = ~n16508 & ~n16509;
  assign n16511 = ~po11  & n16504;
  assign n16512 = ~n16510 & ~n16511;
  assign n16513 = ~n16505 & ~n16512;
  assign n16514 = po12  & ~n16513;
  assign n16515 = ~po12  & ~n16505;
  assign n16516 = ~n16512 & n16515;
  assign n16517 = ~n15950 & ~n15951;
  assign n16518 = po5  & n16517;
  assign n16519 = n15956 & n16518;
  assign n16520 = ~n15956 & ~n16518;
  assign n16521 = ~n16519 & ~n16520;
  assign n16522 = ~n16516 & n16521;
  assign n16523 = ~n16514 & ~n16522;
  assign n16524 = po13  & ~n16523;
  assign n16525 = ~n15959 & ~n15961;
  assign n16526 = po5  & n16525;
  assign n16527 = n15966 & ~n16526;
  assign n16528 = ~n15966 & n16526;
  assign n16529 = ~n16527 & ~n16528;
  assign n16530 = ~po13  & n16523;
  assign n16531 = ~n16529 & ~n16530;
  assign n16532 = ~n16524 & ~n16531;
  assign n16533 = po14  & ~n16532;
  assign n16534 = ~po14  & ~n16524;
  assign n16535 = ~n16531 & n16534;
  assign n16536 = ~n15969 & ~n15970;
  assign n16537 = po5  & n16536;
  assign n16538 = ~n15975 & ~n16537;
  assign n16539 = n15975 & n16537;
  assign n16540 = ~n16538 & ~n16539;
  assign n16541 = ~n16535 & n16540;
  assign n16542 = ~n16533 & ~n16541;
  assign n16543 = po15  & ~n16542;
  assign n16544 = ~n15978 & ~n15980;
  assign n16545 = po5  & n16544;
  assign n16546 = n15985 & ~n16545;
  assign n16547 = ~n15985 & n16545;
  assign n16548 = ~n16546 & ~n16547;
  assign n16549 = ~po15  & n16542;
  assign n16550 = ~n16548 & ~n16549;
  assign n16551 = ~n16543 & ~n16550;
  assign n16552 = po16  & ~n16551;
  assign n16553 = ~n15988 & ~n15989;
  assign n16554 = po5  & n16553;
  assign n16555 = n15994 & ~n16554;
  assign n16556 = ~n15994 & n16554;
  assign n16557 = ~n16555 & ~n16556;
  assign n16558 = ~po16  & ~n16543;
  assign n16559 = ~n16550 & n16558;
  assign n16560 = ~n16557 & ~n16559;
  assign n16561 = ~n16552 & ~n16560;
  assign n16562 = po17  & ~n16561;
  assign n16563 = ~n15997 & ~n15999;
  assign n16564 = po5  & n16563;
  assign n16565 = n16004 & ~n16564;
  assign n16566 = ~n16004 & n16564;
  assign n16567 = ~n16565 & ~n16566;
  assign n16568 = ~po17  & n16561;
  assign n16569 = ~n16567 & ~n16568;
  assign n16570 = ~n16562 & ~n16569;
  assign n16571 = po18  & ~n16570;
  assign n16572 = ~po18  & ~n16562;
  assign n16573 = ~n16569 & n16572;
  assign n16574 = ~n16007 & po5 ;
  assign n16575 = ~n16013 & n16574;
  assign n16576 = n16012 & ~n16575;
  assign n16577 = n16014 & n16574;
  assign n16578 = ~n16576 & ~n16577;
  assign n16579 = ~n16573 & n16578;
  assign n16580 = ~n16571 & ~n16579;
  assign n16581 = po19  & ~n16580;
  assign n16582 = ~n16016 & ~n16018;
  assign n16583 = po5  & n16582;
  assign n16584 = n16023 & ~n16583;
  assign n16585 = ~n16023 & n16583;
  assign n16586 = ~n16584 & ~n16585;
  assign n16587 = ~po19  & n16580;
  assign n16588 = ~n16586 & ~n16587;
  assign n16589 = ~n16581 & ~n16588;
  assign n16590 = po20  & ~n16589;
  assign n16591 = ~n16026 & ~n16027;
  assign n16592 = po5  & n16591;
  assign n16593 = n16032 & ~n16592;
  assign n16594 = ~n16032 & n16592;
  assign n16595 = ~n16593 & ~n16594;
  assign n16596 = ~po20  & ~n16581;
  assign n16597 = ~n16588 & n16596;
  assign n16598 = ~n16595 & ~n16597;
  assign n16599 = ~n16590 & ~n16598;
  assign n16600 = po21  & ~n16599;
  assign n16601 = ~n16035 & ~n16037;
  assign n16602 = po5  & n16601;
  assign n16603 = n16042 & ~n16602;
  assign n16604 = ~n16042 & n16602;
  assign n16605 = ~n16603 & ~n16604;
  assign n16606 = ~po21  & n16599;
  assign n16607 = ~n16605 & ~n16606;
  assign n16608 = ~n16600 & ~n16607;
  assign n16609 = po22  & ~n16608;
  assign n16610 = ~po22  & ~n16600;
  assign n16611 = ~n16607 & n16610;
  assign n16612 = ~n16045 & po5 ;
  assign n16613 = ~n16051 & n16612;
  assign n16614 = n16050 & ~n16613;
  assign n16615 = n16052 & n16612;
  assign n16616 = ~n16614 & ~n16615;
  assign n16617 = ~n16611 & n16616;
  assign n16618 = ~n16609 & ~n16617;
  assign n16619 = po23  & ~n16618;
  assign n16620 = ~n16054 & ~n16056;
  assign n16621 = po5  & n16620;
  assign n16622 = n16061 & ~n16621;
  assign n16623 = ~n16061 & n16621;
  assign n16624 = ~n16622 & ~n16623;
  assign n16625 = ~po23  & n16618;
  assign n16626 = ~n16624 & ~n16625;
  assign n16627 = ~n16619 & ~n16626;
  assign n16628 = po24  & ~n16627;
  assign n16629 = ~n16064 & ~n16065;
  assign n16630 = po5  & n16629;
  assign n16631 = n16070 & ~n16630;
  assign n16632 = ~n16070 & n16630;
  assign n16633 = ~n16631 & ~n16632;
  assign n16634 = ~po24  & ~n16619;
  assign n16635 = ~n16626 & n16634;
  assign n16636 = ~n16633 & ~n16635;
  assign n16637 = ~n16628 & ~n16636;
  assign n16638 = po25  & ~n16637;
  assign n16639 = ~n16073 & ~n16075;
  assign n16640 = po5  & n16639;
  assign n16641 = n16080 & ~n16640;
  assign n16642 = ~n16080 & n16640;
  assign n16643 = ~n16641 & ~n16642;
  assign n16644 = ~po25  & n16637;
  assign n16645 = ~n16643 & ~n16644;
  assign n16646 = ~n16638 & ~n16645;
  assign n16647 = po26  & ~n16646;
  assign n16648 = ~po26  & ~n16638;
  assign n16649 = ~n16645 & n16648;
  assign n16650 = ~n16083 & po5 ;
  assign n16651 = ~n16089 & n16650;
  assign n16652 = n16088 & ~n16651;
  assign n16653 = n16090 & n16650;
  assign n16654 = ~n16652 & ~n16653;
  assign n16655 = ~n16649 & n16654;
  assign n16656 = ~n16647 & ~n16655;
  assign n16657 = po27  & ~n16656;
  assign n16658 = ~n16092 & ~n16094;
  assign n16659 = po5  & n16658;
  assign n16660 = n16099 & ~n16659;
  assign n16661 = ~n16099 & n16659;
  assign n16662 = ~n16660 & ~n16661;
  assign n16663 = ~po27  & n16656;
  assign n16664 = ~n16662 & ~n16663;
  assign n16665 = ~n16657 & ~n16664;
  assign n16666 = po28  & ~n16665;
  assign n16667 = ~n16102 & ~n16103;
  assign n16668 = po5  & n16667;
  assign n16669 = n16108 & ~n16668;
  assign n16670 = ~n16108 & n16668;
  assign n16671 = ~n16669 & ~n16670;
  assign n16672 = ~po28  & ~n16657;
  assign n16673 = ~n16664 & n16672;
  assign n16674 = ~n16671 & ~n16673;
  assign n16675 = ~n16666 & ~n16674;
  assign n16676 = po29  & ~n16675;
  assign n16677 = ~n16111 & ~n16113;
  assign n16678 = po5  & n16677;
  assign n16679 = n16118 & ~n16678;
  assign n16680 = ~n16118 & n16678;
  assign n16681 = ~n16679 & ~n16680;
  assign n16682 = ~po29  & n16675;
  assign n16683 = ~n16681 & ~n16682;
  assign n16684 = ~n16676 & ~n16683;
  assign n16685 = po30  & ~n16684;
  assign n16686 = ~po30  & ~n16676;
  assign n16687 = ~n16683 & n16686;
  assign n16688 = ~n16121 & po5 ;
  assign n16689 = ~n16127 & n16688;
  assign n16690 = n16126 & ~n16689;
  assign n16691 = n16128 & n16688;
  assign n16692 = ~n16690 & ~n16691;
  assign n16693 = ~n16687 & n16692;
  assign n16694 = ~n16685 & ~n16693;
  assign n16695 = po31  & ~n16694;
  assign n16696 = ~n16130 & ~n16132;
  assign n16697 = po5  & n16696;
  assign n16698 = n16137 & ~n16697;
  assign n16699 = ~n16137 & n16697;
  assign n16700 = ~n16698 & ~n16699;
  assign n16701 = ~po31  & n16694;
  assign n16702 = ~n16700 & ~n16701;
  assign n16703 = ~n16695 & ~n16702;
  assign n16704 = po32  & ~n16703;
  assign n16705 = ~n16140 & ~n16141;
  assign n16706 = po5  & n16705;
  assign n16707 = n16146 & ~n16706;
  assign n16708 = ~n16146 & n16706;
  assign n16709 = ~n16707 & ~n16708;
  assign n16710 = ~po32  & ~n16695;
  assign n16711 = ~n16702 & n16710;
  assign n16712 = ~n16709 & ~n16711;
  assign n16713 = ~n16704 & ~n16712;
  assign n16714 = po33  & ~n16713;
  assign n16715 = ~n16149 & ~n16151;
  assign n16716 = po5  & n16715;
  assign n16717 = n16156 & ~n16716;
  assign n16718 = ~n16156 & n16716;
  assign n16719 = ~n16717 & ~n16718;
  assign n16720 = ~po33  & n16713;
  assign n16721 = ~n16719 & ~n16720;
  assign n16722 = ~n16714 & ~n16721;
  assign n16723 = po34  & ~n16722;
  assign n16724 = ~po34  & ~n16714;
  assign n16725 = ~n16721 & n16724;
  assign n16726 = ~n16159 & po5 ;
  assign n16727 = ~n16165 & n16726;
  assign n16728 = n16164 & ~n16727;
  assign n16729 = n16166 & n16726;
  assign n16730 = ~n16728 & ~n16729;
  assign n16731 = ~n16725 & n16730;
  assign n16732 = ~n16723 & ~n16731;
  assign n16733 = po35  & ~n16732;
  assign n16734 = ~n16168 & ~n16170;
  assign n16735 = po5  & n16734;
  assign n16736 = n16175 & ~n16735;
  assign n16737 = ~n16175 & n16735;
  assign n16738 = ~n16736 & ~n16737;
  assign n16739 = ~po35  & n16732;
  assign n16740 = ~n16738 & ~n16739;
  assign n16741 = ~n16733 & ~n16740;
  assign n16742 = po36  & ~n16741;
  assign n16743 = ~n16178 & ~n16179;
  assign n16744 = po5  & n16743;
  assign n16745 = n16184 & ~n16744;
  assign n16746 = ~n16184 & n16744;
  assign n16747 = ~n16745 & ~n16746;
  assign n16748 = ~po36  & ~n16733;
  assign n16749 = ~n16740 & n16748;
  assign n16750 = ~n16747 & ~n16749;
  assign n16751 = ~n16742 & ~n16750;
  assign n16752 = po37  & ~n16751;
  assign n16753 = ~n16187 & ~n16189;
  assign n16754 = po5  & n16753;
  assign n16755 = n16194 & ~n16754;
  assign n16756 = ~n16194 & n16754;
  assign n16757 = ~n16755 & ~n16756;
  assign n16758 = ~po37  & n16751;
  assign n16759 = ~n16757 & ~n16758;
  assign n16760 = ~n16752 & ~n16759;
  assign n16761 = po38  & ~n16760;
  assign n16762 = ~po38  & ~n16752;
  assign n16763 = ~n16759 & n16762;
  assign n16764 = ~n16197 & po5 ;
  assign n16765 = ~n16203 & n16764;
  assign n16766 = n16202 & ~n16765;
  assign n16767 = n16204 & n16764;
  assign n16768 = ~n16766 & ~n16767;
  assign n16769 = ~n16763 & n16768;
  assign n16770 = ~n16761 & ~n16769;
  assign n16771 = po39  & ~n16770;
  assign n16772 = ~n16206 & ~n16208;
  assign n16773 = po5  & n16772;
  assign n16774 = n16213 & ~n16773;
  assign n16775 = ~n16213 & n16773;
  assign n16776 = ~n16774 & ~n16775;
  assign n16777 = ~po39  & n16770;
  assign n16778 = ~n16776 & ~n16777;
  assign n16779 = ~n16771 & ~n16778;
  assign n16780 = po40  & ~n16779;
  assign n16781 = ~n16216 & ~n16217;
  assign n16782 = po5  & n16781;
  assign n16783 = n16222 & ~n16782;
  assign n16784 = ~n16222 & n16782;
  assign n16785 = ~n16783 & ~n16784;
  assign n16786 = ~po40  & ~n16771;
  assign n16787 = ~n16778 & n16786;
  assign n16788 = ~n16785 & ~n16787;
  assign n16789 = ~n16780 & ~n16788;
  assign n16790 = po41  & ~n16789;
  assign n16791 = ~n16225 & ~n16227;
  assign n16792 = po5  & n16791;
  assign n16793 = n16232 & ~n16792;
  assign n16794 = ~n16232 & n16792;
  assign n16795 = ~n16793 & ~n16794;
  assign n16796 = ~po41  & n16789;
  assign n16797 = ~n16795 & ~n16796;
  assign n16798 = ~n16790 & ~n16797;
  assign n16799 = po42  & ~n16798;
  assign n16800 = ~po42  & ~n16790;
  assign n16801 = ~n16797 & n16800;
  assign n16802 = ~n16235 & po5 ;
  assign n16803 = ~n16241 & n16802;
  assign n16804 = n16240 & ~n16803;
  assign n16805 = n16242 & n16802;
  assign n16806 = ~n16804 & ~n16805;
  assign n16807 = ~n16801 & n16806;
  assign n16808 = ~n16799 & ~n16807;
  assign n16809 = po43  & ~n16808;
  assign n16810 = ~n16244 & ~n16246;
  assign n16811 = po5  & n16810;
  assign n16812 = n16251 & ~n16811;
  assign n16813 = ~n16251 & n16811;
  assign n16814 = ~n16812 & ~n16813;
  assign n16815 = ~po43  & n16808;
  assign n16816 = ~n16814 & ~n16815;
  assign n16817 = ~n16809 & ~n16816;
  assign n16818 = po44  & ~n16817;
  assign n16819 = ~n16254 & ~n16255;
  assign n16820 = po5  & n16819;
  assign n16821 = n16260 & ~n16820;
  assign n16822 = ~n16260 & n16820;
  assign n16823 = ~n16821 & ~n16822;
  assign n16824 = ~po44  & ~n16809;
  assign n16825 = ~n16816 & n16824;
  assign n16826 = ~n16823 & ~n16825;
  assign n16827 = ~n16818 & ~n16826;
  assign n16828 = po45  & ~n16827;
  assign n16829 = ~n16263 & ~n16265;
  assign n16830 = po5  & n16829;
  assign n16831 = n16270 & ~n16830;
  assign n16832 = ~n16270 & n16830;
  assign n16833 = ~n16831 & ~n16832;
  assign n16834 = ~po45  & n16827;
  assign n16835 = ~n16833 & ~n16834;
  assign n16836 = ~n16828 & ~n16835;
  assign n16837 = po46  & ~n16836;
  assign n16838 = ~po46  & ~n16828;
  assign n16839 = ~n16835 & n16838;
  assign n16840 = ~n16273 & po5 ;
  assign n16841 = ~n16279 & n16840;
  assign n16842 = n16278 & ~n16841;
  assign n16843 = n16280 & n16840;
  assign n16844 = ~n16842 & ~n16843;
  assign n16845 = ~n16839 & n16844;
  assign n16846 = ~n16837 & ~n16845;
  assign n16847 = po47  & ~n16846;
  assign n16848 = ~n16282 & ~n16284;
  assign n16849 = po5  & n16848;
  assign n16850 = n16289 & ~n16849;
  assign n16851 = ~n16289 & n16849;
  assign n16852 = ~n16850 & ~n16851;
  assign n16853 = ~po47  & n16846;
  assign n16854 = ~n16852 & ~n16853;
  assign n16855 = ~n16847 & ~n16854;
  assign n16856 = po48  & ~n16855;
  assign n16857 = ~n16292 & ~n16293;
  assign n16858 = po5  & n16857;
  assign n16859 = n16298 & ~n16858;
  assign n16860 = ~n16298 & n16858;
  assign n16861 = ~n16859 & ~n16860;
  assign n16862 = ~po48  & ~n16847;
  assign n16863 = ~n16854 & n16862;
  assign n16864 = ~n16861 & ~n16863;
  assign n16865 = ~n16856 & ~n16864;
  assign n16866 = po49  & ~n16865;
  assign n16867 = ~n16301 & ~n16303;
  assign n16868 = po5  & n16867;
  assign n16869 = n16308 & ~n16868;
  assign n16870 = ~n16308 & n16868;
  assign n16871 = ~n16869 & ~n16870;
  assign n16872 = ~po49  & n16865;
  assign n16873 = ~n16871 & ~n16872;
  assign n16874 = ~n16866 & ~n16873;
  assign n16875 = po50  & ~n16874;
  assign n16876 = ~po50  & ~n16866;
  assign n16877 = ~n16873 & n16876;
  assign n16878 = ~n16311 & po5 ;
  assign n16879 = ~n16317 & n16878;
  assign n16880 = n16316 & ~n16879;
  assign n16881 = n16318 & n16878;
  assign n16882 = ~n16880 & ~n16881;
  assign n16883 = ~n16877 & n16882;
  assign n16884 = ~n16875 & ~n16883;
  assign n16885 = po51  & ~n16884;
  assign n16886 = ~n16320 & ~n16322;
  assign n16887 = po5  & n16886;
  assign n16888 = n16327 & ~n16887;
  assign n16889 = ~n16327 & n16887;
  assign n16890 = ~n16888 & ~n16889;
  assign n16891 = ~po51  & n16884;
  assign n16892 = ~n16890 & ~n16891;
  assign n16893 = ~n16885 & ~n16892;
  assign n16894 = po52  & ~n16893;
  assign n16895 = ~n16330 & ~n16331;
  assign n16896 = po5  & n16895;
  assign n16897 = n16336 & ~n16896;
  assign n16898 = ~n16336 & n16896;
  assign n16899 = ~n16897 & ~n16898;
  assign n16900 = ~po52  & ~n16885;
  assign n16901 = ~n16892 & n16900;
  assign n16902 = ~n16899 & ~n16901;
  assign n16903 = ~n16894 & ~n16902;
  assign n16904 = po53  & ~n16903;
  assign n16905 = ~n16339 & ~n16341;
  assign n16906 = po5  & n16905;
  assign n16907 = n16346 & ~n16906;
  assign n16908 = ~n16346 & n16906;
  assign n16909 = ~n16907 & ~n16908;
  assign n16910 = ~po53  & n16903;
  assign n16911 = ~n16909 & ~n16910;
  assign n16912 = ~n16904 & ~n16911;
  assign n16913 = po54  & ~n16912;
  assign n16914 = ~po54  & ~n16904;
  assign n16915 = ~n16911 & n16914;
  assign n16916 = ~n16349 & po5 ;
  assign n16917 = ~n16355 & n16916;
  assign n16918 = n16354 & ~n16917;
  assign n16919 = n16356 & n16916;
  assign n16920 = ~n16918 & ~n16919;
  assign n16921 = ~n16915 & n16920;
  assign n16922 = ~n16913 & ~n16921;
  assign n16923 = po55  & ~n16922;
  assign n16924 = ~n16358 & ~n16360;
  assign n16925 = po5  & n16924;
  assign n16926 = n16365 & ~n16925;
  assign n16927 = ~n16365 & n16925;
  assign n16928 = ~n16926 & ~n16927;
  assign n16929 = ~po55  & n16922;
  assign n16930 = ~n16928 & ~n16929;
  assign n16931 = ~n16923 & ~n16930;
  assign n16932 = po56  & ~n16931;
  assign n16933 = ~n16368 & ~n16369;
  assign n16934 = po5  & n16933;
  assign n16935 = n16374 & ~n16934;
  assign n16936 = ~n16374 & n16934;
  assign n16937 = ~n16935 & ~n16936;
  assign n16938 = ~po56  & ~n16923;
  assign n16939 = ~n16930 & n16938;
  assign n16940 = ~n16937 & ~n16939;
  assign n16941 = ~n16932 & ~n16940;
  assign n16942 = ~po57  & n16941;
  assign n16943 = ~n16377 & po5 ;
  assign n16944 = ~n16384 & n16943;
  assign n16945 = n16382 & ~n16944;
  assign n16946 = n16385 & n16943;
  assign n16947 = ~n16945 & ~n16946;
  assign n16948 = ~n16942 & n16947;
  assign n16949 = po57  & ~n16941;
  assign n16950 = ~n16948 & ~n16949;
  assign n16951 = po58  & ~n16950;
  assign n16952 = ~n16387 & ~n16389;
  assign n16953 = po5  & n16952;
  assign n16954 = n15908 & ~n16953;
  assign n16955 = ~n15908 & n16953;
  assign n16956 = ~n16954 & ~n16955;
  assign n16957 = ~po58  & ~n16949;
  assign n16958 = ~n16948 & n16957;
  assign n16959 = n16956 & ~n16958;
  assign n16960 = ~n16951 & ~n16959;
  assign n16961 = ~po59  & n16960;
  assign n16962 = po59  & ~n16960;
  assign n16963 = ~n16454 & ~n16961;
  assign n16964 = ~n16962 & ~n16963;
  assign n16965 = po60  & ~n16964;
  assign n16966 = ~po60  & ~n16962;
  assign n16967 = ~n16963 & n16966;
  assign n16968 = ~n16396 & po5 ;
  assign n16969 = ~n16402 & n16968;
  assign n16970 = n16401 & ~n16969;
  assign n16971 = n16403 & n16968;
  assign n16972 = ~n16970 & ~n16971;
  assign n16973 = ~n16967 & n16972;
  assign n16974 = ~n16965 & ~n16973;
  assign n16975 = po61  & ~n16974;
  assign n16976 = ~n16405 & ~n16407;
  assign n16977 = po5  & n16976;
  assign n16978 = n16412 & ~n16977;
  assign n16979 = ~n16412 & n16977;
  assign n16980 = ~n16978 & ~n16979;
  assign n16981 = ~po61  & n16974;
  assign n16982 = ~n16980 & ~n16981;
  assign n16983 = ~n16975 & ~n16982;
  assign n16984 = po62  & ~n16983;
  assign n16985 = ~po62  & ~n16975;
  assign n16986 = ~n16982 & n16985;
  assign n16987 = ~n16415 & po5 ;
  assign n16988 = ~n16421 & n16987;
  assign n16989 = n16420 & ~n16988;
  assign n16990 = n16422 & n16987;
  assign n16991 = ~n16989 & ~n16990;
  assign n16992 = ~n16986 & n16991;
  assign n16993 = ~n16984 & ~n16992;
  assign n16994 = n16442 & po5 ;
  assign n16995 = ~n16433 & n16994;
  assign n16996 = ~n16424 & ~n16426;
  assign n16997 = po5  & n16996;
  assign n16998 = n16431 & ~n16997;
  assign n16999 = ~n16431 & n16997;
  assign n17000 = ~n16998 & ~n16999;
  assign n17001 = ~n16446 & ~n16995;
  assign n17002 = ~n17000 & n17001;
  assign n17003 = ~n16993 & n17002;
  assign n17004 = ~po63  & ~n17003;
  assign n17005 = n16993 & n17000;
  assign n17006 = n16433 & ~n16994;
  assign n17007 = ~n16433 & n16442;
  assign n17008 = po63  & ~n17007;
  assign n17009 = ~n17006 & n17008;
  assign n17010 = ~n17005 & ~n17009;
  assign po4  = n17004 | ~n17010;
  assign n17012 = ~n16962 & po4 ;
  assign n17013 = ~n16961 & n17012;
  assign n17014 = n16454 & ~n17013;
  assign n17015 = n16963 & n17012;
  assign n17016 = ~n17014 & ~n17015;
  assign n17017 = pi8  & po4 ;
  assign n17018 = ~pi6  & ~pi7 ;
  assign n17019 = ~pi8  & n17018;
  assign n17020 = ~n17017 & ~n17019;
  assign n17021 = po5  & ~n17020;
  assign n17022 = ~pi8  & po4 ;
  assign n17023 = pi9  & ~n17022;
  assign n17024 = ~pi9  & n17022;
  assign n17025 = ~n17023 & ~n17024;
  assign n17026 = ~po5  & n17020;
  assign n17027 = n17025 & ~n17026;
  assign n17028 = ~n17021 & ~n17027;
  assign n17029 = po6  & ~n17028;
  assign n17030 = ~po6  & ~n17021;
  assign n17031 = ~n17027 & n17030;
  assign n17032 = po5  & ~po4 ;
  assign n17033 = ~n17024 & ~n17032;
  assign n17034 = pi10  & ~n17033;
  assign n17035 = ~pi10  & n17033;
  assign n17036 = ~n17034 & ~n17035;
  assign n17037 = ~n17031 & ~n17036;
  assign n17038 = ~n17029 & ~n17037;
  assign n17039 = po7  & ~n17038;
  assign n17040 = ~po7  & n17038;
  assign n17041 = ~n16459 & ~n16460;
  assign n17042 = po4  & n17041;
  assign n17043 = n16464 & ~n17042;
  assign n17044 = ~n16464 & n17042;
  assign n17045 = ~n17043 & ~n17044;
  assign n17046 = ~n17040 & ~n17045;
  assign n17047 = ~n17039 & ~n17046;
  assign n17048 = po8  & ~n17047;
  assign n17049 = ~po8  & ~n17039;
  assign n17050 = ~n17046 & n17049;
  assign n17051 = ~n16467 & po4 ;
  assign n17052 = ~n16473 & n17051;
  assign n17053 = n16472 & ~n17052;
  assign n17054 = n16474 & n17051;
  assign n17055 = ~n17053 & ~n17054;
  assign n17056 = ~n17050 & n17055;
  assign n17057 = ~n17048 & ~n17056;
  assign n17058 = po9  & ~n17057;
  assign n17059 = ~po9  & n17057;
  assign n17060 = ~n16476 & ~n16478;
  assign n17061 = po4  & n17060;
  assign n17062 = n16483 & ~n17061;
  assign n17063 = ~n16483 & n17061;
  assign n17064 = ~n17062 & ~n17063;
  assign n17065 = ~n17059 & n17064;
  assign n17066 = ~n17058 & ~n17065;
  assign n17067 = po10  & ~n17066;
  assign n17068 = ~po10  & ~n17058;
  assign n17069 = ~n17065 & n17068;
  assign n17070 = ~n16486 & po4 ;
  assign n17071 = ~n16492 & n17070;
  assign n17072 = n16491 & ~n17071;
  assign n17073 = n16493 & n17070;
  assign n17074 = ~n17072 & ~n17073;
  assign n17075 = ~n17069 & n17074;
  assign n17076 = ~n17067 & ~n17075;
  assign n17077 = po11  & ~n17076;
  assign n17078 = ~po11  & n17076;
  assign n17079 = ~n16495 & ~n16497;
  assign n17080 = po4  & n17079;
  assign n17081 = n16502 & n17080;
  assign n17082 = ~n16502 & ~n17080;
  assign n17083 = ~n17081 & ~n17082;
  assign n17084 = ~n17078 & n17083;
  assign n17085 = ~n17077 & ~n17084;
  assign n17086 = po12  & ~n17085;
  assign n17087 = ~po12  & ~n17077;
  assign n17088 = ~n17084 & n17087;
  assign n17089 = ~n16505 & po4 ;
  assign n17090 = ~n16511 & n17089;
  assign n17091 = n16510 & ~n17090;
  assign n17092 = n16512 & n17089;
  assign n17093 = ~n17091 & ~n17092;
  assign n17094 = ~n17088 & n17093;
  assign n17095 = ~n17086 & ~n17094;
  assign n17096 = po13  & ~n17095;
  assign n17097 = ~po13  & n17095;
  assign n17098 = ~n16514 & ~n16516;
  assign n17099 = po4  & n17098;
  assign n17100 = ~n16521 & ~n17099;
  assign n17101 = n16521 & n17099;
  assign n17102 = ~n17100 & ~n17101;
  assign n17103 = ~n17097 & n17102;
  assign n17104 = ~n17096 & ~n17103;
  assign n17105 = po14  & ~n17104;
  assign n17106 = ~po14  & ~n17096;
  assign n17107 = ~n17103 & n17106;
  assign n17108 = ~n16524 & po4 ;
  assign n17109 = ~n16530 & n17108;
  assign n17110 = n16529 & ~n17109;
  assign n17111 = n16531 & n17108;
  assign n17112 = ~n17110 & ~n17111;
  assign n17113 = ~n17107 & n17112;
  assign n17114 = ~n17105 & ~n17113;
  assign n17115 = po15  & ~n17114;
  assign n17116 = ~n16533 & ~n16535;
  assign n17117 = po4  & n17116;
  assign n17118 = n16540 & ~n17117;
  assign n17119 = ~n16540 & n17117;
  assign n17120 = ~n17118 & ~n17119;
  assign n17121 = ~po15  & n17114;
  assign n17122 = ~n17120 & ~n17121;
  assign n17123 = ~n17115 & ~n17122;
  assign n17124 = po16  & ~n17123;
  assign n17125 = ~po16  & ~n17115;
  assign n17126 = ~n17122 & n17125;
  assign n17127 = ~n16543 & po4 ;
  assign n17128 = ~n16549 & n17127;
  assign n17129 = n16548 & ~n17128;
  assign n17130 = n16550 & n17127;
  assign n17131 = ~n17129 & ~n17130;
  assign n17132 = ~n17126 & n17131;
  assign n17133 = ~n17124 & ~n17132;
  assign n17134 = po17  & ~n17133;
  assign n17135 = ~po17  & n17133;
  assign n17136 = ~n16552 & po4 ;
  assign n17137 = ~n16559 & n17136;
  assign n17138 = n16557 & ~n17137;
  assign n17139 = n16560 & n17136;
  assign n17140 = ~n17138 & ~n17139;
  assign n17141 = ~n17135 & n17140;
  assign n17142 = ~n17134 & ~n17141;
  assign n17143 = po18  & ~n17142;
  assign n17144 = ~po18  & ~n17134;
  assign n17145 = ~n17141 & n17144;
  assign n17146 = ~n16562 & po4 ;
  assign n17147 = ~n16568 & n17146;
  assign n17148 = n16567 & ~n17147;
  assign n17149 = n16569 & n17146;
  assign n17150 = ~n17148 & ~n17149;
  assign n17151 = ~n17145 & n17150;
  assign n17152 = ~n17143 & ~n17151;
  assign n17153 = po19  & ~n17152;
  assign n17154 = ~n16571 & ~n16573;
  assign n17155 = po4  & n17154;
  assign n17156 = n16578 & ~n17155;
  assign n17157 = ~n16578 & n17155;
  assign n17158 = ~n17156 & ~n17157;
  assign n17159 = ~po19  & n17152;
  assign n17160 = ~n17158 & ~n17159;
  assign n17161 = ~n17153 & ~n17160;
  assign n17162 = po20  & ~n17161;
  assign n17163 = ~po20  & ~n17153;
  assign n17164 = ~n17160 & n17163;
  assign n17165 = ~n16581 & po4 ;
  assign n17166 = ~n16587 & n17165;
  assign n17167 = n16586 & ~n17166;
  assign n17168 = n16588 & n17165;
  assign n17169 = ~n17167 & ~n17168;
  assign n17170 = ~n17164 & n17169;
  assign n17171 = ~n17162 & ~n17170;
  assign n17172 = po21  & ~n17171;
  assign n17173 = ~po21  & n17171;
  assign n17174 = ~n16590 & po4 ;
  assign n17175 = ~n16597 & n17174;
  assign n17176 = n16595 & ~n17175;
  assign n17177 = n16598 & n17174;
  assign n17178 = ~n17176 & ~n17177;
  assign n17179 = ~n17173 & n17178;
  assign n17180 = ~n17172 & ~n17179;
  assign n17181 = po22  & ~n17180;
  assign n17182 = ~po22  & ~n17172;
  assign n17183 = ~n17179 & n17182;
  assign n17184 = ~n16600 & po4 ;
  assign n17185 = ~n16606 & n17184;
  assign n17186 = n16605 & ~n17185;
  assign n17187 = n16607 & n17184;
  assign n17188 = ~n17186 & ~n17187;
  assign n17189 = ~n17183 & n17188;
  assign n17190 = ~n17181 & ~n17189;
  assign n17191 = po23  & ~n17190;
  assign n17192 = ~n16609 & ~n16611;
  assign n17193 = po4  & n17192;
  assign n17194 = n16616 & ~n17193;
  assign n17195 = ~n16616 & n17193;
  assign n17196 = ~n17194 & ~n17195;
  assign n17197 = ~po23  & n17190;
  assign n17198 = ~n17196 & ~n17197;
  assign n17199 = ~n17191 & ~n17198;
  assign n17200 = po24  & ~n17199;
  assign n17201 = ~po24  & ~n17191;
  assign n17202 = ~n17198 & n17201;
  assign n17203 = ~n16619 & po4 ;
  assign n17204 = ~n16625 & n17203;
  assign n17205 = n16624 & ~n17204;
  assign n17206 = n16626 & n17203;
  assign n17207 = ~n17205 & ~n17206;
  assign n17208 = ~n17202 & n17207;
  assign n17209 = ~n17200 & ~n17208;
  assign n17210 = po25  & ~n17209;
  assign n17211 = ~po25  & n17209;
  assign n17212 = ~n16628 & po4 ;
  assign n17213 = ~n16635 & n17212;
  assign n17214 = n16633 & ~n17213;
  assign n17215 = n16636 & n17212;
  assign n17216 = ~n17214 & ~n17215;
  assign n17217 = ~n17211 & n17216;
  assign n17218 = ~n17210 & ~n17217;
  assign n17219 = po26  & ~n17218;
  assign n17220 = ~po26  & ~n17210;
  assign n17221 = ~n17217 & n17220;
  assign n17222 = ~n16638 & po4 ;
  assign n17223 = ~n16644 & n17222;
  assign n17224 = n16643 & ~n17223;
  assign n17225 = n16645 & n17222;
  assign n17226 = ~n17224 & ~n17225;
  assign n17227 = ~n17221 & n17226;
  assign n17228 = ~n17219 & ~n17227;
  assign n17229 = po27  & ~n17228;
  assign n17230 = ~n16647 & ~n16649;
  assign n17231 = po4  & n17230;
  assign n17232 = n16654 & ~n17231;
  assign n17233 = ~n16654 & n17231;
  assign n17234 = ~n17232 & ~n17233;
  assign n17235 = ~po27  & n17228;
  assign n17236 = ~n17234 & ~n17235;
  assign n17237 = ~n17229 & ~n17236;
  assign n17238 = po28  & ~n17237;
  assign n17239 = ~po28  & ~n17229;
  assign n17240 = ~n17236 & n17239;
  assign n17241 = ~n16657 & po4 ;
  assign n17242 = ~n16663 & n17241;
  assign n17243 = n16662 & ~n17242;
  assign n17244 = n16664 & n17241;
  assign n17245 = ~n17243 & ~n17244;
  assign n17246 = ~n17240 & n17245;
  assign n17247 = ~n17238 & ~n17246;
  assign n17248 = po29  & ~n17247;
  assign n17249 = ~po29  & n17247;
  assign n17250 = ~n16666 & po4 ;
  assign n17251 = ~n16673 & n17250;
  assign n17252 = n16671 & ~n17251;
  assign n17253 = n16674 & n17250;
  assign n17254 = ~n17252 & ~n17253;
  assign n17255 = ~n17249 & n17254;
  assign n17256 = ~n17248 & ~n17255;
  assign n17257 = po30  & ~n17256;
  assign n17258 = ~po30  & ~n17248;
  assign n17259 = ~n17255 & n17258;
  assign n17260 = ~n16676 & po4 ;
  assign n17261 = ~n16682 & n17260;
  assign n17262 = n16681 & ~n17261;
  assign n17263 = n16683 & n17260;
  assign n17264 = ~n17262 & ~n17263;
  assign n17265 = ~n17259 & n17264;
  assign n17266 = ~n17257 & ~n17265;
  assign n17267 = po31  & ~n17266;
  assign n17268 = ~n16685 & ~n16687;
  assign n17269 = po4  & n17268;
  assign n17270 = n16692 & ~n17269;
  assign n17271 = ~n16692 & n17269;
  assign n17272 = ~n17270 & ~n17271;
  assign n17273 = ~po31  & n17266;
  assign n17274 = ~n17272 & ~n17273;
  assign n17275 = ~n17267 & ~n17274;
  assign n17276 = po32  & ~n17275;
  assign n17277 = ~po32  & ~n17267;
  assign n17278 = ~n17274 & n17277;
  assign n17279 = ~n16695 & po4 ;
  assign n17280 = ~n16701 & n17279;
  assign n17281 = n16700 & ~n17280;
  assign n17282 = n16702 & n17279;
  assign n17283 = ~n17281 & ~n17282;
  assign n17284 = ~n17278 & n17283;
  assign n17285 = ~n17276 & ~n17284;
  assign n17286 = po33  & ~n17285;
  assign n17287 = ~po33  & n17285;
  assign n17288 = ~n16704 & po4 ;
  assign n17289 = ~n16711 & n17288;
  assign n17290 = n16709 & ~n17289;
  assign n17291 = n16712 & n17288;
  assign n17292 = ~n17290 & ~n17291;
  assign n17293 = ~n17287 & n17292;
  assign n17294 = ~n17286 & ~n17293;
  assign n17295 = po34  & ~n17294;
  assign n17296 = ~po34  & ~n17286;
  assign n17297 = ~n17293 & n17296;
  assign n17298 = ~n16714 & po4 ;
  assign n17299 = ~n16720 & n17298;
  assign n17300 = n16719 & ~n17299;
  assign n17301 = n16721 & n17298;
  assign n17302 = ~n17300 & ~n17301;
  assign n17303 = ~n17297 & n17302;
  assign n17304 = ~n17295 & ~n17303;
  assign n17305 = po35  & ~n17304;
  assign n17306 = ~n16723 & ~n16725;
  assign n17307 = po4  & n17306;
  assign n17308 = n16730 & ~n17307;
  assign n17309 = ~n16730 & n17307;
  assign n17310 = ~n17308 & ~n17309;
  assign n17311 = ~po35  & n17304;
  assign n17312 = ~n17310 & ~n17311;
  assign n17313 = ~n17305 & ~n17312;
  assign n17314 = po36  & ~n17313;
  assign n17315 = ~po36  & ~n17305;
  assign n17316 = ~n17312 & n17315;
  assign n17317 = ~n16733 & po4 ;
  assign n17318 = ~n16739 & n17317;
  assign n17319 = n16738 & ~n17318;
  assign n17320 = n16740 & n17317;
  assign n17321 = ~n17319 & ~n17320;
  assign n17322 = ~n17316 & n17321;
  assign n17323 = ~n17314 & ~n17322;
  assign n17324 = po37  & ~n17323;
  assign n17325 = ~po37  & n17323;
  assign n17326 = ~n16742 & po4 ;
  assign n17327 = ~n16749 & n17326;
  assign n17328 = n16747 & ~n17327;
  assign n17329 = n16750 & n17326;
  assign n17330 = ~n17328 & ~n17329;
  assign n17331 = ~n17325 & n17330;
  assign n17332 = ~n17324 & ~n17331;
  assign n17333 = po38  & ~n17332;
  assign n17334 = ~po38  & ~n17324;
  assign n17335 = ~n17331 & n17334;
  assign n17336 = ~n16752 & po4 ;
  assign n17337 = ~n16758 & n17336;
  assign n17338 = n16757 & ~n17337;
  assign n17339 = n16759 & n17336;
  assign n17340 = ~n17338 & ~n17339;
  assign n17341 = ~n17335 & n17340;
  assign n17342 = ~n17333 & ~n17341;
  assign n17343 = po39  & ~n17342;
  assign n17344 = ~n16761 & ~n16763;
  assign n17345 = po4  & n17344;
  assign n17346 = n16768 & ~n17345;
  assign n17347 = ~n16768 & n17345;
  assign n17348 = ~n17346 & ~n17347;
  assign n17349 = ~po39  & n17342;
  assign n17350 = ~n17348 & ~n17349;
  assign n17351 = ~n17343 & ~n17350;
  assign n17352 = po40  & ~n17351;
  assign n17353 = ~po40  & ~n17343;
  assign n17354 = ~n17350 & n17353;
  assign n17355 = ~n16771 & po4 ;
  assign n17356 = ~n16777 & n17355;
  assign n17357 = n16776 & ~n17356;
  assign n17358 = n16778 & n17355;
  assign n17359 = ~n17357 & ~n17358;
  assign n17360 = ~n17354 & n17359;
  assign n17361 = ~n17352 & ~n17360;
  assign n17362 = po41  & ~n17361;
  assign n17363 = ~po41  & n17361;
  assign n17364 = ~n16780 & po4 ;
  assign n17365 = ~n16787 & n17364;
  assign n17366 = n16785 & ~n17365;
  assign n17367 = n16788 & n17364;
  assign n17368 = ~n17366 & ~n17367;
  assign n17369 = ~n17363 & n17368;
  assign n17370 = ~n17362 & ~n17369;
  assign n17371 = po42  & ~n17370;
  assign n17372 = ~po42  & ~n17362;
  assign n17373 = ~n17369 & n17372;
  assign n17374 = ~n16790 & po4 ;
  assign n17375 = ~n16796 & n17374;
  assign n17376 = n16795 & ~n17375;
  assign n17377 = n16797 & n17374;
  assign n17378 = ~n17376 & ~n17377;
  assign n17379 = ~n17373 & n17378;
  assign n17380 = ~n17371 & ~n17379;
  assign n17381 = po43  & ~n17380;
  assign n17382 = ~n16799 & ~n16801;
  assign n17383 = po4  & n17382;
  assign n17384 = n16806 & ~n17383;
  assign n17385 = ~n16806 & n17383;
  assign n17386 = ~n17384 & ~n17385;
  assign n17387 = ~po43  & n17380;
  assign n17388 = ~n17386 & ~n17387;
  assign n17389 = ~n17381 & ~n17388;
  assign n17390 = po44  & ~n17389;
  assign n17391 = ~po44  & ~n17381;
  assign n17392 = ~n17388 & n17391;
  assign n17393 = ~n16809 & po4 ;
  assign n17394 = ~n16815 & n17393;
  assign n17395 = n16814 & ~n17394;
  assign n17396 = n16816 & n17393;
  assign n17397 = ~n17395 & ~n17396;
  assign n17398 = ~n17392 & n17397;
  assign n17399 = ~n17390 & ~n17398;
  assign n17400 = po45  & ~n17399;
  assign n17401 = ~po45  & n17399;
  assign n17402 = ~n16818 & po4 ;
  assign n17403 = ~n16825 & n17402;
  assign n17404 = n16823 & ~n17403;
  assign n17405 = n16826 & n17402;
  assign n17406 = ~n17404 & ~n17405;
  assign n17407 = ~n17401 & n17406;
  assign n17408 = ~n17400 & ~n17407;
  assign n17409 = po46  & ~n17408;
  assign n17410 = ~po46  & ~n17400;
  assign n17411 = ~n17407 & n17410;
  assign n17412 = ~n16828 & po4 ;
  assign n17413 = ~n16834 & n17412;
  assign n17414 = n16833 & ~n17413;
  assign n17415 = n16835 & n17412;
  assign n17416 = ~n17414 & ~n17415;
  assign n17417 = ~n17411 & n17416;
  assign n17418 = ~n17409 & ~n17417;
  assign n17419 = po47  & ~n17418;
  assign n17420 = ~n16837 & ~n16839;
  assign n17421 = po4  & n17420;
  assign n17422 = n16844 & ~n17421;
  assign n17423 = ~n16844 & n17421;
  assign n17424 = ~n17422 & ~n17423;
  assign n17425 = ~po47  & n17418;
  assign n17426 = ~n17424 & ~n17425;
  assign n17427 = ~n17419 & ~n17426;
  assign n17428 = po48  & ~n17427;
  assign n17429 = ~po48  & ~n17419;
  assign n17430 = ~n17426 & n17429;
  assign n17431 = ~n16847 & po4 ;
  assign n17432 = ~n16853 & n17431;
  assign n17433 = n16852 & ~n17432;
  assign n17434 = n16854 & n17431;
  assign n17435 = ~n17433 & ~n17434;
  assign n17436 = ~n17430 & n17435;
  assign n17437 = ~n17428 & ~n17436;
  assign n17438 = po49  & ~n17437;
  assign n17439 = ~po49  & n17437;
  assign n17440 = ~n16856 & po4 ;
  assign n17441 = ~n16863 & n17440;
  assign n17442 = n16861 & ~n17441;
  assign n17443 = n16864 & n17440;
  assign n17444 = ~n17442 & ~n17443;
  assign n17445 = ~n17439 & n17444;
  assign n17446 = ~n17438 & ~n17445;
  assign n17447 = po50  & ~n17446;
  assign n17448 = ~po50  & ~n17438;
  assign n17449 = ~n17445 & n17448;
  assign n17450 = ~n16866 & po4 ;
  assign n17451 = ~n16872 & n17450;
  assign n17452 = n16871 & ~n17451;
  assign n17453 = n16873 & n17450;
  assign n17454 = ~n17452 & ~n17453;
  assign n17455 = ~n17449 & n17454;
  assign n17456 = ~n17447 & ~n17455;
  assign n17457 = po51  & ~n17456;
  assign n17458 = ~n16875 & ~n16877;
  assign n17459 = po4  & n17458;
  assign n17460 = n16882 & ~n17459;
  assign n17461 = ~n16882 & n17459;
  assign n17462 = ~n17460 & ~n17461;
  assign n17463 = ~po51  & n17456;
  assign n17464 = ~n17462 & ~n17463;
  assign n17465 = ~n17457 & ~n17464;
  assign n17466 = po52  & ~n17465;
  assign n17467 = ~po52  & ~n17457;
  assign n17468 = ~n17464 & n17467;
  assign n17469 = ~n16885 & po4 ;
  assign n17470 = ~n16891 & n17469;
  assign n17471 = n16890 & ~n17470;
  assign n17472 = n16892 & n17469;
  assign n17473 = ~n17471 & ~n17472;
  assign n17474 = ~n17468 & n17473;
  assign n17475 = ~n17466 & ~n17474;
  assign n17476 = po53  & ~n17475;
  assign n17477 = ~po53  & n17475;
  assign n17478 = ~n16894 & po4 ;
  assign n17479 = ~n16901 & n17478;
  assign n17480 = n16899 & ~n17479;
  assign n17481 = n16902 & n17478;
  assign n17482 = ~n17480 & ~n17481;
  assign n17483 = ~n17477 & n17482;
  assign n17484 = ~n17476 & ~n17483;
  assign n17485 = po54  & ~n17484;
  assign n17486 = ~po54  & ~n17476;
  assign n17487 = ~n17483 & n17486;
  assign n17488 = ~n16904 & po4 ;
  assign n17489 = ~n16910 & n17488;
  assign n17490 = n16909 & ~n17489;
  assign n17491 = n16911 & n17488;
  assign n17492 = ~n17490 & ~n17491;
  assign n17493 = ~n17487 & n17492;
  assign n17494 = ~n17485 & ~n17493;
  assign n17495 = po55  & ~n17494;
  assign n17496 = ~n16913 & ~n16915;
  assign n17497 = po4  & n17496;
  assign n17498 = n16920 & ~n17497;
  assign n17499 = ~n16920 & n17497;
  assign n17500 = ~n17498 & ~n17499;
  assign n17501 = ~po55  & n17494;
  assign n17502 = ~n17500 & ~n17501;
  assign n17503 = ~n17495 & ~n17502;
  assign n17504 = po56  & ~n17503;
  assign n17505 = ~po56  & ~n17495;
  assign n17506 = ~n17502 & n17505;
  assign n17507 = ~n16923 & po4 ;
  assign n17508 = ~n16929 & n17507;
  assign n17509 = n16928 & ~n17508;
  assign n17510 = n16930 & n17507;
  assign n17511 = ~n17509 & ~n17510;
  assign n17512 = ~n17506 & n17511;
  assign n17513 = ~n17504 & ~n17512;
  assign n17514 = po57  & ~n17513;
  assign n17515 = ~po57  & n17513;
  assign n17516 = ~n16932 & po4 ;
  assign n17517 = ~n16939 & n17516;
  assign n17518 = n16937 & ~n17517;
  assign n17519 = n16940 & n17516;
  assign n17520 = ~n17518 & ~n17519;
  assign n17521 = ~n17515 & n17520;
  assign n17522 = ~n17514 & ~n17521;
  assign n17523 = po58  & ~n17522;
  assign n17524 = ~n16942 & ~n16949;
  assign n17525 = po4  & n17524;
  assign n17526 = n16947 & ~n17525;
  assign n17527 = ~n16947 & n17525;
  assign n17528 = ~n17526 & ~n17527;
  assign n17529 = ~po58  & ~n17514;
  assign n17530 = ~n17521 & n17529;
  assign n17531 = ~n17528 & ~n17530;
  assign n17532 = ~n17523 & ~n17531;
  assign n17533 = ~po59  & n17532;
  assign n17534 = ~n16951 & ~n16958;
  assign n17535 = po4  & n17534;
  assign n17536 = n16956 & n17535;
  assign n17537 = ~n16956 & ~n17535;
  assign n17538 = ~n17536 & ~n17537;
  assign n17539 = ~n17533 & n17538;
  assign n17540 = po59  & ~n17532;
  assign n17541 = ~po60  & ~n17540;
  assign n17542 = ~n17539 & n17541;
  assign n17543 = ~n17539 & ~n17540;
  assign n17544 = po60  & ~n17543;
  assign n17545 = n17016 & ~n17542;
  assign n17546 = ~n17544 & ~n17545;
  assign n17547 = po61  & ~n17546;
  assign n17548 = ~n16965 & ~n16967;
  assign n17549 = po4  & n17548;
  assign n17550 = n16972 & ~n17549;
  assign n17551 = ~n16972 & n17549;
  assign n17552 = ~n17550 & ~n17551;
  assign n17553 = ~po61  & n17546;
  assign n17554 = ~n17552 & ~n17553;
  assign n17555 = ~n17547 & ~n17554;
  assign n17556 = po62  & ~n17555;
  assign n17557 = ~po62  & ~n17547;
  assign n17558 = ~n17554 & n17557;
  assign n17559 = ~n16975 & po4 ;
  assign n17560 = ~n16981 & n17559;
  assign n17561 = n16980 & ~n17560;
  assign n17562 = n16982 & n17559;
  assign n17563 = ~n17561 & ~n17562;
  assign n17564 = ~n17558 & n17563;
  assign n17565 = ~n17556 & ~n17564;
  assign n17566 = ~n16984 & ~n16986;
  assign n17567 = po4  & n17566;
  assign n17568 = n16991 & ~n17567;
  assign n17569 = ~n16991 & n17567;
  assign n17570 = ~n17568 & ~n17569;
  assign n17571 = n16993 & po4 ;
  assign n17572 = ~n17000 & ~n17571;
  assign n17573 = ~n17005 & ~n17572;
  assign n17574 = po4  & ~n17573;
  assign n17575 = ~n17570 & ~n17574;
  assign n17576 = ~n17565 & n17575;
  assign n17577 = ~po63  & ~n17576;
  assign n17578 = n17565 & n17570;
  assign n17579 = po63  & n17573;
  assign n17580 = ~n17578 & ~n17579;
  assign po3  = n17577 | ~n17580;
  assign n17582 = ~n17542 & ~n17544;
  assign n17583 = po3  & n17582;
  assign n17584 = n17016 & ~n17583;
  assign n17585 = ~n17016 & n17583;
  assign n17586 = ~n17584 & ~n17585;
  assign n17587 = pi6  & po3 ;
  assign n17588 = ~pi4  & ~pi5 ;
  assign n17589 = ~pi6  & n17588;
  assign n17590 = ~n17587 & ~n17589;
  assign n17591 = po4  & ~n17590;
  assign n17592 = ~po4  & n17590;
  assign n17593 = ~pi6  & po3 ;
  assign n17594 = pi7  & ~n17593;
  assign n17595 = ~pi7  & n17593;
  assign n17596 = ~n17594 & ~n17595;
  assign n17597 = ~n17592 & n17596;
  assign n17598 = ~n17591 & ~n17597;
  assign n17599 = po5  & ~n17598;
  assign n17600 = po4  & ~po3 ;
  assign n17601 = ~n17595 & ~n17600;
  assign n17602 = pi8  & ~n17601;
  assign n17603 = ~pi8  & n17601;
  assign n17604 = ~n17602 & ~n17603;
  assign n17605 = ~po5  & n17598;
  assign n17606 = ~n17604 & ~n17605;
  assign n17607 = ~n17599 & ~n17606;
  assign n17608 = po6  & ~n17607;
  assign n17609 = ~po6  & ~n17599;
  assign n17610 = ~n17606 & n17609;
  assign n17611 = ~n17021 & ~n17026;
  assign n17612 = po3  & n17611;
  assign n17613 = n17025 & ~n17612;
  assign n17614 = ~n17025 & n17612;
  assign n17615 = ~n17613 & ~n17614;
  assign n17616 = ~n17610 & ~n17615;
  assign n17617 = ~n17608 & ~n17616;
  assign n17618 = po7  & ~n17617;
  assign n17619 = ~n17029 & ~n17031;
  assign n17620 = po3  & n17619;
  assign n17621 = ~n17036 & ~n17620;
  assign n17622 = n17036 & n17620;
  assign n17623 = ~n17621 & ~n17622;
  assign n17624 = ~po7  & n17617;
  assign n17625 = ~n17623 & ~n17624;
  assign n17626 = ~n17618 & ~n17625;
  assign n17627 = po8  & ~n17626;
  assign n17628 = ~po8  & ~n17618;
  assign n17629 = ~n17625 & n17628;
  assign n17630 = ~n17039 & ~n17040;
  assign n17631 = po3  & n17630;
  assign n17632 = n17045 & ~n17631;
  assign n17633 = ~n17045 & n17631;
  assign n17634 = ~n17632 & ~n17633;
  assign n17635 = ~n17629 & n17634;
  assign n17636 = ~n17627 & ~n17635;
  assign n17637 = po9  & ~n17636;
  assign n17638 = ~n17048 & ~n17050;
  assign n17639 = po3  & n17638;
  assign n17640 = n17055 & ~n17639;
  assign n17641 = ~n17055 & n17639;
  assign n17642 = ~n17640 & ~n17641;
  assign n17643 = ~po9  & n17636;
  assign n17644 = ~n17642 & ~n17643;
  assign n17645 = ~n17637 & ~n17644;
  assign n17646 = po10  & ~n17645;
  assign n17647 = ~po10  & ~n17637;
  assign n17648 = ~n17644 & n17647;
  assign n17649 = ~n17058 & ~n17059;
  assign n17650 = po3  & n17649;
  assign n17651 = n17064 & n17650;
  assign n17652 = ~n17064 & ~n17650;
  assign n17653 = ~n17651 & ~n17652;
  assign n17654 = ~n17648 & n17653;
  assign n17655 = ~n17646 & ~n17654;
  assign n17656 = po11  & ~n17655;
  assign n17657 = ~n17067 & ~n17069;
  assign n17658 = po3  & n17657;
  assign n17659 = n17074 & ~n17658;
  assign n17660 = ~n17074 & n17658;
  assign n17661 = ~n17659 & ~n17660;
  assign n17662 = ~po11  & n17655;
  assign n17663 = ~n17661 & ~n17662;
  assign n17664 = ~n17656 & ~n17663;
  assign n17665 = po12  & ~n17664;
  assign n17666 = ~po12  & ~n17656;
  assign n17667 = ~n17663 & n17666;
  assign n17668 = ~n17077 & ~n17078;
  assign n17669 = po3  & n17668;
  assign n17670 = ~n17083 & ~n17669;
  assign n17671 = n17083 & n17669;
  assign n17672 = ~n17670 & ~n17671;
  assign n17673 = ~n17667 & n17672;
  assign n17674 = ~n17665 & ~n17673;
  assign n17675 = po13  & ~n17674;
  assign n17676 = ~n17086 & ~n17088;
  assign n17677 = po3  & n17676;
  assign n17678 = n17093 & ~n17677;
  assign n17679 = ~n17093 & n17677;
  assign n17680 = ~n17678 & ~n17679;
  assign n17681 = ~po13  & n17674;
  assign n17682 = ~n17680 & ~n17681;
  assign n17683 = ~n17675 & ~n17682;
  assign n17684 = po14  & ~n17683;
  assign n17685 = ~n17096 & ~n17097;
  assign n17686 = po3  & n17685;
  assign n17687 = n17102 & ~n17686;
  assign n17688 = ~n17102 & n17686;
  assign n17689 = ~n17687 & ~n17688;
  assign n17690 = ~po14  & ~n17675;
  assign n17691 = ~n17682 & n17690;
  assign n17692 = ~n17689 & ~n17691;
  assign n17693 = ~n17684 & ~n17692;
  assign n17694 = po15  & ~n17693;
  assign n17695 = ~n17105 & ~n17107;
  assign n17696 = po3  & n17695;
  assign n17697 = n17112 & ~n17696;
  assign n17698 = ~n17112 & n17696;
  assign n17699 = ~n17697 & ~n17698;
  assign n17700 = ~po15  & n17693;
  assign n17701 = ~n17699 & ~n17700;
  assign n17702 = ~n17694 & ~n17701;
  assign n17703 = po16  & ~n17702;
  assign n17704 = ~po16  & ~n17694;
  assign n17705 = ~n17701 & n17704;
  assign n17706 = ~n17115 & po3 ;
  assign n17707 = ~n17121 & n17706;
  assign n17708 = n17120 & ~n17707;
  assign n17709 = n17122 & n17706;
  assign n17710 = ~n17708 & ~n17709;
  assign n17711 = ~n17705 & n17710;
  assign n17712 = ~n17703 & ~n17711;
  assign n17713 = po17  & ~n17712;
  assign n17714 = ~n17124 & ~n17126;
  assign n17715 = po3  & n17714;
  assign n17716 = n17131 & ~n17715;
  assign n17717 = ~n17131 & n17715;
  assign n17718 = ~n17716 & ~n17717;
  assign n17719 = ~po17  & n17712;
  assign n17720 = ~n17718 & ~n17719;
  assign n17721 = ~n17713 & ~n17720;
  assign n17722 = po18  & ~n17721;
  assign n17723 = ~n17134 & ~n17135;
  assign n17724 = po3  & n17723;
  assign n17725 = n17140 & ~n17724;
  assign n17726 = ~n17140 & n17724;
  assign n17727 = ~n17725 & ~n17726;
  assign n17728 = ~po18  & ~n17713;
  assign n17729 = ~n17720 & n17728;
  assign n17730 = ~n17727 & ~n17729;
  assign n17731 = ~n17722 & ~n17730;
  assign n17732 = po19  & ~n17731;
  assign n17733 = ~n17143 & ~n17145;
  assign n17734 = po3  & n17733;
  assign n17735 = n17150 & ~n17734;
  assign n17736 = ~n17150 & n17734;
  assign n17737 = ~n17735 & ~n17736;
  assign n17738 = ~po19  & n17731;
  assign n17739 = ~n17737 & ~n17738;
  assign n17740 = ~n17732 & ~n17739;
  assign n17741 = po20  & ~n17740;
  assign n17742 = ~po20  & ~n17732;
  assign n17743 = ~n17739 & n17742;
  assign n17744 = ~n17153 & po3 ;
  assign n17745 = ~n17159 & n17744;
  assign n17746 = n17158 & ~n17745;
  assign n17747 = n17160 & n17744;
  assign n17748 = ~n17746 & ~n17747;
  assign n17749 = ~n17743 & n17748;
  assign n17750 = ~n17741 & ~n17749;
  assign n17751 = po21  & ~n17750;
  assign n17752 = ~n17162 & ~n17164;
  assign n17753 = po3  & n17752;
  assign n17754 = n17169 & ~n17753;
  assign n17755 = ~n17169 & n17753;
  assign n17756 = ~n17754 & ~n17755;
  assign n17757 = ~po21  & n17750;
  assign n17758 = ~n17756 & ~n17757;
  assign n17759 = ~n17751 & ~n17758;
  assign n17760 = po22  & ~n17759;
  assign n17761 = ~n17172 & ~n17173;
  assign n17762 = po3  & n17761;
  assign n17763 = n17178 & ~n17762;
  assign n17764 = ~n17178 & n17762;
  assign n17765 = ~n17763 & ~n17764;
  assign n17766 = ~po22  & ~n17751;
  assign n17767 = ~n17758 & n17766;
  assign n17768 = ~n17765 & ~n17767;
  assign n17769 = ~n17760 & ~n17768;
  assign n17770 = po23  & ~n17769;
  assign n17771 = ~n17181 & ~n17183;
  assign n17772 = po3  & n17771;
  assign n17773 = n17188 & ~n17772;
  assign n17774 = ~n17188 & n17772;
  assign n17775 = ~n17773 & ~n17774;
  assign n17776 = ~po23  & n17769;
  assign n17777 = ~n17775 & ~n17776;
  assign n17778 = ~n17770 & ~n17777;
  assign n17779 = po24  & ~n17778;
  assign n17780 = ~po24  & ~n17770;
  assign n17781 = ~n17777 & n17780;
  assign n17782 = ~n17191 & po3 ;
  assign n17783 = ~n17197 & n17782;
  assign n17784 = n17196 & ~n17783;
  assign n17785 = n17198 & n17782;
  assign n17786 = ~n17784 & ~n17785;
  assign n17787 = ~n17781 & n17786;
  assign n17788 = ~n17779 & ~n17787;
  assign n17789 = po25  & ~n17788;
  assign n17790 = ~n17200 & ~n17202;
  assign n17791 = po3  & n17790;
  assign n17792 = n17207 & ~n17791;
  assign n17793 = ~n17207 & n17791;
  assign n17794 = ~n17792 & ~n17793;
  assign n17795 = ~po25  & n17788;
  assign n17796 = ~n17794 & ~n17795;
  assign n17797 = ~n17789 & ~n17796;
  assign n17798 = po26  & ~n17797;
  assign n17799 = ~n17210 & ~n17211;
  assign n17800 = po3  & n17799;
  assign n17801 = n17216 & ~n17800;
  assign n17802 = ~n17216 & n17800;
  assign n17803 = ~n17801 & ~n17802;
  assign n17804 = ~po26  & ~n17789;
  assign n17805 = ~n17796 & n17804;
  assign n17806 = ~n17803 & ~n17805;
  assign n17807 = ~n17798 & ~n17806;
  assign n17808 = po27  & ~n17807;
  assign n17809 = ~n17219 & ~n17221;
  assign n17810 = po3  & n17809;
  assign n17811 = n17226 & ~n17810;
  assign n17812 = ~n17226 & n17810;
  assign n17813 = ~n17811 & ~n17812;
  assign n17814 = ~po27  & n17807;
  assign n17815 = ~n17813 & ~n17814;
  assign n17816 = ~n17808 & ~n17815;
  assign n17817 = po28  & ~n17816;
  assign n17818 = ~po28  & ~n17808;
  assign n17819 = ~n17815 & n17818;
  assign n17820 = ~n17229 & po3 ;
  assign n17821 = ~n17235 & n17820;
  assign n17822 = n17234 & ~n17821;
  assign n17823 = n17236 & n17820;
  assign n17824 = ~n17822 & ~n17823;
  assign n17825 = ~n17819 & n17824;
  assign n17826 = ~n17817 & ~n17825;
  assign n17827 = po29  & ~n17826;
  assign n17828 = ~n17238 & ~n17240;
  assign n17829 = po3  & n17828;
  assign n17830 = n17245 & ~n17829;
  assign n17831 = ~n17245 & n17829;
  assign n17832 = ~n17830 & ~n17831;
  assign n17833 = ~po29  & n17826;
  assign n17834 = ~n17832 & ~n17833;
  assign n17835 = ~n17827 & ~n17834;
  assign n17836 = po30  & ~n17835;
  assign n17837 = ~n17248 & ~n17249;
  assign n17838 = po3  & n17837;
  assign n17839 = n17254 & ~n17838;
  assign n17840 = ~n17254 & n17838;
  assign n17841 = ~n17839 & ~n17840;
  assign n17842 = ~po30  & ~n17827;
  assign n17843 = ~n17834 & n17842;
  assign n17844 = ~n17841 & ~n17843;
  assign n17845 = ~n17836 & ~n17844;
  assign n17846 = po31  & ~n17845;
  assign n17847 = ~n17257 & ~n17259;
  assign n17848 = po3  & n17847;
  assign n17849 = n17264 & ~n17848;
  assign n17850 = ~n17264 & n17848;
  assign n17851 = ~n17849 & ~n17850;
  assign n17852 = ~po31  & n17845;
  assign n17853 = ~n17851 & ~n17852;
  assign n17854 = ~n17846 & ~n17853;
  assign n17855 = po32  & ~n17854;
  assign n17856 = ~po32  & ~n17846;
  assign n17857 = ~n17853 & n17856;
  assign n17858 = ~n17267 & po3 ;
  assign n17859 = ~n17273 & n17858;
  assign n17860 = n17272 & ~n17859;
  assign n17861 = n17274 & n17858;
  assign n17862 = ~n17860 & ~n17861;
  assign n17863 = ~n17857 & n17862;
  assign n17864 = ~n17855 & ~n17863;
  assign n17865 = po33  & ~n17864;
  assign n17866 = ~n17276 & ~n17278;
  assign n17867 = po3  & n17866;
  assign n17868 = n17283 & ~n17867;
  assign n17869 = ~n17283 & n17867;
  assign n17870 = ~n17868 & ~n17869;
  assign n17871 = ~po33  & n17864;
  assign n17872 = ~n17870 & ~n17871;
  assign n17873 = ~n17865 & ~n17872;
  assign n17874 = po34  & ~n17873;
  assign n17875 = ~n17286 & ~n17287;
  assign n17876 = po3  & n17875;
  assign n17877 = n17292 & ~n17876;
  assign n17878 = ~n17292 & n17876;
  assign n17879 = ~n17877 & ~n17878;
  assign n17880 = ~po34  & ~n17865;
  assign n17881 = ~n17872 & n17880;
  assign n17882 = ~n17879 & ~n17881;
  assign n17883 = ~n17874 & ~n17882;
  assign n17884 = po35  & ~n17883;
  assign n17885 = ~n17295 & ~n17297;
  assign n17886 = po3  & n17885;
  assign n17887 = n17302 & ~n17886;
  assign n17888 = ~n17302 & n17886;
  assign n17889 = ~n17887 & ~n17888;
  assign n17890 = ~po35  & n17883;
  assign n17891 = ~n17889 & ~n17890;
  assign n17892 = ~n17884 & ~n17891;
  assign n17893 = po36  & ~n17892;
  assign n17894 = ~po36  & ~n17884;
  assign n17895 = ~n17891 & n17894;
  assign n17896 = ~n17305 & po3 ;
  assign n17897 = ~n17311 & n17896;
  assign n17898 = n17310 & ~n17897;
  assign n17899 = n17312 & n17896;
  assign n17900 = ~n17898 & ~n17899;
  assign n17901 = ~n17895 & n17900;
  assign n17902 = ~n17893 & ~n17901;
  assign n17903 = po37  & ~n17902;
  assign n17904 = ~n17314 & ~n17316;
  assign n17905 = po3  & n17904;
  assign n17906 = n17321 & ~n17905;
  assign n17907 = ~n17321 & n17905;
  assign n17908 = ~n17906 & ~n17907;
  assign n17909 = ~po37  & n17902;
  assign n17910 = ~n17908 & ~n17909;
  assign n17911 = ~n17903 & ~n17910;
  assign n17912 = po38  & ~n17911;
  assign n17913 = ~n17324 & ~n17325;
  assign n17914 = po3  & n17913;
  assign n17915 = n17330 & ~n17914;
  assign n17916 = ~n17330 & n17914;
  assign n17917 = ~n17915 & ~n17916;
  assign n17918 = ~po38  & ~n17903;
  assign n17919 = ~n17910 & n17918;
  assign n17920 = ~n17917 & ~n17919;
  assign n17921 = ~n17912 & ~n17920;
  assign n17922 = po39  & ~n17921;
  assign n17923 = ~n17333 & ~n17335;
  assign n17924 = po3  & n17923;
  assign n17925 = n17340 & ~n17924;
  assign n17926 = ~n17340 & n17924;
  assign n17927 = ~n17925 & ~n17926;
  assign n17928 = ~po39  & n17921;
  assign n17929 = ~n17927 & ~n17928;
  assign n17930 = ~n17922 & ~n17929;
  assign n17931 = po40  & ~n17930;
  assign n17932 = ~po40  & ~n17922;
  assign n17933 = ~n17929 & n17932;
  assign n17934 = ~n17343 & po3 ;
  assign n17935 = ~n17349 & n17934;
  assign n17936 = n17348 & ~n17935;
  assign n17937 = n17350 & n17934;
  assign n17938 = ~n17936 & ~n17937;
  assign n17939 = ~n17933 & n17938;
  assign n17940 = ~n17931 & ~n17939;
  assign n17941 = po41  & ~n17940;
  assign n17942 = ~n17352 & ~n17354;
  assign n17943 = po3  & n17942;
  assign n17944 = n17359 & ~n17943;
  assign n17945 = ~n17359 & n17943;
  assign n17946 = ~n17944 & ~n17945;
  assign n17947 = ~po41  & n17940;
  assign n17948 = ~n17946 & ~n17947;
  assign n17949 = ~n17941 & ~n17948;
  assign n17950 = po42  & ~n17949;
  assign n17951 = ~n17362 & ~n17363;
  assign n17952 = po3  & n17951;
  assign n17953 = n17368 & ~n17952;
  assign n17954 = ~n17368 & n17952;
  assign n17955 = ~n17953 & ~n17954;
  assign n17956 = ~po42  & ~n17941;
  assign n17957 = ~n17948 & n17956;
  assign n17958 = ~n17955 & ~n17957;
  assign n17959 = ~n17950 & ~n17958;
  assign n17960 = po43  & ~n17959;
  assign n17961 = ~n17371 & ~n17373;
  assign n17962 = po3  & n17961;
  assign n17963 = n17378 & ~n17962;
  assign n17964 = ~n17378 & n17962;
  assign n17965 = ~n17963 & ~n17964;
  assign n17966 = ~po43  & n17959;
  assign n17967 = ~n17965 & ~n17966;
  assign n17968 = ~n17960 & ~n17967;
  assign n17969 = po44  & ~n17968;
  assign n17970 = ~po44  & ~n17960;
  assign n17971 = ~n17967 & n17970;
  assign n17972 = ~n17381 & po3 ;
  assign n17973 = ~n17387 & n17972;
  assign n17974 = n17386 & ~n17973;
  assign n17975 = n17388 & n17972;
  assign n17976 = ~n17974 & ~n17975;
  assign n17977 = ~n17971 & n17976;
  assign n17978 = ~n17969 & ~n17977;
  assign n17979 = po45  & ~n17978;
  assign n17980 = ~n17390 & ~n17392;
  assign n17981 = po3  & n17980;
  assign n17982 = n17397 & ~n17981;
  assign n17983 = ~n17397 & n17981;
  assign n17984 = ~n17982 & ~n17983;
  assign n17985 = ~po45  & n17978;
  assign n17986 = ~n17984 & ~n17985;
  assign n17987 = ~n17979 & ~n17986;
  assign n17988 = po46  & ~n17987;
  assign n17989 = ~n17400 & ~n17401;
  assign n17990 = po3  & n17989;
  assign n17991 = n17406 & ~n17990;
  assign n17992 = ~n17406 & n17990;
  assign n17993 = ~n17991 & ~n17992;
  assign n17994 = ~po46  & ~n17979;
  assign n17995 = ~n17986 & n17994;
  assign n17996 = ~n17993 & ~n17995;
  assign n17997 = ~n17988 & ~n17996;
  assign n17998 = po47  & ~n17997;
  assign n17999 = ~n17409 & ~n17411;
  assign n18000 = po3  & n17999;
  assign n18001 = n17416 & ~n18000;
  assign n18002 = ~n17416 & n18000;
  assign n18003 = ~n18001 & ~n18002;
  assign n18004 = ~po47  & n17997;
  assign n18005 = ~n18003 & ~n18004;
  assign n18006 = ~n17998 & ~n18005;
  assign n18007 = po48  & ~n18006;
  assign n18008 = ~po48  & ~n17998;
  assign n18009 = ~n18005 & n18008;
  assign n18010 = ~n17419 & po3 ;
  assign n18011 = ~n17425 & n18010;
  assign n18012 = n17424 & ~n18011;
  assign n18013 = n17426 & n18010;
  assign n18014 = ~n18012 & ~n18013;
  assign n18015 = ~n18009 & n18014;
  assign n18016 = ~n18007 & ~n18015;
  assign n18017 = po49  & ~n18016;
  assign n18018 = ~n17428 & ~n17430;
  assign n18019 = po3  & n18018;
  assign n18020 = n17435 & ~n18019;
  assign n18021 = ~n17435 & n18019;
  assign n18022 = ~n18020 & ~n18021;
  assign n18023 = ~po49  & n18016;
  assign n18024 = ~n18022 & ~n18023;
  assign n18025 = ~n18017 & ~n18024;
  assign n18026 = po50  & ~n18025;
  assign n18027 = ~n17438 & ~n17439;
  assign n18028 = po3  & n18027;
  assign n18029 = n17444 & ~n18028;
  assign n18030 = ~n17444 & n18028;
  assign n18031 = ~n18029 & ~n18030;
  assign n18032 = ~po50  & ~n18017;
  assign n18033 = ~n18024 & n18032;
  assign n18034 = ~n18031 & ~n18033;
  assign n18035 = ~n18026 & ~n18034;
  assign n18036 = po51  & ~n18035;
  assign n18037 = ~n17447 & ~n17449;
  assign n18038 = po3  & n18037;
  assign n18039 = n17454 & ~n18038;
  assign n18040 = ~n17454 & n18038;
  assign n18041 = ~n18039 & ~n18040;
  assign n18042 = ~po51  & n18035;
  assign n18043 = ~n18041 & ~n18042;
  assign n18044 = ~n18036 & ~n18043;
  assign n18045 = po52  & ~n18044;
  assign n18046 = ~po52  & ~n18036;
  assign n18047 = ~n18043 & n18046;
  assign n18048 = ~n17457 & po3 ;
  assign n18049 = ~n17463 & n18048;
  assign n18050 = n17462 & ~n18049;
  assign n18051 = n17464 & n18048;
  assign n18052 = ~n18050 & ~n18051;
  assign n18053 = ~n18047 & n18052;
  assign n18054 = ~n18045 & ~n18053;
  assign n18055 = po53  & ~n18054;
  assign n18056 = ~n17466 & ~n17468;
  assign n18057 = po3  & n18056;
  assign n18058 = n17473 & ~n18057;
  assign n18059 = ~n17473 & n18057;
  assign n18060 = ~n18058 & ~n18059;
  assign n18061 = ~po53  & n18054;
  assign n18062 = ~n18060 & ~n18061;
  assign n18063 = ~n18055 & ~n18062;
  assign n18064 = po54  & ~n18063;
  assign n18065 = ~n17476 & ~n17477;
  assign n18066 = po3  & n18065;
  assign n18067 = n17482 & ~n18066;
  assign n18068 = ~n17482 & n18066;
  assign n18069 = ~n18067 & ~n18068;
  assign n18070 = ~po54  & ~n18055;
  assign n18071 = ~n18062 & n18070;
  assign n18072 = ~n18069 & ~n18071;
  assign n18073 = ~n18064 & ~n18072;
  assign n18074 = po55  & ~n18073;
  assign n18075 = ~n17485 & ~n17487;
  assign n18076 = po3  & n18075;
  assign n18077 = n17492 & ~n18076;
  assign n18078 = ~n17492 & n18076;
  assign n18079 = ~n18077 & ~n18078;
  assign n18080 = ~po55  & n18073;
  assign n18081 = ~n18079 & ~n18080;
  assign n18082 = ~n18074 & ~n18081;
  assign n18083 = po56  & ~n18082;
  assign n18084 = ~po56  & ~n18074;
  assign n18085 = ~n18081 & n18084;
  assign n18086 = ~n17495 & po3 ;
  assign n18087 = ~n17501 & n18086;
  assign n18088 = n17500 & ~n18087;
  assign n18089 = n17502 & n18086;
  assign n18090 = ~n18088 & ~n18089;
  assign n18091 = ~n18085 & n18090;
  assign n18092 = ~n18083 & ~n18091;
  assign n18093 = po57  & ~n18092;
  assign n18094 = ~n17504 & ~n17506;
  assign n18095 = po3  & n18094;
  assign n18096 = n17511 & ~n18095;
  assign n18097 = ~n17511 & n18095;
  assign n18098 = ~n18096 & ~n18097;
  assign n18099 = ~po57  & n18092;
  assign n18100 = ~n18098 & ~n18099;
  assign n18101 = ~n18093 & ~n18100;
  assign n18102 = po58  & ~n18101;
  assign n18103 = ~n17514 & ~n17515;
  assign n18104 = po3  & n18103;
  assign n18105 = n17520 & ~n18104;
  assign n18106 = ~n17520 & n18104;
  assign n18107 = ~n18105 & ~n18106;
  assign n18108 = ~po58  & ~n18093;
  assign n18109 = ~n18100 & n18108;
  assign n18110 = ~n18107 & ~n18109;
  assign n18111 = ~n18102 & ~n18110;
  assign n18112 = ~po59  & n18111;
  assign n18113 = ~n17523 & po3 ;
  assign n18114 = ~n17530 & n18113;
  assign n18115 = n17528 & ~n18114;
  assign n18116 = n17531 & n18113;
  assign n18117 = ~n18115 & ~n18116;
  assign n18118 = ~n18112 & n18117;
  assign n18119 = po59  & ~n18111;
  assign n18120 = ~n18118 & ~n18119;
  assign n18121 = po60  & ~n18120;
  assign n18122 = ~n17533 & ~n17540;
  assign n18123 = po3  & n18122;
  assign n18124 = ~n17538 & ~n18123;
  assign n18125 = n17538 & n18123;
  assign n18126 = ~n18124 & ~n18125;
  assign n18127 = ~po60  & ~n18119;
  assign n18128 = ~n18118 & n18127;
  assign n18129 = n18126 & ~n18128;
  assign n18130 = ~n18121 & ~n18129;
  assign n18131 = ~po61  & n18130;
  assign n18132 = po61  & ~n18130;
  assign n18133 = ~n17586 & ~n18131;
  assign n18134 = ~n18132 & ~n18133;
  assign n18135 = po62  & ~n18134;
  assign n18136 = ~po62  & ~n18132;
  assign n18137 = ~n18133 & n18136;
  assign n18138 = ~n17547 & po3 ;
  assign n18139 = ~n17553 & n18138;
  assign n18140 = n17552 & ~n18139;
  assign n18141 = n17554 & n18138;
  assign n18142 = ~n18140 & ~n18141;
  assign n18143 = ~n18137 & n18142;
  assign n18144 = ~n18135 & ~n18143;
  assign n18145 = ~n17556 & ~n17558;
  assign n18146 = po3  & n18145;
  assign n18147 = n17563 & ~n18146;
  assign n18148 = ~n17563 & n18146;
  assign n18149 = ~n18147 & ~n18148;
  assign n18150 = n17565 & po3 ;
  assign n18151 = ~n17570 & ~n18150;
  assign n18152 = ~n17578 & ~n18151;
  assign n18153 = po3  & ~n18152;
  assign n18154 = ~n18149 & ~n18153;
  assign n18155 = ~n18144 & n18154;
  assign n18156 = ~po63  & ~n18155;
  assign n18157 = n18144 & n18149;
  assign n18158 = po63  & n18152;
  assign n18159 = ~n18157 & ~n18158;
  assign po2  = n18156 | ~n18159;
  assign n18161 = ~n18132 & po2 ;
  assign n18162 = ~n18131 & n18161;
  assign n18163 = n17586 & ~n18162;
  assign n18164 = n18133 & n18161;
  assign n18165 = ~n18163 & ~n18164;
  assign n18166 = ~n18121 & ~n18128;
  assign n18167 = po2  & n18166;
  assign n18168 = n18126 & ~n18167;
  assign n18169 = ~n18126 & n18167;
  assign n18170 = ~n18168 & ~n18169;
  assign n18171 = pi4  & po2 ;
  assign n18172 = ~pi2  & ~pi3 ;
  assign n18173 = ~pi4  & n18172;
  assign n18174 = ~n18171 & ~n18173;
  assign n18175 = po3  & ~n18174;
  assign n18176 = ~pi4  & po2 ;
  assign n18177 = pi5  & ~n18176;
  assign n18178 = ~pi5  & n18176;
  assign n18179 = ~n18177 & ~n18178;
  assign n18180 = ~po3  & n18174;
  assign n18181 = n18179 & ~n18180;
  assign n18182 = ~n18175 & ~n18181;
  assign n18183 = po4  & ~n18182;
  assign n18184 = ~po4  & ~n18175;
  assign n18185 = ~n18181 & n18184;
  assign n18186 = po3  & ~po2 ;
  assign n18187 = ~n18178 & ~n18186;
  assign n18188 = pi6  & ~n18187;
  assign n18189 = ~pi6  & n18187;
  assign n18190 = ~n18188 & ~n18189;
  assign n18191 = ~n18185 & ~n18190;
  assign n18192 = ~n18183 & ~n18191;
  assign n18193 = po5  & ~n18192;
  assign n18194 = ~po5  & n18192;
  assign n18195 = ~n17591 & ~n17592;
  assign n18196 = po2  & n18195;
  assign n18197 = n17596 & ~n18196;
  assign n18198 = ~n17596 & n18196;
  assign n18199 = ~n18197 & ~n18198;
  assign n18200 = ~n18194 & ~n18199;
  assign n18201 = ~n18193 & ~n18200;
  assign n18202 = po6  & ~n18201;
  assign n18203 = ~po6  & ~n18193;
  assign n18204 = ~n18200 & n18203;
  assign n18205 = ~n17599 & po2 ;
  assign n18206 = ~n17605 & n18205;
  assign n18207 = n17604 & ~n18206;
  assign n18208 = n17606 & n18205;
  assign n18209 = ~n18207 & ~n18208;
  assign n18210 = ~n18204 & n18209;
  assign n18211 = ~n18202 & ~n18210;
  assign n18212 = po7  & ~n18211;
  assign n18213 = ~po7  & n18211;
  assign n18214 = ~n17608 & ~n17610;
  assign n18215 = po2  & n18214;
  assign n18216 = n17615 & ~n18215;
  assign n18217 = ~n17615 & n18215;
  assign n18218 = ~n18216 & ~n18217;
  assign n18219 = ~n18213 & n18218;
  assign n18220 = ~n18212 & ~n18219;
  assign n18221 = po8  & ~n18220;
  assign n18222 = ~po8  & ~n18212;
  assign n18223 = ~n18219 & n18222;
  assign n18224 = ~n17618 & po2 ;
  assign n18225 = ~n17624 & n18224;
  assign n18226 = n17623 & ~n18225;
  assign n18227 = n17625 & n18224;
  assign n18228 = ~n18226 & ~n18227;
  assign n18229 = ~n18223 & n18228;
  assign n18230 = ~n18221 & ~n18229;
  assign n18231 = po9  & ~n18230;
  assign n18232 = ~po9  & n18230;
  assign n18233 = ~n17627 & ~n17629;
  assign n18234 = po2  & n18233;
  assign n18235 = n17634 & n18234;
  assign n18236 = ~n17634 & ~n18234;
  assign n18237 = ~n18235 & ~n18236;
  assign n18238 = ~n18232 & n18237;
  assign n18239 = ~n18231 & ~n18238;
  assign n18240 = po10  & ~n18239;
  assign n18241 = ~po10  & ~n18231;
  assign n18242 = ~n18238 & n18241;
  assign n18243 = ~n17637 & po2 ;
  assign n18244 = ~n17643 & n18243;
  assign n18245 = n17642 & ~n18244;
  assign n18246 = n17644 & n18243;
  assign n18247 = ~n18245 & ~n18246;
  assign n18248 = ~n18242 & n18247;
  assign n18249 = ~n18240 & ~n18248;
  assign n18250 = po11  & ~n18249;
  assign n18251 = ~po11  & n18249;
  assign n18252 = ~n17646 & ~n17648;
  assign n18253 = po2  & n18252;
  assign n18254 = ~n17653 & ~n18253;
  assign n18255 = n17653 & n18253;
  assign n18256 = ~n18254 & ~n18255;
  assign n18257 = ~n18251 & n18256;
  assign n18258 = ~n18250 & ~n18257;
  assign n18259 = po12  & ~n18258;
  assign n18260 = ~po12  & ~n18250;
  assign n18261 = ~n18257 & n18260;
  assign n18262 = ~n17656 & po2 ;
  assign n18263 = ~n17662 & n18262;
  assign n18264 = n17661 & ~n18263;
  assign n18265 = n17663 & n18262;
  assign n18266 = ~n18264 & ~n18265;
  assign n18267 = ~n18261 & n18266;
  assign n18268 = ~n18259 & ~n18267;
  assign n18269 = po13  & ~n18268;
  assign n18270 = ~n17665 & ~n17667;
  assign n18271 = po2  & n18270;
  assign n18272 = n17672 & ~n18271;
  assign n18273 = ~n17672 & n18271;
  assign n18274 = ~n18272 & ~n18273;
  assign n18275 = ~po13  & n18268;
  assign n18276 = ~n18274 & ~n18275;
  assign n18277 = ~n18269 & ~n18276;
  assign n18278 = po14  & ~n18277;
  assign n18279 = ~po14  & ~n18269;
  assign n18280 = ~n18276 & n18279;
  assign n18281 = ~n17675 & po2 ;
  assign n18282 = ~n17681 & n18281;
  assign n18283 = n17680 & ~n18282;
  assign n18284 = n17682 & n18281;
  assign n18285 = ~n18283 & ~n18284;
  assign n18286 = ~n18280 & n18285;
  assign n18287 = ~n18278 & ~n18286;
  assign n18288 = po15  & ~n18287;
  assign n18289 = ~po15  & n18287;
  assign n18290 = ~n17684 & po2 ;
  assign n18291 = ~n17691 & n18290;
  assign n18292 = n17689 & ~n18291;
  assign n18293 = n17692 & n18290;
  assign n18294 = ~n18292 & ~n18293;
  assign n18295 = ~n18289 & n18294;
  assign n18296 = ~n18288 & ~n18295;
  assign n18297 = po16  & ~n18296;
  assign n18298 = ~po16  & ~n18288;
  assign n18299 = ~n18295 & n18298;
  assign n18300 = ~n17694 & po2 ;
  assign n18301 = ~n17700 & n18300;
  assign n18302 = n17699 & ~n18301;
  assign n18303 = n17701 & n18300;
  assign n18304 = ~n18302 & ~n18303;
  assign n18305 = ~n18299 & n18304;
  assign n18306 = ~n18297 & ~n18305;
  assign n18307 = po17  & ~n18306;
  assign n18308 = ~n17703 & ~n17705;
  assign n18309 = po2  & n18308;
  assign n18310 = n17710 & ~n18309;
  assign n18311 = ~n17710 & n18309;
  assign n18312 = ~n18310 & ~n18311;
  assign n18313 = ~po17  & n18306;
  assign n18314 = ~n18312 & ~n18313;
  assign n18315 = ~n18307 & ~n18314;
  assign n18316 = po18  & ~n18315;
  assign n18317 = ~po18  & ~n18307;
  assign n18318 = ~n18314 & n18317;
  assign n18319 = ~n17713 & po2 ;
  assign n18320 = ~n17719 & n18319;
  assign n18321 = n17718 & ~n18320;
  assign n18322 = n17720 & n18319;
  assign n18323 = ~n18321 & ~n18322;
  assign n18324 = ~n18318 & n18323;
  assign n18325 = ~n18316 & ~n18324;
  assign n18326 = po19  & ~n18325;
  assign n18327 = ~po19  & n18325;
  assign n18328 = ~n17722 & po2 ;
  assign n18329 = ~n17729 & n18328;
  assign n18330 = n17727 & ~n18329;
  assign n18331 = n17730 & n18328;
  assign n18332 = ~n18330 & ~n18331;
  assign n18333 = ~n18327 & n18332;
  assign n18334 = ~n18326 & ~n18333;
  assign n18335 = po20  & ~n18334;
  assign n18336 = ~po20  & ~n18326;
  assign n18337 = ~n18333 & n18336;
  assign n18338 = ~n17732 & po2 ;
  assign n18339 = ~n17738 & n18338;
  assign n18340 = n17737 & ~n18339;
  assign n18341 = n17739 & n18338;
  assign n18342 = ~n18340 & ~n18341;
  assign n18343 = ~n18337 & n18342;
  assign n18344 = ~n18335 & ~n18343;
  assign n18345 = po21  & ~n18344;
  assign n18346 = ~n17741 & ~n17743;
  assign n18347 = po2  & n18346;
  assign n18348 = n17748 & ~n18347;
  assign n18349 = ~n17748 & n18347;
  assign n18350 = ~n18348 & ~n18349;
  assign n18351 = ~po21  & n18344;
  assign n18352 = ~n18350 & ~n18351;
  assign n18353 = ~n18345 & ~n18352;
  assign n18354 = po22  & ~n18353;
  assign n18355 = ~po22  & ~n18345;
  assign n18356 = ~n18352 & n18355;
  assign n18357 = ~n17751 & po2 ;
  assign n18358 = ~n17757 & n18357;
  assign n18359 = n17756 & ~n18358;
  assign n18360 = n17758 & n18357;
  assign n18361 = ~n18359 & ~n18360;
  assign n18362 = ~n18356 & n18361;
  assign n18363 = ~n18354 & ~n18362;
  assign n18364 = po23  & ~n18363;
  assign n18365 = ~po23  & n18363;
  assign n18366 = ~n17760 & po2 ;
  assign n18367 = ~n17767 & n18366;
  assign n18368 = n17765 & ~n18367;
  assign n18369 = n17768 & n18366;
  assign n18370 = ~n18368 & ~n18369;
  assign n18371 = ~n18365 & n18370;
  assign n18372 = ~n18364 & ~n18371;
  assign n18373 = po24  & ~n18372;
  assign n18374 = ~po24  & ~n18364;
  assign n18375 = ~n18371 & n18374;
  assign n18376 = ~n17770 & po2 ;
  assign n18377 = ~n17776 & n18376;
  assign n18378 = n17775 & ~n18377;
  assign n18379 = n17777 & n18376;
  assign n18380 = ~n18378 & ~n18379;
  assign n18381 = ~n18375 & n18380;
  assign n18382 = ~n18373 & ~n18381;
  assign n18383 = po25  & ~n18382;
  assign n18384 = ~n17779 & ~n17781;
  assign n18385 = po2  & n18384;
  assign n18386 = n17786 & ~n18385;
  assign n18387 = ~n17786 & n18385;
  assign n18388 = ~n18386 & ~n18387;
  assign n18389 = ~po25  & n18382;
  assign n18390 = ~n18388 & ~n18389;
  assign n18391 = ~n18383 & ~n18390;
  assign n18392 = po26  & ~n18391;
  assign n18393 = ~po26  & ~n18383;
  assign n18394 = ~n18390 & n18393;
  assign n18395 = ~n17789 & po2 ;
  assign n18396 = ~n17795 & n18395;
  assign n18397 = n17794 & ~n18396;
  assign n18398 = n17796 & n18395;
  assign n18399 = ~n18397 & ~n18398;
  assign n18400 = ~n18394 & n18399;
  assign n18401 = ~n18392 & ~n18400;
  assign n18402 = po27  & ~n18401;
  assign n18403 = ~po27  & n18401;
  assign n18404 = ~n17798 & po2 ;
  assign n18405 = ~n17805 & n18404;
  assign n18406 = n17803 & ~n18405;
  assign n18407 = n17806 & n18404;
  assign n18408 = ~n18406 & ~n18407;
  assign n18409 = ~n18403 & n18408;
  assign n18410 = ~n18402 & ~n18409;
  assign n18411 = po28  & ~n18410;
  assign n18412 = ~po28  & ~n18402;
  assign n18413 = ~n18409 & n18412;
  assign n18414 = ~n17808 & po2 ;
  assign n18415 = ~n17814 & n18414;
  assign n18416 = n17813 & ~n18415;
  assign n18417 = n17815 & n18414;
  assign n18418 = ~n18416 & ~n18417;
  assign n18419 = ~n18413 & n18418;
  assign n18420 = ~n18411 & ~n18419;
  assign n18421 = po29  & ~n18420;
  assign n18422 = ~n17817 & ~n17819;
  assign n18423 = po2  & n18422;
  assign n18424 = n17824 & ~n18423;
  assign n18425 = ~n17824 & n18423;
  assign n18426 = ~n18424 & ~n18425;
  assign n18427 = ~po29  & n18420;
  assign n18428 = ~n18426 & ~n18427;
  assign n18429 = ~n18421 & ~n18428;
  assign n18430 = po30  & ~n18429;
  assign n18431 = ~po30  & ~n18421;
  assign n18432 = ~n18428 & n18431;
  assign n18433 = ~n17827 & po2 ;
  assign n18434 = ~n17833 & n18433;
  assign n18435 = n17832 & ~n18434;
  assign n18436 = n17834 & n18433;
  assign n18437 = ~n18435 & ~n18436;
  assign n18438 = ~n18432 & n18437;
  assign n18439 = ~n18430 & ~n18438;
  assign n18440 = po31  & ~n18439;
  assign n18441 = ~po31  & n18439;
  assign n18442 = ~n17836 & po2 ;
  assign n18443 = ~n17843 & n18442;
  assign n18444 = n17841 & ~n18443;
  assign n18445 = n17844 & n18442;
  assign n18446 = ~n18444 & ~n18445;
  assign n18447 = ~n18441 & n18446;
  assign n18448 = ~n18440 & ~n18447;
  assign n18449 = po32  & ~n18448;
  assign n18450 = ~po32  & ~n18440;
  assign n18451 = ~n18447 & n18450;
  assign n18452 = ~n17846 & po2 ;
  assign n18453 = ~n17852 & n18452;
  assign n18454 = n17851 & ~n18453;
  assign n18455 = n17853 & n18452;
  assign n18456 = ~n18454 & ~n18455;
  assign n18457 = ~n18451 & n18456;
  assign n18458 = ~n18449 & ~n18457;
  assign n18459 = po33  & ~n18458;
  assign n18460 = ~n17855 & ~n17857;
  assign n18461 = po2  & n18460;
  assign n18462 = n17862 & ~n18461;
  assign n18463 = ~n17862 & n18461;
  assign n18464 = ~n18462 & ~n18463;
  assign n18465 = ~po33  & n18458;
  assign n18466 = ~n18464 & ~n18465;
  assign n18467 = ~n18459 & ~n18466;
  assign n18468 = po34  & ~n18467;
  assign n18469 = ~po34  & ~n18459;
  assign n18470 = ~n18466 & n18469;
  assign n18471 = ~n17865 & po2 ;
  assign n18472 = ~n17871 & n18471;
  assign n18473 = n17870 & ~n18472;
  assign n18474 = n17872 & n18471;
  assign n18475 = ~n18473 & ~n18474;
  assign n18476 = ~n18470 & n18475;
  assign n18477 = ~n18468 & ~n18476;
  assign n18478 = po35  & ~n18477;
  assign n18479 = ~po35  & n18477;
  assign n18480 = ~n17874 & po2 ;
  assign n18481 = ~n17881 & n18480;
  assign n18482 = n17879 & ~n18481;
  assign n18483 = n17882 & n18480;
  assign n18484 = ~n18482 & ~n18483;
  assign n18485 = ~n18479 & n18484;
  assign n18486 = ~n18478 & ~n18485;
  assign n18487 = po36  & ~n18486;
  assign n18488 = ~po36  & ~n18478;
  assign n18489 = ~n18485 & n18488;
  assign n18490 = ~n17884 & po2 ;
  assign n18491 = ~n17890 & n18490;
  assign n18492 = n17889 & ~n18491;
  assign n18493 = n17891 & n18490;
  assign n18494 = ~n18492 & ~n18493;
  assign n18495 = ~n18489 & n18494;
  assign n18496 = ~n18487 & ~n18495;
  assign n18497 = po37  & ~n18496;
  assign n18498 = ~n17893 & ~n17895;
  assign n18499 = po2  & n18498;
  assign n18500 = n17900 & ~n18499;
  assign n18501 = ~n17900 & n18499;
  assign n18502 = ~n18500 & ~n18501;
  assign n18503 = ~po37  & n18496;
  assign n18504 = ~n18502 & ~n18503;
  assign n18505 = ~n18497 & ~n18504;
  assign n18506 = po38  & ~n18505;
  assign n18507 = ~po38  & ~n18497;
  assign n18508 = ~n18504 & n18507;
  assign n18509 = ~n17903 & po2 ;
  assign n18510 = ~n17909 & n18509;
  assign n18511 = n17908 & ~n18510;
  assign n18512 = n17910 & n18509;
  assign n18513 = ~n18511 & ~n18512;
  assign n18514 = ~n18508 & n18513;
  assign n18515 = ~n18506 & ~n18514;
  assign n18516 = po39  & ~n18515;
  assign n18517 = ~po39  & n18515;
  assign n18518 = ~n17912 & po2 ;
  assign n18519 = ~n17919 & n18518;
  assign n18520 = n17917 & ~n18519;
  assign n18521 = n17920 & n18518;
  assign n18522 = ~n18520 & ~n18521;
  assign n18523 = ~n18517 & n18522;
  assign n18524 = ~n18516 & ~n18523;
  assign n18525 = po40  & ~n18524;
  assign n18526 = ~po40  & ~n18516;
  assign n18527 = ~n18523 & n18526;
  assign n18528 = ~n17922 & po2 ;
  assign n18529 = ~n17928 & n18528;
  assign n18530 = n17927 & ~n18529;
  assign n18531 = n17929 & n18528;
  assign n18532 = ~n18530 & ~n18531;
  assign n18533 = ~n18527 & n18532;
  assign n18534 = ~n18525 & ~n18533;
  assign n18535 = po41  & ~n18534;
  assign n18536 = ~n17931 & ~n17933;
  assign n18537 = po2  & n18536;
  assign n18538 = n17938 & ~n18537;
  assign n18539 = ~n17938 & n18537;
  assign n18540 = ~n18538 & ~n18539;
  assign n18541 = ~po41  & n18534;
  assign n18542 = ~n18540 & ~n18541;
  assign n18543 = ~n18535 & ~n18542;
  assign n18544 = po42  & ~n18543;
  assign n18545 = ~po42  & ~n18535;
  assign n18546 = ~n18542 & n18545;
  assign n18547 = ~n17941 & po2 ;
  assign n18548 = ~n17947 & n18547;
  assign n18549 = n17946 & ~n18548;
  assign n18550 = n17948 & n18547;
  assign n18551 = ~n18549 & ~n18550;
  assign n18552 = ~n18546 & n18551;
  assign n18553 = ~n18544 & ~n18552;
  assign n18554 = po43  & ~n18553;
  assign n18555 = ~po43  & n18553;
  assign n18556 = ~n17950 & po2 ;
  assign n18557 = ~n17957 & n18556;
  assign n18558 = n17955 & ~n18557;
  assign n18559 = n17958 & n18556;
  assign n18560 = ~n18558 & ~n18559;
  assign n18561 = ~n18555 & n18560;
  assign n18562 = ~n18554 & ~n18561;
  assign n18563 = po44  & ~n18562;
  assign n18564 = ~po44  & ~n18554;
  assign n18565 = ~n18561 & n18564;
  assign n18566 = ~n17960 & po2 ;
  assign n18567 = ~n17966 & n18566;
  assign n18568 = n17965 & ~n18567;
  assign n18569 = n17967 & n18566;
  assign n18570 = ~n18568 & ~n18569;
  assign n18571 = ~n18565 & n18570;
  assign n18572 = ~n18563 & ~n18571;
  assign n18573 = po45  & ~n18572;
  assign n18574 = ~n17969 & ~n17971;
  assign n18575 = po2  & n18574;
  assign n18576 = n17976 & ~n18575;
  assign n18577 = ~n17976 & n18575;
  assign n18578 = ~n18576 & ~n18577;
  assign n18579 = ~po45  & n18572;
  assign n18580 = ~n18578 & ~n18579;
  assign n18581 = ~n18573 & ~n18580;
  assign n18582 = po46  & ~n18581;
  assign n18583 = ~po46  & ~n18573;
  assign n18584 = ~n18580 & n18583;
  assign n18585 = ~n17979 & po2 ;
  assign n18586 = ~n17985 & n18585;
  assign n18587 = n17984 & ~n18586;
  assign n18588 = n17986 & n18585;
  assign n18589 = ~n18587 & ~n18588;
  assign n18590 = ~n18584 & n18589;
  assign n18591 = ~n18582 & ~n18590;
  assign n18592 = po47  & ~n18591;
  assign n18593 = ~po47  & n18591;
  assign n18594 = ~n17988 & po2 ;
  assign n18595 = ~n17995 & n18594;
  assign n18596 = n17993 & ~n18595;
  assign n18597 = n17996 & n18594;
  assign n18598 = ~n18596 & ~n18597;
  assign n18599 = ~n18593 & n18598;
  assign n18600 = ~n18592 & ~n18599;
  assign n18601 = po48  & ~n18600;
  assign n18602 = ~po48  & ~n18592;
  assign n18603 = ~n18599 & n18602;
  assign n18604 = ~n17998 & po2 ;
  assign n18605 = ~n18004 & n18604;
  assign n18606 = n18003 & ~n18605;
  assign n18607 = n18005 & n18604;
  assign n18608 = ~n18606 & ~n18607;
  assign n18609 = ~n18603 & n18608;
  assign n18610 = ~n18601 & ~n18609;
  assign n18611 = po49  & ~n18610;
  assign n18612 = ~n18007 & ~n18009;
  assign n18613 = po2  & n18612;
  assign n18614 = n18014 & ~n18613;
  assign n18615 = ~n18014 & n18613;
  assign n18616 = ~n18614 & ~n18615;
  assign n18617 = ~po49  & n18610;
  assign n18618 = ~n18616 & ~n18617;
  assign n18619 = ~n18611 & ~n18618;
  assign n18620 = po50  & ~n18619;
  assign n18621 = ~po50  & ~n18611;
  assign n18622 = ~n18618 & n18621;
  assign n18623 = ~n18017 & po2 ;
  assign n18624 = ~n18023 & n18623;
  assign n18625 = n18022 & ~n18624;
  assign n18626 = n18024 & n18623;
  assign n18627 = ~n18625 & ~n18626;
  assign n18628 = ~n18622 & n18627;
  assign n18629 = ~n18620 & ~n18628;
  assign n18630 = po51  & ~n18629;
  assign n18631 = ~po51  & n18629;
  assign n18632 = ~n18026 & po2 ;
  assign n18633 = ~n18033 & n18632;
  assign n18634 = n18031 & ~n18633;
  assign n18635 = n18034 & n18632;
  assign n18636 = ~n18634 & ~n18635;
  assign n18637 = ~n18631 & n18636;
  assign n18638 = ~n18630 & ~n18637;
  assign n18639 = po52  & ~n18638;
  assign n18640 = ~po52  & ~n18630;
  assign n18641 = ~n18637 & n18640;
  assign n18642 = ~n18036 & po2 ;
  assign n18643 = ~n18042 & n18642;
  assign n18644 = n18041 & ~n18643;
  assign n18645 = n18043 & n18642;
  assign n18646 = ~n18644 & ~n18645;
  assign n18647 = ~n18641 & n18646;
  assign n18648 = ~n18639 & ~n18647;
  assign n18649 = po53  & ~n18648;
  assign n18650 = ~n18045 & ~n18047;
  assign n18651 = po2  & n18650;
  assign n18652 = n18052 & ~n18651;
  assign n18653 = ~n18052 & n18651;
  assign n18654 = ~n18652 & ~n18653;
  assign n18655 = ~po53  & n18648;
  assign n18656 = ~n18654 & ~n18655;
  assign n18657 = ~n18649 & ~n18656;
  assign n18658 = po54  & ~n18657;
  assign n18659 = ~po54  & ~n18649;
  assign n18660 = ~n18656 & n18659;
  assign n18661 = ~n18055 & po2 ;
  assign n18662 = ~n18061 & n18661;
  assign n18663 = n18060 & ~n18662;
  assign n18664 = n18062 & n18661;
  assign n18665 = ~n18663 & ~n18664;
  assign n18666 = ~n18660 & n18665;
  assign n18667 = ~n18658 & ~n18666;
  assign n18668 = po55  & ~n18667;
  assign n18669 = ~po55  & n18667;
  assign n18670 = ~n18064 & po2 ;
  assign n18671 = ~n18071 & n18670;
  assign n18672 = n18069 & ~n18671;
  assign n18673 = n18072 & n18670;
  assign n18674 = ~n18672 & ~n18673;
  assign n18675 = ~n18669 & n18674;
  assign n18676 = ~n18668 & ~n18675;
  assign n18677 = po56  & ~n18676;
  assign n18678 = ~po56  & ~n18668;
  assign n18679 = ~n18675 & n18678;
  assign n18680 = ~n18074 & po2 ;
  assign n18681 = ~n18080 & n18680;
  assign n18682 = n18079 & ~n18681;
  assign n18683 = n18081 & n18680;
  assign n18684 = ~n18682 & ~n18683;
  assign n18685 = ~n18679 & n18684;
  assign n18686 = ~n18677 & ~n18685;
  assign n18687 = po57  & ~n18686;
  assign n18688 = ~n18083 & ~n18085;
  assign n18689 = po2  & n18688;
  assign n18690 = n18090 & ~n18689;
  assign n18691 = ~n18090 & n18689;
  assign n18692 = ~n18690 & ~n18691;
  assign n18693 = ~po57  & n18686;
  assign n18694 = ~n18692 & ~n18693;
  assign n18695 = ~n18687 & ~n18694;
  assign n18696 = po58  & ~n18695;
  assign n18697 = ~po58  & ~n18687;
  assign n18698 = ~n18694 & n18697;
  assign n18699 = ~n18093 & po2 ;
  assign n18700 = ~n18099 & n18699;
  assign n18701 = n18098 & ~n18700;
  assign n18702 = n18100 & n18699;
  assign n18703 = ~n18701 & ~n18702;
  assign n18704 = ~n18698 & n18703;
  assign n18705 = ~n18696 & ~n18704;
  assign n18706 = po59  & ~n18705;
  assign n18707 = ~po59  & n18705;
  assign n18708 = ~n18102 & po2 ;
  assign n18709 = ~n18109 & n18708;
  assign n18710 = n18107 & ~n18709;
  assign n18711 = n18110 & n18708;
  assign n18712 = ~n18710 & ~n18711;
  assign n18713 = ~n18707 & n18712;
  assign n18714 = ~n18706 & ~n18713;
  assign n18715 = po60  & ~n18714;
  assign n18716 = ~n18112 & ~n18119;
  assign n18717 = po2  & n18716;
  assign n18718 = n18117 & ~n18717;
  assign n18719 = ~n18117 & n18717;
  assign n18720 = ~n18718 & ~n18719;
  assign n18721 = ~po60  & ~n18706;
  assign n18722 = ~n18713 & n18721;
  assign n18723 = ~n18720 & ~n18722;
  assign n18724 = ~n18715 & ~n18723;
  assign n18725 = ~po61  & n18724;
  assign n18726 = ~n18170 & ~n18725;
  assign n18727 = po61  & ~n18724;
  assign n18728 = ~po62  & ~n18727;
  assign n18729 = ~n18726 & n18728;
  assign n18730 = ~n18726 & ~n18727;
  assign n18731 = po62  & ~n18730;
  assign n18732 = n18165 & ~n18729;
  assign n18733 = ~n18731 & ~n18732;
  assign n18734 = ~n18135 & ~n18137;
  assign n18735 = po2  & n18734;
  assign n18736 = n18142 & ~n18735;
  assign n18737 = ~n18142 & n18735;
  assign n18738 = ~n18736 & ~n18737;
  assign n18739 = n18144 & po2 ;
  assign n18740 = ~n18149 & ~n18739;
  assign n18741 = ~n18157 & ~n18740;
  assign n18742 = po2  & ~n18741;
  assign n18743 = ~n18738 & ~n18742;
  assign n18744 = ~n18733 & n18743;
  assign n18745 = ~po63  & ~n18744;
  assign n18746 = n18733 & n18738;
  assign n18747 = po63  & n18741;
  assign n18748 = ~n18746 & ~n18747;
  assign po1  = n18745 | ~n18748;
  assign n18750 = ~n18729 & ~n18731;
  assign n18751 = po1  & n18750;
  assign n18752 = n18165 & ~n18751;
  assign n18753 = ~n18165 & n18751;
  assign n18754 = ~n18752 & ~n18753;
  assign n18755 = po63  & ~n18754;
  assign n18756 = ~n18725 & ~n18727;
  assign n18757 = po1  & n18756;
  assign n18758 = n18170 & n18757;
  assign n18759 = ~n18170 & ~n18757;
  assign n18760 = ~n18758 & ~n18759;
  assign n18761 = po62  & ~n18760;
  assign n18762 = ~po62  & n18760;
  assign n18763 = ~n18715 & po1 ;
  assign n18764 = ~n18722 & n18763;
  assign n18765 = n18720 & ~n18764;
  assign n18766 = n18723 & n18763;
  assign n18767 = ~n18765 & ~n18766;
  assign n18768 = ~po61  & ~n18767;
  assign n18769 = po61  & n18767;
  assign n18770 = ~n18706 & ~n18707;
  assign n18771 = po1  & n18770;
  assign n18772 = n18712 & ~n18771;
  assign n18773 = ~n18712 & n18771;
  assign n18774 = ~n18772 & ~n18773;
  assign n18775 = po60  & ~n18774;
  assign n18776 = ~po60  & n18774;
  assign n18777 = ~n18696 & ~n18698;
  assign n18778 = po1  & n18777;
  assign n18779 = n18703 & ~n18778;
  assign n18780 = ~n18703 & n18778;
  assign n18781 = ~n18779 & ~n18780;
  assign n18782 = ~po59  & n18781;
  assign n18783 = po59  & ~n18781;
  assign n18784 = ~n18687 & po1 ;
  assign n18785 = ~n18693 & n18784;
  assign n18786 = n18692 & ~n18785;
  assign n18787 = n18694 & n18784;
  assign n18788 = ~n18786 & ~n18787;
  assign n18789 = po58  & n18788;
  assign n18790 = ~po58  & ~n18788;
  assign n18791 = ~n18677 & ~n18679;
  assign n18792 = po1  & n18791;
  assign n18793 = n18684 & ~n18792;
  assign n18794 = ~n18684 & n18792;
  assign n18795 = ~n18793 & ~n18794;
  assign n18796 = ~po57  & n18795;
  assign n18797 = po57  & ~n18795;
  assign n18798 = ~n18668 & ~n18669;
  assign n18799 = po1  & n18798;
  assign n18800 = n18674 & ~n18799;
  assign n18801 = ~n18674 & n18799;
  assign n18802 = ~n18800 & ~n18801;
  assign n18803 = po56  & ~n18802;
  assign n18804 = ~po56  & n18802;
  assign n18805 = ~n18658 & ~n18660;
  assign n18806 = po1  & n18805;
  assign n18807 = n18665 & ~n18806;
  assign n18808 = ~n18665 & n18806;
  assign n18809 = ~n18807 & ~n18808;
  assign n18810 = ~po55  & n18809;
  assign n18811 = po55  & ~n18809;
  assign n18812 = ~n18649 & po1 ;
  assign n18813 = ~n18655 & n18812;
  assign n18814 = n18654 & ~n18813;
  assign n18815 = n18656 & n18812;
  assign n18816 = ~n18814 & ~n18815;
  assign n18817 = po54  & n18816;
  assign n18818 = ~po54  & ~n18816;
  assign n18819 = ~n18639 & ~n18641;
  assign n18820 = po1  & n18819;
  assign n18821 = n18646 & ~n18820;
  assign n18822 = ~n18646 & n18820;
  assign n18823 = ~n18821 & ~n18822;
  assign n18824 = ~po53  & n18823;
  assign n18825 = po53  & ~n18823;
  assign n18826 = ~n18630 & ~n18631;
  assign n18827 = po1  & n18826;
  assign n18828 = n18636 & ~n18827;
  assign n18829 = ~n18636 & n18827;
  assign n18830 = ~n18828 & ~n18829;
  assign n18831 = po52  & ~n18830;
  assign n18832 = ~po52  & n18830;
  assign n18833 = ~n18620 & ~n18622;
  assign n18834 = po1  & n18833;
  assign n18835 = n18627 & ~n18834;
  assign n18836 = ~n18627 & n18834;
  assign n18837 = ~n18835 & ~n18836;
  assign n18838 = ~po51  & n18837;
  assign n18839 = po51  & ~n18837;
  assign n18840 = ~n18611 & po1 ;
  assign n18841 = ~n18617 & n18840;
  assign n18842 = n18616 & ~n18841;
  assign n18843 = n18618 & n18840;
  assign n18844 = ~n18842 & ~n18843;
  assign n18845 = po50  & n18844;
  assign n18846 = ~po50  & ~n18844;
  assign n18847 = ~n18601 & ~n18603;
  assign n18848 = po1  & n18847;
  assign n18849 = n18608 & ~n18848;
  assign n18850 = ~n18608 & n18848;
  assign n18851 = ~n18849 & ~n18850;
  assign n18852 = ~po49  & n18851;
  assign n18853 = po49  & ~n18851;
  assign n18854 = ~n18592 & ~n18593;
  assign n18855 = po1  & n18854;
  assign n18856 = n18598 & ~n18855;
  assign n18857 = ~n18598 & n18855;
  assign n18858 = ~n18856 & ~n18857;
  assign n18859 = po48  & ~n18858;
  assign n18860 = ~po48  & n18858;
  assign n18861 = ~n18582 & ~n18584;
  assign n18862 = po1  & n18861;
  assign n18863 = n18589 & ~n18862;
  assign n18864 = ~n18589 & n18862;
  assign n18865 = ~n18863 & ~n18864;
  assign n18866 = ~po47  & n18865;
  assign n18867 = po47  & ~n18865;
  assign n18868 = ~n18573 & po1 ;
  assign n18869 = ~n18579 & n18868;
  assign n18870 = n18578 & ~n18869;
  assign n18871 = n18580 & n18868;
  assign n18872 = ~n18870 & ~n18871;
  assign n18873 = po46  & n18872;
  assign n18874 = ~po46  & ~n18872;
  assign n18875 = ~n18563 & ~n18565;
  assign n18876 = po1  & n18875;
  assign n18877 = n18570 & ~n18876;
  assign n18878 = ~n18570 & n18876;
  assign n18879 = ~n18877 & ~n18878;
  assign n18880 = ~po45  & n18879;
  assign n18881 = po45  & ~n18879;
  assign n18882 = ~n18554 & ~n18555;
  assign n18883 = po1  & n18882;
  assign n18884 = n18560 & ~n18883;
  assign n18885 = ~n18560 & n18883;
  assign n18886 = ~n18884 & ~n18885;
  assign n18887 = po44  & ~n18886;
  assign n18888 = ~po44  & n18886;
  assign n18889 = ~n18544 & ~n18546;
  assign n18890 = po1  & n18889;
  assign n18891 = n18551 & ~n18890;
  assign n18892 = ~n18551 & n18890;
  assign n18893 = ~n18891 & ~n18892;
  assign n18894 = ~po43  & n18893;
  assign n18895 = po43  & ~n18893;
  assign n18896 = ~n18535 & po1 ;
  assign n18897 = ~n18541 & n18896;
  assign n18898 = n18540 & ~n18897;
  assign n18899 = n18542 & n18896;
  assign n18900 = ~n18898 & ~n18899;
  assign n18901 = po42  & n18900;
  assign n18902 = ~po42  & ~n18900;
  assign n18903 = ~n18525 & ~n18527;
  assign n18904 = po1  & n18903;
  assign n18905 = n18532 & ~n18904;
  assign n18906 = ~n18532 & n18904;
  assign n18907 = ~n18905 & ~n18906;
  assign n18908 = ~po41  & n18907;
  assign n18909 = po41  & ~n18907;
  assign n18910 = ~n18516 & ~n18517;
  assign n18911 = po1  & n18910;
  assign n18912 = n18522 & ~n18911;
  assign n18913 = ~n18522 & n18911;
  assign n18914 = ~n18912 & ~n18913;
  assign n18915 = po40  & ~n18914;
  assign n18916 = ~po40  & n18914;
  assign n18917 = ~n18506 & ~n18508;
  assign n18918 = po1  & n18917;
  assign n18919 = n18513 & ~n18918;
  assign n18920 = ~n18513 & n18918;
  assign n18921 = ~n18919 & ~n18920;
  assign n18922 = ~po39  & n18921;
  assign n18923 = po39  & ~n18921;
  assign n18924 = ~n18497 & po1 ;
  assign n18925 = ~n18503 & n18924;
  assign n18926 = n18502 & ~n18925;
  assign n18927 = n18504 & n18924;
  assign n18928 = ~n18926 & ~n18927;
  assign n18929 = po38  & n18928;
  assign n18930 = ~po38  & ~n18928;
  assign n18931 = ~n18487 & ~n18489;
  assign n18932 = po1  & n18931;
  assign n18933 = n18494 & ~n18932;
  assign n18934 = ~n18494 & n18932;
  assign n18935 = ~n18933 & ~n18934;
  assign n18936 = ~po37  & n18935;
  assign n18937 = po37  & ~n18935;
  assign n18938 = ~n18478 & ~n18479;
  assign n18939 = po1  & n18938;
  assign n18940 = n18484 & ~n18939;
  assign n18941 = ~n18484 & n18939;
  assign n18942 = ~n18940 & ~n18941;
  assign n18943 = po36  & ~n18942;
  assign n18944 = ~po36  & n18942;
  assign n18945 = ~n18468 & ~n18470;
  assign n18946 = po1  & n18945;
  assign n18947 = n18475 & ~n18946;
  assign n18948 = ~n18475 & n18946;
  assign n18949 = ~n18947 & ~n18948;
  assign n18950 = ~po35  & n18949;
  assign n18951 = po35  & ~n18949;
  assign n18952 = ~n18459 & po1 ;
  assign n18953 = ~n18465 & n18952;
  assign n18954 = n18464 & ~n18953;
  assign n18955 = n18466 & n18952;
  assign n18956 = ~n18954 & ~n18955;
  assign n18957 = po34  & n18956;
  assign n18958 = ~po34  & ~n18956;
  assign n18959 = ~n18449 & ~n18451;
  assign n18960 = po1  & n18959;
  assign n18961 = n18456 & ~n18960;
  assign n18962 = ~n18456 & n18960;
  assign n18963 = ~n18961 & ~n18962;
  assign n18964 = ~po33  & n18963;
  assign n18965 = po33  & ~n18963;
  assign n18966 = ~n18440 & ~n18441;
  assign n18967 = po1  & n18966;
  assign n18968 = n18446 & ~n18967;
  assign n18969 = ~n18446 & n18967;
  assign n18970 = ~n18968 & ~n18969;
  assign n18971 = po32  & ~n18970;
  assign n18972 = ~po32  & n18970;
  assign n18973 = ~n18430 & ~n18432;
  assign n18974 = po1  & n18973;
  assign n18975 = n18437 & ~n18974;
  assign n18976 = ~n18437 & n18974;
  assign n18977 = ~n18975 & ~n18976;
  assign n18978 = ~po31  & n18977;
  assign n18979 = po31  & ~n18977;
  assign n18980 = ~n18421 & po1 ;
  assign n18981 = ~n18427 & n18980;
  assign n18982 = n18426 & ~n18981;
  assign n18983 = n18428 & n18980;
  assign n18984 = ~n18982 & ~n18983;
  assign n18985 = po30  & n18984;
  assign n18986 = ~po30  & ~n18984;
  assign n18987 = ~n18411 & ~n18413;
  assign n18988 = po1  & n18987;
  assign n18989 = n18418 & ~n18988;
  assign n18990 = ~n18418 & n18988;
  assign n18991 = ~n18989 & ~n18990;
  assign n18992 = ~po29  & n18991;
  assign n18993 = po29  & ~n18991;
  assign n18994 = ~n18402 & ~n18403;
  assign n18995 = po1  & n18994;
  assign n18996 = n18408 & ~n18995;
  assign n18997 = ~n18408 & n18995;
  assign n18998 = ~n18996 & ~n18997;
  assign n18999 = po28  & ~n18998;
  assign n19000 = ~po28  & n18998;
  assign n19001 = ~n18392 & ~n18394;
  assign n19002 = po1  & n19001;
  assign n19003 = n18399 & ~n19002;
  assign n19004 = ~n18399 & n19002;
  assign n19005 = ~n19003 & ~n19004;
  assign n19006 = ~po27  & n19005;
  assign n19007 = po27  & ~n19005;
  assign n19008 = ~n18383 & po1 ;
  assign n19009 = ~n18389 & n19008;
  assign n19010 = n18388 & ~n19009;
  assign n19011 = n18390 & n19008;
  assign n19012 = ~n19010 & ~n19011;
  assign n19013 = po26  & n19012;
  assign n19014 = ~po26  & ~n19012;
  assign n19015 = ~n18373 & ~n18375;
  assign n19016 = po1  & n19015;
  assign n19017 = n18380 & ~n19016;
  assign n19018 = ~n18380 & n19016;
  assign n19019 = ~n19017 & ~n19018;
  assign n19020 = ~po25  & n19019;
  assign n19021 = po25  & ~n19019;
  assign n19022 = ~n18364 & ~n18365;
  assign n19023 = po1  & n19022;
  assign n19024 = n18370 & ~n19023;
  assign n19025 = ~n18370 & n19023;
  assign n19026 = ~n19024 & ~n19025;
  assign n19027 = po24  & ~n19026;
  assign n19028 = ~po24  & n19026;
  assign n19029 = ~n18354 & ~n18356;
  assign n19030 = po1  & n19029;
  assign n19031 = n18361 & ~n19030;
  assign n19032 = ~n18361 & n19030;
  assign n19033 = ~n19031 & ~n19032;
  assign n19034 = ~po23  & n19033;
  assign n19035 = po23  & ~n19033;
  assign n19036 = ~n18345 & po1 ;
  assign n19037 = ~n18351 & n19036;
  assign n19038 = n18350 & ~n19037;
  assign n19039 = n18352 & n19036;
  assign n19040 = ~n19038 & ~n19039;
  assign n19041 = po22  & n19040;
  assign n19042 = ~po22  & ~n19040;
  assign n19043 = ~n18335 & ~n18337;
  assign n19044 = po1  & n19043;
  assign n19045 = n18342 & ~n19044;
  assign n19046 = ~n18342 & n19044;
  assign n19047 = ~n19045 & ~n19046;
  assign n19048 = ~po21  & n19047;
  assign n19049 = po21  & ~n19047;
  assign n19050 = ~n18326 & ~n18327;
  assign n19051 = po1  & n19050;
  assign n19052 = n18332 & ~n19051;
  assign n19053 = ~n18332 & n19051;
  assign n19054 = ~n19052 & ~n19053;
  assign n19055 = po20  & ~n19054;
  assign n19056 = ~po20  & n19054;
  assign n19057 = ~n18316 & ~n18318;
  assign n19058 = po1  & n19057;
  assign n19059 = n18323 & ~n19058;
  assign n19060 = ~n18323 & n19058;
  assign n19061 = ~n19059 & ~n19060;
  assign n19062 = ~po19  & n19061;
  assign n19063 = po19  & ~n19061;
  assign n19064 = ~n18307 & po1 ;
  assign n19065 = ~n18313 & n19064;
  assign n19066 = n18312 & ~n19065;
  assign n19067 = n18314 & n19064;
  assign n19068 = ~n19066 & ~n19067;
  assign n19069 = po18  & n19068;
  assign n19070 = ~po18  & ~n19068;
  assign n19071 = ~n18297 & ~n18299;
  assign n19072 = po1  & n19071;
  assign n19073 = n18304 & ~n19072;
  assign n19074 = ~n18304 & n19072;
  assign n19075 = ~n19073 & ~n19074;
  assign n19076 = ~po17  & n19075;
  assign n19077 = po17  & ~n19075;
  assign n19078 = ~n18288 & ~n18289;
  assign n19079 = po1  & n19078;
  assign n19080 = n18294 & ~n19079;
  assign n19081 = ~n18294 & n19079;
  assign n19082 = ~n19080 & ~n19081;
  assign n19083 = po16  & ~n19082;
  assign n19084 = ~po16  & n19082;
  assign n19085 = ~n18278 & ~n18280;
  assign n19086 = po1  & n19085;
  assign n19087 = n18285 & ~n19086;
  assign n19088 = ~n18285 & n19086;
  assign n19089 = ~n19087 & ~n19088;
  assign n19090 = ~po15  & n19089;
  assign n19091 = po15  & ~n19089;
  assign n19092 = ~n18269 & po1 ;
  assign n19093 = ~n18275 & n19092;
  assign n19094 = n18274 & ~n19093;
  assign n19095 = n18276 & n19092;
  assign n19096 = ~n19094 & ~n19095;
  assign n19097 = po14  & n19096;
  assign n19098 = ~po14  & ~n19096;
  assign n19099 = ~n18259 & ~n18261;
  assign n19100 = po1  & n19099;
  assign n19101 = n18266 & ~n19100;
  assign n19102 = ~n18266 & n19100;
  assign n19103 = ~n19101 & ~n19102;
  assign n19104 = ~po13  & n19103;
  assign n19105 = po13  & ~n19103;
  assign n19106 = ~n18250 & ~n18251;
  assign n19107 = po1  & n19106;
  assign n19108 = n18256 & ~n19107;
  assign n19109 = ~n18256 & n19107;
  assign n19110 = ~n19108 & ~n19109;
  assign n19111 = po12  & ~n19110;
  assign n19112 = ~po12  & n19110;
  assign n19113 = ~n18240 & ~n18242;
  assign n19114 = po1  & n19113;
  assign n19115 = n18247 & ~n19114;
  assign n19116 = ~n18247 & n19114;
  assign n19117 = ~n19115 & ~n19116;
  assign n19118 = ~po11  & n19117;
  assign n19119 = po11  & ~n19117;
  assign n19120 = ~n18231 & ~n18232;
  assign n19121 = po1  & n19120;
  assign n19122 = ~n18237 & ~n19121;
  assign n19123 = n18237 & n19121;
  assign n19124 = ~n19122 & ~n19123;
  assign n19125 = po10  & n19124;
  assign n19126 = ~po10  & ~n19124;
  assign n19127 = ~n18221 & ~n18223;
  assign n19128 = po1  & n19127;
  assign n19129 = n18228 & ~n19128;
  assign n19130 = ~n18228 & n19128;
  assign n19131 = ~n19129 & ~n19130;
  assign n19132 = ~po9  & n19131;
  assign n19133 = po9  & ~n19131;
  assign n19134 = ~n18212 & ~n18213;
  assign n19135 = po1  & n19134;
  assign n19136 = n18218 & n19135;
  assign n19137 = ~n18218 & ~n19135;
  assign n19138 = ~n19136 & ~n19137;
  assign n19139 = po8  & n19138;
  assign n19140 = ~po8  & ~n19138;
  assign n19141 = ~n18202 & ~n18204;
  assign n19142 = po1  & n19141;
  assign n19143 = n18209 & ~n19142;
  assign n19144 = ~n18209 & n19142;
  assign n19145 = ~n19143 & ~n19144;
  assign n19146 = ~po7  & n19145;
  assign n19147 = po7  & ~n19145;
  assign n19148 = ~n18193 & ~n18194;
  assign n19149 = po1  & n19148;
  assign n19150 = n18199 & ~n19149;
  assign n19151 = ~n18199 & n19149;
  assign n19152 = ~n19150 & ~n19151;
  assign n19153 = po6  & n19152;
  assign n19154 = ~n18183 & ~n18185;
  assign n19155 = po1  & n19154;
  assign n19156 = ~n18190 & ~n19155;
  assign n19157 = n18190 & n19155;
  assign n19158 = ~n19156 & ~n19157;
  assign n19159 = ~po5  & n19158;
  assign n19160 = ~po6  & ~n19152;
  assign n19161 = po5  & ~n19158;
  assign n19162 = ~n18175 & ~n18180;
  assign n19163 = po1  & n19162;
  assign n19164 = n18179 & ~n19163;
  assign n19165 = ~n18179 & n19163;
  assign n19166 = ~n19164 & ~n19165;
  assign n19167 = po4  & ~n19166;
  assign n19168 = po2  & ~po1 ;
  assign n19169 = ~pi2  & po1 ;
  assign n19170 = ~pi3  & n19169;
  assign n19171 = ~n19168 & ~n19170;
  assign n19172 = pi4  & ~n19171;
  assign n19173 = ~pi4  & n19171;
  assign n19174 = ~pi0  & ~pi1 ;
  assign n19175 = ~pi2  & ~n19174;
  assign n19176 = pi2  & ~po1 ;
  assign n19177 = ~n19175 & ~n19176;
  assign n19178 = ~po2  & ~n19177;
  assign n19179 = po2  & n19177;
  assign n19180 = pi3  & ~n19169;
  assign n19181 = ~n19170 & ~n19180;
  assign n19182 = ~n19179 & ~n19181;
  assign n19183 = ~n19178 & ~n19182;
  assign n19184 = po3  & n19183;
  assign n19185 = ~n19172 & ~n19173;
  assign n19186 = ~n19184 & n19185;
  assign n19187 = ~po4  & n19166;
  assign n19188 = ~po3  & ~n19183;
  assign n19189 = ~n19187 & ~n19188;
  assign n19190 = ~n19186 & n19189;
  assign n19191 = ~n19161 & ~n19167;
  assign n19192 = ~n19190 & n19191;
  assign n19193 = ~n19159 & ~n19160;
  assign n19194 = ~n19192 & n19193;
  assign n19195 = ~n19147 & ~n19153;
  assign n19196 = ~n19194 & n19195;
  assign n19197 = ~n19140 & ~n19146;
  assign n19198 = ~n19196 & n19197;
  assign n19199 = ~n19133 & ~n19139;
  assign n19200 = ~n19198 & n19199;
  assign n19201 = ~n19126 & ~n19132;
  assign n19202 = ~n19200 & n19201;
  assign n19203 = ~n19119 & ~n19125;
  assign n19204 = ~n19202 & n19203;
  assign n19205 = ~n19112 & ~n19118;
  assign n19206 = ~n19204 & n19205;
  assign n19207 = ~n19105 & ~n19111;
  assign n19208 = ~n19206 & n19207;
  assign n19209 = ~n19098 & ~n19104;
  assign n19210 = ~n19208 & n19209;
  assign n19211 = ~n19091 & ~n19097;
  assign n19212 = ~n19210 & n19211;
  assign n19213 = ~n19084 & ~n19090;
  assign n19214 = ~n19212 & n19213;
  assign n19215 = ~n19077 & ~n19083;
  assign n19216 = ~n19214 & n19215;
  assign n19217 = ~n19070 & ~n19076;
  assign n19218 = ~n19216 & n19217;
  assign n19219 = ~n19063 & ~n19069;
  assign n19220 = ~n19218 & n19219;
  assign n19221 = ~n19056 & ~n19062;
  assign n19222 = ~n19220 & n19221;
  assign n19223 = ~n19049 & ~n19055;
  assign n19224 = ~n19222 & n19223;
  assign n19225 = ~n19042 & ~n19048;
  assign n19226 = ~n19224 & n19225;
  assign n19227 = ~n19035 & ~n19041;
  assign n19228 = ~n19226 & n19227;
  assign n19229 = ~n19028 & ~n19034;
  assign n19230 = ~n19228 & n19229;
  assign n19231 = ~n19021 & ~n19027;
  assign n19232 = ~n19230 & n19231;
  assign n19233 = ~n19014 & ~n19020;
  assign n19234 = ~n19232 & n19233;
  assign n19235 = ~n19007 & ~n19013;
  assign n19236 = ~n19234 & n19235;
  assign n19237 = ~n19000 & ~n19006;
  assign n19238 = ~n19236 & n19237;
  assign n19239 = ~n18993 & ~n18999;
  assign n19240 = ~n19238 & n19239;
  assign n19241 = ~n18986 & ~n18992;
  assign n19242 = ~n19240 & n19241;
  assign n19243 = ~n18979 & ~n18985;
  assign n19244 = ~n19242 & n19243;
  assign n19245 = ~n18972 & ~n18978;
  assign n19246 = ~n19244 & n19245;
  assign n19247 = ~n18965 & ~n18971;
  assign n19248 = ~n19246 & n19247;
  assign n19249 = ~n18958 & ~n18964;
  assign n19250 = ~n19248 & n19249;
  assign n19251 = ~n18951 & ~n18957;
  assign n19252 = ~n19250 & n19251;
  assign n19253 = ~n18944 & ~n18950;
  assign n19254 = ~n19252 & n19253;
  assign n19255 = ~n18937 & ~n18943;
  assign n19256 = ~n19254 & n19255;
  assign n19257 = ~n18930 & ~n18936;
  assign n19258 = ~n19256 & n19257;
  assign n19259 = ~n18923 & ~n18929;
  assign n19260 = ~n19258 & n19259;
  assign n19261 = ~n18916 & ~n18922;
  assign n19262 = ~n19260 & n19261;
  assign n19263 = ~n18909 & ~n18915;
  assign n19264 = ~n19262 & n19263;
  assign n19265 = ~n18902 & ~n18908;
  assign n19266 = ~n19264 & n19265;
  assign n19267 = ~n18895 & ~n18901;
  assign n19268 = ~n19266 & n19267;
  assign n19269 = ~n18888 & ~n18894;
  assign n19270 = ~n19268 & n19269;
  assign n19271 = ~n18881 & ~n18887;
  assign n19272 = ~n19270 & n19271;
  assign n19273 = ~n18874 & ~n18880;
  assign n19274 = ~n19272 & n19273;
  assign n19275 = ~n18867 & ~n18873;
  assign n19276 = ~n19274 & n19275;
  assign n19277 = ~n18860 & ~n18866;
  assign n19278 = ~n19276 & n19277;
  assign n19279 = ~n18853 & ~n18859;
  assign n19280 = ~n19278 & n19279;
  assign n19281 = ~n18846 & ~n18852;
  assign n19282 = ~n19280 & n19281;
  assign n19283 = ~n18839 & ~n18845;
  assign n19284 = ~n19282 & n19283;
  assign n19285 = ~n18832 & ~n18838;
  assign n19286 = ~n19284 & n19285;
  assign n19287 = ~n18825 & ~n18831;
  assign n19288 = ~n19286 & n19287;
  assign n19289 = ~n18818 & ~n18824;
  assign n19290 = ~n19288 & n19289;
  assign n19291 = ~n18811 & ~n18817;
  assign n19292 = ~n19290 & n19291;
  assign n19293 = ~n18804 & ~n18810;
  assign n19294 = ~n19292 & n19293;
  assign n19295 = ~n18797 & ~n18803;
  assign n19296 = ~n19294 & n19295;
  assign n19297 = ~n18790 & ~n18796;
  assign n19298 = ~n19296 & n19297;
  assign n19299 = ~n18783 & ~n18789;
  assign n19300 = ~n19298 & n19299;
  assign n19301 = ~n18776 & ~n18782;
  assign n19302 = ~n19300 & n19301;
  assign n19303 = ~n18769 & ~n18775;
  assign n19304 = ~n19302 & n19303;
  assign n19305 = ~n18762 & ~n18768;
  assign n19306 = ~n19304 & n19305;
  assign n19307 = ~n18755 & ~n18761;
  assign n19308 = ~n19306 & n19307;
  assign n19309 = n18733 & po1 ;
  assign n19310 = ~n18738 & ~n19309;
  assign n19311 = ~n18746 & ~n19310;
  assign n19312 = po63  & n19311;
  assign n19313 = po1  & ~n19311;
  assign n19314 = ~n18754 & ~n19313;
  assign n19315 = ~po63  & ~n19314;
  assign n19316 = ~n19312 & ~n19315;
  assign po0  = n19308 | ~n19316;
endmodule
