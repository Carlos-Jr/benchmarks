module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24 ;
  wire n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591,
    n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3626, n3627,
    n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651,
    n3652, n3653, n3654, n3655, n3656, n3657,
    n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681,
    n3682, n3683, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927,
    n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951,
    n3952, n3953, n3954, n3955, n3956, n3957,
    n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987,
    n3988, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4017,
    n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047,
    n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077,
    n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101,
    n4102, n4103, n4104, n4105, n4106, n4107,
    n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131,
    n4132, n4133, n4134, n4135, n4136, n4137,
    n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161,
    n4162, n4163, n4164, n4165, n4166, n4167,
    n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191,
    n4192, n4193, n4194, n4195, n4196, n4197,
    n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251,
    n4252, n4253, n4254, n4255, n4256, n4257,
    n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317,
    n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341,
    n4342, n4343, n4344, n4345, n4346, n4347,
    n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4375, n4376, n4377,
    n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395,
    n4396, n4397, n4398, n4399, n4400, n4401,
    n4402, n4403, n4404, n4405, n4406, n4407,
    n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431,
    n4432, n4433, n4434, n4435, n4436, n4437,
    n4438, n4439, n4440, n4441, n4442, n4443,
    n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4455,
    n4456, n4457, n4458, n4459, n4460, n4461,
    n4462, n4463, n4464, n4465, n4466, n4467,
    n4468, n4469, n4470, n4471, n4472, n4473,
    n4474, n4475, n4476, n4477, n4478, n4479,
    n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491,
    n4492, n4493, n4494, n4495, n4496, n4497,
    n4498, n4499, n4500, n4501, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4520, n4521,
    n4522, n4523, n4524, n4525, n4526, n4527,
    n4528, n4529, n4530, n4531, n4532, n4533,
    n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551,
    n4552, n4553, n4554, n4555, n4556, n4557,
    n4558, n4559, n4560, n4561, n4562, n4563,
    n4564, n4565, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581,
    n4582, n4583, n4584, n4585, n4586, n4587,
    n4588, n4589, n4590, n4591, n4592, n4593,
    n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611,
    n4612, n4613, n4614, n4615, n4616, n4617,
    n4618, n4619, n4620, n4621, n4622, n4623,
    n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641,
    n4642, n4643, n4644, n4645, n4646, n4647,
    n4648, n4649, n4650, n4651, n4652, n4653,
    n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671,
    n4672, n4673, n4674, n4675, n4676, n4677,
    n4678, n4679, n4680, n4681, n4682, n4683,
    n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737,
    n4738, n4739, n4740, n4741, n4742, n4743,
    n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4763, n4764, n4765, n4766, n4767,
    n4768, n4769, n4770, n4771, n4772, n4773,
    n4774, n4775, n4776, n4777, n4778, n4779,
    n4780, n4781, n4782, n4783, n4784, n4785,
    n4786, n4787, n4788, n4789, n4790, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797,
    n4798, n4799, n4800, n4801, n4802, n4803,
    n4804, n4805, n4806, n4807, n4808, n4809,
    n4810, n4811, n4812, n4813, n4814, n4815,
    n4816, n4817, n4818, n4819, n4820, n4821,
    n4822, n4823, n4824, n4825, n4826, n4827,
    n4828, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845,
    n4846, n4847, n4848, n4849, n4850, n4851,
    n4852, n4853, n4854, n4855, n4856, n4857,
    n4858, n4859, n4860, n4861, n4862, n4863,
    n4864, n4865, n4866, n4867, n4868, n4869,
    n4870, n4871, n4872, n4873, n4874, n4875,
    n4876, n4877, n4878, n4879, n4880, n4881,
    n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4889, n4890, n4891, n4892, n4893,
    n4894, n4895, n4896, n4897, n4898, n4899,
    n4900, n4901, n4902, n4903, n4904, n4905,
    n4906, n4907, n4908, n4909, n4910, n4911,
    n4912, n4913, n4914, n4915, n4916, n4917,
    n4918, n4919, n4920, n4921, n4922, n4923,
    n4924, n4925, n4926, n4927, n4928, n4929,
    n4930, n4931, n4932, n4933, n4934, n4935,
    n4936, n4937, n4938, n4939, n4940, n4941,
    n4942, n4943, n4944, n4945, n4946, n4947,
    n4948, n4949, n4950, n4951, n4952, n4953,
    n4954, n4955, n4956, n4957, n4958, n4959,
    n4960, n4961, n4962, n4963, n4964, n4965,
    n4966, n4967, n4968, n4969, n4970, n4971,
    n4972, n4973, n4974, n4975, n4976, n4977,
    n4978, n4979, n4980, n4981, n4982, n4983,
    n4984, n4985, n4986, n4987, n4988, n4989,
    n4990, n4991, n4992, n4993, n4994, n4995,
    n4996, n4997, n4998, n4999, n5000, n5001,
    n5002, n5003, n5004, n5005, n5006, n5007,
    n5008, n5009, n5010, n5011, n5012, n5013,
    n5014, n5015, n5016, n5017, n5018, n5019,
    n5020, n5021, n5022, n5023, n5024, n5025,
    n5026, n5027, n5028, n5029, n5030, n5031,
    n5032, n5033, n5034, n5035, n5036, n5037,
    n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049,
    n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061,
    n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151,
    n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217,
    n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5244, n5245, n5246, n5247,
    n5248, n5249, n5250, n5251, n5252, n5253,
    n5254, n5255, n5256, n5257, n5258, n5259,
    n5260, n5261, n5262, n5263, n5264, n5265,
    n5266, n5267, n5268, n5269, n5270, n5271,
    n5272, n5273, n5274, n5275, n5276, n5277,
    n5278, n5279, n5280, n5281, n5282, n5283,
    n5284, n5285, n5286, n5287, n5288, n5289,
    n5290, n5291, n5292, n5293, n5294, n5295,
    n5296, n5297, n5298, n5299, n5300, n5301,
    n5302, n5303, n5304, n5305, n5306, n5307,
    n5308, n5309, n5310, n5311, n5312, n5313,
    n5314, n5315, n5316, n5317, n5318, n5319,
    n5320, n5321, n5322, n5323, n5324, n5325,
    n5326, n5327, n5328, n5329, n5330, n5331,
    n5332, n5333, n5334, n5335, n5336, n5337,
    n5338, n5339, n5340, n5341, n5342, n5343,
    n5344, n5345, n5346, n5347, n5348, n5349,
    n5350, n5351, n5352, n5353, n5354, n5355,
    n5356, n5357, n5358, n5359, n5360, n5361,
    n5362, n5363, n5364, n5365, n5366, n5367,
    n5368, n5369, n5370, n5371, n5372, n5373,
    n5374, n5375, n5376, n5377, n5378, n5379,
    n5380, n5381, n5382, n5383, n5384, n5385,
    n5386, n5387, n5388, n5389, n5390, n5391,
    n5392, n5393, n5394, n5395, n5396, n5397,
    n5398, n5399, n5400, n5401, n5402, n5403,
    n5404, n5405, n5406, n5407, n5408, n5409,
    n5410, n5411, n5412, n5413, n5414, n5415,
    n5416, n5417, n5418, n5419, n5420, n5421,
    n5422, n5423, n5424, n5425, n5426, n5427,
    n5428, n5429, n5430, n5431, n5432, n5433,
    n5434, n5435, n5436, n5437, n5438, n5439,
    n5440, n5441, n5442, n5443, n5444, n5445,
    n5446, n5447, n5448, n5449, n5450, n5451,
    n5452, n5453, n5454, n5455, n5456, n5457,
    n5458, n5459, n5460, n5461, n5462, n5463,
    n5464, n5465, n5466, n5467, n5468, n5469,
    n5470, n5471, n5472, n5473, n5474, n5475,
    n5476, n5477, n5478, n5479, n5480, n5481,
    n5482, n5483, n5484, n5485, n5486, n5487,
    n5488, n5489, n5490, n5491, n5492, n5493,
    n5494, n5495, n5496, n5497, n5498, n5499,
    n5500, n5501, n5502, n5503, n5504, n5505,
    n5506, n5507, n5508, n5509, n5510, n5511,
    n5512, n5513, n5514, n5515, n5516, n5517,
    n5518, n5519, n5520, n5521, n5522, n5523,
    n5524, n5525, n5526, n5527, n5528, n5529,
    n5530, n5531, n5532, n5533, n5534, n5535,
    n5536, n5537, n5538, n5539, n5540, n5541,
    n5542, n5543, n5544, n5545, n5546, n5547,
    n5548, n5549, n5550, n5551, n5552, n5553,
    n5554, n5555, n5556, n5557, n5558, n5559,
    n5560, n5561, n5562, n5563, n5564, n5565,
    n5566, n5567, n5568, n5569, n5570, n5571,
    n5572, n5573, n5574, n5575, n5576, n5577,
    n5578, n5579, n5580, n5581, n5582, n5583,
    n5584, n5585, n5586, n5587, n5588, n5589,
    n5590, n5591, n5592, n5593, n5594, n5595,
    n5596, n5597, n5598, n5599, n5600, n5601,
    n5602, n5603, n5604, n5605, n5606, n5607,
    n5608, n5609, n5610, n5611, n5612, n5613,
    n5614, n5615, n5616, n5617, n5618, n5619,
    n5620, n5621, n5622, n5623, n5624, n5625,
    n5626, n5627, n5628, n5629, n5630, n5631,
    n5632, n5633, n5634, n5635, n5636, n5637,
    n5638, n5639, n5640, n5641, n5642, n5643,
    n5644, n5645, n5646, n5647, n5648, n5649,
    n5650, n5651, n5652, n5653, n5654, n5655,
    n5656, n5657, n5658, n5659, n5660, n5661,
    n5662, n5663, n5664, n5665, n5666, n5667,
    n5668, n5669, n5670, n5671, n5672, n5673,
    n5674, n5675, n5676, n5677, n5678, n5679,
    n5680, n5681, n5682, n5683, n5684, n5685,
    n5686, n5687, n5688, n5689, n5690, n5691,
    n5692, n5693, n5694, n5695, n5696, n5697,
    n5698, n5699, n5700, n5701, n5702, n5703,
    n5704, n5705, n5706, n5707, n5708, n5709,
    n5710, n5711, n5712, n5713, n5714, n5715,
    n5716, n5717, n5718, n5719, n5720, n5721,
    n5722, n5723, n5724, n5725, n5726, n5727,
    n5728, n5729, n5730, n5731, n5732, n5733,
    n5734, n5735, n5736, n5737, n5738, n5739,
    n5740, n5741, n5742, n5743, n5744, n5745,
    n5746, n5747, n5748, n5749, n5750, n5751,
    n5752, n5753, n5754, n5755, n5756, n5757,
    n5758, n5759, n5760, n5761, n5762, n5763,
    n5764, n5765, n5766, n5767, n5768, n5769,
    n5770, n5771, n5772, n5773, n5774, n5775,
    n5776, n5777, n5778, n5779, n5780, n5781,
    n5782, n5783, n5784, n5785, n5786, n5787,
    n5788, n5789, n5790, n5791, n5792, n5793,
    n5794, n5795, n5796, n5797, n5798, n5799,
    n5800, n5801, n5802, n5803, n5804, n5805,
    n5806, n5807, n5808, n5809, n5810, n5811,
    n5812, n5813, n5814, n5815, n5816, n5817,
    n5818, n5819, n5820, n5821, n5822, n5823,
    n5824, n5825, n5826, n5827, n5828, n5829,
    n5830, n5831, n5832, n5833, n5834, n5835,
    n5836, n5837, n5838, n5839, n5840, n5841,
    n5842, n5843, n5844, n5845, n5846, n5847,
    n5848, n5849, n5850, n5851, n5852, n5853,
    n5854, n5855, n5856, n5857, n5858, n5859,
    n5860, n5861, n5862, n5863, n5864, n5865,
    n5866, n5867, n5868, n5869, n5870, n5871,
    n5872, n5873, n5874, n5875, n5876, n5877,
    n5878, n5879, n5880, n5881, n5882, n5883,
    n5884, n5885, n5886, n5887, n5888, n5889,
    n5890, n5891, n5892, n5893, n5894, n5895,
    n5896, n5897, n5898, n5899, n5900, n5901,
    n5902, n5903, n5904, n5905, n5906, n5907,
    n5908, n5909, n5910, n5911, n5912, n5913,
    n5914, n5915, n5916, n5917, n5918, n5919,
    n5920, n5921, n5922, n5923, n5924, n5925,
    n5926, n5927, n5928, n5929, n5930, n5931,
    n5932, n5933, n5934, n5935, n5936, n5937,
    n5938, n5939, n5940, n5941, n5942, n5943,
    n5944, n5945, n5946, n5947, n5948, n5949,
    n5950, n5951, n5952, n5953, n5954, n5955,
    n5956, n5957, n5958, n5959, n5960, n5961,
    n5962, n5963, n5964, n5965, n5966, n5967,
    n5968, n5969, n5970, n5971, n5972, n5973,
    n5974, n5975, n5976, n5977, n5978, n5979,
    n5980, n5981, n5982, n5983, n5984, n5985,
    n5986, n5987, n5988, n5989, n5990, n5991,
    n5992, n5993, n5994, n5995, n5996, n5997,
    n5998, n5999, n6000, n6001, n6002, n6003,
    n6004, n6005, n6006, n6007, n6008, n6009,
    n6010, n6011, n6012, n6013, n6014, n6015,
    n6016, n6017, n6018, n6019, n6020, n6021,
    n6022, n6023, n6024, n6025, n6026, n6027,
    n6028, n6029, n6030, n6031, n6032, n6033,
    n6034, n6035, n6036, n6037, n6038, n6039,
    n6040, n6041, n6042, n6043, n6044, n6045,
    n6046, n6047, n6048, n6049, n6050, n6051,
    n6052, n6053, n6054, n6055, n6056, n6057,
    n6058, n6059, n6060, n6061, n6062, n6063,
    n6064, n6065, n6066, n6067, n6068, n6069,
    n6070, n6071, n6072, n6073, n6074, n6075,
    n6076, n6077, n6078, n6079, n6080, n6081,
    n6082, n6083, n6084, n6085, n6086, n6087,
    n6088, n6089, n6090, n6091, n6092, n6093,
    n6094, n6095, n6096, n6097, n6098, n6099,
    n6100, n6101, n6102, n6103, n6104, n6105,
    n6106, n6107, n6108, n6109, n6110, n6111,
    n6112, n6113, n6114, n6115, n6116, n6117,
    n6118, n6119, n6120, n6121, n6122, n6123,
    n6124, n6125, n6126, n6127, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6139, n6140, n6141,
    n6142, n6143, n6144, n6145, n6146, n6147,
    n6148, n6149, n6150, n6151, n6152, n6153,
    n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6165,
    n6166, n6167, n6168, n6169, n6170, n6171,
    n6172, n6173, n6174, n6175, n6176, n6177,
    n6178, n6179, n6180, n6181, n6182, n6183,
    n6184, n6185, n6186, n6187, n6188, n6189,
    n6190, n6191, n6192, n6193, n6194, n6195,
    n6196, n6197, n6198, n6199, n6200, n6201,
    n6202, n6203, n6204, n6205, n6206, n6207,
    n6208, n6209, n6210, n6211, n6212, n6213,
    n6214, n6215, n6216, n6217, n6218, n6219,
    n6220, n6221, n6222, n6223, n6224, n6225,
    n6226, n6227, n6228, n6229, n6230, n6231,
    n6232, n6233, n6234, n6235, n6236, n6237,
    n6238, n6239, n6240, n6241, n6242, n6243,
    n6244, n6245, n6246, n6247, n6248, n6249,
    n6250, n6251, n6252, n6253, n6254, n6255,
    n6256, n6257, n6258, n6259, n6260, n6261,
    n6262, n6263, n6264, n6265, n6266, n6267,
    n6268, n6269, n6270, n6271, n6272, n6273,
    n6274, n6275, n6276, n6277, n6278, n6279,
    n6280, n6281, n6282, n6283, n6284, n6285,
    n6286, n6287, n6288, n6289, n6290, n6291,
    n6292, n6293, n6294, n6295, n6296, n6297,
    n6298, n6299, n6300, n6301, n6302, n6303,
    n6304, n6305, n6306, n6307, n6308, n6309,
    n6310, n6311, n6312, n6313, n6314, n6315,
    n6316, n6317, n6318, n6319, n6320, n6321,
    n6322, n6323, n6324, n6325, n6326, n6327,
    n6328, n6329, n6330, n6331, n6332, n6333,
    n6334, n6335, n6336, n6337, n6338, n6339,
    n6340, n6341, n6342, n6343, n6344, n6345,
    n6346, n6347, n6348, n6349, n6350, n6351,
    n6352, n6353, n6354, n6355, n6356, n6357,
    n6358, n6359, n6360, n6361, n6362, n6363,
    n6364, n6365, n6366, n6367, n6368, n6369,
    n6370, n6371, n6372, n6373, n6374, n6375,
    n6376, n6377, n6378, n6379, n6380, n6381,
    n6382, n6383, n6384, n6385, n6386, n6387,
    n6388, n6389, n6390, n6391, n6392, n6393,
    n6394, n6395, n6396, n6397, n6398, n6399,
    n6400, n6401, n6402, n6403, n6404, n6405,
    n6406, n6407, n6408, n6409, n6410, n6411,
    n6412, n6413, n6414, n6415, n6416, n6417,
    n6418, n6419, n6420, n6421, n6422, n6423,
    n6424, n6425, n6426, n6427, n6428, n6429,
    n6430, n6431, n6432, n6433, n6434, n6435,
    n6436, n6437, n6438, n6439, n6440, n6441,
    n6442, n6443, n6444, n6445, n6446, n6447,
    n6448, n6449, n6450, n6451, n6452, n6453,
    n6454, n6455, n6456, n6457, n6458, n6459,
    n6460, n6461, n6462, n6463, n6464, n6465,
    n6466, n6467, n6468, n6469, n6470, n6471,
    n6472, n6473, n6474, n6475, n6476, n6477,
    n6478, n6479, n6480, n6481, n6482, n6483,
    n6484, n6485, n6486, n6487, n6488, n6489,
    n6490, n6491, n6492, n6493, n6494, n6495,
    n6496, n6497, n6498, n6499, n6500, n6501,
    n6502, n6503, n6504, n6505, n6506, n6507,
    n6508, n6509, n6510, n6511, n6512, n6513,
    n6514, n6515, n6516, n6517, n6518, n6519,
    n6520, n6521, n6522, n6523, n6524, n6525,
    n6526, n6527, n6528, n6529, n6530, n6531,
    n6532, n6533, n6534, n6535, n6536, n6537,
    n6538, n6539, n6540, n6541, n6542, n6543,
    n6544, n6545, n6546, n6547, n6548, n6549,
    n6550, n6551, n6552, n6553, n6554, n6555,
    n6556, n6557, n6558, n6559, n6560, n6561,
    n6562, n6563, n6564, n6565, n6566, n6567,
    n6568, n6569, n6570, n6571, n6572, n6573,
    n6574, n6575, n6576, n6577, n6578, n6579,
    n6580, n6581, n6582, n6583, n6584, n6585,
    n6586, n6587, n6588, n6589, n6590, n6591,
    n6592, n6593, n6594, n6595, n6596, n6597,
    n6598, n6599, n6600, n6601, n6602, n6603,
    n6604, n6605, n6606, n6607, n6608, n6609,
    n6610, n6611, n6612, n6613, n6614, n6615,
    n6616, n6617, n6618, n6619, n6620, n6621,
    n6622, n6623, n6624, n6625, n6626, n6627,
    n6628, n6629, n6630, n6631, n6632, n6633,
    n6634, n6635, n6636, n6637, n6638, n6639,
    n6640, n6641, n6642, n6643, n6644, n6645,
    n6646, n6647, n6648, n6649, n6650, n6651,
    n6652, n6653, n6654, n6655, n6656, n6657,
    n6658, n6659, n6660, n6661, n6662, n6663,
    n6664, n6665, n6666, n6667, n6668, n6669,
    n6670, n6671, n6672, n6673, n6674, n6675,
    n6676, n6677, n6678, n6679, n6680, n6681,
    n6682, n6683, n6684, n6685, n6686, n6687,
    n6688, n6689, n6690, n6691, n6692, n6693,
    n6694, n6695, n6696, n6697, n6698, n6699,
    n6700, n6701, n6702, n6703, n6704, n6705,
    n6706, n6707, n6708, n6709, n6710, n6711,
    n6712, n6713, n6714, n6715, n6716, n6717,
    n6718, n6719, n6720, n6721, n6722, n6723,
    n6724, n6725, n6726, n6727, n6728, n6729,
    n6730, n6731, n6732, n6733, n6734, n6735,
    n6736, n6737, n6738, n6739, n6740, n6741,
    n6742, n6743, n6744, n6745, n6746, n6747,
    n6748, n6749, n6750, n6751, n6752, n6753,
    n6754, n6755, n6756, n6757, n6758, n6759,
    n6760, n6761, n6762, n6763, n6764, n6765,
    n6766, n6767, n6768, n6769, n6770, n6771,
    n6772, n6773, n6774, n6775, n6776, n6777,
    n6778, n6779, n6780, n6781, n6782, n6783,
    n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801,
    n6802, n6803, n6804, n6805, n6806, n6807,
    n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843,
    n6844, n6845, n6846, n6847, n6848, n6849,
    n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861,
    n6862, n6863, n6864, n6865, n6866, n6867,
    n6868, n6869, n6870, n6871, n6872, n6873,
    n6874, n6875, n6876, n6877, n6878, n6879,
    n6880, n6881, n6882, n6883, n6884, n6885,
    n6886, n6887, n6888, n6889, n6890, n6891,
    n6892, n6893, n6894, n6895, n6896, n6897,
    n6898, n6899, n6900, n6901, n6902, n6903,
    n6904, n6905, n6906, n6907, n6908, n6909,
    n6910, n6911, n6912, n6913, n6914, n6915,
    n6916, n6917, n6918, n6919, n6920, n6921,
    n6922, n6923, n6924, n6925, n6926, n6927,
    n6928, n6929, n6930, n6931, n6932, n6933,
    n6934, n6935, n6936, n6937, n6938, n6939,
    n6940, n6941, n6942, n6943, n6944, n6945,
    n6946, n6947, n6948, n6949, n6950, n6951,
    n6952, n6953, n6954, n6955, n6956, n6957,
    n6958, n6959, n6960, n6961, n6962, n6963,
    n6964, n6965, n6966, n6967, n6968, n6969,
    n6970, n6971, n6972, n6973, n6974, n6975,
    n6976, n6977, n6978, n6979, n6980, n6981,
    n6982, n6983, n6984, n6985, n6986, n6987,
    n6988, n6989, n6990, n6991, n6992, n6993,
    n6994, n6995, n6996, n6997, n6998, n6999,
    n7000, n7001, n7002, n7003, n7004, n7005,
    n7006, n7007, n7008, n7009, n7010, n7011,
    n7012, n7013, n7014, n7015, n7016, n7017,
    n7018, n7019, n7020, n7021, n7022, n7023,
    n7024, n7025, n7026, n7027, n7028, n7029,
    n7030, n7031, n7032, n7033, n7034, n7035,
    n7036, n7037, n7038, n7039, n7040, n7041,
    n7042, n7043, n7044, n7045, n7046, n7047,
    n7048, n7049, n7050, n7051, n7052, n7053,
    n7054, n7055, n7056, n7057, n7058, n7059,
    n7060, n7061, n7062, n7063, n7064, n7065,
    n7066, n7067, n7068, n7069, n7070, n7071,
    n7072, n7073, n7074, n7075, n7076, n7077,
    n7078, n7079, n7080, n7081, n7082, n7083,
    n7084, n7085, n7086, n7087, n7088, n7089,
    n7090, n7091, n7092, n7093, n7094, n7095,
    n7096, n7097, n7098, n7099, n7100, n7101,
    n7102, n7103, n7104, n7105, n7106, n7107,
    n7108, n7109, n7110, n7111, n7112, n7113,
    n7114, n7115, n7116, n7117, n7118, n7119,
    n7120, n7121, n7122, n7123, n7124, n7125,
    n7126, n7127, n7128, n7129, n7130, n7131,
    n7132, n7133, n7134, n7135, n7136, n7137,
    n7138, n7139, n7140, n7141, n7142, n7143,
    n7144, n7145, n7146, n7147, n7148, n7149,
    n7150, n7151, n7152, n7153, n7154, n7155,
    n7156, n7157, n7158, n7159, n7160, n7161,
    n7162, n7163, n7164, n7165, n7166, n7167,
    n7168, n7169, n7170, n7171, n7172, n7173,
    n7174, n7175, n7176, n7177, n7178, n7179,
    n7180, n7181, n7182, n7183, n7184, n7185,
    n7186, n7187, n7188, n7189, n7190, n7191,
    n7192, n7193, n7194, n7195, n7196, n7197,
    n7198, n7199, n7200, n7201, n7202, n7203,
    n7204, n7205, n7206, n7207, n7208, n7209,
    n7210, n7211, n7212, n7213, n7214, n7215,
    n7216, n7217, n7218, n7219, n7220, n7221,
    n7222, n7223, n7224, n7225, n7226, n7227,
    n7228, n7229, n7230, n7231, n7232, n7233,
    n7234, n7235, n7236, n7237, n7238, n7239,
    n7240, n7241, n7242, n7243, n7244, n7245,
    n7246, n7247, n7248, n7249, n7250, n7251,
    n7252, n7253, n7254, n7255, n7256, n7257,
    n7258, n7259, n7260, n7261, n7262, n7263,
    n7264, n7265, n7266, n7267, n7268, n7269,
    n7270, n7271, n7272, n7273, n7274, n7275,
    n7276, n7277, n7278, n7279, n7280, n7281,
    n7282, n7283, n7284, n7285, n7286, n7287,
    n7288, n7289, n7290, n7291, n7292, n7293,
    n7294, n7295, n7296, n7297, n7298, n7299,
    n7300, n7301, n7302, n7303, n7304, n7305,
    n7306, n7307, n7308, n7309, n7310, n7311,
    n7312, n7313, n7314, n7315, n7316, n7317,
    n7318, n7319, n7320, n7321, n7322, n7323,
    n7324, n7325, n7326, n7327, n7328, n7329,
    n7330, n7331, n7332, n7333, n7334, n7335,
    n7336, n7337, n7338, n7339, n7340, n7341,
    n7342, n7343, n7344, n7345, n7346, n7347,
    n7348, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7357, n7358, n7359,
    n7360, n7361, n7362, n7363, n7364, n7365,
    n7366, n7367, n7368, n7369, n7370, n7371,
    n7372, n7373, n7374, n7375, n7376, n7377,
    n7378, n7379, n7380, n7381, n7382, n7383,
    n7384, n7385, n7386, n7387, n7388, n7389,
    n7390, n7391, n7392, n7393, n7394, n7395,
    n7396, n7397, n7398, n7399, n7400, n7401,
    n7402, n7403, n7404, n7405, n7406, n7407,
    n7408, n7409, n7410, n7411, n7412, n7413,
    n7414, n7415, n7416, n7417, n7418, n7419,
    n7420, n7421, n7422, n7423, n7424, n7425,
    n7426, n7427, n7428, n7429, n7430, n7431,
    n7432, n7433, n7434, n7435, n7436, n7437,
    n7438, n7439, n7440, n7441, n7442, n7443,
    n7444, n7445, n7446, n7447, n7448, n7449,
    n7450, n7451, n7452, n7453, n7454, n7455,
    n7456, n7457, n7458, n7459, n7460, n7461,
    n7462, n7463, n7464, n7465, n7466, n7467,
    n7468, n7469, n7470, n7471, n7472, n7473,
    n7474, n7475, n7476, n7477, n7478, n7479,
    n7480, n7481, n7482, n7483, n7484, n7485,
    n7486, n7487, n7488, n7489, n7490, n7491,
    n7492, n7493, n7494, n7495, n7496, n7497,
    n7498, n7499, n7500, n7501, n7502, n7503,
    n7504, n7505, n7506, n7507, n7508, n7509,
    n7510, n7511, n7512, n7513, n7514, n7515,
    n7516, n7517, n7518, n7519, n7520, n7521,
    n7522, n7523, n7524, n7525, n7526, n7527,
    n7528, n7529, n7530, n7531, n7532, n7533,
    n7534, n7535, n7536, n7537, n7538, n7539,
    n7540, n7541, n7542, n7543, n7544, n7545,
    n7546, n7547, n7548, n7549, n7550, n7551,
    n7552, n7553, n7554, n7555, n7556, n7557,
    n7558, n7559, n7560, n7561, n7562, n7563,
    n7564, n7565, n7566, n7567, n7568, n7569,
    n7570, n7571, n7572, n7573, n7574, n7575,
    n7576, n7577, n7578, n7579, n7580, n7581,
    n7582, n7583, n7584, n7585, n7586, n7587,
    n7588, n7589, n7590, n7591, n7592, n7593,
    n7594, n7595, n7596, n7597, n7598, n7599,
    n7600, n7601, n7602, n7603, n7604, n7605,
    n7606, n7607, n7608, n7609, n7610, n7611,
    n7612, n7613, n7614, n7615, n7616, n7617,
    n7618, n7619, n7621, n7622, n7623, n7624,
    n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636,
    n7637, n7638, n7639, n7640, n7641, n7642,
    n7643, n7644, n7645, n7646, n7647, n7648,
    n7649, n7650, n7651, n7652, n7653, n7654,
    n7655, n7656, n7657, n7658, n7659, n7660,
    n7661, n7662, n7663, n7664, n7665, n7666,
    n7667, n7668, n7669, n7670, n7671, n7672,
    n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7684,
    n7685, n7686, n7687, n7688, n7689, n7690,
    n7691, n7692, n7693, n7694, n7695, n7696,
    n7697, n7698, n7699, n7700, n7701, n7702,
    n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714,
    n7715, n7716, n7717, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726,
    n7727, n7728, n7729, n7730, n7731, n7732,
    n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744,
    n7745, n7746, n7747, n7748, n7749, n7750,
    n7751, n7752, n7753, n7754, n7755, n7756,
    n7757, n7758, n7759, n7760, n7761, n7762,
    n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7786,
    n7787, n7788, n7789, n7790, n7791, n7792,
    n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7813, n7814, n7815, n7816,
    n7817, n7818, n7819, n7820, n7821, n7822,
    n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062,
    n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8090, n8091, n8092,
    n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104,
    n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116,
    n8117, n8118, n8119, n8120, n8121, n8122,
    n8123, n8124, n8125, n8126, n8127, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134,
    n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146,
    n8147, n8148, n8149, n8150, n8151, n8152,
    n8153, n8154, n8155, n8156, n8157, n8158,
    n8159, n8160, n8161, n8162, n8163, n8164,
    n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176,
    n8177, n8178, n8179, n8180, n8181, n8182,
    n8183, n8184, n8185, n8186, n8187, n8188,
    n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206,
    n8207, n8208, n8209, n8210, n8211, n8212,
    n8213, n8214, n8215, n8216, n8217, n8218,
    n8219, n8220, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236,
    n8237, n8238, n8239, n8240, n8241, n8242,
    n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8272,
    n8273, n8274, n8275, n8276, n8277, n8278,
    n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296,
    n8297, n8298, n8299, n8300, n8301, n8302,
    n8303, n8304, n8305, n8306, n8307, n8308,
    n8309, n8310, n8311, n8312, n8313, n8314,
    n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326,
    n8327, n8328, n8329, n8330, n8331, n8332,
    n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356,
    n8357, n8358, n8359, n8360, n8361, n8362,
    n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8371, n8372, n8373, n8374,
    n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386,
    n8387, n8388, n8389, n8390, n8391, n8392,
    n8393, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404,
    n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416,
    n8417, n8418, n8419, n8420, n8421, n8422,
    n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434,
    n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446,
    n8447, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476,
    n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8596,
    n8597, n8598, n8599, n8600, n8601, n8602,
    n8603, n8604, n8605, n8606, n8607, n8608,
    n8609, n8610, n8611, n8612, n8613, n8614,
    n8615, n8616, n8617, n8618, n8619, n8620,
    n8621, n8622, n8623, n8624, n8625, n8626,
    n8627, n8628, n8629, n8630, n8631, n8632,
    n8633, n8634, n8635, n8636, n8637, n8638,
    n8639, n8640, n8641, n8642, n8643, n8644,
    n8645, n8646, n8647, n8648, n8649, n8650,
    n8651, n8652, n8653, n8654, n8655, n8656,
    n8657, n8658, n8659, n8660, n8661, n8662,
    n8663, n8664, n8665, n8666, n8667, n8668,
    n8669, n8670, n8671, n8672, n8673, n8674,
    n8675, n8676, n8677, n8678, n8679, n8680,
    n8681, n8682, n8683, n8684, n8685, n8686,
    n8687, n8688, n8689, n8690, n8691, n8692,
    n8693, n8694, n8695, n8696, n8697, n8698,
    n8699, n8700, n8701, n8702, n8703, n8704,
    n8705, n8706, n8707, n8708, n8709, n8710,
    n8711, n8712, n8713, n8714, n8715, n8716,
    n8717, n8718, n8719, n8720, n8721, n8722,
    n8723, n8724, n8725, n8726, n8727, n8728,
    n8729, n8730, n8731, n8732, n8733, n8734,
    n8735, n8736, n8737, n8738, n8739, n8740,
    n8741, n8742, n8743, n8744, n8745, n8746,
    n8747, n8748, n8749, n8750, n8751, n8752,
    n8753, n8754, n8755, n8756, n8757, n8758,
    n8759, n8760, n8761, n8762, n8763, n8764,
    n8765, n8766, n8767, n8768, n8769, n8770,
    n8771, n8772, n8773, n8774, n8775, n8776,
    n8777, n8778, n8779, n8780, n8781, n8782,
    n8783, n8784, n8785, n8786, n8787, n8788,
    n8789, n8790, n8791, n8792, n8793, n8794,
    n8795, n8796, n8797, n8798, n8799, n8800,
    n8801, n8802, n8803, n8804, n8805, n8806,
    n8807, n8808, n8809, n8810, n8811, n8812,
    n8813, n8814, n8815, n8816, n8817, n8818,
    n8819, n8820, n8821, n8822, n8823, n8824,
    n8825, n8826, n8827, n8828, n8829, n8830,
    n8831, n8832, n8833, n8834, n8835, n8836,
    n8837, n8838, n8839, n8840, n8841, n8842,
    n8843, n8844, n8845, n8846, n8847, n8848,
    n8849, n8850, n8851, n8852, n8853, n8854,
    n8855, n8856, n8857, n8858, n8859, n8860,
    n8861, n8862, n8863, n8864, n8865, n8866,
    n8867, n8868, n8869, n8870, n8871, n8872,
    n8873, n8874, n8875, n8876, n8877, n8878,
    n8879, n8880, n8881, n8882, n8883, n8884,
    n8885, n8886, n8887, n8888, n8889, n8890,
    n8891, n8892, n8893, n8894, n8895, n8896,
    n8897, n8898, n8899, n8900, n8901, n8902,
    n8903, n8904, n8905, n8906, n8907, n8908,
    n8909, n8910, n8911, n8912, n8913, n8914,
    n8915, n8916, n8917, n8918, n8919, n8920,
    n8921, n8922, n8923, n8924, n8925, n8926,
    n8927, n8928, n8929, n8930, n8931, n8932,
    n8933, n8934, n8935, n8936, n8937, n8938,
    n8939, n8940, n8941, n8942, n8943, n8944,
    n8945, n8946, n8947, n8948, n8949, n8950,
    n8951, n8952, n8953, n8954, n8955, n8956,
    n8957, n8958, n8959, n8960, n8961, n8962,
    n8963, n8964, n8965, n8966, n8967, n8968,
    n8969, n8970, n8971, n8972, n8973, n8974,
    n8975, n8976, n8977, n8978, n8979, n8980,
    n8981, n8982, n8983, n8984, n8985, n8986,
    n8987, n8988, n8989, n8990, n8991, n8992,
    n8993, n8994, n8995, n8996, n8997, n8998,
    n8999, n9000, n9001, n9002, n9003, n9004,
    n9005, n9006, n9007, n9008, n9009, n9010,
    n9011, n9012, n9013, n9014, n9015, n9016,
    n9017, n9018, n9019, n9020, n9021, n9022,
    n9023, n9024, n9025, n9026, n9027, n9028,
    n9029, n9030, n9031, n9032, n9033, n9034,
    n9035, n9036, n9037, n9038, n9039, n9040,
    n9041, n9042, n9043, n9044, n9045, n9046,
    n9047, n9048, n9049, n9050, n9051, n9052,
    n9053, n9054, n9055, n9056, n9057, n9058,
    n9059, n9060, n9061, n9062, n9063, n9064,
    n9065, n9066, n9067, n9068, n9069, n9070,
    n9071, n9072, n9073, n9074, n9075, n9076,
    n9077, n9078, n9079, n9080, n9081, n9082,
    n9083, n9084, n9085, n9086, n9087, n9088,
    n9089, n9090, n9091, n9092, n9093, n9094,
    n9095, n9096, n9097, n9098, n9099, n9100,
    n9101, n9102, n9103, n9104, n9105, n9106,
    n9107, n9108, n9109, n9110, n9111, n9112,
    n9113, n9114, n9115, n9116, n9117, n9118,
    n9119, n9120, n9121, n9122, n9123, n9124,
    n9125, n9126, n9127, n9128, n9129, n9130,
    n9131, n9132, n9133, n9134, n9135, n9136,
    n9137, n9138, n9139, n9140, n9141, n9142,
    n9143, n9144, n9145, n9146, n9147, n9148,
    n9149, n9150, n9151, n9152, n9153, n9154,
    n9155, n9156, n9157, n9158, n9159, n9160,
    n9161, n9162, n9163, n9164, n9165, n9166,
    n9167, n9168, n9169, n9170, n9171, n9172,
    n9173, n9174, n9175, n9176, n9177, n9178,
    n9179, n9180, n9181, n9182, n9183, n9184,
    n9185, n9186, n9187, n9188, n9189, n9190,
    n9191, n9192, n9193, n9194, n9195, n9196,
    n9197, n9198, n9199, n9200, n9201, n9202,
    n9203, n9204, n9205, n9206, n9207, n9208,
    n9209, n9210, n9211, n9212, n9213, n9214,
    n9215, n9216, n9217, n9218, n9219, n9220,
    n9221, n9222, n9223, n9224, n9225, n9226,
    n9227, n9228, n9229, n9230, n9231, n9232,
    n9233, n9234, n9235, n9236, n9237, n9238,
    n9239, n9240, n9241, n9242, n9243, n9244,
    n9245, n9246, n9247, n9248, n9249, n9250,
    n9251, n9252, n9253, n9254, n9255, n9256,
    n9257, n9258, n9259, n9260, n9261, n9262,
    n9263, n9264, n9265, n9266, n9267, n9268,
    n9269, n9270, n9271, n9272, n9273, n9274,
    n9275, n9276, n9277, n9278, n9279, n9280,
    n9281, n9282, n9283, n9284, n9285, n9287,
    n9288, n9289, n9290, n9291, n9292, n9293,
    n9294, n9295, n9296, n9297, n9298, n9299,
    n9300, n9301, n9302, n9303, n9304, n9305,
    n9306, n9307, n9308, n9309, n9310, n9311,
    n9312, n9313, n9314, n9315, n9316, n9317,
    n9318, n9319, n9320, n9321, n9322, n9323,
    n9324, n9325, n9326, n9327, n9328, n9329,
    n9330, n9331, n9332, n9333, n9334, n9335,
    n9336, n9337, n9338, n9339, n9340, n9341,
    n9342, n9343, n9344, n9345, n9346, n9347,
    n9348, n9349, n9350, n9351, n9352, n9353,
    n9354, n9355, n9356, n9357, n9358, n9359,
    n9360, n9361, n9362, n9363, n9364, n9365,
    n9366, n9367, n9368, n9369, n9370, n9371,
    n9372, n9373, n9374, n9375, n9376, n9377,
    n9378, n9379, n9380, n9381, n9382, n9383,
    n9384, n9385, n9386, n9387, n9388, n9389,
    n9390, n9391, n9392, n9393, n9394, n9395,
    n9396, n9397, n9398, n9399, n9400, n9401,
    n9402, n9403, n9404, n9405, n9406, n9407,
    n9408, n9409, n9410, n9411, n9412, n9413,
    n9414, n9415, n9416, n9417, n9418, n9419,
    n9420, n9421, n9422, n9423, n9424, n9425,
    n9426, n9427, n9428, n9429, n9430, n9431,
    n9432, n9433, n9434, n9435, n9436, n9437,
    n9438, n9439, n9440, n9441, n9442, n9443,
    n9444, n9445, n9446, n9447, n9448, n9449,
    n9450, n9451, n9452, n9453, n9454, n9455,
    n9456, n9457, n9458, n9459, n9460, n9461,
    n9462, n9463, n9464, n9465, n9466, n9467,
    n9468, n9469, n9470, n9471, n9472, n9473,
    n9474, n9475, n9476, n9477, n9478, n9479,
    n9480, n9481, n9482, n9483, n9484, n9485,
    n9486, n9487, n9488, n9489, n9490, n9491,
    n9492, n9493, n9494, n9495, n9496, n9497,
    n9498, n9499, n9500, n9501, n9502, n9503,
    n9504, n9505, n9506, n9507, n9508, n9509,
    n9510, n9511, n9512, n9513, n9514, n9515,
    n9516, n9517, n9518, n9519, n9520, n9521,
    n9522, n9523, n9524, n9525, n9527, n9528,
    n9529, n9530, n9531, n9532, n9533, n9534,
    n9535, n9536, n9537, n9538, n9539, n9540,
    n9541, n9542, n9543, n9544, n9545, n9546,
    n9547, n9548, n9549, n9550, n9551, n9552,
    n9553, n9554, n9555, n9556, n9557, n9558,
    n9559, n9560, n9561, n9562, n9563, n9564,
    n9565, n9566, n9567, n9568, n9569, n9570,
    n9571, n9572, n9573, n9574, n9575, n9576,
    n9577, n9578, n9579, n9580, n9581, n9582,
    n9583, n9584, n9585, n9586, n9587, n9588,
    n9589, n9590, n9591, n9592, n9593, n9594,
    n9595, n9596, n9597, n9598, n9599, n9600,
    n9601, n9602, n9603, n9604, n9605, n9606,
    n9607, n9608, n9609, n9610, n9611, n9612,
    n9613, n9614, n9615, n9616, n9617, n9618,
    n9619, n9620, n9621, n9622, n9623, n9624,
    n9625, n9626, n9627, n9628, n9629, n9630,
    n9631, n9632, n9633, n9634, n9635, n9636,
    n9637, n9638, n9639, n9640, n9641, n9642,
    n9643, n9644, n9645, n9646, n9647, n9648,
    n9649, n9650, n9651, n9652, n9653, n9654,
    n9655, n9656, n9657, n9658, n9659, n9660,
    n9661, n9662, n9663, n9664, n9665, n9666,
    n9667, n9668, n9669, n9670, n9671, n9672,
    n9673, n9674, n9675, n9676, n9677, n9678,
    n9679, n9680, n9681, n9682, n9683, n9684,
    n9685, n9686, n9687, n9688, n9689, n9690,
    n9691, n9692, n9693, n9694, n9695, n9696,
    n9697, n9698, n9699, n9700, n9701, n9702,
    n9703, n9704, n9705, n9706, n9707, n9708,
    n9709, n9710, n9711, n9712, n9713, n9714,
    n9715, n9716, n9717, n9718, n9719, n9720,
    n9721, n9722, n9723, n9724, n9725, n9726,
    n9727, n9728, n9729, n9730, n9731, n9732,
    n9733, n9734, n9735, n9736, n9737, n9738,
    n9739, n9740, n9741, n9742, n9743, n9744,
    n9745, n9746, n9747, n9748, n9749, n9750,
    n9751, n9752, n9753, n9754, n9755, n9756,
    n9757, n9758, n9759, n9760, n9761, n9762,
    n9763, n9764, n9765, n9766, n9767, n9768,
    n9769, n9770, n9771, n9772, n9773, n9774,
    n9775, n9776, n9777, n9778, n9779, n9780,
    n9781, n9782, n9783, n9784, n9785, n9786,
    n9787, n9788, n9789, n9790, n9791, n9792,
    n9793, n9794, n9795, n9796, n9797, n9798,
    n9799, n9800, n9801, n9802, n9803, n9804,
    n9805, n9806, n9807, n9808, n9809, n9810,
    n9811, n9812, n9813, n9814, n9815, n9816,
    n9817, n9818, n9819, n9820, n9821, n9822,
    n9823, n9824, n9825, n9826, n9827, n9828,
    n9829, n9830, n9831, n9832, n9833, n9834,
    n9835, n9836, n9837, n9838, n9839, n9840,
    n9841, n9842, n9843, n9844, n9845, n9846,
    n9847, n9848, n9849, n9850, n9851, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858,
    n9859, n9860, n9861, n9862, n9863, n9864,
    n9865, n9866, n9867, n9868, n9869, n9870,
    n9871, n9872, n9873, n9874, n9875, n9876,
    n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888,
    n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900,
    n9901, n9902, n9903, n9904, n9905, n9906,
    n9907, n9908, n9909, n9910, n9911, n9912,
    n9913, n9914, n9915, n9916, n9917, n9918,
    n9919, n9920, n9921, n9922, n9923, n9924,
    n9925, n9926, n9927, n9928, n9929, n9930,
    n9931, n9932, n9933, n9934, n9935, n9936,
    n9937, n9938, n9939, n9940, n9941, n9942,
    n9943, n9944, n9945, n9946, n9947, n9948,
    n9949, n9950, n9951, n9952, n9953, n9954,
    n9955, n9956, n9957, n9958, n9959, n9960,
    n9961, n9962, n9963, n9964, n9965, n9966,
    n9967, n9968, n9969, n9970, n9971, n9972,
    n9973, n9974, n9975, n9976, n9977, n9978,
    n9979, n9980, n9981, n9982, n9983, n9984,
    n9985, n9986, n9987, n9988, n9989, n9990,
    n9991, n9992, n9993, n9994, n9995, n9996,
    n9997, n9998, n9999, n10000, n10001, n10002,
    n10003, n10004, n10005, n10006, n10007, n10008,
    n10009, n10010, n10011, n10012, n10013, n10014,
    n10015, n10016, n10017, n10018, n10019, n10020,
    n10021, n10022, n10023, n10024, n10025, n10026,
    n10027, n10028, n10029, n10030, n10031, n10032,
    n10033, n10034, n10035, n10036, n10037, n10038,
    n10039, n10040, n10041, n10042, n10043, n10044,
    n10045, n10046, n10047, n10048, n10049, n10050,
    n10051, n10052, n10053, n10054, n10055, n10056,
    n10057, n10058, n10059, n10060, n10061, n10062,
    n10063, n10064, n10065, n10066, n10067, n10068,
    n10069, n10070, n10071, n10072, n10073, n10074,
    n10075, n10076, n10077, n10078, n10079, n10080,
    n10081, n10082, n10083, n10084, n10085, n10086,
    n10087, n10088, n10089, n10090, n10091, n10092,
    n10093, n10094, n10095, n10096, n10097, n10098,
    n10099, n10100, n10101, n10102, n10103, n10104,
    n10105, n10106, n10107, n10108, n10109, n10110,
    n10111, n10112, n10113, n10114, n10115, n10116,
    n10117, n10118, n10119, n10120, n10121, n10122,
    n10123, n10124, n10125, n10126, n10127, n10128,
    n10129, n10130, n10131, n10132, n10133, n10134,
    n10135, n10136, n10137, n10138, n10139, n10140,
    n10141, n10142, n10143, n10144, n10145, n10146,
    n10147, n10148, n10149, n10150, n10151, n10152,
    n10153, n10154, n10155, n10156, n10157, n10158,
    n10159, n10160, n10161, n10162, n10163, n10164,
    n10165, n10166, n10167, n10168, n10169, n10170,
    n10171, n10172, n10173, n10174, n10175, n10176,
    n10177, n10178, n10179, n10180, n10181, n10182,
    n10183, n10184, n10185, n10186, n10187, n10188,
    n10189, n10190, n10191, n10192, n10193, n10194,
    n10195, n10196, n10197, n10198, n10199, n10200,
    n10201, n10202, n10203, n10204, n10205, n10206,
    n10207, n10208, n10209, n10210, n10211, n10212,
    n10213, n10214, n10215, n10216, n10217, n10218,
    n10219, n10220, n10221, n10222, n10223, n10224,
    n10225, n10226, n10227, n10228, n10229, n10230,
    n10231, n10232, n10233, n10234, n10235, n10236,
    n10237, n10238, n10239, n10240, n10241, n10242,
    n10243, n10244, n10245, n10246, n10247, n10248,
    n10249, n10250, n10251, n10252, n10253, n10254,
    n10255, n10256, n10257, n10258, n10259, n10260,
    n10261, n10262, n10263, n10264, n10265, n10266,
    n10267, n10268, n10269, n10270, n10271, n10272,
    n10273, n10274, n10275, n10276, n10277, n10278,
    n10279, n10280, n10281, n10282, n10283, n10284,
    n10285, n10286, n10287, n10288, n10289, n10290,
    n10291, n10292, n10293, n10294, n10295, n10296,
    n10297, n10298, n10299, n10300, n10301, n10302,
    n10303, n10304, n10305, n10306, n10307, n10308,
    n10309, n10310, n10311, n10312, n10313, n10314,
    n10315, n10316, n10317, n10318, n10319, n10320,
    n10321, n10322, n10323, n10324, n10325, n10326,
    n10327, n10328, n10329, n10330, n10331, n10332,
    n10333, n10334, n10335, n10336, n10337, n10338,
    n10339, n10340, n10341, n10342, n10343, n10344,
    n10345, n10346, n10347, n10348, n10349, n10350,
    n10351, n10352, n10353, n10354, n10355, n10356,
    n10357, n10358, n10359, n10360, n10361, n10362,
    n10363, n10364, n10365, n10366, n10367, n10368,
    n10369, n10370, n10371, n10372, n10373, n10374,
    n10375, n10376, n10377, n10378, n10379, n10380,
    n10381, n10382, n10383, n10384, n10385, n10386,
    n10387, n10388, n10389, n10390, n10391, n10392,
    n10393, n10394, n10395, n10396, n10397, n10398,
    n10399, n10400, n10401, n10402, n10403, n10404,
    n10405, n10406, n10407, n10408, n10409, n10410,
    n10411, n10412, n10413, n10414, n10415, n10416,
    n10417, n10418, n10419, n10420, n10421, n10422,
    n10423, n10424, n10425, n10426, n10427, n10428,
    n10429, n10430, n10431, n10432, n10433, n10434,
    n10435, n10436, n10437, n10438, n10439, n10440,
    n10441, n10442, n10443, n10444, n10445, n10446,
    n10447, n10448, n10449, n10450, n10451, n10452,
    n10453, n10454, n10455, n10456, n10457, n10458,
    n10459, n10460, n10461, n10462, n10463, n10464,
    n10465, n10466, n10467, n10468, n10469, n10470,
    n10471, n10472, n10473, n10474, n10475, n10476,
    n10477, n10478, n10479, n10480, n10481, n10482,
    n10483, n10484, n10485, n10486, n10487, n10488,
    n10489, n10490, n10491, n10492, n10493, n10494,
    n10495, n10496, n10497, n10498, n10499, n10500,
    n10501, n10502, n10503, n10504, n10505, n10506,
    n10507, n10508, n10509, n10510, n10511, n10512,
    n10513, n10514, n10515, n10516, n10517, n10518,
    n10519, n10520, n10521, n10522, n10523, n10524,
    n10525, n10526, n10527, n10528, n10529, n10530,
    n10531, n10532, n10533, n10534, n10535, n10536,
    n10537, n10538, n10539, n10540, n10541, n10542,
    n10543, n10544, n10545, n10546, n10547, n10548,
    n10549, n10550, n10551, n10552, n10553, n10554,
    n10555, n10556, n10557, n10558, n10559, n10560,
    n10561, n10562, n10563, n10564, n10565, n10566,
    n10567, n10568, n10569, n10570, n10571, n10572,
    n10573, n10574, n10575, n10576, n10577, n10578,
    n10579, n10580, n10581, n10582, n10583, n10584,
    n10585, n10586, n10587, n10588, n10589, n10590,
    n10591, n10592, n10593, n10594, n10595, n10596,
    n10597, n10598, n10599, n10600, n10601, n10602,
    n10603, n10604, n10605, n10606, n10607, n10608,
    n10609, n10610, n10611, n10612, n10613, n10614,
    n10615, n10616, n10617, n10618, n10619, n10620,
    n10621, n10622, n10623, n10624, n10625, n10626,
    n10627, n10628, n10629, n10630, n10631, n10632,
    n10633, n10634, n10635, n10636, n10637, n10638,
    n10639, n10640, n10641, n10642, n10643, n10644,
    n10645, n10646, n10647;
  assign n50 = ~pi0  & ~pi1 ;
  assign n51 = ~pi1  & ~pi2 ;
  assign n52 = ~pi0  & n51;
  assign n53 = ~pi2  & n50;
  assign n54 = ~pi3  & n9527;
  assign n55 = ~pi4  & n54;
  assign n56 = ~pi22  & ~n55;
  assign n57 = pi5  & ~n56;
  assign n58 = ~pi5  & n56;
  assign n59 = ~pi5  & ~n56;
  assign n60 = pi5  & n56;
  assign n61 = ~n59 & ~n60;
  assign n62 = ~n57 & ~n58;
  assign n63 = ~pi22  & ~n9527;
  assign n64 = pi3  & ~n63;
  assign n65 = ~pi3  & n63;
  assign n66 = ~pi3  & ~n63;
  assign n67 = pi3  & n63;
  assign n68 = ~n66 & ~n67;
  assign n69 = ~n64 & ~n65;
  assign n70 = pi2  & pi22 ;
  assign n71 = pi2  & ~n50;
  assign n72 = n63 & ~n71;
  assign n73 = ~n70 & ~n72;
  assign n74 = n9529 & ~n73;
  assign n75 = ~n9529 & n73;
  assign n76 = ~n9529 & ~n73;
  assign n77 = n9529 & n73;
  assign n78 = ~n76 & ~n77;
  assign n79 = ~n74 & ~n75;
  assign n80 = pi4  & pi22 ;
  assign n81 = pi4  & ~n54;
  assign n82 = n56 & ~n81;
  assign n83 = ~n80 & ~n82;
  assign n84 = n9528 & ~n83;
  assign n85 = ~n9528 & n83;
  assign n86 = ~n9528 & ~n83;
  assign n87 = n9528 & n83;
  assign n88 = ~n86 & ~n87;
  assign n89 = ~n84 & ~n85;
  assign n90 = ~n9530 & ~n9531;
  assign n91 = ~pi5  & n55;
  assign n92 = ~pi6  & n91;
  assign n93 = ~pi7  & n92;
  assign n94 = ~pi8  & n93;
  assign n95 = ~pi9  & n94;
  assign n96 = ~pi10  & n95;
  assign n97 = ~pi11  & n96;
  assign n98 = ~pi12  & n97;
  assign n99 = ~pi13  & n98;
  assign n100 = ~pi14  & n99;
  assign n101 = ~pi22  & ~n100;
  assign n102 = ~pi15  & ~n101;
  assign n103 = pi15  & n101;
  assign n104 = pi15  & ~n101;
  assign n105 = ~pi15  & n101;
  assign n106 = ~n104 & ~n105;
  assign n107 = pi15  & pi22 ;
  assign n108 = ~pi15  & n100;
  assign n109 = ~pi22  & ~n108;
  assign n110 = pi15  & ~n100;
  assign n111 = n109 & ~n110;
  assign n112 = ~n107 & ~n111;
  assign n113 = ~n102 & ~n103;
  assign n114 = pi20  & pi22 ;
  assign n115 = ~pi16  & n108;
  assign n116 = ~pi17  & n115;
  assign n117 = ~pi18  & n116;
  assign n118 = ~pi19  & n117;
  assign n119 = pi20  & ~n118;
  assign n120 = ~pi20  & n118;
  assign n121 = ~pi22  & ~n120;
  assign n122 = ~n119 & ~n120;
  assign n123 = ~pi22  & n122;
  assign n124 = ~n119 & n121;
  assign n125 = ~n114 & ~n9533;
  assign n126 = ~pi21  & ~n121;
  assign n127 = pi21  & n121;
  assign n128 = pi21  & ~n121;
  assign n129 = ~pi21  & ~pi22 ;
  assign n130 = ~n120 & n129;
  assign n131 = ~n128 & ~n130;
  assign n132 = pi21  & pi22 ;
  assign n133 = pi21  & ~n120;
  assign n134 = ~pi21  & n120;
  assign n135 = ~pi22  & ~n134;
  assign n136 = ~n133 & ~n134;
  assign n137 = ~pi22  & n136;
  assign n138 = ~n133 & n135;
  assign n139 = ~n132 & ~n9535;
  assign n140 = ~n126 & ~n127;
  assign n141 = n125 & ~n9534;
  assign n142 = n9532 & n141;
  assign n143 = ~pi22  & ~n115;
  assign n144 = pi17  & ~n143;
  assign n145 = ~pi17  & n143;
  assign n146 = ~n144 & ~n145;
  assign n147 = pi16  & ~n109;
  assign n148 = ~pi16  & n109;
  assign n149 = ~n147 & ~n148;
  assign n150 = n146 & ~n149;
  assign n151 = pi18  & pi22 ;
  assign n152 = ~pi22  & ~n117;
  assign n153 = pi18  & ~n116;
  assign n154 = n152 & ~n153;
  assign n155 = ~n151 & ~n154;
  assign n156 = pi19  & ~n152;
  assign n157 = ~pi19  & n152;
  assign n158 = ~pi19  & ~n152;
  assign n159 = pi19  & n152;
  assign n160 = ~n158 & ~n159;
  assign n161 = ~n156 & ~n157;
  assign n162 = ~n155 & ~n9536;
  assign n163 = n150 & n162;
  assign n164 = n142 & n163;
  assign n165 = n155 & ~n9536;
  assign n166 = ~n146 & ~n149;
  assign n167 = n165 & n166;
  assign n168 = n141 & n167;
  assign n169 = n142 & n167;
  assign n170 = n9532 & n168;
  assign n171 = ~n164 & ~n9537;
  assign n172 = n146 & n149;
  assign n173 = ~n155 & n9536;
  assign n174 = n172 & n173;
  assign n175 = n142 & n174;
  assign n176 = ~n125 & n9534;
  assign n177 = ~n9532 & n176;
  assign n178 = n150 & n173;
  assign n179 = n177 & n178;
  assign n180 = ~n175 & ~n179;
  assign n181 = ~n9537 & ~n175;
  assign n182 = ~n164 & n181;
  assign n183 = ~n179 & n182;
  assign n184 = ~n164 & ~n175;
  assign n185 = ~n9537 & ~n179;
  assign n186 = n184 & n185;
  assign n187 = n171 & n180;
  assign n188 = n165 & n172;
  assign n189 = n9532 & n176;
  assign n190 = n188 & n189;
  assign n191 = n166 & n173;
  assign n192 = n189 & n191;
  assign n193 = n155 & n9536;
  assign n194 = n172 & n193;
  assign n195 = n177 & n194;
  assign n196 = ~n192 & ~n195;
  assign n197 = ~n190 & n196;
  assign n198 = ~n9532 & n141;
  assign n199 = n174 & n198;
  assign n200 = n125 & n9534;
  assign n201 = n9532 & n200;
  assign n202 = n167 & n201;
  assign n203 = ~n199 & ~n202;
  assign n204 = n162 & n166;
  assign n205 = n201 & n204;
  assign n206 = n203 & ~n205;
  assign n207 = n197 & n206;
  assign n208 = n9538 & n206;
  assign n209 = n197 & n208;
  assign n210 = n9538 & n207;
  assign n211 = ~n125 & ~n9534;
  assign n212 = ~n9532 & n211;
  assign n213 = ~n146 & n149;
  assign n214 = n162 & n213;
  assign n215 = n212 & n214;
  assign n216 = n162 & n172;
  assign n217 = n198 & n216;
  assign n218 = n166 & n193;
  assign n219 = n198 & n218;
  assign n220 = ~n217 & ~n219;
  assign n221 = ~n215 & ~n219;
  assign n222 = ~n217 & n221;
  assign n223 = ~n215 & n220;
  assign n224 = n9532 & n211;
  assign n225 = n194 & n224;
  assign n226 = n177 & n191;
  assign n227 = ~n225 & ~n226;
  assign n228 = n167 & n198;
  assign n229 = ~n9532 & n168;
  assign n230 = n174 & n201;
  assign n231 = ~n9541 & ~n230;
  assign n232 = ~n225 & ~n230;
  assign n233 = ~n226 & ~n9541;
  assign n234 = n232 & n233;
  assign n235 = n227 & n231;
  assign n236 = n9540 & ~n225;
  assign n237 = ~n9541 & n236;
  assign n238 = ~n226 & n237;
  assign n239 = ~n230 & n238;
  assign n240 = n9540 & n9542;
  assign n241 = n163 & n198;
  assign n242 = n193 & n213;
  assign n243 = n189 & n242;
  assign n244 = ~n241 & ~n243;
  assign n245 = n141 & n242;
  assign n246 = n198 & n242;
  assign n247 = ~n9532 & n245;
  assign n248 = n173 & n213;
  assign n249 = n142 & n248;
  assign n250 = n194 & n201;
  assign n251 = ~n249 & ~n250;
  assign n252 = ~n9544 & ~n249;
  assign n253 = ~n250 & n252;
  assign n254 = ~n9544 & n251;
  assign n255 = ~n241 & n9545;
  assign n256 = ~n243 & n255;
  assign n257 = n244 & n9545;
  assign n258 = n189 & n194;
  assign n259 = ~n9532 & n200;
  assign n260 = n242 & n259;
  assign n261 = ~n258 & ~n260;
  assign n262 = n191 & n224;
  assign n263 = n150 & n193;
  assign n264 = n189 & n263;
  assign n265 = n177 & n216;
  assign n266 = ~n264 & ~n265;
  assign n267 = ~n262 & n266;
  assign n268 = ~n262 & ~n265;
  assign n269 = ~n258 & n268;
  assign n270 = ~n264 & n269;
  assign n271 = ~n260 & n270;
  assign n272 = ~n260 & ~n264;
  assign n273 = ~n258 & n272;
  assign n274 = n261 & ~n264;
  assign n275 = n268 & n9548;
  assign n276 = n261 & n267;
  assign n277 = n9546 & n9547;
  assign n278 = n9543 & n9547;
  assign n279 = n9546 & n278;
  assign n280 = n9543 & n9546;
  assign n281 = n9547 & n280;
  assign n282 = n9543 & n277;
  assign n283 = n9539 & n9549;
  assign n284 = n218 & n259;
  assign n285 = n141 & n178;
  assign n286 = n142 & n178;
  assign n287 = n9532 & n285;
  assign n288 = n178 & n198;
  assign n289 = ~n9532 & n285;
  assign n290 = ~n284 & ~n9551;
  assign n291 = ~n9550 & n290;
  assign n292 = ~n284 & ~n285;
  assign n293 = n165 & n213;
  assign n294 = n201 & n293;
  assign n295 = n142 & n214;
  assign n296 = n224 & n248;
  assign n297 = ~n295 & ~n296;
  assign n298 = ~n294 & n297;
  assign n299 = n9552 & n298;
  assign n300 = n167 & n259;
  assign n301 = n167 & n177;
  assign n302 = n191 & n200;
  assign n303 = n191 & n259;
  assign n304 = ~n9532 & n302;
  assign n305 = ~n301 & ~n9553;
  assign n306 = ~n300 & ~n9553;
  assign n307 = ~n301 & n306;
  assign n308 = ~n300 & ~n301;
  assign n309 = ~n9553 & n308;
  assign n310 = ~n300 & n305;
  assign n311 = n191 & n212;
  assign n312 = n212 & n242;
  assign n313 = n211 & n218;
  assign n314 = n212 & n218;
  assign n315 = ~n9532 & n313;
  assign n316 = ~n312 & ~n9555;
  assign n317 = ~n311 & ~n9555;
  assign n318 = ~n312 & n317;
  assign n319 = ~n311 & ~n312;
  assign n320 = ~n9555 & n319;
  assign n321 = ~n311 & n316;
  assign n322 = n9554 & n9556;
  assign n323 = n299 & n322;
  assign n324 = n142 & n216;
  assign n325 = n174 & n224;
  assign n326 = ~n324 & ~n325;
  assign n327 = n174 & n212;
  assign n328 = n142 & n218;
  assign n329 = ~n327 & ~n328;
  assign n330 = n326 & n329;
  assign n331 = n201 & n218;
  assign n332 = n177 & n263;
  assign n333 = ~n331 & ~n332;
  assign n334 = n178 & n212;
  assign n335 = n177 & n188;
  assign n336 = ~n334 & ~n335;
  assign n337 = n333 & n336;
  assign n338 = n326 & ~n334;
  assign n339 = ~n327 & n338;
  assign n340 = ~n328 & n339;
  assign n341 = ~n335 & n340;
  assign n342 = ~n332 & n341;
  assign n343 = ~n331 & n342;
  assign n344 = ~n328 & ~n335;
  assign n345 = ~n327 & ~n334;
  assign n346 = n329 & n336;
  assign n347 = n344 & n345;
  assign n348 = n326 & n333;
  assign n349 = n9558 & n348;
  assign n350 = n330 & n337;
  assign n351 = n259 & n293;
  assign n352 = n201 & n214;
  assign n353 = ~n351 & ~n352;
  assign n354 = n163 & n211;
  assign n355 = n191 & n201;
  assign n356 = n9532 & n302;
  assign n357 = ~n354 & ~n9559;
  assign n358 = n353 & ~n9559;
  assign n359 = ~n354 & n358;
  assign n360 = n163 & n212;
  assign n361 = ~n9532 & n354;
  assign n362 = n163 & n224;
  assign n363 = n9532 & n354;
  assign n364 = n353 & ~n9562;
  assign n365 = ~n9561 & n364;
  assign n366 = ~n9559 & n365;
  assign n367 = n353 & n357;
  assign n368 = n9557 & n9560;
  assign n369 = n9552 & n322;
  assign n370 = n9560 & n369;
  assign n371 = n9557 & n370;
  assign n372 = ~n296 & n371;
  assign n373 = ~n295 & n372;
  assign n374 = ~n294 & n373;
  assign n375 = n9554 & n9560;
  assign n376 = n9556 & n375;
  assign n377 = n299 & n9557;
  assign n378 = n376 & n377;
  assign n379 = n323 & n368;
  assign n380 = n177 & n248;
  assign n381 = n163 & n189;
  assign n382 = ~n380 & ~n381;
  assign n383 = n212 & n248;
  assign n384 = n204 & n259;
  assign n385 = ~n383 & ~n384;
  assign n386 = n224 & n242;
  assign n387 = n218 & n224;
  assign n388 = n9532 & n313;
  assign n389 = ~n386 & ~n9564;
  assign n390 = n385 & n389;
  assign n391 = n382 & n389;
  assign n392 = n385 & n391;
  assign n393 = n382 & n390;
  assign n394 = n198 & n248;
  assign n395 = n204 & n211;
  assign n396 = ~n394 & ~n395;
  assign n397 = n189 & n248;
  assign n398 = n214 & n259;
  assign n399 = ~n397 & ~n398;
  assign n400 = n396 & n399;
  assign n401 = n212 & n263;
  assign n402 = n178 & n224;
  assign n403 = ~n401 & ~n402;
  assign n404 = n214 & n224;
  assign n405 = n224 & n263;
  assign n406 = ~n404 & ~n405;
  assign n407 = n403 & n406;
  assign n408 = ~n395 & ~n398;
  assign n409 = ~n394 & ~n401;
  assign n410 = n408 & n409;
  assign n411 = ~n397 & ~n402;
  assign n412 = n406 & n411;
  assign n413 = n410 & n412;
  assign n414 = n204 & n224;
  assign n415 = n204 & n212;
  assign n416 = ~n401 & ~n415;
  assign n417 = ~n414 & n416;
  assign n418 = ~n394 & ~n398;
  assign n419 = n406 & n418;
  assign n420 = n411 & n419;
  assign n421 = n417 & n420;
  assign n422 = n400 & n407;
  assign n423 = n9565 & n411;
  assign n424 = n406 & n423;
  assign n425 = ~n414 & n424;
  assign n426 = ~n415 & n425;
  assign n427 = ~n401 & n426;
  assign n428 = ~n394 & n427;
  assign n429 = ~n398 & n428;
  assign n430 = n9565 & n9566;
  assign n431 = n189 & n216;
  assign n432 = n194 & n212;
  assign n433 = ~n431 & ~n432;
  assign n434 = n9567 & ~n432;
  assign n435 = ~n431 & n434;
  assign n436 = n9567 & n433;
  assign n437 = n9563 & n9568;
  assign n438 = n203 & n9568;
  assign n439 = n197 & n438;
  assign n440 = n9538 & n439;
  assign n441 = n9547 & n440;
  assign n442 = n9543 & n441;
  assign n443 = n9563 & n442;
  assign n444 = n9546 & n443;
  assign n445 = ~n205 & n444;
  assign n446 = n283 & n9563;
  assign n447 = n9568 & n446;
  assign n448 = n283 & n437;
  assign n449 = n142 & n242;
  assign n450 = n9532 & n245;
  assign n451 = ~n175 & ~n9570;
  assign n452 = ~n414 & ~n432;
  assign n453 = ~n295 & ~n381;
  assign n454 = n452 & n453;
  assign n455 = ~n295 & n452;
  assign n456 = ~n9570 & n455;
  assign n457 = ~n175 & n456;
  assign n458 = ~n381 & n457;
  assign n459 = n451 & n452;
  assign n460 = n453 & n459;
  assign n461 = ~n175 & ~n381;
  assign n462 = ~n295 & ~n9570;
  assign n463 = n461 & n462;
  assign n464 = n452 & n463;
  assign n465 = n451 & n454;
  assign n466 = ~n226 & ~n397;
  assign n467 = n142 & n194;
  assign n468 = n167 & n224;
  assign n469 = ~n467 & ~n468;
  assign n470 = n201 & n263;
  assign n471 = ~n205 & ~n470;
  assign n472 = n469 & n471;
  assign n473 = n466 & n471;
  assign n474 = n469 & n473;
  assign n475 = n466 & n472;
  assign n476 = n178 & n201;
  assign n477 = ~n195 & ~n398;
  assign n478 = ~n476 & n477;
  assign n479 = n163 & n259;
  assign n480 = n216 & n259;
  assign n481 = ~n324 & ~n480;
  assign n482 = ~n324 & ~n479;
  assign n483 = ~n480 & n482;
  assign n484 = ~n479 & n481;
  assign n485 = n478 & n9573;
  assign n486 = ~n226 & ~n476;
  assign n487 = ~n205 & ~n397;
  assign n488 = n486 & n487;
  assign n489 = n477 & n488;
  assign n490 = n469 & ~n470;
  assign n491 = n9573 & n490;
  assign n492 = n489 & n491;
  assign n493 = ~n397 & ~n468;
  assign n494 = n477 & n493;
  assign n495 = n486 & n494;
  assign n496 = ~n467 & ~n470;
  assign n497 = ~n205 & n496;
  assign n498 = n9573 & n497;
  assign n499 = n495 & n498;
  assign n500 = n9572 & n485;
  assign n501 = n9573 & n486;
  assign n502 = n9571 & n501;
  assign n503 = n477 & n502;
  assign n504 = ~n468 & n503;
  assign n505 = ~n467 & n504;
  assign n506 = ~n397 & n505;
  assign n507 = ~n205 & n506;
  assign n508 = ~n470 & n507;
  assign n509 = n9571 & n9574;
  assign n510 = ~n225 & ~n250;
  assign n511 = n248 & n259;
  assign n512 = ~n264 & ~n511;
  assign n513 = n189 & n214;
  assign n514 = n150 & n165;
  assign n515 = n177 & n514;
  assign n516 = ~n513 & ~n515;
  assign n517 = n512 & n516;
  assign n518 = ~n225 & ~n515;
  assign n519 = ~n264 & n518;
  assign n520 = ~n513 & n519;
  assign n521 = ~n250 & n520;
  assign n522 = ~n511 & n521;
  assign n523 = ~n250 & ~n264;
  assign n524 = ~n511 & ~n513;
  assign n525 = n518 & n524;
  assign n526 = n523 & n525;
  assign n527 = ~n225 & ~n511;
  assign n528 = ~n250 & ~n515;
  assign n529 = ~n264 & ~n513;
  assign n530 = n528 & n529;
  assign n531 = n527 & n530;
  assign n532 = n510 & n517;
  assign n533 = n174 & n177;
  assign n534 = n177 & n293;
  assign n535 = ~n533 & ~n534;
  assign n536 = n201 & n248;
  assign n537 = ~n351 & ~n536;
  assign n538 = n177 & n204;
  assign n539 = ~n405 & ~n538;
  assign n540 = ~n536 & ~n538;
  assign n541 = ~n351 & ~n405;
  assign n542 = n540 & n541;
  assign n543 = n537 & n539;
  assign n544 = ~n405 & ~n536;
  assign n545 = ~n351 & ~n534;
  assign n546 = ~n533 & ~n538;
  assign n547 = n545 & n546;
  assign n548 = n544 & n547;
  assign n549 = n535 & n9577;
  assign n550 = ~n217 & ~n241;
  assign n551 = ~n335 & n550;
  assign n552 = n259 & n514;
  assign n553 = ~n219 & ~n552;
  assign n554 = n198 & n263;
  assign n555 = ~n243 & ~n554;
  assign n556 = ~n219 & ~n554;
  assign n557 = ~n243 & n556;
  assign n558 = ~n552 & n557;
  assign n559 = ~n243 & ~n552;
  assign n560 = n556 & n559;
  assign n561 = n553 & n555;
  assign n562 = n551 & n9579;
  assign n563 = n9578 & n562;
  assign n564 = n9576 & n551;
  assign n565 = n9579 & n564;
  assign n566 = ~n405 & n565;
  assign n567 = ~n538 & n566;
  assign n568 = ~n533 & n567;
  assign n569 = ~n534 & n568;
  assign n570 = ~n536 & n569;
  assign n571 = ~n351 & n570;
  assign n572 = n9576 & n563;
  assign n573 = n142 & n514;
  assign n574 = n198 & n293;
  assign n575 = ~n9551 & ~n574;
  assign n576 = ~n573 & ~n574;
  assign n577 = ~n9551 & n576;
  assign n578 = ~n9551 & ~n573;
  assign n579 = ~n574 & n578;
  assign n580 = ~n573 & n575;
  assign n581 = n188 & n212;
  assign n582 = n177 & n214;
  assign n583 = n212 & n216;
  assign n584 = ~n582 & ~n583;
  assign n585 = ~n581 & ~n583;
  assign n586 = ~n582 & n585;
  assign n587 = ~n581 & ~n582;
  assign n588 = ~n583 & n587;
  assign n589 = ~n581 & n584;
  assign n590 = ~n249 & ~n394;
  assign n591 = n141 & n248;
  assign n592 = n216 & n224;
  assign n593 = n9583 & ~n592;
  assign n594 = ~n300 & n9583;
  assign n595 = ~n592 & n594;
  assign n596 = ~n300 & ~n592;
  assign n597 = n9583 & n596;
  assign n598 = ~n300 & n593;
  assign n599 = n9582 & n9584;
  assign n600 = n9581 & n9584;
  assign n601 = n9582 & n600;
  assign n602 = n9581 & n599;
  assign n603 = ~n331 & ~n415;
  assign n604 = n198 & n204;
  assign n605 = n167 & n189;
  assign n606 = ~n604 & ~n605;
  assign n607 = n176 & n218;
  assign n608 = n177 & n218;
  assign n609 = ~n9532 & n607;
  assign n610 = ~n9553 & ~n9586;
  assign n611 = n606 & n610;
  assign n612 = ~n415 & ~n604;
  assign n613 = ~n9586 & n612;
  assign n614 = ~n605 & n613;
  assign n615 = ~n331 & n614;
  assign n616 = ~n9553 & n615;
  assign n617 = n603 & n611;
  assign n618 = n201 & n242;
  assign n619 = ~n431 & ~n618;
  assign n620 = n178 & n189;
  assign n621 = ~n230 & ~n620;
  assign n622 = n619 & n621;
  assign n623 = n188 & n259;
  assign n624 = n224 & n514;
  assign n625 = ~n623 & ~n624;
  assign n626 = n188 & n224;
  assign n627 = n167 & n212;
  assign n628 = ~n626 & ~n627;
  assign n629 = n625 & n628;
  assign n630 = ~n624 & ~n626;
  assign n631 = ~n627 & n630;
  assign n632 = ~n431 & n631;
  assign n633 = ~n620 & n632;
  assign n634 = ~n230 & n633;
  assign n635 = ~n618 & n634;
  assign n636 = ~n623 & n635;
  assign n637 = n621 & n628;
  assign n638 = n619 & n625;
  assign n639 = n637 & n638;
  assign n640 = ~n230 & ~n626;
  assign n641 = n619 & n640;
  assign n642 = ~n620 & ~n627;
  assign n643 = n625 & n642;
  assign n644 = n641 & n643;
  assign n645 = n622 & n629;
  assign n646 = n9587 & n9588;
  assign n647 = n9585 & n646;
  assign n648 = n9580 & n647;
  assign n649 = n9581 & n9582;
  assign n650 = n9587 & n649;
  assign n651 = n9575 & n650;
  assign n652 = n9580 & n651;
  assign n653 = n9588 & n652;
  assign n654 = ~n592 & n653;
  assign n655 = ~n249 & n654;
  assign n656 = ~n394 & n655;
  assign n657 = ~n300 & n656;
  assign n658 = n9575 & n648;
  assign n659 = ~n190 & ~n511;
  assign n660 = ~n9555 & ~n384;
  assign n661 = n659 & n660;
  assign n662 = ~n164 & ~n295;
  assign n663 = n212 & n293;
  assign n664 = ~n583 & ~n663;
  assign n665 = n662 & n664;
  assign n666 = n659 & n664;
  assign n667 = ~n9555 & n666;
  assign n668 = ~n295 & n667;
  assign n669 = ~n164 & n668;
  assign n670 = ~n384 & n669;
  assign n671 = n660 & n662;
  assign n672 = n666 & n671;
  assign n673 = n661 & n665;
  assign n674 = n163 & n201;
  assign n675 = ~n241 & ~n674;
  assign n676 = n189 & n204;
  assign n677 = ~n592 & ~n676;
  assign n678 = ~n241 & ~n592;
  assign n679 = ~n674 & ~n676;
  assign n680 = n678 & n679;
  assign n681 = n675 & n677;
  assign n682 = n212 & n514;
  assign n683 = ~n383 & ~n682;
  assign n684 = n389 & n683;
  assign n685 = ~n243 & ~n538;
  assign n686 = ~n296 & ~n468;
  assign n687 = n685 & n686;
  assign n688 = n389 & n686;
  assign n689 = n683 & n685;
  assign n690 = n688 & n689;
  assign n691 = n684 & n687;
  assign n692 = n9591 & n9592;
  assign n693 = n684 & n685;
  assign n694 = n9590 & n693;
  assign n695 = ~n592 & n694;
  assign n696 = ~n468 & n695;
  assign n697 = ~n296 & n696;
  assign n698 = ~n241 & n697;
  assign n699 = ~n676 & n698;
  assign n700 = ~n674 & n699;
  assign n701 = n9590 & n692;
  assign n702 = ~n250 & ~n311;
  assign n703 = ~n311 & n9593;
  assign n704 = ~n250 & n703;
  assign n705 = n9593 & n702;
  assign n706 = ~n394 & ~n536;
  assign n707 = ~n9570 & ~n605;
  assign n708 = ~n9550 & ~n627;
  assign n709 = ~n605 & ~n627;
  assign n710 = ~n9550 & ~n9570;
  assign n711 = n709 & n710;
  assign n712 = n707 & n708;
  assign n713 = n706 & n9595;
  assign n714 = n224 & n293;
  assign n715 = n142 & n293;
  assign n716 = ~n312 & ~n715;
  assign n717 = ~n312 & ~n714;
  assign n718 = ~n715 & n717;
  assign n719 = ~n714 & n716;
  assign n720 = n174 & n189;
  assign n721 = ~n334 & ~n720;
  assign n722 = ~n230 & ~n720;
  assign n723 = ~n334 & n722;
  assign n724 = ~n230 & n721;
  assign n725 = n9596 & n9597;
  assign n726 = ~n226 & ~n401;
  assign n727 = ~n325 & ~n401;
  assign n728 = ~n226 & n727;
  assign n729 = ~n325 & n726;
  assign n730 = n259 & n263;
  assign n731 = ~n192 & ~n730;
  assign n732 = ~n199 & ~n332;
  assign n733 = ~n192 & n732;
  assign n734 = ~n730 & n733;
  assign n735 = ~n332 & ~n730;
  assign n736 = ~n192 & ~n199;
  assign n737 = n735 & n736;
  assign n738 = n731 & n732;
  assign n739 = n9598 & n9599;
  assign n740 = n9597 & n9598;
  assign n741 = n9596 & n740;
  assign n742 = n9599 & n741;
  assign n743 = n9596 & n9599;
  assign n744 = n740 & n743;
  assign n745 = n725 & n739;
  assign n746 = ~n627 & n9600;
  assign n747 = ~n9570 & n746;
  assign n748 = ~n9550 & n747;
  assign n749 = ~n394 & n748;
  assign n750 = ~n605 & n749;
  assign n751 = ~n536 & n750;
  assign n752 = n713 & n9600;
  assign n753 = ~n479 & ~n574;
  assign n754 = n201 & n514;
  assign n755 = ~n618 & ~n754;
  assign n756 = n753 & n755;
  assign n757 = n198 & n514;
  assign n758 = ~n202 & ~n757;
  assign n759 = n382 & n758;
  assign n760 = n753 & n758;
  assign n761 = n382 & n760;
  assign n762 = ~n754 & n761;
  assign n763 = ~n618 & n762;
  assign n764 = n382 & n755;
  assign n765 = n760 & n764;
  assign n766 = n756 & n759;
  assign n767 = ~n533 & n9602;
  assign n768 = ~n534 & n767;
  assign n769 = n535 & n9602;
  assign n770 = n189 & n293;
  assign n771 = ~n265 & ~n770;
  assign n772 = n142 & n263;
  assign n773 = ~n9551 & ~n772;
  assign n774 = n771 & n773;
  assign n775 = ~n327 & ~n554;
  assign n776 = n194 & n198;
  assign n777 = ~n402 & ~n776;
  assign n778 = n775 & n777;
  assign n779 = n774 & n778;
  assign n780 = ~n249 & ~n620;
  assign n781 = n178 & n259;
  assign n782 = ~n300 & ~n781;
  assign n783 = ~n300 & n780;
  assign n784 = ~n781 & n783;
  assign n785 = n780 & n782;
  assign n786 = ~n284 & ~n335;
  assign n787 = ~n262 & ~n552;
  assign n788 = n786 & n787;
  assign n789 = n9604 & n788;
  assign n790 = n268 & n773;
  assign n791 = n268 & n775;
  assign n792 = n773 & n777;
  assign n793 = n791 & n792;
  assign n794 = n773 & n775;
  assign n795 = n268 & n777;
  assign n796 = n794 & n795;
  assign n797 = n778 & n790;
  assign n798 = ~n552 & ~n770;
  assign n799 = ~n335 & ~n552;
  assign n800 = ~n284 & ~n770;
  assign n801 = n799 & n800;
  assign n802 = n786 & n798;
  assign n803 = n9604 & n9606;
  assign n804 = n9605 & n803;
  assign n805 = n779 & n789;
  assign n806 = n9603 & n9607;
  assign n807 = n9601 & n806;
  assign n808 = n9594 & n9603;
  assign n809 = n777 & n808;
  assign n810 = n775 & n809;
  assign n811 = n773 & n810;
  assign n812 = n9601 & n811;
  assign n813 = n9604 & n812;
  assign n814 = ~n335 & n813;
  assign n815 = n268 & n814;
  assign n816 = ~n770 & n815;
  assign n817 = ~n552 & n816;
  assign n818 = ~n284 & n817;
  assign n819 = n9594 & n807;
  assign n820 = ~n9589 & ~n9608;
  assign n821 = ~n9569 & ~n820;
  assign n822 = ~n9551 & ~n627;
  assign n823 = ~n312 & ~n627;
  assign n824 = ~n9551 & n823;
  assign n825 = ~n312 & n822;
  assign n826 = ~n199 & ~n468;
  assign n827 = n389 & n826;
  assign n828 = ~n312 & n827;
  assign n829 = ~n627 & n828;
  assign n830 = ~n9551 & n829;
  assign n831 = ~n312 & n826;
  assign n832 = n389 & n822;
  assign n833 = n831 & n832;
  assign n834 = ~n312 & n389;
  assign n835 = n822 & n826;
  assign n836 = n834 & n835;
  assign n837 = n9609 & n827;
  assign n838 = ~n175 & ~n9550;
  assign n839 = ~n9550 & n9610;
  assign n840 = ~n175 & n839;
  assign n841 = n9610 & n838;
  assign n842 = ~n467 & ~n776;
  assign n843 = ~n415 & ~n467;
  assign n844 = ~n776 & n843;
  assign n845 = ~n415 & n842;
  assign n846 = ~n215 & ~n772;
  assign n847 = ~n414 & ~n592;
  assign n848 = ~n215 & n847;
  assign n849 = ~n772 & n848;
  assign n850 = ~n414 & ~n772;
  assign n851 = ~n215 & ~n592;
  assign n852 = n850 & n851;
  assign n853 = ~n215 & ~n414;
  assign n854 = ~n592 & ~n772;
  assign n855 = n853 & n854;
  assign n856 = n846 & n847;
  assign n857 = ~n554 & ~n583;
  assign n858 = n9613 & n857;
  assign n859 = n9612 & n9613;
  assign n860 = ~n583 & n859;
  assign n861 = ~n554 & n860;
  assign n862 = n9612 & n857;
  assign n863 = n9613 & n862;
  assign n864 = n9612 & n858;
  assign n865 = ~n296 & ~n624;
  assign n866 = ~n334 & ~n581;
  assign n867 = ~n581 & ~n624;
  assign n868 = ~n296 & ~n334;
  assign n869 = n867 & n868;
  assign n870 = n865 & n866;
  assign n871 = n191 & n198;
  assign n872 = ~n626 & ~n871;
  assign n873 = n403 & n872;
  assign n874 = ~n334 & ~n401;
  assign n875 = ~n296 & ~n402;
  assign n876 = n874 & n875;
  assign n877 = n867 & n872;
  assign n878 = n876 & n877;
  assign n879 = ~n334 & ~n402;
  assign n880 = n867 & n879;
  assign n881 = ~n296 & ~n401;
  assign n882 = n872 & n881;
  assign n883 = n880 & n882;
  assign n884 = n9615 & n873;
  assign n885 = n9614 & n9616;
  assign n886 = n9611 & n872;
  assign n887 = n9614 & n886;
  assign n888 = ~n624 & n887;
  assign n889 = ~n402 & n888;
  assign n890 = ~n296 & n889;
  assign n891 = ~n334 & n890;
  assign n892 = ~n581 & n891;
  assign n893 = ~n401 & n892;
  assign n894 = n9611 & n9616;
  assign n895 = n9614 & n894;
  assign n896 = n9611 & n885;
  assign n897 = n142 & n204;
  assign n898 = n198 & n214;
  assign n899 = ~n897 & ~n898;
  assign n900 = ~n9562 & ~n404;
  assign n901 = n899 & n900;
  assign n902 = ~n245 & ~n432;
  assign n903 = ~n219 & ~n405;
  assign n904 = ~n245 & ~n405;
  assign n905 = ~n219 & ~n432;
  assign n906 = n904 & n905;
  assign n907 = n902 & n903;
  assign n908 = ~n225 & ~n328;
  assign n909 = ~n9561 & ~n604;
  assign n910 = n908 & n909;
  assign n911 = n9618 & n910;
  assign n912 = n406 & n899;
  assign n913 = n899 & n908;
  assign n914 = n909 & n913;
  assign n915 = n406 & n914;
  assign n916 = n910 & n912;
  assign n917 = ~n9562 & n9619;
  assign n918 = ~n432 & n917;
  assign n919 = ~n245 & n918;
  assign n920 = ~n219 & n919;
  assign n921 = ~n219 & ~n245;
  assign n922 = ~n9562 & ~n432;
  assign n923 = n921 & n922;
  assign n924 = n9619 & n923;
  assign n925 = ~n245 & n908;
  assign n926 = n899 & n925;
  assign n927 = ~n219 & ~n9562;
  assign n928 = ~n432 & n927;
  assign n929 = n406 & n909;
  assign n930 = n928 & n929;
  assign n931 = n926 & n930;
  assign n932 = n901 & n911;
  assign n933 = n142 & n191;
  assign n934 = ~n9555 & ~n933;
  assign n935 = ~n327 & n9583;
  assign n936 = ~n325 & n9583;
  assign n937 = ~n327 & n936;
  assign n938 = ~n325 & n935;
  assign n939 = ~n9555 & ~n325;
  assign n940 = ~n327 & n939;
  assign n941 = ~n933 & n940;
  assign n942 = ~n249 & n941;
  assign n943 = ~n394 & n942;
  assign n944 = ~n327 & ~n394;
  assign n945 = ~n249 & ~n325;
  assign n946 = n934 & n945;
  assign n947 = n944 & n946;
  assign n948 = n934 & n9621;
  assign n949 = ~n191 & ~n293;
  assign n950 = ~n262 & ~n663;
  assign n951 = ~n311 & ~n714;
  assign n952 = n950 & n951;
  assign n953 = n211 & ~n949;
  assign n954 = n683 & n9623;
  assign n955 = n9622 & n954;
  assign n956 = n9620 & n955;
  assign n957 = n683 & n9622;
  assign n958 = n9617 & n957;
  assign n959 = n9620 & n958;
  assign n960 = ~n714 & n959;
  assign n961 = ~n262 & n960;
  assign n962 = ~n663 & n961;
  assign n963 = ~n311 & n962;
  assign n964 = n9617 & n956;
  assign n965 = ~pi22  & ~n94;
  assign n966 = pi9  & ~n965;
  assign n967 = ~pi9  & n965;
  assign n968 = ~pi9  & ~n965;
  assign n969 = pi9  & n965;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~n966 & ~n967;
  assign n972 = ~n9624 & n9625;
  assign n973 = ~n821 & n972;
  assign n974 = pi10  & pi22 ;
  assign n975 = ~pi22  & ~n96;
  assign n976 = pi10  & ~n95;
  assign n977 = n975 & ~n976;
  assign n978 = ~n974 & ~n977;
  assign n979 = ~n9624 & ~n978;
  assign n980 = n821 & ~n972;
  assign n981 = ~n973 & ~n980;
  assign n982 = n979 & n981;
  assign n983 = ~n973 & ~n982;
  assign n984 = pi11  & ~n975;
  assign n985 = ~pi11  & n975;
  assign n986 = ~pi11  & ~n975;
  assign n987 = pi11  & n975;
  assign n988 = ~n986 & ~n987;
  assign n989 = ~n984 & ~n985;
  assign n990 = n142 & n188;
  assign n991 = ~n574 & ~n757;
  assign n992 = ~n990 & n991;
  assign n993 = ~n9541 & ~n715;
  assign n994 = ~n192 & ~n295;
  assign n995 = n188 & n198;
  assign n996 = ~n720 & ~n995;
  assign n997 = n994 & n996;
  assign n998 = n993 & n996;
  assign n999 = n994 & n998;
  assign n1000 = n993 & n997;
  assign n1001 = ~n720 & ~n990;
  assign n1002 = ~n995 & n1001;
  assign n1003 = n991 & n994;
  assign n1004 = n993 & n994;
  assign n1005 = n991 & n1004;
  assign n1006 = n993 & n1003;
  assign n1007 = n1002 & n9628;
  assign n1008 = n992 & n9627;
  assign n1009 = ~n179 & ~n533;
  assign n1010 = ~n620 & n1009;
  assign n1011 = ~n380 & ~n607;
  assign n1012 = ~n607 & n1010;
  assign n1013 = ~n380 & n1012;
  assign n1014 = n1010 & n1011;
  assign n1015 = n177 & n242;
  assign n1016 = ~n9537 & ~n573;
  assign n1017 = ~n573 & ~n1015;
  assign n1018 = ~n9537 & n1017;
  assign n1019 = ~n1015 & n1016;
  assign n1020 = ~n226 & n9631;
  assign n1021 = ~n397 & n1020;
  assign n1022 = ~n9537 & ~n226;
  assign n1023 = ~n397 & ~n573;
  assign n1024 = ~n1015 & n1023;
  assign n1025 = n1022 & n1024;
  assign n1026 = ~n1015 & n1022;
  assign n1027 = n1023 & n1026;
  assign n1028 = n466 & n9631;
  assign n1029 = n9630 & n9632;
  assign n1030 = n9628 & n9632;
  assign n1031 = n9630 & n1030;
  assign n1032 = ~n990 & n1031;
  assign n1033 = ~n995 & n1032;
  assign n1034 = ~n720 & n1033;
  assign n1035 = n9629 & n1029;
  assign n1036 = ~n164 & ~n324;
  assign n1037 = n174 & n259;
  assign n1038 = ~n781 & ~n1037;
  assign n1039 = n1036 & n1038;
  assign n1040 = n659 & n1038;
  assign n1041 = n1036 & n1040;
  assign n1042 = n659 & n1036;
  assign n1043 = n1038 & n1042;
  assign n1044 = n659 & n1039;
  assign n1045 = ~n302 & ~n536;
  assign n1046 = ~n9559 & ~n536;
  assign n1047 = ~n9553 & ~n476;
  assign n1048 = n1046 & n1047;
  assign n1049 = ~n476 & n1045;
  assign n1050 = n551 & n9635;
  assign n1051 = n551 & n1038;
  assign n1052 = n659 & n1051;
  assign n1053 = n1036 & n1052;
  assign n1054 = ~n536 & n1053;
  assign n1055 = ~n9559 & n1054;
  assign n1056 = ~n476 & n1055;
  assign n1057 = ~n9553 & n1056;
  assign n1058 = n9634 & n1050;
  assign n1059 = ~n284 & ~n331;
  assign n1060 = ~n230 & ~n260;
  assign n1061 = ~n230 & ~n331;
  assign n1062 = ~n260 & ~n284;
  assign n1063 = n1061 & n1062;
  assign n1064 = n1059 & n1060;
  assign n1065 = ~n230 & n9636;
  assign n1066 = ~n331 & n1065;
  assign n1067 = ~n284 & n1066;
  assign n1068 = ~n260 & n1067;
  assign n1069 = n9636 & n9637;
  assign n1070 = n194 & n259;
  assign n1071 = ~n470 & ~n1070;
  assign n1072 = ~n618 & ~n730;
  assign n1073 = n1071 & n1072;
  assign n1074 = n9638 & n1073;
  assign n1075 = n9638 & ~n1070;
  assign n1076 = n9633 & n1075;
  assign n1077 = ~n618 & n1076;
  assign n1078 = ~n470 & n1077;
  assign n1079 = ~n730 & n1078;
  assign n1080 = n9633 & n1073;
  assign n1081 = n9638 & n1080;
  assign n1082 = n9633 & n1074;
  assign n1083 = n163 & n177;
  assign n1084 = ~n676 & ~n1083;
  assign n1085 = ~n513 & ~n676;
  assign n1086 = ~n1083 & n1085;
  assign n1087 = ~n513 & n1084;
  assign n1088 = ~n195 & ~n582;
  assign n1089 = ~n195 & ~n264;
  assign n1090 = ~n582 & n1089;
  assign n1091 = ~n264 & n1088;
  assign n1092 = ~n258 & ~n332;
  assign n1093 = n685 & n1092;
  assign n1094 = n9641 & n1093;
  assign n1095 = n685 & n9640;
  assign n1096 = ~n582 & n1095;
  assign n1097 = ~n195 & n1096;
  assign n1098 = ~n332 & n1097;
  assign n1099 = ~n258 & n1098;
  assign n1100 = ~n264 & n1099;
  assign n1101 = n9640 & n1094;
  assign n1102 = n550 & n1036;
  assign n1103 = n9642 & n1102;
  assign n1104 = n9633 & n9642;
  assign n1105 = n550 & n1104;
  assign n1106 = n1036 & n1105;
  assign n1107 = n9633 & n1103;
  assign n1108 = n189 & n514;
  assign n1109 = ~n605 & ~n1108;
  assign n1110 = ~n515 & n1109;
  assign n1111 = ~n265 & ~n1108;
  assign n1112 = ~n515 & n1111;
  assign n1113 = ~n770 & n1112;
  assign n1114 = ~n605 & n1113;
  assign n1115 = ~n515 & ~n770;
  assign n1116 = ~n265 & n1115;
  assign n1117 = n1109 & n1116;
  assign n1118 = ~n605 & ~n770;
  assign n1119 = ~n515 & ~n605;
  assign n1120 = ~n770 & n1119;
  assign n1121 = ~n515 & n1118;
  assign n1122 = n1111 & n9645;
  assign n1123 = n771 & n1110;
  assign n1124 = ~n301 & ~n431;
  assign n1125 = ~n301 & ~n534;
  assign n1126 = ~n431 & n1125;
  assign n1127 = ~n534 & n1124;
  assign n1128 = ~n301 & n9644;
  assign n1129 = ~n534 & n1128;
  assign n1130 = ~n431 & n1129;
  assign n1131 = n9644 & n9646;
  assign n1132 = ~n381 & n9647;
  assign n1133 = n9643 & n9647;
  assign n1134 = ~n381 & n1133;
  assign n1135 = n9643 & n1132;
  assign n1136 = ~n9639 & ~n9648;
  assign n1137 = n9639 & n9648;
  assign n1138 = n9639 & ~n9648;
  assign n1139 = ~n9639 & n9648;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = ~n1136 & ~n1137;
  assign n1142 = n9624 & n9649;
  assign n1143 = ~n9626 & n1142;
  assign n1144 = n9626 & n1137;
  assign n1145 = pi12  & pi22 ;
  assign n1146 = ~pi22  & ~n98;
  assign n1147 = pi12  & ~n97;
  assign n1148 = n1146 & ~n1147;
  assign n1149 = ~n1145 & ~n1148;
  assign n1150 = ~n9624 & ~n1149;
  assign n1151 = n9624 & n1149;
  assign n1152 = ~n1150 & ~n1151;
  assign n1153 = ~n9649 & n1149;
  assign n1154 = ~n9649 & ~n1152;
  assign n1155 = ~n1144 & ~n9650;
  assign n1156 = ~n1143 & ~n1144;
  assign n1157 = ~n9650 & n1156;
  assign n1158 = ~n1143 & n1155;
  assign n1159 = pi14  & pi22 ;
  assign n1160 = pi14  & ~n99;
  assign n1161 = ~n100 & ~n1160;
  assign n1162 = ~pi22  & n1161;
  assign n1163 = n101 & ~n1160;
  assign n1164 = ~n1159 & ~n9652;
  assign n1165 = ~n215 & ~n401;
  assign n1166 = ~n335 & ~n352;
  assign n1167 = ~n335 & ~n401;
  assign n1168 = ~n215 & ~n352;
  assign n1169 = n1167 & n1168;
  assign n1170 = n1165 & n1166;
  assign n1171 = ~n195 & ~n513;
  assign n1172 = ~n480 & ~n536;
  assign n1173 = n406 & n1172;
  assign n1174 = n406 & n1171;
  assign n1175 = n1172 & n1174;
  assign n1176 = n1171 & n1173;
  assign n1177 = ~n215 & n1173;
  assign n1178 = ~n401 & n1177;
  assign n1179 = ~n335 & n1178;
  assign n1180 = ~n195 & n1179;
  assign n1181 = ~n513 & n1180;
  assign n1182 = ~n352 & n1181;
  assign n1183 = ~n195 & ~n215;
  assign n1184 = ~n352 & ~n513;
  assign n1185 = n1183 & n1184;
  assign n1186 = n406 & n1167;
  assign n1187 = n1172 & n1186;
  assign n1188 = n1185 & n1187;
  assign n1189 = n9653 & n9654;
  assign n1190 = n201 & n216;
  assign n1191 = ~n479 & ~n1190;
  assign n1192 = ~n9537 & ~n1037;
  assign n1193 = ~n217 & ~n995;
  assign n1194 = n1192 & n1193;
  assign n1195 = ~n217 & ~n479;
  assign n1196 = ~n995 & ~n1190;
  assign n1197 = n1195 & n1196;
  assign n1198 = n1192 & n1197;
  assign n1199 = n1191 & n1194;
  assign n1200 = ~n225 & ~n258;
  assign n1201 = ~n225 & ~n624;
  assign n1202 = ~n258 & n1201;
  assign n1203 = ~n258 & ~n624;
  assign n1204 = ~n225 & n1203;
  assign n1205 = ~n624 & n1200;
  assign n1206 = ~n9562 & ~n581;
  assign n1207 = ~n332 & ~n415;
  assign n1208 = ~n415 & n1206;
  assign n1209 = ~n332 & n1208;
  assign n1210 = n1206 & n1207;
  assign n1211 = n9657 & n9658;
  assign n1212 = n9656 & n1211;
  assign n1213 = n9655 & n1212;
  assign n1214 = n9594 & n9658;
  assign n1215 = n1192 & n1214;
  assign n1216 = n9657 & n1215;
  assign n1217 = n9655 & n1216;
  assign n1218 = ~n217 & n1217;
  assign n1219 = ~n995 & n1218;
  assign n1220 = ~n1190 & n1219;
  assign n1221 = ~n479 & n1220;
  assign n1222 = n9594 & n1213;
  assign n1223 = ~n573 & ~n871;
  assign n1224 = ~n9561 & ~n402;
  assign n1225 = ~n9553 & ~n398;
  assign n1226 = ~n398 & ~n402;
  assign n1227 = ~n9553 & ~n9561;
  assign n1228 = n1226 & n1227;
  assign n1229 = n1224 & n1225;
  assign n1230 = n1223 & n9660;
  assign n1231 = n9596 & n1223;
  assign n1232 = ~n402 & n1231;
  assign n1233 = ~n9561 & n1232;
  assign n1234 = ~n9553 & n1233;
  assign n1235 = ~n398 & n1234;
  assign n1236 = n9596 & n1230;
  assign n1237 = ~n627 & ~n757;
  assign n1238 = ~n627 & n9661;
  assign n1239 = ~n757 & n1238;
  assign n1240 = n9661 & n1237;
  assign n1241 = ~n327 & ~n574;
  assign n1242 = ~n262 & ~n582;
  assign n1243 = ~n262 & ~n327;
  assign n1244 = ~n574 & ~n582;
  assign n1245 = n1243 & n1244;
  assign n1246 = n1241 & n1242;
  assign n1247 = ~n626 & ~n933;
  assign n1248 = ~n264 & ~n334;
  assign n1249 = n1247 & n1248;
  assign n1250 = ~n262 & n1249;
  assign n1251 = ~n327 & n1250;
  assign n1252 = ~n574 & n1251;
  assign n1253 = ~n582 & n1252;
  assign n1254 = n9663 & n1249;
  assign n1255 = n452 & ~n781;
  assign n1256 = ~n205 & ~n9559;
  assign n1257 = n326 & n1256;
  assign n1258 = ~n9541 & ~n1083;
  assign n1259 = ~n476 & ~n990;
  assign n1260 = n1258 & n1259;
  assign n1261 = ~n9541 & ~n9559;
  assign n1262 = ~n205 & ~n1083;
  assign n1263 = n1261 & n1262;
  assign n1264 = n326 & n1259;
  assign n1265 = n1263 & n1264;
  assign n1266 = n1257 & n1260;
  assign n1267 = n1255 & n9665;
  assign n1268 = n9664 & n1267;
  assign n1269 = n9662 & n1268;
  assign n1270 = n326 & n9662;
  assign n1271 = n1255 & n1270;
  assign n1272 = n1259 & n1271;
  assign n1273 = n9664 & n1272;
  assign n1274 = n9659 & n1273;
  assign n1275 = n1258 & n1274;
  assign n1276 = ~n205 & n1275;
  assign n1277 = ~n9559 & n1276;
  assign n1278 = n9659 & n1269;
  assign n1279 = ~n9569 & ~n9666;
  assign n1280 = n9569 & n9666;
  assign n1281 = n9569 & ~n9666;
  assign n1282 = ~n9569 & n9666;
  assign n1283 = ~n1281 & ~n1282;
  assign n1284 = ~n1279 & ~n1280;
  assign n1285 = n9639 & ~n1280;
  assign n1286 = ~n9667 & ~n1285;
  assign n1287 = ~n9639 & ~n9667;
  assign n1288 = ~n1164 & n9668;
  assign n1289 = ~n9639 & ~n1279;
  assign n1290 = ~n9667 & ~n1289;
  assign n1291 = n9639 & ~n9667;
  assign n1292 = n1164 & n9669;
  assign n1293 = ~n1288 & ~n1292;
  assign n1294 = pi13  & ~n1146;
  assign n1295 = ~pi13  & n1146;
  assign n1296 = ~pi13  & ~n1146;
  assign n1297 = pi13  & n1146;
  assign n1298 = ~n1296 & ~n1297;
  assign n1299 = ~n1294 & ~n1295;
  assign n1300 = n9639 & ~n9666;
  assign n1301 = n9667 & ~n1285;
  assign n1302 = n9667 & ~n1300;
  assign n1303 = n9670 & n9671;
  assign n1304 = n9667 & ~n1289;
  assign n1305 = ~n9670 & n1304;
  assign n1306 = ~n1303 & ~n1305;
  assign n1307 = ~n1292 & n1306;
  assign n1308 = ~n1288 & n1307;
  assign n1309 = n1293 & n1306;
  assign n1310 = n9651 & n9672;
  assign n1311 = n9589 & n9608;
  assign n1312 = n9589 & ~n9608;
  assign n1313 = ~n9589 & n9608;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = ~n820 & ~n1311;
  assign n1316 = ~n1164 & n9673;
  assign n1317 = ~n821 & ~n9673;
  assign n1318 = n9569 & ~n9673;
  assign n1319 = ~n821 & n1164;
  assign n1320 = ~n9674 & ~n1319;
  assign n1321 = ~n821 & ~n1316;
  assign n1322 = n9569 & ~n9608;
  assign n1323 = n9569 & ~n1311;
  assign n1324 = n9673 & ~n1323;
  assign n1325 = n9673 & ~n1322;
  assign n1326 = ~n1164 & n9676;
  assign n1327 = n9675 & ~n1326;
  assign n1328 = ~n972 & n1327;
  assign n1329 = n972 & ~n1327;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = n9668 & n9670;
  assign n1332 = n9669 & ~n9670;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = ~n1149 & n9671;
  assign n1335 = n1149 & n1304;
  assign n1336 = ~n1334 & ~n1335;
  assign n1337 = ~n1332 & n1336;
  assign n1338 = ~n1331 & n1337;
  assign n1339 = n1333 & n1336;
  assign n1340 = n1330 & n9677;
  assign n1341 = ~n1328 & ~n1340;
  assign n1342 = ~n9651 & ~n9672;
  assign n1343 = ~n1310 & ~n1342;
  assign n1344 = ~n1341 & n1343;
  assign n1345 = ~n1310 & ~n1344;
  assign n1346 = ~n983 & ~n1345;
  assign n1347 = ~n9624 & n9626;
  assign n1348 = ~n1164 & n9667;
  assign n1349 = n1164 & ~n1289;
  assign n1350 = ~n9669 & ~n1349;
  assign n1351 = ~n1289 & ~n1348;
  assign n1352 = ~n1164 & n9671;
  assign n1353 = n9678 & ~n1352;
  assign n1354 = ~n1347 & n1353;
  assign n1355 = n1347 & ~n1353;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = n1142 & n1149;
  assign n1358 = n1137 & ~n1149;
  assign n1359 = ~n9624 & n9670;
  assign n1360 = n9624 & ~n9670;
  assign n1361 = ~n1359 & ~n1360;
  assign n1362 = ~n9649 & ~n9670;
  assign n1363 = ~n9649 & ~n1361;
  assign n1364 = ~n1358 & ~n9679;
  assign n1365 = ~n1357 & ~n1358;
  assign n1366 = ~n9679 & n1365;
  assign n1367 = ~n1357 & n1364;
  assign n1368 = n1356 & n9680;
  assign n1369 = ~n1356 & ~n9680;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = n983 & n1345;
  assign n1372 = ~n983 & ~n1346;
  assign n1373 = ~n983 & n1345;
  assign n1374 = ~n1345 & ~n1346;
  assign n1375 = n983 & ~n1345;
  assign n1376 = ~n9681 & ~n9682;
  assign n1377 = ~n1346 & ~n1371;
  assign n1378 = n1370 & ~n9683;
  assign n1379 = ~n1346 & ~n1378;
  assign n1380 = ~n1354 & ~n1368;
  assign n1381 = n1142 & ~n9670;
  assign n1382 = n1137 & n9670;
  assign n1383 = ~n9624 & n1164;
  assign n1384 = n9624 & ~n1164;
  assign n1385 = ~n1383 & ~n1384;
  assign n1386 = ~n9649 & n1164;
  assign n1387 = ~n9649 & n1385;
  assign n1388 = ~n1382 & ~n9684;
  assign n1389 = ~n1381 & ~n1382;
  assign n1390 = ~n9684 & n1389;
  assign n1391 = ~n1381 & n1388;
  assign n1392 = ~n1380 & n9685;
  assign n1393 = n1380 & ~n9685;
  assign n1394 = ~n1392 & ~n1393;
  assign n1395 = ~n1289 & ~n1347;
  assign n1396 = n1150 & n1395;
  assign n1397 = ~n1150 & ~n1395;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = n1394 & n1398;
  assign n1400 = ~n1394 & ~n1398;
  assign n1401 = ~n1399 & ~n1400;
  assign n1402 = ~n1379 & n1401;
  assign n1403 = ~pi22  & ~n92;
  assign n1404 = pi7  & ~n1403;
  assign n1405 = ~pi7  & n1403;
  assign n1406 = ~pi7  & ~n1403;
  assign n1407 = pi7  & n1403;
  assign n1408 = ~n1406 & ~n1407;
  assign n1409 = ~n1404 & ~n1405;
  assign n1410 = ~n9624 & n9686;
  assign n1411 = ~n192 & ~n715;
  assign n1412 = ~n715 & ~n1070;
  assign n1413 = ~n192 & n1412;
  assign n1414 = ~n470 & n1413;
  assign n1415 = n1071 & n1411;
  assign n1416 = ~n296 & ~n325;
  assign n1417 = ~n179 & ~n262;
  assign n1418 = ~n262 & n1416;
  assign n1419 = ~n179 & n1418;
  assign n1420 = ~n262 & ~n325;
  assign n1421 = ~n179 & ~n296;
  assign n1422 = n1420 & n1421;
  assign n1423 = n1416 & n1417;
  assign n1424 = ~n714 & ~n730;
  assign n1425 = ~n215 & ~n730;
  assign n1426 = ~n714 & n1425;
  assign n1427 = ~n215 & n1424;
  assign n1428 = n9688 & n9689;
  assign n1429 = n9687 & n9689;
  assign n1430 = n9688 & n1429;
  assign n1431 = n9687 & n1428;
  assign n1432 = ~n592 & ~n624;
  assign n1433 = ~n9550 & ~n432;
  assign n1434 = ~n311 & ~n432;
  assign n1435 = ~n9550 & n1434;
  assign n1436 = ~n311 & n1433;
  assign n1437 = ~n311 & n1432;
  assign n1438 = ~n432 & n1437;
  assign n1439 = ~n9550 & n1438;
  assign n1440 = n1432 & n9691;
  assign n1441 = n336 & n1223;
  assign n1442 = n336 & n780;
  assign n1443 = n1223 & n1442;
  assign n1444 = n780 & n1441;
  assign n1445 = n9692 & n9693;
  assign n1446 = n1223 & n9688;
  assign n1447 = n9692 & n1446;
  assign n1448 = n9687 & n1447;
  assign n1449 = ~n714 & n1448;
  assign n1450 = ~n334 & n1449;
  assign n1451 = ~n215 & n1450;
  assign n1452 = ~n335 & n1451;
  assign n1453 = n780 & n1452;
  assign n1454 = ~n730 & n1453;
  assign n1455 = n9690 & n1445;
  assign n1456 = ~n225 & ~n327;
  assign n1457 = ~n205 & ~n250;
  assign n1458 = n1456 & n1457;
  assign n1459 = ~n225 & n9694;
  assign n1460 = ~n327 & n1459;
  assign n1461 = ~n205 & n1460;
  assign n1462 = ~n250 & n1461;
  assign n1463 = n9694 & n1458;
  assign n1464 = n189 & n218;
  assign n1465 = n9532 & n607;
  assign n1466 = ~n582 & ~n9696;
  assign n1467 = ~n328 & n1466;
  assign n1468 = ~n217 & ~n331;
  assign n1469 = ~n217 & n1467;
  assign n1470 = ~n331 & n1469;
  assign n1471 = n1467 & n1468;
  assign n1472 = ~n9559 & ~n772;
  assign n1473 = ~n264 & ~n772;
  assign n1474 = ~n9559 & n1473;
  assign n1475 = ~n264 & n1472;
  assign n1476 = n406 & n9698;
  assign n1477 = n9590 & n1476;
  assign n1478 = n9697 & n1477;
  assign n1479 = ~n394 & ~n467;
  assign n1480 = ~n618 & n1479;
  assign n1481 = ~n897 & ~n995;
  assign n1482 = ~n260 & ~n9553;
  assign n1483 = ~n402 & ~n605;
  assign n1484 = n1482 & n1483;
  assign n1485 = n1481 & n1483;
  assign n1486 = n1482 & n1485;
  assign n1487 = n1481 & n1484;
  assign n1488 = n1480 & n1482;
  assign n1489 = ~n402 & n1488;
  assign n1490 = ~n897 & n1489;
  assign n1491 = ~n995 & n1490;
  assign n1492 = ~n605 & n1491;
  assign n1493 = n1480 & n9699;
  assign n1494 = ~n9541 & ~n332;
  assign n1495 = ~n332 & ~n9586;
  assign n1496 = ~n9541 & n1495;
  assign n1497 = ~n9586 & n1494;
  assign n1498 = ~n383 & ~n676;
  assign n1499 = n1124 & n1498;
  assign n1500 = n451 & n1498;
  assign n1501 = n1124 & n1500;
  assign n1502 = ~n175 & ~n383;
  assign n1503 = ~n301 & ~n9570;
  assign n1504 = ~n431 & ~n676;
  assign n1505 = n1503 & n1504;
  assign n1506 = n1502 & n1505;
  assign n1507 = n451 & n1499;
  assign n1508 = ~n383 & n9701;
  assign n1509 = ~n9570 & n1508;
  assign n1510 = ~n175 & n1509;
  assign n1511 = ~n301 & n1510;
  assign n1512 = ~n431 & n1511;
  assign n1513 = ~n676 & n1512;
  assign n1514 = n9701 & n9702;
  assign n1515 = n9700 & n9703;
  assign n1516 = n1478 & n1515;
  assign n1517 = n9695 & n9697;
  assign n1518 = n406 & n1517;
  assign n1519 = n9700 & n1518;
  assign n1520 = n9703 & n1519;
  assign n1521 = n9590 & n1520;
  assign n1522 = ~n772 & n1521;
  assign n1523 = ~n264 & n1522;
  assign n1524 = ~n9559 & n1523;
  assign n1525 = n9695 & n1516;
  assign n1526 = ~n296 & ~n663;
  assign n1527 = ~n296 & ~n898;
  assign n1528 = ~n663 & n1527;
  assign n1529 = ~n898 & n1526;
  assign n1530 = ~n258 & ~n605;
  assign n1531 = ~n226 & ~n9561;
  assign n1532 = ~n604 & ~n933;
  assign n1533 = ~n226 & ~n933;
  assign n1534 = n909 & n1533;
  assign n1535 = n1531 & n1532;
  assign n1536 = n1530 & n1532;
  assign n1537 = n1531 & n1536;
  assign n1538 = n1530 & n1531;
  assign n1539 = n1532 & n1538;
  assign n1540 = n1530 & n9706;
  assign n1541 = n9705 & n1530;
  assign n1542 = n909 & n1541;
  assign n1543 = ~n933 & n1542;
  assign n1544 = ~n226 & n1543;
  assign n1545 = n9705 & n9707;
  assign n1546 = ~n230 & ~n328;
  assign n1547 = ~n9570 & n625;
  assign n1548 = ~n624 & n1546;
  assign n1549 = ~n9570 & n1548;
  assign n1550 = ~n623 & n1549;
  assign n1551 = n1546 & n1547;
  assign n1552 = ~n205 & ~n284;
  assign n1553 = ~n205 & ~n351;
  assign n1554 = ~n284 & n1553;
  assign n1555 = ~n284 & ~n351;
  assign n1556 = ~n205 & n1555;
  assign n1557 = ~n351 & n1552;
  assign n1558 = ~n620 & ~n995;
  assign n1559 = n411 & n1558;
  assign n1560 = ~n205 & n1559;
  assign n1561 = ~n351 & n1560;
  assign n1562 = ~n284 & n1561;
  assign n1563 = n9710 & n1559;
  assign n1564 = ~n199 & ~n538;
  assign n1565 = ~n262 & ~n515;
  assign n1566 = ~n199 & ~n262;
  assign n1567 = ~n515 & ~n538;
  assign n1568 = n1566 & n1567;
  assign n1569 = n1564 & n1565;
  assign n1570 = ~n582 & ~n720;
  assign n1571 = ~n384 & ~n9564;
  assign n1572 = n1570 & n1571;
  assign n1573 = ~n9564 & ~n538;
  assign n1574 = n1565 & n1573;
  assign n1575 = ~n199 & ~n384;
  assign n1576 = n1570 & n1575;
  assign n1577 = n1574 & n1576;
  assign n1578 = n1566 & n1571;
  assign n1579 = n1567 & n1570;
  assign n1580 = n1578 & n1579;
  assign n1581 = n9712 & n1572;
  assign n1582 = n9711 & n9713;
  assign n1583 = n9709 & n9713;
  assign n1584 = n9711 & n1583;
  assign n1585 = n9709 & n1582;
  assign n1586 = n9709 & n1570;
  assign n1587 = n9708 & n1586;
  assign n1588 = n9711 & n1587;
  assign n1589 = ~n9564 & n1588;
  assign n1590 = ~n262 & n1589;
  assign n1591 = ~n199 & n1590;
  assign n1592 = ~n538 & n1591;
  assign n1593 = ~n515 & n1592;
  assign n1594 = ~n384 & n1593;
  assign n1595 = n9708 & n9714;
  assign n1596 = ~n243 & ~n9559;
  assign n1597 = ~n202 & ~n312;
  assign n1598 = ~n243 & ~n312;
  assign n1599 = ~n202 & ~n9559;
  assign n1600 = n1598 & n1599;
  assign n1601 = n1596 & n1597;
  assign n1602 = ~n312 & n9612;
  assign n1603 = ~n243 & n1602;
  assign n1604 = ~n202 & n1603;
  assign n1605 = ~n9559 & n1604;
  assign n1606 = n9612 & n9716;
  assign n1607 = ~n627 & ~n772;
  assign n1608 = ~n381 & ~n627;
  assign n1609 = ~n772 & n1608;
  assign n1610 = ~n381 & n1607;
  assign n1611 = ~n405 & ~n897;
  assign n1612 = n1248 & n1611;
  assign n1613 = n9718 & n1612;
  assign n1614 = n9554 & n9687;
  assign n1615 = n1613 & n1614;
  assign n1616 = n9554 & n1248;
  assign n1617 = n1611 & n1616;
  assign n1618 = n9717 & n1617;
  assign n1619 = n9687 & n1618;
  assign n1620 = ~n627 & n1619;
  assign n1621 = ~n772 & n1620;
  assign n1622 = ~n381 & n1621;
  assign n1623 = n9717 & n1615;
  assign n1624 = ~n250 & ~n383;
  assign n1625 = ~n383 & ~n583;
  assign n1626 = ~n250 & n1625;
  assign n1627 = ~n250 & ~n583;
  assign n1628 = ~n383 & n1627;
  assign n1629 = ~n583 & n1624;
  assign n1630 = ~n311 & ~n9696;
  assign n1631 = ~n511 & n1630;
  assign n1632 = n9540 & n1631;
  assign n1633 = n9540 & n9720;
  assign n1634 = n1631 & n1633;
  assign n1635 = n9720 & n1632;
  assign n1636 = ~n9544 & ~n394;
  assign n1637 = ~n552 & n1636;
  assign n1638 = ~n175 & ~n581;
  assign n1639 = ~n324 & ~n1037;
  assign n1640 = n1638 & n1639;
  assign n1641 = ~n324 & ~n581;
  assign n1642 = ~n175 & n1641;
  assign n1643 = ~n9544 & n1642;
  assign n1644 = ~n394 & n1643;
  assign n1645 = ~n552 & n1644;
  assign n1646 = ~n1037 & n1645;
  assign n1647 = ~n1037 & n1636;
  assign n1648 = ~n324 & ~n552;
  assign n1649 = n1638 & n1648;
  assign n1650 = n1647 & n1649;
  assign n1651 = ~n175 & ~n1037;
  assign n1652 = ~n552 & n1651;
  assign n1653 = ~n324 & ~n394;
  assign n1654 = ~n9544 & ~n581;
  assign n1655 = n1653 & n1654;
  assign n1656 = n1652 & n1655;
  assign n1657 = n1637 & n1640;
  assign n1658 = ~n294 & ~n574;
  assign n1659 = ~n554 & ~n1108;
  assign n1660 = n1658 & n1659;
  assign n1661 = n188 & n201;
  assign n1662 = ~n754 & ~n1661;
  assign n1663 = ~n265 & ~n871;
  assign n1664 = n1662 & n1663;
  assign n1665 = ~n554 & ~n1661;
  assign n1666 = ~n754 & ~n1108;
  assign n1667 = n1665 & n1666;
  assign n1668 = n1658 & n1663;
  assign n1669 = n1667 & n1668;
  assign n1670 = ~n871 & ~n1108;
  assign n1671 = n1665 & n1670;
  assign n1672 = ~n265 & ~n754;
  assign n1673 = n1658 & n1672;
  assign n1674 = n1671 & n1673;
  assign n1675 = ~n754 & ~n871;
  assign n1676 = n1658 & n1675;
  assign n1677 = n1111 & n1665;
  assign n1678 = n1676 & n1677;
  assign n1679 = n1660 & n1664;
  assign n1680 = n9722 & n9723;
  assign n1681 = n9721 & n1680;
  assign n1682 = n9719 & n1681;
  assign n1683 = n9540 & n1111;
  assign n1684 = n9720 & n1683;
  assign n1685 = n1631 & n1684;
  assign n1686 = n1665 & n1685;
  assign n1687 = n9722 & n1686;
  assign n1688 = n9719 & n1687;
  assign n1689 = n9715 & n1688;
  assign n1690 = ~n574 & n1689;
  assign n1691 = ~n871 & n1690;
  assign n1692 = ~n754 & n1691;
  assign n1693 = ~n294 & n1692;
  assign n1694 = n9715 & n1682;
  assign n1695 = ~n9704 & ~n9724;
  assign n1696 = ~n9589 & ~n1695;
  assign n1697 = n1410 & ~n1696;
  assign n1698 = ~n1410 & n1696;
  assign n1699 = ~n1697 & ~n1698;
  assign n1700 = pi8  & pi22 ;
  assign n1701 = pi8  & ~n93;
  assign n1702 = n965 & ~n1701;
  assign n1703 = ~n1700 & ~n1702;
  assign n1704 = ~n9624 & ~n1703;
  assign n1705 = n1699 & ~n1703;
  assign n1706 = ~n9624 & n1705;
  assign n1707 = n1699 & n1704;
  assign n1708 = ~n1697 & ~n9725;
  assign n1709 = n978 & n1142;
  assign n1710 = ~n978 & n1137;
  assign n1711 = n9624 & ~n9626;
  assign n1712 = ~n1347 & ~n1711;
  assign n1713 = ~n9626 & ~n9649;
  assign n1714 = ~n9649 & ~n1712;
  assign n1715 = ~n1710 & ~n9726;
  assign n1716 = ~n1709 & ~n1710;
  assign n1717 = ~n9726 & n1716;
  assign n1718 = ~n1709 & n1715;
  assign n1719 = ~n1708 & n9727;
  assign n1720 = n1164 & n9674;
  assign n1721 = ~n9673 & ~n1323;
  assign n1722 = ~n9569 & ~n9673;
  assign n1723 = ~n1164 & n9728;
  assign n1724 = ~n1720 & ~n1723;
  assign n1725 = n9670 & n9676;
  assign n1726 = ~n821 & n9673;
  assign n1727 = ~n9670 & n1726;
  assign n1728 = ~n1725 & ~n1727;
  assign n1729 = ~n1720 & n1728;
  assign n1730 = ~n1723 & n1729;
  assign n1731 = ~n1720 & ~n1725;
  assign n1732 = ~n1723 & ~n1727;
  assign n1733 = n1731 & n1732;
  assign n1734 = n1724 & n1728;
  assign n1735 = ~n1149 & n9668;
  assign n1736 = n1149 & n9669;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = n9626 & n9671;
  assign n1739 = ~n9626 & n1304;
  assign n1740 = ~n1738 & ~n1739;
  assign n1741 = ~n1736 & n1740;
  assign n1742 = ~n1735 & n1741;
  assign n1743 = n1737 & n1740;
  assign n1744 = n9729 & n9730;
  assign n1745 = ~n9729 & ~n9730;
  assign n1746 = n9729 & ~n9730;
  assign n1747 = ~n9729 & n9730;
  assign n1748 = ~n1746 & ~n1747;
  assign n1749 = ~n1744 & ~n1745;
  assign n1750 = ~n9625 & n1142;
  assign n1751 = n9625 & n1137;
  assign n1752 = n9624 & n978;
  assign n1753 = ~n979 & ~n1752;
  assign n1754 = n978 & ~n9649;
  assign n1755 = ~n9649 & ~n1753;
  assign n1756 = ~n1751 & ~n9732;
  assign n1757 = ~n1750 & ~n1751;
  assign n1758 = ~n9732 & n1757;
  assign n1759 = ~n1750 & n1756;
  assign n1760 = ~n9731 & n9733;
  assign n1761 = ~n1744 & ~n1760;
  assign n1762 = n1708 & ~n9727;
  assign n1763 = n9727 & ~n1719;
  assign n1764 = ~n1708 & ~n1719;
  assign n1765 = ~n1763 & ~n1764;
  assign n1766 = ~n1719 & ~n1762;
  assign n1767 = ~n1761 & ~n9734;
  assign n1768 = ~n1719 & ~n1767;
  assign n1769 = ~n979 & ~n981;
  assign n1770 = ~n982 & ~n1769;
  assign n1771 = ~n1768 & n1770;
  assign n1772 = n1768 & ~n1770;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = n1341 & ~n1343;
  assign n1775 = ~n1344 & ~n1774;
  assign n1776 = n1773 & n1775;
  assign n1777 = ~n1771 & ~n1776;
  assign n1778 = ~n1370 & n9683;
  assign n1779 = ~n9683 & ~n1378;
  assign n1780 = ~n1370 & ~n9683;
  assign n1781 = n1370 & ~n1378;
  assign n1782 = n1370 & n9683;
  assign n1783 = ~n9735 & ~n9736;
  assign n1784 = ~n1378 & ~n1778;
  assign n1785 = ~n1777 & ~n9737;
  assign n1786 = n1142 & n1703;
  assign n1787 = n1137 & ~n1703;
  assign n1788 = n9624 & ~n9625;
  assign n1789 = ~n972 & ~n1788;
  assign n1790 = ~n9625 & ~n9649;
  assign n1791 = ~n9649 & ~n1789;
  assign n1792 = ~n1787 & ~n9738;
  assign n1793 = ~n1786 & ~n1787;
  assign n1794 = ~n9738 & n1793;
  assign n1795 = ~n1786 & n1792;
  assign n1796 = n9626 & n9668;
  assign n1797 = ~n9626 & n9669;
  assign n1798 = ~n1796 & ~n1797;
  assign n1799 = ~n978 & n9671;
  assign n1800 = n978 & n1304;
  assign n1801 = ~n1799 & ~n1800;
  assign n1802 = ~n1797 & n1801;
  assign n1803 = ~n1796 & n1802;
  assign n1804 = n1798 & n1801;
  assign n1805 = n9739 & n9740;
  assign n1806 = ~n9739 & ~n9740;
  assign n1807 = ~n1805 & ~n1806;
  assign n1808 = ~n9537 & ~n327;
  assign n1809 = ~n264 & ~n476;
  assign n1810 = ~n264 & n1808;
  assign n1811 = ~n476 & n1810;
  assign n1812 = n1808 & n1809;
  assign n1813 = ~n249 & ~n995;
  assign n1814 = ~n249 & ~n294;
  assign n1815 = ~n995 & n1814;
  assign n1816 = ~n294 & n1813;
  assign n1817 = ~n295 & ~n515;
  assign n1818 = ~n1108 & n1817;
  assign n1819 = n9742 & n1818;
  assign n1820 = n9741 & n9742;
  assign n1821 = n1818 & n1820;
  assign n1822 = n9741 & n1819;
  assign n1823 = ~n226 & ~n897;
  assign n1824 = ~n260 & ~n262;
  assign n1825 = ~n226 & ~n262;
  assign n1826 = ~n260 & ~n897;
  assign n1827 = n1825 & n1826;
  assign n1828 = n1823 & n1824;
  assign n1829 = n382 & n9744;
  assign n1830 = n9692 & n1829;
  assign n1831 = n9692 & n9743;
  assign n1832 = n382 & n1831;
  assign n1833 = ~n262 & n1832;
  assign n1834 = ~n897 & n1833;
  assign n1835 = ~n226 & n1834;
  assign n1836 = ~n260 & n1835;
  assign n1837 = n9743 & n1830;
  assign n1838 = ~n730 & ~n1190;
  assign n1839 = ~n404 & ~n776;
  assign n1840 = ~n205 & ~n554;
  assign n1841 = n1839 & n1840;
  assign n1842 = n1838 & n1841;
  assign n1843 = ~n394 & ~n620;
  assign n1844 = ~n534 & n1843;
  assign n1845 = ~n468 & ~n1661;
  assign n1846 = n664 & n1845;
  assign n1847 = n1844 & n1846;
  assign n1848 = n664 & n1838;
  assign n1849 = n1838 & n1839;
  assign n1850 = n664 & n1849;
  assign n1851 = ~n404 & ~n583;
  assign n1852 = ~n663 & ~n776;
  assign n1853 = n1838 & n1852;
  assign n1854 = n1851 & n1853;
  assign n1855 = n1839 & n1848;
  assign n1856 = ~n468 & ~n534;
  assign n1857 = ~n205 & n1856;
  assign n1858 = n1665 & n1843;
  assign n1859 = ~n205 & ~n468;
  assign n1860 = ~n394 & n1859;
  assign n1861 = ~n534 & ~n620;
  assign n1862 = n1665 & n1861;
  assign n1863 = n1860 & n1862;
  assign n1864 = n1857 & n1858;
  assign n1865 = n9746 & n9747;
  assign n1866 = n1842 & n1847;
  assign n1867 = ~n245 & ~n511;
  assign n1868 = ~n265 & ~n1015;
  assign n1869 = ~n607 & n1868;
  assign n1870 = ~n265 & ~n511;
  assign n1871 = ~n245 & ~n265;
  assign n1872 = ~n511 & n1871;
  assign n1873 = ~n245 & n1870;
  assign n1874 = ~n607 & n9749;
  assign n1875 = ~n1015 & n1874;
  assign n1876 = ~n607 & ~n1015;
  assign n1877 = n9749 & n1876;
  assign n1878 = n1867 & n1869;
  assign n1879 = n9560 & n9750;
  assign n1880 = n9560 & n9747;
  assign n1881 = n9746 & n9750;
  assign n1882 = n1880 & n1881;
  assign n1883 = n9748 & n1879;
  assign n1884 = ~n217 & ~n284;
  assign n1885 = ~n195 & ~n772;
  assign n1886 = n1884 & n1885;
  assign n1887 = n326 & n753;
  assign n1888 = ~n415 & ~n533;
  assign n1889 = n1570 & n1888;
  assign n1890 = n1887 & n1889;
  assign n1891 = n326 & n1570;
  assign n1892 = n753 & n1891;
  assign n1893 = ~n415 & n1892;
  assign n1894 = ~n772 & n1893;
  assign n1895 = ~n217 & n1894;
  assign n1896 = ~n195 & n1895;
  assign n1897 = ~n533 & n1896;
  assign n1898 = ~n284 & n1897;
  assign n1899 = ~n284 & ~n533;
  assign n1900 = ~n195 & ~n415;
  assign n1901 = n1899 & n1900;
  assign n1902 = ~n217 & ~n772;
  assign n1903 = n753 & n1902;
  assign n1904 = n1891 & n1903;
  assign n1905 = n1901 & n1904;
  assign n1906 = ~n284 & ~n772;
  assign n1907 = n1900 & n1906;
  assign n1908 = ~n217 & ~n533;
  assign n1909 = n753 & n1908;
  assign n1910 = n1891 & n1909;
  assign n1911 = n1907 & n1910;
  assign n1912 = n1885 & n1899;
  assign n1913 = ~n217 & ~n415;
  assign n1914 = n326 & n1913;
  assign n1915 = n753 & n1570;
  assign n1916 = n1914 & n1915;
  assign n1917 = n1912 & n1916;
  assign n1918 = n1886 & n1890;
  assign n1919 = ~n334 & ~n1070;
  assign n1920 = ~n538 & n1919;
  assign n1921 = ~n623 & ~n770;
  assign n1922 = n993 & n1921;
  assign n1923 = n1638 & n1922;
  assign n1924 = n993 & ~n1070;
  assign n1925 = ~n334 & n1924;
  assign n1926 = ~n581 & n1925;
  assign n1927 = ~n175 & n1926;
  assign n1928 = ~n538 & n1927;
  assign n1929 = ~n770 & n1928;
  assign n1930 = ~n623 & n1929;
  assign n1931 = ~n334 & ~n770;
  assign n1932 = ~n1070 & n1931;
  assign n1933 = ~n538 & ~n623;
  assign n1934 = n993 & n1933;
  assign n1935 = n1638 & n1934;
  assign n1936 = n1932 & n1935;
  assign n1937 = ~n770 & ~n1070;
  assign n1938 = ~n538 & n1937;
  assign n1939 = ~n175 & ~n623;
  assign n1940 = n866 & n1939;
  assign n1941 = n993 & n1940;
  assign n1942 = n1938 & n1941;
  assign n1943 = n1920 & n1923;
  assign n1944 = n9752 & n9753;
  assign n1945 = n9751 & n1944;
  assign n1946 = n9560 & n9746;
  assign n1947 = n1665 & n1946;
  assign n1948 = n9753 & n1947;
  assign n1949 = n9750 & n1948;
  assign n1950 = n9752 & n1949;
  assign n1951 = n9745 & n1950;
  assign n1952 = ~n468 & n1951;
  assign n1953 = ~n394 & n1952;
  assign n1954 = ~n534 & n1953;
  assign n1955 = ~n620 & n1954;
  assign n1956 = ~n205 & n1955;
  assign n1957 = n9745 & n1945;
  assign n1958 = ~n296 & ~n9561;
  assign n1959 = ~n990 & n1958;
  assign n1960 = n1255 & n1959;
  assign n1961 = n9720 & n1960;
  assign n1962 = ~n215 & ~n311;
  assign n1963 = n991 & n1962;
  assign n1964 = n775 & n1838;
  assign n1965 = n991 & n1838;
  assign n1966 = n775 & n1965;
  assign n1967 = ~n215 & n1966;
  assign n1968 = ~n311 & n1967;
  assign n1969 = n775 & n1962;
  assign n1970 = n1965 & n1969;
  assign n1971 = n1963 & n1964;
  assign n1972 = ~n262 & ~n332;
  assign n1973 = ~n386 & ~n674;
  assign n1974 = n606 & n1973;
  assign n1975 = n1972 & n1974;
  assign n1976 = n9750 & n1975;
  assign n1977 = n9755 & n1976;
  assign n1978 = n1255 & n9720;
  assign n1979 = n909 & n1978;
  assign n1980 = n9750 & n1979;
  assign n1981 = n9755 & n1980;
  assign n1982 = ~n296 & n1981;
  assign n1983 = ~n262 & n1982;
  assign n1984 = ~n386 & n1983;
  assign n1985 = ~n990 & n1984;
  assign n1986 = ~n332 & n1985;
  assign n1987 = ~n605 & n1986;
  assign n1988 = ~n674 & n1987;
  assign n1989 = ~n296 & ~n605;
  assign n1990 = ~n990 & n1989;
  assign n1991 = n1255 & n1990;
  assign n1992 = n9720 & n1991;
  assign n1993 = n909 & n1973;
  assign n1994 = n1972 & n1993;
  assign n1995 = n9750 & n1994;
  assign n1996 = n9755 & n1995;
  assign n1997 = n1992 & n1996;
  assign n1998 = ~n990 & n1973;
  assign n1999 = n1255 & n1998;
  assign n2000 = n9720 & n1999;
  assign n2001 = n909 & n1989;
  assign n2002 = n1972 & n2001;
  assign n2003 = n9750 & n2002;
  assign n2004 = n9755 & n2003;
  assign n2005 = n2000 & n2004;
  assign n2006 = ~n605 & ~n990;
  assign n2007 = ~n674 & n2006;
  assign n2008 = n1255 & n2007;
  assign n2009 = n9720 & n2008;
  assign n2010 = ~n296 & ~n386;
  assign n2011 = n1972 & n2010;
  assign n2012 = n909 & n2011;
  assign n2013 = n9750 & n2012;
  assign n2014 = n9755 & n2013;
  assign n2015 = n2009 & n2014;
  assign n2016 = n1961 & n1977;
  assign n2017 = ~n295 & ~n581;
  assign n2018 = ~n552 & ~n682;
  assign n2019 = ~n581 & ~n682;
  assign n2020 = ~n295 & ~n552;
  assign n2021 = n2019 & n2020;
  assign n2022 = n2017 & n2018;
  assign n2023 = ~n205 & ~n772;
  assign n2024 = n1247 & n1546;
  assign n2025 = n2023 & n2024;
  assign n2026 = n1247 & n2019;
  assign n2027 = ~n682 & n2024;
  assign n2028 = ~n581 & n2027;
  assign n2029 = n1546 & n2026;
  assign n2030 = ~n295 & n9758;
  assign n2031 = ~n772 & n2030;
  assign n2032 = ~n205 & n2031;
  assign n2033 = ~n552 & n2032;
  assign n2034 = ~n295 & ~n772;
  assign n2035 = ~n205 & ~n552;
  assign n2036 = n2034 & n2035;
  assign n2037 = n9758 & n2036;
  assign n2038 = n9757 & n2025;
  assign n2039 = ~n623 & ~n776;
  assign n2040 = n550 & n2039;
  assign n2041 = n9552 & n1662;
  assign n2042 = n2040 & n2041;
  assign n2043 = ~n384 & ~n480;
  assign n2044 = ~n219 & n2043;
  assign n2045 = n1480 & n2044;
  assign n2046 = ~n219 & ~n623;
  assign n2047 = n550 & n2046;
  assign n2048 = n2041 & n2047;
  assign n2049 = ~n480 & ~n776;
  assign n2050 = ~n384 & n2049;
  assign n2051 = n1480 & n2050;
  assign n2052 = n2048 & n2051;
  assign n2053 = ~n219 & ~n384;
  assign n2054 = ~n480 & ~n754;
  assign n2055 = n2053 & n2054;
  assign n2056 = n550 & n2055;
  assign n2057 = ~n776 & ~n1661;
  assign n2058 = ~n623 & n2057;
  assign n2059 = n9552 & n2058;
  assign n2060 = n1480 & n2059;
  assign n2061 = n2056 & n2060;
  assign n2062 = n2042 & n2045;
  assign n2063 = n9552 & n1480;
  assign n2064 = ~n1661 & n2063;
  assign n2065 = n9759 & n2064;
  assign n2066 = n550 & n2065;
  assign n2067 = ~n219 & n2066;
  assign n2068 = ~n776 & n2067;
  assign n2069 = ~n754 & n2068;
  assign n2070 = ~n623 & n2069;
  assign n2071 = ~n384 & n2070;
  assign n2072 = ~n480 & n2071;
  assign n2073 = n9759 & n9760;
  assign n2074 = ~n397 & ~n592;
  assign n2075 = ~n720 & n2074;
  assign n2076 = ~n9562 & ~n1108;
  assign n2077 = ~n9564 & ~n627;
  assign n2078 = n2076 & n2077;
  assign n2079 = n1010 & n2078;
  assign n2080 = ~n397 & ~n720;
  assign n2081 = ~n9562 & ~n592;
  assign n2082 = ~n397 & n2081;
  assign n2083 = ~n720 & n2082;
  assign n2084 = ~n9562 & ~n720;
  assign n2085 = n2074 & n2084;
  assign n2086 = n2080 & n2081;
  assign n2087 = ~n1108 & n2077;
  assign n2088 = n1010 & n2087;
  assign n2089 = n9762 & n2088;
  assign n2090 = n2075 & n2079;
  assign n2091 = ~n431 & ~n770;
  assign n2092 = ~n190 & ~n676;
  assign n2093 = n2091 & n2092;
  assign n2094 = ~n431 & n1258;
  assign n2095 = ~n770 & n2094;
  assign n2096 = ~n676 & n2095;
  assign n2097 = ~n190 & n2096;
  assign n2098 = ~n190 & ~n9541;
  assign n2099 = n1084 & n2098;
  assign n2100 = n1258 & n2092;
  assign n2101 = n2091 & n9765;
  assign n2102 = n1258 & n2093;
  assign n2103 = n406 & n685;
  assign n2104 = n486 & n685;
  assign n2105 = n406 & n2104;
  assign n2106 = n486 & n2103;
  assign n2107 = n9764 & n9766;
  assign n2108 = n9763 & n2107;
  assign n2109 = n9761 & n2108;
  assign n2110 = n486 & n9762;
  assign n2111 = n1010 & n2110;
  assign n2112 = n685 & n2111;
  assign n2113 = n9764 & n2112;
  assign n2114 = n406 & n2113;
  assign n2115 = n9761 & n2114;
  assign n2116 = n9756 & n2115;
  assign n2117 = ~n9564 & n2116;
  assign n2118 = ~n627 & n2117;
  assign n2119 = ~n1108 & n2118;
  assign n2120 = n9756 & n2108;
  assign n2121 = n9761 & n2120;
  assign n2122 = n9756 & n2109;
  assign n2123 = ~n9754 & ~n9767;
  assign n2124 = ~n9724 & ~n2123;
  assign n2125 = n9754 & ~n2124;
  assign n2126 = n9724 & n9754;
  assign n2127 = pi6  & pi22 ;
  assign n2128 = pi6  & ~n91;
  assign n2129 = n1403 & ~n2128;
  assign n2130 = ~n2127 & ~n2129;
  assign n2131 = ~n9624 & ~n2130;
  assign n2132 = ~n9724 & n9767;
  assign n2133 = ~n9754 & n9767;
  assign n2134 = ~n9724 & n2133;
  assign n2135 = ~n9754 & n2124;
  assign n2136 = ~n9754 & n2132;
  assign n2137 = n2131 & ~n9769;
  assign n2138 = ~n9768 & n2131;
  assign n2139 = ~n9769 & n2138;
  assign n2140 = ~n9768 & ~n2139;
  assign n2141 = ~n9768 & ~n2137;
  assign n2142 = n1807 & ~n9770;
  assign n2143 = ~n1805 & ~n2142;
  assign n2144 = n9704 & n9724;
  assign n2145 = ~n9704 & n9724;
  assign n2146 = n9704 & ~n9724;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~n1695 & ~n2144;
  assign n2149 = ~n1164 & n9771;
  assign n2150 = ~n1696 & ~n9771;
  assign n2151 = n9589 & ~n9771;
  assign n2152 = n1164 & ~n1696;
  assign n2153 = ~n9772 & ~n2152;
  assign n2154 = ~n1696 & ~n2149;
  assign n2155 = n9589 & ~n2144;
  assign n2156 = n9771 & ~n2155;
  assign n2157 = ~n1164 & n2156;
  assign n2158 = n2149 & ~n2155;
  assign n2159 = n9773 & ~n9774;
  assign n2160 = ~n1410 & n2159;
  assign n2161 = n1410 & ~n2159;
  assign n2162 = ~n2160 & ~n2161;
  assign n2163 = ~n9670 & n9674;
  assign n2164 = n9670 & n9728;
  assign n2165 = ~n2163 & ~n2164;
  assign n2166 = ~n1149 & n9676;
  assign n2167 = n1149 & n1726;
  assign n2168 = ~n2166 & ~n2167;
  assign n2169 = ~n2163 & n2168;
  assign n2170 = ~n2164 & n2169;
  assign n2171 = ~n2163 & ~n2166;
  assign n2172 = ~n2164 & ~n2167;
  assign n2173 = n2171 & n2172;
  assign n2174 = n2165 & n2168;
  assign n2175 = n2162 & n9775;
  assign n2176 = ~n2160 & ~n2175;
  assign n2177 = ~n2143 & ~n2176;
  assign n2178 = ~n1699 & ~n1704;
  assign n2179 = ~n9624 & ~n9725;
  assign n2180 = ~n1703 & n2179;
  assign n2181 = n1704 & ~n9725;
  assign n2182 = n1699 & ~n9725;
  assign n2183 = ~n9776 & ~n2182;
  assign n2184 = ~n9725 & ~n2178;
  assign n2185 = n2143 & n2176;
  assign n2186 = ~n2143 & ~n2177;
  assign n2187 = ~n2143 & n2176;
  assign n2188 = ~n2176 & ~n2177;
  assign n2189 = n2143 & ~n2176;
  assign n2190 = ~n9778 & ~n9779;
  assign n2191 = ~n2177 & ~n2185;
  assign n2192 = ~n9777 & ~n9780;
  assign n2193 = ~n2177 & ~n2192;
  assign n2194 = ~n1330 & ~n9677;
  assign n2195 = ~n1340 & ~n2194;
  assign n2196 = ~n2193 & n2195;
  assign n2197 = n2193 & ~n2195;
  assign n2198 = ~n2196 & ~n2197;
  assign n2199 = n1761 & n9734;
  assign n2200 = ~n1761 & ~n1767;
  assign n2201 = ~n9734 & ~n1767;
  assign n2202 = ~n2200 & ~n2201;
  assign n2203 = ~n1767 & ~n2199;
  assign n2204 = n2198 & ~n9781;
  assign n2205 = ~n2196 & ~n2204;
  assign n2206 = ~n1773 & ~n1775;
  assign n2207 = ~n1776 & ~n2206;
  assign n2208 = ~n2205 & n2207;
  assign n2209 = ~n2198 & n9781;
  assign n2210 = n2198 & ~n2204;
  assign n2211 = ~n9781 & ~n2204;
  assign n2212 = ~n2210 & ~n2211;
  assign n2213 = ~n2204 & ~n2209;
  assign n2214 = n1142 & ~n9686;
  assign n2215 = n1137 & n9686;
  assign n2216 = n9624 & n1703;
  assign n2217 = ~n1704 & ~n2216;
  assign n2218 = ~n9649 & n1703;
  assign n2219 = ~n9649 & ~n2217;
  assign n2220 = ~n2215 & ~n9783;
  assign n2221 = ~n2214 & ~n2215;
  assign n2222 = ~n9783 & n2221;
  assign n2223 = ~n2214 & n2220;
  assign n2224 = ~n978 & n9668;
  assign n2225 = n978 & n9669;
  assign n2226 = ~n2224 & ~n2225;
  assign n2227 = n9625 & n9671;
  assign n2228 = ~n9625 & n1304;
  assign n2229 = ~n2227 & ~n2228;
  assign n2230 = ~n2225 & n2229;
  assign n2231 = ~n2224 & n2230;
  assign n2232 = n2226 & n2229;
  assign n2233 = n9784 & n9785;
  assign n2234 = ~n9784 & ~n9785;
  assign n2235 = ~n9784 & n9785;
  assign n2236 = n9784 & ~n9785;
  assign n2237 = ~n2235 & ~n2236;
  assign n2238 = ~n2233 & ~n2234;
  assign n2239 = ~n9771 & ~n2155;
  assign n2240 = ~n9589 & ~n9771;
  assign n2241 = ~n1164 & n9787;
  assign n2242 = n1164 & n9772;
  assign n2243 = ~n2241 & ~n2242;
  assign n2244 = n9670 & n2156;
  assign n2245 = ~n1696 & n9771;
  assign n2246 = ~n9670 & n2245;
  assign n2247 = ~n2244 & ~n2246;
  assign n2248 = ~n2242 & n2247;
  assign n2249 = ~n2241 & n2248;
  assign n2250 = n2243 & n2247;
  assign n2251 = ~n9786 & n9788;
  assign n2252 = ~n2233 & ~n2251;
  assign n2253 = ~n2162 & ~n9775;
  assign n2254 = ~n2175 & ~n2253;
  assign n2255 = ~n2252 & n2254;
  assign n2256 = ~n1807 & n9770;
  assign n2257 = ~n2142 & ~n2256;
  assign n2258 = n2252 & ~n2254;
  assign n2259 = ~n2252 & ~n2255;
  assign n2260 = n2254 & ~n2255;
  assign n2261 = ~n2259 & ~n2260;
  assign n2262 = ~n2255 & ~n2258;
  assign n2263 = n2257 & ~n9789;
  assign n2264 = ~n2255 & ~n2263;
  assign n2265 = n9731 & ~n9733;
  assign n2266 = n9733 & ~n1760;
  assign n2267 = n9731 & n9733;
  assign n2268 = ~n9731 & ~n1760;
  assign n2269 = ~n9731 & ~n9733;
  assign n2270 = ~n9790 & ~n9791;
  assign n2271 = ~n1760 & ~n2265;
  assign n2272 = n2264 & n9792;
  assign n2273 = ~n2264 & ~n9792;
  assign n2274 = n9777 & n9780;
  assign n2275 = ~n9780 & ~n2192;
  assign n2276 = n9777 & ~n9780;
  assign n2277 = ~n9777 & ~n2192;
  assign n2278 = ~n9777 & n9780;
  assign n2279 = ~n9793 & ~n9794;
  assign n2280 = ~n2192 & ~n2274;
  assign n2281 = ~n2273 & n9795;
  assign n2282 = ~n2264 & ~n2273;
  assign n2283 = ~n9792 & ~n2273;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = ~n2272 & ~n2273;
  assign n2286 = ~n9795 & ~n9796;
  assign n2287 = ~n2273 & ~n2286;
  assign n2288 = ~n2272 & ~n2281;
  assign n2289 = ~n9782 & ~n9797;
  assign n2290 = ~n9768 & ~n9769;
  assign n2291 = n2131 & ~n2139;
  assign n2292 = n2131 & ~n2290;
  assign n2293 = ~n9769 & n9770;
  assign n2294 = ~n2137 & n2290;
  assign n2295 = ~n9798 & ~n9799;
  assign n2296 = n1149 & n9674;
  assign n2297 = ~n1149 & n9728;
  assign n2298 = ~n2296 & ~n2297;
  assign n2299 = n9626 & n9676;
  assign n2300 = ~n9626 & n1726;
  assign n2301 = ~n2299 & ~n2300;
  assign n2302 = ~n2296 & n2301;
  assign n2303 = ~n2297 & n2302;
  assign n2304 = ~n2296 & ~n2299;
  assign n2305 = ~n2297 & ~n2300;
  assign n2306 = n2304 & n2305;
  assign n2307 = n2298 & n2301;
  assign n2308 = ~n2295 & n9800;
  assign n2309 = n9528 & ~n9624;
  assign n2310 = ~n9754 & n2309;
  assign n2311 = n9754 & ~n2309;
  assign n2312 = ~n2310 & ~n2311;
  assign n2313 = n9754 & n9767;
  assign n2314 = n9754 & ~n9767;
  assign n2315 = ~n2133 & ~n2314;
  assign n2316 = ~n2123 & ~n2313;
  assign n2317 = ~n1164 & n9801;
  assign n2318 = ~n2124 & ~n9801;
  assign n2319 = n9724 & ~n9801;
  assign n2320 = n1164 & ~n2124;
  assign n2321 = ~n9802 & ~n2320;
  assign n2322 = ~n2124 & ~n2317;
  assign n2323 = n9724 & ~n2313;
  assign n2324 = n9801 & ~n2323;
  assign n2325 = ~n1164 & n2324;
  assign n2326 = n2317 & ~n2323;
  assign n2327 = n9803 & ~n9804;
  assign n2328 = ~n2310 & n2327;
  assign n2329 = ~n2311 & n2328;
  assign n2330 = n2312 & n2327;
  assign n2331 = ~n2310 & ~n9805;
  assign n2332 = n2295 & ~n9800;
  assign n2333 = ~n2308 & ~n2332;
  assign n2334 = ~n2331 & n2333;
  assign n2335 = ~n2308 & ~n2334;
  assign n2336 = n9670 & n9787;
  assign n2337 = ~n9670 & n9772;
  assign n2338 = ~n2336 & ~n2337;
  assign n2339 = ~n1149 & n2156;
  assign n2340 = n1149 & n2245;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = ~n2337 & n2341;
  assign n2343 = ~n2336 & n2342;
  assign n2344 = n2338 & n2341;
  assign n2345 = ~n9626 & n9674;
  assign n2346 = n9626 & n9728;
  assign n2347 = ~n2345 & ~n2346;
  assign n2348 = ~n978 & n9676;
  assign n2349 = n978 & n1726;
  assign n2350 = ~n2348 & ~n2349;
  assign n2351 = ~n2345 & n2350;
  assign n2352 = ~n2346 & n2351;
  assign n2353 = ~n2345 & ~n2348;
  assign n2354 = ~n2346 & ~n2349;
  assign n2355 = n2353 & n2354;
  assign n2356 = n2347 & n2350;
  assign n2357 = n9806 & n9807;
  assign n2358 = ~n9806 & ~n9807;
  assign n2359 = n9806 & ~n9807;
  assign n2360 = ~n9806 & n9807;
  assign n2361 = ~n2359 & ~n2360;
  assign n2362 = ~n2357 & ~n2358;
  assign n2363 = n9625 & n9668;
  assign n2364 = ~n9625 & n9669;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = n9671 & ~n1703;
  assign n2367 = n1304 & n1703;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = ~n2364 & n2368;
  assign n2370 = ~n2363 & n2369;
  assign n2371 = n2365 & n2368;
  assign n2372 = ~n9808 & n9809;
  assign n2373 = ~n2357 & ~n2372;
  assign n2374 = n9786 & ~n9788;
  assign n2375 = ~n2251 & ~n2374;
  assign n2376 = ~n2373 & n2375;
  assign n2377 = ~n83 & ~n9624;
  assign n2378 = ~n9754 & n2377;
  assign n2379 = n9754 & ~n2377;
  assign n2380 = ~n2378 & ~n2379;
  assign n2381 = ~n9801 & ~n2323;
  assign n2382 = ~n9724 & ~n9801;
  assign n2383 = ~n1164 & n9810;
  assign n2384 = n1164 & n9802;
  assign n2385 = ~n2383 & ~n2384;
  assign n2386 = n9670 & n2324;
  assign n2387 = ~n2124 & n9801;
  assign n2388 = ~n2132 & n9801;
  assign n2389 = ~n9670 & n9811;
  assign n2390 = ~n2386 & ~n2389;
  assign n2391 = ~n2384 & n2390;
  assign n2392 = ~n2383 & n2391;
  assign n2393 = n2385 & n2390;
  assign n2394 = ~n2378 & n9812;
  assign n2395 = ~n2379 & n2394;
  assign n2396 = n2380 & n9812;
  assign n2397 = ~n2378 & ~n9813;
  assign n2398 = n1142 & n2130;
  assign n2399 = n1137 & ~n2130;
  assign n2400 = n9624 & ~n9686;
  assign n2401 = ~n1410 & ~n2400;
  assign n2402 = ~n9649 & ~n9686;
  assign n2403 = ~n9649 & ~n2401;
  assign n2404 = ~n2399 & ~n9814;
  assign n2405 = ~n2398 & ~n2399;
  assign n2406 = ~n9814 & n2405;
  assign n2407 = ~n2398 & n2404;
  assign n2408 = ~n2397 & n9815;
  assign n2409 = n2397 & ~n9815;
  assign n2410 = ~n2408 & ~n2409;
  assign n2411 = n978 & n9674;
  assign n2412 = ~n978 & n9728;
  assign n2413 = ~n2411 & ~n2412;
  assign n2414 = n9625 & n9676;
  assign n2415 = ~n9625 & n1726;
  assign n2416 = ~n2414 & ~n2415;
  assign n2417 = ~n2411 & n2416;
  assign n2418 = ~n2412 & n2417;
  assign n2419 = ~n2411 & ~n2414;
  assign n2420 = ~n2412 & ~n2415;
  assign n2421 = n2419 & n2420;
  assign n2422 = n2413 & n2416;
  assign n2423 = ~n1149 & n9787;
  assign n2424 = n1149 & n9772;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = n9626 & n2156;
  assign n2427 = ~n9626 & n2245;
  assign n2428 = ~n2426 & ~n2427;
  assign n2429 = ~n2424 & n2428;
  assign n2430 = ~n2423 & n2429;
  assign n2431 = n2425 & n2428;
  assign n2432 = n9816 & n9817;
  assign n2433 = ~n9816 & ~n9817;
  assign n2434 = ~n9816 & n9817;
  assign n2435 = n9816 & ~n9817;
  assign n2436 = ~n2434 & ~n2435;
  assign n2437 = ~n2432 & ~n2433;
  assign n2438 = n9668 & ~n1703;
  assign n2439 = n9669 & n1703;
  assign n2440 = ~n2438 & ~n2439;
  assign n2441 = n9671 & n9686;
  assign n2442 = n1304 & ~n9686;
  assign n2443 = ~n2441 & ~n2442;
  assign n2444 = ~n2439 & n2443;
  assign n2445 = ~n2438 & n2444;
  assign n2446 = n2440 & n2443;
  assign n2447 = ~n9818 & n9819;
  assign n2448 = ~n2432 & ~n2447;
  assign n2449 = n2410 & ~n2448;
  assign n2450 = ~n2408 & ~n2449;
  assign n2451 = n2373 & ~n2375;
  assign n2452 = ~n2376 & ~n2451;
  assign n2453 = ~n2450 & n2452;
  assign n2454 = ~n2376 & ~n2453;
  assign n2455 = ~n2335 & ~n2454;
  assign n2456 = ~n2257 & n9789;
  assign n2457 = n2257 & ~n2263;
  assign n2458 = ~n9789 & ~n2263;
  assign n2459 = ~n2457 & ~n2458;
  assign n2460 = ~n2263 & ~n2456;
  assign n2461 = n2335 & n2454;
  assign n2462 = ~n2335 & ~n2455;
  assign n2463 = ~n2335 & n2454;
  assign n2464 = ~n2454 & ~n2455;
  assign n2465 = n2335 & ~n2454;
  assign n2466 = ~n9821 & ~n9822;
  assign n2467 = ~n2455 & ~n2461;
  assign n2468 = ~n9820 & ~n9823;
  assign n2469 = ~n2455 & ~n2468;
  assign n2470 = n9795 & ~n9796;
  assign n2471 = ~n9795 & n9796;
  assign n2472 = ~n2470 & ~n2471;
  assign n2473 = ~n2469 & ~n2472;
  assign n2474 = ~n2312 & ~n2327;
  assign n2475 = ~n2311 & n2331;
  assign n2476 = n2327 & ~n9805;
  assign n2477 = ~n2475 & ~n2476;
  assign n2478 = ~n9805 & ~n2474;
  assign n2479 = n9808 & ~n9809;
  assign n2480 = n9809 & ~n2372;
  assign n2481 = n9808 & n9809;
  assign n2482 = ~n9808 & ~n2372;
  assign n2483 = ~n9808 & ~n9809;
  assign n2484 = ~n9825 & ~n9826;
  assign n2485 = ~n2372 & ~n2479;
  assign n2486 = ~n9824 & ~n9827;
  assign n2487 = n9529 & ~n9624;
  assign n2488 = ~n225 & ~n9559;
  assign n2489 = n683 & n2488;
  assign n2490 = n1259 & n1479;
  assign n2491 = n2489 & n2490;
  assign n2492 = ~n215 & ~n9570;
  assign n2493 = ~n605 & n2492;
  assign n2494 = ~n215 & ~n605;
  assign n2495 = ~n9570 & n2494;
  assign n2496 = ~n215 & n707;
  assign n2497 = ~n9550 & ~n581;
  assign n2498 = ~n301 & n2497;
  assign n2499 = n9538 & n2498;
  assign n2500 = n9828 & n2499;
  assign n2501 = n9538 & n683;
  assign n2502 = n9828 & n2501;
  assign n2503 = n1479 & n2502;
  assign n2504 = n1259 & n2503;
  assign n2505 = ~n225 & n2504;
  assign n2506 = ~n581 & n2505;
  assign n2507 = ~n9550 & n2506;
  assign n2508 = ~n301 & n2507;
  assign n2509 = ~n9559 & n2508;
  assign n2510 = ~n225 & ~n581;
  assign n2511 = n683 & n2510;
  assign n2512 = n2490 & n2511;
  assign n2513 = ~n9550 & ~n9559;
  assign n2514 = ~n301 & n2513;
  assign n2515 = n9538 & n2514;
  assign n2516 = n9828 & n2515;
  assign n2517 = n2512 & n2516;
  assign n2518 = ~n301 & ~n581;
  assign n2519 = n683 & n2518;
  assign n2520 = n2490 & n2519;
  assign n2521 = ~n9550 & n2488;
  assign n2522 = n9538 & n2521;
  assign n2523 = n9828 & n2522;
  assign n2524 = n2520 & n2523;
  assign n2525 = n2491 & n2500;
  assign n2526 = ~n325 & ~n1083;
  assign n2527 = ~n265 & n2526;
  assign n2528 = ~n9562 & ~n754;
  assign n2529 = n1172 & n2528;
  assign n2530 = n1191 & n2529;
  assign n2531 = ~n325 & ~n9562;
  assign n2532 = ~n1083 & n2531;
  assign n2533 = n1172 & n1191;
  assign n2534 = n1672 & n2533;
  assign n2535 = n2532 & n2534;
  assign n2536 = ~n754 & ~n1083;
  assign n2537 = ~n1190 & n2536;
  assign n2538 = ~n265 & ~n325;
  assign n2539 = ~n9562 & ~n479;
  assign n2540 = n2538 & n2539;
  assign n2541 = n1172 & n2540;
  assign n2542 = n2537 & n2541;
  assign n2543 = n2527 & n2530;
  assign n2544 = n9610 & n9830;
  assign n2545 = ~n9541 & ~n384;
  assign n2546 = ~n995 & n2545;
  assign n2547 = ~n190 & ~n264;
  assign n2548 = ~n243 & ~n335;
  assign n2549 = ~n1037 & ~n1661;
  assign n2550 = n2548 & n2549;
  assign n2551 = n2547 & n2549;
  assign n2552 = n2548 & n2551;
  assign n2553 = n2547 & n2550;
  assign n2554 = ~n9541 & ~n1661;
  assign n2555 = ~n995 & n2554;
  assign n2556 = ~n335 & n2555;
  assign n2557 = ~n264 & n2556;
  assign n2558 = ~n190 & n2557;
  assign n2559 = ~n243 & n2558;
  assign n2560 = ~n1037 & n2559;
  assign n2561 = ~n384 & n2560;
  assign n2562 = ~n995 & ~n1037;
  assign n2563 = ~n1661 & n2562;
  assign n2564 = ~n264 & ~n384;
  assign n2565 = n2098 & n2564;
  assign n2566 = n2548 & n2565;
  assign n2567 = n2563 & n2566;
  assign n2568 = ~n9541 & ~n995;
  assign n2569 = ~n264 & n2568;
  assign n2570 = ~n335 & ~n384;
  assign n2571 = ~n243 & ~n1661;
  assign n2572 = ~n190 & ~n1037;
  assign n2573 = n2571 & n2572;
  assign n2574 = n2570 & n2573;
  assign n2575 = n2569 & n2574;
  assign n2576 = n2546 & n9831;
  assign n2577 = ~n192 & ~n328;
  assign n2578 = n1531 & n2577;
  assign n2579 = n758 & n1658;
  assign n2580 = n1840 & n2579;
  assign n2581 = ~n9561 & n758;
  assign n2582 = ~n328 & n2581;
  assign n2583 = ~n574 & n2582;
  assign n2584 = ~n554 & n2583;
  assign n2585 = ~n226 & n2584;
  assign n2586 = ~n192 & n2585;
  assign n2587 = ~n205 & n2586;
  assign n2588 = ~n294 & n2587;
  assign n2589 = n1840 & n2577;
  assign n2590 = n1531 & n2579;
  assign n2591 = n2589 & n2590;
  assign n2592 = ~n192 & ~n205;
  assign n2593 = n1658 & n2592;
  assign n2594 = ~n328 & ~n554;
  assign n2595 = n1531 & n2594;
  assign n2596 = n758 & n2595;
  assign n2597 = n2593 & n2596;
  assign n2598 = n2578 & n2580;
  assign n2599 = n9832 & n9833;
  assign n2600 = n2544 & n2599;
  assign n2601 = n1172 & n9832;
  assign n2602 = n9829 & n2601;
  assign n2603 = n9610 & n2602;
  assign n2604 = n9833 & n2603;
  assign n2605 = ~n325 & n2604;
  assign n2606 = ~n9562 & n2605;
  assign n2607 = ~n265 & n2606;
  assign n2608 = ~n1083 & n2607;
  assign n2609 = ~n754 & n2608;
  assign n2610 = ~n1190 & n2609;
  assign n2611 = ~n479 & n2610;
  assign n2612 = n9829 & n2600;
  assign n2613 = n9754 & ~n9834;
  assign n2614 = ~n9834 & ~n2613;
  assign n2615 = ~n9754 & ~n9834;
  assign n2616 = n1164 & ~n9754;
  assign n2617 = ~n1164 & n9834;
  assign n2618 = ~n9754 & ~n2617;
  assign n2619 = ~n9835 & ~n2616;
  assign n2620 = n2487 & n9836;
  assign n2621 = ~n2487 & ~n9836;
  assign n2622 = ~n2620 & ~n2621;
  assign n2623 = n9670 & n9810;
  assign n2624 = ~n9670 & n9802;
  assign n2625 = ~n2623 & ~n2624;
  assign n2626 = ~n1149 & n2324;
  assign n2627 = n1149 & n9811;
  assign n2628 = ~n2626 & ~n2627;
  assign n2629 = ~n2624 & n2628;
  assign n2630 = ~n2623 & n2629;
  assign n2631 = n2625 & n2628;
  assign n2632 = n2622 & n9837;
  assign n2633 = ~n2620 & ~n2632;
  assign n2634 = ~n9528 & n1142;
  assign n2635 = n9528 & n1137;
  assign n2636 = n9624 & n2130;
  assign n2637 = ~n2131 & ~n2636;
  assign n2638 = ~n9649 & n2130;
  assign n2639 = ~n9649 & ~n2637;
  assign n2640 = ~n2635 & ~n9838;
  assign n2641 = ~n2634 & ~n2635;
  assign n2642 = ~n9838 & n2641;
  assign n2643 = ~n2634 & n2640;
  assign n2644 = ~n2633 & n9839;
  assign n2645 = n2633 & ~n9839;
  assign n2646 = ~n2644 & ~n2645;
  assign n2647 = ~n9625 & n9674;
  assign n2648 = n9625 & n9728;
  assign n2649 = ~n2647 & ~n2648;
  assign n2650 = n9676 & ~n1703;
  assign n2651 = n1703 & n1726;
  assign n2652 = ~n2650 & ~n2651;
  assign n2653 = ~n2647 & n2652;
  assign n2654 = ~n2648 & n2653;
  assign n2655 = ~n2647 & ~n2650;
  assign n2656 = ~n2648 & ~n2651;
  assign n2657 = n2655 & n2656;
  assign n2658 = n2649 & n2652;
  assign n2659 = n9626 & n9787;
  assign n2660 = ~n9626 & n9772;
  assign n2661 = ~n2659 & ~n2660;
  assign n2662 = ~n978 & n2156;
  assign n2663 = n978 & n2245;
  assign n2664 = ~n2662 & ~n2663;
  assign n2665 = ~n2660 & n2664;
  assign n2666 = ~n2659 & n2665;
  assign n2667 = n2661 & n2664;
  assign n2668 = n9840 & n9841;
  assign n2669 = ~n9840 & ~n9841;
  assign n2670 = ~n9840 & n9841;
  assign n2671 = n9840 & ~n9841;
  assign n2672 = ~n2670 & ~n2671;
  assign n2673 = ~n2668 & ~n2669;
  assign n2674 = n9668 & n9686;
  assign n2675 = n9669 & ~n9686;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = n9671 & ~n2130;
  assign n2678 = n1304 & n2130;
  assign n2679 = ~n2677 & ~n2678;
  assign n2680 = ~n2675 & n2679;
  assign n2681 = ~n2674 & n2680;
  assign n2682 = n2676 & n2679;
  assign n2683 = ~n9842 & n9843;
  assign n2684 = ~n2668 & ~n2683;
  assign n2685 = n2646 & ~n2684;
  assign n2686 = ~n2644 & ~n2685;
  assign n2687 = n9824 & n9827;
  assign n2688 = ~n9824 & ~n2486;
  assign n2689 = ~n9824 & n9827;
  assign n2690 = ~n9827 & ~n2486;
  assign n2691 = n9824 & ~n9827;
  assign n2692 = ~n9844 & ~n9845;
  assign n2693 = ~n2486 & ~n2687;
  assign n2694 = ~n2686 & ~n9846;
  assign n2695 = ~n2486 & ~n2694;
  assign n2696 = n2331 & ~n2333;
  assign n2697 = ~n2334 & ~n2696;
  assign n2698 = ~n2695 & n2697;
  assign n2699 = n2695 & ~n2697;
  assign n2700 = ~n2698 & ~n2699;
  assign n2701 = n2450 & ~n2452;
  assign n2702 = ~n2453 & ~n2701;
  assign n2703 = n2700 & n2702;
  assign n2704 = ~n2698 & ~n2703;
  assign n2705 = n9820 & n9823;
  assign n2706 = ~n9823 & ~n2468;
  assign n2707 = n9820 & ~n9823;
  assign n2708 = ~n9820 & ~n2468;
  assign n2709 = ~n9820 & n9823;
  assign n2710 = ~n9847 & ~n9848;
  assign n2711 = ~n2468 & ~n2705;
  assign n2712 = ~n2704 & ~n9849;
  assign n2713 = ~n1164 & ~n9834;
  assign n2714 = n9754 & ~n2713;
  assign n2715 = ~n1164 & n9835;
  assign n2716 = n9670 & n9834;
  assign n2717 = ~n2715 & ~n2716;
  assign n2718 = n1164 & n2613;
  assign n2719 = ~n9670 & ~n9754;
  assign n2720 = n9834 & ~n2719;
  assign n2721 = ~n2718 & ~n2720;
  assign n2722 = ~n2715 & n2721;
  assign n2723 = ~n2714 & n2717;
  assign n2724 = ~n9624 & n9850;
  assign n2725 = n83 & n1142;
  assign n2726 = ~n83 & n1137;
  assign n2727 = ~n9528 & n9624;
  assign n2728 = ~n2309 & ~n2727;
  assign n2729 = ~n9528 & ~n9649;
  assign n2730 = ~n9649 & ~n2728;
  assign n2731 = ~n2726 & ~n9851;
  assign n2732 = ~n2725 & ~n2726;
  assign n2733 = ~n9851 & n2732;
  assign n2734 = ~n2725 & n2731;
  assign n2735 = n2724 & n9852;
  assign n2736 = n9674 & n1703;
  assign n2737 = ~n1703 & n9728;
  assign n2738 = ~n2736 & ~n2737;
  assign n2739 = n9676 & n9686;
  assign n2740 = ~n9686 & n1726;
  assign n2741 = ~n2739 & ~n2740;
  assign n2742 = ~n2736 & n2741;
  assign n2743 = ~n2737 & n2742;
  assign n2744 = ~n2736 & ~n2739;
  assign n2745 = ~n2737 & ~n2740;
  assign n2746 = n2744 & n2745;
  assign n2747 = n2738 & n2741;
  assign n2748 = n9668 & ~n2130;
  assign n2749 = n9669 & n2130;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = n9528 & n9671;
  assign n2752 = ~n9528 & n1304;
  assign n2753 = ~n2751 & ~n2752;
  assign n2754 = ~n2749 & n2753;
  assign n2755 = ~n2748 & n2754;
  assign n2756 = n2750 & n2753;
  assign n2757 = n9853 & n9854;
  assign n2758 = ~n9853 & ~n9854;
  assign n2759 = n9853 & ~n9854;
  assign n2760 = ~n9853 & n9854;
  assign n2761 = ~n2759 & ~n2760;
  assign n2762 = ~n2757 & ~n2758;
  assign n2763 = ~n978 & n9787;
  assign n2764 = n978 & n9772;
  assign n2765 = ~n2763 & ~n2764;
  assign n2766 = n9625 & n2156;
  assign n2767 = ~n9625 & n2245;
  assign n2768 = ~n2766 & ~n2767;
  assign n2769 = ~n2764 & n2768;
  assign n2770 = ~n2763 & n2769;
  assign n2771 = n2765 & n2768;
  assign n2772 = ~n9855 & n9856;
  assign n2773 = ~n2757 & ~n2772;
  assign n2774 = ~n2724 & ~n9852;
  assign n2775 = ~n2735 & ~n2774;
  assign n2776 = ~n2773 & n2775;
  assign n2777 = ~n2735 & ~n2776;
  assign n2778 = ~n2380 & ~n9812;
  assign n2779 = ~n2379 & n2397;
  assign n2780 = n9812 & ~n9813;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = ~n9813 & ~n2778;
  assign n2783 = ~n2777 & ~n9857;
  assign n2784 = n2777 & n9857;
  assign n2785 = n2777 & ~n9857;
  assign n2786 = ~n2777 & n9857;
  assign n2787 = ~n2785 & ~n2786;
  assign n2788 = ~n2783 & ~n2784;
  assign n2789 = n9818 & ~n9819;
  assign n2790 = n9819 & ~n2447;
  assign n2791 = n9818 & n9819;
  assign n2792 = ~n9818 & ~n2447;
  assign n2793 = ~n9818 & ~n9819;
  assign n2794 = ~n9859 & ~n9860;
  assign n2795 = ~n2447 & ~n2789;
  assign n2796 = ~n9858 & ~n9861;
  assign n2797 = ~n2783 & ~n2796;
  assign n2798 = ~n2410 & n2448;
  assign n2799 = ~n2449 & ~n2798;
  assign n2800 = ~n2797 & n2799;
  assign n2801 = n2797 & ~n2799;
  assign n2802 = ~n2800 & ~n2801;
  assign n2803 = n2686 & n9846;
  assign n2804 = ~n2686 & n9846;
  assign n2805 = n2686 & ~n9846;
  assign n2806 = ~n2804 & ~n2805;
  assign n2807 = ~n2694 & ~n2803;
  assign n2808 = n2802 & ~n9862;
  assign n2809 = ~n2800 & ~n2808;
  assign n2810 = ~n2700 & ~n2702;
  assign n2811 = ~n2703 & ~n2810;
  assign n2812 = ~n2809 & n2811;
  assign n2813 = ~n2646 & n2684;
  assign n2814 = ~n2685 & ~n2813;
  assign n2815 = ~n9529 & n1142;
  assign n2816 = n9529 & n1137;
  assign n2817 = n83 & n9624;
  assign n2818 = ~n2377 & ~n2817;
  assign n2819 = n83 & ~n9649;
  assign n2820 = ~n9649 & ~n2818;
  assign n2821 = ~n2816 & ~n9863;
  assign n2822 = ~n2815 & ~n2816;
  assign n2823 = ~n9863 & n2822;
  assign n2824 = ~n2815 & n2821;
  assign n2825 = ~n1149 & n9810;
  assign n2826 = n1149 & n9802;
  assign n2827 = ~n2825 & ~n2826;
  assign n2828 = n9626 & n2324;
  assign n2829 = ~n9626 & n9811;
  assign n2830 = ~n2828 & ~n2829;
  assign n2831 = ~n2826 & n2830;
  assign n2832 = ~n2825 & n2831;
  assign n2833 = n2827 & n2830;
  assign n2834 = n9864 & n9865;
  assign n2835 = n9624 & ~n9850;
  assign n2836 = ~n2724 & ~n2835;
  assign n2837 = ~n9864 & ~n9865;
  assign n2838 = ~n2834 & ~n2837;
  assign n2839 = ~n2834 & n2836;
  assign n2840 = ~n2837 & n2839;
  assign n2841 = n2836 & n2838;
  assign n2842 = ~n2834 & ~n9866;
  assign n2843 = ~n2622 & ~n9837;
  assign n2844 = ~n2632 & ~n2843;
  assign n2845 = n2842 & ~n2844;
  assign n2846 = ~n2842 & n2844;
  assign n2847 = n9842 & ~n9843;
  assign n2848 = n9843 & ~n2683;
  assign n2849 = n9842 & n9843;
  assign n2850 = ~n9842 & ~n2683;
  assign n2851 = ~n9842 & ~n9843;
  assign n2852 = ~n9867 & ~n9868;
  assign n2853 = ~n2683 & ~n2847;
  assign n2854 = ~n2846 & n9869;
  assign n2855 = ~n2845 & ~n9869;
  assign n2856 = ~n2846 & ~n2855;
  assign n2857 = ~n2845 & ~n2846;
  assign n2858 = ~n9869 & n2857;
  assign n2859 = ~n2846 & ~n2858;
  assign n2860 = ~n2845 & ~n2854;
  assign n2861 = n2814 & ~n9870;
  assign n2862 = ~n2814 & n9870;
  assign n2863 = ~n2861 & ~n2862;
  assign n2864 = n9858 & n9861;
  assign n2865 = ~n2796 & ~n2864;
  assign n2866 = n2863 & n2865;
  assign n2867 = ~n2861 & ~n2866;
  assign n2868 = ~n2802 & n9862;
  assign n2869 = ~n2808 & ~n2868;
  assign n2870 = ~n2867 & n2869;
  assign n2871 = n9625 & n9787;
  assign n2872 = ~n9625 & n9772;
  assign n2873 = ~n2871 & ~n2872;
  assign n2874 = ~n1703 & n2156;
  assign n2875 = n1703 & n2245;
  assign n2876 = ~n2874 & ~n2875;
  assign n2877 = ~n2872 & n2876;
  assign n2878 = ~n2871 & n2877;
  assign n2879 = n2873 & n2876;
  assign n2880 = n9674 & ~n9686;
  assign n2881 = n9686 & n9728;
  assign n2882 = ~n2880 & ~n2881;
  assign n2883 = n9676 & ~n2130;
  assign n2884 = n1726 & n2130;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = ~n2880 & n2885;
  assign n2887 = ~n2881 & n2886;
  assign n2888 = ~n2880 & ~n2883;
  assign n2889 = ~n2881 & ~n2884;
  assign n2890 = n2888 & n2889;
  assign n2891 = n2882 & n2885;
  assign n2892 = n9871 & n9872;
  assign n2893 = n9529 & ~n9667;
  assign n2894 = n9529 & n9668;
  assign n2895 = ~n9529 & ~n1289;
  assign n2896 = ~n1304 & ~n2895;
  assign n2897 = ~n2894 & n2896;
  assign n2898 = n1289 & n2897;
  assign n2899 = n1289 & ~n2894;
  assign n2900 = n1289 & ~n2893;
  assign n2901 = ~n1149 & ~n9834;
  assign n2902 = n9754 & ~n2901;
  assign n2903 = ~n1149 & n9835;
  assign n2904 = n9626 & n9834;
  assign n2905 = ~n2903 & ~n2904;
  assign n2906 = n1149 & n2613;
  assign n2907 = ~n9626 & ~n9754;
  assign n2908 = n9834 & ~n2907;
  assign n2909 = ~n2906 & ~n2908;
  assign n2910 = ~n2903 & n2909;
  assign n2911 = ~n2902 & n2905;
  assign n2912 = n9873 & n9874;
  assign n2913 = ~n9871 & ~n9872;
  assign n2914 = n9871 & ~n9872;
  assign n2915 = ~n9871 & n9872;
  assign n2916 = ~n2914 & ~n2915;
  assign n2917 = ~n2892 & ~n2913;
  assign n2918 = n2912 & ~n9875;
  assign n2919 = ~n2892 & ~n2918;
  assign n2920 = n9670 & ~n9834;
  assign n2921 = n9754 & ~n2920;
  assign n2922 = n9670 & n9835;
  assign n2923 = ~n1149 & n9834;
  assign n2924 = ~n2922 & ~n2923;
  assign n2925 = ~n9670 & n2613;
  assign n2926 = n1149 & ~n9754;
  assign n2927 = n9834 & ~n2926;
  assign n2928 = ~n2925 & ~n2927;
  assign n2929 = ~n2922 & n2928;
  assign n2930 = ~n2921 & n2924;
  assign n2931 = n9626 & n9810;
  assign n2932 = ~n9626 & n9802;
  assign n2933 = ~n2931 & ~n2932;
  assign n2934 = ~n978 & n2324;
  assign n2935 = n978 & n9811;
  assign n2936 = ~n2934 & ~n2935;
  assign n2937 = ~n2932 & n2936;
  assign n2938 = ~n2931 & n2937;
  assign n2939 = n2933 & n2936;
  assign n2940 = n9876 & n9877;
  assign n2941 = ~n9876 & ~n9877;
  assign n2942 = n9876 & ~n9877;
  assign n2943 = ~n9876 & n9877;
  assign n2944 = ~n2942 & ~n2943;
  assign n2945 = ~n2940 & ~n2941;
  assign n2946 = n9528 & n9668;
  assign n2947 = ~n9528 & n9669;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = ~n83 & n9671;
  assign n2950 = n83 & n1304;
  assign n2951 = ~n2949 & ~n2950;
  assign n2952 = ~n2947 & n2951;
  assign n2953 = ~n2946 & n2952;
  assign n2954 = n2948 & n2951;
  assign n2955 = ~n9878 & n9879;
  assign n2956 = ~n2940 & ~n2955;
  assign n2957 = ~n2919 & ~n2956;
  assign n2958 = n2919 & n2956;
  assign n2959 = ~n2919 & ~n2957;
  assign n2960 = ~n2919 & n2956;
  assign n2961 = ~n2956 & ~n2957;
  assign n2962 = n2919 & ~n2956;
  assign n2963 = ~n9880 & ~n9881;
  assign n2964 = ~n2957 & ~n2958;
  assign n2965 = n9855 & ~n9856;
  assign n2966 = n9856 & ~n2772;
  assign n2967 = n9855 & n9856;
  assign n2968 = ~n9855 & ~n2772;
  assign n2969 = ~n9855 & ~n9856;
  assign n2970 = ~n9883 & ~n9884;
  assign n2971 = ~n2772 & ~n2965;
  assign n2972 = ~n9882 & ~n9885;
  assign n2973 = ~n2957 & ~n2972;
  assign n2974 = n2773 & ~n2775;
  assign n2975 = ~n2776 & ~n2974;
  assign n2976 = ~n2973 & n2975;
  assign n2977 = n2973 & ~n2975;
  assign n2978 = ~n2976 & ~n2977;
  assign n2979 = n9869 & ~n2857;
  assign n2980 = n2857 & ~n2858;
  assign n2981 = ~n9869 & ~n2858;
  assign n2982 = ~n2980 & ~n2981;
  assign n2983 = ~n2858 & ~n2979;
  assign n2984 = n2978 & ~n9886;
  assign n2985 = ~n2976 & ~n2984;
  assign n2986 = ~n2863 & ~n2865;
  assign n2987 = ~n2866 & ~n2986;
  assign n2988 = ~n2985 & n2987;
  assign n2989 = ~n9529 & n9624;
  assign n2990 = ~n1142 & ~n2989;
  assign n2991 = n9624 & n2990;
  assign n2992 = n9529 & ~n9649;
  assign n2993 = ~n978 & n9810;
  assign n2994 = n978 & n9802;
  assign n2995 = ~n2993 & ~n2994;
  assign n2996 = n9625 & n2324;
  assign n2997 = ~n9625 & n9811;
  assign n2998 = ~n2996 & ~n2997;
  assign n2999 = ~n2994 & n2998;
  assign n3000 = ~n2993 & n2999;
  assign n3001 = n2995 & n2998;
  assign n3002 = n9674 & n2130;
  assign n3003 = n9728 & ~n2130;
  assign n3004 = ~n3002 & ~n3003;
  assign n3005 = n9528 & n9676;
  assign n3006 = ~n9528 & n1726;
  assign n3007 = ~n3005 & ~n3006;
  assign n3008 = ~n3002 & n3007;
  assign n3009 = ~n3003 & n3008;
  assign n3010 = ~n3002 & ~n3005;
  assign n3011 = ~n3003 & ~n3006;
  assign n3012 = n3010 & n3011;
  assign n3013 = n3004 & n3007;
  assign n3014 = n9888 & n9889;
  assign n3015 = ~n9888 & ~n9889;
  assign n3016 = n9888 & ~n9889;
  assign n3017 = ~n9888 & n9889;
  assign n3018 = ~n3016 & ~n3017;
  assign n3019 = ~n3014 & ~n3015;
  assign n3020 = ~n1703 & n9787;
  assign n3021 = n1703 & n9772;
  assign n3022 = ~n3020 & ~n3021;
  assign n3023 = n9686 & n2156;
  assign n3024 = ~n9686 & n2245;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = ~n3021 & n3025;
  assign n3027 = ~n3020 & n3026;
  assign n3028 = n3022 & n3025;
  assign n3029 = ~n9890 & n9891;
  assign n3030 = ~n3014 & ~n3029;
  assign n3031 = n9624 & ~n3030;
  assign n3032 = n2990 & n3031;
  assign n3033 = n9887 & ~n3030;
  assign n3034 = ~n2912 & n9875;
  assign n3035 = ~n2918 & ~n3034;
  assign n3036 = ~n9887 & n3030;
  assign n3037 = n9624 & ~n9892;
  assign n3038 = n2990 & n3037;
  assign n3039 = n9887 & ~n9892;
  assign n3040 = ~n3030 & ~n9892;
  assign n3041 = ~n9893 & ~n3040;
  assign n3042 = ~n9892 & ~n3036;
  assign n3043 = n3035 & ~n9894;
  assign n3044 = ~n9892 & ~n3043;
  assign n3045 = ~n2836 & ~n2838;
  assign n3046 = n2836 & ~n9866;
  assign n3047 = n2836 & ~n2838;
  assign n3048 = ~n2837 & n2842;
  assign n3049 = ~n2836 & n2838;
  assign n3050 = ~n9895 & ~n9896;
  assign n3051 = ~n9866 & ~n3045;
  assign n3052 = ~n3044 & ~n9897;
  assign n3053 = n9882 & n9885;
  assign n3054 = ~n9882 & ~n2972;
  assign n3055 = ~n9885 & ~n2972;
  assign n3056 = ~n3054 & ~n3055;
  assign n3057 = ~n2972 & ~n3053;
  assign n3058 = n3044 & n9897;
  assign n3059 = ~n3044 & n9897;
  assign n3060 = n3044 & ~n9897;
  assign n3061 = ~n3059 & ~n3060;
  assign n3062 = ~n3052 & ~n3058;
  assign n3063 = ~n9898 & ~n9899;
  assign n3064 = ~n3052 & ~n3063;
  assign n3065 = ~n2978 & n9886;
  assign n3066 = ~n2984 & ~n3065;
  assign n3067 = ~n3064 & n3066;
  assign n3068 = n3064 & ~n3066;
  assign n3069 = ~n3067 & ~n3068;
  assign n3070 = n9898 & n9899;
  assign n3071 = ~n3063 & ~n3070;
  assign n3072 = ~n3035 & n9894;
  assign n3073 = ~n9894 & ~n3043;
  assign n3074 = n3035 & ~n3043;
  assign n3075 = ~n3073 & ~n3074;
  assign n3076 = ~n3043 & ~n3072;
  assign n3077 = ~n9873 & ~n9874;
  assign n3078 = ~n2912 & ~n3077;
  assign n3079 = ~n83 & n9668;
  assign n3080 = n83 & n9669;
  assign n3081 = ~n3079 & ~n3080;
  assign n3082 = n9529 & n9671;
  assign n3083 = ~n9529 & n1304;
  assign n3084 = ~n3082 & ~n3083;
  assign n3085 = ~n3080 & n3084;
  assign n3086 = ~n3079 & n3085;
  assign n3087 = n3081 & n3084;
  assign n3088 = n3078 & n9901;
  assign n3089 = n9626 & ~n9834;
  assign n3090 = n9754 & ~n3089;
  assign n3091 = n9626 & n9835;
  assign n3092 = ~n978 & n9834;
  assign n3093 = ~n3091 & ~n3092;
  assign n3094 = ~n9626 & n2613;
  assign n3095 = n978 & ~n9754;
  assign n3096 = n9834 & ~n3095;
  assign n3097 = ~n3094 & ~n3096;
  assign n3098 = ~n3091 & n3097;
  assign n3099 = ~n3090 & n3093;
  assign n3100 = n9625 & n9810;
  assign n3101 = ~n9625 & n9802;
  assign n3102 = ~n3100 & ~n3101;
  assign n3103 = ~n1703 & n2324;
  assign n3104 = n1703 & n9811;
  assign n3105 = ~n3103 & ~n3104;
  assign n3106 = ~n3101 & n3105;
  assign n3107 = ~n3100 & n3106;
  assign n3108 = n3102 & n3105;
  assign n3109 = n9902 & n9903;
  assign n3110 = ~n9902 & ~n9903;
  assign n3111 = n9902 & ~n9903;
  assign n3112 = ~n9902 & n9903;
  assign n3113 = ~n3111 & ~n3112;
  assign n3114 = ~n3109 & ~n3110;
  assign n3115 = n9686 & n9787;
  assign n3116 = ~n9686 & n9772;
  assign n3117 = ~n3115 & ~n3116;
  assign n3118 = ~n2130 & n2156;
  assign n3119 = n2130 & n2245;
  assign n3120 = ~n3118 & ~n3119;
  assign n3121 = ~n3116 & n3120;
  assign n3122 = ~n3115 & n3121;
  assign n3123 = n3117 & n3120;
  assign n3124 = ~n9904 & n9905;
  assign n3125 = ~n3109 & ~n3124;
  assign n3126 = ~n3078 & ~n9901;
  assign n3127 = ~n3078 & n9901;
  assign n3128 = n3078 & ~n9901;
  assign n3129 = ~n3127 & ~n3128;
  assign n3130 = ~n3088 & ~n3126;
  assign n3131 = ~n3125 & ~n9906;
  assign n3132 = ~n3088 & ~n3131;
  assign n3133 = n9878 & ~n9879;
  assign n3134 = n9879 & ~n2955;
  assign n3135 = n9878 & n9879;
  assign n3136 = ~n9878 & ~n2955;
  assign n3137 = ~n9878 & ~n9879;
  assign n3138 = ~n9907 & ~n9908;
  assign n3139 = ~n2955 & ~n3133;
  assign n3140 = ~n3132 & ~n9909;
  assign n3141 = n3132 & n9909;
  assign n3142 = ~n3132 & ~n3140;
  assign n3143 = ~n9909 & ~n3140;
  assign n3144 = ~n3142 & ~n3143;
  assign n3145 = ~n3140 & ~n3141;
  assign n3146 = ~n9900 & ~n9910;
  assign n3147 = n9900 & n9910;
  assign n3148 = ~n3146 & ~n3147;
  assign n3149 = n9529 & ~n9673;
  assign n3150 = n9529 & n9728;
  assign n3151 = ~n9529 & ~n821;
  assign n3152 = ~n1726 & ~n3151;
  assign n3153 = ~n3150 & n3152;
  assign n3154 = n821 & n3153;
  assign n3155 = n821 & ~n3149;
  assign n3156 = ~n978 & ~n9834;
  assign n3157 = n9754 & ~n3156;
  assign n3158 = ~n978 & n9835;
  assign n3159 = n9625 & n9834;
  assign n3160 = ~n3158 & ~n3159;
  assign n3161 = n978 & n2613;
  assign n3162 = ~n9625 & ~n9754;
  assign n3163 = n9834 & ~n3162;
  assign n3164 = ~n3161 & ~n3163;
  assign n3165 = ~n3158 & n3164;
  assign n3166 = ~n3157 & n3160;
  assign n3167 = n9911 & n9912;
  assign n3168 = ~n9528 & n9674;
  assign n3169 = n9528 & n9728;
  assign n3170 = ~n3168 & ~n3169;
  assign n3171 = ~n83 & n9676;
  assign n3172 = n83 & n1726;
  assign n3173 = ~n3171 & ~n3172;
  assign n3174 = ~n3168 & n3173;
  assign n3175 = ~n3169 & n3174;
  assign n3176 = ~n3168 & ~n3171;
  assign n3177 = ~n3169 & ~n3172;
  assign n3178 = n3176 & n3177;
  assign n3179 = n3170 & n3173;
  assign n3180 = n3167 & n9913;
  assign n3181 = ~n3167 & ~n9913;
  assign n3182 = n3167 & ~n9913;
  assign n3183 = ~n3167 & n9913;
  assign n3184 = ~n3182 & ~n3183;
  assign n3185 = ~n3180 & ~n3181;
  assign n3186 = n2893 & ~n9914;
  assign n3187 = ~n3180 & ~n3186;
  assign n3188 = n9890 & ~n9891;
  assign n3189 = ~n3029 & ~n3188;
  assign n3190 = ~n3187 & n3189;
  assign n3191 = n3187 & ~n3189;
  assign n3192 = ~n3190 & ~n3191;
  assign n3193 = n3125 & n9906;
  assign n3194 = ~n3131 & ~n3193;
  assign n3195 = n3192 & n3194;
  assign n3196 = ~n3192 & ~n3194;
  assign n3197 = ~n3195 & ~n3196;
  assign n3198 = n9686 & ~n9834;
  assign n3199 = n9754 & ~n3198;
  assign n3200 = n9686 & n9835;
  assign n3201 = ~n2130 & n9834;
  assign n3202 = ~n3200 & ~n3201;
  assign n3203 = ~n9686 & n2613;
  assign n3204 = ~n9754 & n2130;
  assign n3205 = n9834 & ~n3204;
  assign n3206 = ~n3203 & ~n3205;
  assign n3207 = ~n3200 & n3206;
  assign n3208 = ~n3199 & n3202;
  assign n3209 = n9528 & n9810;
  assign n3210 = ~n9528 & n9802;
  assign n3211 = ~n3209 & ~n3210;
  assign n3212 = ~n83 & n2324;
  assign n3213 = n83 & n9811;
  assign n3214 = ~n3212 & ~n3213;
  assign n3215 = ~n3210 & n3214;
  assign n3216 = ~n3209 & n3215;
  assign n3217 = n3211 & n3214;
  assign n3218 = n9915 & n9916;
  assign n3219 = n9529 & ~n9801;
  assign n3220 = n9529 & n9810;
  assign n3221 = ~n9529 & ~n2124;
  assign n3222 = ~n9811 & ~n3221;
  assign n3223 = ~n3220 & n3222;
  assign n3224 = n2124 & n3223;
  assign n3225 = n2124 & ~n3219;
  assign n3226 = ~n2130 & ~n9834;
  assign n3227 = n9754 & ~n3226;
  assign n3228 = ~n2130 & n9835;
  assign n3229 = n9528 & n9834;
  assign n3230 = ~n3228 & ~n3229;
  assign n3231 = n2130 & n2613;
  assign n3232 = ~n9528 & ~n9754;
  assign n3233 = n9834 & ~n3232;
  assign n3234 = ~n3231 & ~n3233;
  assign n3235 = ~n3228 & n3234;
  assign n3236 = ~n3227 & n3230;
  assign n3237 = n9917 & n9918;
  assign n3238 = ~n9915 & ~n9916;
  assign n3239 = n9915 & ~n9916;
  assign n3240 = ~n9915 & n9916;
  assign n3241 = ~n3239 & ~n3240;
  assign n3242 = ~n3218 & ~n3238;
  assign n3243 = n3237 & ~n9919;
  assign n3244 = ~n3218 & ~n3243;
  assign n3245 = n9529 & ~n9771;
  assign n3246 = n9529 & n9787;
  assign n3247 = ~n9529 & ~n1696;
  assign n3248 = ~n2245 & ~n3247;
  assign n3249 = ~n3246 & n3248;
  assign n3250 = n1696 & n3249;
  assign n3251 = n1696 & ~n3246;
  assign n3252 = n1696 & ~n3245;
  assign n3253 = ~n1703 & ~n9834;
  assign n3254 = n9754 & ~n3253;
  assign n3255 = ~n1703 & n9835;
  assign n3256 = n9686 & n9834;
  assign n3257 = ~n3255 & ~n3256;
  assign n3258 = n1703 & n2613;
  assign n3259 = ~n9686 & ~n9754;
  assign n3260 = n9834 & ~n3259;
  assign n3261 = ~n3258 & ~n3260;
  assign n3262 = ~n3255 & n3261;
  assign n3263 = ~n3254 & n3257;
  assign n3264 = n9920 & n9921;
  assign n3265 = ~n9920 & ~n9921;
  assign n3266 = ~n3264 & ~n3265;
  assign n3267 = ~n2130 & n9810;
  assign n3268 = n2130 & n9802;
  assign n3269 = ~n3267 & ~n3268;
  assign n3270 = ~n9528 & n9811;
  assign n3271 = n9528 & n2324;
  assign n3272 = ~n3270 & ~n3271;
  assign n3273 = ~n3268 & n3272;
  assign n3274 = ~n3267 & n3273;
  assign n3275 = n3269 & n3272;
  assign n3276 = ~n83 & n9787;
  assign n3277 = n83 & n9772;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = ~n9529 & n2245;
  assign n3280 = n9529 & n2156;
  assign n3281 = ~n3279 & ~n3280;
  assign n3282 = ~n3277 & n3281;
  assign n3283 = ~n3276 & n3282;
  assign n3284 = n3278 & n3281;
  assign n3285 = n9922 & n9923;
  assign n3286 = ~n9922 & ~n9923;
  assign n3287 = ~n3285 & ~n3286;
  assign n3288 = n3266 & ~n3285;
  assign n3289 = ~n3286 & n3288;
  assign n3290 = n3266 & n3287;
  assign n3291 = ~n3266 & ~n3287;
  assign n3292 = n3266 & ~n9924;
  assign n3293 = n3266 & ~n3287;
  assign n3294 = ~n3285 & ~n9924;
  assign n3295 = ~n3286 & n3294;
  assign n3296 = ~n3266 & n3287;
  assign n3297 = ~n9925 & ~n9926;
  assign n3298 = ~n9924 & ~n3291;
  assign n3299 = n3244 & n9927;
  assign n3300 = ~n3237 & n9919;
  assign n3301 = ~n3243 & ~n3300;
  assign n3302 = ~n83 & n9810;
  assign n3303 = n83 & n9802;
  assign n3304 = ~n3302 & ~n3303;
  assign n3305 = n9529 & n2324;
  assign n3306 = ~n9529 & n9811;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = n3304 & n3307;
  assign n3309 = ~n9917 & ~n9918;
  assign n3310 = ~n3237 & ~n3309;
  assign n3311 = ~n83 & ~n9834;
  assign n3312 = ~n9529 & ~n9754;
  assign n3313 = ~n3311 & n3312;
  assign n3314 = ~n3219 & ~n3313;
  assign n3315 = n9528 & ~n9834;
  assign n3316 = n9754 & ~n3315;
  assign n3317 = n9528 & n9835;
  assign n3318 = ~n83 & n9834;
  assign n3319 = ~n3317 & ~n3318;
  assign n3320 = n9754 & n9834;
  assign n3321 = n83 & ~n3320;
  assign n3322 = ~n3311 & ~n3321;
  assign n3323 = ~n9528 & n2613;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = ~n3317 & n3324;
  assign n3326 = ~n3317 & ~n3323;
  assign n3327 = ~n3322 & n3326;
  assign n3328 = ~n3316 & n3319;
  assign n3329 = ~n3313 & ~n9928;
  assign n3330 = ~n9917 & ~n3329;
  assign n3331 = n3222 & n3330;
  assign n3332 = n3219 & n9928;
  assign n3333 = ~n3313 & ~n9929;
  assign n3334 = ~n3219 & ~n9928;
  assign n3335 = ~n3333 & ~n3334;
  assign n3336 = n3313 & n9928;
  assign n3337 = ~n9929 & ~n3336;
  assign n3338 = ~n3314 & n9928;
  assign n3339 = n3310 & n9930;
  assign n3340 = ~n3308 & ~n3339;
  assign n3341 = ~n3310 & ~n9930;
  assign n3342 = n3308 & n3310;
  assign n3343 = ~n9930 & ~n3342;
  assign n3344 = ~n3308 & ~n3310;
  assign n3345 = ~n3343 & ~n3344;
  assign n3346 = ~n3306 & ~n3341;
  assign n3347 = ~n3305 & n3346;
  assign n3348 = ~n3303 & n3347;
  assign n3349 = ~n3302 & n3348;
  assign n3350 = n3308 & ~n3341;
  assign n3351 = ~n3339 & ~n9932;
  assign n3352 = ~n3340 & ~n3341;
  assign n3353 = n3245 & n9931;
  assign n3354 = ~n3301 & ~n3353;
  assign n3355 = ~n3245 & ~n9931;
  assign n3356 = ~n3243 & ~n3355;
  assign n3357 = ~n3300 & n3356;
  assign n3358 = n3301 & ~n3355;
  assign n3359 = ~n3353 & ~n9933;
  assign n3360 = ~n3354 & ~n3355;
  assign n3361 = n3245 & n3301;
  assign n3362 = ~n9931 & ~n3361;
  assign n3363 = ~n3245 & ~n3301;
  assign n3364 = ~n3299 & ~n3363;
  assign n3365 = ~n3362 & n3364;
  assign n3366 = ~n3299 & ~n9934;
  assign n3367 = ~n9911 & n3264;
  assign n3368 = n3152 & n3367;
  assign n3369 = n3149 & n3264;
  assign n3370 = ~n3149 & ~n3264;
  assign n3371 = n3264 & ~n9936;
  assign n3372 = ~n3149 & n3264;
  assign n3373 = n3149 & ~n9936;
  assign n3374 = ~n9911 & ~n9936;
  assign n3375 = n3152 & n3374;
  assign n3376 = n3149 & ~n3264;
  assign n3377 = ~n9937 & ~n9938;
  assign n3378 = ~n9936 & ~n3370;
  assign n3379 = ~n3294 & ~n9939;
  assign n3380 = n3294 & n9939;
  assign n3381 = ~n3294 & ~n3379;
  assign n3382 = ~n9939 & ~n3379;
  assign n3383 = ~n3381 & ~n3382;
  assign n3384 = ~n3379 & ~n3380;
  assign n3385 = n9625 & ~n9834;
  assign n3386 = n9754 & ~n3385;
  assign n3387 = n9625 & n9835;
  assign n3388 = ~n1703 & n9834;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = ~n9625 & n2613;
  assign n3391 = n1703 & ~n9754;
  assign n3392 = n9834 & ~n3391;
  assign n3393 = ~n3390 & ~n3392;
  assign n3394 = ~n3387 & n3393;
  assign n3395 = ~n3386 & n3389;
  assign n3396 = n9686 & n9810;
  assign n3397 = ~n9686 & n9802;
  assign n3398 = ~n3396 & ~n3397;
  assign n3399 = ~n2130 & n2324;
  assign n3400 = n2130 & n9811;
  assign n3401 = ~n3399 & ~n3400;
  assign n3402 = ~n3397 & n3401;
  assign n3403 = ~n3396 & n3402;
  assign n3404 = n3398 & n3401;
  assign n3405 = n9941 & n9942;
  assign n3406 = ~n9941 & ~n9942;
  assign n3407 = n9941 & ~n9942;
  assign n3408 = ~n9941 & n9942;
  assign n3409 = ~n3407 & ~n3408;
  assign n3410 = ~n3405 & ~n3406;
  assign n3411 = n9528 & n9787;
  assign n3412 = ~n9528 & n9772;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = ~n83 & n2156;
  assign n3415 = n83 & n2245;
  assign n3416 = ~n3414 & ~n3415;
  assign n3417 = ~n3412 & n3416;
  assign n3418 = ~n3411 & n3417;
  assign n3419 = n3413 & n3416;
  assign n3420 = ~n9943 & n9944;
  assign n3421 = n9943 & ~n9944;
  assign n3422 = ~n3420 & ~n3421;
  assign n3423 = ~n9940 & n3422;
  assign n3424 = ~n3244 & ~n9927;
  assign n3425 = ~n3423 & ~n3424;
  assign n3426 = n9934 & ~n3424;
  assign n3427 = n9927 & n9934;
  assign n3428 = ~n3244 & ~n3427;
  assign n3429 = ~n9927 & ~n9934;
  assign n3430 = ~n3428 & ~n3429;
  assign n3431 = ~n3299 & ~n3426;
  assign n3432 = ~n3423 & n9945;
  assign n3433 = ~n9935 & n3425;
  assign n3434 = ~n9911 & ~n9912;
  assign n3435 = ~n3167 & ~n3434;
  assign n3436 = ~n3405 & ~n3420;
  assign n3437 = n3435 & ~n3436;
  assign n3438 = ~n3435 & n3436;
  assign n3439 = ~n3437 & ~n3438;
  assign n3440 = ~n1703 & n9810;
  assign n3441 = n1703 & n9802;
  assign n3442 = ~n3440 & ~n3441;
  assign n3443 = n9686 & n2324;
  assign n3444 = ~n9686 & n9811;
  assign n3445 = ~n3443 & ~n3444;
  assign n3446 = ~n3441 & n3445;
  assign n3447 = ~n3440 & n3446;
  assign n3448 = n3442 & n3445;
  assign n3449 = ~n2130 & n9787;
  assign n3450 = n2130 & n9772;
  assign n3451 = ~n3449 & ~n3450;
  assign n3452 = n9528 & n2156;
  assign n3453 = ~n9528 & n2245;
  assign n3454 = ~n3452 & ~n3453;
  assign n3455 = ~n3450 & n3454;
  assign n3456 = ~n3449 & n3455;
  assign n3457 = n3451 & n3454;
  assign n3458 = n9947 & n9948;
  assign n3459 = ~n9947 & ~n9948;
  assign n3460 = n9947 & ~n9948;
  assign n3461 = ~n9947 & n9948;
  assign n3462 = ~n3460 & ~n3461;
  assign n3463 = ~n3458 & ~n3459;
  assign n3464 = n83 & n9674;
  assign n3465 = ~n83 & n9728;
  assign n3466 = ~n3464 & ~n3465;
  assign n3467 = n9529 & n9676;
  assign n3468 = ~n9529 & n1726;
  assign n3469 = ~n3467 & ~n3468;
  assign n3470 = ~n3464 & n3469;
  assign n3471 = ~n3465 & n3470;
  assign n3472 = ~n3465 & ~n3467;
  assign n3473 = ~n3464 & ~n3468;
  assign n3474 = n3472 & n3473;
  assign n3475 = n3466 & n3469;
  assign n3476 = ~n9949 & n9950;
  assign n3477 = n9949 & ~n9950;
  assign n3478 = n9950 & ~n3476;
  assign n3479 = n9949 & n9950;
  assign n3480 = ~n9949 & ~n3476;
  assign n3481 = ~n9949 & ~n9950;
  assign n3482 = ~n9951 & ~n9952;
  assign n3483 = ~n3476 & ~n3477;
  assign n3484 = n3439 & ~n9953;
  assign n3485 = ~n3439 & n9953;
  assign n3486 = ~n3484 & ~n3485;
  assign n3487 = ~n9936 & ~n3379;
  assign n3488 = ~n3486 & n3487;
  assign n3489 = n9940 & ~n3422;
  assign n3490 = ~n3488 & ~n3489;
  assign n3491 = n9940 & n9945;
  assign n3492 = ~n3420 & ~n3491;
  assign n3493 = ~n3421 & n3492;
  assign n3494 = n3422 & ~n3491;
  assign n3495 = ~n9940 & ~n9945;
  assign n3496 = ~n9954 & ~n3495;
  assign n3497 = ~n9946 & ~n3489;
  assign n3498 = ~n3488 & ~n9955;
  assign n3499 = ~n9946 & n3490;
  assign n3500 = n3486 & ~n3487;
  assign n3501 = ~n3437 & ~n3484;
  assign n3502 = ~n2893 & n9914;
  assign n3503 = ~n3186 & ~n3502;
  assign n3504 = ~n3458 & ~n3476;
  assign n3505 = n9904 & ~n9905;
  assign n3506 = ~n3124 & ~n3505;
  assign n3507 = ~n3504 & n3506;
  assign n3508 = n3504 & ~n3506;
  assign n3509 = ~n3504 & ~n3507;
  assign n3510 = n3506 & ~n3507;
  assign n3511 = ~n3509 & ~n3510;
  assign n3512 = ~n3507 & ~n3508;
  assign n3513 = n3503 & ~n9957;
  assign n3514 = ~n3503 & n9957;
  assign n3515 = ~n3513 & ~n3514;
  assign n3516 = ~n3501 & n3515;
  assign n3517 = ~n3500 & ~n3516;
  assign n3518 = ~n9956 & n3517;
  assign n3519 = n3501 & ~n3515;
  assign n3520 = ~n3487 & ~n9955;
  assign n3521 = n3487 & n9955;
  assign n3522 = n3486 & ~n3521;
  assign n3523 = ~n3520 & ~n3522;
  assign n3524 = n3486 & ~n9955;
  assign n3525 = n3487 & ~n3524;
  assign n3526 = ~n3486 & n9955;
  assign n3527 = ~n3525 & ~n3526;
  assign n3528 = ~n9956 & ~n3500;
  assign n3529 = n3515 & ~n9958;
  assign n3530 = n3501 & ~n3529;
  assign n3531 = ~n3515 & n9958;
  assign n3532 = ~n3530 & ~n3531;
  assign n3533 = ~n3501 & ~n9958;
  assign n3534 = n3501 & n9958;
  assign n3535 = n3515 & ~n3534;
  assign n3536 = ~n3533 & ~n3535;
  assign n3537 = ~n3518 & ~n3519;
  assign n3538 = n3197 & n9959;
  assign n3539 = ~n3507 & ~n3513;
  assign n3540 = ~n3538 & n3539;
  assign n3541 = ~n3197 & ~n9959;
  assign n3542 = ~n9959 & n3539;
  assign n3543 = ~n3195 & ~n3542;
  assign n3544 = ~n3196 & n3543;
  assign n3545 = n3197 & ~n3542;
  assign n3546 = n9959 & ~n3539;
  assign n3547 = ~n9960 & ~n3546;
  assign n3548 = ~n3540 & ~n3541;
  assign n3549 = n3148 & ~n9961;
  assign n3550 = ~n3190 & ~n3195;
  assign n3551 = ~n3549 & n3550;
  assign n3552 = ~n3148 & n9961;
  assign n3553 = ~n9961 & ~n3550;
  assign n3554 = n9961 & n3550;
  assign n3555 = n3148 & ~n3554;
  assign n3556 = ~n3553 & ~n3555;
  assign n3557 = ~n3551 & ~n3552;
  assign n3558 = n3071 & ~n9962;
  assign n3559 = ~n3140 & ~n3146;
  assign n3560 = ~n3558 & n3559;
  assign n3561 = ~n3071 & n9962;
  assign n3562 = n9962 & n3559;
  assign n3563 = ~n3070 & ~n3562;
  assign n3564 = ~n3063 & n3563;
  assign n3565 = n3071 & ~n3562;
  assign n3566 = ~n9962 & ~n3559;
  assign n3567 = ~n9963 & ~n3566;
  assign n3568 = ~n3560 & ~n3561;
  assign n3569 = n3069 & ~n9964;
  assign n3570 = ~n3067 & ~n3569;
  assign n3571 = n2985 & ~n2987;
  assign n3572 = ~n2988 & ~n3571;
  assign n3573 = ~n3570 & n3572;
  assign n3574 = ~n2988 & ~n3573;
  assign n3575 = n2867 & ~n2869;
  assign n3576 = ~n2870 & ~n3575;
  assign n3577 = ~n3574 & n3576;
  assign n3578 = ~n2870 & ~n3577;
  assign n3579 = n2809 & ~n2811;
  assign n3580 = ~n2812 & ~n3579;
  assign n3581 = ~n3578 & n3580;
  assign n3582 = ~n2812 & ~n3581;
  assign n3583 = n2704 & n9849;
  assign n3584 = ~n2704 & n9849;
  assign n3585 = n2704 & ~n9849;
  assign n3586 = ~n3584 & ~n3585;
  assign n3587 = ~n2712 & ~n3583;
  assign n3588 = ~n3582 & ~n9965;
  assign n3589 = ~n2712 & ~n3588;
  assign n3590 = n2469 & n2472;
  assign n3591 = ~n2473 & ~n3590;
  assign n3592 = ~n3589 & n3591;
  assign n3593 = ~n2473 & ~n3592;
  assign n3594 = n9782 & n9797;
  assign n3595 = ~n9782 & ~n2289;
  assign n3596 = ~n9797 & ~n2289;
  assign n3597 = ~n3595 & ~n3596;
  assign n3598 = ~n2289 & ~n3594;
  assign n3599 = ~n3593 & ~n9966;
  assign n3600 = ~n2289 & ~n3599;
  assign n3601 = n2205 & ~n2207;
  assign n3602 = ~n2208 & ~n3601;
  assign n3603 = ~n3600 & n3602;
  assign n3604 = ~n2208 & ~n3603;
  assign n3605 = n1777 & n9737;
  assign n3606 = ~n1777 & n9737;
  assign n3607 = n1777 & ~n9737;
  assign n3608 = ~n3606 & ~n3607;
  assign n3609 = ~n1785 & ~n3605;
  assign n3610 = ~n3604 & ~n9967;
  assign n3611 = ~n1785 & ~n3610;
  assign n3612 = n1379 & ~n1401;
  assign n3613 = ~n1402 & ~n3612;
  assign n3614 = ~n3611 & n3613;
  assign n3615 = ~n1402 & ~n3614;
  assign n3616 = ~n1392 & ~n1399;
  assign n3617 = ~n1347 & ~n1396;
  assign n3618 = n9624 & n1164;
  assign n3619 = n9649 & ~n1164;
  assign n3620 = n9624 & ~n3619;
  assign n3621 = n9649 & ~n3618;
  assign n3622 = n1137 & ~n1164;
  assign n3623 = ~n9968 & ~n3622;
  assign n3624 = ~n1359 & n3623;
  assign n3625 = n1359 & ~n3623;
  assign n3626 = ~n3624 & ~n3625;
  assign n3627 = ~n3617 & ~n3624;
  assign n3628 = ~n3625 & n3627;
  assign n3629 = ~n3617 & n3626;
  assign n3630 = n3617 & ~n3626;
  assign n3631 = ~n3617 & ~n9969;
  assign n3632 = ~n3624 & ~n9969;
  assign n3633 = ~n3625 & n3632;
  assign n3634 = ~n3631 & ~n3633;
  assign n3635 = ~n9969 & ~n3630;
  assign n3636 = ~n3616 & ~n9970;
  assign n3637 = n3616 & n9970;
  assign n3638 = ~n3616 & n9970;
  assign n3639 = n3616 & ~n9970;
  assign n3640 = ~n3638 & ~n3639;
  assign n3641 = ~n3636 & ~n3637;
  assign n3642 = ~n3615 & ~n9971;
  assign n3643 = n3615 & n9971;
  assign n3644 = ~n3642 & ~n3643;
  assign n3645 = ~n676 & ~n772;
  assign n3646 = ~n404 & ~n757;
  assign n3647 = ~n294 & ~n381;
  assign n3648 = n3646 & n3647;
  assign n3649 = ~n381 & ~n757;
  assign n3650 = ~n294 & ~n404;
  assign n3651 = n3645 & n3650;
  assign n3652 = n3649 & n3651;
  assign n3653 = ~n381 & ~n404;
  assign n3654 = ~n294 & ~n757;
  assign n3655 = n3645 & n3654;
  assign n3656 = n3653 & n3655;
  assign n3657 = n3645 & n3648;
  assign n3658 = ~n404 & n9599;
  assign n3659 = ~n772 & n3658;
  assign n3660 = ~n757 & n3659;
  assign n3661 = ~n676 & n3660;
  assign n3662 = ~n381 & n3661;
  assign n3663 = ~n294 & n3662;
  assign n3664 = n9599 & n9972;
  assign n3665 = n389 & n899;
  assign n3666 = n481 & n777;
  assign n3667 = n389 & n481;
  assign n3668 = n777 & n899;
  assign n3669 = n3667 & n3668;
  assign n3670 = n3665 & n3666;
  assign n3671 = ~n401 & ~n627;
  assign n3672 = ~n401 & ~n1070;
  assign n3673 = ~n627 & n3672;
  assign n3674 = ~n1070 & n3671;
  assign n3675 = ~n9559 & ~n714;
  assign n3676 = ~n432 & ~n538;
  assign n3677 = ~n432 & ~n714;
  assign n3678 = ~n9559 & ~n538;
  assign n3679 = n3677 & n3678;
  assign n3680 = n3675 & n3676;
  assign n3681 = n9975 & n9976;
  assign n3682 = n777 & n3676;
  assign n3683 = n3665 & n3682;
  assign n3684 = n481 & n3675;
  assign n3685 = n9975 & n3684;
  assign n3686 = n3683 & n3685;
  assign n3687 = n9974 & n3681;
  assign n3688 = n9587 & n9977;
  assign n3689 = n9973 & n3688;
  assign n3690 = n551 & n9688;
  assign n3691 = ~n397 & ~n1083;
  assign n3692 = ~n1083 & n1479;
  assign n3693 = ~n397 & n3692;
  assign n3694 = n1479 & n3691;
  assign n3695 = n1818 & n9978;
  assign n3696 = n3690 & n3695;
  assign n3697 = ~n190 & ~n533;
  assign n3698 = ~n533 & ~n626;
  assign n3699 = ~n190 & n3698;
  assign n3700 = ~n626 & n3697;
  assign n3701 = ~n626 & n1206;
  assign n3702 = ~n533 & n3701;
  assign n3703 = ~n190 & n3702;
  assign n3704 = n1206 & n9979;
  assign n3705 = n353 & ~n384;
  assign n3706 = ~n384 & n477;
  assign n3707 = n353 & n3706;
  assign n3708 = n477 & n3705;
  assign n3709 = n9980 & n9981;
  assign n3710 = n353 & n9978;
  assign n3711 = n551 & n3710;
  assign n3712 = n1818 & n3711;
  assign n3713 = n9980 & n3712;
  assign n3714 = n9688 & n3713;
  assign n3715 = n477 & n3714;
  assign n3716 = ~n384 & n3715;
  assign n3717 = n3696 & n3709;
  assign n3718 = ~n164 & ~n674;
  assign n3719 = ~n770 & ~n1037;
  assign n3720 = ~n573 & n3719;
  assign n3721 = ~n164 & ~n573;
  assign n3722 = ~n770 & n3721;
  assign n3723 = ~n674 & n3722;
  assign n3724 = ~n1037 & n3723;
  assign n3725 = ~n573 & ~n674;
  assign n3726 = ~n164 & ~n1037;
  assign n3727 = ~n164 & ~n770;
  assign n3728 = ~n1037 & n3727;
  assign n3729 = ~n770 & n3726;
  assign n3730 = n3725 & n9984;
  assign n3731 = n3718 & n3720;
  assign n3732 = ~n202 & ~n534;
  assign n3733 = ~n9696 & n3732;
  assign n3734 = ~n175 & ~n249;
  assign n3735 = n553 & n3734;
  assign n3736 = n486 & n3735;
  assign n3737 = ~n202 & ~n249;
  assign n3738 = ~n9696 & n3737;
  assign n3739 = ~n534 & ~n552;
  assign n3740 = ~n175 & ~n219;
  assign n3741 = n3739 & n3740;
  assign n3742 = n486 & n3741;
  assign n3743 = n3738 & n3742;
  assign n3744 = ~n552 & n3737;
  assign n3745 = ~n219 & ~n9696;
  assign n3746 = ~n175 & ~n534;
  assign n3747 = n3745 & n3746;
  assign n3748 = n486 & n3747;
  assign n3749 = n3744 & n3748;
  assign n3750 = n3733 & n3736;
  assign n3751 = n486 & n9983;
  assign n3752 = ~n249 & n3751;
  assign n3753 = ~n175 & n3752;
  assign n3754 = ~n219 & n3753;
  assign n3755 = ~n534 & n3754;
  assign n3756 = ~n9696 & n3755;
  assign n3757 = ~n202 & n3756;
  assign n3758 = ~n552 & n3757;
  assign n3759 = n9983 & n9985;
  assign n3760 = n9982 & n9986;
  assign n3761 = n389 & n777;
  assign n3762 = n899 & n3761;
  assign n3763 = n9587 & n3762;
  assign n3764 = n9973 & n3763;
  assign n3765 = n9982 & n3764;
  assign n3766 = n9986 & n3765;
  assign n3767 = n9975 & n3766;
  assign n3768 = ~n714 & n3767;
  assign n3769 = ~n432 & n3768;
  assign n3770 = ~n324 & n3769;
  assign n3771 = ~n538 & n3770;
  assign n3772 = ~n9559 & n3771;
  assign n3773 = ~n480 & n3772;
  assign n3774 = n3689 & n3760;
  assign n3775 = ~n3644 & ~n9987;
  assign n3776 = n3611 & ~n3613;
  assign n3777 = ~n3614 & ~n3776;
  assign n3778 = n659 & n1247;
  assign n3779 = ~n300 & ~n533;
  assign n3780 = n411 & n3779;
  assign n3781 = n3778 & n3780;
  assign n3782 = ~n331 & ~n770;
  assign n3783 = ~n757 & n3782;
  assign n3784 = n9705 & n3783;
  assign n3785 = n9579 & n9597;
  assign n3786 = n3784 & n3785;
  assign n3787 = ~n331 & ~n533;
  assign n3788 = n659 & n3787;
  assign n3789 = n411 & n1247;
  assign n3790 = n3788 & n3789;
  assign n3791 = ~n300 & ~n757;
  assign n3792 = ~n770 & n3791;
  assign n3793 = n9579 & n3792;
  assign n3794 = n9597 & n9705;
  assign n3795 = n3793 & n3794;
  assign n3796 = n3790 & n3795;
  assign n3797 = ~n300 & ~n331;
  assign n3798 = n411 & n3797;
  assign n3799 = n3778 & n3798;
  assign n3800 = ~n533 & ~n770;
  assign n3801 = ~n757 & n3800;
  assign n3802 = n9705 & n3801;
  assign n3803 = n3785 & n3802;
  assign n3804 = n3799 & n3803;
  assign n3805 = n3781 & n3786;
  assign n3806 = n9655 & n9703;
  assign n3807 = n9988 & n3806;
  assign n3808 = n411 & n9597;
  assign n3809 = n9705 & n3808;
  assign n3810 = n659 & n3809;
  assign n3811 = n1247 & n3810;
  assign n3812 = n9579 & n3811;
  assign n3813 = n9703 & n3812;
  assign n3814 = n9655 & n3813;
  assign n3815 = n9745 & n3814;
  assign n3816 = ~n757 & n3815;
  assign n3817 = ~n533 & n3816;
  assign n3818 = ~n770 & n3817;
  assign n3819 = ~n331 & n3818;
  assign n3820 = ~n300 & n3819;
  assign n3821 = n9745 & n3807;
  assign n3822 = ~n3777 & ~n9989;
  assign n3823 = n3604 & n9967;
  assign n3824 = ~n3610 & ~n3823;
  assign n3825 = ~n164 & ~n714;
  assign n3826 = ~n714 & ~n871;
  assign n3827 = ~n164 & n3826;
  assign n3828 = ~n871 & n3825;
  assign n3829 = ~n9551 & ~n9561;
  assign n3830 = ~n311 & ~n534;
  assign n3831 = ~n9551 & ~n534;
  assign n3832 = ~n311 & ~n9561;
  assign n3833 = n3831 & n3832;
  assign n3834 = ~n9561 & ~n534;
  assign n3835 = ~n9551 & ~n311;
  assign n3836 = n3834 & n3835;
  assign n3837 = n3829 & n3830;
  assign n3838 = n9990 & n9991;
  assign n3839 = n9975 & n9978;
  assign n3840 = n9978 & n9991;
  assign n3841 = n9975 & n9990;
  assign n3842 = n3840 & n3841;
  assign n3843 = n3838 & n3839;
  assign n3844 = ~n301 & ~n511;
  assign n3845 = n753 & n1247;
  assign n3846 = n753 & n3844;
  assign n3847 = n1247 & n3846;
  assign n3848 = n3844 & n3845;
  assign n3849 = n9546 & n9993;
  assign n3850 = n9978 & n9990;
  assign n3851 = n3844 & n3850;
  assign n3852 = n753 & n3851;
  assign n3853 = n1247 & n3852;
  assign n3854 = n9975 & n3853;
  assign n3855 = n9546 & n3854;
  assign n3856 = ~n9561 & n3855;
  assign n3857 = ~n311 & n3856;
  assign n3858 = ~n9551 & n3857;
  assign n3859 = ~n534 & n3858;
  assign n3860 = n9992 & n3849;
  assign n3861 = ~n351 & ~n381;
  assign n3862 = ~n9586 & n3861;
  assign n3863 = ~n573 & ~n720;
  assign n3864 = n1558 & n3863;
  assign n3865 = ~n573 & n1558;
  assign n3866 = ~n9586 & n3865;
  assign n3867 = ~n381 & n3866;
  assign n3868 = ~n720 & n3867;
  assign n3869 = ~n351 & n3868;
  assign n3870 = ~n381 & ~n573;
  assign n3871 = ~n720 & n3870;
  assign n3872 = ~n351 & ~n9586;
  assign n3873 = n1558 & n3872;
  assign n3874 = n3871 & n3873;
  assign n3875 = ~n351 & ~n573;
  assign n3876 = ~n9586 & n3875;
  assign n3877 = ~n381 & ~n720;
  assign n3878 = n1558 & n3877;
  assign n3879 = n3876 & n3878;
  assign n3880 = n3862 & n3864;
  assign n3881 = ~n9555 & ~n554;
  assign n3882 = ~n9550 & ~n552;
  assign n3883 = n3881 & n3882;
  assign n3884 = n9658 & n3883;
  assign n3885 = n9547 & n3884;
  assign n3886 = n9547 & n9658;
  assign n3887 = n9995 & n3886;
  assign n3888 = ~n9555 & n3887;
  assign n3889 = ~n9550 & n3888;
  assign n3890 = ~n554 & n3889;
  assign n3891 = ~n552 & n3890;
  assign n3892 = n9995 & n3885;
  assign n3893 = ~n470 & ~n604;
  assign n3894 = ~n582 & ~n604;
  assign n3895 = ~n470 & n3894;
  assign n3896 = ~n582 & n3893;
  assign n3897 = ~n325 & ~n513;
  assign n3898 = ~n9553 & ~n513;
  assign n3899 = ~n325 & n3898;
  assign n3900 = ~n9553 & ~n325;
  assign n3901 = ~n513 & n3900;
  assign n3902 = ~n9553 & n3897;
  assign n3903 = ~n352 & n1852;
  assign n3904 = n9998 & n3903;
  assign n3905 = n9997 & n3903;
  assign n3906 = n9998 & n3905;
  assign n3907 = n9997 & n3904;
  assign n3908 = n385 & n1038;
  assign n3909 = n1259 & n3908;
  assign n3910 = n9543 & n3909;
  assign n3911 = ~n352 & n385;
  assign n3912 = n9998 & n3911;
  assign n3913 = n9997 & n3912;
  assign n3914 = n1038 & n1259;
  assign n3915 = n1852 & n3914;
  assign n3916 = n9543 & n3915;
  assign n3917 = n3913 & n3916;
  assign n3918 = n9999 & n3910;
  assign n3919 = n9996 & n10000;
  assign n3920 = n1038 & n9997;
  assign n3921 = n9998 & n3920;
  assign n3922 = n385 & n3921;
  assign n3923 = n9543 & n3922;
  assign n3924 = n1259 & n3923;
  assign n3925 = n9996 & n3924;
  assign n3926 = n9994 & n3925;
  assign n3927 = ~n663 & n3926;
  assign n3928 = ~n776 & n3927;
  assign n3929 = ~n352 & n3928;
  assign n3930 = n9994 & n10000;
  assign n3931 = n9996 & n3930;
  assign n3932 = n9994 & n3919;
  assign n3933 = ~n3824 & ~n10001;
  assign n3934 = n3600 & ~n3602;
  assign n3935 = ~n3603 & ~n3934;
  assign n3936 = ~n284 & ~n480;
  assign n3937 = ~n9564 & ~n480;
  assign n3938 = ~n284 & n3937;
  assign n3939 = ~n9564 & n3936;
  assign n3940 = ~n9564 & n9994;
  assign n3941 = ~n284 & n3940;
  assign n3942 = ~n480 & n3941;
  assign n3943 = n9994 & n10002;
  assign n3944 = n686 & n3897;
  assign n3945 = ~n405 & ~n431;
  assign n3946 = ~n1108 & ~n1190;
  assign n3947 = n3945 & n3946;
  assign n3948 = n3944 & n3947;
  assign n3949 = ~n302 & n908;
  assign n3950 = n1010 & n3949;
  assign n3951 = n908 & n9998;
  assign n3952 = n1010 & n3951;
  assign n3953 = ~n405 & n3952;
  assign n3954 = ~n468 & n3953;
  assign n3955 = ~n296 & n3954;
  assign n3956 = ~n431 & n3955;
  assign n3957 = ~n1108 & n3956;
  assign n3958 = ~n9559 & n3957;
  assign n3959 = ~n1190 & n3958;
  assign n3960 = n686 & n3945;
  assign n3961 = n686 & n908;
  assign n3962 = n3945 & n3961;
  assign n3963 = n908 & n3960;
  assign n3964 = ~n9559 & ~n1190;
  assign n3965 = ~n9559 & ~n1108;
  assign n3966 = ~n1190 & n3965;
  assign n3967 = ~n1108 & n3964;
  assign n3968 = n1010 & n10006;
  assign n3969 = n9998 & n3968;
  assign n3970 = n10005 & n3969;
  assign n3971 = ~n405 & ~n1108;
  assign n3972 = n686 & n3971;
  assign n3973 = n908 & n3972;
  assign n3974 = ~n9559 & ~n431;
  assign n3975 = ~n1190 & n3974;
  assign n3976 = n1010 & n3975;
  assign n3977 = n9998 & n3976;
  assign n3978 = n3973 & n3977;
  assign n3979 = n3948 & n3950;
  assign n3980 = ~n9537 & ~n604;
  assign n3981 = ~n9541 & n3980;
  assign n3982 = ~n168 & ~n604;
  assign n3983 = ~n219 & ~n334;
  assign n3984 = ~n168 & ~n219;
  assign n3985 = ~n334 & ~n604;
  assign n3986 = n3984 & n3985;
  assign n3987 = n10007 & n3983;
  assign n3988 = n1432 & n1665;
  assign n3989 = n10008 & n3988;
  assign n3990 = ~n205 & ~n300;
  assign n3991 = ~n205 & ~n9586;
  assign n3992 = ~n300 & n3991;
  assign n3993 = ~n300 & ~n9586;
  assign n3994 = ~n205 & n3993;
  assign n3995 = ~n9586 & n3990;
  assign n3996 = n9828 & n10009;
  assign n3997 = n1665 & n3983;
  assign n3998 = n1432 & n3997;
  assign n3999 = n9828 & n10007;
  assign n4000 = n10009 & n3999;
  assign n4001 = n3998 & n4000;
  assign n4002 = n3989 & n3996;
  assign n4003 = n9973 & n10010;
  assign n4004 = n10004 & n4003;
  assign n4005 = n9828 & n10003;
  assign n4006 = n10009 & n4005;
  assign n4007 = n1665 & n4006;
  assign n4008 = n9973 & n4007;
  assign n4009 = n10004 & n4008;
  assign n4010 = n1432 & n4009;
  assign n4011 = ~n334 & n4010;
  assign n4012 = ~n9537 & n4011;
  assign n4013 = ~n219 & n4012;
  assign n4014 = ~n9541 & n4013;
  assign n4015 = ~n604 & n4014;
  assign n4016 = n10003 & n4004;
  assign n4017 = ~n3935 & ~n10011;
  assign n4018 = n3593 & n9966;
  assign n4019 = ~n3599 & ~n4018;
  assign n4020 = ~n536 & ~n674;
  assign n4021 = ~n536 & n9715;
  assign n4022 = ~n674 & n4021;
  assign n4023 = n9715 & n4020;
  assign n4024 = ~n312 & ~n618;
  assign n4025 = ~n192 & ~n757;
  assign n4026 = n4024 & n4025;
  assign n4027 = n406 & n1259;
  assign n4028 = ~n225 & ~n9586;
  assign n4029 = n1838 & n4028;
  assign n4030 = n4027 & n4029;
  assign n4031 = n406 & n4025;
  assign n4032 = n1259 & n1838;
  assign n4033 = n4024 & n4028;
  assign n4034 = n4032 & n4033;
  assign n4035 = n4031 & n4034;
  assign n4036 = ~n192 & ~n225;
  assign n4037 = ~n9586 & ~n757;
  assign n4038 = n4036 & n4037;
  assign n4039 = n406 & n4024;
  assign n4040 = n4032 & n4039;
  assign n4041 = n4038 & n4040;
  assign n4042 = n4026 & n4030;
  assign n4043 = n406 & n1838;
  assign n4044 = n9722 & n4043;
  assign n4045 = n1259 & n4044;
  assign n4046 = n4024 & n4045;
  assign n4047 = ~n225 & n4046;
  assign n4048 = ~n757 & n4047;
  assign n4049 = ~n9586 & n4048;
  assign n4050 = ~n192 & n4049;
  assign n4051 = n9722 & n10013;
  assign n4052 = ~n380 & ~n479;
  assign n4053 = ~n241 & ~n432;
  assign n4054 = ~n260 & n4053;
  assign n4055 = ~n380 & n4053;
  assign n4056 = ~n479 & n4055;
  assign n4057 = ~n260 & n4056;
  assign n4058 = ~n241 & ~n479;
  assign n4059 = ~n380 & ~n432;
  assign n4060 = ~n260 & n4059;
  assign n4061 = n4058 & n4060;
  assign n4062 = ~n260 & n4052;
  assign n4063 = n4053 & n4062;
  assign n4064 = n4052 & n4054;
  assign n4065 = ~n331 & ~n676;
  assign n4066 = ~n301 & ~n414;
  assign n4067 = ~n301 & ~n676;
  assign n4068 = ~n331 & ~n414;
  assign n4069 = n4067 & n4068;
  assign n4070 = n4065 & n4066;
  assign n4071 = n2548 & n3881;
  assign n4072 = ~n9555 & ~n414;
  assign n4073 = ~n554 & n4072;
  assign n4074 = ~n335 & n4073;
  assign n4075 = ~n301 & n4074;
  assign n4076 = ~n676 & n4075;
  assign n4077 = ~n243 & n4076;
  assign n4078 = ~n331 & n4077;
  assign n4079 = ~n243 & ~n414;
  assign n4080 = n4067 & n4079;
  assign n4081 = ~n331 & ~n335;
  assign n4082 = n3881 & n4081;
  assign n4083 = n4080 & n4082;
  assign n4084 = n10016 & n4071;
  assign n4085 = ~n592 & ~n627;
  assign n4086 = ~n470 & ~n682;
  assign n4087 = n4085 & n4086;
  assign n4088 = ~n195 & ~n714;
  assign n4089 = n1009 & n4088;
  assign n4090 = ~n470 & ~n592;
  assign n4091 = ~n682 & ~n714;
  assign n4092 = n4090 & n4091;
  assign n4093 = ~n195 & ~n627;
  assign n4094 = n1009 & n4093;
  assign n4095 = n4092 & n4094;
  assign n4096 = n4088 & n4090;
  assign n4097 = ~n627 & ~n682;
  assign n4098 = n1009 & n4097;
  assign n4099 = n4096 & n4098;
  assign n4100 = n4087 & n4089;
  assign n4101 = n10017 & n10018;
  assign n4102 = n10015 & n4101;
  assign n4103 = n10014 & n4102;
  assign n4104 = n10012 & n10015;
  assign n4105 = n10014 & n4104;
  assign n4106 = n10017 & n4105;
  assign n4107 = ~n714 & n4106;
  assign n4108 = ~n592 & n4107;
  assign n4109 = ~n682 & n4108;
  assign n4110 = ~n627 & n4109;
  assign n4111 = ~n195 & n4110;
  assign n4112 = n1009 & n4111;
  assign n4113 = ~n470 & n4112;
  assign n4114 = n10012 & n4103;
  assign n4115 = ~n4019 & ~n10019;
  assign n4116 = n3589 & ~n3591;
  assign n4117 = ~n3592 & ~n4116;
  assign n4118 = ~n623 & ~n990;
  assign n4119 = ~n552 & ~n623;
  assign n4120 = ~n990 & n4119;
  assign n4121 = ~n552 & n4118;
  assign n4122 = ~n990 & n9640;
  assign n4123 = ~n552 & n4122;
  assign n4124 = ~n623 & n4123;
  assign n4125 = n9640 & n10020;
  assign n4126 = ~n380 & ~n414;
  assign n4127 = ~n241 & ~n515;
  assign n4128 = n1867 & n4127;
  assign n4129 = n4126 & n4128;
  assign n4130 = n9717 & n4129;
  assign n4131 = n10021 & n4130;
  assign n4132 = n1092 & n1570;
  assign n4133 = ~n260 & ~n674;
  assign n4134 = n1611 & n4133;
  assign n4135 = n1092 & n1611;
  assign n4136 = n1570 & n4133;
  assign n4137 = n4135 & n4136;
  assign n4138 = n1092 & n4133;
  assign n4139 = n1570 & n1611;
  assign n4140 = n4138 & n4139;
  assign n4141 = n4132 & n4134;
  assign n4142 = n9573 & n1570;
  assign n4143 = n1611 & n4142;
  assign n4144 = ~n332 & n4143;
  assign n4145 = ~n258 & n4144;
  assign n4146 = ~n674 & n4145;
  assign n4147 = ~n260 & n4146;
  assign n4148 = n9573 & n10022;
  assign n4149 = ~n295 & ~n536;
  assign n4150 = ~n351 & n4149;
  assign n4151 = ~n295 & n537;
  assign n4152 = ~n265 & ~n9564;
  assign n4153 = n1192 & n4152;
  assign n4154 = n683 & n909;
  assign n4155 = n4153 & n4154;
  assign n4156 = n10024 & n4155;
  assign n4157 = n10023 & n4156;
  assign n4158 = n1192 & n1867;
  assign n4159 = n4126 & n4158;
  assign n4160 = n9717 & n4159;
  assign n4161 = n10021 & n4160;
  assign n4162 = n4127 & n4152;
  assign n4163 = n4154 & n4162;
  assign n4164 = n10024 & n4163;
  assign n4165 = n10023 & n4164;
  assign n4166 = n4161 & n4165;
  assign n4167 = n909 & n1192;
  assign n4168 = n683 & n4126;
  assign n4169 = n4167 & n4168;
  assign n4170 = n9717 & n4169;
  assign n4171 = n10021 & n4170;
  assign n4172 = ~n241 & ~n9564;
  assign n4173 = ~n515 & n4172;
  assign n4174 = n9749 & n4173;
  assign n4175 = n10024 & n4174;
  assign n4176 = n10023 & n4175;
  assign n4177 = n4171 & n4176;
  assign n4178 = n4131 & n4157;
  assign n4179 = n683 & n10024;
  assign n4180 = n4126 & n4179;
  assign n4181 = n9749 & n4180;
  assign n4182 = n1192 & n4181;
  assign n4183 = n909 & n4182;
  assign n4184 = n10023 & n4183;
  assign n4185 = n9694 & n4184;
  assign n4186 = n9717 & n4185;
  assign n4187 = n10021 & n4186;
  assign n4188 = ~n9564 & n4187;
  assign n4189 = ~n241 & n4188;
  assign n4190 = ~n515 & n4189;
  assign n4191 = n9694 & n10025;
  assign n4192 = ~n4117 & ~n10026;
  assign n4193 = n3582 & n9965;
  assign n4194 = ~n3588 & ~n4193;
  assign n4195 = ~n9559 & ~n715;
  assign n4196 = ~n715 & n4024;
  assign n4197 = ~n9559 & n4196;
  assign n4198 = n4024 & n4195;
  assign n4199 = ~n730 & n1172;
  assign n4200 = ~n328 & ~n380;
  assign n4201 = ~n394 & n4200;
  assign n4202 = ~n380 & ~n394;
  assign n4203 = ~n328 & ~n730;
  assign n4204 = ~n380 & ~n730;
  assign n4205 = ~n328 & ~n394;
  assign n4206 = n4204 & n4205;
  assign n4207 = ~n394 & ~n730;
  assign n4208 = n4200 & n4207;
  assign n4209 = n4202 & n4203;
  assign n4210 = n1172 & n10028;
  assign n4211 = n4199 & n4201;
  assign n4212 = n10027 & n10029;
  assign n4213 = n9546 & n9764;
  assign n4214 = n1172 & n10027;
  assign n4215 = n9764 & n4214;
  assign n4216 = n9546 & n4215;
  assign n4217 = ~n328 & n4216;
  assign n4218 = ~n394 & n4217;
  assign n4219 = ~n380 & n4218;
  assign n4220 = ~n730 & n4219;
  assign n4221 = n4212 & n4213;
  assign n4222 = n385 & ~n9570;
  assign n4223 = n385 & n10030;
  assign n4224 = ~n9570 & n4223;
  assign n4225 = n10030 & n4222;
  assign n4226 = ~n179 & ~n871;
  assign n4227 = ~n179 & ~n352;
  assign n4228 = ~n871 & n4227;
  assign n4229 = ~n352 & n4226;
  assign n4230 = ~n468 & ~n897;
  assign n4231 = ~n217 & ~n264;
  assign n4232 = n4230 & n4231;
  assign n4233 = ~n300 & ~n682;
  assign n4234 = n662 & n4233;
  assign n4235 = ~n164 & ~n897;
  assign n4236 = ~n264 & ~n295;
  assign n4237 = n4235 & n4236;
  assign n4238 = ~n217 & ~n468;
  assign n4239 = n4233 & n4238;
  assign n4240 = n4237 & n4239;
  assign n4241 = n4232 & n4234;
  assign n4242 = n10032 & n10033;
  assign n4243 = n10032 & n4233;
  assign n4244 = n9711 & n4243;
  assign n4245 = ~n468 & n4244;
  assign n4246 = ~n897 & n4245;
  assign n4247 = ~n295 & n4246;
  assign n4248 = ~n164 & n4247;
  assign n4249 = ~n217 & n4248;
  assign n4250 = ~n264 & n4249;
  assign n4251 = n9711 & n4242;
  assign n4252 = ~n9550 & ~n511;
  assign n4253 = ~n294 & ~n1015;
  assign n4254 = n4252 & n4253;
  assign n4255 = n406 & n1532;
  assign n4256 = n406 & ~n933;
  assign n4257 = ~n9550 & n4256;
  assign n4258 = ~n604 & n4257;
  assign n4259 = ~n1015 & n4258;
  assign n4260 = ~n294 & n4259;
  assign n4261 = ~n511 & n4260;
  assign n4262 = ~n9550 & ~n294;
  assign n4263 = n1532 & n4262;
  assign n4264 = ~n511 & ~n1015;
  assign n4265 = n406 & n4264;
  assign n4266 = n4263 & n4265;
  assign n4267 = n4254 & n4255;
  assign n4268 = ~n219 & ~n9561;
  assign n4269 = n191 & n211;
  assign n4270 = ~n607 & ~n4269;
  assign n4271 = ~n192 & n4270;
  assign n4272 = n4268 & n4271;
  assign n4273 = ~n192 & ~n262;
  assign n4274 = ~n311 & n4273;
  assign n4275 = ~n476 & ~n607;
  assign n4276 = n477 & n4275;
  assign n4277 = n4268 & n4276;
  assign n4278 = n4274 & n4277;
  assign n4279 = ~n192 & ~n9561;
  assign n4280 = ~n311 & ~n476;
  assign n4281 = n4279 & n4280;
  assign n4282 = ~n219 & ~n262;
  assign n4283 = ~n607 & n4282;
  assign n4284 = n477 & n4283;
  assign n4285 = n4281 & n4284;
  assign n4286 = n478 & n4272;
  assign n4287 = n10035 & n10036;
  assign n4288 = n10034 & n4287;
  assign n4289 = ~n607 & n10031;
  assign n4290 = n10034 & n4289;
  assign n4291 = n477 & n4290;
  assign n4292 = n10035 & n4291;
  assign n4293 = ~n262 & n4292;
  assign n4294 = ~n9561 & n4293;
  assign n4295 = ~n311 & n4294;
  assign n4296 = ~n219 & n4295;
  assign n4297 = ~n192 & n4296;
  assign n4298 = ~n476 & n4297;
  assign n4299 = n10031 & n4288;
  assign n4300 = ~n4194 & ~n10037;
  assign n4301 = n3578 & ~n3580;
  assign n4302 = ~n3581 & ~n4301;
  assign n4303 = ~n258 & ~n674;
  assign n4304 = ~n9541 & ~n730;
  assign n4305 = ~n674 & ~n730;
  assign n4306 = ~n9541 & ~n258;
  assign n4307 = n4305 & n4306;
  assign n4308 = ~n258 & ~n730;
  assign n4309 = ~n9541 & ~n674;
  assign n4310 = n4308 & n4309;
  assign n4311 = n4303 & n4304;
  assign n4312 = n1558 & n10038;
  assign n4313 = n9556 & n9613;
  assign n4314 = n9997 & n4313;
  assign n4315 = n9556 & n9997;
  assign n4316 = n1558 & n4315;
  assign n4317 = n9613 & n4316;
  assign n4318 = ~n9541 & n4317;
  assign n4319 = ~n258 & n4318;
  assign n4320 = ~n674 & n4319;
  assign n4321 = ~n730 & n4320;
  assign n4322 = n4312 & n4314;
  assign n4323 = ~n301 & ~n627;
  assign n4324 = ~n352 & n4323;
  assign n4325 = ~n754 & ~n776;
  assign n4326 = ~n284 & ~n1037;
  assign n4327 = n4325 & n4326;
  assign n4328 = ~n301 & ~n352;
  assign n4329 = ~n1037 & n4328;
  assign n4330 = ~n627 & ~n754;
  assign n4331 = ~n284 & ~n776;
  assign n4332 = n4330 & n4331;
  assign n4333 = n4329 & n4332;
  assign n4334 = n4324 & n4327;
  assign n4335 = n9688 & n10040;
  assign n4336 = ~n195 & ~n9559;
  assign n4337 = n872 & n4336;
  assign n4338 = n1036 & n1868;
  assign n4339 = n872 & n1036;
  assign n4340 = ~n195 & n4339;
  assign n4341 = ~n265 & n4340;
  assign n4342 = ~n1015 & n4341;
  assign n4343 = ~n9559 & n4342;
  assign n4344 = n1868 & n4336;
  assign n4345 = n4339 & n4344;
  assign n4346 = n4337 & n4338;
  assign n4347 = ~n249 & ~n432;
  assign n4348 = n203 & n382;
  assign n4349 = n4347 & n4348;
  assign n4350 = n10041 & n4349;
  assign n4351 = ~n776 & ~n1037;
  assign n4352 = ~n352 & n4351;
  assign n4353 = ~n301 & ~n432;
  assign n4354 = ~n284 & ~n754;
  assign n4355 = n4353 & n4354;
  assign n4356 = n4352 & n4355;
  assign n4357 = n9688 & n4356;
  assign n4358 = ~n249 & ~n627;
  assign n4359 = n382 & n4358;
  assign n4360 = n203 & n4359;
  assign n4361 = n10041 & n4360;
  assign n4362 = n4357 & n4361;
  assign n4363 = n4335 & n4350;
  assign n4364 = n9580 & n10042;
  assign n4365 = n203 & n10041;
  assign n4366 = n10039 & n4365;
  assign n4367 = n9580 & n4366;
  assign n4368 = n9688 & n4367;
  assign n4369 = n382 & n4368;
  assign n4370 = ~n432 & n4369;
  assign n4371 = ~n627 & n4370;
  assign n4372 = ~n249 & n4371;
  assign n4373 = ~n776 & n4372;
  assign n4374 = ~n301 & n4373;
  assign n4375 = ~n754 & n4374;
  assign n4376 = ~n352 & n4375;
  assign n4377 = ~n1037 & n4376;
  assign n4378 = ~n284 & n4377;
  assign n4379 = n10039 & n4364;
  assign n4380 = ~n4302 & ~n10043;
  assign n4381 = n3574 & ~n3576;
  assign n4382 = ~n3577 & ~n4381;
  assign n4383 = n9687 & n4199;
  assign n4384 = n10009 & n4383;
  assign n4385 = ~n294 & ~n1190;
  assign n4386 = ~n1108 & n4385;
  assign n4387 = ~n294 & n3946;
  assign n4388 = ~n720 & ~n781;
  assign n4389 = ~n720 & n10044;
  assign n4390 = ~n781 & n4389;
  assign n4391 = ~n720 & ~n1108;
  assign n4392 = ~n1108 & n4388;
  assign n4393 = ~n781 & n4391;
  assign n4394 = n4385 & n10046;
  assign n4395 = n10044 & n4388;
  assign n4396 = ~n476 & n2091;
  assign n4397 = ~n179 & ~n284;
  assign n4398 = n1482 & n4397;
  assign n4399 = n4396 & n4398;
  assign n4400 = n10021 & n4399;
  assign n4401 = n10045 & n4400;
  assign n4402 = n10045 & n4398;
  assign n4403 = n10009 & n4402;
  assign n4404 = n1172 & n4403;
  assign n4405 = n10021 & n4404;
  assign n4406 = n9687 & n4405;
  assign n4407 = ~n431 & n4406;
  assign n4408 = ~n770 & n4407;
  assign n4409 = ~n476 & n4408;
  assign n4410 = ~n730 & n4409;
  assign n4411 = ~n476 & ~n730;
  assign n4412 = n1172 & n4411;
  assign n4413 = n9687 & n4412;
  assign n4414 = n10009 & n4413;
  assign n4415 = n1482 & n2091;
  assign n4416 = n4397 & n4415;
  assign n4417 = n10021 & n4416;
  assign n4418 = n10045 & n4417;
  assign n4419 = n4414 & n4418;
  assign n4420 = ~n730 & ~n770;
  assign n4421 = ~n431 & ~n476;
  assign n4422 = n2091 & n4411;
  assign n4423 = n4420 & n4421;
  assign n4424 = n9687 & n10048;
  assign n4425 = n10009 & n4424;
  assign n4426 = n1172 & n1482;
  assign n4427 = n4397 & n4426;
  assign n4428 = n10021 & n4427;
  assign n4429 = n10045 & n4428;
  assign n4430 = n4425 & n4429;
  assign n4431 = n4384 & n4401;
  assign n4432 = ~n250 & ~n538;
  assign n4433 = n773 & n908;
  assign n4434 = n4432 & n4433;
  assign n4435 = ~n9541 & ~n581;
  assign n4436 = ~n351 & n4435;
  assign n4437 = ~n467 & ~n714;
  assign n4438 = n1665 & n4437;
  assign n4439 = ~n9541 & n4437;
  assign n4440 = ~n351 & ~n581;
  assign n4441 = n1665 & n4440;
  assign n4442 = n4439 & n4441;
  assign n4443 = n4436 & n4438;
  assign n4444 = n908 & n1665;
  assign n4445 = n4432 & n4444;
  assign n4446 = ~n581 & ~n714;
  assign n4447 = ~n9541 & n4446;
  assign n4448 = ~n351 & ~n467;
  assign n4449 = n773 & n4448;
  assign n4450 = n4447 & n4449;
  assign n4451 = n4445 & n4450;
  assign n4452 = n4434 & n10049;
  assign n4453 = n9692 & n10041;
  assign n4454 = n10050 & n4453;
  assign n4455 = n9567 & n9708;
  assign n4456 = n9708 & n4454;
  assign n4457 = n9567 & n4456;
  assign n4458 = n4454 & n4455;
  assign n4459 = n10041 & n4434;
  assign n4460 = n1665 & n4459;
  assign n4461 = n9708 & n4460;
  assign n4462 = n9692 & n4461;
  assign n4463 = n10047 & n4462;
  assign n4464 = n9567 & n4463;
  assign n4465 = ~n714 & n4464;
  assign n4466 = ~n581 & n4465;
  assign n4467 = ~n467 & n4466;
  assign n4468 = ~n9541 & n4467;
  assign n4469 = ~n351 & n4468;
  assign n4470 = n10047 & n10051;
  assign n4471 = ~n4382 & ~n10052;
  assign n4472 = n3570 & ~n3572;
  assign n4473 = ~n3573 & ~n4472;
  assign n4474 = n659 & n1223;
  assign n4475 = n1223 & n4397;
  assign n4476 = n659 & n4475;
  assign n4477 = n4397 & n4474;
  assign n4478 = ~n9544 & ~n676;
  assign n4479 = ~n470 & ~n1015;
  assign n4480 = ~n470 & ~n676;
  assign n4481 = ~n9544 & ~n1015;
  assign n4482 = n4480 & n4481;
  assign n4483 = n4478 & n4479;
  assign n4484 = ~n9562 & ~n401;
  assign n4485 = ~n225 & ~n554;
  assign n4486 = n4484 & n4485;
  assign n4487 = ~n225 & ~n1015;
  assign n4488 = n4480 & n4487;
  assign n4489 = ~n401 & ~n554;
  assign n4490 = ~n9544 & ~n9562;
  assign n4491 = n4489 & n4490;
  assign n4492 = n4488 & n4491;
  assign n4493 = n10054 & n4486;
  assign n4494 = n9604 & n10055;
  assign n4495 = n4475 & n4484;
  assign n4496 = n659 & n4485;
  assign n4497 = n10054 & n4496;
  assign n4498 = n9604 & n4497;
  assign n4499 = n4495 & n4498;
  assign n4500 = n10053 & n4494;
  assign n4501 = ~n192 & ~n313;
  assign n4502 = ~n192 & ~n352;
  assign n4503 = ~n313 & n4502;
  assign n4504 = ~n352 & n4501;
  assign n4505 = ~n9564 & n1839;
  assign n4506 = ~n9555 & n4505;
  assign n4507 = ~n192 & n4506;
  assign n4508 = ~n352 & n4507;
  assign n4509 = n1839 & n10057;
  assign n4510 = ~n334 & ~n1083;
  assign n4511 = n142 & ~n949;
  assign n4512 = ~n398 & ~n4511;
  assign n4513 = ~n334 & ~n933;
  assign n4514 = ~n715 & n4513;
  assign n4515 = ~n1083 & n4514;
  assign n4516 = ~n398 & n4515;
  assign n4517 = ~n334 & ~n398;
  assign n4518 = ~n933 & ~n1083;
  assign n4519 = ~n715 & n4518;
  assign n4520 = ~n1083 & ~n4511;
  assign n4521 = n4517 & n10060;
  assign n4522 = n4510 & n4512;
  assign n4523 = n200 & n204;
  assign n4524 = ~n9537 & ~n4523;
  assign n4525 = ~n431 & ~n757;
  assign n4526 = ~n431 & ~n4523;
  assign n4527 = ~n9537 & ~n757;
  assign n4528 = n4526 & n4527;
  assign n4529 = ~n9537 & ~n384;
  assign n4530 = ~n205 & n4525;
  assign n4531 = n4529 & n4530;
  assign n4532 = n4524 & n4525;
  assign n4533 = n10059 & n10061;
  assign n4534 = n10058 & n10059;
  assign n4535 = ~n9537 & n4534;
  assign n4536 = ~n757 & n4535;
  assign n4537 = ~n431 & n4536;
  assign n4538 = ~n205 & n4537;
  assign n4539 = ~n384 & n4538;
  assign n4540 = n10058 & n10061;
  assign n4541 = n10059 & n4540;
  assign n4542 = n10058 & n4533;
  assign n4543 = n10023 & n10062;
  assign n4544 = n10023 & n10053;
  assign n4545 = n10062 & n4544;
  assign n4546 = n9604 & n4545;
  assign n4547 = ~n225 & n4546;
  assign n4548 = ~n9562 & n4547;
  assign n4549 = ~n401 & n4548;
  assign n4550 = ~n9544 & n4549;
  assign n4551 = ~n554 & n4550;
  assign n4552 = ~n1015 & n4551;
  assign n4553 = ~n676 & n4552;
  assign n4554 = ~n470 & n4553;
  assign n4555 = n10023 & n10056;
  assign n4556 = n10062 & n4555;
  assign n4557 = n10056 & n4543;
  assign n4558 = ~n4473 & ~n10063;
  assign n4559 = ~n3069 & n9964;
  assign n4560 = ~n9964 & ~n3569;
  assign n4561 = n3069 & ~n3569;
  assign n4562 = ~n4560 & ~n4561;
  assign n4563 = ~n3569 & ~n4559;
  assign n4564 = n9579 & n9581;
  assign n4565 = n9741 & n4564;
  assign n4566 = ~n9550 & ~n770;
  assign n4567 = ~n1190 & n4566;
  assign n4568 = ~n9544 & ~n9696;
  assign n4569 = n1172 & n4568;
  assign n4570 = n4567 & n4569;
  assign n4571 = n9709 & n4570;
  assign n4572 = n4565 & n4571;
  assign n4573 = n9982 & n4572;
  assign n4574 = n9581 & n9741;
  assign n4575 = n9709 & n4574;
  assign n4576 = n1172 & n4575;
  assign n4577 = n10039 & n4576;
  assign n4578 = n9579 & n4577;
  assign n4579 = n9982 & n4578;
  assign n4580 = ~n9550 & n4579;
  assign n4581 = ~n9544 & n4580;
  assign n4582 = ~n770 & n4581;
  assign n4583 = ~n9696 & n4582;
  assign n4584 = ~n1190 & n4583;
  assign n4585 = n10039 & n4573;
  assign n4586 = ~n10064 & n10065;
  assign n4587 = n4473 & n10063;
  assign n4588 = ~n4558 & ~n4587;
  assign n4589 = ~n4558 & ~n4586;
  assign n4590 = ~n4587 & n4589;
  assign n4591 = ~n4586 & n4588;
  assign n4592 = ~n4558 & ~n10066;
  assign n4593 = n4382 & n10052;
  assign n4594 = ~n4471 & ~n4593;
  assign n4595 = ~n4471 & ~n4592;
  assign n4596 = ~n4593 & n4595;
  assign n4597 = ~n4592 & n4594;
  assign n4598 = ~n4471 & ~n10067;
  assign n4599 = n4302 & n10043;
  assign n4600 = ~n4380 & ~n4599;
  assign n4601 = ~n4598 & n4600;
  assign n4602 = ~n4380 & ~n4601;
  assign n4603 = n4194 & n10037;
  assign n4604 = ~n4300 & ~n4603;
  assign n4605 = ~n4602 & n4604;
  assign n4606 = ~n4300 & ~n4605;
  assign n4607 = n4117 & n10026;
  assign n4608 = ~n4192 & ~n4607;
  assign n4609 = ~n4192 & ~n4606;
  assign n4610 = ~n4607 & n4609;
  assign n4611 = ~n4606 & n4608;
  assign n4612 = ~n4192 & ~n10068;
  assign n4613 = n4019 & n10019;
  assign n4614 = ~n10019 & ~n4115;
  assign n4615 = ~n4019 & ~n4115;
  assign n4616 = ~n4614 & ~n4615;
  assign n4617 = ~n4115 & ~n4613;
  assign n4618 = ~n4612 & ~n10069;
  assign n4619 = ~n4115 & ~n4618;
  assign n4620 = n3935 & n10011;
  assign n4621 = ~n4017 & ~n4620;
  assign n4622 = ~n4017 & ~n4619;
  assign n4623 = ~n4620 & n4622;
  assign n4624 = ~n4619 & n4621;
  assign n4625 = ~n4017 & ~n10070;
  assign n4626 = n3824 & n10001;
  assign n4627 = ~n3933 & ~n4626;
  assign n4628 = ~n4625 & n4627;
  assign n4629 = ~n3933 & ~n4628;
  assign n4630 = n3777 & n9989;
  assign n4631 = ~n3822 & ~n4630;
  assign n4632 = ~n3822 & ~n4629;
  assign n4633 = ~n4630 & n4632;
  assign n4634 = ~n4629 & n4631;
  assign n4635 = ~n3822 & ~n10071;
  assign n4636 = n3644 & n9987;
  assign n4637 = ~n3775 & ~n4636;
  assign n4638 = ~n4635 & n4637;
  assign n4639 = ~n3775 & ~n4638;
  assign n4640 = ~n386 & ~n623;
  assign n4641 = ~n467 & ~n754;
  assign n4642 = n4640 & n4641;
  assign n4643 = n1665 & n4484;
  assign n4644 = n994 & n1192;
  assign n4645 = n1192 & n4484;
  assign n4646 = n994 & n1665;
  assign n4647 = n4645 & n4646;
  assign n4648 = n4643 & n4644;
  assign n4649 = n4642 & n4643;
  assign n4650 = n4644 & n4649;
  assign n4651 = n4484 & n4641;
  assign n4652 = n1192 & n1665;
  assign n4653 = n994 & n4640;
  assign n4654 = n4652 & n4653;
  assign n4655 = n4651 & n4654;
  assign n4656 = n4642 & n10072;
  assign n4657 = ~n776 & ~n1108;
  assign n4658 = ~n468 & ~n776;
  assign n4659 = ~n1108 & n4658;
  assign n4660 = ~n468 & n4657;
  assign n4661 = ~n225 & ~n468;
  assign n4662 = ~n327 & n4661;
  assign n4663 = ~n776 & n4662;
  assign n4664 = ~n1108 & n4663;
  assign n4665 = ~n327 & ~n468;
  assign n4666 = ~n225 & n4657;
  assign n4667 = n4665 & n4666;
  assign n4668 = n1456 & n10074;
  assign n4669 = ~n331 & ~n897;
  assign n4670 = ~n674 & ~n897;
  assign n4671 = ~n331 & n4670;
  assign n4672 = ~n331 & ~n674;
  assign n4673 = ~n897 & n4672;
  assign n4674 = ~n674 & n4669;
  assign n4675 = ~n897 & n9990;
  assign n4676 = ~n331 & n4675;
  assign n4677 = ~n674 & n4676;
  assign n4678 = n9990 & n10076;
  assign n4679 = n10075 & n10077;
  assign n4680 = n10073 & n4679;
  assign n4681 = n9708 & n9752;
  assign n4682 = n4680 & n4681;
  assign n4683 = n994 & n10031;
  assign n4684 = n4640 & n4683;
  assign n4685 = n4641 & n4684;
  assign n4686 = n1192 & n4685;
  assign n4687 = n10075 & n4686;
  assign n4688 = n10077 & n4687;
  assign n4689 = n1665 & n4688;
  assign n4690 = n9708 & n4689;
  assign n4691 = n9752 & n4690;
  assign n4692 = ~n9562 & n4691;
  assign n4693 = ~n401 & n4692;
  assign n4694 = n10031 & n4682;
  assign n4695 = ~n1164 & n9670;
  assign n4696 = n1164 & ~n9670;
  assign n4697 = ~n1164 & ~n9670;
  assign n4698 = n1164 & n9670;
  assign n4699 = ~n4697 & ~n4698;
  assign n4700 = ~n4695 & ~n4696;
  assign n4701 = ~n1136 & ~n10079;
  assign n4702 = ~n1136 & n10079;
  assign n4703 = n1136 & ~n10079;
  assign n4704 = n1136 & n10079;
  assign n4705 = ~n4701 & ~n4704;
  assign n4706 = ~n4702 & ~n4703;
  assign n4707 = ~n9624 & n10080;
  assign n4708 = ~n9624 & ~n4701;
  assign n4709 = ~n3636 & ~n3642;
  assign n4710 = ~n3632 & n4709;
  assign n4711 = n3632 & ~n4709;
  assign n4712 = ~n4710 & ~n4711;
  assign n4713 = n10081 & n4712;
  assign n4714 = ~n10081 & ~n4712;
  assign n4715 = ~n4713 & ~n4714;
  assign n4716 = ~n10078 & ~n4715;
  assign n4717 = n10078 & n4715;
  assign n4718 = ~n4716 & ~n4717;
  assign n4719 = n4639 & ~n4718;
  assign n4720 = ~n4639 & ~n4716;
  assign n4721 = ~n4717 & n4720;
  assign n4722 = ~n4639 & n4718;
  assign n4723 = ~n4639 & ~n10082;
  assign n4724 = ~n4639 & ~n4717;
  assign n4725 = ~n4716 & ~n10082;
  assign n4726 = ~n4716 & ~n4724;
  assign n4727 = ~n4717 & n10083;
  assign n4728 = ~n4723 & ~n4727;
  assign n4729 = ~n4719 & ~n10082;
  assign n4730 = n4635 & ~n4637;
  assign n4731 = ~n4638 & ~n4730;
  assign n4732 = ~n10084 & n4731;
  assign n4733 = n4629 & ~n4631;
  assign n4734 = ~n4629 & ~n10071;
  assign n4735 = ~n4630 & n4635;
  assign n4736 = ~n4734 & ~n4735;
  assign n4737 = ~n10071 & ~n4733;
  assign n4738 = n4731 & ~n10085;
  assign n4739 = n4625 & ~n4627;
  assign n4740 = ~n4628 & ~n4739;
  assign n4741 = ~n10085 & n4740;
  assign n4742 = n4619 & ~n4621;
  assign n4743 = ~n4619 & ~n10070;
  assign n4744 = ~n4620 & n4625;
  assign n4745 = ~n4743 & ~n4744;
  assign n4746 = ~n10070 & ~n4742;
  assign n4747 = n4740 & ~n10086;
  assign n4748 = n4612 & n10069;
  assign n4749 = ~n4612 & ~n4618;
  assign n4750 = ~n10069 & ~n4618;
  assign n4751 = ~n4749 & ~n4750;
  assign n4752 = ~n4618 & ~n4748;
  assign n4753 = ~n10086 & ~n10087;
  assign n4754 = n4606 & ~n4608;
  assign n4755 = ~n4606 & ~n10068;
  assign n4756 = ~n4607 & n4612;
  assign n4757 = ~n4755 & ~n4756;
  assign n4758 = ~n10068 & ~n4754;
  assign n4759 = ~n10087 & ~n10088;
  assign n4760 = n4602 & ~n4604;
  assign n4761 = ~n4605 & ~n4760;
  assign n4762 = ~n10088 & n4761;
  assign n4763 = n4598 & ~n4600;
  assign n4764 = ~n4601 & ~n4763;
  assign n4765 = n4761 & n4764;
  assign n4766 = n4592 & ~n4594;
  assign n4767 = ~n4592 & ~n10067;
  assign n4768 = ~n4593 & n4598;
  assign n4769 = ~n4767 & ~n4768;
  assign n4770 = ~n10067 & ~n4766;
  assign n4771 = n4764 & ~n10089;
  assign n4772 = ~n4764 & n10089;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = n10064 & ~n10065;
  assign n4775 = ~n4586 & ~n4774;
  assign n4776 = n10089 & n4775;
  assign n4777 = n4586 & ~n4588;
  assign n4778 = ~n4586 & ~n10066;
  assign n4779 = ~n4587 & n4592;
  assign n4780 = ~n4778 & ~n4779;
  assign n4781 = ~n10066 & ~n4777;
  assign n4782 = ~n10089 & ~n10090;
  assign n4783 = ~n4775 & ~n10090;
  assign n4784 = n10089 & n4783;
  assign n4785 = ~n4782 & ~n4784;
  assign n4786 = ~n4776 & ~n10090;
  assign n4787 = ~n4772 & ~n10091;
  assign n4788 = ~n4771 & n4787;
  assign n4789 = n4773 & ~n10091;
  assign n4790 = ~n4771 & ~n10092;
  assign n4791 = ~n4761 & ~n4764;
  assign n4792 = ~n4765 & ~n4791;
  assign n4793 = ~n4790 & ~n4791;
  assign n4794 = ~n4765 & n4793;
  assign n4795 = ~n4790 & n4792;
  assign n4796 = ~n4765 & ~n10093;
  assign n4797 = n10088 & ~n4761;
  assign n4798 = ~n4762 & ~n4797;
  assign n4799 = ~n4796 & n4798;
  assign n4800 = ~n4762 & ~n4799;
  assign n4801 = n10087 & n10088;
  assign n4802 = ~n4759 & ~n4801;
  assign n4803 = ~n4800 & n4802;
  assign n4804 = ~n4759 & ~n4803;
  assign n4805 = n10086 & n10087;
  assign n4806 = ~n4753 & ~n4805;
  assign n4807 = ~n4804 & n4806;
  assign n4808 = ~n4753 & ~n4807;
  assign n4809 = ~n4740 & n10086;
  assign n4810 = ~n4747 & ~n4809;
  assign n4811 = ~n4808 & n4810;
  assign n4812 = ~n4747 & ~n4811;
  assign n4813 = n10085 & ~n4740;
  assign n4814 = ~n4741 & ~n4813;
  assign n4815 = ~n4812 & n4814;
  assign n4816 = ~n4741 & ~n4815;
  assign n4817 = ~n4731 & n10085;
  assign n4818 = ~n4738 & ~n4817;
  assign n4819 = ~n4816 & n4818;
  assign n4820 = ~n4738 & ~n4819;
  assign n4821 = n10084 & ~n4731;
  assign n4822 = ~n4732 & ~n4821;
  assign n4823 = ~n4820 & n4822;
  assign n4824 = ~n4732 & ~n4823;
  assign n4825 = ~n352 & ~n730;
  assign n4826 = n1630 & n2023;
  assign n4827 = n4825 & n4826;
  assign n4828 = n382 & n1038;
  assign n4829 = n1818 & n4828;
  assign n4830 = n1630 & n4828;
  assign n4831 = ~n730 & ~n772;
  assign n4832 = ~n205 & ~n352;
  assign n4833 = n4831 & n4832;
  assign n4834 = n1818 & n4833;
  assign n4835 = n4830 & n4834;
  assign n4836 = n4827 & n4829;
  assign n4837 = n9661 & n10094;
  assign n4838 = ~n328 & ~n468;
  assign n4839 = ~n9555 & ~n618;
  assign n4840 = ~n592 & n4839;
  assign n4841 = ~n468 & ~n618;
  assign n4842 = ~n9555 & ~n592;
  assign n4843 = ~n9555 & ~n328;
  assign n4844 = ~n592 & n4843;
  assign n4845 = ~n328 & n4842;
  assign n4846 = n4841 & n10095;
  assign n4847 = n4838 & n4840;
  assign n4848 = ~n592 & n9598;
  assign n4849 = ~n468 & n4848;
  assign n4850 = ~n9555 & n4849;
  assign n4851 = ~n328 & n4850;
  assign n4852 = ~n618 & n4851;
  assign n4853 = n9598 & n10096;
  assign n4854 = n10023 & n10097;
  assign n4855 = n4837 & n4854;
  assign n4856 = n1038 & n1818;
  assign n4857 = n10023 & n4856;
  assign n4858 = n9829 & n4857;
  assign n4859 = n10097 & n4858;
  assign n4860 = n9661 & n4859;
  assign n4861 = n382 & n4860;
  assign n4862 = ~n772 & n4861;
  assign n4863 = n1630 & n4862;
  assign n4864 = ~n205 & n4863;
  assign n4865 = ~n352 & n4864;
  assign n4866 = ~n730 & n4865;
  assign n4867 = n9829 & n4855;
  assign n4868 = n10083 & n10098;
  assign n4869 = ~n10083 & ~n10098;
  assign n4870 = ~n4868 & ~n4869;
  assign n4871 = ~n10084 & ~n4870;
  assign n4872 = n10084 & n4870;
  assign n4873 = ~n4871 & ~n4872;
  assign n4874 = ~n4824 & n4873;
  assign n4875 = n4824 & ~n4873;
  assign n4876 = ~n4874 & ~n4875;
  assign n4877 = n90 & n4876;
  assign n4878 = ~n9530 & n9531;
  assign n4879 = ~n4870 & n4878;
  assign n4880 = n9529 & ~n83;
  assign n4881 = ~n9529 & n83;
  assign n4882 = ~n9529 & ~n83;
  assign n4883 = n9529 & n83;
  assign n4884 = ~n4882 & ~n4883;
  assign n4885 = ~n4880 & ~n4881;
  assign n4886 = n9530 & ~n10099;
  assign n4887 = ~n10084 & n4886;
  assign n4888 = n9530 & ~n9531;
  assign n4889 = n9530 & n10099;
  assign n4890 = ~n9531 & n4889;
  assign n4891 = n10099 & n4888;
  assign n4892 = n4731 & n10100;
  assign n4893 = ~n4887 & ~n4892;
  assign n4894 = ~n4879 & ~n4892;
  assign n4895 = ~n4887 & n4894;
  assign n4896 = ~n4879 & n4893;
  assign n4897 = ~n4877 & n10101;
  assign n4898 = n9528 & ~n4897;
  assign n4899 = ~n9528 & n4897;
  assign n4900 = ~n4898 & ~n4899;
  assign n4901 = ~n978 & n9626;
  assign n4902 = n978 & ~n9626;
  assign n4903 = ~n978 & ~n9626;
  assign n4904 = n978 & n9626;
  assign n4905 = ~n4903 & ~n4904;
  assign n4906 = ~n4901 & ~n4902;
  assign n4907 = n9625 & ~n1703;
  assign n4908 = ~n9625 & n1703;
  assign n4909 = ~n9625 & ~n1703;
  assign n4910 = n9625 & n1703;
  assign n4911 = ~n4909 & ~n4910;
  assign n4912 = ~n4907 & ~n4908;
  assign n4913 = ~n10102 & ~n10103;
  assign n4914 = n4790 & ~n4792;
  assign n4915 = ~n4790 & ~n10093;
  assign n4916 = ~n4791 & n4796;
  assign n4917 = ~n4915 & ~n4916;
  assign n4918 = ~n10093 & ~n4914;
  assign n4919 = n4913 & ~n10104;
  assign n4920 = n10102 & ~n10103;
  assign n4921 = n4761 & n4920;
  assign n4922 = n9625 & ~n978;
  assign n4923 = ~n9625 & n978;
  assign n4924 = ~n9625 & ~n978;
  assign n4925 = n9625 & n978;
  assign n4926 = ~n4924 & ~n4925;
  assign n4927 = ~n4922 & ~n4923;
  assign n4928 = ~n10102 & n10103;
  assign n4929 = n10103 & n10105;
  assign n4930 = ~n10102 & n4929;
  assign n4931 = n10105 & n4928;
  assign n4932 = ~n10089 & n10106;
  assign n4933 = n10103 & ~n10105;
  assign n4934 = n4764 & n4933;
  assign n4935 = ~n4932 & ~n4934;
  assign n4936 = ~n4921 & ~n4934;
  assign n4937 = ~n4932 & n4936;
  assign n4938 = ~n4921 & n4935;
  assign n4939 = ~n4913 & n10107;
  assign n4940 = n10104 & n10107;
  assign n4941 = ~n4939 & ~n4940;
  assign n4942 = ~n4919 & n10107;
  assign n4943 = ~n9626 & ~n10108;
  assign n4944 = n9626 & n10108;
  assign n4945 = ~n4943 & ~n4944;
  assign n4946 = n9626 & ~n1149;
  assign n4947 = ~n9626 & n1149;
  assign n4948 = ~n9626 & ~n1149;
  assign n4949 = n9626 & n1149;
  assign n4950 = ~n4948 & ~n4949;
  assign n4951 = ~n4946 & ~n4947;
  assign n4952 = ~n1164 & ~n4775;
  assign n4953 = ~n10109 & n4952;
  assign n4954 = ~n4775 & n10090;
  assign n4955 = n4775 & ~n10090;
  assign n4956 = ~n4588 & n4775;
  assign n4957 = ~n4954 & ~n10110;
  assign n4958 = ~n10079 & ~n10109;
  assign n4959 = ~n4957 & n4958;
  assign n4960 = ~n1149 & n9670;
  assign n4961 = n1149 & ~n9670;
  assign n4962 = ~n1149 & ~n9670;
  assign n4963 = n1149 & n9670;
  assign n4964 = ~n4962 & ~n4963;
  assign n4965 = ~n4960 & ~n4961;
  assign n4966 = n10109 & ~n10111;
  assign n4967 = ~n4775 & n4966;
  assign n4968 = n10079 & ~n10109;
  assign n4969 = ~n10090 & n4968;
  assign n4970 = ~n4967 & ~n4969;
  assign n4971 = ~n4959 & n4970;
  assign n4972 = n4953 & ~n4971;
  assign n4973 = ~n4953 & n4971;
  assign n4974 = ~n4775 & ~n10109;
  assign n4975 = n4971 & ~n4974;
  assign n4976 = ~n1164 & ~n4974;
  assign n4977 = ~n1164 & ~n4971;
  assign n4978 = ~n1164 & ~n4977;
  assign n4979 = ~n4971 & ~n4977;
  assign n4980 = ~n4978 & ~n4979;
  assign n4981 = n4976 & ~n4980;
  assign n4982 = ~n1164 & n4975;
  assign n4983 = ~n4976 & n4980;
  assign n4984 = ~n10112 & ~n4983;
  assign n4985 = ~n4972 & ~n4973;
  assign n4986 = n4945 & n10113;
  assign n4987 = n4913 & ~n4957;
  assign n4988 = ~n4775 & n4933;
  assign n4989 = ~n10090 & n4920;
  assign n4990 = ~n4988 & ~n4989;
  assign n4991 = ~n4987 & n4990;
  assign n4992 = ~n4775 & ~n10103;
  assign n4993 = n9626 & ~n4992;
  assign n4994 = n9626 & ~n4991;
  assign n4995 = ~n9626 & n4991;
  assign n4996 = ~n4994 & ~n4995;
  assign n4997 = n4993 & n4996;
  assign n4998 = n4991 & n4993;
  assign n4999 = ~n10089 & ~n10110;
  assign n5000 = n10089 & n10110;
  assign n5001 = n10089 & ~n10110;
  assign n5002 = ~n10089 & n10110;
  assign n5003 = ~n5001 & ~n5002;
  assign n5004 = ~n4999 & ~n5000;
  assign n5005 = n4913 & n10115;
  assign n5006 = ~n10089 & n4920;
  assign n5007 = ~n4775 & n10106;
  assign n5008 = ~n10090 & n4933;
  assign n5009 = ~n5007 & ~n5008;
  assign n5010 = ~n5006 & n5009;
  assign n5011 = ~n4913 & n5010;
  assign n5012 = ~n10115 & n5010;
  assign n5013 = ~n5011 & ~n5012;
  assign n5014 = ~n5005 & n5010;
  assign n5015 = ~n9626 & ~n10116;
  assign n5016 = n9626 & n10116;
  assign n5017 = ~n5015 & ~n5016;
  assign n5018 = n10114 & n5017;
  assign n5019 = n10114 & ~n10116;
  assign n5020 = n4974 & n10117;
  assign n5021 = ~n4773 & n10091;
  assign n5022 = ~n10091 & ~n10092;
  assign n5023 = ~n4772 & n4790;
  assign n5024 = ~n5022 & ~n5023;
  assign n5025 = ~n10092 & ~n5021;
  assign n5026 = n4913 & ~n10118;
  assign n5027 = n4764 & n4920;
  assign n5028 = ~n10089 & n4933;
  assign n5029 = ~n10090 & n10106;
  assign n5030 = ~n5028 & ~n5029;
  assign n5031 = ~n5027 & ~n5029;
  assign n5032 = ~n5028 & n5031;
  assign n5033 = ~n5027 & n5030;
  assign n5034 = ~n5026 & n10119;
  assign n5035 = n9626 & ~n5034;
  assign n5036 = ~n9626 & n5034;
  assign n5037 = ~n5035 & ~n5036;
  assign n5038 = ~n4974 & ~n10117;
  assign n5039 = n10117 & ~n5020;
  assign n5040 = ~n4974 & n10117;
  assign n5041 = n4974 & ~n5020;
  assign n5042 = n4974 & ~n10117;
  assign n5043 = ~n10120 & ~n10121;
  assign n5044 = ~n5020 & ~n5038;
  assign n5045 = n5037 & ~n10122;
  assign n5046 = ~n5020 & ~n5045;
  assign n5047 = ~n4945 & ~n10113;
  assign n5048 = ~n4986 & ~n5047;
  assign n5049 = ~n5046 & n5048;
  assign n5050 = ~n4986 & ~n5049;
  assign n5051 = n4796 & ~n4798;
  assign n5052 = ~n4799 & ~n5051;
  assign n5053 = n4913 & n5052;
  assign n5054 = ~n10088 & n4920;
  assign n5055 = n4764 & n10106;
  assign n5056 = n4761 & n4933;
  assign n5057 = ~n5055 & ~n5056;
  assign n5058 = ~n5054 & n5057;
  assign n5059 = ~n5053 & n5058;
  assign n5060 = n9626 & ~n5059;
  assign n5061 = ~n9626 & n5059;
  assign n5062 = ~n5060 & ~n5061;
  assign n5063 = ~n1164 & ~n4975;
  assign n5064 = n4958 & n10115;
  assign n5065 = ~n10089 & n4968;
  assign n5066 = n10109 & n10111;
  assign n5067 = ~n10079 & n10109;
  assign n5068 = n10111 & n5067;
  assign n5069 = ~n10079 & n5066;
  assign n5070 = ~n4775 & n10123;
  assign n5071 = ~n10090 & n4966;
  assign n5072 = ~n5070 & ~n5071;
  assign n5073 = ~n5065 & n5072;
  assign n5074 = ~n4958 & n5073;
  assign n5075 = ~n10115 & n5073;
  assign n5076 = ~n5074 & ~n5075;
  assign n5077 = ~n5064 & n5073;
  assign n5078 = n5063 & n10124;
  assign n5079 = ~n5063 & ~n10124;
  assign n5080 = n4975 & ~n10124;
  assign n5081 = ~n1164 & n5080;
  assign n5082 = n1164 & ~n10124;
  assign n5083 = ~n1164 & n10124;
  assign n5084 = ~n5082 & ~n5083;
  assign n5085 = n10112 & n5084;
  assign n5086 = n10112 & ~n10124;
  assign n5087 = ~n10112 & ~n5084;
  assign n5088 = ~n10125 & ~n5087;
  assign n5089 = ~n5078 & ~n5079;
  assign n5090 = n5062 & n10126;
  assign n5091 = ~n5062 & ~n10126;
  assign n5092 = ~n5090 & ~n5091;
  assign n5093 = n5050 & ~n5092;
  assign n5094 = ~n5050 & n5092;
  assign n5095 = ~n5093 & ~n5094;
  assign n5096 = n9528 & ~n2130;
  assign n5097 = ~n9528 & n2130;
  assign n5098 = ~n9528 & ~n2130;
  assign n5099 = n9528 & n2130;
  assign n5100 = ~n5098 & ~n5099;
  assign n5101 = ~n5096 & ~n5097;
  assign n5102 = n9686 & ~n1703;
  assign n5103 = ~n9686 & n1703;
  assign n5104 = ~n9686 & ~n1703;
  assign n5105 = n9686 & n1703;
  assign n5106 = ~n5104 & ~n5105;
  assign n5107 = ~n5102 & ~n5103;
  assign n5108 = ~n10127 & ~n10128;
  assign n5109 = n4808 & ~n4810;
  assign n5110 = ~n4811 & ~n5109;
  assign n5111 = n5108 & n5110;
  assign n5112 = ~n10127 & n10128;
  assign n5113 = n4740 & n5112;
  assign n5114 = n9686 & ~n2130;
  assign n5115 = ~n9686 & n2130;
  assign n5116 = ~n9686 & ~n2130;
  assign n5117 = n9686 & n2130;
  assign n5118 = ~n5116 & ~n5117;
  assign n5119 = ~n5114 & ~n5115;
  assign n5120 = n10127 & ~n10129;
  assign n5121 = ~n10086 & n5120;
  assign n5122 = n10127 & n10129;
  assign n5123 = n10127 & ~n10128;
  assign n5124 = n10129 & n5123;
  assign n5125 = ~n10128 & n5122;
  assign n5126 = ~n10087 & n10130;
  assign n5127 = ~n5121 & ~n5126;
  assign n5128 = ~n5113 & ~n5126;
  assign n5129 = ~n5121 & n5128;
  assign n5130 = ~n5113 & n5127;
  assign n5131 = ~n5110 & n10131;
  assign n5132 = ~n5108 & n10131;
  assign n5133 = ~n5131 & ~n5132;
  assign n5134 = ~n5111 & n10131;
  assign n5135 = n1703 & ~n10132;
  assign n5136 = ~n1703 & n10132;
  assign n5137 = ~n5135 & ~n5136;
  assign n5138 = n5095 & n5137;
  assign n5139 = ~n5095 & ~n5137;
  assign n5140 = n5095 & ~n5138;
  assign n5141 = n5137 & ~n5138;
  assign n5142 = ~n5140 & ~n5141;
  assign n5143 = ~n5138 & ~n5139;
  assign n5144 = n4804 & ~n4806;
  assign n5145 = ~n4807 & ~n5144;
  assign n5146 = n5108 & n5145;
  assign n5147 = ~n10086 & n5112;
  assign n5148 = ~n10088 & n10130;
  assign n5149 = ~n10087 & n5120;
  assign n5150 = ~n5148 & ~n5149;
  assign n5151 = ~n5147 & n5150;
  assign n5152 = ~n5146 & n5151;
  assign n5153 = ~n1703 & ~n5152;
  assign n5154 = ~n5152 & ~n5153;
  assign n5155 = n1703 & ~n5152;
  assign n5156 = ~n1703 & ~n5153;
  assign n5157 = ~n1703 & n5152;
  assign n5158 = ~n10134 & ~n10135;
  assign n5159 = n5046 & ~n5048;
  assign n5160 = ~n5049 & ~n5159;
  assign n5161 = n5158 & ~n5160;
  assign n5162 = ~n5158 & n5160;
  assign n5163 = n4800 & ~n4802;
  assign n5164 = ~n4803 & ~n5163;
  assign n5165 = n5108 & n5164;
  assign n5166 = ~n10087 & n5112;
  assign n5167 = n4761 & n10130;
  assign n5168 = ~n10088 & n5120;
  assign n5169 = ~n5167 & ~n5168;
  assign n5170 = ~n5166 & n5169;
  assign n5171 = ~n5164 & n5170;
  assign n5172 = ~n5108 & n5170;
  assign n5173 = ~n5171 & ~n5172;
  assign n5174 = ~n5165 & n5170;
  assign n5175 = n1703 & ~n10136;
  assign n5176 = ~n1703 & n10136;
  assign n5177 = ~n5175 & ~n5176;
  assign n5178 = ~n5037 & n10122;
  assign n5179 = ~n10122 & ~n5045;
  assign n5180 = ~n5037 & ~n10122;
  assign n5181 = n5037 & ~n5045;
  assign n5182 = n5037 & n10122;
  assign n5183 = ~n10137 & ~n10138;
  assign n5184 = ~n5045 & ~n5178;
  assign n5185 = n5177 & ~n10139;
  assign n5186 = ~n5177 & n10139;
  assign n5187 = ~n10139 & ~n5185;
  assign n5188 = ~n5177 & ~n10139;
  assign n5189 = n5177 & ~n5185;
  assign n5190 = n5177 & n10139;
  assign n5191 = ~n10140 & ~n10141;
  assign n5192 = ~n5185 & ~n5186;
  assign n5193 = n5052 & n5108;
  assign n5194 = ~n10088 & n5112;
  assign n5195 = n4764 & n10130;
  assign n5196 = n4761 & n5120;
  assign n5197 = ~n5195 & ~n5196;
  assign n5198 = ~n5194 & n5197;
  assign n5199 = ~n5193 & n5198;
  assign n5200 = ~n1703 & ~n5199;
  assign n5201 = ~n5199 & ~n5200;
  assign n5202 = n1703 & ~n5199;
  assign n5203 = ~n1703 & ~n5200;
  assign n5204 = ~n1703 & n5199;
  assign n5205 = ~n10143 & ~n10144;
  assign n5206 = n9626 & ~n10114;
  assign n5207 = n10116 & n5206;
  assign n5208 = ~n10116 & ~n5206;
  assign n5209 = ~n10114 & ~n5017;
  assign n5210 = ~n10117 & ~n5209;
  assign n5211 = ~n5207 & ~n5208;
  assign n5212 = n5205 & ~n10145;
  assign n5213 = ~n5205 & n10145;
  assign n5214 = ~n10104 & n5108;
  assign n5215 = n4761 & n5112;
  assign n5216 = ~n10089 & n10130;
  assign n5217 = n4764 & n5120;
  assign n5218 = ~n5216 & ~n5217;
  assign n5219 = ~n5215 & ~n5217;
  assign n5220 = ~n5216 & n5219;
  assign n5221 = ~n5215 & n5218;
  assign n5222 = ~n5108 & n10146;
  assign n5223 = n10104 & n10146;
  assign n5224 = ~n5222 & ~n5223;
  assign n5225 = ~n5214 & n10146;
  assign n5226 = n1703 & ~n10147;
  assign n5227 = ~n1703 & n10147;
  assign n5228 = ~n5226 & ~n5227;
  assign n5229 = n9626 & n4992;
  assign n5230 = ~n4991 & n5229;
  assign n5231 = n4991 & ~n5229;
  assign n5232 = ~n4993 & ~n4996;
  assign n5233 = ~n10114 & ~n5232;
  assign n5234 = ~n5230 & ~n5231;
  assign n5235 = n5228 & n10148;
  assign n5236 = ~n4957 & n5108;
  assign n5237 = ~n4775 & n5120;
  assign n5238 = ~n10090 & n5112;
  assign n5239 = ~n5237 & ~n5238;
  assign n5240 = ~n5236 & n5239;
  assign n5241 = ~n4775 & ~n10127;
  assign n5242 = ~n1703 & ~n5241;
  assign n5243 = ~n1703 & ~n5240;
  assign n5244 = ~n1703 & ~n5243;
  assign n5245 = ~n5240 & ~n5243;
  assign n5246 = ~n5244 & ~n5245;
  assign n5247 = n5242 & ~n5246;
  assign n5248 = n5240 & n5242;
  assign n5249 = n10115 & n5108;
  assign n5250 = ~n10089 & n5112;
  assign n5251 = ~n4775 & n10130;
  assign n5252 = ~n10090 & n5120;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = ~n5250 & n5253;
  assign n5255 = ~n10115 & n5254;
  assign n5256 = ~n5108 & n5254;
  assign n5257 = ~n5255 & ~n5256;
  assign n5258 = ~n5249 & n5254;
  assign n5259 = n1703 & ~n10150;
  assign n5260 = ~n1703 & n10150;
  assign n5261 = ~n5259 & ~n5260;
  assign n5262 = n10149 & n5261;
  assign n5263 = n10149 & ~n10150;
  assign n5264 = n4992 & n10151;
  assign n5265 = ~n10118 & n5108;
  assign n5266 = n4764 & n5112;
  assign n5267 = ~n10089 & n5120;
  assign n5268 = ~n10090 & n10130;
  assign n5269 = ~n5267 & ~n5268;
  assign n5270 = ~n5266 & ~n5268;
  assign n5271 = ~n5267 & n5270;
  assign n5272 = ~n5266 & n5269;
  assign n5273 = ~n5265 & n10152;
  assign n5274 = ~n1703 & ~n5273;
  assign n5275 = ~n1703 & ~n5274;
  assign n5276 = ~n1703 & n5273;
  assign n5277 = ~n5273 & ~n5274;
  assign n5278 = n1703 & ~n5273;
  assign n5279 = ~n10153 & ~n10154;
  assign n5280 = ~n4992 & ~n10151;
  assign n5281 = n10151 & ~n5264;
  assign n5282 = ~n4992 & n10151;
  assign n5283 = n4992 & ~n5264;
  assign n5284 = n4992 & ~n10151;
  assign n5285 = ~n10155 & ~n10156;
  assign n5286 = ~n5264 & ~n5280;
  assign n5287 = ~n5279 & ~n10157;
  assign n5288 = ~n5264 & ~n5287;
  assign n5289 = ~n5228 & ~n10148;
  assign n5290 = ~n5235 & ~n5289;
  assign n5291 = ~n5288 & n5290;
  assign n5292 = ~n5235 & ~n5291;
  assign n5293 = ~n5213 & n5292;
  assign n5294 = ~n5205 & ~n5213;
  assign n5295 = n10145 & ~n5213;
  assign n5296 = ~n5294 & ~n5295;
  assign n5297 = ~n5212 & ~n5213;
  assign n5298 = ~n5292 & ~n10158;
  assign n5299 = ~n5213 & ~n5298;
  assign n5300 = ~n5212 & ~n5293;
  assign n5301 = ~n10142 & ~n10159;
  assign n5302 = ~n5185 & ~n5301;
  assign n5303 = ~n5162 & n5302;
  assign n5304 = ~n5158 & ~n5162;
  assign n5305 = n5160 & ~n5162;
  assign n5306 = ~n5304 & ~n5305;
  assign n5307 = ~n5161 & ~n5162;
  assign n5308 = ~n5302 & ~n10160;
  assign n5309 = ~n5162 & ~n5308;
  assign n5310 = ~n5161 & ~n5303;
  assign n5311 = ~n10133 & ~n10161;
  assign n5312 = ~n5138 & ~n5311;
  assign n5313 = ~n5090 & ~n5094;
  assign n5314 = n4913 & n5164;
  assign n5315 = ~n10087 & n4920;
  assign n5316 = n4761 & n10106;
  assign n5317 = ~n10088 & n4933;
  assign n5318 = ~n5316 & ~n5317;
  assign n5319 = ~n5315 & n5318;
  assign n5320 = ~n5314 & n5319;
  assign n5321 = n9626 & ~n5320;
  assign n5322 = ~n9626 & n5320;
  assign n5323 = ~n5321 & ~n5322;
  assign n5324 = ~n4952 & ~n10125;
  assign n5325 = n4952 & n5080;
  assign n5326 = n4952 & n10125;
  assign n5327 = ~n4775 & n10125;
  assign n5328 = ~n5324 & ~n10162;
  assign n5329 = ~n1164 & ~n5328;
  assign n5330 = n4958 & ~n10118;
  assign n5331 = n4764 & n4968;
  assign n5332 = ~n10089 & n4966;
  assign n5333 = ~n10090 & n10123;
  assign n5334 = ~n5332 & ~n5333;
  assign n5335 = ~n5331 & ~n5333;
  assign n5336 = ~n5332 & n5335;
  assign n5337 = ~n5331 & n5334;
  assign n5338 = ~n5330 & n10163;
  assign n5339 = n5329 & ~n5338;
  assign n5340 = ~n5329 & n5338;
  assign n5341 = ~n1164 & ~n5338;
  assign n5342 = ~n5338 & ~n5341;
  assign n5343 = n1164 & ~n5338;
  assign n5344 = ~n1164 & ~n5341;
  assign n5345 = ~n1164 & n5338;
  assign n5346 = ~n10164 & ~n10165;
  assign n5347 = ~n10162 & ~n5346;
  assign n5348 = ~n5324 & n5347;
  assign n5349 = n5328 & ~n5346;
  assign n5350 = ~n5328 & n5346;
  assign n5351 = ~n10166 & ~n5350;
  assign n5352 = ~n5346 & ~n10166;
  assign n5353 = ~n10162 & ~n10166;
  assign n5354 = ~n5324 & n5338;
  assign n5355 = ~n5324 & n10168;
  assign n5356 = ~n5352 & ~n5355;
  assign n5357 = ~n5339 & ~n5340;
  assign n5358 = n5323 & n10167;
  assign n5359 = ~n5323 & ~n10167;
  assign n5360 = n5323 & ~n5358;
  assign n5361 = n10167 & ~n5358;
  assign n5362 = ~n5360 & ~n5361;
  assign n5363 = ~n5358 & ~n5359;
  assign n5364 = n5313 & n10169;
  assign n5365 = ~n5313 & ~n10169;
  assign n5366 = ~n5364 & ~n5365;
  assign n5367 = n4812 & ~n4814;
  assign n5368 = ~n4815 & ~n5367;
  assign n5369 = n5108 & n5368;
  assign n5370 = ~n10085 & n5112;
  assign n5371 = ~n10086 & n10130;
  assign n5372 = n4740 & n5120;
  assign n5373 = ~n5371 & ~n5372;
  assign n5374 = ~n5370 & n5373;
  assign n5375 = ~n5368 & n5374;
  assign n5376 = ~n5108 & n5374;
  assign n5377 = ~n5375 & ~n5376;
  assign n5378 = ~n5369 & n5374;
  assign n5379 = n1703 & ~n10170;
  assign n5380 = ~n1703 & n10170;
  assign n5381 = ~n5379 & ~n5380;
  assign n5382 = n5366 & n5381;
  assign n5383 = ~n5366 & ~n5381;
  assign n5384 = n5366 & ~n5382;
  assign n5385 = n5381 & ~n5382;
  assign n5386 = ~n5384 & ~n5385;
  assign n5387 = ~n5382 & ~n5383;
  assign n5388 = ~n5312 & ~n10171;
  assign n5389 = n5312 & n10171;
  assign n5390 = ~n5312 & ~n5388;
  assign n5391 = ~n10171 & ~n5388;
  assign n5392 = ~n5390 & ~n5391;
  assign n5393 = ~n5388 & ~n5389;
  assign n5394 = n4900 & ~n10172;
  assign n5395 = n4820 & ~n4822;
  assign n5396 = ~n4823 & ~n5395;
  assign n5397 = n90 & n5396;
  assign n5398 = ~n10084 & n4878;
  assign n5399 = ~n10085 & n10100;
  assign n5400 = n4731 & n4886;
  assign n5401 = ~n5399 & ~n5400;
  assign n5402 = ~n5398 & n5401;
  assign n5403 = ~n5397 & n5402;
  assign n5404 = n9528 & ~n5403;
  assign n5405 = ~n9528 & n5403;
  assign n5406 = ~n5404 & ~n5405;
  assign n5407 = n10133 & n10161;
  assign n5408 = ~n10161 & ~n5311;
  assign n5409 = ~n10133 & ~n5311;
  assign n5410 = ~n5408 & ~n5409;
  assign n5411 = ~n5311 & ~n5407;
  assign n5412 = n5406 & ~n10173;
  assign n5413 = n4816 & ~n4818;
  assign n5414 = ~n4819 & ~n5413;
  assign n5415 = n90 & n5414;
  assign n5416 = n4731 & n4878;
  assign n5417 = ~n10085 & n4886;
  assign n5418 = n4740 & n10100;
  assign n5419 = ~n5417 & ~n5418;
  assign n5420 = ~n5416 & ~n5418;
  assign n5421 = ~n5417 & n5420;
  assign n5422 = ~n5416 & n5419;
  assign n5423 = ~n90 & n10174;
  assign n5424 = ~n5414 & n10174;
  assign n5425 = ~n5423 & ~n5424;
  assign n5426 = ~n5415 & n10174;
  assign n5427 = ~n9528 & ~n10175;
  assign n5428 = n9528 & n10175;
  assign n5429 = ~n5427 & ~n5428;
  assign n5430 = n5302 & ~n10160;
  assign n5431 = ~n5302 & n10160;
  assign n5432 = ~n5430 & ~n5431;
  assign n5433 = n5429 & ~n5432;
  assign n5434 = n90 & n5368;
  assign n5435 = ~n10085 & n4878;
  assign n5436 = ~n10086 & n10100;
  assign n5437 = n4740 & n4886;
  assign n5438 = ~n5436 & ~n5437;
  assign n5439 = ~n5435 & n5438;
  assign n5440 = ~n90 & n5439;
  assign n5441 = ~n5368 & n5439;
  assign n5442 = ~n5440 & ~n5441;
  assign n5443 = ~n5434 & n5439;
  assign n5444 = ~n9528 & ~n10176;
  assign n5445 = n9528 & n10176;
  assign n5446 = ~n5444 & ~n5445;
  assign n5447 = n10142 & n10159;
  assign n5448 = ~n10159 & ~n5301;
  assign n5449 = n10142 & ~n10159;
  assign n5450 = ~n10142 & ~n5301;
  assign n5451 = ~n10142 & n10159;
  assign n5452 = ~n10177 & ~n10178;
  assign n5453 = ~n5301 & ~n5447;
  assign n5454 = n5446 & ~n10179;
  assign n5455 = n90 & n5110;
  assign n5456 = n4740 & n4878;
  assign n5457 = ~n10086 & n4886;
  assign n5458 = ~n10087 & n10100;
  assign n5459 = ~n5457 & ~n5458;
  assign n5460 = ~n5456 & ~n5458;
  assign n5461 = ~n5457 & n5460;
  assign n5462 = ~n5456 & n5459;
  assign n5463 = ~n90 & n10180;
  assign n5464 = ~n5110 & n10180;
  assign n5465 = ~n5463 & ~n5464;
  assign n5466 = ~n5455 & n10180;
  assign n5467 = ~n9528 & ~n10181;
  assign n5468 = n9528 & n10181;
  assign n5469 = ~n5467 & ~n5468;
  assign n5470 = n5292 & ~n10158;
  assign n5471 = ~n5292 & n10158;
  assign n5472 = ~n5470 & ~n5471;
  assign n5473 = n5469 & ~n5472;
  assign n5474 = n90 & n5145;
  assign n5475 = ~n10086 & n4878;
  assign n5476 = ~n10088 & n10100;
  assign n5477 = ~n10087 & n4886;
  assign n5478 = ~n5476 & ~n5477;
  assign n5479 = ~n5475 & n5478;
  assign n5480 = ~n5474 & n5479;
  assign n5481 = n9528 & ~n5480;
  assign n5482 = ~n9528 & n5480;
  assign n5483 = ~n5481 & ~n5482;
  assign n5484 = n5288 & ~n5290;
  assign n5485 = ~n5291 & ~n5484;
  assign n5486 = n5483 & n5485;
  assign n5487 = n90 & n5164;
  assign n5488 = ~n10087 & n4878;
  assign n5489 = n4761 & n10100;
  assign n5490 = ~n10088 & n4886;
  assign n5491 = ~n5489 & ~n5490;
  assign n5492 = ~n5488 & n5491;
  assign n5493 = ~n90 & n5492;
  assign n5494 = ~n5164 & n5492;
  assign n5495 = ~n5493 & ~n5494;
  assign n5496 = ~n5487 & n5492;
  assign n5497 = ~n9528 & ~n10182;
  assign n5498 = n9528 & n10182;
  assign n5499 = ~n5497 & ~n5498;
  assign n5500 = n5279 & n10157;
  assign n5501 = ~n10157 & ~n5287;
  assign n5502 = ~n5279 & ~n5287;
  assign n5503 = ~n5501 & ~n5502;
  assign n5504 = ~n5287 & ~n5500;
  assign n5505 = n5499 & ~n10183;
  assign n5506 = n90 & n5052;
  assign n5507 = ~n10088 & n4878;
  assign n5508 = n4764 & n10100;
  assign n5509 = n4761 & n4886;
  assign n5510 = ~n5508 & ~n5509;
  assign n5511 = ~n5507 & n5510;
  assign n5512 = ~n5506 & n5511;
  assign n5513 = n9528 & ~n5512;
  assign n5514 = ~n9528 & n5512;
  assign n5515 = ~n5513 & ~n5514;
  assign n5516 = ~n1703 & ~n10149;
  assign n5517 = n10150 & n5516;
  assign n5518 = ~n10150 & ~n5516;
  assign n5519 = ~n10149 & ~n5261;
  assign n5520 = ~n10151 & ~n5519;
  assign n5521 = ~n5517 & ~n5518;
  assign n5522 = n5515 & n10184;
  assign n5523 = n90 & ~n10104;
  assign n5524 = n4761 & n4878;
  assign n5525 = ~n10089 & n10100;
  assign n5526 = n4764 & n4886;
  assign n5527 = ~n5525 & ~n5526;
  assign n5528 = ~n5524 & ~n5526;
  assign n5529 = ~n5525 & n5528;
  assign n5530 = ~n5524 & n5527;
  assign n5531 = ~n90 & n10185;
  assign n5532 = n10104 & n10185;
  assign n5533 = ~n5531 & ~n5532;
  assign n5534 = ~n5523 & n10185;
  assign n5535 = ~n9528 & ~n10186;
  assign n5536 = n9528 & n10186;
  assign n5537 = ~n5535 & ~n5536;
  assign n5538 = ~n1703 & n5241;
  assign n5539 = ~n5240 & n5538;
  assign n5540 = n5240 & ~n5538;
  assign n5541 = ~n5242 & n5246;
  assign n5542 = ~n10149 & ~n5541;
  assign n5543 = ~n5539 & ~n5540;
  assign n5544 = n5537 & n10187;
  assign n5545 = n90 & ~n4957;
  assign n5546 = ~n4775 & n4886;
  assign n5547 = ~n10090 & n4878;
  assign n5548 = ~n5546 & ~n5547;
  assign n5549 = ~n5545 & n5548;
  assign n5550 = ~n9530 & ~n4775;
  assign n5551 = n9528 & ~n5550;
  assign n5552 = n9528 & ~n5549;
  assign n5553 = ~n9528 & n5549;
  assign n5554 = ~n5552 & ~n5553;
  assign n5555 = n5551 & n5554;
  assign n5556 = n5549 & n5551;
  assign n5557 = n90 & n10115;
  assign n5558 = ~n10089 & n4878;
  assign n5559 = ~n4775 & n10100;
  assign n5560 = ~n10090 & n4886;
  assign n5561 = ~n5559 & ~n5560;
  assign n5562 = ~n5558 & n5561;
  assign n5563 = ~n90 & n5562;
  assign n5564 = ~n10115 & n5562;
  assign n5565 = ~n5563 & ~n5564;
  assign n5566 = ~n5557 & n5562;
  assign n5567 = ~n9528 & ~n10189;
  assign n5568 = n9528 & n10189;
  assign n5569 = ~n5567 & ~n5568;
  assign n5570 = n10188 & n5569;
  assign n5571 = n10188 & ~n10189;
  assign n5572 = n5241 & n10190;
  assign n5573 = n90 & ~n10118;
  assign n5574 = n4764 & n4878;
  assign n5575 = ~n10089 & n4886;
  assign n5576 = ~n10090 & n10100;
  assign n5577 = ~n5575 & ~n5576;
  assign n5578 = ~n5574 & ~n5576;
  assign n5579 = ~n5575 & n5578;
  assign n5580 = ~n5574 & n5577;
  assign n5581 = ~n5573 & n10191;
  assign n5582 = n9528 & ~n5581;
  assign n5583 = ~n9528 & n5581;
  assign n5584 = ~n5582 & ~n5583;
  assign n5585 = ~n5241 & ~n10190;
  assign n5586 = n10190 & ~n5572;
  assign n5587 = ~n5241 & n10190;
  assign n5588 = n5241 & ~n5572;
  assign n5589 = n5241 & ~n10190;
  assign n5590 = ~n10192 & ~n10193;
  assign n5591 = ~n5572 & ~n5585;
  assign n5592 = n5584 & ~n10194;
  assign n5593 = ~n5572 & ~n5592;
  assign n5594 = ~n5537 & ~n10187;
  assign n5595 = ~n5544 & ~n5594;
  assign n5596 = ~n5593 & n5595;
  assign n5597 = ~n5544 & ~n5596;
  assign n5598 = ~n5515 & ~n10184;
  assign n5599 = ~n5522 & ~n5598;
  assign n5600 = ~n5597 & n5599;
  assign n5601 = ~n5522 & ~n5600;
  assign n5602 = ~n5499 & n10183;
  assign n5603 = ~n10183 & ~n5505;
  assign n5604 = n5499 & ~n5505;
  assign n5605 = ~n5603 & ~n5604;
  assign n5606 = ~n5505 & ~n5602;
  assign n5607 = ~n5601 & ~n10195;
  assign n5608 = ~n5505 & ~n5607;
  assign n5609 = ~n5483 & ~n5485;
  assign n5610 = ~n5486 & ~n5609;
  assign n5611 = ~n5608 & n5610;
  assign n5612 = ~n5486 & ~n5611;
  assign n5613 = ~n5469 & n5472;
  assign n5614 = ~n5472 & ~n5473;
  assign n5615 = n5469 & ~n5473;
  assign n5616 = ~n5614 & ~n5615;
  assign n5617 = ~n5473 & ~n5613;
  assign n5618 = ~n5612 & ~n10196;
  assign n5619 = ~n5473 & ~n5618;
  assign n5620 = ~n5446 & n10179;
  assign n5621 = ~n10179 & ~n5454;
  assign n5622 = ~n5446 & ~n10179;
  assign n5623 = n5446 & ~n5454;
  assign n5624 = n5446 & n10179;
  assign n5625 = ~n10197 & ~n10198;
  assign n5626 = ~n5454 & ~n5620;
  assign n5627 = ~n5619 & ~n10199;
  assign n5628 = ~n5454 & ~n5627;
  assign n5629 = ~n5429 & n5432;
  assign n5630 = ~n5433 & ~n5629;
  assign n5631 = ~n5628 & n5630;
  assign n5632 = ~n5433 & ~n5631;
  assign n5633 = ~n5406 & n10173;
  assign n5634 = n5406 & ~n5412;
  assign n5635 = ~n10173 & ~n5412;
  assign n5636 = ~n5634 & ~n5635;
  assign n5637 = ~n5412 & ~n5633;
  assign n5638 = ~n5632 & ~n10200;
  assign n5639 = ~n5412 & ~n5638;
  assign n5640 = ~n4900 & n10172;
  assign n5641 = n4900 & ~n5394;
  assign n5642 = ~n10172 & ~n5394;
  assign n5643 = ~n5641 & ~n5642;
  assign n5644 = ~n5394 & ~n5640;
  assign n5645 = ~n5639 & ~n10201;
  assign n5646 = ~n5394 & ~n5645;
  assign n5647 = ~n4871 & ~n4874;
  assign n5648 = ~n574 & ~n674;
  assign n5649 = ~n574 & n777;
  assign n5650 = ~n674 & n5649;
  assign n5651 = n777 & n5648;
  assign n5652 = ~n626 & ~n715;
  assign n5653 = ~n9586 & ~n990;
  assign n5654 = n5652 & n5653;
  assign n5655 = n9975 & n5654;
  assign n5656 = n10202 & n5655;
  assign n5657 = ~n217 & ~n682;
  assign n5658 = ~n217 & ~n262;
  assign n5659 = ~n682 & n5658;
  assign n5660 = ~n262 & n5657;
  assign n5661 = ~n9544 & ~n682;
  assign n5662 = ~n262 & ~n682;
  assign n5663 = ~n9544 & n5662;
  assign n5664 = ~n262 & n5661;
  assign n5665 = ~n217 & n10204;
  assign n5666 = ~n9696 & n5665;
  assign n5667 = ~n217 & ~n9696;
  assign n5668 = n10204 & n5667;
  assign n5669 = n4568 & n10203;
  assign n5670 = ~n1037 & ~n1108;
  assign n5671 = ~n258 & ~n536;
  assign n5672 = ~n249 & ~n770;
  assign n5673 = n5671 & n5672;
  assign n5674 = n5670 & n5673;
  assign n5675 = n10205 & n5674;
  assign n5676 = n10202 & n10205;
  assign n5677 = n9975 & n5676;
  assign n5678 = ~n626 & n5677;
  assign n5679 = ~n249 & n5678;
  assign n5680 = ~n990 & n5679;
  assign n5681 = ~n715 & n5680;
  assign n5682 = ~n9586 & n5681;
  assign n5683 = ~n1108 & n5682;
  assign n5684 = ~n258 & n5683;
  assign n5685 = ~n770 & n5684;
  assign n5686 = ~n536 & n5685;
  assign n5687 = ~n1037 & n5686;
  assign n5688 = ~n626 & ~n770;
  assign n5689 = n5653 & n5688;
  assign n5690 = n9975 & n5689;
  assign n5691 = n10202 & n5690;
  assign n5692 = ~n249 & ~n715;
  assign n5693 = n5671 & n5692;
  assign n5694 = n5670 & n5693;
  assign n5695 = n10205 & n5694;
  assign n5696 = n5691 & n5695;
  assign n5697 = ~n770 & ~n990;
  assign n5698 = n5692 & n5697;
  assign n5699 = n9975 & n5698;
  assign n5700 = n10202 & n5699;
  assign n5701 = ~n9586 & ~n626;
  assign n5702 = n5671 & n5701;
  assign n5703 = n5670 & n5702;
  assign n5704 = n10205 & n5703;
  assign n5705 = n5700 & n5704;
  assign n5706 = ~n715 & ~n770;
  assign n5707 = n5701 & n5706;
  assign n5708 = n9975 & n5707;
  assign n5709 = n10202 & n5708;
  assign n5710 = ~n249 & ~n990;
  assign n5711 = n5670 & n5710;
  assign n5712 = n5671 & n5711;
  assign n5713 = n10205 & n5712;
  assign n5714 = n5709 & n5713;
  assign n5715 = n5656 & n5675;
  assign n5716 = ~n9562 & ~n534;
  assign n5717 = ~n9562 & ~n898;
  assign n5718 = ~n534 & n5717;
  assign n5719 = ~n534 & ~n898;
  assign n5720 = ~n9562 & n5719;
  assign n5721 = ~n898 & n5716;
  assign n5722 = ~n215 & ~n9555;
  assign n5723 = ~n781 & ~n995;
  assign n5724 = n5722 & n5723;
  assign n5725 = n10032 & n5724;
  assign n5726 = n10207 & n5725;
  assign n5727 = ~n199 & ~n386;
  assign n5728 = n385 & n4510;
  assign n5729 = n5727 & n5728;
  assign n5730 = n9576 & n5729;
  assign n5731 = ~n995 & ~n1083;
  assign n5732 = n5722 & n5731;
  assign n5733 = n10032 & n5732;
  assign n5734 = n10207 & n5733;
  assign n5735 = ~n334 & ~n781;
  assign n5736 = n385 & n5735;
  assign n5737 = n5727 & n5736;
  assign n5738 = n9576 & n5737;
  assign n5739 = n5734 & n5738;
  assign n5740 = ~n9555 & ~n1083;
  assign n5741 = n5723 & n5740;
  assign n5742 = n10207 & n5741;
  assign n5743 = n10032 & n5742;
  assign n5744 = ~n334 & ~n386;
  assign n5745 = ~n199 & ~n215;
  assign n5746 = n5744 & n5745;
  assign n5747 = n385 & n5746;
  assign n5748 = n9576 & n5747;
  assign n5749 = n5743 & n5748;
  assign n5750 = n5726 & n5730;
  assign n5751 = n9575 & n10208;
  assign n5752 = n9576 & n10032;
  assign n5753 = n385 & n5752;
  assign n5754 = n9575 & n5753;
  assign n5755 = n10206 & n5754;
  assign n5756 = n10207 & n5755;
  assign n5757 = ~n386 & n5756;
  assign n5758 = ~n334 & n5757;
  assign n5759 = ~n215 & n5758;
  assign n5760 = ~n9555 & n5759;
  assign n5761 = ~n199 & n5760;
  assign n5762 = ~n995 & n5761;
  assign n5763 = ~n1083 & n5762;
  assign n5764 = ~n781 & n5763;
  assign n5765 = n10206 & n5751;
  assign n5766 = n4868 & n10209;
  assign n5767 = ~n4868 & ~n10209;
  assign n5768 = ~n4868 & n10209;
  assign n5769 = n4868 & ~n10209;
  assign n5770 = ~n5768 & ~n5769;
  assign n5771 = ~n5766 & ~n5767;
  assign n5772 = ~n4870 & n10210;
  assign n5773 = n4870 & ~n10210;
  assign n5774 = n4870 & n10209;
  assign n5775 = ~n5772 & ~n10211;
  assign n5776 = ~n5647 & n5775;
  assign n5777 = n5647 & ~n5775;
  assign n5778 = ~n5776 & ~n5777;
  assign n5779 = n90 & n5778;
  assign n5780 = n4878 & n10210;
  assign n5781 = ~n10084 & n10100;
  assign n5782 = ~n4870 & n4886;
  assign n5783 = ~n5781 & ~n5782;
  assign n5784 = ~n5780 & n5783;
  assign n5785 = ~n5779 & n5784;
  assign n5786 = n9528 & ~n5785;
  assign n5787 = ~n9528 & n5785;
  assign n5788 = ~n5786 & ~n5787;
  assign n5789 = ~n5382 & ~n5388;
  assign n5790 = n5108 & n5414;
  assign n5791 = n4731 & n5112;
  assign n5792 = ~n10085 & n5120;
  assign n5793 = n4740 & n10130;
  assign n5794 = ~n5792 & ~n5793;
  assign n5795 = ~n5791 & ~n5793;
  assign n5796 = ~n5792 & n5795;
  assign n5797 = ~n5791 & n5794;
  assign n5798 = ~n5414 & n10212;
  assign n5799 = ~n5108 & n10212;
  assign n5800 = ~n5798 & ~n5799;
  assign n5801 = ~n5790 & n10212;
  assign n5802 = n1703 & ~n10213;
  assign n5803 = ~n1703 & n10213;
  assign n5804 = ~n5802 & ~n5803;
  assign n5805 = ~n5358 & ~n5365;
  assign n5806 = n4913 & n5145;
  assign n5807 = ~n10086 & n4920;
  assign n5808 = ~n10088 & n10106;
  assign n5809 = ~n10087 & n4933;
  assign n5810 = ~n5808 & ~n5809;
  assign n5811 = ~n5807 & n5810;
  assign n5812 = ~n5806 & n5811;
  assign n5813 = n9626 & ~n5812;
  assign n5814 = ~n9626 & n5812;
  assign n5815 = ~n5813 & ~n5814;
  assign n5816 = ~n1164 & n10090;
  assign n5817 = ~n10104 & n4958;
  assign n5818 = n4761 & n4968;
  assign n5819 = ~n10089 & n10123;
  assign n5820 = n4764 & n4966;
  assign n5821 = ~n5819 & ~n5820;
  assign n5822 = ~n5818 & ~n5820;
  assign n5823 = ~n5819 & n5822;
  assign n5824 = ~n5818 & n5821;
  assign n5825 = ~n5817 & n10214;
  assign n5826 = n5816 & ~n5825;
  assign n5827 = ~n5816 & n5825;
  assign n5828 = ~n1164 & ~n10090;
  assign n5829 = ~n1164 & ~n5825;
  assign n5830 = n5828 & ~n5829;
  assign n5831 = n5825 & n5828;
  assign n5832 = n5828 & ~n10215;
  assign n5833 = n1164 & n5825;
  assign n5834 = ~n5829 & ~n5833;
  assign n5835 = ~n10215 & n5834;
  assign n5836 = ~n5832 & ~n5835;
  assign n5837 = ~n5826 & ~n5827;
  assign n5838 = ~n10168 & ~n10216;
  assign n5839 = n10168 & n10216;
  assign n5840 = ~n10168 & ~n5838;
  assign n5841 = ~n10216 & ~n5838;
  assign n5842 = ~n5840 & ~n5841;
  assign n5843 = ~n5838 & ~n5839;
  assign n5844 = n5815 & ~n10217;
  assign n5845 = ~n5815 & n10217;
  assign n5846 = n5815 & ~n5844;
  assign n5847 = ~n10217 & ~n5844;
  assign n5848 = ~n5846 & ~n5847;
  assign n5849 = ~n5844 & ~n5845;
  assign n5850 = ~n5805 & ~n10218;
  assign n5851 = n5805 & n10218;
  assign n5852 = ~n5805 & n10218;
  assign n5853 = n5805 & ~n10218;
  assign n5854 = ~n5852 & ~n5853;
  assign n5855 = ~n5850 & ~n5851;
  assign n5856 = n5804 & ~n10219;
  assign n5857 = ~n5804 & n10219;
  assign n5858 = ~n5856 & ~n5857;
  assign n5859 = ~n5789 & n5858;
  assign n5860 = n5789 & ~n5858;
  assign n5861 = ~n5859 & ~n5860;
  assign n5862 = n5788 & n5861;
  assign n5863 = ~n5788 & ~n5861;
  assign n5864 = ~n5862 & ~n5863;
  assign n5865 = ~n5646 & n5864;
  assign n5866 = n5646 & ~n5864;
  assign n5867 = ~n5865 & ~n5866;
  assign n5868 = pi0  & ~pi22 ;
  assign n5869 = pi1  & ~n5868;
  assign n5870 = ~pi1  & n5868;
  assign n5871 = ~n5869 & ~n5870;
  assign n5872 = n73 & n5871;
  assign n5873 = ~n73 & ~n5871;
  assign n5874 = ~n73 & n5871;
  assign n5875 = n73 & ~n5871;
  assign n5876 = ~n5874 & ~n5875;
  assign n5877 = ~n5872 & ~n5873;
  assign n5878 = pi0  & ~n10220;
  assign n5879 = ~n226 & ~n538;
  assign n5880 = n4385 & n5879;
  assign n5881 = n758 & n1466;
  assign n5882 = n1662 & n3779;
  assign n5883 = n5881 & n5882;
  assign n5884 = n758 & n5879;
  assign n5885 = n1466 & n1662;
  assign n5886 = n3779 & n4385;
  assign n5887 = n5885 & n5886;
  assign n5888 = n5884 & n5887;
  assign n5889 = ~n226 & ~n300;
  assign n5890 = n546 & n5889;
  assign n5891 = n1662 & n4385;
  assign n5892 = n5881 & n5891;
  assign n5893 = n5890 & n5892;
  assign n5894 = ~n533 & ~n754;
  assign n5895 = ~n538 & ~n1661;
  assign n5896 = n5894 & n5895;
  assign n5897 = n758 & n5889;
  assign n5898 = n1466 & n4385;
  assign n5899 = n5897 & n5898;
  assign n5900 = n5896 & n5899;
  assign n5901 = n5880 & n5883;
  assign n5902 = n9995 & n10021;
  assign n5903 = n10221 & n5902;
  assign n5904 = n9636 & n5903;
  assign n5905 = n758 & ~n1661;
  assign n5906 = n9636 & n5905;
  assign n5907 = n9617 & n5906;
  assign n5908 = n9995 & n5907;
  assign n5909 = n10021 & n5908;
  assign n5910 = n4385 & n5909;
  assign n5911 = n1466 & n5910;
  assign n5912 = ~n538 & n5911;
  assign n5913 = ~n533 & n5912;
  assign n5914 = ~n226 & n5913;
  assign n5915 = ~n754 & n5914;
  assign n5916 = ~n300 & n5915;
  assign n5917 = n9617 & n5904;
  assign n5918 = n5766 & n10222;
  assign n5919 = ~n5766 & ~n10222;
  assign n5920 = ~n5918 & ~n5919;
  assign n5921 = ~n401 & ~n583;
  assign n5922 = n909 & n994;
  assign n5923 = n5921 & n5922;
  assign n5924 = ~n404 & n899;
  assign n5925 = n9762 & n5924;
  assign n5926 = n901 & n2075;
  assign n5927 = n899 & n994;
  assign n5928 = n5921 & n5927;
  assign n5929 = ~n404 & n909;
  assign n5930 = n9762 & n5929;
  assign n5931 = n5928 & n5930;
  assign n5932 = n5923 & n10223;
  assign n5933 = n9622 & n9630;
  assign n5934 = n10224 & n5933;
  assign n5935 = n9611 & n9636;
  assign n5936 = n9647 & n5935;
  assign n5937 = n9611 & n994;
  assign n5938 = n9762 & n5937;
  assign n5939 = n899 & n5938;
  assign n5940 = n9622 & n5939;
  assign n5941 = n909 & n5940;
  assign n5942 = n9636 & n5941;
  assign n5943 = n9647 & n5942;
  assign n5944 = n9630 & n5943;
  assign n5945 = n5921 & n5944;
  assign n5946 = ~n404 & n5945;
  assign n5947 = n5934 & n5936;
  assign n5948 = n5918 & n10225;
  assign n5949 = ~n5918 & ~n10225;
  assign n5950 = ~n5918 & n10225;
  assign n5951 = n5918 & ~n10225;
  assign n5952 = ~n5950 & ~n5951;
  assign n5953 = ~n5948 & ~n5949;
  assign n5954 = ~n5920 & n10226;
  assign n5955 = n10210 & ~n5920;
  assign n5956 = ~n5772 & ~n5776;
  assign n5957 = ~n10210 & n5920;
  assign n5958 = ~n10210 & n10222;
  assign n5959 = ~n5955 & ~n10227;
  assign n5960 = ~n5956 & n5959;
  assign n5961 = ~n5955 & ~n5960;
  assign n5962 = n5920 & ~n10226;
  assign n5963 = n5920 & n10225;
  assign n5964 = ~n5954 & ~n10228;
  assign n5965 = ~n5961 & n5964;
  assign n5966 = ~n5954 & ~n5965;
  assign n5967 = n9614 & n9636;
  assign n5968 = n9642 & n5967;
  assign n5969 = ~n295 & n9647;
  assign n5970 = ~n381 & n5969;
  assign n5971 = n453 & n9647;
  assign n5972 = ~n468 & ~n627;
  assign n5973 = n167 & n211;
  assign n5974 = ~n1015 & n10230;
  assign n5975 = n9620 & n5974;
  assign n5976 = n10229 & n5975;
  assign n5977 = n9642 & n10229;
  assign n5978 = n9636 & n5977;
  assign n5979 = n9614 & n5978;
  assign n5980 = n9620 & n5979;
  assign n5981 = ~n468 & n5980;
  assign n5982 = ~n627 & n5981;
  assign n5983 = ~n1015 & n5982;
  assign n5984 = n5968 & n5976;
  assign n5985 = ~n5948 & ~n10231;
  assign n5986 = n5948 & n10231;
  assign n5987 = ~n5985 & ~n5986;
  assign n5988 = n10226 & ~n5987;
  assign n5989 = ~n10226 & n5987;
  assign n5990 = ~n10226 & n10231;
  assign n5991 = ~n5988 & ~n10232;
  assign n5992 = ~n5966 & n5991;
  assign n5993 = n5966 & ~n5991;
  assign n5994 = ~n5992 & ~n5993;
  assign n5995 = n5878 & n5994;
  assign n5996 = pi0  & n10220;
  assign n5997 = ~n5987 & n5996;
  assign n5998 = n50 & ~n10220;
  assign n5999 = pi2  & n50;
  assign n6000 = ~n5920 & n10233;
  assign n6001 = ~pi0  & ~n5871;
  assign n6002 = n10226 & n6001;
  assign n6003 = ~n6000 & ~n6002;
  assign n6004 = ~n5997 & n6003;
  assign n6005 = ~n5878 & n6004;
  assign n6006 = ~n5994 & n6004;
  assign n6007 = ~n6005 & ~n6006;
  assign n6008 = ~n5995 & n6004;
  assign n6009 = n73 & ~n10234;
  assign n6010 = ~n73 & n10234;
  assign n6011 = ~n6009 & ~n6010;
  assign n6012 = n5867 & n6011;
  assign n6013 = n5639 & n10201;
  assign n6014 = ~n5645 & ~n6013;
  assign n6015 = n5961 & ~n5964;
  assign n6016 = ~n5965 & ~n6015;
  assign n6017 = n5878 & n6016;
  assign n6018 = n10226 & n5996;
  assign n6019 = n10210 & n10233;
  assign n6020 = ~n5920 & n6001;
  assign n6021 = ~n6019 & ~n6020;
  assign n6022 = ~n6018 & n6021;
  assign n6023 = ~n5878 & n6022;
  assign n6024 = ~n6016 & n6022;
  assign n6025 = ~n6023 & ~n6024;
  assign n6026 = ~n6017 & n6022;
  assign n6027 = n73 & ~n10235;
  assign n6028 = ~n73 & n10235;
  assign n6029 = ~n6027 & ~n6028;
  assign n6030 = n6014 & n6029;
  assign n6031 = n5632 & n10200;
  assign n6032 = ~n5638 & ~n6031;
  assign n6033 = n5956 & ~n5959;
  assign n6034 = ~n5960 & ~n6033;
  assign n6035 = n5878 & n6034;
  assign n6036 = ~n5920 & n5996;
  assign n6037 = ~n4870 & n10233;
  assign n6038 = n10210 & n6001;
  assign n6039 = ~n6037 & ~n6038;
  assign n6040 = ~n6036 & n6039;
  assign n6041 = ~n5878 & n6040;
  assign n6042 = ~n6034 & n6040;
  assign n6043 = ~n6041 & ~n6042;
  assign n6044 = ~n6035 & n6040;
  assign n6045 = n73 & ~n10236;
  assign n6046 = ~n73 & n10236;
  assign n6047 = ~n6045 & ~n6046;
  assign n6048 = n6032 & n6047;
  assign n6049 = ~n6032 & ~n6047;
  assign n6050 = n6032 & ~n6048;
  assign n6051 = n6047 & ~n6048;
  assign n6052 = ~n6050 & ~n6051;
  assign n6053 = ~n6048 & ~n6049;
  assign n6054 = n5628 & ~n5630;
  assign n6055 = ~n5631 & ~n6054;
  assign n6056 = n5619 & n10199;
  assign n6057 = ~n5627 & ~n6056;
  assign n6058 = n4876 & n5878;
  assign n6059 = ~n10084 & n6001;
  assign n6060 = ~n4870 & n5996;
  assign n6061 = ~n6059 & ~n6060;
  assign n6062 = ~n6058 & n6061;
  assign n6063 = n4731 & n10233;
  assign n6064 = ~n73 & ~n6063;
  assign n6065 = n6062 & ~n6064;
  assign n6066 = ~n73 & ~n6062;
  assign n6067 = n6062 & n6064;
  assign n6068 = n73 & ~n6062;
  assign n6069 = ~n6067 & ~n6068;
  assign n6070 = ~n6059 & ~n6063;
  assign n6071 = ~n6060 & ~n6063;
  assign n6072 = ~n6059 & n6071;
  assign n6073 = ~n6060 & n6070;
  assign n6074 = ~n6058 & n10239;
  assign n6075 = ~n73 & ~n6074;
  assign n6076 = n73 & n6074;
  assign n6077 = ~n6075 & ~n6076;
  assign n6078 = ~n6065 & ~n6066;
  assign n6079 = n6057 & ~n10238;
  assign n6080 = ~n6057 & n10238;
  assign n6081 = n5612 & n10196;
  assign n6082 = ~n5618 & ~n6081;
  assign n6083 = n5396 & n5878;
  assign n6084 = ~n10084 & n5996;
  assign n6085 = ~n10085 & n10233;
  assign n6086 = n4731 & n6001;
  assign n6087 = ~n6085 & ~n6086;
  assign n6088 = ~n6084 & n6087;
  assign n6089 = ~n6083 & n6088;
  assign n6090 = n73 & ~n6089;
  assign n6091 = ~n73 & n6089;
  assign n6092 = ~n6090 & ~n6091;
  assign n6093 = ~n6082 & n6092;
  assign n6094 = n5608 & ~n5610;
  assign n6095 = ~n5611 & ~n6094;
  assign n6096 = n5414 & n5878;
  assign n6097 = n4731 & n5996;
  assign n6098 = ~n10085 & n6001;
  assign n6099 = n4740 & n10233;
  assign n6100 = ~n6098 & ~n6099;
  assign n6101 = ~n6097 & ~n6099;
  assign n6102 = ~n6098 & n6101;
  assign n6103 = ~n6097 & n6100;
  assign n6104 = n73 & n10240;
  assign n6105 = ~n6096 & n10240;
  assign n6106 = n73 & n6105;
  assign n6107 = ~n6096 & n6104;
  assign n6108 = ~n73 & ~n10240;
  assign n6109 = ~n73 & n5878;
  assign n6110 = n5414 & n6109;
  assign n6111 = ~n6108 & ~n6110;
  assign n6112 = ~n6097 & ~n6098;
  assign n6113 = ~n6096 & n6112;
  assign n6114 = ~n73 & ~n6099;
  assign n6115 = n6113 & ~n6114;
  assign n6116 = ~n73 & ~n6113;
  assign n6117 = ~n6115 & ~n6116;
  assign n6118 = n6113 & n6114;
  assign n6119 = n73 & ~n6113;
  assign n6120 = ~n6118 & ~n6119;
  assign n6121 = ~n10241 & n6111;
  assign n6122 = ~n6095 & ~n10242;
  assign n6123 = n5597 & ~n5599;
  assign n6124 = ~n5600 & ~n6123;
  assign n6125 = n4740 & n5996;
  assign n6126 = ~n10087 & n10233;
  assign n6127 = ~n10086 & n6001;
  assign n6128 = ~n6126 & ~n6127;
  assign n6129 = ~n6125 & ~n6126;
  assign n6130 = ~n6127 & n6129;
  assign n6131 = ~n6125 & n6128;
  assign n6132 = ~n73 & ~n10243;
  assign n6133 = n5110 & n6109;
  assign n6134 = n5110 & n5878;
  assign n6135 = ~n6125 & ~n6127;
  assign n6136 = ~n6134 & n6135;
  assign n6137 = ~n6126 & n6136;
  assign n6138 = n10243 & ~n6134;
  assign n6139 = ~n73 & ~n10244;
  assign n6140 = ~n6132 & ~n6133;
  assign n6141 = n73 & n10243;
  assign n6142 = n73 & n6136;
  assign n6143 = n73 & n10244;
  assign n6144 = ~n6134 & n6141;
  assign n6145 = ~n73 & ~n6126;
  assign n6146 = n6136 & ~n6145;
  assign n6147 = ~n73 & ~n6136;
  assign n6148 = ~n6146 & ~n6147;
  assign n6149 = ~n10245 & ~n10246;
  assign n6150 = n6124 & n10247;
  assign n6151 = n5593 & ~n5595;
  assign n6152 = ~n5596 & ~n6151;
  assign n6153 = ~n5584 & n10194;
  assign n6154 = ~n10194 & ~n5592;
  assign n6155 = n5584 & ~n5592;
  assign n6156 = ~n6154 & ~n6155;
  assign n6157 = ~n5592 & ~n6153;
  assign n6158 = n9528 & ~n10188;
  assign n6159 = n10189 & n6158;
  assign n6160 = ~n10189 & ~n6158;
  assign n6161 = ~n10188 & ~n5569;
  assign n6162 = ~n10190 & ~n6161;
  assign n6163 = ~n6159 & ~n6160;
  assign n6164 = n9528 & n5550;
  assign n6165 = ~n5549 & n6164;
  assign n6166 = n5549 & ~n6164;
  assign n6167 = ~n5551 & ~n5554;
  assign n6168 = ~n10188 & ~n6167;
  assign n6169 = ~n6165 & ~n6166;
  assign n6170 = n10089 & n4957;
  assign n6171 = n5878 & ~n6170;
  assign n6172 = n10089 & n10090;
  assign n6173 = n5996 & ~n6172;
  assign n6174 = ~n10090 & n6001;
  assign n6175 = ~n9527 & ~n4775;
  assign n6176 = ~n73 & ~n6175;
  assign n6177 = ~n6174 & n6176;
  assign n6178 = ~n6173 & n6177;
  assign n6179 = pi0  & ~n4775;
  assign n6180 = n10115 & n6109;
  assign n6181 = ~n10089 & n5996;
  assign n6182 = ~n4775 & n10233;
  assign n6183 = ~n6174 & ~n6182;
  assign n6184 = ~n6181 & n6183;
  assign n6185 = ~n73 & ~n6184;
  assign n6186 = ~n4957 & n6109;
  assign n6187 = ~n10090 & n5996;
  assign n6188 = ~n4775 & n6001;
  assign n6189 = ~n73 & ~n6188;
  assign n6190 = ~n6187 & n6189;
  assign n6191 = ~n6186 & n6190;
  assign n6192 = ~n6185 & n6191;
  assign n6193 = ~n6180 & n6192;
  assign n6194 = ~n6179 & n6193;
  assign n6195 = ~n50 & ~n4775;
  assign n6196 = ~n73 & ~n6179;
  assign n6197 = ~n6188 & n6196;
  assign n6198 = ~n73 & ~n6195;
  assign n6199 = ~n6187 & n10252;
  assign n6200 = ~n6186 & n6199;
  assign n6201 = ~n6185 & n6200;
  assign n6202 = ~n6180 & n6201;
  assign n6203 = ~n6180 & n6200;
  assign n6204 = ~n6185 & n6203;
  assign n6205 = ~n6171 & n6178;
  assign n6206 = ~n5550 & ~n10251;
  assign n6207 = ~n10118 & n5878;
  assign n6208 = n4764 & n5996;
  assign n6209 = ~n10089 & n6001;
  assign n6210 = ~n10090 & n10233;
  assign n6211 = ~n6209 & ~n6210;
  assign n6212 = ~n6208 & ~n6210;
  assign n6213 = ~n6209 & n6212;
  assign n6214 = ~n6208 & n6211;
  assign n6215 = ~n6207 & n10253;
  assign n6216 = ~n73 & n6215;
  assign n6217 = n73 & ~n6215;
  assign n6218 = n73 & n6215;
  assign n6219 = ~n73 & ~n6215;
  assign n6220 = ~n6218 & ~n6219;
  assign n6221 = ~n6216 & ~n6217;
  assign n6222 = ~n6206 & ~n6219;
  assign n6223 = ~n6218 & n6222;
  assign n6224 = ~n6206 & n10254;
  assign n6225 = n10250 & n10255;
  assign n6226 = ~n10250 & ~n10255;
  assign n6227 = n4761 & n5996;
  assign n6228 = ~n10089 & n10233;
  assign n6229 = n4764 & n6001;
  assign n6230 = ~n6228 & ~n6229;
  assign n6231 = ~n6227 & ~n6229;
  assign n6232 = ~n6228 & n6231;
  assign n6233 = ~n6227 & n6230;
  assign n6234 = ~n73 & ~n10256;
  assign n6235 = ~n10104 & n6109;
  assign n6236 = ~n10104 & n5878;
  assign n6237 = n10256 & ~n6236;
  assign n6238 = ~n73 & ~n6237;
  assign n6239 = ~n6234 & ~n6235;
  assign n6240 = n73 & n10256;
  assign n6241 = n73 & n6237;
  assign n6242 = ~n6236 & n6240;
  assign n6243 = ~n10257 & ~n10258;
  assign n6244 = ~n6226 & ~n6235;
  assign n6245 = ~n10258 & n6244;
  assign n6246 = ~n6234 & n6245;
  assign n6247 = ~n6226 & n6243;
  assign n6248 = ~n6225 & ~n10259;
  assign n6249 = ~n10249 & n6248;
  assign n6250 = n10249 & ~n6248;
  assign n6251 = n5052 & n5878;
  assign n6252 = ~n10088 & n5996;
  assign n6253 = n4764 & n10233;
  assign n6254 = n4761 & n6001;
  assign n6255 = ~n6253 & ~n6254;
  assign n6256 = ~n6252 & n6255;
  assign n6257 = ~n6251 & n6256;
  assign n6258 = ~n73 & ~n6257;
  assign n6259 = ~n6257 & ~n6258;
  assign n6260 = n73 & ~n6257;
  assign n6261 = ~n73 & ~n6258;
  assign n6262 = ~n73 & n6257;
  assign n6263 = ~n10260 & ~n10261;
  assign n6264 = ~n6250 & n6263;
  assign n6265 = n6248 & n6263;
  assign n6266 = ~n10190 & ~n6265;
  assign n6267 = ~n6161 & n6266;
  assign n6268 = n10249 & ~n6265;
  assign n6269 = ~n6248 & ~n6263;
  assign n6270 = ~n10262 & ~n6269;
  assign n6271 = ~n6249 & ~n6264;
  assign n6272 = n10248 & n10263;
  assign n6273 = ~n10248 & ~n10263;
  assign n6274 = n5164 & n5878;
  assign n6275 = ~n10087 & n5996;
  assign n6276 = n4761 & n10233;
  assign n6277 = ~n10088 & n6001;
  assign n6278 = ~n6276 & ~n6277;
  assign n6279 = ~n6275 & n6278;
  assign n6280 = n73 & n6279;
  assign n6281 = ~n6274 & n6279;
  assign n6282 = n73 & n6281;
  assign n6283 = ~n6274 & n6280;
  assign n6284 = ~n73 & ~n6279;
  assign n6285 = n5164 & n6109;
  assign n6286 = ~n6284 & ~n6285;
  assign n6287 = n73 & ~n6281;
  assign n6288 = ~n73 & n6281;
  assign n6289 = ~n6287 & ~n6288;
  assign n6290 = ~n10264 & n6286;
  assign n6291 = ~n6273 & n10265;
  assign n6292 = ~n6272 & ~n6285;
  assign n6293 = ~n10264 & n6292;
  assign n6294 = ~n6284 & n6293;
  assign n6295 = ~n6272 & ~n10265;
  assign n6296 = ~n6273 & ~n10266;
  assign n6297 = ~n6272 & ~n6291;
  assign n6298 = n6152 & ~n10267;
  assign n6299 = n5145 & n5878;
  assign n6300 = ~n10086 & n5996;
  assign n6301 = ~n10088 & n10233;
  assign n6302 = ~n10087 & n6001;
  assign n6303 = ~n6301 & ~n6302;
  assign n6304 = ~n6300 & n6303;
  assign n6305 = ~n6299 & n6304;
  assign n6306 = ~n73 & ~n6305;
  assign n6307 = ~n6305 & ~n6306;
  assign n6308 = n73 & ~n6305;
  assign n6309 = ~n73 & ~n6306;
  assign n6310 = ~n73 & n6305;
  assign n6311 = ~n10268 & ~n10269;
  assign n6312 = ~n6298 & n6311;
  assign n6313 = ~n6152 & n10267;
  assign n6314 = ~n6124 & ~n10247;
  assign n6315 = ~n6313 & ~n6314;
  assign n6316 = ~n6312 & n6315;
  assign n6317 = n10267 & n6311;
  assign n6318 = ~n5596 & ~n6317;
  assign n6319 = ~n6151 & n6318;
  assign n6320 = n6152 & ~n6317;
  assign n6321 = ~n10267 & ~n6311;
  assign n6322 = ~n10270 & ~n6321;
  assign n6323 = ~n6124 & n6322;
  assign n6324 = ~n6133 & ~n6323;
  assign n6325 = ~n10246 & n6324;
  assign n6326 = ~n6132 & n6325;
  assign n6327 = n10247 & ~n6323;
  assign n6328 = n6124 & ~n6322;
  assign n6329 = ~n10271 & ~n6328;
  assign n6330 = ~n6150 & ~n6316;
  assign n6331 = n5601 & n10195;
  assign n6332 = ~n5601 & ~n5607;
  assign n6333 = ~n10195 & ~n5607;
  assign n6334 = ~n6332 & ~n6333;
  assign n6335 = ~n5607 & ~n6331;
  assign n6336 = n10272 & n10273;
  assign n6337 = ~n10085 & n5996;
  assign n6338 = ~n10086 & n10233;
  assign n6339 = n4740 & n6001;
  assign n6340 = ~n6338 & ~n6339;
  assign n6341 = ~n6337 & n6340;
  assign n6342 = ~n73 & ~n6341;
  assign n6343 = n5368 & n6109;
  assign n6344 = n5368 & n5878;
  assign n6345 = n6341 & ~n6344;
  assign n6346 = ~n73 & ~n6345;
  assign n6347 = ~n6342 & ~n6343;
  assign n6348 = n73 & n6341;
  assign n6349 = n73 & n6345;
  assign n6350 = ~n6344 & n6348;
  assign n6351 = ~n10274 & ~n10275;
  assign n6352 = ~n6336 & ~n6343;
  assign n6353 = ~n10275 & n6352;
  assign n6354 = ~n6342 & n6353;
  assign n6355 = ~n6336 & n6351;
  assign n6356 = ~n10272 & ~n10273;
  assign n6357 = n6095 & n10242;
  assign n6358 = ~n6356 & ~n6357;
  assign n6359 = ~n10276 & n6358;
  assign n6360 = ~n10276 & ~n6356;
  assign n6361 = ~n10242 & n6360;
  assign n6362 = n10242 & ~n6360;
  assign n6363 = ~n6095 & ~n6362;
  assign n6364 = ~n6361 & ~n6363;
  assign n6365 = ~n6095 & n6360;
  assign n6366 = ~n6110 & ~n6365;
  assign n6367 = ~n10241 & n6366;
  assign n6368 = ~n6108 & n6367;
  assign n6369 = n10242 & ~n6365;
  assign n6370 = n6095 & ~n6360;
  assign n6371 = ~n10278 & ~n6370;
  assign n6372 = ~n6122 & ~n6359;
  assign n6373 = ~n6093 & n10277;
  assign n6374 = n6082 & ~n6092;
  assign n6375 = n6082 & n10277;
  assign n6376 = n6092 & ~n6375;
  assign n6377 = ~n6082 & ~n10277;
  assign n6378 = ~n6376 & ~n6377;
  assign n6379 = ~n6373 & ~n6374;
  assign n6380 = ~n6080 & ~n6377;
  assign n6381 = ~n6376 & n6380;
  assign n6382 = ~n6080 & n10279;
  assign n6383 = ~n6057 & ~n10279;
  assign n6384 = ~n10238 & ~n6383;
  assign n6385 = n6057 & n10279;
  assign n6386 = ~n6384 & ~n6385;
  assign n6387 = ~n6079 & ~n10280;
  assign n6388 = ~n6055 & n10281;
  assign n6389 = n6055 & ~n10281;
  assign n6390 = n5778 & n5878;
  assign n6391 = n10210 & n5996;
  assign n6392 = ~n10084 & n10233;
  assign n6393 = ~n4870 & n6001;
  assign n6394 = ~n6392 & ~n6393;
  assign n6395 = ~n6391 & n6394;
  assign n6396 = ~n6390 & n6395;
  assign n6397 = ~n73 & ~n6396;
  assign n6398 = ~n6396 & ~n6397;
  assign n6399 = n73 & ~n6396;
  assign n6400 = ~n73 & ~n6397;
  assign n6401 = ~n73 & n6396;
  assign n6402 = ~n10282 & ~n10283;
  assign n6403 = ~n6389 & n6402;
  assign n6404 = n10281 & n6402;
  assign n6405 = ~n5631 & ~n6404;
  assign n6406 = ~n6054 & n6405;
  assign n6407 = n6055 & ~n6404;
  assign n6408 = ~n10281 & ~n6402;
  assign n6409 = ~n10284 & ~n6408;
  assign n6410 = ~n6388 & ~n6403;
  assign n6411 = ~n10237 & ~n10285;
  assign n6412 = ~n6048 & ~n6411;
  assign n6413 = ~n6014 & ~n6029;
  assign n6414 = n6014 & ~n6030;
  assign n6415 = n6029 & ~n6030;
  assign n6416 = ~n6414 & ~n6415;
  assign n6417 = ~n6030 & ~n6413;
  assign n6418 = ~n6412 & ~n10286;
  assign n6419 = ~n6030 & ~n6418;
  assign n6420 = ~n5867 & ~n6011;
  assign n6421 = ~n6012 & ~n6420;
  assign n6422 = ~n6419 & n6421;
  assign n6423 = ~n6012 & ~n6422;
  assign n6424 = ~n5988 & ~n5992;
  assign n6425 = ~n554 & ~n898;
  assign n6426 = ~n260 & ~n9570;
  assign n6427 = ~n9570 & ~n554;
  assign n6428 = ~n260 & ~n898;
  assign n6429 = n6427 & n6428;
  assign n6430 = n6425 & n6426;
  assign n6431 = ~n300 & ~n351;
  assign n6432 = n203 & n3893;
  assign n6433 = n6431 & n6432;
  assign n6434 = n203 & n6431;
  assign n6435 = ~n9570 & n6434;
  assign n6436 = ~n554 & n6435;
  assign n6437 = ~n604 & n6436;
  assign n6438 = ~n898 & n6437;
  assign n6439 = ~n470 & n6438;
  assign n6440 = ~n260 & n6439;
  assign n6441 = ~n9570 & ~n604;
  assign n6442 = ~n260 & ~n470;
  assign n6443 = n6441 & n6442;
  assign n6444 = n6425 & n6431;
  assign n6445 = n203 & n6444;
  assign n6446 = n6443 & n6445;
  assign n6447 = n10287 & n6433;
  assign n6448 = ~n324 & ~n624;
  assign n6449 = n1191 & n6448;
  assign n6450 = ~n175 & ~n663;
  assign n6451 = n4825 & n6450;
  assign n6452 = n6449 & n6451;
  assign n6453 = ~n294 & ~n1070;
  assign n6454 = ~n398 & n6453;
  assign n6455 = n9545 & n6454;
  assign n6456 = ~n398 & ~n624;
  assign n6457 = n482 & n6456;
  assign n6458 = n4385 & n4825;
  assign n6459 = n6457 & n6458;
  assign n6460 = ~n1070 & n6450;
  assign n6461 = n9545 & n6460;
  assign n6462 = n6459 & n6461;
  assign n6463 = ~n175 & ~n479;
  assign n6464 = ~n624 & ~n730;
  assign n6465 = n6463 & n6464;
  assign n6466 = ~n324 & ~n398;
  assign n6467 = n4385 & n6466;
  assign n6468 = n6465 & n6467;
  assign n6469 = ~n663 & ~n1070;
  assign n6470 = ~n352 & n6469;
  assign n6471 = n9545 & n6470;
  assign n6472 = n6468 & n6471;
  assign n6473 = n6452 & n6455;
  assign n6474 = n10077 & n10289;
  assign n6475 = n10288 & n6474;
  assign n6476 = n9545 & ~n1070;
  assign n6477 = n10077 & n6476;
  assign n6478 = n9761 & n6477;
  assign n6479 = n10288 & n6478;
  assign n6480 = n4385 & n6479;
  assign n6481 = ~n624 & n6480;
  assign n6482 = ~n663 & n6481;
  assign n6483 = ~n324 & n6482;
  assign n6484 = ~n175 & n6483;
  assign n6485 = ~n352 & n6484;
  assign n6486 = ~n479 & n6485;
  assign n6487 = ~n398 & n6486;
  assign n6488 = ~n730 & n6487;
  assign n6489 = n9761 & n6475;
  assign n6490 = ~n5986 & ~n10290;
  assign n6491 = n5986 & ~n10290;
  assign n6492 = ~n10290 & ~n6491;
  assign n6493 = ~n5987 & n6492;
  assign n6494 = ~n5987 & n6490;
  assign n6495 = n5987 & ~n6492;
  assign n6496 = n5987 & n10290;
  assign n6497 = ~n10291 & ~n10292;
  assign n6498 = ~n6424 & n6497;
  assign n6499 = n6424 & ~n6497;
  assign n6500 = ~n6498 & ~n6499;
  assign n6501 = n5878 & n6500;
  assign n6502 = n5996 & n6492;
  assign n6503 = n5996 & n6490;
  assign n6504 = n10226 & n10233;
  assign n6505 = ~n5987 & n6001;
  assign n6506 = ~n6504 & ~n6505;
  assign n6507 = ~n10293 & n6506;
  assign n6508 = ~n6501 & n6507;
  assign n6509 = ~n73 & ~n6508;
  assign n6510 = ~n6508 & ~n6509;
  assign n6511 = n73 & ~n6508;
  assign n6512 = ~n73 & ~n6509;
  assign n6513 = ~n73 & n6508;
  assign n6514 = ~n10294 & ~n10295;
  assign n6515 = ~n5862 & ~n5865;
  assign n6516 = ~n5856 & ~n5859;
  assign n6517 = n5108 & n5396;
  assign n6518 = ~n10084 & n5112;
  assign n6519 = ~n10085 & n10130;
  assign n6520 = n4731 & n5120;
  assign n6521 = ~n6519 & ~n6520;
  assign n6522 = ~n6518 & n6521;
  assign n6523 = ~n6517 & n6522;
  assign n6524 = ~n1703 & ~n6523;
  assign n6525 = ~n6523 & ~n6524;
  assign n6526 = n1703 & ~n6523;
  assign n6527 = ~n1703 & ~n6524;
  assign n6528 = ~n1703 & n6523;
  assign n6529 = ~n10296 & ~n10297;
  assign n6530 = ~n5844 & ~n5850;
  assign n6531 = ~n1164 & n10089;
  assign n6532 = n4958 & n5052;
  assign n6533 = ~n10088 & n4968;
  assign n6534 = n4764 & n10123;
  assign n6535 = n4761 & n4966;
  assign n6536 = ~n6534 & ~n6535;
  assign n6537 = ~n6533 & n6536;
  assign n6538 = ~n6532 & n6537;
  assign n6539 = n6531 & ~n6538;
  assign n6540 = ~n6531 & n6538;
  assign n6541 = ~n6539 & ~n6540;
  assign n6542 = ~n10215 & ~n5838;
  assign n6543 = n6541 & ~n6542;
  assign n6544 = ~n6541 & n6542;
  assign n6545 = ~n6543 & ~n6544;
  assign n6546 = n4913 & n5110;
  assign n6547 = n4740 & n4920;
  assign n6548 = ~n10086 & n4933;
  assign n6549 = ~n10087 & n10106;
  assign n6550 = ~n6548 & ~n6549;
  assign n6551 = ~n6547 & ~n6549;
  assign n6552 = ~n6548 & n6551;
  assign n6553 = ~n6547 & n6550;
  assign n6554 = ~n4913 & n10298;
  assign n6555 = ~n5110 & n10298;
  assign n6556 = ~n6554 & ~n6555;
  assign n6557 = ~n6546 & n10298;
  assign n6558 = ~n9626 & ~n10299;
  assign n6559 = n9626 & n10299;
  assign n6560 = ~n6558 & ~n6559;
  assign n6561 = n6545 & n6560;
  assign n6562 = ~n6545 & ~n6560;
  assign n6563 = n6545 & ~n6561;
  assign n6564 = n6560 & ~n6561;
  assign n6565 = ~n6563 & ~n6564;
  assign n6566 = ~n6561 & ~n6562;
  assign n6567 = ~n6530 & ~n10300;
  assign n6568 = n6530 & n10300;
  assign n6569 = ~n6530 & ~n6567;
  assign n6570 = ~n10300 & ~n6567;
  assign n6571 = ~n6569 & ~n6570;
  assign n6572 = ~n6567 & ~n6568;
  assign n6573 = ~n6529 & ~n10301;
  assign n6574 = n6529 & n10301;
  assign n6575 = ~n6529 & ~n6573;
  assign n6576 = ~n10301 & ~n6573;
  assign n6577 = ~n6575 & ~n6576;
  assign n6578 = ~n6573 & ~n6574;
  assign n6579 = n6516 & n10302;
  assign n6580 = ~n6516 & ~n10302;
  assign n6581 = ~n6579 & ~n6580;
  assign n6582 = n90 & n6034;
  assign n6583 = n4878 & ~n5920;
  assign n6584 = ~n4870 & n10100;
  assign n6585 = n4886 & n10210;
  assign n6586 = ~n6584 & ~n6585;
  assign n6587 = ~n6583 & n6586;
  assign n6588 = ~n90 & n6587;
  assign n6589 = ~n6034 & n6587;
  assign n6590 = ~n6588 & ~n6589;
  assign n6591 = ~n6582 & n6587;
  assign n6592 = ~n9528 & ~n10303;
  assign n6593 = n9528 & n10303;
  assign n6594 = ~n6592 & ~n6593;
  assign n6595 = n6581 & n6594;
  assign n6596 = ~n6581 & ~n6594;
  assign n6597 = n6581 & ~n6595;
  assign n6598 = n6594 & ~n6595;
  assign n6599 = ~n6597 & ~n6598;
  assign n6600 = ~n6595 & ~n6596;
  assign n6601 = ~n6515 & ~n10304;
  assign n6602 = n6515 & n10304;
  assign n6603 = ~n6515 & ~n6601;
  assign n6604 = ~n10304 & ~n6601;
  assign n6605 = ~n6603 & ~n6604;
  assign n6606 = ~n6601 & ~n6602;
  assign n6607 = ~n6514 & ~n10305;
  assign n6608 = n6514 & n10305;
  assign n6609 = ~n6514 & ~n6607;
  assign n6610 = ~n10305 & ~n6607;
  assign n6611 = ~n6609 & ~n6610;
  assign n6612 = ~n6607 & ~n6608;
  assign n6613 = n6423 & n10306;
  assign n6614 = ~n6423 & ~n10306;
  assign n6615 = ~n6613 & ~n6614;
  assign n6616 = n9742 & n9828;
  assign n6617 = n9742 & n10207;
  assign n6618 = n9828 & n6617;
  assign n6619 = n10207 & n6616;
  assign n6620 = ~n623 & ~n871;
  assign n6621 = ~n381 & ~n623;
  assign n6622 = ~n871 & n6621;
  assign n6623 = ~n381 & ~n871;
  assign n6624 = ~n623 & n6623;
  assign n6625 = ~n381 & n6620;
  assign n6626 = n773 & n6431;
  assign n6627 = n10308 & n6626;
  assign n6628 = n9664 & n6627;
  assign n6629 = n10307 & n6628;
  assign n6630 = n9593 & n6629;
  assign n6631 = n9742 & n6431;
  assign n6632 = n773 & n6631;
  assign n6633 = n9828 & n6632;
  assign n6634 = n10014 & n6633;
  assign n6635 = n9664 & n6634;
  assign n6636 = n9593 & n6635;
  assign n6637 = n10207 & n6636;
  assign n6638 = ~n871 & n6637;
  assign n6639 = ~n381 & n6638;
  assign n6640 = ~n623 & n6639;
  assign n6641 = n10014 & n6630;
  assign n6642 = ~n6615 & n10309;
  assign n6643 = n6615 & ~n10309;
  assign n6644 = ~n6642 & ~n6643;
  assign n6645 = n6419 & ~n6421;
  assign n6646 = ~n6422 & ~n6645;
  assign n6647 = ~n9555 & ~n730;
  assign n6648 = ~n9551 & ~n1015;
  assign n6649 = ~n9551 & ~n730;
  assign n6650 = ~n9555 & ~n1015;
  assign n6651 = n6649 & n6650;
  assign n6652 = n6647 & n6648;
  assign n6653 = ~n249 & ~n9551;
  assign n6654 = ~n9555 & ~n432;
  assign n6655 = ~n249 & n6654;
  assign n6656 = ~n9551 & n6655;
  assign n6657 = n6653 & n6654;
  assign n6658 = ~n1015 & n10311;
  assign n6659 = ~n730 & n6658;
  assign n6660 = ~n730 & ~n1015;
  assign n6661 = n10311 & n6660;
  assign n6662 = n4347 & n10310;
  assign n6663 = ~n215 & ~n624;
  assign n6664 = ~n175 & ~n627;
  assign n6665 = n6663 & n6664;
  assign n6666 = ~n9561 & ~n480;
  assign n6667 = n244 & n6666;
  assign n6668 = n3844 & n6431;
  assign n6669 = n6667 & n6668;
  assign n6670 = ~n175 & ~n480;
  assign n6671 = ~n215 & ~n9561;
  assign n6672 = n6670 & n6671;
  assign n6673 = ~n624 & ~n627;
  assign n6674 = n244 & n6673;
  assign n6675 = n6668 & n6674;
  assign n6676 = n6672 & n6675;
  assign n6677 = ~n215 & ~n627;
  assign n6678 = ~n9561 & ~n624;
  assign n6679 = n6677 & n6678;
  assign n6680 = ~n243 & ~n480;
  assign n6681 = ~n175 & ~n241;
  assign n6682 = n6680 & n6681;
  assign n6683 = n6668 & n6682;
  assign n6684 = n6679 & n6683;
  assign n6685 = n6665 & n6669;
  assign n6686 = n10312 & n6668;
  assign n6687 = ~n624 & n6686;
  assign n6688 = ~n9561 & n6687;
  assign n6689 = ~n215 & n6688;
  assign n6690 = ~n627 & n6689;
  assign n6691 = ~n175 & n6690;
  assign n6692 = ~n241 & n6691;
  assign n6693 = ~n243 & n6692;
  assign n6694 = ~n480 & n6693;
  assign n6695 = n10312 & n10313;
  assign n6696 = ~n226 & ~n479;
  assign n6697 = ~n581 & ~n990;
  assign n6698 = ~n226 & ~n990;
  assign n6699 = ~n479 & ~n581;
  assign n6700 = n6698 & n6699;
  assign n6701 = n6696 & n6697;
  assign n6702 = ~n581 & n10314;
  assign n6703 = ~n990 & n6702;
  assign n6704 = ~n226 & n6703;
  assign n6705 = ~n479 & n6704;
  assign n6706 = n10314 & n10315;
  assign n6707 = ~n219 & ~n620;
  assign n6708 = n826 & n6707;
  assign n6709 = n9557 & n6708;
  assign n6710 = n826 & n10205;
  assign n6711 = n9557 & n6710;
  assign n6712 = ~n219 & n6711;
  assign n6713 = ~n620 & n6712;
  assign n6714 = n10205 & n6709;
  assign n6715 = n1223 & n4641;
  assign n6716 = ~n536 & ~n720;
  assign n6717 = ~n258 & ~n265;
  assign n6718 = n6716 & n6717;
  assign n6719 = n6715 & n6718;
  assign n6720 = ~n312 & ~n554;
  assign n6721 = ~n296 & n6720;
  assign n6722 = n10207 & n6721;
  assign n6723 = ~n265 & n10207;
  assign n6724 = ~n296 & ~n554;
  assign n6725 = ~n312 & ~n720;
  assign n6726 = ~n554 & ~n720;
  assign n6727 = ~n296 & ~n312;
  assign n6728 = n6726 & n6727;
  assign n6729 = ~n296 & ~n720;
  assign n6730 = n6720 & n6729;
  assign n6731 = n6724 & n6725;
  assign n6732 = n5671 & n6715;
  assign n6733 = n10318 & n6732;
  assign n6734 = n6723 & n6733;
  assign n6735 = n6719 & n6722;
  assign n6736 = n9567 & n10319;
  assign n6737 = n10317 & n6736;
  assign n6738 = n10316 & n6715;
  assign n6739 = n10207 & n6738;
  assign n6740 = n10317 & n6739;
  assign n6741 = n9567 & n6740;
  assign n6742 = ~n296 & n6741;
  assign n6743 = ~n312 & n6742;
  assign n6744 = ~n554 & n6743;
  assign n6745 = ~n265 & n6744;
  assign n6746 = ~n258 & n6745;
  assign n6747 = ~n720 & n6746;
  assign n6748 = ~n536 & n6747;
  assign n6749 = n10316 & n6737;
  assign n6750 = ~n6646 & n10320;
  assign n6751 = n6646 & ~n10320;
  assign n6752 = n6412 & ~n6415;
  assign n6753 = ~n6414 & n6752;
  assign n6754 = n6412 & n10286;
  assign n6755 = ~n6418 & ~n10321;
  assign n6756 = ~n480 & ~n871;
  assign n6757 = n685 & n6756;
  assign n6758 = n4127 & n6757;
  assign n6759 = ~n9553 & ~n470;
  assign n6760 = ~n294 & ~n470;
  assign n6761 = ~n9553 & n6760;
  assign n6762 = ~n294 & n6759;
  assign n6763 = n10027 & n10322;
  assign n6764 = n4127 & n6759;
  assign n6765 = n685 & n6764;
  assign n6766 = ~n294 & ~n480;
  assign n6767 = ~n871 & n6766;
  assign n6768 = n10027 & n6767;
  assign n6769 = n6765 & n6768;
  assign n6770 = ~n241 & ~n480;
  assign n6771 = ~n470 & ~n871;
  assign n6772 = n6770 & n6771;
  assign n6773 = n685 & n6772;
  assign n6774 = ~n9553 & ~n515;
  assign n6775 = ~n294 & n6774;
  assign n6776 = n10027 & n6775;
  assign n6777 = n6773 & n6776;
  assign n6778 = n6758 & n6763;
  assign n6779 = n685 & n10027;
  assign n6780 = n9755 & n6779;
  assign n6781 = ~n241 & n6780;
  assign n6782 = ~n871 & n6781;
  assign n6783 = ~n515 & n6782;
  assign n6784 = ~n294 & n6783;
  assign n6785 = ~n470 & n6784;
  assign n6786 = ~n9553 & n6785;
  assign n6787 = ~n480 & n6786;
  assign n6788 = n9755 & n10323;
  assign n6789 = ~n195 & ~n9550;
  assign n6790 = n9604 & n6789;
  assign n6791 = n9604 & n10324;
  assign n6792 = ~n9550 & n6791;
  assign n6793 = ~n195 & n6792;
  assign n6794 = n10324 & n6790;
  assign n6795 = ~n513 & ~n552;
  assign n6796 = ~n258 & ~n284;
  assign n6797 = ~n284 & ~n384;
  assign n6798 = ~n258 & n6797;
  assign n6799 = ~n384 & n6796;
  assign n6800 = ~n258 & ~n513;
  assign n6801 = ~n552 & n6800;
  assign n6802 = ~n284 & n6801;
  assign n6803 = ~n384 & n6802;
  assign n6804 = ~n258 & ~n384;
  assign n6805 = ~n284 & ~n513;
  assign n6806 = ~n552 & n6805;
  assign n6807 = n6804 & n6806;
  assign n6808 = n6795 & n10326;
  assign n6809 = ~n397 & ~n604;
  assign n6810 = n706 & n6809;
  assign n6811 = n773 & n3945;
  assign n6812 = n5727 & n6811;
  assign n6813 = n773 & n6809;
  assign n6814 = n706 & n3945;
  assign n6815 = n5727 & n6814;
  assign n6816 = n6813 & n6815;
  assign n6817 = n3945 & n6809;
  assign n6818 = n706 & n773;
  assign n6819 = n5727 & n6818;
  assign n6820 = n6817 & n6819;
  assign n6821 = ~n431 & ~n604;
  assign n6822 = n5727 & n6821;
  assign n6823 = ~n397 & ~n405;
  assign n6824 = n706 & n6823;
  assign n6825 = n773 & n6824;
  assign n6826 = n6822 & n6825;
  assign n6827 = n6810 & n6812;
  assign n6828 = n773 & n10327;
  assign n6829 = ~n405 & n6828;
  assign n6830 = ~n386 & n6829;
  assign n6831 = ~n199 & n6830;
  assign n6832 = ~n604 & n6831;
  assign n6833 = ~n394 & n6832;
  assign n6834 = ~n431 & n6833;
  assign n6835 = ~n397 & n6834;
  assign n6836 = ~n536 & n6835;
  assign n6837 = n10327 & n10328;
  assign n6838 = ~n230 & ~n380;
  assign n6839 = ~n573 & n6838;
  assign n6840 = n1432 & n1888;
  assign n6841 = n1481 & n5670;
  assign n6842 = n6840 & n6841;
  assign n6843 = ~n415 & ~n573;
  assign n6844 = ~n380 & n6843;
  assign n6845 = ~n230 & ~n533;
  assign n6846 = n1432 & n6845;
  assign n6847 = n6841 & n6846;
  assign n6848 = n6844 & n6847;
  assign n6849 = ~n230 & n5670;
  assign n6850 = ~n533 & ~n573;
  assign n6851 = n1481 & n6850;
  assign n6852 = ~n380 & ~n415;
  assign n6853 = n1432 & n6852;
  assign n6854 = n6851 & n6853;
  assign n6855 = n6849 & n6854;
  assign n6856 = n6839 & n6842;
  assign n6857 = n10058 & n10330;
  assign n6858 = n10329 & n6857;
  assign n6859 = n10058 & n10325;
  assign n6860 = n10329 & n6859;
  assign n6861 = n1432 & n6860;
  assign n6862 = ~n415 & n6861;
  assign n6863 = ~n573 & n6862;
  assign n6864 = ~n897 & n6863;
  assign n6865 = ~n995 & n6864;
  assign n6866 = ~n380 & n6865;
  assign n6867 = ~n533 & n6866;
  assign n6868 = ~n1108 & n6867;
  assign n6869 = ~n230 & n6868;
  assign n6870 = ~n1037 & n6869;
  assign n6871 = n10325 & n6858;
  assign n6872 = ~n6755 & n10331;
  assign n6873 = n6755 & ~n10331;
  assign n6874 = n10237 & n10285;
  assign n6875 = ~n383 & ~n415;
  assign n6876 = n10075 & n6875;
  assign n6877 = n9602 & n10075;
  assign n6878 = ~n415 & n6877;
  assign n6879 = ~n383 & n6878;
  assign n6880 = n9602 & n6875;
  assign n6881 = n10075 & n6880;
  assign n6882 = n9602 & n6876;
  assign n6883 = ~n402 & ~n781;
  assign n6884 = n899 & n6883;
  assign n6885 = ~n190 & ~n402;
  assign n6886 = ~n264 & ~n781;
  assign n6887 = n6885 & n6886;
  assign n6888 = n899 & n6887;
  assign n6889 = n2547 & n6884;
  assign n6890 = n10009 & n10333;
  assign n6891 = n899 & n10009;
  assign n6892 = n10017 & n6891;
  assign n6893 = ~n402 & n6892;
  assign n6894 = ~n264 & n6893;
  assign n6895 = ~n190 & n6894;
  assign n6896 = ~n781 & n6895;
  assign n6897 = n10017 & n6890;
  assign n6898 = n628 & n4397;
  assign n6899 = n4432 & n6450;
  assign n6900 = n628 & n4432;
  assign n6901 = n4397 & n6450;
  assign n6902 = n6900 & n6901;
  assign n6903 = n6898 & n6899;
  assign n6904 = ~n386 & ~n582;
  assign n6905 = ~n328 & n6904;
  assign n6906 = n993 & n1192;
  assign n6907 = n6905 & n6906;
  assign n6908 = n4397 & n4432;
  assign n6909 = n993 & n4397;
  assign n6910 = n4432 & n6909;
  assign n6911 = n1192 & n6910;
  assign n6912 = n6906 & n6908;
  assign n6913 = ~n582 & ~n663;
  assign n6914 = ~n626 & n6913;
  assign n6915 = ~n328 & ~n386;
  assign n6916 = n6664 & n6915;
  assign n6917 = n628 & n6450;
  assign n6918 = n6905 & n6917;
  assign n6919 = n6914 & n6916;
  assign n6920 = n10336 & n10337;
  assign n6921 = n10335 & n6907;
  assign n6922 = n10035 & n10338;
  assign n6923 = n10334 & n6922;
  assign n6924 = n10332 & n10336;
  assign n6925 = n10334 & n6924;
  assign n6926 = n10035 & n6925;
  assign n6927 = ~n626 & n6926;
  assign n6928 = ~n386 & n6927;
  assign n6929 = ~n663 & n6928;
  assign n6930 = ~n627 & n6929;
  assign n6931 = ~n328 & n6930;
  assign n6932 = ~n175 & n6931;
  assign n6933 = ~n582 & n6932;
  assign n6934 = n10332 & n6922;
  assign n6935 = n10334 & n6934;
  assign n6936 = n10332 & n6923;
  assign n6937 = ~n6411 & ~n10339;
  assign n6938 = ~n6411 & ~n6874;
  assign n6939 = ~n10339 & n6938;
  assign n6940 = ~n6874 & n6937;
  assign n6941 = ~n6873 & ~n10340;
  assign n6942 = ~n6755 & ~n10340;
  assign n6943 = ~n10331 & ~n6942;
  assign n6944 = n6755 & n10340;
  assign n6945 = ~n6943 & ~n6944;
  assign n6946 = ~n6872 & ~n6941;
  assign n6947 = ~n6751 & n10341;
  assign n6948 = ~n6750 & ~n10341;
  assign n6949 = ~n6751 & ~n6948;
  assign n6950 = ~n10320 & ~n6751;
  assign n6951 = n6646 & ~n6751;
  assign n6952 = ~n6950 & ~n6951;
  assign n6953 = ~n6750 & ~n6751;
  assign n6954 = ~n10341 & ~n10343;
  assign n6955 = ~n6751 & ~n6954;
  assign n6956 = ~n6750 & ~n6947;
  assign n6957 = n6644 & ~n10342;
  assign n6958 = ~n6644 & n10342;
  assign n6959 = ~n6957 & ~n6958;
  assign n6960 = ~n10343 & ~n6954;
  assign n6961 = n10341 & ~n10343;
  assign n6962 = ~n10341 & ~n6954;
  assign n6963 = ~n10341 & n10343;
  assign n6964 = n10341 & n10343;
  assign n6965 = ~n6954 & ~n6964;
  assign n6966 = ~n10344 & ~n10345;
  assign n6967 = n6959 & n10346;
  assign n6968 = ~n6959 & ~n10346;
  assign n6969 = n6959 & ~n6967;
  assign n6970 = n6959 & ~n10346;
  assign n6971 = n10346 & ~n6967;
  assign n6972 = ~n6959 & n10346;
  assign n6973 = ~n10347 & ~n10348;
  assign n6974 = ~n6967 & ~n6968;
  assign n6975 = pi22  & ~pi23 ;
  assign n6976 = ~pi22  & pi23 ;
  assign n6977 = ~pi22  & ~pi23 ;
  assign n6978 = pi22  & pi23 ;
  assign n6979 = ~n6977 & ~n6978;
  assign n6980 = ~n6975 & ~n6976;
  assign n6981 = ~n10349 & n10350;
  assign n6982 = ~n6643 & ~n6957;
  assign n6983 = ~n6607 & ~n6614;
  assign n6984 = ~n10291 & ~n6498;
  assign n6985 = ~n265 & ~n620;
  assign n6986 = n333 & n6985;
  assign n6987 = n477 & n3844;
  assign n6988 = n4432 & n6987;
  assign n6989 = n477 & n6985;
  assign n6990 = n333 & n3844;
  assign n6991 = n4432 & n6990;
  assign n6992 = n6989 & n6991;
  assign n6993 = n6986 & n6988;
  assign n6994 = n3844 & n4432;
  assign n6995 = n9632 & n6994;
  assign n6996 = n477 & n6995;
  assign n6997 = ~n332 & n6996;
  assign n6998 = ~n265 & n6997;
  assign n6999 = ~n620 & n6998;
  assign n7000 = ~n331 & n6999;
  assign n7001 = n9632 & n10351;
  assign n7002 = n1466 & n1530;
  assign n7003 = ~n230 & ~n674;
  assign n7004 = ~n515 & n7003;
  assign n7005 = ~n9559 & ~n674;
  assign n7006 = ~n230 & ~n515;
  assign n7007 = n7005 & n7006;
  assign n7008 = n353 & n7007;
  assign n7009 = n358 & n7004;
  assign n7010 = n353 & n1530;
  assign n7011 = n1466 & n7010;
  assign n7012 = n7007 & n7011;
  assign n7013 = n7002 & n10353;
  assign n7014 = n9603 & n10354;
  assign n7015 = n9832 & n7014;
  assign n7016 = n10352 & n7015;
  assign n7017 = n9603 & n7010;
  assign n7018 = n9832 & n7017;
  assign n7019 = n10352 & n7018;
  assign n7020 = n10047 & n7019;
  assign n7021 = n1466 & n7020;
  assign n7022 = ~n515 & n7021;
  assign n7023 = ~n230 & n7022;
  assign n7024 = ~n9559 & n7023;
  assign n7025 = ~n674 & n7024;
  assign n7026 = n10047 & n7016;
  assign n7027 = ~n6492 & n10355;
  assign n7028 = ~n6490 & n10355;
  assign n7029 = n6492 & ~n10355;
  assign n7030 = n6490 & ~n10355;
  assign n7031 = ~n6492 & ~n10355;
  assign n7032 = n6492 & n10355;
  assign n7033 = ~n7031 & ~n7032;
  assign n7034 = ~n10356 & ~n10357;
  assign n7035 = ~n6984 & ~n10358;
  assign n7036 = n6984 & n10358;
  assign n7037 = ~n7035 & ~n7036;
  assign n7038 = n5878 & n7037;
  assign n7039 = n5996 & ~n10355;
  assign n7040 = ~n5987 & n10233;
  assign n7041 = n6001 & n6492;
  assign n7042 = n6001 & n6490;
  assign n7043 = ~n7040 & ~n10359;
  assign n7044 = ~n7039 & n7043;
  assign n7045 = ~n7038 & n7044;
  assign n7046 = ~n73 & ~n7045;
  assign n7047 = ~n7045 & ~n7046;
  assign n7048 = n73 & ~n7045;
  assign n7049 = ~n73 & ~n7046;
  assign n7050 = ~n73 & n7045;
  assign n7051 = ~n10360 & ~n10361;
  assign n7052 = ~n6595 & ~n6601;
  assign n7053 = ~n6573 & ~n6580;
  assign n7054 = n4876 & n5108;
  assign n7055 = ~n4870 & n5112;
  assign n7056 = ~n10084 & n5120;
  assign n7057 = n4731 & n10130;
  assign n7058 = ~n7056 & ~n7057;
  assign n7059 = ~n7055 & ~n7057;
  assign n7060 = ~n7056 & n7059;
  assign n7061 = ~n7055 & n7058;
  assign n7062 = ~n7054 & n10362;
  assign n7063 = ~n1703 & ~n7062;
  assign n7064 = ~n7062 & ~n7063;
  assign n7065 = n1703 & ~n7062;
  assign n7066 = ~n1703 & ~n7063;
  assign n7067 = ~n1703 & n7062;
  assign n7068 = ~n10363 & ~n10364;
  assign n7069 = ~n6561 & ~n6567;
  assign n7070 = n4913 & n5368;
  assign n7071 = ~n10085 & n4920;
  assign n7072 = ~n10086 & n10106;
  assign n7073 = n4740 & n4933;
  assign n7074 = ~n7072 & ~n7073;
  assign n7075 = ~n7071 & n7074;
  assign n7076 = ~n4913 & n7075;
  assign n7077 = ~n5368 & n7075;
  assign n7078 = ~n7076 & ~n7077;
  assign n7079 = ~n7070 & n7075;
  assign n7080 = ~n9626 & ~n10365;
  assign n7081 = n9626 & n10365;
  assign n7082 = ~n7080 & ~n7081;
  assign n7083 = ~n1164 & ~n4764;
  assign n7084 = n4958 & n5164;
  assign n7085 = ~n10087 & n4968;
  assign n7086 = n4761 & n10123;
  assign n7087 = ~n10088 & n4966;
  assign n7088 = ~n7086 & ~n7087;
  assign n7089 = ~n7085 & n7088;
  assign n7090 = ~n7084 & n7089;
  assign n7091 = n7083 & ~n7090;
  assign n7092 = ~n7083 & n7090;
  assign n7093 = ~n7091 & ~n7092;
  assign n7094 = ~n1164 & ~n10089;
  assign n7095 = n6538 & n7094;
  assign n7096 = ~n6543 & ~n7095;
  assign n7097 = n7093 & ~n7096;
  assign n7098 = ~n7093 & n7096;
  assign n7099 = ~n7096 & ~n7097;
  assign n7100 = ~n7093 & ~n7096;
  assign n7101 = n7093 & ~n7097;
  assign n7102 = n7093 & n7096;
  assign n7103 = ~n10366 & ~n10367;
  assign n7104 = ~n7097 & ~n7098;
  assign n7105 = n7082 & ~n10368;
  assign n7106 = ~n7082 & n10368;
  assign n7107 = ~n10368 & ~n7105;
  assign n7108 = ~n7082 & ~n10368;
  assign n7109 = n7082 & ~n7105;
  assign n7110 = n7082 & n10368;
  assign n7111 = ~n10369 & ~n10370;
  assign n7112 = ~n7105 & ~n7106;
  assign n7113 = ~n7069 & ~n10371;
  assign n7114 = n7069 & n10371;
  assign n7115 = ~n7069 & ~n7113;
  assign n7116 = ~n7069 & n10371;
  assign n7117 = ~n10371 & ~n7113;
  assign n7118 = n7069 & ~n10371;
  assign n7119 = ~n10372 & ~n10373;
  assign n7120 = ~n7113 & ~n7114;
  assign n7121 = ~n7068 & ~n10374;
  assign n7122 = n7068 & n10374;
  assign n7123 = ~n7068 & ~n7121;
  assign n7124 = ~n10374 & ~n7121;
  assign n7125 = ~n7123 & ~n7124;
  assign n7126 = ~n7121 & ~n7122;
  assign n7127 = n7053 & n10375;
  assign n7128 = ~n7053 & ~n10375;
  assign n7129 = ~n7127 & ~n7128;
  assign n7130 = n90 & n6016;
  assign n7131 = n4878 & n10226;
  assign n7132 = n10100 & n10210;
  assign n7133 = n4886 & ~n5920;
  assign n7134 = ~n7132 & ~n7133;
  assign n7135 = ~n7131 & n7134;
  assign n7136 = ~n90 & n7135;
  assign n7137 = ~n6016 & n7135;
  assign n7138 = ~n7136 & ~n7137;
  assign n7139 = ~n7130 & n7135;
  assign n7140 = ~n9528 & ~n10376;
  assign n7141 = n9528 & n10376;
  assign n7142 = ~n7140 & ~n7141;
  assign n7143 = n7129 & n7142;
  assign n7144 = ~n7129 & ~n7142;
  assign n7145 = n7129 & ~n7143;
  assign n7146 = n7142 & ~n7143;
  assign n7147 = ~n7145 & ~n7146;
  assign n7148 = ~n7143 & ~n7144;
  assign n7149 = ~n7052 & ~n10377;
  assign n7150 = n7052 & n10377;
  assign n7151 = ~n7052 & ~n7149;
  assign n7152 = ~n10377 & ~n7149;
  assign n7153 = ~n7151 & ~n7152;
  assign n7154 = ~n7149 & ~n7150;
  assign n7155 = ~n7051 & ~n10378;
  assign n7156 = n7051 & n10378;
  assign n7157 = ~n7051 & ~n7155;
  assign n7158 = ~n10378 & ~n7155;
  assign n7159 = ~n7157 & ~n7158;
  assign n7160 = ~n7155 & ~n7156;
  assign n7161 = n6983 & n10379;
  assign n7162 = ~n6983 & ~n10379;
  assign n7163 = ~n7161 & ~n7162;
  assign n7164 = ~n404 & ~n754;
  assign n7165 = ~n583 & n7164;
  assign n7166 = ~n1083 & n7165;
  assign n7167 = ~n1083 & n1851;
  assign n7168 = ~n754 & n7167;
  assign n7169 = ~n583 & ~n1083;
  assign n7170 = n7164 & n7169;
  assign n7171 = n1851 & n2536;
  assign n7172 = ~n897 & n10202;
  assign n7173 = n6723 & n7172;
  assign n7174 = n10380 & n7173;
  assign n7175 = ~n327 & n4126;
  assign n7176 = ~n217 & ~n383;
  assign n7177 = ~n470 & n7176;
  assign n7178 = n477 & n1247;
  assign n7179 = n7177 & n7178;
  assign n7180 = n7175 & n7179;
  assign n7181 = n10004 & n7180;
  assign n7182 = ~n265 & ~n383;
  assign n7183 = n1247 & n7182;
  assign n7184 = n477 & n4126;
  assign n7185 = n7183 & n7184;
  assign n7186 = ~n217 & ~n327;
  assign n7187 = ~n470 & ~n897;
  assign n7188 = n7186 & n7187;
  assign n7189 = n10207 & n7188;
  assign n7190 = n10202 & n10380;
  assign n7191 = n7189 & n7190;
  assign n7192 = n7174 & n7180;
  assign n7193 = ~n327 & ~n383;
  assign n7194 = ~n897 & n7193;
  assign n7195 = n10202 & n7194;
  assign n7196 = n10380 & n7195;
  assign n7197 = ~n217 & ~n470;
  assign n7198 = n477 & n7197;
  assign n7199 = n1247 & n4126;
  assign n7200 = n7198 & n7199;
  assign n7201 = n6723 & n7200;
  assign n7202 = n7196 & n7201;
  assign n7203 = n7185 & n7191;
  assign n7204 = n10004 & n10381;
  assign n7205 = n7174 & n7181;
  assign n7206 = n10004 & n7199;
  assign n7207 = n10314 & n7206;
  assign n7208 = n477 & n7207;
  assign n7209 = n10380 & n7208;
  assign n7210 = n10207 & n7209;
  assign n7211 = n10202 & n7210;
  assign n7212 = ~n327 & n7211;
  assign n7213 = ~n383 & n7212;
  assign n7214 = ~n897 & n7213;
  assign n7215 = ~n217 & n7214;
  assign n7216 = ~n265 & n7215;
  assign n7217 = ~n470 & n7216;
  assign n7218 = n10004 & n10314;
  assign n7219 = n10381 & n7218;
  assign n7220 = n10314 & n10381;
  assign n7221 = n10004 & n7220;
  assign n7222 = n10314 & n10382;
  assign n7223 = ~n7163 & n10383;
  assign n7224 = n7163 & ~n10383;
  assign n7225 = ~n7223 & ~n7224;
  assign n7226 = ~n6982 & n7225;
  assign n7227 = n6982 & ~n7225;
  assign n7228 = ~n7226 & ~n7227;
  assign n7229 = n6967 & n7228;
  assign n7230 = ~n6967 & ~n7228;
  assign n7231 = ~n7229 & ~n7230;
  assign n7232 = n6981 & ~n7231;
  assign n7233 = n6981 & ~n7228;
  assign n7234 = ~n6981 & n7231;
  assign n7235 = ~n10384 & ~n7234;
  assign n7236 = ~n7224 & ~n7226;
  assign n7237 = ~n7155 & ~n7162;
  assign n7238 = n10355 & n7035;
  assign n7239 = ~n6492 & ~n6498;
  assign n7240 = ~n6490 & ~n6498;
  assign n7241 = ~n10355 & n10385;
  assign n7242 = ~n6492 & ~n7035;
  assign n7243 = ~n10355 & ~n7242;
  assign n7244 = n10355 & ~n7035;
  assign n7245 = ~n7243 & ~n7244;
  assign n7246 = ~n7238 & ~n7241;
  assign n7247 = n5878 & n10386;
  assign n7248 = n10233 & n6492;
  assign n7249 = n10233 & n6490;
  assign n7250 = n6001 & ~n10355;
  assign n7251 = ~n10387 & ~n7250;
  assign n7252 = ~n7247 & n7251;
  assign n7253 = ~n73 & ~n7252;
  assign n7254 = ~n7252 & ~n7253;
  assign n7255 = n73 & ~n7252;
  assign n7256 = ~n73 & ~n7253;
  assign n7257 = ~n73 & n7252;
  assign n7258 = ~n10388 & ~n10389;
  assign n7259 = ~n7143 & ~n7149;
  assign n7260 = ~n7121 & ~n7128;
  assign n7261 = n5108 & n5778;
  assign n7262 = n5112 & n10210;
  assign n7263 = ~n10084 & n10130;
  assign n7264 = ~n4870 & n5120;
  assign n7265 = ~n7263 & ~n7264;
  assign n7266 = ~n7262 & n7265;
  assign n7267 = ~n7261 & n7266;
  assign n7268 = ~n1703 & ~n7267;
  assign n7269 = ~n7267 & ~n7268;
  assign n7270 = n1703 & ~n7267;
  assign n7271 = ~n1703 & ~n7268;
  assign n7272 = ~n1703 & n7267;
  assign n7273 = ~n10390 & ~n10391;
  assign n7274 = ~n7105 & ~n7113;
  assign n7275 = n4913 & n5414;
  assign n7276 = n4731 & n4920;
  assign n7277 = ~n10085 & n4933;
  assign n7278 = n4740 & n10106;
  assign n7279 = ~n7277 & ~n7278;
  assign n7280 = ~n7276 & ~n7278;
  assign n7281 = ~n7277 & n7280;
  assign n7282 = ~n7276 & n7279;
  assign n7283 = ~n4913 & n10392;
  assign n7284 = ~n5414 & n10392;
  assign n7285 = ~n7283 & ~n7284;
  assign n7286 = ~n7275 & n10392;
  assign n7287 = ~n9626 & ~n10393;
  assign n7288 = n9626 & n10393;
  assign n7289 = ~n7287 & ~n7288;
  assign n7290 = ~n1164 & ~n4761;
  assign n7291 = n4958 & n5145;
  assign n7292 = ~n10086 & n4968;
  assign n7293 = ~n10088 & n10123;
  assign n7294 = ~n10087 & n4966;
  assign n7295 = ~n7293 & ~n7294;
  assign n7296 = ~n7292 & n7295;
  assign n7297 = ~n7291 & n7296;
  assign n7298 = n7290 & ~n7297;
  assign n7299 = ~n7290 & n7297;
  assign n7300 = ~n7298 & ~n7299;
  assign n7301 = ~n1164 & n4764;
  assign n7302 = ~n1164 & n7090;
  assign n7303 = n4764 & n7302;
  assign n7304 = n7090 & n7301;
  assign n7305 = ~n7097 & ~n10394;
  assign n7306 = n7300 & ~n7305;
  assign n7307 = ~n7300 & n7305;
  assign n7308 = ~n7305 & ~n7306;
  assign n7309 = ~n7300 & ~n7305;
  assign n7310 = n7300 & ~n7306;
  assign n7311 = n7300 & n7305;
  assign n7312 = ~n10395 & ~n10396;
  assign n7313 = ~n7306 & ~n7307;
  assign n7314 = n7289 & ~n10397;
  assign n7315 = ~n7289 & n10397;
  assign n7316 = ~n10397 & ~n7314;
  assign n7317 = ~n7289 & ~n10397;
  assign n7318 = n7289 & ~n7314;
  assign n7319 = n7289 & n10397;
  assign n7320 = ~n10398 & ~n10399;
  assign n7321 = ~n7314 & ~n7315;
  assign n7322 = ~n7274 & ~n10400;
  assign n7323 = n7274 & n10400;
  assign n7324 = ~n7274 & ~n7322;
  assign n7325 = ~n7274 & n10400;
  assign n7326 = ~n10400 & ~n7322;
  assign n7327 = n7274 & ~n10400;
  assign n7328 = ~n10401 & ~n10402;
  assign n7329 = ~n7322 & ~n7323;
  assign n7330 = ~n7273 & ~n10403;
  assign n7331 = n7273 & n10403;
  assign n7332 = ~n7273 & ~n7330;
  assign n7333 = ~n10403 & ~n7330;
  assign n7334 = ~n7332 & ~n7333;
  assign n7335 = ~n7330 & ~n7331;
  assign n7336 = n7260 & n10404;
  assign n7337 = ~n7260 & ~n10404;
  assign n7338 = ~n7336 & ~n7337;
  assign n7339 = n90 & n5994;
  assign n7340 = n4878 & ~n5987;
  assign n7341 = n10100 & ~n5920;
  assign n7342 = n4886 & n10226;
  assign n7343 = ~n7341 & ~n7342;
  assign n7344 = ~n7340 & n7343;
  assign n7345 = ~n90 & n7344;
  assign n7346 = ~n5994 & n7344;
  assign n7347 = ~n7345 & ~n7346;
  assign n7348 = ~n7339 & n7344;
  assign n7349 = ~n9528 & ~n10405;
  assign n7350 = n9528 & n10405;
  assign n7351 = ~n7349 & ~n7350;
  assign n7352 = n7338 & n7351;
  assign n7353 = ~n7338 & ~n7351;
  assign n7354 = n7338 & ~n7352;
  assign n7355 = n7351 & ~n7352;
  assign n7356 = ~n7354 & ~n7355;
  assign n7357 = ~n7352 & ~n7353;
  assign n7358 = ~n7259 & ~n10406;
  assign n7359 = n7259 & n10406;
  assign n7360 = ~n7259 & ~n7358;
  assign n7361 = ~n10406 & ~n7358;
  assign n7362 = ~n7360 & ~n7361;
  assign n7363 = ~n7358 & ~n7359;
  assign n7364 = ~n7258 & ~n10407;
  assign n7365 = n7258 & n10407;
  assign n7366 = ~n7258 & ~n7364;
  assign n7367 = ~n10407 & ~n7364;
  assign n7368 = ~n7366 & ~n7367;
  assign n7369 = ~n7364 & ~n7365;
  assign n7370 = ~n7237 & ~n10408;
  assign n7371 = n7237 & n10408;
  assign n7372 = ~n7237 & n10408;
  assign n7373 = n7237 & ~n10408;
  assign n7374 = ~n7372 & ~n7373;
  assign n7375 = ~n7370 & ~n7371;
  assign n7376 = ~n296 & ~n432;
  assign n7377 = ~n398 & ~n432;
  assign n7378 = ~n296 & n7377;
  assign n7379 = ~n398 & n7376;
  assign n7380 = n2074 & n4640;
  assign n7381 = ~n592 & n4640;
  assign n7382 = ~n296 & n7381;
  assign n7383 = ~n432 & n7382;
  assign n7384 = ~n397 & n7383;
  assign n7385 = ~n398 & n7384;
  assign n7386 = ~n397 & ~n432;
  assign n7387 = ~n592 & n7386;
  assign n7388 = ~n296 & ~n398;
  assign n7389 = n4640 & n7388;
  assign n7390 = n7387 & n7389;
  assign n7391 = n10410 & n7380;
  assign n7392 = ~n604 & ~n674;
  assign n7393 = n872 & n7392;
  assign n7394 = n1171 & n7393;
  assign n7395 = ~n380 & ~n757;
  assign n7396 = ~n538 & n7395;
  assign n7397 = n9657 & n7396;
  assign n7398 = ~n538 & ~n604;
  assign n7399 = n872 & n7398;
  assign n7400 = n1171 & n7399;
  assign n7401 = ~n674 & n7395;
  assign n7402 = n9657 & n7401;
  assign n7403 = n7400 & n7402;
  assign n7404 = ~n195 & ~n380;
  assign n7405 = n7392 & n7404;
  assign n7406 = n872 & n7405;
  assign n7407 = ~n538 & ~n757;
  assign n7408 = ~n513 & n7407;
  assign n7409 = n9657 & n7408;
  assign n7410 = n7406 & n7409;
  assign n7411 = n7394 & n7397;
  assign n7412 = n10411 & n10412;
  assign n7413 = n9601 & n7412;
  assign n7414 = n872 & n9657;
  assign n7415 = n9601 & n7414;
  assign n7416 = n10411 & n7415;
  assign n7417 = n10334 & n7416;
  assign n7418 = ~n604 & n7417;
  assign n7419 = ~n757 & n7418;
  assign n7420 = ~n538 & n7419;
  assign n7421 = ~n195 & n7420;
  assign n7422 = ~n380 & n7421;
  assign n7423 = ~n513 & n7422;
  assign n7424 = ~n674 & n7423;
  assign n7425 = n10334 & n7413;
  assign n7426 = ~n10409 & ~n10413;
  assign n7427 = n10409 & n10413;
  assign n7428 = ~n7426 & ~n7427;
  assign n7429 = ~n7236 & ~n7427;
  assign n7430 = ~n7426 & n7429;
  assign n7431 = ~n7236 & n7428;
  assign n7432 = n7236 & ~n7428;
  assign n7433 = ~n7236 & ~n10414;
  assign n7434 = ~n7426 & ~n10414;
  assign n7435 = ~n7427 & n7434;
  assign n7436 = ~n7433 & ~n7435;
  assign n7437 = ~n10414 & ~n7432;
  assign n7438 = ~n7229 & n10415;
  assign n7439 = n7229 & ~n10415;
  assign n7440 = ~n7438 & ~n7439;
  assign n7441 = n10349 & ~n7231;
  assign n7442 = n10350 & ~n7441;
  assign n7443 = n7440 & ~n7442;
  assign n7444 = ~n7440 & n7442;
  assign n7445 = ~n7443 & ~n7444;
  assign n7446 = ~n7440 & n7441;
  assign n7447 = n10350 & ~n7446;
  assign n7448 = ~n7364 & ~n7370;
  assign n7449 = ~n7352 & ~n7358;
  assign n7450 = n5878 & ~n10385;
  assign n7451 = ~n10233 & ~n7450;
  assign n7452 = n10233 & ~n10355;
  assign n7453 = n5878 & n7243;
  assign n7454 = ~n7452 & ~n7453;
  assign n7455 = ~n10355 & ~n7451;
  assign n7456 = ~n73 & ~n10416;
  assign n7457 = ~n10416 & ~n7456;
  assign n7458 = n73 & ~n10416;
  assign n7459 = ~n73 & ~n7456;
  assign n7460 = ~n73 & n10416;
  assign n7461 = ~n10417 & ~n10418;
  assign n7462 = ~n7330 & ~n7337;
  assign n7463 = n5108 & n6034;
  assign n7464 = n5112 & ~n5920;
  assign n7465 = ~n4870 & n10130;
  assign n7466 = n5120 & n10210;
  assign n7467 = ~n7465 & ~n7466;
  assign n7468 = ~n7464 & n7467;
  assign n7469 = ~n7463 & n7468;
  assign n7470 = ~n1703 & ~n7469;
  assign n7471 = ~n7469 & ~n7470;
  assign n7472 = n1703 & ~n7469;
  assign n7473 = ~n1703 & ~n7470;
  assign n7474 = ~n1703 & n7469;
  assign n7475 = ~n10419 & ~n10420;
  assign n7476 = ~n7314 & ~n7322;
  assign n7477 = n4913 & n5396;
  assign n7478 = ~n10084 & n4920;
  assign n7479 = ~n10085 & n10106;
  assign n7480 = n4731 & n4933;
  assign n7481 = ~n7479 & ~n7480;
  assign n7482 = ~n7478 & n7481;
  assign n7483 = ~n4913 & n7482;
  assign n7484 = ~n5396 & n7482;
  assign n7485 = ~n7483 & ~n7484;
  assign n7486 = ~n7477 & n7482;
  assign n7487 = ~n9626 & ~n10421;
  assign n7488 = n9626 & n10421;
  assign n7489 = ~n7487 & ~n7488;
  assign n7490 = ~n1164 & n10088;
  assign n7491 = n4958 & n5110;
  assign n7492 = n4740 & n4968;
  assign n7493 = ~n10086 & n4966;
  assign n7494 = ~n10087 & n10123;
  assign n7495 = ~n7493 & ~n7494;
  assign n7496 = ~n7492 & ~n7494;
  assign n7497 = ~n7493 & n7496;
  assign n7498 = ~n7492 & n7495;
  assign n7499 = ~n7491 & n10422;
  assign n7500 = n7490 & ~n7499;
  assign n7501 = ~n7490 & n7499;
  assign n7502 = ~n7500 & ~n7501;
  assign n7503 = ~n1164 & n4761;
  assign n7504 = ~n1164 & n7297;
  assign n7505 = n4761 & n7504;
  assign n7506 = n7297 & n7503;
  assign n7507 = ~n7306 & ~n10423;
  assign n7508 = n7502 & ~n7507;
  assign n7509 = ~n7502 & n7507;
  assign n7510 = ~n7507 & ~n7508;
  assign n7511 = ~n7502 & ~n7507;
  assign n7512 = n7502 & ~n7508;
  assign n7513 = n7502 & n7507;
  assign n7514 = ~n10424 & ~n10425;
  assign n7515 = ~n7508 & ~n7509;
  assign n7516 = n7489 & ~n10426;
  assign n7517 = ~n7489 & n10426;
  assign n7518 = ~n7516 & ~n7517;
  assign n7519 = ~n7476 & n7518;
  assign n7520 = n7476 & ~n7518;
  assign n7521 = ~n7519 & ~n7520;
  assign n7522 = ~n7475 & n7521;
  assign n7523 = n7475 & ~n7521;
  assign n7524 = ~n7475 & ~n7522;
  assign n7525 = n7521 & ~n7522;
  assign n7526 = ~n7524 & ~n7525;
  assign n7527 = ~n7522 & ~n7523;
  assign n7528 = n7462 & n10427;
  assign n7529 = ~n7462 & ~n10427;
  assign n7530 = ~n7528 & ~n7529;
  assign n7531 = n90 & n6500;
  assign n7532 = n4878 & n6492;
  assign n7533 = n4878 & n6490;
  assign n7534 = n10100 & n10226;
  assign n7535 = n4886 & ~n5987;
  assign n7536 = ~n7534 & ~n7535;
  assign n7537 = ~n10428 & n7536;
  assign n7538 = ~n90 & n7537;
  assign n7539 = ~n6500 & n7537;
  assign n7540 = ~n7538 & ~n7539;
  assign n7541 = ~n7531 & n7537;
  assign n7542 = ~n9528 & ~n10429;
  assign n7543 = n9528 & n10429;
  assign n7544 = ~n7542 & ~n7543;
  assign n7545 = n7530 & n7544;
  assign n7546 = ~n7530 & ~n7544;
  assign n7547 = ~n7545 & ~n7546;
  assign n7548 = ~n7461 & n7547;
  assign n7549 = n7461 & ~n7547;
  assign n7550 = ~n7548 & ~n7549;
  assign n7551 = ~n7449 & n7550;
  assign n7552 = n7449 & ~n7550;
  assign n7553 = ~n7551 & ~n7552;
  assign n7554 = ~n7448 & n7553;
  assign n7555 = n7448 & ~n7553;
  assign n7556 = ~n7554 & ~n7555;
  assign n7557 = n9546 & n9588;
  assign n7558 = n10327 & n7557;
  assign n7559 = ~n715 & ~n720;
  assign n7560 = ~n351 & n7559;
  assign n7561 = ~n663 & ~n754;
  assign n7562 = n899 & n7561;
  assign n7563 = ~n663 & ~n715;
  assign n7564 = ~n351 & n7563;
  assign n7565 = ~n720 & ~n754;
  assign n7566 = n899 & n7565;
  assign n7567 = n7564 & n7566;
  assign n7568 = n7560 & n7562;
  assign n7569 = n1631 & n7175;
  assign n7570 = ~n351 & ~n715;
  assign n7571 = n899 & n7570;
  assign n7572 = n4126 & n7571;
  assign n7573 = ~n327 & ~n663;
  assign n7574 = n7565 & n7573;
  assign n7575 = n1631 & n7574;
  assign n7576 = n7572 & n7575;
  assign n7577 = ~n327 & ~n720;
  assign n7578 = n899 & n7577;
  assign n7579 = n4126 & n7578;
  assign n7580 = ~n351 & ~n754;
  assign n7581 = n7563 & n7580;
  assign n7582 = n1631 & n7581;
  assign n7583 = n7579 & n7582;
  assign n7584 = n10430 & n7569;
  assign n7585 = n9973 & n10431;
  assign n7586 = n7558 & n7585;
  assign n7587 = n4126 & n10327;
  assign n7588 = n899 & n7587;
  assign n7589 = n1631 & n7588;
  assign n7590 = n9973 & n7589;
  assign n7591 = n9829 & n7590;
  assign n7592 = n9588 & n7591;
  assign n7593 = n9546 & n7592;
  assign n7594 = ~n663 & n7593;
  assign n7595 = ~n327 & n7594;
  assign n7596 = ~n715 & n7595;
  assign n7597 = ~n720 & n7596;
  assign n7598 = ~n754 & n7597;
  assign n7599 = ~n351 & n7598;
  assign n7600 = n9829 & n7586;
  assign n7601 = n7556 & ~n10432;
  assign n7602 = ~n7556 & n10432;
  assign n7603 = ~n10432 & ~n7601;
  assign n7604 = n7556 & ~n7601;
  assign n7605 = ~n7603 & ~n7604;
  assign n7606 = ~n7601 & ~n7602;
  assign n7607 = ~n7434 & ~n10433;
  assign n7608 = n7434 & ~n7604;
  assign n7609 = ~n7603 & n7608;
  assign n7610 = n7434 & n10433;
  assign n7611 = ~n7607 & ~n10434;
  assign n7612 = n7439 & n7611;
  assign n7613 = ~n7439 & ~n7611;
  assign n7614 = n7611 & ~n7612;
  assign n7615 = n7439 & ~n7612;
  assign n7616 = ~n7614 & ~n7615;
  assign n7617 = ~n7612 & ~n7613;
  assign n7618 = n7447 & ~n10435;
  assign n7619 = ~n7447 & n10435;
  assign po3  = ~n7618 & ~n7619;
  assign n7621 = ~n7601 & ~n7607;
  assign n7622 = ~n7551 & ~n7554;
  assign n7623 = ~n7545 & ~n7548;
  assign n7624 = ~n7522 & ~n7529;
  assign n7625 = n5108 & n6016;
  assign n7626 = n5112 & n10226;
  assign n7627 = n10130 & n10210;
  assign n7628 = n5120 & ~n5920;
  assign n7629 = ~n7627 & ~n7628;
  assign n7630 = ~n7626 & n7629;
  assign n7631 = ~n7625 & n7630;
  assign n7632 = ~n1703 & ~n7631;
  assign n7633 = ~n1703 & ~n7632;
  assign n7634 = ~n1703 & n7631;
  assign n7635 = ~n7631 & ~n7632;
  assign n7636 = n1703 & ~n7631;
  assign n7637 = ~n10436 & ~n10437;
  assign n7638 = ~n7516 & ~n7519;
  assign n7639 = n4876 & n4913;
  assign n7640 = ~n4870 & n4920;
  assign n7641 = ~n10084 & n4933;
  assign n7642 = n4731 & n10106;
  assign n7643 = ~n7641 & ~n7642;
  assign n7644 = ~n7640 & ~n7642;
  assign n7645 = ~n7641 & n7644;
  assign n7646 = ~n7640 & n7643;
  assign n7647 = ~n7639 & n10438;
  assign n7648 = n9626 & ~n7647;
  assign n7649 = ~n9626 & n7647;
  assign n7650 = ~n7648 & ~n7649;
  assign n7651 = n4958 & n5368;
  assign n7652 = ~n10085 & n4968;
  assign n7653 = ~n10086 & n10123;
  assign n7654 = n4740 & n4966;
  assign n7655 = ~n7653 & ~n7654;
  assign n7656 = ~n7652 & n7655;
  assign n7657 = ~n7651 & n7656;
  assign n7658 = ~n1164 & ~n7657;
  assign n7659 = ~n7657 & ~n7658;
  assign n7660 = n1164 & ~n7657;
  assign n7661 = ~n1164 & ~n7658;
  assign n7662 = ~n1164 & n7657;
  assign n7663 = ~n10439 & ~n10440;
  assign n7664 = ~n73 & ~n1164;
  assign n7665 = ~n1164 & ~n10087;
  assign n7666 = ~n73 & n7665;
  assign n7667 = ~n10087 & n7664;
  assign n7668 = n73 & ~n7665;
  assign n7669 = ~n73 & ~n10441;
  assign n7670 = ~n10087 & ~n10441;
  assign n7671 = ~n1164 & n7670;
  assign n7672 = n7665 & ~n10441;
  assign n7673 = ~n7669 & ~n10442;
  assign n7674 = ~n10441 & ~n7668;
  assign n7675 = ~n7663 & ~n10443;
  assign n7676 = n7663 & n10443;
  assign n7677 = ~n7663 & ~n7675;
  assign n7678 = ~n10443 & ~n7675;
  assign n7679 = ~n7677 & ~n7678;
  assign n7680 = ~n7675 & ~n7676;
  assign n7681 = ~n1164 & ~n10088;
  assign n7682 = n7499 & n7681;
  assign n7683 = ~n7508 & ~n7682;
  assign n7684 = ~n10444 & ~n7683;
  assign n7685 = n10444 & n7683;
  assign n7686 = n10444 & ~n7683;
  assign n7687 = ~n10444 & n7683;
  assign n7688 = ~n7686 & ~n7687;
  assign n7689 = ~n7684 & ~n7685;
  assign n7690 = n7650 & ~n10445;
  assign n7691 = ~n7650 & n10445;
  assign n7692 = ~n10445 & ~n7690;
  assign n7693 = ~n7650 & ~n10445;
  assign n7694 = n7650 & ~n7690;
  assign n7695 = n7650 & n10445;
  assign n7696 = ~n10446 & ~n10447;
  assign n7697 = ~n7690 & ~n7691;
  assign n7698 = ~n7638 & ~n10448;
  assign n7699 = n7638 & n10448;
  assign n7700 = ~n7638 & n10448;
  assign n7701 = n7638 & ~n10448;
  assign n7702 = ~n7700 & ~n7701;
  assign n7703 = ~n7698 & ~n7699;
  assign n7704 = ~n7637 & ~n10449;
  assign n7705 = n7637 & n10449;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = ~n7624 & n7706;
  assign n7708 = n7624 & ~n7706;
  assign n7709 = ~n7707 & ~n7708;
  assign n7710 = n90 & n7037;
  assign n7711 = n4878 & ~n10355;
  assign n7712 = n10100 & ~n5987;
  assign n7713 = n4886 & n6492;
  assign n7714 = n4886 & n6490;
  assign n7715 = ~n7712 & ~n10450;
  assign n7716 = ~n7711 & n7715;
  assign n7717 = ~n7710 & n7716;
  assign n7718 = n9528 & ~n7717;
  assign n7719 = ~n9528 & n7717;
  assign n7720 = ~n7718 & ~n7719;
  assign n7721 = n7709 & n7720;
  assign n7722 = ~n7709 & ~n7720;
  assign n7723 = ~n7721 & ~n7722;
  assign n7724 = ~n7623 & n7723;
  assign n7725 = n7623 & ~n7723;
  assign n7726 = ~n7724 & ~n7725;
  assign n7727 = n7622 & ~n7726;
  assign n7728 = ~n7622 & n7726;
  assign n7729 = ~n7727 & ~n7728;
  assign n7730 = n753 & n4640;
  assign n7731 = n1259 & n7730;
  assign n7732 = ~n325 & ~n682;
  assign n7733 = ~n202 & ~n265;
  assign n7734 = n7732 & n7733;
  assign n7735 = n10044 & n7734;
  assign n7736 = n1111 & n4385;
  assign n7737 = n4640 & n7736;
  assign n7738 = ~n202 & ~n325;
  assign n7739 = ~n682 & n7738;
  assign n7740 = ~n202 & n7732;
  assign n7741 = n753 & n1259;
  assign n7742 = n10451 & n7741;
  assign n7743 = n7737 & n7742;
  assign n7744 = n1111 & n1259;
  assign n7745 = n4385 & n7744;
  assign n7746 = n7730 & n10451;
  assign n7747 = n7745 & n7746;
  assign n7748 = n7731 & n7735;
  assign n7749 = n9700 & n10452;
  assign n7750 = n10062 & n7749;
  assign n7751 = n1111 & n4640;
  assign n7752 = n753 & n7751;
  assign n7753 = n10062 & n7752;
  assign n7754 = n9700 & n7753;
  assign n7755 = n9580 & n7754;
  assign n7756 = n1259 & n7755;
  assign n7757 = n4385 & n7756;
  assign n7758 = ~n325 & n7757;
  assign n7759 = ~n682 & n7758;
  assign n7760 = ~n202 & n7759;
  assign n7761 = n9580 & n7749;
  assign n7762 = n10062 & n7761;
  assign n7763 = n9580 & n7750;
  assign n7764 = ~n7729 & n10453;
  assign n7765 = n7729 & ~n10453;
  assign n7766 = ~n7764 & ~n7765;
  assign n7767 = ~n7621 & n7766;
  assign n7768 = n7621 & ~n7766;
  assign n7769 = ~n7767 & ~n7768;
  assign n7770 = ~n7612 & ~n7769;
  assign n7771 = n7612 & n7769;
  assign n7772 = ~n7770 & ~n7771;
  assign n7773 = n7446 & n10435;
  assign n7774 = n10350 & ~n7773;
  assign n7775 = n7772 & ~n7774;
  assign n7776 = ~n7772 & n7774;
  assign n7777 = ~n7775 & ~n7776;
  assign n7778 = ~n7765 & ~n7767;
  assign n7779 = ~n7724 & ~n7728;
  assign n7780 = ~n7707 & ~n7721;
  assign n7781 = n90 & n10386;
  assign n7782 = n10100 & n6492;
  assign n7783 = n10100 & n6490;
  assign n7784 = n4886 & ~n10355;
  assign n7785 = ~n10454 & ~n7784;
  assign n7786 = ~n7781 & n7785;
  assign n7787 = n9528 & ~n7786;
  assign n7788 = ~n9528 & n7786;
  assign n7789 = ~n7787 & ~n7788;
  assign n7790 = ~n7698 & ~n7704;
  assign n7791 = n5108 & n5994;
  assign n7792 = n5112 & ~n5987;
  assign n7793 = n10130 & ~n5920;
  assign n7794 = n5120 & n10226;
  assign n7795 = ~n7793 & ~n7794;
  assign n7796 = ~n7792 & n7795;
  assign n7797 = ~n7791 & n7796;
  assign n7798 = ~n1703 & ~n7797;
  assign n7799 = ~n7797 & ~n7798;
  assign n7800 = n1703 & ~n7797;
  assign n7801 = ~n1703 & ~n7798;
  assign n7802 = ~n1703 & n7797;
  assign n7803 = ~n10455 & ~n10456;
  assign n7804 = ~n7684 & ~n7690;
  assign n7805 = n4913 & n5778;
  assign n7806 = n4920 & n10210;
  assign n7807 = ~n10084 & n10106;
  assign n7808 = ~n4870 & n4933;
  assign n7809 = ~n7807 & ~n7808;
  assign n7810 = ~n7806 & n7809;
  assign n7811 = ~n7805 & n7810;
  assign n7812 = n9626 & ~n7811;
  assign n7813 = ~n9626 & n7811;
  assign n7814 = ~n7812 & ~n7813;
  assign n7815 = n4958 & n5414;
  assign n7816 = n4731 & n4968;
  assign n7817 = ~n10085 & n4966;
  assign n7818 = n4740 & n10123;
  assign n7819 = ~n7817 & ~n7818;
  assign n7820 = ~n7816 & ~n7818;
  assign n7821 = ~n7817 & n7820;
  assign n7822 = ~n7816 & n7819;
  assign n7823 = ~n4958 & n10457;
  assign n7824 = ~n5414 & n10457;
  assign n7825 = ~n7823 & ~n7824;
  assign n7826 = ~n7815 & n10457;
  assign n7827 = n1164 & ~n10458;
  assign n7828 = ~n1164 & n10458;
  assign n7829 = ~n7827 & ~n7828;
  assign n7830 = ~n10441 & ~n7675;
  assign n7831 = ~n1164 & ~n10086;
  assign n7832 = ~n73 & n7831;
  assign n7833 = ~n10086 & n7664;
  assign n7834 = n73 & ~n7831;
  assign n7835 = ~n73 & ~n10459;
  assign n7836 = ~n10086 & ~n10459;
  assign n7837 = ~n1164 & n7836;
  assign n7838 = n7831 & ~n10459;
  assign n7839 = ~n7835 & ~n10460;
  assign n7840 = ~n10459 & ~n7834;
  assign n7841 = ~n7830 & ~n10461;
  assign n7842 = n7830 & n10461;
  assign n7843 = ~n7830 & ~n7841;
  assign n7844 = ~n10461 & ~n7841;
  assign n7845 = ~n7843 & ~n7844;
  assign n7846 = ~n7841 & ~n7842;
  assign n7847 = n7829 & ~n10462;
  assign n7848 = ~n7829 & n10462;
  assign n7849 = ~n10462 & ~n7847;
  assign n7850 = n7829 & ~n7847;
  assign n7851 = ~n7849 & ~n7850;
  assign n7852 = ~n7847 & ~n7848;
  assign n7853 = n7814 & ~n10463;
  assign n7854 = ~n7814 & ~n7850;
  assign n7855 = ~n7849 & n7854;
  assign n7856 = ~n7814 & n10463;
  assign n7857 = ~n7853 & ~n10464;
  assign n7858 = ~n7804 & n7857;
  assign n7859 = n7804 & ~n7857;
  assign n7860 = ~n7804 & ~n7858;
  assign n7861 = n7857 & ~n7858;
  assign n7862 = ~n7860 & ~n7861;
  assign n7863 = ~n7858 & ~n7859;
  assign n7864 = ~n7803 & ~n10465;
  assign n7865 = n7803 & ~n7861;
  assign n7866 = ~n7860 & n7865;
  assign n7867 = n7803 & n10465;
  assign n7868 = ~n7864 & ~n10466;
  assign n7869 = ~n7790 & n7868;
  assign n7870 = n7790 & ~n7868;
  assign n7871 = ~n7790 & ~n7869;
  assign n7872 = n7868 & ~n7869;
  assign n7873 = ~n7871 & ~n7872;
  assign n7874 = ~n7869 & ~n7870;
  assign n7875 = n7789 & ~n10467;
  assign n7876 = ~n7789 & ~n7872;
  assign n7877 = ~n7871 & n7876;
  assign n7878 = ~n7789 & n10467;
  assign n7879 = ~n7875 & ~n10468;
  assign n7880 = ~n7780 & n7879;
  assign n7881 = n7780 & ~n7879;
  assign n7882 = ~n7880 & ~n7881;
  assign n7883 = ~n7779 & n7882;
  assign n7884 = n7779 & ~n7882;
  assign n7885 = ~n7883 & ~n7884;
  assign n7886 = ~n325 & ~n772;
  assign n7887 = ~n9550 & ~n300;
  assign n7888 = ~n300 & ~n325;
  assign n7889 = ~n9550 & ~n772;
  assign n7890 = n7888 & n7889;
  assign n7891 = n7886 & n7887;
  assign n7892 = n775 & n909;
  assign n7893 = n10469 & n7892;
  assign n7894 = ~n618 & n831;
  assign n7895 = n826 & n4024;
  assign n7896 = ~n431 & ~n663;
  assign n7897 = ~n663 & n4421;
  assign n7898 = ~n476 & n7896;
  assign n7899 = n10470 & n10471;
  assign n7900 = n7893 & n7899;
  assign n7901 = n10015 & n10380;
  assign n7902 = n7893 & n10471;
  assign n7903 = n10470 & n7901;
  assign n7904 = n7902 & n7903;
  assign n7905 = n10380 & n10469;
  assign n7906 = n10471 & n7905;
  assign n7907 = n826 & n909;
  assign n7908 = n775 & n4024;
  assign n7909 = n7892 & n10470;
  assign n7910 = n7907 & n7908;
  assign n7911 = n10015 & n10473;
  assign n7912 = n7906 & n7911;
  assign n7913 = n7900 & n7901;
  assign n7914 = n10206 & n10472;
  assign n7915 = n775 & n826;
  assign n7916 = n10471 & n7915;
  assign n7917 = n10015 & n7916;
  assign n7918 = n909 & n7917;
  assign n7919 = n10352 & n7918;
  assign n7920 = n10206 & n7919;
  assign n7921 = n10380 & n7920;
  assign n7922 = n4024 & n7921;
  assign n7923 = ~n325 & n7922;
  assign n7924 = ~n9550 & n7923;
  assign n7925 = ~n772 & n7924;
  assign n7926 = ~n300 & n7925;
  assign n7927 = n10206 & n10352;
  assign n7928 = n10472 & n7927;
  assign n7929 = n10352 & n7914;
  assign n7930 = ~n7885 & n10474;
  assign n7931 = n7885 & ~n10474;
  assign n7932 = ~n7930 & ~n7931;
  assign n7933 = ~n7778 & n7932;
  assign n7934 = n7778 & ~n7932;
  assign n7935 = ~n7933 & ~n7934;
  assign n7936 = ~n7771 & ~n7935;
  assign n7937 = n7771 & n7935;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = ~n7772 & n7773;
  assign n7940 = n10350 & ~n7939;
  assign n7941 = n7938 & ~n7940;
  assign n7942 = ~n7938 & n7940;
  assign n7943 = ~n7941 & ~n7942;
  assign n7944 = ~n7931 & ~n7933;
  assign n7945 = ~n7880 & ~n7883;
  assign n7946 = ~n7869 & ~n7875;
  assign n7947 = ~n7858 & ~n7864;
  assign n7948 = n90 & ~n10385;
  assign n7949 = ~n10100 & ~n7948;
  assign n7950 = n10100 & ~n10355;
  assign n7951 = n90 & n7243;
  assign n7952 = ~n7950 & ~n7951;
  assign n7953 = ~n10355 & ~n7949;
  assign n7954 = ~n9528 & ~n10475;
  assign n7955 = n9528 & n10475;
  assign n7956 = ~n7954 & ~n7955;
  assign n7957 = ~n7947 & ~n7956;
  assign n7958 = n7947 & n7956;
  assign n7959 = ~n7957 & ~n7958;
  assign n7960 = n5108 & n6500;
  assign n7961 = n5112 & n6492;
  assign n7962 = n5112 & n6490;
  assign n7963 = n10130 & n10226;
  assign n7964 = n5120 & ~n5987;
  assign n7965 = ~n7963 & ~n7964;
  assign n7966 = ~n10476 & n7965;
  assign n7967 = ~n7960 & n7966;
  assign n7968 = ~n1703 & ~n7967;
  assign n7969 = ~n7967 & ~n7968;
  assign n7970 = n1703 & ~n7967;
  assign n7971 = ~n1703 & ~n7968;
  assign n7972 = ~n1703 & n7967;
  assign n7973 = ~n10477 & ~n10478;
  assign n7974 = ~n7847 & ~n7853;
  assign n7975 = n4913 & n6034;
  assign n7976 = n4920 & ~n5920;
  assign n7977 = ~n4870 & n10106;
  assign n7978 = n4933 & n10210;
  assign n7979 = ~n7977 & ~n7978;
  assign n7980 = ~n7976 & n7979;
  assign n7981 = ~n7975 & n7980;
  assign n7982 = n9626 & ~n7981;
  assign n7983 = ~n9626 & n7981;
  assign n7984 = ~n7982 & ~n7983;
  assign n7985 = n4958 & n5396;
  assign n7986 = ~n10084 & n4968;
  assign n7987 = ~n10085 & n10123;
  assign n7988 = n4731 & n4966;
  assign n7989 = ~n7987 & ~n7988;
  assign n7990 = ~n7986 & n7989;
  assign n7991 = ~n4958 & n7990;
  assign n7992 = ~n5396 & n7990;
  assign n7993 = ~n7991 & ~n7992;
  assign n7994 = ~n7985 & n7990;
  assign n7995 = n1164 & ~n10479;
  assign n7996 = ~n1164 & n10479;
  assign n7997 = ~n7995 & ~n7996;
  assign n7998 = ~n10459 & ~n7841;
  assign n7999 = ~n1164 & n4740;
  assign n8000 = ~n73 & n7999;
  assign n8001 = n4740 & n7664;
  assign n8002 = n73 & ~n7999;
  assign n8003 = ~n73 & ~n10480;
  assign n8004 = n4740 & ~n10480;
  assign n8005 = ~n1164 & n8004;
  assign n8006 = n7999 & ~n10480;
  assign n8007 = ~n8003 & ~n10481;
  assign n8008 = ~n10480 & ~n8002;
  assign n8009 = ~n7998 & ~n10482;
  assign n8010 = n7998 & n10482;
  assign n8011 = ~n7998 & ~n8009;
  assign n8012 = ~n10482 & ~n8009;
  assign n8013 = ~n8011 & ~n8012;
  assign n8014 = ~n8009 & ~n8010;
  assign n8015 = n7997 & ~n10483;
  assign n8016 = ~n7997 & n10483;
  assign n8017 = ~n10483 & ~n8015;
  assign n8018 = n7997 & ~n8015;
  assign n8019 = ~n8017 & ~n8018;
  assign n8020 = ~n8015 & ~n8016;
  assign n8021 = n7984 & ~n10484;
  assign n8022 = ~n7984 & ~n8018;
  assign n8023 = ~n8017 & n8022;
  assign n8024 = ~n7984 & n10484;
  assign n8025 = ~n8021 & ~n10485;
  assign n8026 = ~n7974 & n8025;
  assign n8027 = n7974 & ~n8025;
  assign n8028 = ~n7974 & ~n8026;
  assign n8029 = n8025 & ~n8026;
  assign n8030 = ~n8028 & ~n8029;
  assign n8031 = ~n8026 & ~n8027;
  assign n8032 = ~n7973 & ~n10486;
  assign n8033 = n7973 & ~n8029;
  assign n8034 = ~n8028 & n8033;
  assign n8035 = n7973 & n10486;
  assign n8036 = ~n8032 & ~n10487;
  assign n8037 = n7959 & n8036;
  assign n8038 = ~n7959 & ~n8036;
  assign n8039 = ~n8037 & ~n8038;
  assign n8040 = ~n7946 & n8039;
  assign n8041 = n7946 & ~n8039;
  assign n8042 = ~n8040 & ~n8041;
  assign n8043 = ~n7945 & n8042;
  assign n8044 = n7945 & ~n8042;
  assign n8045 = ~n8043 & ~n8044;
  assign n8046 = n385 & ~n676;
  assign n8047 = n197 & n8046;
  assign n8048 = n7002 & n8047;
  assign n8049 = n1839 & n4024;
  assign n8050 = n4024 & n4126;
  assign n8051 = n1839 & n8050;
  assign n8052 = n4126 & n8049;
  assign n8053 = n10045 & n10488;
  assign n8054 = n1530 & n1839;
  assign n8055 = n197 & n8054;
  assign n8056 = n10045 & n8055;
  assign n8057 = n4126 & n8056;
  assign n8058 = n385 & n8057;
  assign n8059 = n4024 & n8058;
  assign n8060 = n1466 & n8059;
  assign n8061 = ~n676 & n8060;
  assign n8062 = n1530 & n4024;
  assign n8063 = n8046 & n8062;
  assign n8064 = n197 & n8063;
  assign n8065 = n1466 & n1839;
  assign n8066 = n4126 & n8065;
  assign n8067 = n10045 & n8066;
  assign n8068 = n8064 & n8067;
  assign n8069 = n8048 & n8053;
  assign n8070 = n1482 & n4028;
  assign n8071 = n5921 & n8070;
  assign n8072 = ~n335 & ~n386;
  assign n8073 = ~n332 & ~n381;
  assign n8074 = ~n335 & ~n381;
  assign n8075 = ~n332 & ~n386;
  assign n8076 = n8074 & n8075;
  assign n8077 = n8072 & n8073;
  assign n8078 = n10059 & n10490;
  assign n8079 = ~n332 & ~n335;
  assign n8080 = n4028 & n8079;
  assign n8081 = ~n381 & ~n386;
  assign n8082 = n1482 & n8081;
  assign n8083 = n5921 & n8082;
  assign n8084 = n8080 & n8083;
  assign n8085 = n10059 & n8084;
  assign n8086 = n8071 & n8078;
  assign n8087 = n10489 & n10491;
  assign n8088 = n1482 & n10316;
  assign n8089 = n10059 & n8088;
  assign n8090 = n5921 & n8089;
  assign n8091 = n10489 & n8090;
  assign n8092 = ~n225 & n8091;
  assign n8093 = ~n386 & n8092;
  assign n8094 = ~n335 & n8093;
  assign n8095 = ~n332 & n8094;
  assign n8096 = ~n9586 & n8095;
  assign n8097 = ~n381 & n8096;
  assign n8098 = n10316 & n8087;
  assign n8099 = ~n8045 & n10492;
  assign n8100 = n8045 & ~n10492;
  assign n8101 = ~n8099 & ~n8100;
  assign n8102 = ~n7944 & n8101;
  assign n8103 = n7944 & ~n8101;
  assign n8104 = ~n8102 & ~n8103;
  assign n8105 = ~n7937 & ~n8104;
  assign n8106 = n7937 & n8104;
  assign n8107 = ~n8105 & ~n8106;
  assign n8108 = ~n7938 & n7939;
  assign n8109 = n10350 & ~n8108;
  assign n8110 = n8107 & ~n8109;
  assign n8111 = ~n8107 & n8109;
  assign n8112 = ~n8110 & ~n8111;
  assign n8113 = ~n8100 & ~n8102;
  assign n8114 = ~n8040 & ~n8043;
  assign n8115 = ~n7957 & ~n8037;
  assign n8116 = ~n8026 & ~n8032;
  assign n8117 = n5108 & n7037;
  assign n8118 = n5112 & ~n10355;
  assign n8119 = n10130 & ~n5987;
  assign n8120 = n5120 & n6492;
  assign n8121 = n5120 & n6490;
  assign n8122 = ~n8119 & ~n10493;
  assign n8123 = ~n8118 & n8122;
  assign n8124 = ~n7037 & n8123;
  assign n8125 = ~n5108 & n8123;
  assign n8126 = ~n8124 & ~n8125;
  assign n8127 = ~n8117 & n8123;
  assign n8128 = n1703 & ~n10494;
  assign n8129 = ~n1703 & n10494;
  assign n8130 = ~n8128 & ~n8129;
  assign n8131 = ~n8116 & n8130;
  assign n8132 = n8116 & ~n8130;
  assign n8133 = ~n8131 & ~n8132;
  assign n8134 = ~n8015 & ~n8021;
  assign n8135 = n4913 & n6016;
  assign n8136 = n4920 & n10226;
  assign n8137 = n10106 & n10210;
  assign n8138 = n4933 & ~n5920;
  assign n8139 = ~n8137 & ~n8138;
  assign n8140 = ~n8136 & n8139;
  assign n8141 = ~n4913 & n8140;
  assign n8142 = ~n6016 & n8140;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = ~n8135 & n8140;
  assign n8145 = ~n9626 & ~n10495;
  assign n8146 = n9626 & n10495;
  assign n8147 = ~n8145 & ~n8146;
  assign n8148 = ~n10480 & ~n8009;
  assign n8149 = n4876 & n4958;
  assign n8150 = ~n4870 & n4968;
  assign n8151 = ~n10084 & n4966;
  assign n8152 = n4731 & n10123;
  assign n8153 = ~n8151 & ~n8152;
  assign n8154 = ~n8150 & ~n8152;
  assign n8155 = ~n8151 & n8154;
  assign n8156 = ~n8150 & n8153;
  assign n8157 = ~n8149 & n10496;
  assign n8158 = ~n1164 & ~n8157;
  assign n8159 = ~n8157 & ~n8158;
  assign n8160 = n1164 & ~n8157;
  assign n8161 = ~n1164 & ~n8158;
  assign n8162 = ~n1164 & n8157;
  assign n8163 = ~n10497 & ~n10498;
  assign n8164 = ~n1164 & ~n10085;
  assign n8165 = ~n9528 & n73;
  assign n8166 = n9528 & ~n73;
  assign n8167 = ~n8165 & ~n8166;
  assign n8168 = n8164 & n8167;
  assign n8169 = ~n8164 & ~n8167;
  assign n8170 = ~n8168 & ~n8169;
  assign n8171 = ~n8163 & n8170;
  assign n8172 = n8163 & ~n8170;
  assign n8173 = ~n8163 & ~n8171;
  assign n8174 = ~n8163 & ~n8170;
  assign n8175 = n8170 & ~n8171;
  assign n8176 = n8163 & n8170;
  assign n8177 = ~n10499 & ~n10500;
  assign n8178 = ~n8171 & ~n8172;
  assign n8179 = ~n8148 & ~n10501;
  assign n8180 = n8148 & n10501;
  assign n8181 = ~n8148 & n10501;
  assign n8182 = n8148 & ~n10501;
  assign n8183 = ~n8181 & ~n8182;
  assign n8184 = ~n8179 & ~n8180;
  assign n8185 = n8147 & ~n10502;
  assign n8186 = ~n8147 & n10502;
  assign n8187 = ~n10502 & ~n8185;
  assign n8188 = n8147 & ~n8185;
  assign n8189 = ~n8187 & ~n8188;
  assign n8190 = ~n8185 & ~n8186;
  assign n8191 = ~n8134 & ~n10503;
  assign n8192 = n8134 & n10503;
  assign n8193 = ~n8134 & ~n8191;
  assign n8194 = ~n10503 & ~n8191;
  assign n8195 = ~n8193 & ~n8194;
  assign n8196 = ~n8191 & ~n8192;
  assign n8197 = n8133 & ~n10504;
  assign n8198 = ~n8133 & n10504;
  assign n8199 = n8133 & ~n8197;
  assign n8200 = ~n10504 & ~n8197;
  assign n8201 = ~n8199 & ~n8200;
  assign n8202 = ~n8197 & ~n8198;
  assign n8203 = ~n8115 & ~n10505;
  assign n8204 = n8115 & n10505;
  assign n8205 = ~n8115 & n10505;
  assign n8206 = n8115 & ~n10505;
  assign n8207 = ~n8205 & ~n8206;
  assign n8208 = ~n8203 & ~n8204;
  assign n8209 = n8114 & n10506;
  assign n8210 = ~n8114 & ~n10506;
  assign n8211 = ~n8209 & ~n8210;
  assign n8212 = n758 & n1611;
  assign n8213 = ~n175 & ~n682;
  assign n8214 = n1817 & n8213;
  assign n8215 = n8212 & n8214;
  assign n8216 = ~n296 & ~n470;
  assign n8217 = n603 & n8216;
  assign n8218 = n10471 & n8217;
  assign n8219 = ~n296 & ~n415;
  assign n8220 = n758 & n8219;
  assign n8221 = n1611 & n1817;
  assign n8222 = n8220 & n8221;
  assign n8223 = ~n331 & ~n682;
  assign n8224 = ~n175 & ~n470;
  assign n8225 = n8223 & n8224;
  assign n8226 = n10471 & n8225;
  assign n8227 = n8222 & n8226;
  assign n8228 = n8215 & n8218;
  assign n8229 = n10489 & n10507;
  assign n8230 = n1611 & n10003;
  assign n8231 = n10471 & n8230;
  assign n8232 = n758 & n8231;
  assign n8233 = n10489 & n8232;
  assign n8234 = ~n296 & n8233;
  assign n8235 = ~n682 & n8234;
  assign n8236 = ~n415 & n8235;
  assign n8237 = ~n175 & n8236;
  assign n8238 = n1817 & n8237;
  assign n8239 = ~n331 & n8238;
  assign n8240 = ~n470 & n8239;
  assign n8241 = n10003 & n8229;
  assign n8242 = n8211 & ~n10508;
  assign n8243 = ~n8211 & n10508;
  assign n8244 = ~n8242 & ~n8243;
  assign n8245 = ~n8113 & n8244;
  assign n8246 = n8113 & ~n8244;
  assign n8247 = ~n8245 & ~n8246;
  assign n8248 = n8106 & n8247;
  assign n8249 = ~n8106 & ~n8247;
  assign n8250 = ~n8248 & ~n8249;
  assign n8251 = ~n8107 & n8108;
  assign n8252 = n10350 & ~n8251;
  assign n8253 = n8250 & ~n8252;
  assign n8254 = ~n8250 & n8252;
  assign n8255 = ~n8253 & ~n8254;
  assign n8256 = ~n8242 & ~n8245;
  assign n8257 = ~n8203 & ~n8210;
  assign n8258 = ~n8131 & ~n8197;
  assign n8259 = n5108 & n10386;
  assign n8260 = n10130 & n6492;
  assign n8261 = n10130 & n6490;
  assign n8262 = n5120 & ~n10355;
  assign n8263 = ~n10509 & ~n8262;
  assign n8264 = ~n8259 & n8263;
  assign n8265 = ~n1703 & ~n8264;
  assign n8266 = ~n8264 & ~n8265;
  assign n8267 = n1703 & ~n8264;
  assign n8268 = ~n1703 & ~n8265;
  assign n8269 = ~n1703 & n8264;
  assign n8270 = ~n10510 & ~n10511;
  assign n8271 = ~n8185 & ~n8191;
  assign n8272 = n4913 & n5994;
  assign n8273 = n4920 & ~n5987;
  assign n8274 = n10106 & ~n5920;
  assign n8275 = n4933 & n10226;
  assign n8276 = ~n8274 & ~n8275;
  assign n8277 = ~n8273 & n8276;
  assign n8278 = ~n8272 & n8277;
  assign n8279 = n9626 & ~n8278;
  assign n8280 = ~n9626 & n8278;
  assign n8281 = ~n8279 & ~n8280;
  assign n8282 = ~n8171 & ~n8179;
  assign n8283 = n4958 & n5778;
  assign n8284 = n4968 & n10210;
  assign n8285 = ~n10084 & n10123;
  assign n8286 = ~n4870 & n4966;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = ~n8284 & n8287;
  assign n8289 = ~n4958 & n8288;
  assign n8290 = ~n5778 & n8288;
  assign n8291 = ~n8289 & ~n8290;
  assign n8292 = ~n8283 & n8288;
  assign n8293 = n1164 & ~n10512;
  assign n8294 = ~n1164 & n10512;
  assign n8295 = ~n8293 & ~n8294;
  assign n8296 = ~n1164 & n4731;
  assign n8297 = ~n8165 & ~n8168;
  assign n8298 = ~n8296 & ~n8297;
  assign n8299 = n8296 & n8297;
  assign n8300 = ~n8296 & ~n8298;
  assign n8301 = ~n8296 & n8297;
  assign n8302 = ~n8297 & ~n8298;
  assign n8303 = n8296 & ~n8297;
  assign n8304 = ~n10513 & ~n10514;
  assign n8305 = ~n8298 & ~n8299;
  assign n8306 = n8295 & ~n10515;
  assign n8307 = ~n8295 & n10515;
  assign n8308 = ~n8306 & ~n8307;
  assign n8309 = ~n8282 & n8308;
  assign n8310 = n8282 & ~n8308;
  assign n8311 = ~n8282 & ~n8309;
  assign n8312 = n8308 & ~n8309;
  assign n8313 = ~n8311 & ~n8312;
  assign n8314 = ~n8309 & ~n8310;
  assign n8315 = n8281 & ~n10516;
  assign n8316 = ~n8281 & ~n8312;
  assign n8317 = ~n8311 & n8316;
  assign n8318 = ~n8281 & n10516;
  assign n8319 = ~n8315 & ~n10517;
  assign n8320 = ~n8271 & n8319;
  assign n8321 = n8271 & ~n8319;
  assign n8322 = ~n8320 & ~n8321;
  assign n8323 = ~n8270 & n8322;
  assign n8324 = n8270 & ~n8322;
  assign n8325 = ~n8323 & ~n8324;
  assign n8326 = ~n8258 & n8325;
  assign n8327 = n8258 & ~n8325;
  assign n8328 = ~n8326 & ~n8327;
  assign n8329 = ~n8257 & n8328;
  assign n8330 = n8257 & ~n8328;
  assign n8331 = ~n8329 & ~n8330;
  assign n8332 = ~n479 & n822;
  assign n8333 = n664 & n996;
  assign n8334 = n4268 & n8333;
  assign n8335 = ~n479 & n664;
  assign n8336 = n822 & n996;
  assign n8337 = n4268 & n8336;
  assign n8338 = n8335 & n8337;
  assign n8339 = ~n995 & n3829;
  assign n8340 = ~n219 & ~n720;
  assign n8341 = ~n479 & ~n627;
  assign n8342 = n8340 & n8341;
  assign n8343 = n664 & n8342;
  assign n8344 = n8339 & n8343;
  assign n8345 = n8332 & n8334;
  assign n8346 = n9980 & n10518;
  assign n8347 = n664 & n9980;
  assign n8348 = n9567 & n8347;
  assign n8349 = ~n9561 & n8348;
  assign n8350 = ~n627 & n8349;
  assign n8351 = ~n219 & n8350;
  assign n8352 = ~n9551 & n8351;
  assign n8353 = ~n995 & n8352;
  assign n8354 = ~n720 & n8353;
  assign n8355 = ~n479 & n8354;
  assign n8356 = n9567 & n8346;
  assign n8357 = ~n592 & ~n898;
  assign n8358 = ~n1015 & n8357;
  assign n8359 = ~n467 & ~n1083;
  assign n8360 = n4133 & n8359;
  assign n8361 = ~n898 & ~n1083;
  assign n8362 = ~n1015 & n8361;
  assign n8363 = ~n467 & ~n592;
  assign n8364 = n4133 & n8363;
  assign n8365 = n8362 & n8364;
  assign n8366 = ~n592 & ~n1083;
  assign n8367 = ~n260 & n8366;
  assign n8368 = ~n898 & ~n1015;
  assign n8369 = ~n467 & ~n674;
  assign n8370 = n8368 & n8369;
  assign n8371 = n8367 & n8370;
  assign n8372 = n8358 & n8360;
  assign n8373 = n9701 & n10024;
  assign n8374 = n10520 & n8373;
  assign n8375 = n9697 & n8374;
  assign n8376 = n10325 & n8375;
  assign n8377 = n9697 & n8373;
  assign n8378 = n10325 & n8377;
  assign n8379 = n10519 & n8378;
  assign n8380 = ~n592 & n8379;
  assign n8381 = ~n467 & n8380;
  assign n8382 = ~n898 & n8381;
  assign n8383 = ~n1083 & n8382;
  assign n8384 = ~n1015 & n8383;
  assign n8385 = ~n674 & n8384;
  assign n8386 = ~n260 & n8385;
  assign n8387 = n10519 & n8376;
  assign n8388 = ~n8331 & n10521;
  assign n8389 = n8331 & ~n10521;
  assign n8390 = ~n8388 & ~n8389;
  assign n8391 = ~n8256 & n8390;
  assign n8392 = n8256 & ~n8390;
  assign n8393 = ~n8391 & ~n8392;
  assign n8394 = ~n8248 & ~n8393;
  assign n8395 = n8248 & n8393;
  assign n8396 = ~n8394 & ~n8395;
  assign n8397 = ~n8250 & n8251;
  assign n8398 = n10350 & ~n8397;
  assign n8399 = n8396 & ~n8398;
  assign n8400 = ~n8396 & n8398;
  assign n8401 = ~n8399 & ~n8400;
  assign n8402 = ~n8389 & ~n8391;
  assign n8403 = ~n8326 & ~n8329;
  assign n8404 = ~n8320 & ~n8323;
  assign n8405 = ~n8309 & ~n8315;
  assign n8406 = n5108 & ~n10385;
  assign n8407 = ~n10130 & ~n8406;
  assign n8408 = n10130 & ~n10355;
  assign n8409 = n5108 & n7243;
  assign n8410 = ~n8408 & ~n8409;
  assign n8411 = ~n10355 & ~n8407;
  assign n8412 = ~n1703 & n10522;
  assign n8413 = n1703 & ~n10522;
  assign n8414 = ~n8412 & ~n8413;
  assign n8415 = ~n8405 & ~n8414;
  assign n8416 = n8405 & n8414;
  assign n8417 = ~n8415 & ~n8416;
  assign n8418 = n4913 & n6500;
  assign n8419 = n4920 & n6492;
  assign n8420 = n4920 & n6490;
  assign n8421 = n10106 & n10226;
  assign n8422 = n4933 & ~n5987;
  assign n8423 = ~n8421 & ~n8422;
  assign n8424 = ~n10523 & n8423;
  assign n8425 = ~n8418 & n8424;
  assign n8426 = n9626 & ~n8425;
  assign n8427 = ~n9626 & n8425;
  assign n8428 = ~n8426 & ~n8427;
  assign n8429 = ~n8298 & ~n8306;
  assign n8430 = n4958 & n6034;
  assign n8431 = n4968 & ~n5920;
  assign n8432 = ~n4870 & n10123;
  assign n8433 = n4966 & n10210;
  assign n8434 = ~n8432 & ~n8433;
  assign n8435 = ~n8431 & n8434;
  assign n8436 = ~n8430 & n8435;
  assign n8437 = ~n1164 & ~n8436;
  assign n8438 = ~n8436 & ~n8437;
  assign n8439 = n1164 & ~n8436;
  assign n8440 = ~n1164 & ~n8437;
  assign n8441 = ~n1164 & n8436;
  assign n8442 = ~n10524 & ~n10525;
  assign n8443 = ~n1164 & n4822;
  assign n8444 = ~n8442 & ~n8443;
  assign n8445 = n8442 & n8443;
  assign n8446 = ~n8442 & ~n8444;
  assign n8447 = ~n8443 & ~n8444;
  assign n8448 = ~n8446 & ~n8447;
  assign n8449 = ~n8444 & ~n8445;
  assign n8450 = ~n8429 & ~n10526;
  assign n8451 = n8429 & n10526;
  assign n8452 = ~n8429 & n10526;
  assign n8453 = n8429 & ~n10526;
  assign n8454 = ~n8452 & ~n8453;
  assign n8455 = ~n8450 & ~n8451;
  assign n8456 = n8428 & ~n10527;
  assign n8457 = ~n8428 & n10527;
  assign n8458 = ~n10527 & ~n8456;
  assign n8459 = n8428 & ~n8456;
  assign n8460 = ~n8458 & ~n8459;
  assign n8461 = ~n8456 & ~n8457;
  assign n8462 = n8417 & ~n10528;
  assign n8463 = ~n8417 & n10528;
  assign n8464 = ~n10528 & ~n8462;
  assign n8465 = n8417 & ~n8462;
  assign n8466 = ~n8464 & ~n8465;
  assign n8467 = ~n8462 & ~n8463;
  assign n8468 = ~n8404 & ~n10529;
  assign n8469 = n8404 & n10529;
  assign n8470 = ~n8404 & n10529;
  assign n8471 = n8404 & ~n10529;
  assign n8472 = ~n8470 & ~n8471;
  assign n8473 = ~n8468 & ~n8469;
  assign n8474 = n8403 & n10530;
  assign n8475 = ~n8403 & ~n10530;
  assign n8476 = ~n8474 & ~n8475;
  assign n8477 = ~n190 & ~n243;
  assign n8478 = ~n9551 & ~n301;
  assign n8479 = n8477 & n8478;
  assign n8480 = ~n225 & ~n394;
  assign n8481 = n758 & n8480;
  assign n8482 = n5921 & n8481;
  assign n8483 = ~n190 & ~n394;
  assign n8484 = n8478 & n8483;
  assign n8485 = ~n225 & ~n243;
  assign n8486 = n758 & n8485;
  assign n8487 = n5921 & n8486;
  assign n8488 = n8484 & n8487;
  assign n8489 = n8479 & n8482;
  assign n8490 = n9571 & n7172;
  assign n8491 = ~n243 & ~n394;
  assign n8492 = n8478 & n8491;
  assign n8493 = n758 & n5921;
  assign n8494 = n8492 & n8493;
  assign n8495 = ~n225 & ~n897;
  assign n8496 = ~n190 & n8495;
  assign n8497 = n10202 & n8496;
  assign n8498 = ~n9551 & ~n394;
  assign n8499 = n8485 & n8498;
  assign n8500 = n8493 & n8499;
  assign n8501 = ~n190 & ~n301;
  assign n8502 = ~n897 & n8501;
  assign n8503 = n10202 & n8502;
  assign n8504 = n8500 & n8503;
  assign n8505 = n8494 & n8497;
  assign n8506 = n9571 & n10532;
  assign n8507 = n10531 & n8490;
  assign n8508 = n10317 & n10533;
  assign n8509 = n9571 & n758;
  assign n8510 = n10317 & n8509;
  assign n8511 = n10202 & n8510;
  assign n8512 = n10047 & n8511;
  assign n8513 = n5921 & n8512;
  assign n8514 = ~n225 & n8513;
  assign n8515 = ~n897 & n8514;
  assign n8516 = ~n9551 & n8515;
  assign n8517 = ~n394 & n8516;
  assign n8518 = ~n301 & n8517;
  assign n8519 = ~n190 & n8518;
  assign n8520 = ~n243 & n8519;
  assign n8521 = n10047 & n8508;
  assign n8522 = ~n8476 & n10534;
  assign n8523 = n8476 & ~n10534;
  assign n8524 = ~n8522 & ~n8523;
  assign n8525 = ~n8402 & n8524;
  assign n8526 = n8402 & ~n8524;
  assign n8527 = ~n8525 & ~n8526;
  assign n8528 = ~n8395 & ~n8527;
  assign n8529 = n8395 & n8527;
  assign n8530 = ~n8528 & ~n8529;
  assign n8531 = ~n8396 & n8397;
  assign n8532 = n10350 & ~n8531;
  assign n8533 = n8530 & ~n8532;
  assign n8534 = ~n8530 & n8532;
  assign n8535 = ~n8533 & ~n8534;
  assign n8536 = ~n8523 & ~n8525;
  assign n8537 = ~n8468 & ~n8475;
  assign n8538 = ~n8415 & ~n8462;
  assign n8539 = ~n8450 & ~n8456;
  assign n8540 = n4913 & n7037;
  assign n8541 = n4920 & ~n10355;
  assign n8542 = n10106 & ~n5987;
  assign n8543 = n4933 & n6492;
  assign n8544 = n4933 & n6490;
  assign n8545 = ~n8542 & ~n10535;
  assign n8546 = ~n8541 & n8545;
  assign n8547 = ~n4913 & n8546;
  assign n8548 = ~n7037 & n8546;
  assign n8549 = ~n8547 & ~n8548;
  assign n8550 = ~n8540 & n8546;
  assign n8551 = ~n9626 & ~n10536;
  assign n8552 = n9626 & n10536;
  assign n8553 = ~n8551 & ~n8552;
  assign n8554 = ~n8539 & n8553;
  assign n8555 = n8539 & ~n8553;
  assign n8556 = ~n8539 & ~n8554;
  assign n8557 = n8553 & ~n8554;
  assign n8558 = ~n8556 & ~n8557;
  assign n8559 = ~n8554 & ~n8555;
  assign n8560 = n4958 & n6016;
  assign n8561 = n4968 & n10226;
  assign n8562 = n10123 & n10210;
  assign n8563 = n4966 & ~n5920;
  assign n8564 = ~n8562 & ~n8563;
  assign n8565 = ~n8561 & n8564;
  assign n8566 = ~n8560 & n8565;
  assign n8567 = ~n1164 & ~n8566;
  assign n8568 = ~n1164 & ~n8567;
  assign n8569 = ~n1164 & n8566;
  assign n8570 = ~n8566 & ~n8567;
  assign n8571 = n1164 & ~n8566;
  assign n8572 = ~n10538 & ~n10539;
  assign n8573 = ~n1164 & ~n4870;
  assign n8574 = ~n1703 & ~n8573;
  assign n8575 = n1703 & n8573;
  assign n8576 = ~n8574 & ~n8575;
  assign n8577 = n8296 & ~n8574;
  assign n8578 = n8296 & ~n8575;
  assign n8579 = ~n8574 & n8578;
  assign n8580 = ~n8575 & n8577;
  assign n8581 = n8296 & ~n10540;
  assign n8582 = n8296 & ~n8576;
  assign n8583 = ~n8296 & ~n8575;
  assign n8584 = ~n8575 & ~n10540;
  assign n8585 = ~n8574 & ~n8583;
  assign n8586 = ~n8574 & n10542;
  assign n8587 = ~n8296 & n8576;
  assign n8588 = ~n10541 & ~n10543;
  assign n8589 = ~n1164 & ~n8296;
  assign n8590 = ~n1164 & ~n4731;
  assign n8591 = ~n10084 & ~n8296;
  assign n8592 = ~n1164 & n8591;
  assign n8593 = ~n10084 & n10544;
  assign n8594 = ~n8444 & ~n10545;
  assign n8595 = ~n8588 & ~n8594;
  assign n8596 = n8588 & n8594;
  assign n8597 = ~n8594 & ~n8595;
  assign n8598 = ~n8588 & ~n8595;
  assign n8599 = ~n8597 & ~n8598;
  assign n8600 = ~n8595 & ~n8596;
  assign n8601 = n8572 & n10546;
  assign n8602 = ~n8572 & ~n10546;
  assign n8603 = ~n10546 & ~n8602;
  assign n8604 = ~n8572 & ~n8602;
  assign n8605 = ~n8603 & ~n8604;
  assign n8606 = ~n8601 & ~n8602;
  assign n8607 = ~n10537 & ~n10547;
  assign n8608 = ~n8557 & n10547;
  assign n8609 = ~n8556 & n8608;
  assign n8610 = ~n8556 & n10547;
  assign n8611 = ~n8557 & n8610;
  assign n8612 = n10537 & n10547;
  assign n8613 = ~n8607 & ~n10548;
  assign n8614 = ~n8538 & n8613;
  assign n8615 = n8538 & ~n8613;
  assign n8616 = ~n8614 & ~n8615;
  assign n8617 = ~n8537 & n8616;
  assign n8618 = n8537 & ~n8616;
  assign n8619 = ~n8617 & ~n8618;
  assign n8620 = n685 & n4641;
  assign n8621 = n5921 & n8620;
  assign n8622 = ~n605 & ~n933;
  assign n8623 = ~n9544 & ~n605;
  assign n8624 = ~n933 & n8623;
  assign n8625 = ~n9544 & ~n933;
  assign n8626 = ~n605 & n8625;
  assign n8627 = ~n9544 & n8622;
  assign n8628 = n551 & n10549;
  assign n8629 = n1467 & n10207;
  assign n8630 = n10207 & n10549;
  assign n8631 = n551 & n1467;
  assign n8632 = n8630 & n8631;
  assign n8633 = n8628 & n8629;
  assign n8634 = n8621 & n10550;
  assign n8635 = n9662 & n8634;
  assign n8636 = n9745 & n10329;
  assign n8637 = n9662 & n4641;
  assign n8638 = n551 & n8637;
  assign n8639 = n685 & n8638;
  assign n8640 = n10207 & n8639;
  assign n8641 = n10329 & n8640;
  assign n8642 = n9745 & n8641;
  assign n8643 = n5921 & n8642;
  assign n8644 = n1467 & n8643;
  assign n8645 = ~n933 & n8644;
  assign n8646 = ~n9544 & n8645;
  assign n8647 = ~n605 & n8646;
  assign n8648 = n8635 & n8636;
  assign n8649 = ~n8619 & n10551;
  assign n8650 = n8619 & ~n10551;
  assign n8651 = ~n8649 & ~n8650;
  assign n8652 = ~n8536 & n8651;
  assign n8653 = n8536 & ~n8651;
  assign n8654 = ~n8652 & ~n8653;
  assign n8655 = ~n8529 & ~n8654;
  assign n8656 = n8529 & n8654;
  assign n8657 = ~n8655 & ~n8656;
  assign n8658 = ~n8530 & n8531;
  assign n8659 = n10350 & ~n8658;
  assign n8660 = n8657 & ~n8659;
  assign n8661 = ~n8657 & n8659;
  assign n8662 = ~n8660 & ~n8661;
  assign n8663 = ~n8650 & ~n8652;
  assign n8664 = ~n8614 & ~n8617;
  assign n8665 = ~n8554 & ~n8607;
  assign n8666 = n4913 & n10386;
  assign n8667 = n10106 & n6492;
  assign n8668 = n10106 & n6490;
  assign n8669 = n4933 & ~n10355;
  assign n8670 = ~n10552 & ~n8669;
  assign n8671 = ~n8666 & n8670;
  assign n8672 = n9626 & ~n8671;
  assign n8673 = ~n9626 & n8671;
  assign n8674 = ~n8672 & ~n8673;
  assign n8675 = n4958 & n5994;
  assign n8676 = n4968 & ~n5987;
  assign n8677 = n10123 & ~n5920;
  assign n8678 = n4966 & n10226;
  assign n8679 = ~n8677 & ~n8678;
  assign n8680 = ~n8676 & n8679;
  assign n8681 = ~n4958 & n8680;
  assign n8682 = ~n5994 & n8680;
  assign n8683 = ~n8681 & ~n8682;
  assign n8684 = ~n8675 & n8680;
  assign n8685 = n1164 & ~n10553;
  assign n8686 = ~n1164 & n10553;
  assign n8687 = ~n8685 & ~n8686;
  assign n8688 = ~n1164 & n10210;
  assign n8689 = ~n10542 & ~n8688;
  assign n8690 = n10542 & n8688;
  assign n8691 = ~n10542 & n8688;
  assign n8692 = n10542 & ~n8688;
  assign n8693 = ~n8691 & ~n8692;
  assign n8694 = ~n8689 & ~n8690;
  assign n8695 = n8687 & ~n10554;
  assign n8696 = ~n8687 & n10554;
  assign n8697 = ~n8695 & ~n8696;
  assign n8698 = ~n8572 & ~n8596;
  assign n8699 = n8572 & ~n8595;
  assign n8700 = ~n8596 & ~n8699;
  assign n8701 = ~n8595 & ~n8602;
  assign n8702 = ~n8595 & ~n8698;
  assign n8703 = n8697 & n10555;
  assign n8704 = ~n8697 & ~n10555;
  assign n8705 = n10555 & ~n8703;
  assign n8706 = n8697 & ~n8703;
  assign n8707 = ~n8705 & ~n8706;
  assign n8708 = ~n8703 & ~n8704;
  assign n8709 = n8674 & ~n10556;
  assign n8710 = ~n8674 & ~n8706;
  assign n8711 = ~n8705 & n8710;
  assign n8712 = ~n8674 & n10556;
  assign n8713 = ~n8709 & ~n10557;
  assign n8714 = ~n8665 & n8713;
  assign n8715 = n8665 & ~n8713;
  assign n8716 = ~n8714 & ~n8715;
  assign n8717 = ~n8664 & n8716;
  assign n8718 = n8664 & ~n8716;
  assign n8719 = ~n8717 & ~n8718;
  assign n8720 = ~n776 & n1546;
  assign n8721 = n1480 & n8720;
  assign n8722 = n9630 & n8721;
  assign n8723 = n9644 & n8722;
  assign n8724 = n10288 & n8723;
  assign n8725 = n1480 & n1546;
  assign n8726 = n9644 & n8725;
  assign n8727 = n10288 & n8726;
  assign n8728 = n9659 & n8727;
  assign n8729 = n9630 & n8728;
  assign n8730 = ~n776 & n8729;
  assign n8731 = n9659 & n8724;
  assign n8732 = ~n8719 & n10558;
  assign n8733 = n8719 & ~n10558;
  assign n8734 = ~n8732 & ~n8733;
  assign n8735 = ~n8663 & n8734;
  assign n8736 = n8663 & ~n8734;
  assign n8737 = ~n8735 & ~n8736;
  assign n8738 = ~n8656 & ~n8737;
  assign n8739 = n8656 & n8737;
  assign n8740 = ~n8738 & ~n8739;
  assign n8741 = ~n8657 & n8658;
  assign n8742 = n10350 & ~n8741;
  assign n8743 = n8740 & ~n8742;
  assign n8744 = ~n8740 & n8742;
  assign n8745 = ~n8743 & ~n8744;
  assign n8746 = ~n8733 & ~n8735;
  assign n8747 = ~n8714 & ~n8717;
  assign n8748 = ~n8703 & ~n8709;
  assign n8749 = ~n8689 & ~n8695;
  assign n8750 = ~n1164 & ~n5920;
  assign n8751 = ~n8688 & n8750;
  assign n8752 = ~n10210 & n8750;
  assign n8753 = n8688 & ~n8750;
  assign n8754 = n5920 & n8688;
  assign n8755 = ~n10559 & ~n10560;
  assign n8756 = ~n8749 & ~n10560;
  assign n8757 = ~n10559 & n8756;
  assign n8758 = ~n8749 & n8755;
  assign n8759 = n8749 & ~n8755;
  assign n8760 = ~n8749 & ~n10561;
  assign n8761 = ~n10560 & ~n10561;
  assign n8762 = ~n10559 & n8761;
  assign n8763 = ~n8760 & ~n8762;
  assign n8764 = ~n10561 & ~n8759;
  assign n8765 = n4958 & n6500;
  assign n8766 = n4968 & n6492;
  assign n8767 = n4968 & n6490;
  assign n8768 = n10123 & n10226;
  assign n8769 = n4966 & ~n5987;
  assign n8770 = ~n8768 & ~n8769;
  assign n8771 = ~n10563 & n8770;
  assign n8772 = ~n8765 & n8771;
  assign n8773 = ~n1164 & ~n8772;
  assign n8774 = ~n1164 & ~n8773;
  assign n8775 = ~n1164 & n8772;
  assign n8776 = ~n8772 & ~n8773;
  assign n8777 = n1164 & ~n8772;
  assign n8778 = ~n10564 & ~n10565;
  assign n8779 = n4913 & ~n10385;
  assign n8780 = ~n10106 & ~n8779;
  assign n8781 = n10106 & ~n10355;
  assign n8782 = n4913 & n7243;
  assign n8783 = ~n8781 & ~n8782;
  assign n8784 = ~n10355 & ~n8780;
  assign n8785 = ~n9626 & ~n10566;
  assign n8786 = n9626 & n10566;
  assign n8787 = n9626 & ~n10566;
  assign n8788 = ~n9626 & n10566;
  assign n8789 = ~n8787 & ~n8788;
  assign n8790 = ~n8785 & ~n8786;
  assign n8791 = ~n8778 & n10567;
  assign n8792 = n8778 & ~n10567;
  assign n8793 = n10567 & ~n8791;
  assign n8794 = ~n8778 & ~n8791;
  assign n8795 = ~n8793 & ~n8794;
  assign n8796 = ~n8791 & ~n8792;
  assign n8797 = ~n10562 & ~n10568;
  assign n8798 = n10562 & n10568;
  assign n8799 = n10562 & ~n10568;
  assign n8800 = ~n10562 & n10568;
  assign n8801 = ~n8799 & ~n8800;
  assign n8802 = ~n8797 & ~n8798;
  assign n8803 = ~n8748 & ~n10569;
  assign n8804 = n8748 & n10569;
  assign n8805 = ~n8803 & ~n8804;
  assign n8806 = ~n8747 & n8805;
  assign n8807 = n8747 & ~n8805;
  assign n8808 = ~n8806 & ~n8807;
  assign n8809 = ~n898 & ~n1108;
  assign n8810 = ~n199 & ~n324;
  assign n8811 = ~n301 & n8810;
  assign n8812 = ~n898 & n8810;
  assign n8813 = ~n301 & n8812;
  assign n8814 = ~n1108 & n8813;
  assign n8815 = ~n324 & ~n1108;
  assign n8816 = ~n199 & ~n898;
  assign n8817 = ~n301 & n8816;
  assign n8818 = n8815 & n8817;
  assign n8819 = ~n301 & ~n898;
  assign n8820 = ~n1108 & n8819;
  assign n8821 = n8810 & n8820;
  assign n8822 = n8809 & n8811;
  assign n8823 = ~n401 & ~n405;
  assign n8824 = n211 & n263;
  assign n8825 = ~n479 & n10571;
  assign n8826 = n4233 & n8825;
  assign n8827 = n1631 & n8826;
  assign n8828 = n10411 & n8827;
  assign n8829 = n10411 & n10570;
  assign n8830 = n8827 & n8829;
  assign n8831 = n10570 & n8828;
  assign n8832 = n10030 & n10572;
  assign n8833 = n4233 & n10570;
  assign n8834 = n1631 & n8833;
  assign n8835 = n10411 & n8834;
  assign n8836 = n9996 & n8835;
  assign n8837 = n10030 & n8836;
  assign n8838 = ~n405 & n8837;
  assign n8839 = ~n401 & n8838;
  assign n8840 = ~n479 & n8839;
  assign n8841 = n9996 & n10572;
  assign n8842 = n10030 & n8841;
  assign n8843 = n9996 & n8832;
  assign n8844 = ~n8808 & n10573;
  assign n8845 = n8808 & ~n10573;
  assign n8846 = ~n8844 & ~n8845;
  assign n8847 = ~n8746 & n8846;
  assign n8848 = n8746 & ~n8846;
  assign n8849 = ~n8847 & ~n8848;
  assign n8850 = ~n8739 & ~n8849;
  assign n8851 = n8739 & n8849;
  assign n8852 = ~n8850 & ~n8851;
  assign n8853 = ~n8740 & n8741;
  assign n8854 = n10350 & ~n8853;
  assign n8855 = n8852 & ~n8854;
  assign n8856 = ~n8852 & n8854;
  assign n8857 = ~n8855 & ~n8856;
  assign n8858 = ~n8845 & ~n8847;
  assign n8859 = ~n8803 & ~n8806;
  assign n8860 = ~n8791 & ~n8797;
  assign n8861 = n4958 & n7037;
  assign n8862 = n4968 & ~n10355;
  assign n8863 = n10123 & ~n5987;
  assign n8864 = n4966 & n6492;
  assign n8865 = n4966 & n6490;
  assign n8866 = ~n8863 & ~n10574;
  assign n8867 = ~n8862 & n8866;
  assign n8868 = ~n8861 & n8867;
  assign n8869 = ~n1164 & ~n8868;
  assign n8870 = ~n8868 & ~n8869;
  assign n8871 = n1164 & ~n8868;
  assign n8872 = ~n1164 & ~n8869;
  assign n8873 = ~n1164 & n8868;
  assign n8874 = ~n10575 & ~n10576;
  assign n8875 = ~n9626 & n8750;
  assign n8876 = n9626 & ~n8750;
  assign n8877 = ~n8875 & ~n8876;
  assign n8878 = ~n1164 & n10226;
  assign n8879 = n8877 & n8878;
  assign n8880 = ~n8877 & ~n8878;
  assign n8881 = ~n8879 & ~n8880;
  assign n8882 = ~n8874 & n8881;
  assign n8883 = n8874 & ~n8881;
  assign n8884 = ~n8874 & ~n8882;
  assign n8885 = ~n8874 & ~n8881;
  assign n8886 = n8881 & ~n8882;
  assign n8887 = n8874 & n8881;
  assign n8888 = ~n10577 & ~n10578;
  assign n8889 = ~n8882 & ~n8883;
  assign n8890 = ~n8761 & ~n10579;
  assign n8891 = n8761 & n10579;
  assign n8892 = ~n8761 & n10579;
  assign n8893 = n8761 & ~n10579;
  assign n8894 = ~n8892 & ~n8893;
  assign n8895 = ~n8890 & ~n8891;
  assign n8896 = ~n8860 & ~n10580;
  assign n8897 = n8860 & n10580;
  assign n8898 = ~n8896 & ~n8897;
  assign n8899 = ~n8859 & n8898;
  assign n8900 = n8859 & ~n8898;
  assign n8901 = ~n8899 & ~n8900;
  assign n8902 = ~n9541 & ~n682;
  assign n8903 = ~n311 & n8902;
  assign n8904 = ~n311 & ~n682;
  assign n8905 = ~n871 & n8904;
  assign n8906 = ~n9541 & n8905;
  assign n8907 = ~n265 & n8906;
  assign n8908 = ~n265 & ~n311;
  assign n8909 = ~n871 & n8902;
  assign n8910 = n8908 & n8909;
  assign n8911 = ~n265 & ~n682;
  assign n8912 = ~n9541 & ~n871;
  assign n8913 = ~n311 & n8912;
  assign n8914 = n8911 & n8913;
  assign n8915 = n1663 & n8903;
  assign n8916 = n385 & n1432;
  assign n8917 = n1972 & n8359;
  assign n8918 = n8916 & n8917;
  assign n8919 = ~n9537 & ~n250;
  assign n8920 = ~n230 & ~n397;
  assign n8921 = n8919 & n8920;
  assign n8922 = n7165 & n8921;
  assign n8923 = ~n230 & ~n250;
  assign n8924 = n385 & n8923;
  assign n8925 = n1432 & n1972;
  assign n8926 = n8924 & n8925;
  assign n8927 = ~n397 & ~n467;
  assign n8928 = ~n9537 & n8927;
  assign n8929 = n10380 & n8928;
  assign n8930 = n8926 & n8929;
  assign n8931 = ~n332 & ~n397;
  assign n8932 = ~n262 & ~n467;
  assign n8933 = n8931 & n8932;
  assign n8934 = n8916 & n8933;
  assign n8935 = ~n230 & n8919;
  assign n8936 = n10380 & n8935;
  assign n8937 = n8934 & n8936;
  assign n8938 = n8918 & n8922;
  assign n8939 = n10581 & n10582;
  assign n8940 = n9752 & n8939;
  assign n8941 = n9986 & n10334;
  assign n8942 = n385 & n10581;
  assign n8943 = n10380 & n8942;
  assign n8944 = n9752 & n8943;
  assign n8945 = n9986 & n8944;
  assign n8946 = n1432 & n8945;
  assign n8947 = n10334 & n8946;
  assign n8948 = ~n262 & n8947;
  assign n8949 = ~n9537 & n8948;
  assign n8950 = ~n467 & n8949;
  assign n8951 = ~n332 & n8950;
  assign n8952 = ~n397 & n8951;
  assign n8953 = ~n230 & n8952;
  assign n8954 = ~n250 & n8953;
  assign n8955 = n8940 & n8941;
  assign n8956 = n8901 & ~n10583;
  assign n8957 = ~n8901 & n10583;
  assign n8958 = ~n8956 & ~n8957;
  assign n8959 = ~n8858 & ~n8957;
  assign n8960 = ~n8956 & n8959;
  assign n8961 = ~n8858 & n8958;
  assign n8962 = n8858 & ~n8958;
  assign n8963 = ~n8858 & ~n10584;
  assign n8964 = ~n8956 & ~n10584;
  assign n8965 = ~n8957 & n8964;
  assign n8966 = ~n8963 & ~n8965;
  assign n8967 = ~n10584 & ~n8962;
  assign n8968 = ~n8851 & n10585;
  assign n8969 = n8851 & ~n10585;
  assign n8970 = ~n8968 & ~n8969;
  assign n8971 = ~n8852 & n8853;
  assign n8972 = n10350 & ~n8971;
  assign n8973 = n8970 & ~n8972;
  assign n8974 = ~n8970 & n8972;
  assign n8975 = ~n8973 & ~n8974;
  assign n8976 = ~n8896 & ~n8899;
  assign n8977 = ~n8882 & ~n8890;
  assign n8978 = n4958 & n10386;
  assign n8979 = n10123 & n6492;
  assign n8980 = n10123 & n6490;
  assign n8981 = n4966 & ~n10355;
  assign n8982 = ~n10586 & ~n8981;
  assign n8983 = ~n4958 & n8982;
  assign n8984 = ~n10386 & n8982;
  assign n8985 = ~n8983 & ~n8984;
  assign n8986 = ~n8978 & n8982;
  assign n8987 = n1164 & ~n10587;
  assign n8988 = ~n1164 & n10587;
  assign n8989 = ~n8987 & ~n8988;
  assign n8990 = ~n1164 & ~n5987;
  assign n8991 = ~n8875 & ~n8879;
  assign n8992 = ~n8990 & ~n8991;
  assign n8993 = n8990 & n8991;
  assign n8994 = ~n8990 & ~n8992;
  assign n8995 = ~n8990 & n8991;
  assign n8996 = ~n8991 & ~n8992;
  assign n8997 = n8990 & ~n8991;
  assign n8998 = ~n10588 & ~n10589;
  assign n8999 = ~n8992 & ~n8993;
  assign n9000 = n8989 & ~n10590;
  assign n9001 = ~n8989 & n10590;
  assign n9002 = ~n9000 & ~n9001;
  assign n9003 = ~n8977 & n9002;
  assign n9004 = n8977 & ~n9002;
  assign n9005 = ~n9003 & ~n9004;
  assign n9006 = ~n8976 & n9005;
  assign n9007 = n8976 & ~n9005;
  assign n9008 = ~n9006 & ~n9007;
  assign n9009 = n716 & n4233;
  assign n9010 = n4432 & n5921;
  assign n9011 = n9009 & n9010;
  assign n9012 = ~n334 & ~n414;
  assign n9013 = ~n513 & n9012;
  assign n9014 = ~n9537 & ~n776;
  assign n9015 = n1036 & n9014;
  assign n9016 = n9013 & n9015;
  assign n9017 = n1036 & n4233;
  assign n9018 = n9010 & n9017;
  assign n9019 = ~n9537 & ~n715;
  assign n9020 = ~n513 & n9019;
  assign n9021 = ~n312 & ~n414;
  assign n9022 = ~n334 & ~n776;
  assign n9023 = n9021 & n9022;
  assign n9024 = ~n9537 & n9022;
  assign n9025 = ~n414 & ~n513;
  assign n9026 = n716 & n9025;
  assign n9027 = n9024 & n9026;
  assign n9028 = n9020 & n9023;
  assign n9029 = n9018 & n10591;
  assign n9030 = n9011 & n9016;
  assign n9031 = n9692 & n10592;
  assign n9032 = n9703 & n9833;
  assign n9033 = n9031 & n9032;
  assign n9034 = n4233 & n4432;
  assign n9035 = n1036 & n9034;
  assign n9036 = n9703 & n9035;
  assign n9037 = n9982 & n9036;
  assign n9038 = n9833 & n9037;
  assign n9039 = n9692 & n9038;
  assign n9040 = n5921 & n9039;
  assign n9041 = ~n414 & n9040;
  assign n9042 = ~n334 & n9041;
  assign n9043 = ~n312 & n9042;
  assign n9044 = ~n9537 & n9043;
  assign n9045 = ~n715 & n9044;
  assign n9046 = ~n776 & n9045;
  assign n9047 = ~n513 & n9046;
  assign n9048 = n9982 & n9033;
  assign n9049 = ~n9008 & n10593;
  assign n9050 = n9008 & ~n10593;
  assign n9051 = ~n9049 & ~n9050;
  assign n9052 = ~n8964 & n9051;
  assign n9053 = n8964 & ~n9051;
  assign n9054 = ~n9052 & ~n9053;
  assign n9055 = ~n8969 & ~n9054;
  assign n9056 = n8969 & n9054;
  assign n9057 = ~n9055 & ~n9056;
  assign n9058 = ~n8970 & n8971;
  assign n9059 = n10350 & ~n9058;
  assign n9060 = n9057 & ~n9059;
  assign n9061 = ~n9057 & n9059;
  assign n9062 = ~n9060 & ~n9061;
  assign n9063 = ~n9050 & ~n9052;
  assign n9064 = ~n8992 & ~n9000;
  assign n9065 = n4958 & ~n10385;
  assign n9066 = ~n10123 & ~n9065;
  assign n9067 = n10123 & ~n10355;
  assign n9068 = n4958 & n7243;
  assign n9069 = ~n9067 & ~n9068;
  assign n9070 = ~n10355 & ~n9066;
  assign n9071 = ~n1164 & ~n10594;
  assign n9072 = n6497 & n9071;
  assign n9073 = ~n1164 & ~n6497;
  assign n9074 = n10594 & ~n9073;
  assign n9075 = ~n10594 & ~n9071;
  assign n9076 = n1164 & ~n10594;
  assign n9077 = ~n1164 & ~n9071;
  assign n9078 = ~n1164 & n10594;
  assign n9079 = ~n10595 & ~n10596;
  assign n9080 = ~n1164 & n6497;
  assign n9081 = ~n9079 & ~n9080;
  assign n9082 = ~n9071 & ~n9074;
  assign n9083 = ~n9079 & ~n10597;
  assign n9084 = n6497 & n10596;
  assign n9085 = n9079 & ~n9080;
  assign n9086 = ~n9080 & ~n10597;
  assign n9087 = ~n10598 & ~n10599;
  assign n9088 = ~n9072 & ~n10597;
  assign n9089 = n9064 & n10600;
  assign n9090 = ~n9064 & ~n10600;
  assign n9091 = ~n9089 & ~n9090;
  assign n9092 = ~n9003 & ~n9006;
  assign n9093 = ~n9091 & n9092;
  assign n9094 = n9091 & ~n9092;
  assign n9095 = ~n9093 & ~n9094;
  assign n9096 = ~n225 & ~n714;
  assign n9097 = ~n225 & ~n573;
  assign n9098 = ~n714 & n9097;
  assign n9099 = ~n573 & ~n714;
  assign n9100 = ~n225 & n9099;
  assign n9101 = ~n573 & n9096;
  assign n9102 = ~n225 & n9756;
  assign n9103 = ~n714 & n9102;
  assign n9104 = ~n573 & n9103;
  assign n9105 = n9756 & n10601;
  assign n9106 = ~n241 & ~n249;
  assign n9107 = ~n190 & ~n312;
  assign n9108 = ~n190 & ~n249;
  assign n9109 = ~n241 & ~n312;
  assign n9110 = n9108 & n9109;
  assign n9111 = n9106 & n9107;
  assign n9112 = n1192 & n1482;
  assign n9113 = n6795 & n9112;
  assign n9114 = n6795 & n9108;
  assign n9115 = n1192 & n9109;
  assign n9116 = n1482 & n9115;
  assign n9117 = n9114 & n9116;
  assign n9118 = n10603 & n9113;
  assign n9119 = n10570 & n10604;
  assign n9120 = n9753 & n9119;
  assign n9121 = n10034 & n9120;
  assign n9122 = n1482 & n10602;
  assign n9123 = n1192 & n9122;
  assign n9124 = n10570 & n9123;
  assign n9125 = n10034 & n9124;
  assign n9126 = n9753 & n9125;
  assign n9127 = ~n312 & n9126;
  assign n9128 = ~n249 & n9127;
  assign n9129 = ~n241 & n9128;
  assign n9130 = ~n190 & n9129;
  assign n9131 = ~n513 & n9130;
  assign n9132 = ~n552 & n9131;
  assign n9133 = n10602 & n9121;
  assign n9134 = n9095 & ~n10605;
  assign n9135 = ~n9095 & n10605;
  assign n9136 = ~n9134 & ~n9135;
  assign n9137 = ~n9063 & ~n9135;
  assign n9138 = ~n9134 & n9137;
  assign n9139 = ~n9063 & n9136;
  assign n9140 = n9063 & ~n9136;
  assign n9141 = ~n9063 & ~n10606;
  assign n9142 = ~n9134 & ~n10606;
  assign n9143 = ~n9135 & n9142;
  assign n9144 = ~n9141 & ~n9143;
  assign n9145 = ~n10606 & ~n9140;
  assign n9146 = ~n9056 & n10607;
  assign n9147 = n9056 & ~n10607;
  assign n9148 = ~n9146 & ~n9147;
  assign n9149 = ~n9057 & n9058;
  assign n9150 = n10350 & ~n9149;
  assign n9151 = n9148 & ~n9150;
  assign n9152 = ~n9148 & n9150;
  assign n9153 = ~n9151 & ~n9152;
  assign n9154 = ~n9562 & ~n781;
  assign n9155 = ~n9586 & ~n781;
  assign n9156 = ~n9562 & n9155;
  assign n9157 = ~n9562 & ~n9586;
  assign n9158 = ~n781 & n9157;
  assign n9159 = ~n9586 & n9154;
  assign n9160 = n550 & n1248;
  assign n9161 = n10608 & n9160;
  assign n9162 = n9998 & n9161;
  assign n9163 = n10312 & n10581;
  assign n9164 = n9162 & n9163;
  assign n9165 = n10332 & n9164;
  assign n9166 = n1248 & n10012;
  assign n9167 = n9998 & n9166;
  assign n9168 = n10581 & n9167;
  assign n9169 = n10312 & n9168;
  assign n9170 = n550 & n9169;
  assign n9171 = n10332 & n9170;
  assign n9172 = ~n9562 & n9171;
  assign n9173 = ~n9586 & n9172;
  assign n9174 = ~n781 & n9173;
  assign n9175 = n10012 & n9165;
  assign n9176 = ~n1164 & n6492;
  assign n9177 = ~n1164 & ~n10290;
  assign n9178 = n6492 & ~n8990;
  assign n9179 = ~n1164 & n9178;
  assign n9180 = ~n8990 & n10610;
  assign n9181 = n5987 & n10610;
  assign n9182 = ~n10597 & ~n10611;
  assign n9183 = ~n9090 & ~n9094;
  assign n9184 = ~n5987 & n10355;
  assign n9185 = n5987 & ~n10355;
  assign n9186 = ~n10355 & ~n8990;
  assign n9187 = ~n1164 & ~n9186;
  assign n9188 = ~n1164 & ~n9185;
  assign n9189 = n10355 & ~n8990;
  assign n9190 = ~n10355 & n8990;
  assign n9191 = n10355 & n8990;
  assign n9192 = ~n9186 & ~n9191;
  assign n9193 = ~n9189 & ~n9190;
  assign n9194 = ~n1164 & n10613;
  assign n9195 = n10612 & ~n9191;
  assign n9196 = ~n9184 & n10612;
  assign n9197 = n9183 & ~n10614;
  assign n9198 = ~n9183 & n10614;
  assign n9199 = ~n9197 & ~n9198;
  assign n9200 = n9182 & n9199;
  assign n9201 = ~n9182 & ~n9199;
  assign n9202 = n9182 & ~n9183;
  assign n9203 = ~n9182 & n9183;
  assign n9204 = ~n9202 & ~n9203;
  assign n9205 = ~n10614 & n9204;
  assign n9206 = n10614 & ~n9204;
  assign n9207 = ~n9205 & ~n9206;
  assign n9208 = ~n9200 & ~n9201;
  assign n9209 = ~n10609 & ~n10615;
  assign n9210 = n10609 & n10615;
  assign n9211 = ~n9209 & ~n9210;
  assign n9212 = n9142 & ~n9211;
  assign n9213 = ~n9142 & ~n9210;
  assign n9214 = ~n9209 & n9213;
  assign n9215 = ~n9142 & ~n9209;
  assign n9216 = ~n9210 & n9215;
  assign n9217 = ~n9142 & n9211;
  assign n9218 = ~n9142 & ~n10616;
  assign n9219 = ~n9142 & ~n9211;
  assign n9220 = n9142 & ~n9209;
  assign n9221 = ~n9209 & ~n10616;
  assign n9222 = ~n9210 & ~n9220;
  assign n9223 = ~n9210 & n10618;
  assign n9224 = n9142 & n9211;
  assign n9225 = ~n10617 & ~n10619;
  assign n9226 = ~n9212 & ~n10616;
  assign n9227 = ~n9147 & n10620;
  assign n9228 = n9147 & ~n10620;
  assign n9229 = ~n9227 & ~n9228;
  assign n9230 = ~n9148 & n9149;
  assign n9231 = n10350 & ~n9230;
  assign n9232 = n9229 & ~n9231;
  assign n9233 = ~n9229 & n9231;
  assign n9234 = ~n9232 & ~n9233;
  assign n9235 = ~n9229 & n9230;
  assign n9236 = n10350 & ~n9235;
  assign n9237 = ~n533 & ~n898;
  assign n9238 = n4641 & n9237;
  assign n9239 = n1432 & n1558;
  assign n9240 = n9238 & n9239;
  assign n9241 = ~n480 & ~n618;
  assign n9242 = ~n405 & n9241;
  assign n9243 = n9582 & n9242;
  assign n9244 = ~n405 & ~n533;
  assign n9245 = n1558 & n9244;
  assign n9246 = n1432 & n4641;
  assign n9247 = n9245 & n9246;
  assign n9248 = ~n898 & n9241;
  assign n9249 = n9582 & n9248;
  assign n9250 = n9247 & n9249;
  assign n9251 = ~n405 & ~n898;
  assign n9252 = n4641 & n9251;
  assign n9253 = n9239 & n9252;
  assign n9254 = ~n480 & ~n533;
  assign n9255 = ~n618 & n9254;
  assign n9256 = n9582 & n9255;
  assign n9257 = n9253 & n9256;
  assign n9258 = n9240 & n9243;
  assign n9259 = n9565 & n10621;
  assign n9260 = n9563 & n9259;
  assign n9261 = n9565 & n9582;
  assign n9262 = n1558 & n9261;
  assign n9263 = n4641 & n9262;
  assign n9264 = n10206 & n9263;
  assign n9265 = n9563 & n9264;
  assign n9266 = n1432 & n9265;
  assign n9267 = ~n405 & n9266;
  assign n9268 = ~n898 & n9267;
  assign n9269 = ~n533 & n9268;
  assign n9270 = ~n618 & n9269;
  assign n9271 = ~n480 & n9270;
  assign n9272 = n10206 & n9260;
  assign n9273 = ~n10618 & ~n10622;
  assign n9274 = n10618 & n10622;
  assign n9275 = ~n9273 & ~n9274;
  assign n9276 = n9228 & n9275;
  assign n9277 = ~n9228 & ~n9275;
  assign n9278 = ~n9276 & ~n9277;
  assign n9279 = ~n9228 & n9275;
  assign n9280 = n9228 & ~n9275;
  assign n9281 = ~n9279 & ~n9280;
  assign n9282 = n9236 & ~n9281;
  assign n9283 = n9236 & n9278;
  assign n9284 = ~n9236 & n9281;
  assign n9285 = ~n9236 & ~n9278;
  assign po17  = ~n10623 & ~n10624;
  assign n9287 = n9235 & ~n9278;
  assign n9288 = n10350 & ~n9287;
  assign n9289 = ~n676 & ~n898;
  assign n9290 = ~n9555 & ~n334;
  assign n9291 = ~n351 & n9290;
  assign n9292 = ~n334 & ~n351;
  assign n9293 = ~n9555 & ~n676;
  assign n9294 = ~n898 & n9293;
  assign n9295 = n9292 & n9294;
  assign n9296 = ~n334 & ~n898;
  assign n9297 = ~n9555 & ~n351;
  assign n9298 = ~n676 & n9297;
  assign n9299 = n9296 & n9298;
  assign n9300 = n9289 & n9291;
  assign n9301 = n9657 & n9688;
  assign n9302 = n10625 & n9301;
  assign n9303 = n9750 & n9983;
  assign n9304 = n9302 & n9303;
  assign n9305 = n9759 & n9304;
  assign n9306 = n9568 & n10324;
  assign n9307 = n9568 & n9983;
  assign n9308 = n9657 & n9307;
  assign n9309 = n9759 & n9308;
  assign n9310 = n9750 & n9309;
  assign n9311 = n9688 & n9310;
  assign n9312 = n10324 & n9311;
  assign n9313 = ~n334 & n9312;
  assign n9314 = ~n9555 & n9313;
  assign n9315 = ~n898 & n9314;
  assign n9316 = ~n676 & n9315;
  assign n9317 = ~n351 & n9316;
  assign n9318 = n10324 & n9305;
  assign n9319 = n9568 & n9318;
  assign n9320 = n9305 & n9306;
  assign n9321 = n9273 & ~n10626;
  assign n9322 = ~n9273 & n10626;
  assign n9323 = ~n9321 & ~n9322;
  assign n9324 = ~n9276 & ~n9323;
  assign n9325 = n9276 & ~n9322;
  assign n9326 = ~n9273 & ~n9276;
  assign n9327 = n10626 & ~n9326;
  assign n9328 = ~n10626 & n9326;
  assign n9329 = ~n9327 & ~n9328;
  assign n9330 = ~n9324 & ~n9325;
  assign n9331 = n9235 & n9281;
  assign n9332 = n10350 & ~n9331;
  assign n9333 = n10627 & n9332;
  assign n9334 = n9288 & n10627;
  assign n9335 = ~n10627 & ~n9332;
  assign n9336 = ~n9288 & ~n10627;
  assign n9337 = ~n10628 & ~n10629;
  assign n9338 = ~n195 & ~n404;
  assign n9339 = n1172 & n9338;
  assign n9340 = n5716 & n9339;
  assign n9341 = ~n9564 & ~n402;
  assign n9342 = ~n995 & n9341;
  assign n9343 = n10471 & n9342;
  assign n9344 = n5716 & n9341;
  assign n9345 = n1172 & n9344;
  assign n9346 = ~n995 & n9338;
  assign n9347 = n10471 & n9346;
  assign n9348 = n9345 & n9347;
  assign n9349 = ~n402 & ~n404;
  assign n9350 = ~n9564 & ~n534;
  assign n9351 = n9349 & n9350;
  assign n9352 = n1172 & n9351;
  assign n9353 = ~n195 & ~n9562;
  assign n9354 = ~n995 & n9353;
  assign n9355 = n10471 & n9354;
  assign n9356 = n9352 & n9355;
  assign n9357 = n9340 & n9343;
  assign n9358 = n10097 & n10630;
  assign n9359 = n9719 & n9358;
  assign n9360 = n10471 & n10602;
  assign n9361 = n1172 & n9360;
  assign n9362 = n10097 & n9361;
  assign n9363 = n9719 & n9362;
  assign n9364 = ~n402 & n9363;
  assign n9365 = ~n9564 & n9364;
  assign n9366 = ~n9562 & n9365;
  assign n9367 = ~n404 & n9366;
  assign n9368 = ~n995 & n9367;
  assign n9369 = ~n195 & n9368;
  assign n9370 = ~n534 & n9369;
  assign n9371 = n10602 & n9359;
  assign n9372 = ~n9321 & n10631;
  assign n9373 = n9321 & ~n10631;
  assign n9374 = ~n9372 & ~n9373;
  assign n9375 = n9276 & ~n10626;
  assign n9376 = ~n9374 & ~n9375;
  assign n9377 = n9374 & n9375;
  assign n9378 = ~n9376 & ~n9377;
  assign n9379 = n9287 & n10627;
  assign n9380 = n10350 & ~n9379;
  assign n9381 = ~n9325 & ~n9374;
  assign n9382 = n9325 & n9374;
  assign n9383 = ~n9381 & ~n9382;
  assign n9384 = n10627 & n9331;
  assign n9385 = n10350 & ~n9384;
  assign n9386 = n9383 & ~n9385;
  assign n9387 = n9378 & ~n9380;
  assign n9388 = ~n9383 & n9385;
  assign n9389 = ~n9378 & n9380;
  assign n9390 = ~n10632 & ~n10633;
  assign n9391 = ~n9378 & n9379;
  assign n9392 = n10350 & ~n9391;
  assign n9393 = ~n226 & ~n352;
  assign n9394 = n934 & n9393;
  assign n9395 = n8213 & n9394;
  assign n9396 = n992 & n10470;
  assign n9397 = n992 & n9395;
  assign n9398 = n10470 & n9397;
  assign n9399 = n991 & n6698;
  assign n9400 = n8213 & n9399;
  assign n9401 = ~n352 & n934;
  assign n9402 = n10470 & n9401;
  assign n9403 = n9400 & n9402;
  assign n9404 = n991 & n10470;
  assign n9405 = ~n226 & ~n682;
  assign n9406 = ~n175 & ~n990;
  assign n9407 = n9405 & n9406;
  assign n9408 = n9401 & n9407;
  assign n9409 = n9404 & n9408;
  assign n9410 = n9395 & n9396;
  assign n9411 = n9647 & n10634;
  assign n9412 = n9695 & n9411;
  assign n9413 = n826 & n991;
  assign n9414 = n9695 & n9413;
  assign n9415 = n9647 & n9414;
  assign n9416 = n10519 & n9415;
  assign n9417 = n4024 & n9416;
  assign n9418 = ~n682 & n9417;
  assign n9419 = ~n9555 & n9418;
  assign n9420 = ~n933 & n9419;
  assign n9421 = ~n175 & n9420;
  assign n9422 = ~n990 & n9421;
  assign n9423 = ~n226 & n9422;
  assign n9424 = ~n352 & n9423;
  assign n9425 = n10519 & n9412;
  assign n9426 = n9373 & ~n10635;
  assign n9427 = ~n9373 & n10635;
  assign n9428 = ~n9426 & ~n9427;
  assign n9429 = ~n9382 & ~n9428;
  assign n9430 = n9382 & ~n9427;
  assign n9431 = ~n9373 & ~n9377;
  assign n9432 = n10635 & ~n9431;
  assign n9433 = ~n10635 & n9431;
  assign n9434 = ~n9432 & ~n9433;
  assign n9435 = ~n9429 & ~n9430;
  assign n9436 = ~n9383 & n9384;
  assign n9437 = n10350 & ~n9436;
  assign n9438 = n10636 & n9437;
  assign n9439 = n9392 & n10636;
  assign n9440 = ~n10636 & ~n9437;
  assign n9441 = ~n9392 & ~n10636;
  assign n9442 = ~n10637 & ~n10638;
  assign n9443 = ~n168 & n9638;
  assign n9444 = n10229 & n9443;
  assign n9445 = n9638 & n10229;
  assign n9446 = n9624 & n9445;
  assign n9447 = ~n9537 & n9446;
  assign n9448 = ~n9541 & n9447;
  assign n9449 = n9624 & n9444;
  assign n9450 = ~n9426 & n10639;
  assign n9451 = n9426 & ~n10639;
  assign n9452 = ~n9450 & ~n9451;
  assign n9453 = n9377 & ~n10635;
  assign n9454 = ~n9452 & ~n9453;
  assign n9455 = n9452 & n9453;
  assign n9456 = ~n9454 & ~n9455;
  assign n9457 = n9391 & n10636;
  assign n9458 = n10636 & n9436;
  assign n9459 = n10350 & ~n9458;
  assign n9460 = n10350 & ~n9457;
  assign n9461 = ~n9430 & ~n9452;
  assign n9462 = n9430 & n9452;
  assign n9463 = ~n9461 & ~n9462;
  assign n9464 = ~n10640 & n9463;
  assign n9465 = n9456 & ~n10640;
  assign n9466 = n10640 & ~n9463;
  assign n9467 = ~n9456 & n10640;
  assign n9468 = ~n10641 & ~n10642;
  assign n9469 = ~n9456 & n9457;
  assign n9470 = n10350 & ~n9469;
  assign n9471 = n9624 & n9643;
  assign n9472 = ~n9451 & ~n9455;
  assign n9473 = ~n9471 & ~n9472;
  assign n9474 = n9471 & n9472;
  assign n9475 = ~n9473 & ~n9474;
  assign n9476 = n9471 & ~n9472;
  assign n9477 = ~n9471 & n9472;
  assign n9478 = ~n9476 & ~n9477;
  assign n9479 = n9470 & n9478;
  assign n9480 = n9451 & ~n9471;
  assign n9481 = ~n9451 & n9471;
  assign n9482 = ~n9480 & ~n9481;
  assign n9483 = ~n9462 & ~n9482;
  assign n9484 = n9462 & ~n9481;
  assign n9485 = ~n9483 & ~n9484;
  assign n9486 = n9458 & ~n9463;
  assign n9487 = n10350 & ~n9486;
  assign n9488 = ~n9485 & n9487;
  assign n9489 = n9470 & ~n9475;
  assign n9490 = ~n9470 & ~n9478;
  assign n9491 = n9485 & ~n9487;
  assign n9492 = ~n9470 & n9475;
  assign n9493 = ~n10643 & ~n10644;
  assign n9494 = n9469 & ~n9475;
  assign n9495 = n10350 & ~n9473;
  assign n9496 = ~n9494 & n9495;
  assign n9497 = ~n9470 & n9473;
  assign n9498 = ~pi22  & n134;
  assign n9499 = n120 & n129;
  assign n9500 = ~n9497 & ~n10645;
  assign n9501 = ~n9480 & ~n9484;
  assign n9502 = ~n9485 & n9486;
  assign n9503 = n10350 & ~n9502;
  assign n9504 = n9501 & n9503;
  assign n9505 = ~n9501 & ~n9503;
  assign n9506 = ~n9504 & ~n9505;
  assign n9507 = ~n10645 & n9506;
  assign n9508 = n9469 & n9478;
  assign n9509 = n10350 & ~n9508;
  assign n9510 = ~n9473 & n9509;
  assign n9511 = n9473 & ~n9509;
  assign n9512 = ~n10645 & ~n9511;
  assign n9513 = ~n9510 & n9512;
  assign n9514 = ~n10645 & ~n9505;
  assign n9515 = ~n9504 & n9514;
  assign n9516 = ~n9496 & n9500;
  assign n9517 = n9469 & n9473;
  assign n9518 = ~n10645 & ~n9517;
  assign n9519 = ~n9501 & n9502;
  assign n9520 = n9502 & ~n9519;
  assign n9521 = ~n10645 & n9520;
  assign n9522 = n9508 & n9518;
  assign n9523 = ~n10645 & ~n9519;
  assign n9524 = n9502 & n9523;
  assign n9525 = n9494 & n9518;
  assign po24  = n10350 & ~n10647;
  assign n9527 = n52 | n53;
  assign n9528 = n61 | ~n62;
  assign n9529 = n68 | ~n69;
  assign n9530 = n78 | ~n79;
  assign n9531 = n88 | ~n89;
  assign n9532 = ~n113 | n106 | n112;
  assign n9533 = n123 | n124;
  assign n9534 = ~n140 | n131 | n139;
  assign n9535 = n137 | n138;
  assign n9536 = n160 | ~n161;
  assign n9537 = n169 | n170;
  assign n9538 = n187 | n183 | n186;
  assign n9539 = n209 | n210;
  assign n9540 = n222 | n223;
  assign n9541 = n228 | n229;
  assign n9542 = n234 | n235;
  assign n9543 = n239 | n240;
  assign n9544 = n246 | n247;
  assign n9545 = n253 | n254;
  assign n9546 = n256 | n257;
  assign n9547 = n276 | n271 | n275;
  assign n9548 = n273 | n274;
  assign n9549 = n282 | n279 | n281;
  assign n9550 = n286 | n287;
  assign n9551 = n288 | n289;
  assign n9552 = n291 | n292;
  assign n9553 = n303 | n304;
  assign n9554 = n310 | n307 | n309;
  assign n9555 = n314 | n315;
  assign n9556 = n321 | n318 | n320;
  assign n9557 = n350 | n343 | n349;
  assign n9558 = n346 | n347;
  assign n9559 = n355 | n356;
  assign n9560 = n367 | n359 | n366;
  assign n9561 = n360 | n361;
  assign n9562 = n362 | n363;
  assign n9563 = n379 | n374 | n378;
  assign n9564 = n387 | n388;
  assign n9565 = n392 | n393;
  assign n9566 = n422 | n413 | n421;
  assign n9567 = n429 | n430;
  assign n9568 = n435 | n436;
  assign n9569 = n448 | n445 | n447;
  assign n9570 = n449 | n450;
  assign n9571 = n458 | n460 | n464 | n465;
  assign n9572 = n474 | n475;
  assign n9573 = n483 | n484;
  assign n9574 = n500 | n492 | n499;
  assign n9575 = n508 | n509;
  assign n9576 = n522 | n526 | n531 | n532;
  assign n9577 = n542 | n543;
  assign n9578 = n548 | n549;
  assign n9579 = n561 | n558 | n560;
  assign n9580 = n571 | n572;
  assign n9581 = n580 | n577 | n579;
  assign n9582 = n589 | n586 | n588;
  assign n9583 = n590 | ~n591;
  assign n9584 = n598 | n595 | n597;
  assign n9585 = n601 | n602;
  assign n9586 = n608 | n609;
  assign n9587 = n616 | n617;
  assign n9588 = n636 | n639 | n644 | n645;
  assign n9589 = n657 | n658;
  assign n9590 = n673 | n670 | n672;
  assign n9591 = n680 | n681;
  assign n9592 = n690 | n691;
  assign n9593 = n700 | n701;
  assign n9594 = n704 | n705;
  assign n9595 = n711 | n712;
  assign n9596 = n718 | n719;
  assign n9597 = n723 | n724;
  assign n9598 = n728 | n729;
  assign n9599 = n738 | n734 | n737;
  assign n9600 = n745 | n742 | n744;
  assign n9601 = n751 | n752;
  assign n9602 = n766 | n763 | n765;
  assign n9603 = n768 | n769;
  assign n9604 = n784 | n785;
  assign n9605 = n797 | n793 | n796;
  assign n9606 = n801 | n802;
  assign n9607 = n804 | n805;
  assign n9608 = n818 | n819;
  assign n9609 = n824 | n825;
  assign n9610 = n830 | n833 | n836 | n837;
  assign n9611 = n840 | n841;
  assign n9612 = n844 | n845;
  assign n9613 = n849 | n852 | n855 | n856;
  assign n9614 = n864 | n861 | n863;
  assign n9615 = n869 | n870;
  assign n9616 = n884 | n878 | n883;
  assign n9617 = n896 | n893 | n895;
  assign n9618 = n906 | n907;
  assign n9619 = n915 | n916;
  assign n9620 = n920 | n924 | n931 | n932;
  assign n9621 = n937 | n938;
  assign n9622 = n948 | n943 | n947;
  assign n9623 = n952 | ~n953;
  assign n9624 = n963 | n964;
  assign n9625 = n970 | ~n971;
  assign n9626 = n988 | ~n989;
  assign n9627 = n999 | n1000;
  assign n9628 = n1005 | n1006;
  assign n9629 = n1007 | n1008;
  assign n9630 = n1013 | n1014;
  assign n9631 = n1018 | n1019;
  assign n9632 = n1021 | n1025 | n1027 | n1028;
  assign n9633 = n1034 | n1035;
  assign n9634 = n1044 | n1041 | n1043;
  assign n9635 = n1048 | n1049;
  assign n9636 = n1057 | n1058;
  assign n9637 = n1063 | n1064;
  assign n9638 = n1068 | n1069;
  assign n9639 = n1082 | n1079 | n1081;
  assign n9640 = n1086 | n1087;
  assign n9641 = n1090 | n1091;
  assign n9642 = n1100 | n1101;
  assign n9643 = n1106 | n1107;
  assign n9644 = n1114 | n1117 | n1122 | n1123;
  assign n9645 = n1120 | n1121;
  assign n9646 = n1126 | n1127;
  assign n9647 = n1130 | n1131;
  assign n9648 = n1134 | n1135;
  assign n9649 = n1140 | ~n1141;
  assign n9650 = n1153 | n1154;
  assign n9651 = n1157 | n1158;
  assign n9652 = n1162 | n1163;
  assign n9653 = n1169 | n1170;
  assign n9654 = n1175 | n1176;
  assign n9655 = n1189 | n1182 | n1188;
  assign n9656 = n1198 | n1199;
  assign n9657 = n1205 | n1202 | n1204;
  assign n9658 = n1209 | n1210;
  assign n9659 = n1221 | n1222;
  assign n9660 = n1228 | n1229;
  assign n9661 = n1235 | n1236;
  assign n9662 = n1239 | n1240;
  assign n9663 = n1245 | n1246;
  assign n9664 = n1253 | n1254;
  assign n9665 = n1265 | n1266;
  assign n9666 = n1277 | n1278;
  assign n9667 = n1283 | ~n1284;
  assign n9668 = n1286 | n1287;
  assign n9669 = n1290 | n1291;
  assign n9670 = n1298 | ~n1299;
  assign n9671 = n1301 | n1302;
  assign n9672 = n1308 | n1309;
  assign n9673 = n1314 | ~n1315;
  assign n9674 = n1317 | n1318;
  assign n9675 = n1320 | ~n1321;
  assign n9676 = n1324 | n1325;
  assign n9677 = n1338 | n1339;
  assign n9678 = n1350 | ~n1351;
  assign n9679 = n1362 | n1363;
  assign n9680 = n1366 | n1367;
  assign n9681 = n1372 | n1373;
  assign n9682 = n1374 | n1375;
  assign n9683 = n1376 | ~n1377;
  assign n9684 = n1386 | n1387;
  assign n9685 = n1390 | n1391;
  assign n9686 = n1408 | ~n1409;
  assign n9687 = n1414 | n1415;
  assign n9688 = n1423 | n1419 | n1422;
  assign n9689 = n1426 | n1427;
  assign n9690 = n1430 | n1431;
  assign n9691 = n1435 | n1436;
  assign n9692 = n1439 | n1440;
  assign n9693 = n1443 | n1444;
  assign n9694 = n1454 | n1455;
  assign n9695 = n1462 | n1463;
  assign n9696 = n1464 | n1465;
  assign n9697 = n1470 | n1471;
  assign n9698 = n1474 | n1475;
  assign n9699 = n1486 | n1487;
  assign n9700 = n1492 | n1493;
  assign n9701 = n1496 | n1497;
  assign n9702 = n1507 | n1501 | n1506;
  assign n9703 = n1513 | n1514;
  assign n9704 = n1524 | n1525;
  assign n9705 = n1528 | n1529;
  assign n9706 = n1534 | n1535;
  assign n9707 = n1540 | n1537 | n1539;
  assign n9708 = n1544 | n1545;
  assign n9709 = n1550 | n1551;
  assign n9710 = n1557 | n1554 | n1556;
  assign n9711 = n1562 | n1563;
  assign n9712 = n1568 | n1569;
  assign n9713 = n1581 | n1577 | n1580;
  assign n9714 = n1584 | n1585;
  assign n9715 = n1594 | n1595;
  assign n9716 = n1600 | n1601;
  assign n9717 = n1605 | n1606;
  assign n9718 = n1609 | n1610;
  assign n9719 = n1622 | n1623;
  assign n9720 = n1629 | n1626 | n1628;
  assign n9721 = n1634 | n1635;
  assign n9722 = n1646 | n1650 | n1656 | n1657;
  assign n9723 = n1669 | n1674 | n1678 | n1679;
  assign n9724 = n1693 | n1694;
  assign n9725 = n1706 | n1707;
  assign n9726 = n1713 | n1714;
  assign n9727 = n1717 | n1718;
  assign n9728 = n1721 | n1722;
  assign n9729 = n1734 | n1730 | n1733;
  assign n9730 = n1742 | n1743;
  assign n9731 = n1748 | ~n1749;
  assign n9732 = n1754 | n1755;
  assign n9733 = n1758 | n1759;
  assign n9734 = n1765 | ~n1766;
  assign n9735 = n1779 | n1780;
  assign n9736 = n1781 | n1782;
  assign n9737 = n1783 | ~n1784;
  assign n9738 = n1790 | n1791;
  assign n9739 = n1794 | n1795;
  assign n9740 = n1803 | n1804;
  assign n9741 = n1811 | n1812;
  assign n9742 = n1815 | n1816;
  assign n9743 = n1821 | n1822;
  assign n9744 = n1827 | n1828;
  assign n9745 = n1836 | n1837;
  assign n9746 = n1855 | n1850 | n1854;
  assign n9747 = n1863 | n1864;
  assign n9748 = n1865 | n1866;
  assign n9749 = n1872 | n1873;
  assign n9750 = n1878 | n1875 | n1877;
  assign n9751 = n1882 | n1883;
  assign n9752 = n1911 | n1898 | n1905 | n1917 | n1918;
  assign n9753 = n1930 | n1936 | n1942 | n1943;
  assign n9754 = n1956 | n1957;
  assign n9755 = n1971 | n1968 | n1970;
  assign n9756 = n2005 | n1988 | n1997 | n2015 | n2016;
  assign n9757 = n2021 | n2022;
  assign n9758 = n2028 | n2029;
  assign n9759 = n2038 | n2033 | n2037;
  assign n9760 = n2062 | n2052 | n2061;
  assign n9761 = n2072 | n2073;
  assign n9762 = n2086 | n2083 | n2085;
  assign n9763 = n2089 | n2090;
  assign n9764 = n2102 | n2097 | n2101;
  assign n9765 = n2099 | n2100;
  assign n9766 = n2105 | n2106;
  assign n9767 = n2122 | n2119 | n2121;
  assign n9768 = n2125 | n2126;
  assign n9769 = n2136 | n2134 | n2135;
  assign n9770 = n2140 | n2141;
  assign n9771 = n2147 | ~n2148;
  assign n9772 = n2150 | n2151;
  assign n9773 = n2153 | ~n2154;
  assign n9774 = n2157 | n2158;
  assign n9775 = n2174 | n2170 | n2173;
  assign n9776 = n2180 | n2181;
  assign n9777 = n2183 | ~n2184;
  assign n9778 = n2186 | n2187;
  assign n9779 = n2188 | n2189;
  assign n9780 = n2190 | ~n2191;
  assign n9781 = n2202 | ~n2203;
  assign n9782 = n2212 | ~n2213;
  assign n9783 = n2218 | n2219;
  assign n9784 = n2222 | n2223;
  assign n9785 = n2231 | n2232;
  assign n9786 = n2237 | ~n2238;
  assign n9787 = n2239 | n2240;
  assign n9788 = n2249 | n2250;
  assign n9789 = n2261 | ~n2262;
  assign n9790 = n2266 | n2267;
  assign n9791 = n2268 | n2269;
  assign n9792 = n2270 | ~n2271;
  assign n9793 = n2275 | n2276;
  assign n9794 = n2277 | n2278;
  assign n9795 = n2279 | ~n2280;
  assign n9796 = n2284 | ~n2285;
  assign n9797 = n2287 | ~n2288;
  assign n9798 = n2291 | n2292;
  assign n9799 = n2293 | n2294;
  assign n9800 = n2307 | n2303 | n2306;
  assign n9801 = n2315 | ~n2316;
  assign n9802 = n2318 | n2319;
  assign n9803 = n2321 | ~n2322;
  assign n9804 = n2325 | n2326;
  assign n9805 = n2329 | n2330;
  assign n9806 = n2343 | n2344;
  assign n9807 = n2356 | n2352 | n2355;
  assign n9808 = n2361 | ~n2362;
  assign n9809 = n2370 | n2371;
  assign n9810 = n2381 | n2382;
  assign n9811 = n2387 | n2388;
  assign n9812 = n2392 | n2393;
  assign n9813 = n2395 | n2396;
  assign n9814 = n2402 | n2403;
  assign n9815 = n2406 | n2407;
  assign n9816 = n2422 | n2418 | n2421;
  assign n9817 = n2430 | n2431;
  assign n9818 = n2436 | ~n2437;
  assign n9819 = n2445 | n2446;
  assign n9820 = n2459 | ~n2460;
  assign n9821 = n2462 | n2463;
  assign n9822 = n2464 | n2465;
  assign n9823 = n2466 | ~n2467;
  assign n9824 = n2477 | ~n2478;
  assign n9825 = n2480 | n2481;
  assign n9826 = n2482 | n2483;
  assign n9827 = n2484 | ~n2485;
  assign n9828 = n2496 | n2493 | n2495;
  assign n9829 = n2509 | n2517 | n2524 | n2525;
  assign n9830 = n2543 | n2535 | n2542;
  assign n9831 = n2552 | n2553;
  assign n9832 = n2561 | n2567 | n2575 | n2576;
  assign n9833 = n2588 | n2591 | n2597 | n2598;
  assign n9834 = n2611 | n2612;
  assign n9835 = n2614 | n2615;
  assign n9836 = n2618 | ~n2619;
  assign n9837 = n2630 | n2631;
  assign n9838 = n2638 | n2639;
  assign n9839 = n2642 | n2643;
  assign n9840 = n2658 | n2654 | n2657;
  assign n9841 = n2666 | n2667;
  assign n9842 = n2672 | ~n2673;
  assign n9843 = n2681 | n2682;
  assign n9844 = n2688 | n2689;
  assign n9845 = n2690 | n2691;
  assign n9846 = n2692 | ~n2693;
  assign n9847 = n2706 | n2707;
  assign n9848 = n2708 | n2709;
  assign n9849 = n2710 | ~n2711;
  assign n9850 = n2722 | n2723;
  assign n9851 = n2729 | n2730;
  assign n9852 = n2733 | n2734;
  assign n9853 = n2747 | n2743 | n2746;
  assign n9854 = n2755 | n2756;
  assign n9855 = n2761 | ~n2762;
  assign n9856 = n2770 | n2771;
  assign n9857 = n2781 | ~n2782;
  assign n9858 = n2787 | ~n2788;
  assign n9859 = n2790 | n2791;
  assign n9860 = n2792 | n2793;
  assign n9861 = n2794 | ~n2795;
  assign n9862 = n2806 | ~n2807;
  assign n9863 = n2819 | n2820;
  assign n9864 = n2823 | n2824;
  assign n9865 = n2832 | n2833;
  assign n9866 = n2840 | n2841;
  assign n9867 = n2848 | n2849;
  assign n9868 = n2850 | n2851;
  assign n9869 = n2852 | ~n2853;
  assign n9870 = ~n2860 | n2856 | n2859;
  assign n9871 = n2878 | n2879;
  assign n9872 = n2891 | n2887 | n2890;
  assign n9873 = n2900 | n2898 | n2899;
  assign n9874 = n2910 | n2911;
  assign n9875 = n2916 | ~n2917;
  assign n9876 = n2929 | n2930;
  assign n9877 = n2938 | n2939;
  assign n9878 = n2944 | ~n2945;
  assign n9879 = n2953 | n2954;
  assign n9880 = n2959 | n2960;
  assign n9881 = n2961 | n2962;
  assign n9882 = n2963 | ~n2964;
  assign n9883 = n2966 | n2967;
  assign n9884 = n2968 | n2969;
  assign n9885 = n2970 | ~n2971;
  assign n9886 = n2982 | ~n2983;
  assign n9887 = n2991 | n2992;
  assign n9888 = n3000 | n3001;
  assign n9889 = n3013 | n3009 | n3012;
  assign n9890 = n3018 | ~n3019;
  assign n9891 = n3027 | n3028;
  assign n9892 = n3032 | n3033;
  assign n9893 = n3038 | n3039;
  assign n9894 = n3041 | ~n3042;
  assign n9895 = n3046 | n3047;
  assign n9896 = n3048 | n3049;
  assign n9897 = n3050 | ~n3051;
  assign n9898 = n3056 | ~n3057;
  assign n9899 = n3061 | ~n3062;
  assign n9900 = n3075 | ~n3076;
  assign n9901 = n3086 | n3087;
  assign n9902 = n3098 | n3099;
  assign n9903 = n3107 | n3108;
  assign n9904 = n3113 | ~n3114;
  assign n9905 = n3122 | n3123;
  assign n9906 = n3129 | ~n3130;
  assign n9907 = n3134 | n3135;
  assign n9908 = n3136 | n3137;
  assign n9909 = n3138 | ~n3139;
  assign n9910 = n3144 | ~n3145;
  assign n9911 = n3154 | n3155;
  assign n9912 = n3165 | n3166;
  assign n9913 = n3179 | n3175 | n3178;
  assign n9914 = n3184 | ~n3185;
  assign n9915 = n3207 | n3208;
  assign n9916 = n3216 | n3217;
  assign n9917 = n3224 | n3225;
  assign n9918 = n3235 | n3236;
  assign n9919 = n3241 | ~n3242;
  assign n9920 = n3252 | n3250 | n3251;
  assign n9921 = n3262 | n3263;
  assign n9922 = n3274 | n3275;
  assign n9923 = n3283 | n3284;
  assign n9924 = n3289 | n3290;
  assign n9925 = n3292 | n3293;
  assign n9926 = n3295 | n3296;
  assign n9927 = n3297 | ~n3298;
  assign n9928 = n3328 | n3325 | n3327;
  assign n9929 = n3331 | n3332;
  assign n9930 = n3338 | n3335 | ~n3337;
  assign n9931 = n3352 | n3345 | ~n3351;
  assign n9932 = n3349 | n3350;
  assign n9933 = n3357 | n3358;
  assign n9934 = n3359 | ~n3360;
  assign n9935 = n3365 | n3366;
  assign n9936 = n3368 | n3369;
  assign n9937 = n3371 | n3372;
  assign n9938 = n3376 | n3373 | n3375;
  assign n9939 = n3377 | ~n3378;
  assign n9940 = n3383 | ~n3384;
  assign n9941 = n3394 | n3395;
  assign n9942 = n3403 | n3404;
  assign n9943 = n3409 | ~n3410;
  assign n9944 = n3418 | n3419;
  assign n9945 = n3430 | ~n3431;
  assign n9946 = n3432 | n3433;
  assign n9947 = n3447 | n3448;
  assign n9948 = n3456 | n3457;
  assign n9949 = n3462 | ~n3463;
  assign n9950 = n3475 | n3471 | n3474;
  assign n9951 = n3478 | n3479;
  assign n9952 = n3480 | n3481;
  assign n9953 = n3482 | ~n3483;
  assign n9954 = n3493 | n3494;
  assign n9955 = n3496 | ~n3497;
  assign n9956 = n3498 | n3499;
  assign n9957 = n3511 | ~n3512;
  assign n9958 = n3528 | n3523 | ~n3527;
  assign n9959 = n3537 | n3532 | ~n3536;
  assign n9960 = n3544 | n3545;
  assign n9961 = n3547 | ~n3548;
  assign n9962 = n3556 | ~n3557;
  assign n9963 = n3564 | n3565;
  assign n9964 = n3567 | ~n3568;
  assign n9965 = n3586 | ~n3587;
  assign n9966 = n3597 | ~n3598;
  assign n9967 = n3608 | ~n3609;
  assign n9968 = n3620 | ~n3621;
  assign n9969 = n3628 | n3629;
  assign n9970 = n3634 | ~n3635;
  assign n9971 = n3640 | ~n3641;
  assign n9972 = n3657 | n3652 | n3656;
  assign n9973 = n3663 | n3664;
  assign n9974 = n3669 | n3670;
  assign n9975 = n3673 | n3674;
  assign n9976 = n3679 | n3680;
  assign n9977 = n3686 | n3687;
  assign n9978 = n3693 | n3694;
  assign n9979 = n3699 | n3700;
  assign n9980 = n3703 | n3704;
  assign n9981 = n3707 | n3708;
  assign n9982 = n3716 | n3717;
  assign n9983 = n3731 | n3724 | n3730;
  assign n9984 = n3728 | n3729;
  assign n9985 = n3750 | n3743 | n3749;
  assign n9986 = n3758 | n3759;
  assign n9987 = n3773 | n3774;
  assign n9988 = n3805 | n3796 | n3804;
  assign n9989 = n3820 | n3821;
  assign n9990 = n3827 | n3828;
  assign n9991 = n3837 | n3833 | n3836;
  assign n9992 = n3842 | n3843;
  assign n9993 = n3847 | n3848;
  assign n9994 = n3859 | n3860;
  assign n9995 = n3869 | n3874 | n3879 | n3880;
  assign n9996 = n3891 | n3892;
  assign n9997 = n3895 | n3896;
  assign n9998 = n3902 | n3899 | n3901;
  assign n9999 = n3906 | n3907;
  assign n10000 = n3917 | n3918;
  assign n10001 = n3932 | n3929 | n3931;
  assign n10002 = n3938 | n3939;
  assign n10003 = n3942 | n3943;
  assign n10004 = n3959 | n3970 | n3978 | n3979;
  assign n10005 = n3962 | n3963;
  assign n10006 = n3966 | n3967;
  assign n10007 = n3981 | n3982;
  assign n10008 = n3986 | n3987;
  assign n10009 = n3995 | n3992 | n3994;
  assign n10010 = n4001 | n4002;
  assign n10011 = n4015 | n4016;
  assign n10012 = n4022 | n4023;
  assign n10013 = n4042 | n4035 | n4041;
  assign n10014 = n4050 | n4051;
  assign n10015 = n4057 | n4061 | n4063 | n4064;
  assign n10016 = n4069 | n4070;
  assign n10017 = n4084 | n4078 | n4083;
  assign n10018 = n4100 | n4095 | n4099;
  assign n10019 = n4113 | n4114;
  assign n10020 = n4120 | n4121;
  assign n10021 = n4124 | n4125;
  assign n10022 = n4141 | n4137 | n4140;
  assign n10023 = n4147 | n4148;
  assign n10024 = n4150 | n4151;
  assign n10025 = n4178 | n4166 | n4177;
  assign n10026 = n4190 | n4191;
  assign n10027 = n4197 | n4198;
  assign n10028 = n4209 | n4206 | n4208;
  assign n10029 = n4210 | n4211;
  assign n10030 = n4220 | n4221;
  assign n10031 = n4224 | n4225;
  assign n10032 = n4228 | n4229;
  assign n10033 = n4240 | n4241;
  assign n10034 = n4250 | n4251;
  assign n10035 = n4267 | n4261 | n4266;
  assign n10036 = n4286 | n4278 | n4285;
  assign n10037 = n4298 | n4299;
  assign n10038 = n4311 | n4307 | n4310;
  assign n10039 = n4321 | n4322;
  assign n10040 = n4333 | n4334;
  assign n10041 = n4346 | n4343 | n4345;
  assign n10042 = n4362 | n4363;
  assign n10043 = n4378 | n4379;
  assign n10044 = n4386 | n4387;
  assign n10045 = n4395 | n4390 | n4394;
  assign n10046 = n4392 | n4393;
  assign n10047 = n4410 | n4419 | n4430 | n4431;
  assign n10048 = n4422 | n4423;
  assign n10049 = n4442 | n4443;
  assign n10050 = n4451 | n4452;
  assign n10051 = n4457 | n4458;
  assign n10052 = n4469 | n4470;
  assign n10053 = n4476 | n4477;
  assign n10054 = n4482 | n4483;
  assign n10055 = n4492 | n4493;
  assign n10056 = n4499 | n4500;
  assign n10057 = n4503 | n4504;
  assign n10058 = n4508 | n4509;
  assign n10059 = n4522 | n4516 | n4521;
  assign n10060 = n4519 | n4520;
  assign n10061 = n4532 | n4528 | n4531;
  assign n10062 = n4542 | n4539 | n4541;
  assign n10063 = n4557 | n4554 | n4556;
  assign n10064 = n4562 | ~n4563;
  assign n10065 = n4584 | n4585;
  assign n10066 = n4590 | n4591;
  assign n10067 = n4596 | n4597;
  assign n10068 = n4610 | n4611;
  assign n10069 = n4616 | ~n4617;
  assign n10070 = n4623 | n4624;
  assign n10071 = n4633 | n4634;
  assign n10072 = n4647 | n4648;
  assign n10073 = n4656 | n4650 | n4655;
  assign n10074 = n4659 | n4660;
  assign n10075 = n4668 | n4664 | n4667;
  assign n10076 = n4674 | n4671 | n4673;
  assign n10077 = n4677 | n4678;
  assign n10078 = n4693 | n4694;
  assign n10079 = n4699 | ~n4700;
  assign n10080 = n4705 | ~n4706;
  assign n10081 = n4707 | n4708;
  assign n10082 = n4721 | n4722;
  assign n10083 = n4725 | n4726;
  assign n10084 = n4728 | ~n4729;
  assign n10085 = n4736 | ~n4737;
  assign n10086 = n4745 | ~n4746;
  assign n10087 = n4751 | ~n4752;
  assign n10088 = n4757 | ~n4758;
  assign n10089 = n4769 | ~n4770;
  assign n10090 = n4780 | ~n4781;
  assign n10091 = n4785 | ~n4786;
  assign n10092 = n4788 | n4789;
  assign n10093 = n4794 | n4795;
  assign n10094 = n4835 | n4836;
  assign n10095 = n4844 | n4845;
  assign n10096 = n4846 | n4847;
  assign n10097 = n4852 | n4853;
  assign n10098 = n4866 | n4867;
  assign n10099 = n4884 | ~n4885;
  assign n10100 = n4890 | n4891;
  assign n10101 = n4895 | n4896;
  assign n10102 = n4905 | ~n4906;
  assign n10103 = n4911 | ~n4912;
  assign n10104 = n4917 | ~n4918;
  assign n10105 = n4926 | ~n4927;
  assign n10106 = n4930 | n4931;
  assign n10107 = n4937 | n4938;
  assign n10108 = n4941 | ~n4942;
  assign n10109 = n4950 | ~n4951;
  assign n10110 = n4955 | n4956;
  assign n10111 = n4964 | ~n4965;
  assign n10112 = n4981 | n4982;
  assign n10113 = n4984 | n4985;
  assign n10114 = n4997 | n4998;
  assign n10115 = n5003 | ~n5004;
  assign n10116 = n5013 | ~n5014;
  assign n10117 = n5018 | n5019;
  assign n10118 = n5024 | ~n5025;
  assign n10119 = n5032 | n5033;
  assign n10120 = n5039 | n5040;
  assign n10121 = n5041 | n5042;
  assign n10122 = n5043 | ~n5044;
  assign n10123 = n5068 | n5069;
  assign n10124 = n5076 | ~n5077;
  assign n10125 = n5086 | n5081 | n5085;
  assign n10126 = n5088 | n5089;
  assign n10127 = n5100 | ~n5101;
  assign n10128 = n5106 | ~n5107;
  assign n10129 = n5118 | ~n5119;
  assign n10130 = n5124 | n5125;
  assign n10131 = n5129 | n5130;
  assign n10132 = n5133 | ~n5134;
  assign n10133 = n5142 | ~n5143;
  assign n10134 = n5154 | n5155;
  assign n10135 = n5156 | n5157;
  assign n10136 = n5173 | ~n5174;
  assign n10137 = n5179 | n5180;
  assign n10138 = n5181 | n5182;
  assign n10139 = n5183 | ~n5184;
  assign n10140 = n5187 | n5188;
  assign n10141 = n5189 | n5190;
  assign n10142 = n5191 | ~n5192;
  assign n10143 = n5201 | n5202;
  assign n10144 = n5203 | n5204;
  assign n10145 = n5210 | n5211;
  assign n10146 = n5220 | n5221;
  assign n10147 = n5224 | ~n5225;
  assign n10148 = n5233 | n5234;
  assign n10149 = n5247 | n5248;
  assign n10150 = n5257 | ~n5258;
  assign n10151 = n5262 | n5263;
  assign n10152 = n5271 | n5272;
  assign n10153 = n5275 | n5276;
  assign n10154 = n5277 | n5278;
  assign n10155 = n5281 | n5282;
  assign n10156 = n5283 | n5284;
  assign n10157 = n5285 | ~n5286;
  assign n10158 = n5296 | ~n5297;
  assign n10159 = n5299 | ~n5300;
  assign n10160 = n5306 | ~n5307;
  assign n10161 = n5309 | ~n5310;
  assign n10162 = n5327 | n5325 | n5326;
  assign n10163 = n5336 | n5337;
  assign n10164 = n5342 | n5343;
  assign n10165 = n5344 | n5345;
  assign n10166 = n5348 | n5349;
  assign n10167 = n5357 | n5351 | ~n5356;
  assign n10168 = n5353 | ~n5354;
  assign n10169 = n5362 | ~n5363;
  assign n10170 = n5377 | ~n5378;
  assign n10171 = n5386 | ~n5387;
  assign n10172 = n5392 | ~n5393;
  assign n10173 = n5410 | ~n5411;
  assign n10174 = n5421 | n5422;
  assign n10175 = n5425 | ~n5426;
  assign n10176 = n5442 | ~n5443;
  assign n10177 = n5448 | n5449;
  assign n10178 = n5450 | n5451;
  assign n10179 = n5452 | ~n5453;
  assign n10180 = n5461 | n5462;
  assign n10181 = n5465 | ~n5466;
  assign n10182 = n5495 | ~n5496;
  assign n10183 = n5503 | ~n5504;
  assign n10184 = n5520 | n5521;
  assign n10185 = n5529 | n5530;
  assign n10186 = n5533 | ~n5534;
  assign n10187 = n5542 | n5543;
  assign n10188 = n5555 | n5556;
  assign n10189 = n5565 | ~n5566;
  assign n10190 = n5570 | n5571;
  assign n10191 = n5579 | n5580;
  assign n10192 = n5586 | n5587;
  assign n10193 = n5588 | n5589;
  assign n10194 = n5590 | ~n5591;
  assign n10195 = n5605 | ~n5606;
  assign n10196 = n5616 | ~n5617;
  assign n10197 = n5621 | n5622;
  assign n10198 = n5623 | n5624;
  assign n10199 = n5625 | ~n5626;
  assign n10200 = n5636 | ~n5637;
  assign n10201 = n5643 | ~n5644;
  assign n10202 = n5650 | n5651;
  assign n10203 = n5659 | n5660;
  assign n10204 = n5663 | n5664;
  assign n10205 = n5669 | n5666 | n5668;
  assign n10206 = n5705 | n5687 | n5696 | n5714 | n5715;
  assign n10207 = n5721 | n5718 | n5720;
  assign n10208 = n5750 | n5739 | n5749;
  assign n10209 = n5764 | n5765;
  assign n10210 = n5770 | ~n5771;
  assign n10211 = n5773 | n5774;
  assign n10212 = n5796 | n5797;
  assign n10213 = n5800 | ~n5801;
  assign n10214 = n5823 | n5824;
  assign n10215 = n5830 | n5831;
  assign n10216 = n5836 | ~n5837;
  assign n10217 = n5842 | ~n5843;
  assign n10218 = n5848 | ~n5849;
  assign n10219 = n5854 | ~n5855;
  assign n10220 = n5876 | ~n5877;
  assign n10221 = n5888 | n5893 | n5900 | n5901;
  assign n10222 = n5916 | n5917;
  assign n10223 = n5925 | n5926;
  assign n10224 = n5931 | n5932;
  assign n10225 = n5946 | n5947;
  assign n10226 = n5952 | ~n5953;
  assign n10227 = n5957 | n5958;
  assign n10228 = n5962 | n5963;
  assign n10229 = n5970 | n5971;
  assign n10230 = n5972 | ~n5973;
  assign n10231 = n5983 | n5984;
  assign n10232 = n5989 | n5990;
  assign n10233 = n5998 | n5999;
  assign n10234 = n6007 | ~n6008;
  assign n10235 = n6025 | ~n6026;
  assign n10236 = n6043 | ~n6044;
  assign n10237 = n6052 | ~n6053;
  assign n10238 = ~n6078 | n6069 | ~n6077;
  assign n10239 = n6072 | n6073;
  assign n10240 = n6102 | n6103;
  assign n10241 = n6106 | n6107;
  assign n10242 = n6121 | n6117 | ~n6120;
  assign n10243 = n6130 | n6131;
  assign n10244 = n6137 | n6138;
  assign n10245 = n6139 | ~n6140;
  assign n10246 = n6144 | n6142 | n6143;
  assign n10247 = n6148 | n6149;
  assign n10248 = n6156 | ~n6157;
  assign n10249 = n6162 | n6163;
  assign n10250 = n6168 | n6169;
  assign n10251 = n6194 | n6202 | n6204 | n6205;
  assign n10252 = n6197 | n6198;
  assign n10253 = n6213 | n6214;
  assign n10254 = n6220 | ~n6221;
  assign n10255 = n6223 | n6224;
  assign n10256 = n6232 | n6233;
  assign n10257 = n6238 | ~n6239;
  assign n10258 = n6241 | n6242;
  assign n10259 = n6246 | n6247;
  assign n10260 = n6259 | n6260;
  assign n10261 = n6261 | n6262;
  assign n10262 = n6267 | n6268;
  assign n10263 = n6270 | ~n6271;
  assign n10264 = n6282 | n6283;
  assign n10265 = n6289 | ~n6290;
  assign n10266 = n6294 | n6295;
  assign n10267 = n6296 | ~n6297;
  assign n10268 = n6307 | n6308;
  assign n10269 = n6309 | n6310;
  assign n10270 = n6319 | n6320;
  assign n10271 = n6326 | n6327;
  assign n10272 = n6329 | n6330;
  assign n10273 = n6334 | ~n6335;
  assign n10274 = n6346 | ~n6347;
  assign n10275 = n6349 | n6350;
  assign n10276 = n6354 | n6355;
  assign n10277 = n6372 | n6364 | ~n6371;
  assign n10278 = n6368 | n6369;
  assign n10279 = n6378 | ~n6379;
  assign n10280 = n6381 | n6382;
  assign n10281 = n6386 | n6387;
  assign n10282 = n6398 | n6399;
  assign n10283 = n6400 | n6401;
  assign n10284 = n6406 | n6407;
  assign n10285 = n6409 | ~n6410;
  assign n10286 = n6416 | ~n6417;
  assign n10287 = n6429 | n6430;
  assign n10288 = n6447 | n6440 | n6446;
  assign n10289 = n6473 | n6462 | n6472;
  assign n10290 = n6488 | n6489;
  assign n10291 = n6493 | n6494;
  assign n10292 = n6495 | n6496;
  assign n10293 = n6502 | n6503;
  assign n10294 = n6510 | n6511;
  assign n10295 = n6512 | n6513;
  assign n10296 = n6525 | n6526;
  assign n10297 = n6527 | n6528;
  assign n10298 = n6552 | n6553;
  assign n10299 = n6556 | ~n6557;
  assign n10300 = n6565 | ~n6566;
  assign n10301 = n6571 | ~n6572;
  assign n10302 = n6577 | ~n6578;
  assign n10303 = n6590 | ~n6591;
  assign n10304 = n6599 | ~n6600;
  assign n10305 = n6605 | ~n6606;
  assign n10306 = n6611 | ~n6612;
  assign n10307 = n6618 | n6619;
  assign n10308 = n6625 | n6622 | n6624;
  assign n10309 = n6640 | n6641;
  assign n10310 = n6651 | n6652;
  assign n10311 = n6656 | n6657;
  assign n10312 = n6662 | n6659 | n6661;
  assign n10313 = n6685 | n6676 | n6684;
  assign n10314 = n6694 | n6695;
  assign n10315 = n6700 | n6701;
  assign n10316 = n6705 | n6706;
  assign n10317 = n6713 | n6714;
  assign n10318 = n6731 | n6728 | n6730;
  assign n10319 = n6734 | n6735;
  assign n10320 = n6748 | n6749;
  assign n10321 = n6753 | n6754;
  assign n10322 = n6761 | n6762;
  assign n10323 = n6778 | n6769 | n6777;
  assign n10324 = n6787 | n6788;
  assign n10325 = n6793 | n6794;
  assign n10326 = n6798 | n6799;
  assign n10327 = n6808 | n6803 | n6807;
  assign n10328 = n6816 | n6820 | n6826 | n6827;
  assign n10329 = n6836 | n6837;
  assign n10330 = n6856 | n6848 | n6855;
  assign n10331 = n6870 | n6871;
  assign n10332 = n6882 | n6879 | n6881;
  assign n10333 = n6888 | n6889;
  assign n10334 = n6896 | n6897;
  assign n10335 = n6902 | n6903;
  assign n10336 = n6911 | n6912;
  assign n10337 = n6918 | n6919;
  assign n10338 = n6920 | n6921;
  assign n10339 = n6936 | n6933 | n6935;
  assign n10340 = n6939 | n6940;
  assign n10341 = n6945 | ~n6946;
  assign n10342 = ~n6956 | n6949 | n6955;
  assign n10343 = n6952 | ~n6953;
  assign n10344 = n6960 | n6961;
  assign n10345 = n6962 | n6963;
  assign n10346 = n6965 | ~n6966;
  assign n10347 = n6969 | n6970;
  assign n10348 = n6971 | n6972;
  assign n10349 = n6973 | ~n6974;
  assign n10350 = n6979 | ~n6980;
  assign n10351 = n6992 | n6993;
  assign n10352 = n7000 | n7001;
  assign n10353 = n7008 | n7009;
  assign n10354 = n7012 | n7013;
  assign n10355 = n7025 | n7026;
  assign n10356 = n7027 | n7028;
  assign n10357 = n7029 | n7030;
  assign n10358 = n7033 | ~n7034;
  assign n10359 = n7041 | n7042;
  assign n10360 = n7047 | n7048;
  assign n10361 = n7049 | n7050;
  assign n10362 = n7060 | n7061;
  assign n10363 = n7064 | n7065;
  assign n10364 = n7066 | n7067;
  assign n10365 = n7078 | ~n7079;
  assign n10366 = n7099 | n7100;
  assign n10367 = n7101 | n7102;
  assign n10368 = n7103 | ~n7104;
  assign n10369 = n7107 | n7108;
  assign n10370 = n7109 | n7110;
  assign n10371 = n7111 | ~n7112;
  assign n10372 = n7115 | n7116;
  assign n10373 = n7117 | n7118;
  assign n10374 = n7119 | ~n7120;
  assign n10375 = n7125 | ~n7126;
  assign n10376 = n7138 | ~n7139;
  assign n10377 = n7147 | ~n7148;
  assign n10378 = n7153 | ~n7154;
  assign n10379 = n7159 | ~n7160;
  assign n10380 = n7166 | n7168 | n7170 | n7171;
  assign n10381 = n7203 | n7192 | n7202;
  assign n10382 = n7204 | n7205;
  assign n10383 = n7217 | n7219 | n7221 | n7222;
  assign n10384 = n7232 | n7233;
  assign n10385 = n7239 | n7240;
  assign n10386 = n7245 | ~n7246;
  assign n10387 = n7248 | n7249;
  assign n10388 = n7254 | n7255;
  assign n10389 = n7256 | n7257;
  assign n10390 = n7269 | n7270;
  assign n10391 = n7271 | n7272;
  assign n10392 = n7281 | n7282;
  assign n10393 = n7285 | ~n7286;
  assign n10394 = n7303 | n7304;
  assign n10395 = n7308 | n7309;
  assign n10396 = n7310 | n7311;
  assign n10397 = n7312 | ~n7313;
  assign n10398 = n7316 | n7317;
  assign n10399 = n7318 | n7319;
  assign n10400 = n7320 | ~n7321;
  assign n10401 = n7324 | n7325;
  assign n10402 = n7326 | n7327;
  assign n10403 = n7328 | ~n7329;
  assign n10404 = n7334 | ~n7335;
  assign n10405 = n7347 | ~n7348;
  assign n10406 = n7356 | ~n7357;
  assign n10407 = n7362 | ~n7363;
  assign n10408 = n7368 | ~n7369;
  assign n10409 = n7374 | ~n7375;
  assign n10410 = n7378 | n7379;
  assign n10411 = n7391 | n7385 | n7390;
  assign n10412 = n7411 | n7403 | n7410;
  assign n10413 = n7424 | n7425;
  assign n10414 = n7430 | n7431;
  assign n10415 = n7436 | ~n7437;
  assign n10416 = n7454 | ~n7455;
  assign n10417 = n7457 | n7458;
  assign n10418 = n7459 | n7460;
  assign n10419 = n7471 | n7472;
  assign n10420 = n7473 | n7474;
  assign n10421 = n7485 | ~n7486;
  assign n10422 = n7497 | n7498;
  assign n10423 = n7505 | n7506;
  assign n10424 = n7510 | n7511;
  assign n10425 = n7512 | n7513;
  assign n10426 = n7514 | ~n7515;
  assign n10427 = n7526 | ~n7527;
  assign n10428 = n7532 | n7533;
  assign n10429 = n7540 | ~n7541;
  assign n10430 = n7567 | n7568;
  assign n10431 = n7584 | n7576 | n7583;
  assign n10432 = n7599 | n7600;
  assign n10433 = n7605 | ~n7606;
  assign n10434 = n7609 | n7610;
  assign n10435 = n7616 | ~n7617;
  assign n10436 = n7633 | n7634;
  assign n10437 = n7635 | n7636;
  assign n10438 = n7645 | n7646;
  assign n10439 = n7659 | n7660;
  assign n10440 = n7661 | n7662;
  assign n10441 = n7666 | n7667;
  assign n10442 = n7671 | n7672;
  assign n10443 = n7673 | ~n7674;
  assign n10444 = n7679 | ~n7680;
  assign n10445 = n7688 | ~n7689;
  assign n10446 = n7692 | n7693;
  assign n10447 = n7694 | n7695;
  assign n10448 = n7696 | ~n7697;
  assign n10449 = n7702 | ~n7703;
  assign n10450 = n7713 | n7714;
  assign n10451 = n7739 | n7740;
  assign n10452 = n7748 | n7743 | n7747;
  assign n10453 = n7763 | n7760 | n7762;
  assign n10454 = n7782 | n7783;
  assign n10455 = n7799 | n7800;
  assign n10456 = n7801 | n7802;
  assign n10457 = n7821 | n7822;
  assign n10458 = n7825 | ~n7826;
  assign n10459 = n7832 | n7833;
  assign n10460 = n7837 | n7838;
  assign n10461 = n7839 | ~n7840;
  assign n10462 = n7845 | ~n7846;
  assign n10463 = n7851 | ~n7852;
  assign n10464 = n7855 | n7856;
  assign n10465 = n7862 | ~n7863;
  assign n10466 = n7866 | n7867;
  assign n10467 = n7873 | ~n7874;
  assign n10468 = n7877 | n7878;
  assign n10469 = n7890 | n7891;
  assign n10470 = n7894 | n7895;
  assign n10471 = n7897 | n7898;
  assign n10472 = n7913 | n7904 | n7912;
  assign n10473 = n7909 | n7910;
  assign n10474 = n7929 | n7926 | n7928;
  assign n10475 = n7952 | ~n7953;
  assign n10476 = n7961 | n7962;
  assign n10477 = n7969 | n7970;
  assign n10478 = n7971 | n7972;
  assign n10479 = n7993 | ~n7994;
  assign n10480 = n8000 | n8001;
  assign n10481 = n8005 | n8006;
  assign n10482 = n8007 | ~n8008;
  assign n10483 = n8013 | ~n8014;
  assign n10484 = n8019 | ~n8020;
  assign n10485 = n8023 | n8024;
  assign n10486 = n8030 | ~n8031;
  assign n10487 = n8034 | n8035;
  assign n10488 = n8051 | n8052;
  assign n10489 = n8069 | n8061 | n8068;
  assign n10490 = n8076 | n8077;
  assign n10491 = n8085 | n8086;
  assign n10492 = n8097 | n8098;
  assign n10493 = n8120 | n8121;
  assign n10494 = n8126 | ~n8127;
  assign n10495 = n8143 | ~n8144;
  assign n10496 = n8155 | n8156;
  assign n10497 = n8159 | n8160;
  assign n10498 = n8161 | n8162;
  assign n10499 = n8173 | n8174;
  assign n10500 = n8175 | n8176;
  assign n10501 = n8177 | ~n8178;
  assign n10502 = n8183 | ~n8184;
  assign n10503 = n8189 | ~n8190;
  assign n10504 = n8195 | ~n8196;
  assign n10505 = n8201 | ~n8202;
  assign n10506 = n8207 | ~n8208;
  assign n10507 = n8227 | n8228;
  assign n10508 = n8240 | n8241;
  assign n10509 = n8260 | n8261;
  assign n10510 = n8266 | n8267;
  assign n10511 = n8268 | n8269;
  assign n10512 = n8291 | ~n8292;
  assign n10513 = n8300 | n8301;
  assign n10514 = n8302 | n8303;
  assign n10515 = n8304 | ~n8305;
  assign n10516 = n8313 | ~n8314;
  assign n10517 = n8317 | n8318;
  assign n10518 = n8345 | n8338 | n8344;
  assign n10519 = n8355 | n8356;
  assign n10520 = n8372 | n8365 | n8371;
  assign n10521 = n8386 | n8387;
  assign n10522 = n8410 | ~n8411;
  assign n10523 = n8419 | n8420;
  assign n10524 = n8438 | n8439;
  assign n10525 = n8440 | n8441;
  assign n10526 = n8448 | ~n8449;
  assign n10527 = n8454 | ~n8455;
  assign n10528 = n8460 | ~n8461;
  assign n10529 = n8466 | ~n8467;
  assign n10530 = n8472 | ~n8473;
  assign n10531 = n8488 | n8489;
  assign n10532 = n8504 | n8505;
  assign n10533 = n8506 | n8507;
  assign n10534 = n8520 | n8521;
  assign n10535 = n8543 | n8544;
  assign n10536 = n8549 | ~n8550;
  assign n10537 = n8558 | ~n8559;
  assign n10538 = n8568 | n8569;
  assign n10539 = n8570 | n8571;
  assign n10540 = n8579 | n8580;
  assign n10541 = n8581 | n8582;
  assign n10542 = n8584 | ~n8585;
  assign n10543 = n8586 | n8587;
  assign n10544 = n8589 | n8590;
  assign n10545 = n8592 | n8593;
  assign n10546 = n8599 | ~n8600;
  assign n10547 = n8605 | ~n8606;
  assign n10548 = n8612 | n8609 | n8611;
  assign n10549 = n8627 | n8624 | n8626;
  assign n10550 = n8632 | n8633;
  assign n10551 = n8647 | n8648;
  assign n10552 = n8667 | n8668;
  assign n10553 = n8683 | ~n8684;
  assign n10554 = n8693 | ~n8694;
  assign n10555 = ~n8702 | n8700 | ~n8701;
  assign n10556 = n8707 | ~n8708;
  assign n10557 = n8711 | n8712;
  assign n10558 = n8730 | n8731;
  assign n10559 = n8751 | n8752;
  assign n10560 = n8753 | n8754;
  assign n10561 = n8757 | n8758;
  assign n10562 = n8763 | ~n8764;
  assign n10563 = n8766 | n8767;
  assign n10564 = n8774 | n8775;
  assign n10565 = n8776 | n8777;
  assign n10566 = n8783 | ~n8784;
  assign n10567 = n8789 | ~n8790;
  assign n10568 = n8795 | ~n8796;
  assign n10569 = n8801 | ~n8802;
  assign n10570 = n8814 | n8818 | n8821 | n8822;
  assign n10571 = n8823 | ~n8824;
  assign n10572 = n8830 | n8831;
  assign n10573 = n8843 | n8840 | n8842;
  assign n10574 = n8864 | n8865;
  assign n10575 = n8870 | n8871;
  assign n10576 = n8872 | n8873;
  assign n10577 = n8884 | n8885;
  assign n10578 = n8886 | n8887;
  assign n10579 = n8888 | ~n8889;
  assign n10580 = n8894 | ~n8895;
  assign n10581 = n8907 | n8910 | n8914 | n8915;
  assign n10582 = n8938 | n8930 | n8937;
  assign n10583 = n8954 | n8955;
  assign n10584 = n8960 | n8961;
  assign n10585 = n8966 | ~n8967;
  assign n10586 = n8979 | n8980;
  assign n10587 = n8985 | ~n8986;
  assign n10588 = n8994 | n8995;
  assign n10589 = n8996 | n8997;
  assign n10590 = n8998 | ~n8999;
  assign n10591 = n9027 | n9028;
  assign n10592 = n9029 | n9030;
  assign n10593 = n9047 | n9048;
  assign n10594 = n9069 | ~n9070;
  assign n10595 = n9075 | n9076;
  assign n10596 = n9077 | n9078;
  assign n10597 = n9081 | n9082;
  assign n10598 = n9083 | n9084;
  assign n10599 = n9085 | n9086;
  assign n10600 = n9087 | ~n9088;
  assign n10601 = n9101 | n9098 | n9100;
  assign n10602 = n9104 | n9105;
  assign n10603 = n9110 | n9111;
  assign n10604 = n9117 | n9118;
  assign n10605 = n9132 | n9133;
  assign n10606 = n9138 | n9139;
  assign n10607 = n9144 | ~n9145;
  assign n10608 = n9159 | n9156 | n9158;
  assign n10609 = n9174 | n9175;
  assign n10610 = n9176 | n9177;
  assign n10611 = n9181 | n9179 | n9180;
  assign n10612 = n9187 | n9188;
  assign n10613 = n9192 | ~n9193;
  assign n10614 = n9196 | n9194 | n9195;
  assign n10615 = n9207 | ~n9208;
  assign n10616 = n9217 | n9214 | n9216;
  assign n10617 = n9218 | n9219;
  assign n10618 = n9221 | ~n9222;
  assign n10619 = n9223 | n9224;
  assign n10620 = n9225 | ~n9226;
  assign n10621 = n9258 | n9250 | n9257;
  assign n10622 = n9271 | n9272;
  assign n10623 = n9282 | n9283;
  assign n10624 = n9284 | n9285;
  assign n10625 = n9300 | n9295 | n9299;
  assign n10626 = n9320 | n9317 | n9319;
  assign n10627 = n9329 | ~n9330;
  assign n10628 = n9333 | n9334;
  assign n10629 = n9335 | n9336;
  assign n10630 = n9357 | n9348 | n9356;
  assign n10631 = n9370 | n9371;
  assign n10632 = n9386 | n9387;
  assign n10633 = n9388 | n9389;
  assign n10634 = n9398 | n9403 | n9409 | n9410;
  assign n10635 = n9424 | n9425;
  assign n10636 = n9434 | ~n9435;
  assign n10637 = n9438 | n9439;
  assign n10638 = n9440 | n9441;
  assign n10639 = n9448 | n9449;
  assign n10640 = n9459 | n9460;
  assign n10641 = n9464 | n9465;
  assign n10642 = n9466 | n9467;
  assign n10643 = n9489 | n9479 | n9488;
  assign n10644 = n9492 | n9490 | n9491;
  assign n10645 = n9498 | n9499;
  assign n10646 = n9507 | n9513 | n9515 | n9516;
  assign n10647 = n9521 | n9522 | n9524 | n9525;
  assign po0  = ~n10349;
  assign po1  = ~n7235;
  assign po2  = ~n7445;
  assign po4  = ~n7777;
  assign po5  = ~n7943;
  assign po6  = ~n8112;
  assign po7  = ~n8255;
  assign po8  = ~n8401;
  assign po9  = ~n8535;
  assign po10  = ~n8662;
  assign po11  = ~n8745;
  assign po12  = ~n8857;
  assign po13  = ~n8975;
  assign po14  = ~n9062;
  assign po15  = ~n9153;
  assign po16  = ~n9234;
  assign po18  = ~n9337;
  assign po19  = ~n9390;
  assign po20  = ~n9442;
  assign po21  = ~n9468;
  assign po22  = ~n9493;
  assign po23  = ~n10646;
endmodule
