module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n412,
    n413, n414, n415, n416, n417, n418, n419,
    n420, n421, n422, n424, n425, n426, n427,
    n428, n429, n430, n431, n432, n434, n435,
    n436, n437, n438, n439, n440, n441, n442,
    n443, n444, n445, n447, n448, n449, n450,
    n451, n452, n453, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n475, n476, n477, n478, n479, n480, n481,
    n483, n484, n485, n486, n487, n488, n489,
    n491, n492, n493, n494, n495, n496, n497,
    n498, n500, n501, n502, n503, n504, n506,
    n507, n508, n509, n510, n511, n512, n514,
    n515, n516, n517, n518, n519, n520, n521,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n552, n553, n554, n555, n556, n558, n559,
    n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n570, n571, n572, n573, n574,
    n575, n577, n578, n579, n580, n581, n583,
    n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n603, n604, n605,
    n606, n607, n608, n609, n610, n611, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n622, n623, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n686, n687,
    n688, n689, n690, n691, n692, n693, n695,
    n696, n697, n698, n699, n700, n701, n702,
    n703, n704, n705, n706, n707, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n778, n779, n780, n781, n782,
    n783, n785, n786, n787, n788, n789, n790,
    n792, n793, n794, n795, n796, n797, n799,
    n800, n801, n802, n803, n804, n806, n807,
    n808, n809, n810, n811, n813, n814, n815,
    n816, n817, n818, n820, n821, n822, n823,
    n824, n825, n827, n828, n829, n830, n831,
    n832, n834, n835, n836, n837, n838, n839,
    n840, n841, n842, n843, n844, n845, n846,
    n847, n848, n849, n850, n851, n852, n853,
    n855, n856, n857, n858, n859, n860, n861,
    n863, n864, n865, n866, n867, n868, n869,
    n870, n871, n872, n873, n874, n875, n877,
    n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n888, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906,
    n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n921, n922,
    n923, n924, n925, n926, n927, n928, n930,
    n931, n932, n933, n934, n935, n936, n937,
    n938, n939, n940, n941, n942, n943, n944,
    n945, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n960,
    n961, n962, n963, n964, n965, n966, n967,
    n968, n969, n970, n971, n972, n974, n975,
    n976, n977, n978, n979, n980, n981, n982,
    n983, n984, n985, n986, n987, n988, n989,
    n990, n992, n993, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1002, n1003,
    n1004, n1005, n1006, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1021, n1022, n1023,
    n1025, n1026, n1027, n1029, n1030, n1031,
    n1032, n1033, n1034, n1035, n1036, n1037,
    n1038, n1039, n1041, n1042, n1045, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1067, n1068, n1069, n1070, n1071, n1072,
    n1073, n1074, n1075, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1084, n1085,
    n1086, n1087, n1088, n1089, n1091, n1092,
    n1093, n1094, n1095, n1096, n1097, n1098,
    n1099, n1100, n1101, n1102, n1103, n1104,
    n1105, n1106, n1107, n1108, n1109, n1110,
    n1112, n1113, n1114, n1116, n1117, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1129, n1130, n1131, n1132,
    n1134, n1135, n1136, n1137, n1139, n1140,
    n1141, n1142, n1144, n1145, n1146, n1147,
    n1148, n1150, n1151, n1152, n1154, n1155,
    n1156, n1157, n1159, n1160, n1161, n1162,
    n1164, n1165, n1166, n1167, n1169, n1170,
    n1171, n1172, n1174, n1175, n1176, n1178,
    n1179, n1180, n1182, n1183, n1184, n1186,
    n1187, n1188, n1190, n1191, n1192, n1194,
    n1195, n1196, n1198, n1199, n1200, n1201,
    n1202, n1204, n1205, n1206, n1208, n1209,
    n1210, n1212, n1213, n1214, n1216, n1217,
    n1218, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1229, n1230,
    n1231, n1232, n1233, n1234, n1235, n1236,
    n1237, n1239, n1240, n1241, n1243, n1244,
    n1245, n1246, n1248, n1249, n1250, n1252,
    n1253, n1254, n1256, n1257, n1258, n1259,
    n1260, n1262, n1263, n1264, n1266, n1267,
    n1268, n1270, n1271, n1272, n1274, n1275,
    n1276, n1278, n1279, n1280, n1282, n1283,
    n1284, n1285, n1286, n1287, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1297,
    n1298, n1299, n1301, n1302, n1303, n1305,
    n1306, n1307, n1309, n1310, n1311, n1313,
    n1314, n1315, n1317, n1318, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345,
    n1346, n1347, n1348, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1380, n1381, n1382, n1383, n1384,
    n1385, n1386, n1387, n1388, n1389, n1390,
    n1391, n1392, n1393, n1394, n1395, n1396,
    n1398, n1399, n1400, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410,
    n1411, n1412, n1413, n1414, n1415, n1416,
    n1417, n1418, n1420, n1421, n1422, n1423,
    n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435,
    n1436, n1438, n1439, n1440, n1442, n1443,
    n1445, n1446, n1447, n1448, n1450, n1451,
    n1452, n1454, n1455, n1456, n1457, n1459,
    n1460, n1461, n1463, n1464, n1465, n1466,
    n1469, n1470, n1471, n1472, n1475, n1476,
    n1478, n1483, n1484, n1486;
  assign n291 = ~pi4 & ~pi19;
  assign n292 = ~pi18 & n291;
  assign n293 = ~pi16 & n292;
  assign n294 = ~pi9 & ~pi11;
  assign n295 = ~pi13 & ~pi14;
  assign n296 = ~pi5 & ~pi22;
  assign n297 = ~pi17 & ~pi21;
  assign n298 = ~pi8 & n297;
  assign n299 = ~pi7 & ~pi12;
  assign n300 = ~pi6 & n294;
  assign n301 = n295 & n296;
  assign n302 = n299 & n301;
  assign n303 = n298 & n300;
  assign n304 = n302 & n303;
  assign n305 = n293 & n304;
  assign n306 = pi54 & ~n305;
  assign n307 = ~pi0 & ~n306;
  assign n308 = ~pi56 & ~n294;
  assign n309 = n296 & n308;
  assign n310 = ~pi56 & ~n296;
  assign n311 = ~pi8 & ~pi21;
  assign n312 = ~pi7 & pi13;
  assign n313 = n311 & n312;
  assign n314 = pi7 & ~n311;
  assign n315 = ~pi7 & n311;
  assign n316 = pi8 & pi21;
  assign n317 = ~pi13 & ~n316;
  assign n318 = ~n314 & n317;
  assign n319 = ~n315 & n318;
  assign n320 = ~n313 & ~n319;
  assign n321 = ~pi14 & ~n320;
  assign n322 = ~pi13 & pi14;
  assign n323 = n315 & n322;
  assign n324 = ~n321 & ~n323;
  assign n325 = ~pi10 & ~n324;
  assign n326 = pi10 & n295;
  assign n327 = n315 & n326;
  assign n328 = ~n325 & ~n327;
  assign n329 = ~pi6 & ~pi12;
  assign n330 = ~pi17 & n296;
  assign n331 = n329 & n330;
  assign n332 = n293 & n331;
  assign n333 = ~n328 & n332;
  assign n334 = ~n310 & ~n333;
  assign n335 = n294 & ~n334;
  assign n336 = ~n309 & ~n335;
  assign n337 = pi54 & ~n336;
  assign n338 = ~n307 & ~n337;
  assign n339 = ~pi3 & ~pi129;
  assign po15 = n338 | ~n339;
  assign n341 = ~pi7 & ~pi13;
  assign n342 = ~pi5 & ~pi6;
  assign n343 = n341 & n342;
  assign n344 = ~pi11 & ~pi12;
  assign n345 = ~pi10 & ~pi22;
  assign n346 = ~pi14 & n311;
  assign n347 = n344 & n345;
  assign n348 = n346 & n347;
  assign n349 = n343 & n348;
  assign n350 = n293 & n349;
  assign n351 = ~pi17 & pi54;
  assign n352 = ~n350 & n351;
  assign n353 = ~pi1 & ~n352;
  assign n354 = pi5 & ~n329;
  assign n355 = ~pi5 & n329;
  assign n356 = pi6 & pi12;
  assign n357 = ~pi7 & ~n356;
  assign n358 = ~n354 & n357;
  assign n359 = ~n355 & n358;
  assign n360 = pi7 & n355;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~pi13 & ~n361;
  assign n363 = n312 & n355;
  assign n364 = ~n362 & ~n363;
  assign n365 = ~pi9 & ~n364;
  assign n366 = n341 & n355;
  assign n367 = pi9 & n366;
  assign n368 = ~n365 & ~n367;
  assign n369 = ~pi8 & ~pi11;
  assign n370 = n297 & n369;
  assign n371 = ~pi14 & pi54;
  assign n372 = n345 & n371;
  assign n373 = n370 & n372;
  assign n374 = n293 & n373;
  assign n375 = ~n368 & n374;
  assign n376 = ~n353 & ~n375;
  assign po16 = ~n339 | n376;
  assign n378 = ~pi15 & ~pi20;
  assign n379 = ~pi24 & ~pi49;
  assign n380 = n378 & n379;
  assign n381 = ~pi47 & ~pi48;
  assign n382 = ~pi2 & ~pi45;
  assign n383 = n381 & n382;
  assign n384 = n380 & n383;
  assign n385 = ~pi41 & ~pi46;
  assign n386 = ~pi38 & ~pi50;
  assign n387 = n385 & n386;
  assign n388 = ~pi42 & ~pi44;
  assign n389 = ~pi40 & n388;
  assign n390 = ~pi43 & n387;
  assign n391 = n389 & n390;
  assign n392 = n384 & n391;
  assign n393 = pi82 & ~n392;
  assign n394 = pi122 & pi127;
  assign n395 = ~pi65 & ~n394;
  assign n396 = ~n393 & n395;
  assign n397 = ~pi38 & ~pi40;
  assign n398 = n388 & n397;
  assign n399 = ~pi46 & ~pi50;
  assign n400 = ~pi41 & n399;
  assign n401 = n398 & n400;
  assign n402 = ~pi43 & n401;
  assign n403 = ~pi45 & n381;
  assign n404 = n380 & n403;
  assign n405 = n402 & n404;
  assign n406 = pi82 & ~n405;
  assign n407 = ~pi82 & n394;
  assign n408 = ~n406 & ~n407;
  assign n409 = pi2 & ~n408;
  assign n410 = ~n396 & ~n409;
  assign po17 = ~pi129 & ~n410;
  assign n412 = ~pi12 & n370;
  assign n413 = ~pi9 & ~pi14;
  assign n414 = n345 & n413;
  assign n415 = n343 & n414;
  assign n416 = n293 & n412;
  assign n417 = n415 & n416;
  assign n418 = ~pi61 & ~pi118;
  assign n419 = ~n417 & n418;
  assign n420 = pi0 & ~pi113;
  assign n421 = ~pi123 & n420;
  assign n422 = ~n419 & ~n421;
  assign po18 = ~pi129 & ~n422;
  assign n424 = ~pi16 & pi54;
  assign n425 = n292 & n424;
  assign n426 = n370 & n425;
  assign n427 = pi10 & ~pi22;
  assign n428 = n413 & n427;
  assign n429 = n366 & n428;
  assign n430 = n426 & n429;
  assign n431 = pi4 & ~pi54;
  assign n432 = ~n430 & ~n431;
  assign po19 = n339 & ~n432;
  assign n434 = pi5 & ~pi54;
  assign n435 = ~pi13 & n414;
  assign n436 = ~pi59 & n370;
  assign n437 = n435 & n436;
  assign n438 = n299 & n342;
  assign n439 = n424 & n438;
  assign n440 = ~pi25 & pi28;
  assign n441 = ~pi29 & n440;
  assign n442 = n292 & n441;
  assign n443 = n439 & n442;
  assign n444 = n437 & n443;
  assign n445 = ~n434 & ~n444;
  assign po20 = n339 & ~n445;
  assign n447 = pi6 & ~pi54;
  assign n448 = ~pi28 & ~pi29;
  assign n449 = pi25 & n448;
  assign n450 = n292 & n449;
  assign n451 = n439 & n450;
  assign n452 = n437 & n451;
  assign n453 = ~n447 & ~n452;
  assign po21 = n339 & ~n453;
  assign n455 = pi7 & ~pi54;
  assign n456 = ~pi11 & n438;
  assign n457 = n291 & n424;
  assign n458 = pi8 & ~pi17;
  assign n459 = ~pi18 & ~pi21;
  assign n460 = n458 & n459;
  assign n461 = n457 & n460;
  assign n462 = n435 & n461;
  assign n463 = n456 & n462;
  assign n464 = ~n455 & ~n463;
  assign po22 = n339 & ~n464;
  assign n466 = pi8 & ~pi54;
  assign n467 = n366 & n414;
  assign n468 = ~pi17 & ~pi18;
  assign n469 = pi21 & n369;
  assign n470 = n468 & n469;
  assign n471 = n457 & n470;
  assign n472 = n467 & n471;
  assign n473 = ~n466 & ~n472;
  assign po23 = n339 & ~n473;
  assign n475 = pi9 & ~pi54;
  assign n476 = ~pi18 & n298;
  assign n477 = pi11 & n438;
  assign n478 = n457 & n477;
  assign n479 = n435 & n476;
  assign n480 = n478 & n479;
  assign n481 = ~n475 & ~n480;
  assign po24 = n339 & ~n481;
  assign n483 = pi10 & ~pi54;
  assign n484 = ~pi9 & n345;
  assign n485 = n476 & n484;
  assign n486 = n322 & n457;
  assign n487 = n456 & n486;
  assign n488 = n485 & n487;
  assign n489 = ~n483 & ~n488;
  assign po25 = n339 & ~n489;
  assign n491 = pi11 & ~pi54;
  assign n492 = ~pi10 & ~pi11;
  assign n493 = pi22 & n492;
  assign n494 = n413 & n493;
  assign n495 = n457 & n494;
  assign n496 = n366 & n476;
  assign n497 = n495 & n496;
  assign n498 = ~n491 & ~n497;
  assign po26 = n339 & ~n498;
  assign n500 = pi12 & ~pi54;
  assign n501 = pi18 & n457;
  assign n502 = n412 & n501;
  assign n503 = n415 & n502;
  assign n504 = ~n500 & ~n503;
  assign po27 = n339 & ~n504;
  assign n506 = pi13 & ~pi54;
  assign n507 = ~pi25 & ~pi28;
  assign n508 = pi29 & n507;
  assign n509 = n425 & n508;
  assign n510 = n436 & n509;
  assign n511 = n467 & n510;
  assign n512 = ~n506 & ~n511;
  assign po28 = n339 & ~n512;
  assign n514 = pi14 & ~pi54;
  assign n515 = ~pi9 & pi13;
  assign n516 = ~pi16 & n515;
  assign n517 = n291 & n516;
  assign n518 = n372 & n517;
  assign n519 = n456 & n476;
  assign n520 = n518 & n519;
  assign n521 = ~n514 & ~n520;
  assign po29 = n339 & ~n521;
  assign n523 = ~pi43 & ~pi47;
  assign n524 = ~pi48 & n523;
  assign n525 = n400 & n524;
  assign n526 = n398 & n525;
  assign n527 = ~pi45 & n379;
  assign n528 = n526 & n527;
  assign n529 = pi15 & ~n528;
  assign n530 = ~pi15 & n379;
  assign n531 = ~pi2 & ~pi20;
  assign n532 = n403 & ~n531;
  assign n533 = n530 & n532;
  assign n534 = n402 & n533;
  assign n535 = ~n529 & ~n534;
  assign n536 = pi82 & ~n535;
  assign n537 = ~pi46 & n386;
  assign n538 = n389 & n537;
  assign n539 = ~pi45 & ~pi48;
  assign n540 = ~pi41 & ~pi43;
  assign n541 = ~pi47 & n540;
  assign n542 = n539 & n541;
  assign n543 = n538 & n542;
  assign n544 = n530 & n543;
  assign n545 = pi82 & ~n544;
  assign n546 = ~pi70 & ~n394;
  assign n547 = ~n545 & n546;
  assign n548 = pi15 & n407;
  assign n549 = ~n547 & ~n548;
  assign n550 = ~n536 & n549;
  assign po30 = ~pi129 & ~n550;
  assign n552 = pi16 & ~pi54;
  assign n553 = pi6 & n414;
  assign n554 = n426 & n553;
  assign n555 = n362 & n554;
  assign n556 = ~n552 & ~n555;
  assign po31 = n339 & ~n556;
  assign n558 = pi17 & ~pi54;
  assign n559 = ~pi11 & n311;
  assign n560 = ~pi16 & ~pi25;
  assign n561 = pi59 & n560;
  assign n562 = n351 & n448;
  assign n563 = n561 & n562;
  assign n564 = n292 & n438;
  assign n565 = n559 & n564;
  assign n566 = n435 & n563;
  assign n567 = n565 & n566;
  assign n568 = ~n558 & ~n567;
  assign po32 = n339 & ~n568;
  assign n570 = pi18 & ~pi54;
  assign n571 = pi16 & pi54;
  assign n572 = n292 & n571;
  assign n573 = n370 & n572;
  assign n574 = n467 & n573;
  assign n575 = ~n570 & ~n574;
  assign po33 = n339 & ~n575;
  assign n577 = pi19 & ~pi54;
  assign n578 = pi17 & n559;
  assign n579 = n425 & n578;
  assign n580 = n467 & n579;
  assign n581 = ~n577 & ~n580;
  assign po34 = n339 & ~n581;
  assign n583 = n385 & n523;
  assign n584 = n539 & n583;
  assign n585 = ~pi24 & n584;
  assign n586 = ~pi15 & ~pi49;
  assign n587 = ~pi50 & n398;
  assign n588 = n586 & n587;
  assign n589 = n585 & n588;
  assign n590 = pi20 & ~n589;
  assign n591 = ~pi20 & n585;
  assign n592 = n588 & n591;
  assign n593 = pi2 & n592;
  assign n594 = ~n590 & ~n593;
  assign n595 = pi82 & ~n594;
  assign n596 = pi82 & ~n592;
  assign n597 = ~pi71 & ~n394;
  assign n598 = ~n596 & n597;
  assign n599 = pi20 & n407;
  assign n600 = ~n598 & ~n599;
  assign n601 = ~n595 & n600;
  assign po35 = ~pi129 & ~n601;
  assign n603 = pi21 & ~pi54;
  assign n604 = ~pi4 & ~pi16;
  assign n605 = pi19 & ~pi21;
  assign n606 = pi54 & n605;
  assign n607 = n369 & n604;
  assign n608 = n468 & n607;
  assign n609 = n606 & n608;
  assign n610 = n467 & n609;
  assign n611 = ~n603 & ~n610;
  assign po36 = n339 & ~n611;
  assign n613 = pi22 & ~pi54;
  assign n614 = pi5 & ~pi6;
  assign n615 = ~pi7 & n614;
  assign n616 = n295 & n344;
  assign n617 = n615 & n616;
  assign n618 = n457 & n617;
  assign n619 = n485 & n618;
  assign n620 = ~n613 & ~n619;
  assign po37 = n339 & ~n620;
  assign n622 = ~pi23 & pi55;
  assign n623 = pi61 & ~pi129;
  assign po38 = ~n622 & n623;
  assign n625 = n531 & n586;
  assign n626 = n383 & n625;
  assign n627 = n402 & n626;
  assign n628 = pi82 & ~n627;
  assign n629 = pi63 & ~n394;
  assign n630 = ~n628 & n629;
  assign n631 = pi82 & ~n543;
  assign n632 = pi82 & ~n625;
  assign n633 = n394 & ~n632;
  assign n634 = ~n631 & ~n633;
  assign n635 = ~pi24 & ~n634;
  assign n636 = pi24 & pi82;
  assign n637 = n584 & n636;
  assign n638 = n587 & n637;
  assign n639 = ~pi129 & ~n638;
  assign n640 = ~n630 & n639;
  assign po39 = ~n635 & n640;
  assign n642 = pi85 & pi116;
  assign n643 = ~pi85 & ~pi110;
  assign n644 = ~pi96 & n643;
  assign n645 = ~n642 & ~n644;
  assign n646 = pi100 & ~n645;
  assign n647 = pi25 & ~pi116;
  assign n648 = pi85 & n647;
  assign n649 = ~n646 & ~n648;
  assign n650 = ~pi26 & ~n649;
  assign n651 = ~pi95 & ~pi100;
  assign n652 = ~pi97 & n651;
  assign n653 = ~pi110 & ~n652;
  assign n654 = pi25 & ~n653;
  assign n655 = pi26 & pi116;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~pi39 & ~pi52;
  assign n658 = ~pi51 & n657;
  assign n659 = ~n656 & ~n658;
  assign n660 = pi26 & n647;
  assign n661 = ~n659 & ~n660;
  assign n662 = ~pi85 & ~n661;
  assign n663 = ~n650 & ~n662;
  assign n664 = ~pi27 & ~n663;
  assign n665 = pi116 & n658;
  assign n666 = ~n647 & ~n665;
  assign n667 = pi27 & ~n666;
  assign n668 = n654 & n658;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~pi26 & ~pi85;
  assign n671 = ~n669 & n670;
  assign n672 = ~n664 & ~n671;
  assign n673 = ~pi53 & ~n672;
  assign n674 = ~pi26 & n647;
  assign n675 = pi53 & ~pi85;
  assign n676 = ~pi27 & n675;
  assign n677 = n674 & n676;
  assign n678 = ~n673 & ~n677;
  assign n679 = ~pi58 & ~n678;
  assign n680 = ~pi27 & ~pi85;
  assign n681 = ~pi53 & pi58;
  assign n682 = n680 & n681;
  assign n683 = n674 & n682;
  assign n684 = ~n679 & ~n683;
  assign po40 = n339 & ~n684;
  assign n686 = pi100 & ~n655;
  assign n687 = ~n645 & n686;
  assign n688 = ~pi85 & ~n665;
  assign n689 = pi26 & n688;
  assign n690 = ~n687 & ~n689;
  assign n691 = ~pi53 & ~pi58;
  assign n692 = ~pi27 & n691;
  assign n693 = n339 & n692;
  assign po41 = ~n690 & n693;
  assign n695 = pi85 & ~pi116;
  assign n696 = pi95 & ~pi96;
  assign n697 = pi27 & pi116;
  assign n698 = ~pi110 & ~n695;
  assign n699 = n696 & ~n697;
  assign n700 = n698 & n699;
  assign n701 = ~pi27 & n642;
  assign n702 = ~n700 & ~n701;
  assign n703 = ~pi100 & ~n702;
  assign n704 = pi27 & n688;
  assign n705 = ~n703 & ~n704;
  assign n706 = ~pi26 & n691;
  assign n707 = n339 & n706;
  assign po42 = ~n705 & n707;
  assign n709 = ~pi26 & ~n658;
  assign n710 = ~pi27 & n658;
  assign n711 = ~n709 & ~n710;
  assign n712 = ~n653 & ~n711;
  assign n713 = pi26 & ~pi27;
  assign n714 = ~pi26 & pi27;
  assign n715 = ~n713 & ~n714;
  assign n716 = ~pi116 & ~n715;
  assign n717 = ~n712 & ~n716;
  assign n718 = pi28 & ~n717;
  assign n719 = ~pi26 & ~pi100;
  assign n720 = ~pi110 & n719;
  assign n721 = n696 & n720;
  assign n722 = n655 & n658;
  assign n723 = ~n721 & ~n722;
  assign n724 = ~pi27 & ~n723;
  assign n725 = n697 & n709;
  assign n726 = ~n724 & ~n725;
  assign n727 = ~n718 & n726;
  assign n728 = ~pi85 & ~n727;
  assign n729 = pi28 & ~pi116;
  assign n730 = ~pi100 & pi116;
  assign n731 = ~n729 & ~n730;
  assign n732 = ~pi26 & ~pi27;
  assign n733 = pi85 & n732;
  assign n734 = ~n731 & n733;
  assign n735 = ~n728 & ~n734;
  assign n736 = ~pi53 & ~n735;
  assign n737 = ~pi27 & pi28;
  assign n738 = ~pi116 & n737;
  assign n739 = ~pi26 & n675;
  assign n740 = n738 & n739;
  assign n741 = ~n736 & ~n740;
  assign n742 = ~pi58 & ~n741;
  assign n743 = n670 & n681;
  assign n744 = n738 & n743;
  assign n745 = ~n742 & ~n744;
  assign po43 = n339 & ~n745;
  assign n747 = pi29 & pi110;
  assign n748 = ~pi96 & pi97;
  assign n749 = ~pi110 & n748;
  assign n750 = pi29 & ~pi97;
  assign n751 = ~n749 & ~n750;
  assign n752 = n651 & ~n751;
  assign n753 = ~n747 & ~n752;
  assign n754 = ~pi58 & ~n753;
  assign n755 = pi97 & pi116;
  assign n756 = pi29 & ~pi116;
  assign n757 = ~n755 & ~n756;
  assign n758 = pi58 & ~n757;
  assign n759 = ~n754 & ~n758;
  assign n760 = ~pi53 & ~n759;
  assign n761 = pi53 & ~pi58;
  assign n762 = n756 & n761;
  assign n763 = ~n760 & ~n762;
  assign n764 = ~pi27 & ~n763;
  assign n765 = pi27 & n691;
  assign n766 = n756 & n765;
  assign n767 = ~n764 & ~n766;
  assign n768 = ~pi85 & ~n767;
  assign n769 = pi85 & n756;
  assign n770 = n692 & n769;
  assign n771 = ~n768 & ~n770;
  assign n772 = ~pi26 & ~n771;
  assign n773 = ~pi85 & n691;
  assign n774 = n713 & n773;
  assign n775 = n756 & n774;
  assign n776 = ~n772 & ~n775;
  assign po44 = n339 & ~n776;
  assign n778 = pi30 & ~pi109;
  assign n779 = pi60 & pi109;
  assign n780 = ~n778 & ~n779;
  assign n781 = ~pi106 & ~n780;
  assign n782 = pi88 & pi106;
  assign n783 = ~n781 & ~n782;
  assign po45 = ~pi129 & ~n783;
  assign n785 = pi89 & pi106;
  assign n786 = pi30 & pi109;
  assign n787 = pi31 & ~pi109;
  assign n788 = ~n786 & ~n787;
  assign n789 = ~pi106 & ~n788;
  assign n790 = ~n785 & ~n789;
  assign po46 = ~pi129 & ~n790;
  assign n792 = pi99 & pi106;
  assign n793 = pi31 & pi109;
  assign n794 = pi32 & ~pi109;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~pi106 & ~n795;
  assign n797 = ~n792 & ~n796;
  assign po47 = ~pi129 & ~n797;
  assign n799 = pi90 & pi106;
  assign n800 = pi32 & pi109;
  assign n801 = pi33 & ~pi109;
  assign n802 = ~n800 & ~n801;
  assign n803 = ~pi106 & ~n802;
  assign n804 = ~n799 & ~n803;
  assign po48 = ~pi129 & ~n804;
  assign n806 = pi91 & pi106;
  assign n807 = pi33 & pi109;
  assign n808 = pi34 & ~pi109;
  assign n809 = ~n807 & ~n808;
  assign n810 = ~pi106 & ~n809;
  assign n811 = ~n806 & ~n810;
  assign po49 = ~pi129 & ~n811;
  assign n813 = pi92 & pi106;
  assign n814 = pi34 & pi109;
  assign n815 = pi35 & ~pi109;
  assign n816 = ~n814 & ~n815;
  assign n817 = ~pi106 & ~n816;
  assign n818 = ~n813 & ~n817;
  assign po50 = ~pi129 & ~n818;
  assign n820 = pi98 & pi106;
  assign n821 = pi35 & pi109;
  assign n822 = pi36 & ~pi109;
  assign n823 = ~n821 & ~n822;
  assign n824 = ~pi106 & ~n823;
  assign n825 = ~n820 & ~n824;
  assign po51 = ~pi129 & ~n825;
  assign n827 = pi93 & pi106;
  assign n828 = pi36 & pi109;
  assign n829 = pi37 & ~pi109;
  assign n830 = ~n828 & ~n829;
  assign n831 = ~pi106 & ~n830;
  assign n832 = ~n827 & ~n831;
  assign po52 = ~pi129 & ~n832;
  assign n834 = pi82 & ~n389;
  assign n835 = n380 & n382;
  assign n836 = n525 & n835;
  assign n837 = pi82 & ~n836;
  assign n838 = n394 & ~n837;
  assign n839 = ~n834 & ~n838;
  assign n840 = ~pi38 & ~n839;
  assign n841 = ~pi48 & n835;
  assign n842 = n583 & n841;
  assign n843 = ~pi50 & n389;
  assign n844 = n842 & n843;
  assign n845 = pi82 & ~n844;
  assign n846 = pi74 & ~n394;
  assign n847 = ~n845 & n846;
  assign n848 = ~pi40 & ~pi42;
  assign n849 = ~pi44 & pi82;
  assign n850 = n848 & n849;
  assign n851 = pi38 & n850;
  assign n852 = ~pi129 & ~n851;
  assign n853 = ~n840 & n852;
  assign po53 = ~n847 & n853;
  assign n855 = ~pi51 & ~pi52;
  assign n856 = pi109 & n855;
  assign n857 = pi39 & ~n856;
  assign n858 = ~pi51 & pi109;
  assign n859 = n657 & n858;
  assign n860 = ~pi106 & ~n859;
  assign n861 = ~n857 & n860;
  assign po54 = ~pi129 & ~n861;
  assign n863 = pi82 & ~n388;
  assign n864 = n524 & n835;
  assign n865 = n387 & n864;
  assign n866 = pi82 & ~n865;
  assign n867 = n394 & ~n866;
  assign n868 = ~n863 & ~n867;
  assign n869 = ~pi40 & ~n868;
  assign n870 = pi73 & ~n394;
  assign n871 = ~n863 & n870;
  assign n872 = ~n866 & n871;
  assign n873 = n834 & ~n863;
  assign n874 = ~pi129 & ~n873;
  assign n875 = ~n872 & n874;
  assign po55 = ~n869 & n875;
  assign n877 = pi82 & ~n538;
  assign n878 = pi82 & ~n864;
  assign n879 = n394 & ~n878;
  assign n880 = ~n877 & ~n879;
  assign n881 = ~pi41 & ~n880;
  assign n882 = pi76 & ~n394;
  assign n883 = ~n877 & n882;
  assign n884 = ~n878 & n883;
  assign n885 = pi41 & pi82;
  assign n886 = n538 & n885;
  assign n887 = ~pi129 & ~n886;
  assign n888 = ~n884 & n887;
  assign po56 = ~n881 & n888;
  assign n890 = pi44 & pi82;
  assign n891 = n541 & n841;
  assign n892 = n397 & n399;
  assign n893 = n891 & n892;
  assign n894 = pi82 & ~n893;
  assign n895 = n394 & ~n894;
  assign n896 = ~n890 & ~n895;
  assign n897 = ~pi42 & ~n896;
  assign n898 = ~pi44 & ~pi50;
  assign n899 = n397 & n898;
  assign n900 = n842 & n899;
  assign n901 = pi82 & ~n900;
  assign n902 = pi72 & ~n394;
  assign n903 = ~n901 & n902;
  assign n904 = pi42 & n849;
  assign n905 = ~pi129 & ~n904;
  assign n906 = ~n903 & n905;
  assign po57 = ~n897 & n906;
  assign n908 = pi82 & ~n401;
  assign n909 = pi82 & ~n384;
  assign n910 = n394 & ~n909;
  assign n911 = ~n908 & ~n910;
  assign n912 = ~pi43 & ~n911;
  assign n913 = pi77 & ~n394;
  assign n914 = ~n908 & n913;
  assign n915 = ~n909 & n914;
  assign n916 = pi43 & n387;
  assign n917 = n850 & n916;
  assign n918 = ~pi129 & ~n917;
  assign n919 = ~n915 & n918;
  assign po58 = ~n912 & n919;
  assign n921 = ~pi38 & n848;
  assign n922 = n836 & n921;
  assign n923 = pi82 & ~n922;
  assign n924 = pi67 & ~n394;
  assign n925 = ~pi44 & n394;
  assign n926 = ~n924 & ~n925;
  assign n927 = ~n923 & ~n926;
  assign n928 = ~pi129 & ~n890;
  assign po59 = ~n927 & n928;
  assign n930 = ~pi2 & n381;
  assign n931 = n380 & n930;
  assign n932 = n402 & n931;
  assign n933 = pi82 & ~n932;
  assign n934 = pi68 & ~n394;
  assign n935 = ~n933 & n934;
  assign n936 = pi82 & ~n526;
  assign n937 = n394 & ~n636;
  assign n938 = ~n632 & n937;
  assign n939 = ~n936 & ~n938;
  assign n940 = ~pi45 & ~n939;
  assign n941 = pi45 & n849;
  assign n942 = n921 & n941;
  assign n943 = n525 & n942;
  assign n944 = ~pi129 & ~n943;
  assign n945 = ~n935 & n944;
  assign po60 = ~n940 & n945;
  assign n947 = pi82 & ~n587;
  assign n948 = pi82 & ~n891;
  assign n949 = n394 & ~n948;
  assign n950 = ~n947 & ~n949;
  assign n951 = ~pi46 & ~n950;
  assign n952 = pi75 & ~n394;
  assign n953 = ~n947 & n952;
  assign n954 = ~n948 & n953;
  assign n955 = pi46 & pi82;
  assign n956 = n587 & n955;
  assign n957 = ~pi129 & ~n956;
  assign n958 = ~n954 & n957;
  assign po61 = ~n951 & n958;
  assign n960 = pi82 & ~n402;
  assign n961 = pi82 & ~n841;
  assign n962 = n394 & ~n961;
  assign n963 = ~n960 & ~n962;
  assign n964 = ~pi47 & ~n963;
  assign n965 = pi64 & ~n394;
  assign n966 = ~n960 & n965;
  assign n967 = ~n961 & n966;
  assign n968 = pi47 & n540;
  assign n969 = n537 & n968;
  assign n970 = n850 & n969;
  assign n971 = ~pi129 & ~n970;
  assign n972 = ~n967 & n971;
  assign po62 = ~n964 & n972;
  assign n974 = ~pi47 & n835;
  assign n975 = n402 & n974;
  assign n976 = pi82 & ~n975;
  assign n977 = pi62 & ~n394;
  assign n978 = ~n976 & n977;
  assign n979 = n583 & n587;
  assign n980 = pi82 & ~n979;
  assign n981 = pi82 & ~n835;
  assign n982 = n394 & ~n981;
  assign n983 = ~n980 & ~n982;
  assign n984 = ~pi48 & ~n983;
  assign n985 = pi48 & n523;
  assign n986 = n849 & n985;
  assign n987 = n400 & n921;
  assign n988 = n986 & n987;
  assign n989 = ~pi129 & ~n988;
  assign n990 = ~n978 & n989;
  assign po63 = ~n984 & n990;
  assign n992 = n585 & n587;
  assign n993 = pi49 & ~n992;
  assign n994 = n379 & n587;
  assign n995 = ~pi2 & n378;
  assign n996 = n584 & ~n995;
  assign n997 = n994 & n996;
  assign n998 = ~n993 & ~n997;
  assign n999 = pi82 & ~n998;
  assign n1000 = n584 & n994;
  assign n1001 = pi82 & ~n1000;
  assign n1002 = ~pi69 & ~n394;
  assign n1003 = ~n1001 & n1002;
  assign n1004 = pi49 & n407;
  assign n1005 = ~n1003 & ~n1004;
  assign n1006 = ~n999 & n1005;
  assign po64 = ~pi129 & ~n1006;
  assign n1008 = pi82 & ~n398;
  assign n1009 = pi82 & ~n842;
  assign n1010 = n394 & ~n1009;
  assign n1011 = ~n1008 & ~n1010;
  assign n1012 = ~pi50 & ~n1011;
  assign n1013 = pi66 & ~n394;
  assign n1014 = ~n1008 & n1013;
  assign n1015 = ~n1009 & n1014;
  assign n1016 = pi50 & n849;
  assign n1017 = n921 & n1016;
  assign n1018 = ~pi129 & ~n1017;
  assign n1019 = ~n1015 & n1018;
  assign po65 = ~n1012 & n1019;
  assign n1021 = pi51 & ~pi109;
  assign n1022 = ~pi106 & ~n858;
  assign n1023 = ~n1021 & n1022;
  assign po66 = ~pi129 & ~n1023;
  assign n1025 = pi52 & ~n858;
  assign n1026 = ~pi106 & ~n856;
  assign n1027 = ~n1025 & n1026;
  assign po67 = ~pi129 & ~n1027;
  assign n1029 = pi58 & pi116;
  assign n1030 = ~pi58 & ~pi96;
  assign n1031 = ~pi110 & n1030;
  assign n1032 = n651 & n1031;
  assign n1033 = ~n1029 & ~n1032;
  assign n1034 = ~pi53 & pi97;
  assign n1035 = ~n1033 & n1034;
  assign n1036 = ~pi116 & n761;
  assign n1037 = ~n1035 & ~n1036;
  assign n1038 = ~pi26 & n339;
  assign n1039 = n680 & n1038;
  assign po68 = ~n1037 & n1039;
  assign n1041 = ~n394 & ~n909;
  assign n1042 = ~n960 & n1041;
  assign po69 = pi129 | n1042;
  assign po129 = pi123 | pi129;
  assign n1045 = pi114 & ~pi122;
  assign po70 = ~po129 & n1045;
  assign n1047 = ~pi26 & pi58;
  assign n1048 = ~pi58 & n655;
  assign n1049 = ~n1047 & ~n1048;
  assign n1050 = pi94 & ~n1049;
  assign n1051 = pi58 & ~pi116;
  assign n1052 = pi37 & ~pi116;
  assign n1053 = ~n1047 & ~n1052;
  assign n1054 = ~n1051 & ~n1053;
  assign n1055 = ~n1050 & ~n1054;
  assign n1056 = ~pi53 & ~n1055;
  assign n1057 = ~pi26 & pi37;
  assign n1058 = ~pi58 & n1057;
  assign n1059 = ~n1056 & ~n1058;
  assign n1060 = ~pi85 & ~n1059;
  assign n1061 = n691 & n1057;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~pi27 & ~n1062;
  assign n1064 = n773 & n1057;
  assign n1065 = ~n1063 & ~n1064;
  assign po71 = n339 & ~n1065;
  assign n1067 = ~pi26 & ~pi53;
  assign n1068 = ~pi53 & ~pi85;
  assign n1069 = ~n670 & ~n1067;
  assign n1070 = ~n1068 & n1069;
  assign n1071 = ~pi58 & ~n1070;
  assign n1072 = ~pi85 & n1067;
  assign n1073 = ~pi116 & n1072;
  assign n1074 = ~n1071 & ~n1073;
  assign n1075 = pi57 & ~n1074;
  assign n1076 = pi60 & n1029;
  assign n1077 = n1072 & n1076;
  assign n1078 = ~n1075 & ~n1077;
  assign n1079 = ~pi27 & ~n1078;
  assign n1080 = pi57 & ~pi58;
  assign n1081 = n1072 & n1080;
  assign n1082 = ~n1079 & ~n1081;
  assign po72 = n339 & ~n1082;
  assign n1084 = n732 & n1051;
  assign n1085 = ~pi58 & pi116;
  assign n1086 = n658 & n1085;
  assign n1087 = ~n715 & n1086;
  assign n1088 = ~n1084 & ~n1087;
  assign n1089 = n339 & n1068;
  assign po73 = ~n1088 & n1089;
  assign n1091 = ~n681 & ~n761;
  assign n1092 = ~pi116 & ~n1091;
  assign n1093 = ~n653 & n691;
  assign n1094 = ~n1092 & ~n1093;
  assign n1095 = pi59 & ~n1094;
  assign n1096 = pi96 & n691;
  assign n1097 = n653 & n1096;
  assign n1098 = ~n1095 & ~n1097;
  assign n1099 = ~pi85 & ~n1098;
  assign n1100 = pi59 & ~pi116;
  assign n1101 = pi85 & n691;
  assign n1102 = n1100 & n1101;
  assign n1103 = ~n1099 & ~n1102;
  assign n1104 = ~pi27 & ~n1103;
  assign n1105 = pi27 & n1100;
  assign n1106 = n773 & n1105;
  assign n1107 = ~n1104 & ~n1106;
  assign n1108 = ~pi26 & ~n1107;
  assign n1109 = n774 & n1100;
  assign n1110 = ~n1108 & ~n1109;
  assign po74 = n339 & ~n1110;
  assign n1112 = ~pi117 & ~pi122;
  assign n1113 = pi60 & ~n1112;
  assign n1114 = pi123 & n1112;
  assign po75 = n1113 | n1114;
  assign n1116 = ~pi114 & ~pi122;
  assign n1117 = pi123 & ~pi129;
  assign po76 = n1116 & n1117;
  assign n1119 = pi136 & ~pi137;
  assign n1120 = pi131 & pi132;
  assign n1121 = pi133 & n1120;
  assign n1122 = ~pi138 & n1121;
  assign n1123 = n1119 & n1122;
  assign n1124 = pi62 & ~n1123;
  assign n1125 = ~pi140 & n1119;
  assign n1126 = n1122 & n1125;
  assign n1127 = ~n1124 & ~n1126;
  assign po77 = pi129 | n1127;
  assign n1129 = pi63 & ~n1123;
  assign n1130 = ~pi142 & n1119;
  assign n1131 = n1122 & n1130;
  assign n1132 = ~n1129 & ~n1131;
  assign po78 = pi129 | n1132;
  assign n1134 = pi64 & ~n1123;
  assign n1135 = ~pi139 & n1119;
  assign n1136 = n1122 & n1135;
  assign n1137 = ~n1134 & ~n1136;
  assign po79 = pi129 | n1137;
  assign n1139 = pi65 & ~n1123;
  assign n1140 = ~pi146 & n1119;
  assign n1141 = n1122 & n1140;
  assign n1142 = ~n1139 & ~n1141;
  assign po80 = pi129 | n1142;
  assign n1144 = ~pi136 & ~pi137;
  assign n1145 = n1122 & n1144;
  assign n1146 = pi66 & ~n1145;
  assign n1147 = ~pi143 & n1145;
  assign n1148 = ~n1146 & ~n1147;
  assign po81 = pi129 | n1148;
  assign n1150 = pi67 & ~n1145;
  assign n1151 = ~pi139 & n1145;
  assign n1152 = ~n1150 & ~n1151;
  assign po82 = pi129 | n1152;
  assign n1154 = pi68 & ~n1123;
  assign n1155 = ~pi141 & n1119;
  assign n1156 = n1122 & n1155;
  assign n1157 = ~n1154 & ~n1156;
  assign po83 = pi129 | n1157;
  assign n1159 = pi69 & ~n1123;
  assign n1160 = ~pi143 & n1119;
  assign n1161 = n1122 & n1160;
  assign n1162 = ~n1159 & ~n1161;
  assign po84 = pi129 | n1162;
  assign n1164 = pi70 & ~n1123;
  assign n1165 = ~pi144 & n1119;
  assign n1166 = n1122 & n1165;
  assign n1167 = ~n1164 & ~n1166;
  assign po85 = pi129 | n1167;
  assign n1169 = pi71 & ~n1123;
  assign n1170 = ~pi145 & n1119;
  assign n1171 = n1122 & n1170;
  assign n1172 = ~n1169 & ~n1171;
  assign po86 = pi129 | n1172;
  assign n1174 = pi72 & ~n1145;
  assign n1175 = ~pi140 & n1145;
  assign n1176 = ~n1174 & ~n1175;
  assign po87 = pi129 | n1176;
  assign n1178 = pi73 & ~n1145;
  assign n1179 = ~pi141 & n1145;
  assign n1180 = ~n1178 & ~n1179;
  assign po88 = pi129 | n1180;
  assign n1182 = pi74 & ~n1145;
  assign n1183 = ~pi142 & n1145;
  assign n1184 = ~n1182 & ~n1183;
  assign po89 = pi129 | n1184;
  assign n1186 = pi75 & ~n1145;
  assign n1187 = ~pi144 & n1145;
  assign n1188 = ~n1186 & ~n1187;
  assign po90 = pi129 | n1188;
  assign n1190 = pi76 & ~n1145;
  assign n1191 = ~pi145 & n1145;
  assign n1192 = ~n1190 & ~n1191;
  assign po91 = pi129 | n1192;
  assign n1194 = pi77 & ~n1145;
  assign n1195 = ~pi146 & n1145;
  assign n1196 = ~n1194 & ~n1195;
  assign po92 = pi129 | n1196;
  assign n1198 = ~pi136 & pi137;
  assign n1199 = n1122 & n1198;
  assign n1200 = pi78 & ~n1199;
  assign n1201 = pi142 & n1199;
  assign n1202 = ~n1200 & ~n1201;
  assign po93 = ~pi129 & ~n1202;
  assign n1204 = pi79 & ~n1199;
  assign n1205 = pi143 & n1199;
  assign n1206 = ~n1204 & ~n1205;
  assign po94 = ~pi129 & ~n1206;
  assign n1208 = pi80 & ~n1199;
  assign n1209 = pi144 & n1199;
  assign n1210 = ~n1208 & ~n1209;
  assign po95 = ~pi129 & ~n1210;
  assign n1212 = pi81 & ~n1199;
  assign n1213 = pi145 & n1199;
  assign n1214 = ~n1212 & ~n1213;
  assign po96 = ~pi129 & ~n1214;
  assign n1216 = pi82 & ~n1199;
  assign n1217 = pi146 & n1199;
  assign n1218 = ~n1216 & ~n1217;
  assign po97 = ~pi129 & ~n1218;
  assign n1220 = pi89 & pi138;
  assign n1221 = ~pi62 & ~pi138;
  assign n1222 = ~n1220 & ~n1221;
  assign n1223 = pi136 & ~n1222;
  assign n1224 = pi119 & pi138;
  assign n1225 = ~pi72 & ~pi138;
  assign n1226 = ~n1224 & ~n1225;
  assign n1227 = ~pi136 & ~n1226;
  assign n1228 = ~n1223 & ~n1227;
  assign n1229 = ~pi137 & ~n1228;
  assign n1230 = ~pi115 & pi138;
  assign n1231 = pi87 & ~pi138;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = ~pi136 & ~n1232;
  assign n1234 = pi136 & ~pi138;
  assign n1235 = pi31 & n1234;
  assign n1236 = ~n1233 & ~n1235;
  assign n1237 = pi137 & ~n1236;
  assign po98 = n1229 | n1237;
  assign n1239 = pi84 & ~n1199;
  assign n1240 = pi141 & n1199;
  assign n1241 = ~n1239 & ~n1240;
  assign po99 = ~pi129 & ~n1241;
  assign n1243 = n643 & ~n652;
  assign n1244 = pi96 & n1243;
  assign n1245 = ~n695 & ~n1244;
  assign n1246 = n692 & n1038;
  assign po100 = ~n1245 & n1246;
  assign n1248 = pi86 & ~n1199;
  assign n1249 = pi139 & n1199;
  assign n1250 = ~n1248 & ~n1249;
  assign po101 = ~pi129 & ~n1250;
  assign n1252 = pi87 & ~n1199;
  assign n1253 = pi140 & n1199;
  assign n1254 = ~n1252 & ~n1253;
  assign po102 = ~pi129 & ~n1254;
  assign n1256 = pi136 & pi137;
  assign n1257 = n1122 & n1256;
  assign n1258 = pi88 & ~n1257;
  assign n1259 = pi139 & n1257;
  assign n1260 = ~n1258 & ~n1259;
  assign po103 = ~pi129 & ~n1260;
  assign n1262 = pi89 & ~n1257;
  assign n1263 = pi140 & n1257;
  assign n1264 = ~n1262 & ~n1263;
  assign po104 = ~pi129 & ~n1264;
  assign n1266 = pi90 & ~n1257;
  assign n1267 = pi142 & n1257;
  assign n1268 = ~n1266 & ~n1267;
  assign po105 = ~pi129 & ~n1268;
  assign n1270 = pi91 & ~n1257;
  assign n1271 = pi143 & n1257;
  assign n1272 = ~n1270 & ~n1271;
  assign po106 = ~pi129 & ~n1272;
  assign n1274 = pi92 & ~n1257;
  assign n1275 = pi144 & n1257;
  assign n1276 = ~n1274 & ~n1275;
  assign po107 = ~pi129 & ~n1276;
  assign n1278 = pi93 & ~n1257;
  assign n1279 = pi146 & n1257;
  assign n1280 = ~n1278 & ~n1279;
  assign po108 = ~pi129 & ~n1280;
  assign n1282 = pi82 & pi138;
  assign n1283 = n1144 & n1282;
  assign n1284 = n1121 & n1283;
  assign n1285 = pi94 & ~n1284;
  assign n1286 = pi142 & n1284;
  assign n1287 = ~n1285 & ~n1286;
  assign po109 = ~pi129 & ~n1287;
  assign n1289 = ~pi3 & ~pi110;
  assign n1290 = ~n1121 & n1289;
  assign n1291 = n1121 & ~n1283;
  assign n1292 = ~n1290 & ~n1291;
  assign n1293 = pi95 & ~n1292;
  assign n1294 = pi143 & n1284;
  assign n1295 = ~n1293 & ~n1294;
  assign po110 = ~pi129 & ~n1295;
  assign n1297 = pi96 & ~n1292;
  assign n1298 = pi146 & n1284;
  assign n1299 = ~n1297 & ~n1298;
  assign po111 = ~pi129 & ~n1299;
  assign n1301 = pi97 & ~n1292;
  assign n1302 = pi145 & n1284;
  assign n1303 = ~n1301 & ~n1302;
  assign po112 = ~pi129 & ~n1303;
  assign n1305 = pi98 & ~n1257;
  assign n1306 = pi145 & n1257;
  assign n1307 = ~n1305 & ~n1306;
  assign po113 = ~pi129 & ~n1307;
  assign n1309 = pi99 & ~n1257;
  assign n1310 = pi141 & n1257;
  assign n1311 = ~n1309 & ~n1310;
  assign po114 = ~pi129 & ~n1311;
  assign n1313 = pi100 & ~n1292;
  assign n1314 = pi144 & n1284;
  assign n1315 = ~n1313 & ~n1314;
  assign po115 = ~pi129 & ~n1315;
  assign n1317 = pi124 & pi138;
  assign n1318 = ~pi77 & ~pi138;
  assign n1319 = ~n1317 & ~n1318;
  assign n1320 = ~pi136 & ~n1319;
  assign n1321 = ~pi65 & ~pi138;
  assign n1322 = pi93 & pi138;
  assign n1323 = ~n1321 & ~n1322;
  assign n1324 = pi136 & ~n1323;
  assign n1325 = ~n1320 & ~n1324;
  assign n1326 = ~pi137 & ~n1325;
  assign n1327 = pi37 & n1234;
  assign n1328 = pi96 & pi138;
  assign n1329 = pi82 & ~pi138;
  assign n1330 = ~n1328 & ~n1329;
  assign n1331 = ~pi136 & ~n1330;
  assign n1332 = ~n1327 & ~n1331;
  assign n1333 = pi137 & ~n1332;
  assign po116 = n1326 | n1333;
  assign n1335 = pi91 & n1119;
  assign n1336 = pi95 & n1198;
  assign n1337 = ~n1335 & ~n1336;
  assign n1338 = pi138 & ~n1337;
  assign n1339 = pi79 & ~pi136;
  assign n1340 = pi34 & pi136;
  assign n1341 = ~n1339 & ~n1340;
  assign n1342 = pi137 & ~n1341;
  assign n1343 = ~pi69 & pi136;
  assign n1344 = ~pi66 & ~pi136;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = ~pi137 & ~n1345;
  assign n1347 = ~n1342 & ~n1346;
  assign n1348 = ~pi138 & ~n1347;
  assign po117 = n1338 | n1348;
  assign n1350 = pi90 & n1119;
  assign n1351 = pi94 & n1198;
  assign n1352 = ~n1350 & ~n1351;
  assign n1353 = pi138 & ~n1352;
  assign n1354 = pi78 & ~pi136;
  assign n1355 = pi33 & pi136;
  assign n1356 = ~n1354 & ~n1355;
  assign n1357 = pi137 & ~n1356;
  assign n1358 = ~pi63 & pi136;
  assign n1359 = ~pi74 & ~pi136;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = ~pi137 & ~n1360;
  assign n1362 = ~n1357 & ~n1361;
  assign n1363 = ~pi138 & ~n1362;
  assign po118 = n1353 | n1363;
  assign n1365 = pi99 & n1119;
  assign n1366 = ~pi112 & n1198;
  assign n1367 = ~n1365 & ~n1366;
  assign n1368 = pi138 & ~n1367;
  assign n1369 = ~pi68 & pi136;
  assign n1370 = ~pi73 & ~pi136;
  assign n1371 = ~n1369 & ~n1370;
  assign n1372 = ~pi137 & ~n1371;
  assign n1373 = pi84 & ~pi136;
  assign n1374 = pi32 & pi136;
  assign n1375 = ~n1373 & ~n1374;
  assign n1376 = pi137 & ~n1375;
  assign n1377 = ~n1372 & ~n1376;
  assign n1378 = ~pi138 & ~n1377;
  assign po119 = n1368 | n1378;
  assign n1380 = pi92 & pi138;
  assign n1381 = ~pi70 & ~pi138;
  assign n1382 = ~n1380 & ~n1381;
  assign n1383 = pi136 & ~n1382;
  assign n1384 = pi125 & pi138;
  assign n1385 = ~pi75 & ~pi138;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = ~pi136 & ~n1386;
  assign n1388 = ~n1383 & ~n1387;
  assign n1389 = ~pi137 & ~n1388;
  assign n1390 = pi80 & ~pi138;
  assign n1391 = pi100 & pi138;
  assign n1392 = ~n1390 & ~n1391;
  assign n1393 = ~pi136 & ~n1392;
  assign n1394 = pi35 & n1234;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = pi137 & ~n1395;
  assign po120 = n1389 | n1396;
  assign n1398 = ~pi27 & n706;
  assign n1399 = n1243 & n1398;
  assign n1400 = ~n642 & ~n1399;
  assign po121 = n339 & ~n1400;
  assign n1402 = pi98 & pi138;
  assign n1403 = ~pi71 & ~pi138;
  assign n1404 = ~n1402 & ~n1403;
  assign n1405 = pi136 & ~n1404;
  assign n1406 = ~pi76 & ~pi138;
  assign n1407 = pi23 & pi138;
  assign n1408 = ~n1406 & ~n1407;
  assign n1409 = ~pi136 & ~n1408;
  assign n1410 = ~n1405 & ~n1409;
  assign n1411 = ~pi137 & ~n1410;
  assign n1412 = pi36 & n1234;
  assign n1413 = pi81 & ~pi138;
  assign n1414 = pi97 & pi138;
  assign n1415 = ~n1413 & ~n1414;
  assign n1416 = ~pi136 & ~n1415;
  assign n1417 = ~n1412 & ~n1416;
  assign n1418 = pi137 & ~n1417;
  assign po122 = n1411 | n1418;
  assign n1420 = pi88 & pi138;
  assign n1421 = ~pi64 & ~pi138;
  assign n1422 = ~n1420 & ~n1421;
  assign n1423 = pi136 & ~n1422;
  assign n1424 = pi120 & pi138;
  assign n1425 = ~pi67 & ~pi138;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = ~pi136 & ~n1426;
  assign n1428 = ~n1423 & ~n1427;
  assign n1429 = ~pi137 & ~n1428;
  assign n1430 = pi86 & ~pi138;
  assign n1431 = pi111 & pi138;
  assign n1432 = ~n1430 & ~n1431;
  assign n1433 = ~pi136 & ~n1432;
  assign n1434 = pi30 & n1234;
  assign n1435 = ~n1433 & ~n1434;
  assign n1436 = pi137 & ~n1435;
  assign po123 = n1429 | n1436;
  assign n1438 = ~n658 & n714;
  assign n1439 = ~n713 & ~n1438;
  assign n1440 = pi116 & n339;
  assign po124 = ~n1439 & n1440;
  assign n1442 = ~pi97 & n681;
  assign n1443 = ~n761 & ~n1442;
  assign po125 = n1440 & ~n1443;
  assign n1445 = pi111 & ~n1283;
  assign n1446 = pi139 & n1283;
  assign n1447 = ~n1445 & ~n1446;
  assign n1448 = ~pi129 & n1121;
  assign po126 = ~n1447 & n1448;
  assign n1450 = ~pi112 & ~n1283;
  assign n1451 = pi141 & n1283;
  assign n1452 = ~n1450 & ~n1451;
  assign po127 = n1448 & ~n1452;
  assign n1454 = ~pi54 & ~pi113;
  assign n1455 = ~pi11 & ~pi22;
  assign n1456 = pi54 & ~n1455;
  assign n1457 = ~n1454 & ~n1456;
  assign po128 = n339 & ~n1457;
  assign n1459 = ~pi115 & ~n1283;
  assign n1460 = pi140 & n1283;
  assign n1461 = ~n1459 & ~n1460;
  assign po130 = n1448 & ~n1461;
  assign n1463 = ~pi4 & ~pi7;
  assign n1464 = ~pi9 & ~pi12;
  assign n1465 = n1463 & n1464;
  assign n1466 = pi54 & n339;
  assign po131 = ~n1465 & n1466;
  assign po132 = ~pi122 | pi129;
  assign n1469 = ~pi54 & pi118;
  assign n1470 = pi54 & ~pi59;
  assign n1471 = n508 & n1470;
  assign n1472 = ~n1469 & ~n1471;
  assign po133 = ~pi129 & ~n1472;
  assign po134 = ~pi129 & ~n651;
  assign n1475 = ~pi120 & n1289;
  assign n1476 = ~pi111 & ~pi129;
  assign po135 = ~n1475 & n1476;
  assign n1478 = pi81 & pi120;
  assign po136 = ~pi129 & n1478;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi57 & ~pi129;
  assign n1483 = ~pi96 & pi125;
  assign n1484 = ~pi3 & ~n1483;
  assign po140 = ~pi129 & ~n1484;
  assign n1486 = ~pi126 & pi132;
  assign po141 = pi133 & n1486;
  assign po12 = 1'b1;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
endmodule
