module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n182, n183, n184,
    n185, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n196, n197, n198,
    n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212,
    n213, n214, n215, n216, n217, n218, n219,
    n220, n221, n222, n223, n224, n225, n226,
    n227, n228, n229, n230, n231, n232, n233,
    n234, n235, n236, n237, n238, n239, n240,
    n241, n242, n243, n244, n245, n246, n247,
    n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261,
    n262, n263, n264, n265, n266, n267, n268,
    n269, n270, n271, n272, n273, n274, n275,
    n276, n277, n278, n279, n280, n281, n282,
    n283, n284, n285, n286, n287, n288, n289,
    n290, n291, n292, n293, n294, n295, n296,
    n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310,
    n311, n312, n313, n314, n315, n316, n317,
    n318, n319, n320, n321, n322, n323, n324,
    n325, n326, n327, n328, n329, n330, n331,
    n332, n333, n334, n335, n336, n337, n338,
    n339, n340, n341, n342, n343, n344, n345,
    n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359,
    n360, n361, n362, n363, n364, n365, n366,
    n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380,
    n381, n382, n383, n384, n385, n386, n387,
    n388, n389, n390, n391, n392, n393, n394,
    n395, n396, n397, n398, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408,
    n409, n410, n411, n412, n413, n414, n415,
    n416, n417, n418, n419, n420, n421, n422,
    n423, n424, n425, n426, n427, n428, n429,
    n430, n431, n432, n433, n434, n435, n436,
    n437, n438, n439, n440, n441, n442, n443,
    n444, n445, n446, n447, n448, n449, n450,
    n451, n452, n453, n454, n455, n456, n457,
    n458, n459, n460, n461, n462, n463, n464,
    n465, n466, n467, n468, n469, n470, n471,
    n472, n473, n474, n475, n476, n477, n478,
    n479, n480, n481, n482, n483, n484, n485,
    n486, n487, n488, n489, n490, n491, n492,
    n493, n494, n495, n496, n497, n498, n499,
    n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513,
    n514, n515, n516, n517, n518, n519, n520,
    n521, n522, n523, n524, n525, n526, n527,
    n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541,
    n542, n543, n544, n545, n546, n547, n548,
    n549, n550, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n561, n562,
    n563, n564, n565, n566, n567, n568, n569,
    n570, n571, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590,
    n591, n592, n593, n594, n595, n596, n597,
    n598, n599, n600, n601, n602, n603, n604,
    n605, n606, n607, n608, n609, n610, n611,
    n612, n613, n614, n615, n616, n617, n618,
    n619, n620, n621, n622, n623, n624, n625,
    n626, n627, n628, n629, n630, n631, n632,
    n633, n634, n635, n636, n637, n638, n639,
    n640, n641, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689,
    n690, n691, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731,
    n732, n733, n734, n735, n736, n737, n738,
    n739, n740, n741, n742, n743, n744, n745,
    n746, n747, n748, n749, n750, n751, n752,
    n753, n754, n755, n756, n757, n758, n759,
    n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n770, n771, n772, n773,
    n774, n775, n776, n777, n778, n779, n780,
    n781, n782, n783, n784, n785, n786, n787,
    n788, n789, n790, n791, n792, n793, n794,
    n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815,
    n816, n817, n818, n819, n820, n821, n822,
    n823, n824, n825, n826, n827, n828, n829,
    n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857,
    n858, n859, n860, n861, n862, n863, n864,
    n865, n866, n867, n868, n869, n870, n871,
    n872, n873, n874, n875, n876, n877, n878,
    n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n904, n905, n906,
    n907, n908, n909, n910, n911, n912, n913,
    n914, n915, n916, n917, n918, n919, n920,
    n921, n922, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n934,
    n935, n936, n937, n938, n939, n940, n941,
    n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955,
    n956, n957, n958, n959, n960, n961, n962,
    n963, n964, n965, n966, n967, n968, n969,
    n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990,
    n991, n992, n993, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330;
  assign n23 = pi00 & pi04;
  assign n24 = ~pi08 & pi09;
  assign n25 = pi13 & n24;
  assign n26 = ~pi10 & pi11;
  assign n27 = pi09 & pi11;
  assign n28 = ~pi08 & pi13;
  assign n29 = ~pi08 & pi11;
  assign n30 = pi09 & pi13;
  assign n31 = n29 & n30;
  assign n32 = n27 & n28;
  assign n33 = ~pi10 & n1181;
  assign n34 = n25 & n26;
  assign n35 = n23 & n1182;
  assign n36 = ~pi10 & ~pi13;
  assign n37 = ~pi10 & ~n27;
  assign n38 = ~pi13 & n37;
  assign n39 = ~n27 & n36;
  assign n40 = ~pi08 & ~pi10;
  assign n41 = ~pi13 & ~n27;
  assign n42 = n40 & n41;
  assign n43 = ~pi08 & n1183;
  assign n44 = ~pi00 & n1184;
  assign n45 = ~pi08 & ~pi09;
  assign n46 = pi08 & pi09;
  assign n47 = ~n45 & ~n46;
  assign n48 = pi11 & ~n47;
  assign n49 = ~pi10 & n48;
  assign n50 = n26 & ~n47;
  assign n51 = pi13 & n1185;
  assign n52 = ~pi09 & ~pi11;
  assign n53 = ~pi08 & pi10;
  assign n54 = pi10 & ~pi11;
  assign n55 = ~pi08 & n54;
  assign n56 = ~pi09 & n55;
  assign n57 = n52 & n53;
  assign n58 = ~n51 & ~n1186;
  assign n59 = n23 & ~n58;
  assign n60 = pi08 & pi10;
  assign n61 = ~pi09 & pi11;
  assign n62 = ~pi13 & n61;
  assign n63 = ~pi13 & n60;
  assign n64 = n61 & n63;
  assign n65 = n60 & n62;
  assign n66 = n24 & ~n54;
  assign n67 = pi13 & n66;
  assign n68 = n25 & ~n54;
  assign n69 = n46 & n54;
  assign n70 = ~n1188 & ~n69;
  assign n71 = ~n1187 & ~n1188;
  assign n72 = ~n69 & n71;
  assign n73 = ~n1187 & n70;
  assign n74 = ~pi04 & ~n1189;
  assign n75 = ~pi00 & ~pi04;
  assign n76 = ~pi10 & ~pi11;
  assign n77 = ~pi13 & ~n76;
  assign n78 = ~pi10 & pi13;
  assign n79 = pi08 & ~pi09;
  assign n80 = ~n78 & n79;
  assign n81 = pi10 & pi13;
  assign n82 = ~pi13 & n76;
  assign n83 = ~n81 & ~n82;
  assign n84 = n79 & ~n83;
  assign n85 = ~n77 & n80;
  assign n86 = ~n75 & n1190;
  assign n87 = ~pi00 & ~n54;
  assign n88 = ~pi00 & pi04;
  assign n89 = pi00 & ~pi04;
  assign n90 = ~n88 & ~n89;
  assign n91 = ~n23 & ~n75;
  assign n92 = n25 & ~n1191;
  assign n93 = n54 & n88;
  assign n94 = ~n89 & ~n93;
  assign n95 = pi13 & ~n94;
  assign n96 = n24 & n95;
  assign n97 = ~n87 & n92;
  assign n98 = ~n86 & ~n1192;
  assign n99 = ~n74 & n98;
  assign n100 = ~n59 & n99;
  assign n101 = ~n59 & ~n86;
  assign n102 = ~n44 & ~n74;
  assign n103 = n101 & n102;
  assign n104 = ~n1192 & n103;
  assign n105 = ~n44 & n100;
  assign n106 = ~pi00 & n1193;
  assign n107 = n1181 & ~n106;
  assign n108 = pi13 & n54;
  assign n109 = pi00 & ~n1193;
  assign n110 = pi00 & ~n100;
  assign n111 = n46 & n1194;
  assign n112 = n45 & n1193;
  assign n113 = n23 & n79;
  assign n114 = ~n112 & ~n113;
  assign n115 = ~n111 & ~n113;
  assign n116 = ~n112 & n115;
  assign n117 = ~n111 & n114;
  assign n118 = n108 & ~n1195;
  assign n119 = ~n107 & ~n118;
  assign n120 = pi08 & n54;
  assign n121 = ~pi09 & pi13;
  assign n122 = n120 & n121;
  assign n123 = n79 & n108;
  assign n124 = n119 & n1196;
  assign n125 = ~n35 & ~n124;
  assign n126 = n54 & n79;
  assign n127 = pi10 & n52;
  assign n128 = ~pi09 & n54;
  assign n129 = pi08 & n125;
  assign n130 = n1197 & n129;
  assign n131 = n125 & n126;
  assign n132 = ~pi10 & ~n45;
  assign n133 = ~pi00 & pi11;
  assign n134 = ~pi00 & ~n132;
  assign n135 = pi11 & n134;
  assign n136 = ~n132 & n133;
  assign n137 = ~n1193 & ~n1199;
  assign n138 = ~n1198 & n137;
  assign n139 = pi00 & pi11;
  assign n140 = ~n46 & n139;
  assign n141 = ~n124 & ~n140;
  assign n142 = pi10 & ~n141;
  assign n143 = ~pi10 & n46;
  assign n144 = pi11 & n143;
  assign n145 = n26 & n46;
  assign n146 = pi10 & n24;
  assign n147 = ~pi11 & n146;
  assign n148 = pi09 & n55;
  assign n149 = n24 & n54;
  assign n150 = ~n1200 & ~n1201;
  assign n151 = n1193 & n150;
  assign n152 = ~n142 & n151;
  assign n153 = ~n138 & ~n152;
  assign n154 = pi09 & ~pi10;
  assign n155 = n29 & n154;
  assign n156 = n24 & n26;
  assign n157 = pi09 & n40;
  assign n158 = n125 & n157;
  assign n159 = pi11 & n158;
  assign n160 = n125 & n1202;
  assign n161 = ~pi00 & ~pi08;
  assign n162 = n1197 & n161;
  assign n163 = ~pi00 & n1186;
  assign n164 = ~n119 & ~n1204;
  assign n165 = ~n1203 & n164;
  assign n166 = ~n69 & n119;
  assign n167 = ~n165 & ~n166;
  assign n168 = pi08 & ~pi10;
  assign n169 = pi04 & n168;
  assign n170 = pi00 & ~pi08;
  assign n171 = n119 & n170;
  assign n172 = ~n169 & ~n171;
  assign n173 = n52 & ~n172;
  assign n174 = ~pi09 & n1193;
  assign n175 = pi11 & ~n174;
  assign n176 = pi09 & ~n1193;
  assign n177 = ~pi00 & ~n176;
  assign n178 = n40 & ~n177;
  assign n179 = ~pi11 & ~n177;
  assign n180 = pi00 & ~pi09;
  assign n181 = n1193 & n180;
  assign n182 = ~n179 & ~n181;
  assign n183 = n40 & ~n182;
  assign n184 = n40 & ~n175;
  assign n185 = ~n177 & n184;
  assign n186 = ~n175 & n178;
  assign n187 = pi09 & n60;
  assign n188 = pi10 & n46;
  assign n189 = ~pi00 & n1206;
  assign n190 = pi11 & n189;
  assign n191 = n133 & n1206;
  assign n192 = ~pi09 & n168;
  assign n193 = ~pi10 & ~n1191;
  assign n194 = n79 & n193;
  assign n195 = ~n1191 & n192;
  assign n196 = ~n1207 & ~n1208;
  assign n197 = ~n1205 & n196;
  assign n198 = ~n173 & n197;
  assign n199 = ~n167 & n198;
  assign n200 = ~n1203 & ~n1204;
  assign n201 = ~n119 & ~n200;
  assign n202 = ~n1198 & ~n1199;
  assign n203 = ~n1193 & ~n202;
  assign n204 = ~n142 & n150;
  assign n205 = n1193 & ~n204;
  assign n206 = ~n35 & ~n69;
  assign n207 = n119 & ~n206;
  assign n208 = ~n1207 & ~n207;
  assign n209 = ~n173 & n208;
  assign n210 = ~n205 & n209;
  assign n211 = ~n203 & n210;
  assign n212 = ~n1205 & n211;
  assign n213 = ~n201 & n212;
  assign n214 = ~n1208 & n213;
  assign n215 = n198 & ~n207;
  assign n216 = ~n201 & ~n203;
  assign n217 = n215 & n216;
  assign n218 = ~n205 & n217;
  assign n219 = ~n153 & n199;
  assign n220 = ~pi12 & pi13;
  assign n221 = pi13 & ~n1209;
  assign n222 = ~pi12 & n221;
  assign n223 = ~n1209 & n220;
  assign n224 = pi01 & pi05;
  assign n225 = pi13 & n1197;
  assign n226 = n58 & ~n225;
  assign n227 = ~pi08 & n88;
  assign n228 = n28 & n93;
  assign n229 = n108 & n227;
  assign n230 = n226 & ~n1211;
  assign n231 = n224 & ~n230;
  assign n232 = ~pi05 & ~n1189;
  assign n233 = ~pi09 & pi10;
  assign n234 = n139 & n233;
  assign n235 = ~pi01 & pi05;
  assign n236 = n54 & n235;
  assign n237 = pi01 & ~pi05;
  assign n238 = ~n88 & ~n237;
  assign n239 = ~n236 & n238;
  assign n240 = ~pi01 & ~pi05;
  assign n241 = n88 & ~n240;
  assign n242 = pi09 & ~n241;
  assign n243 = ~n236 & ~n237;
  assign n244 = ~n88 & ~n243;
  assign n245 = n88 & n240;
  assign n246 = ~n244 & ~n245;
  assign n247 = pi09 & ~n246;
  assign n248 = ~n239 & n242;
  assign n249 = ~n234 & ~n1212;
  assign n250 = ~pi08 & ~n249;
  assign n251 = pi13 & n250;
  assign n252 = n28 & ~n249;
  assign n253 = ~pi01 & n1184;
  assign n254 = n1190 & ~n240;
  assign n255 = ~n253 & ~n254;
  assign n256 = ~n1213 & n255;
  assign n257 = ~n232 & ~n253;
  assign n258 = ~n254 & n257;
  assign n259 = ~n1213 & n258;
  assign n260 = ~n232 & n256;
  assign n261 = ~n231 & n1214;
  assign n262 = n1182 & n224;
  assign n263 = ~pi01 & n261;
  assign n264 = ~pi01 & n1214;
  assign n265 = n1181 & ~n1215;
  assign n266 = ~pi05 & ~pi09;
  assign n267 = pi01 & pi08;
  assign n268 = ~n266 & n267;
  assign n269 = ~pi08 & n261;
  assign n270 = ~n268 & ~n269;
  assign n271 = pi09 & n261;
  assign n272 = n108 & ~n271;
  assign n273 = n45 & n261;
  assign n274 = pi09 & ~n261;
  assign n275 = pi05 & ~pi09;
  assign n276 = ~n274 & ~n275;
  assign n277 = pi08 & ~n276;
  assign n278 = pi01 & n277;
  assign n279 = ~n273 & ~n278;
  assign n280 = n108 & ~n279;
  assign n281 = ~n270 & n272;
  assign n282 = ~n265 & ~n1216;
  assign n283 = n1196 & n282;
  assign n284 = ~n262 & ~n283;
  assign n285 = ~n1193 & ~n125;
  assign n286 = ~n284 & n285;
  assign n287 = n284 & ~n285;
  assign n288 = ~n284 & ~n285;
  assign n289 = n284 & n285;
  assign n290 = ~n288 & ~n289;
  assign n291 = ~n286 & ~n287;
  assign n292 = ~n261 & ~n1217;
  assign n293 = n261 & n1217;
  assign n294 = n60 & ~n293;
  assign n295 = ~n261 & n1217;
  assign n296 = n261 & ~n1217;
  assign n297 = ~n295 & ~n296;
  assign n298 = n60 & ~n297;
  assign n299 = ~n292 & n294;
  assign n300 = pi00 & ~n119;
  assign n301 = n282 & ~n300;
  assign n302 = ~n119 & ~n282;
  assign n303 = pi00 & n302;
  assign n304 = n282 & n300;
  assign n305 = ~n282 & ~n300;
  assign n306 = ~n304 & ~n305;
  assign n307 = ~n301 & ~n303;
  assign n308 = pi01 & ~pi08;
  assign n309 = ~pi08 & n1219;
  assign n310 = pi01 & n309;
  assign n311 = n1219 & n308;
  assign n312 = pi05 & n168;
  assign n313 = ~n1220 & ~n312;
  assign n314 = ~n1218 & n313;
  assign n315 = n52 & ~n314;
  assign n316 = n35 & ~n284;
  assign n317 = ~n35 & n284;
  assign n318 = n35 & n284;
  assign n319 = ~n35 & ~n284;
  assign n320 = ~n318 & ~n319;
  assign n321 = ~n316 & ~n317;
  assign n322 = ~n282 & ~n1221;
  assign n323 = n282 & n1221;
  assign n324 = n1202 & ~n323;
  assign n325 = ~n282 & n1221;
  assign n326 = n282 & ~n1221;
  assign n327 = ~n325 & ~n326;
  assign n328 = n1202 & ~n327;
  assign n329 = n1202 & ~n322;
  assign n330 = ~n323 & n329;
  assign n331 = ~n322 & n324;
  assign n332 = pi10 & ~n46;
  assign n333 = ~n45 & ~n332;
  assign n334 = pi11 & ~n333;
  assign n335 = n1194 & ~n261;
  assign n336 = ~n1194 & n261;
  assign n337 = n1194 & n261;
  assign n338 = ~n1194 & ~n261;
  assign n339 = ~n337 & ~n338;
  assign n340 = ~n335 & ~n336;
  assign n341 = n334 & ~n1223;
  assign n342 = n53 & ~n1219;
  assign n343 = n52 & n342;
  assign n344 = n1186 & ~n1219;
  assign n345 = ~n341 & ~n1224;
  assign n346 = ~pi01 & ~n345;
  assign n347 = n119 & n282;
  assign n348 = ~n302 & ~n347;
  assign n349 = n1206 & ~n348;
  assign n350 = n157 & ~n261;
  assign n351 = ~n349 & ~n350;
  assign n352 = ~pi11 & ~n351;
  assign n353 = ~pi10 & n45;
  assign n354 = ~n334 & ~n353;
  assign n355 = ~n54 & ~n333;
  assign n356 = n1223 & ~n1225;
  assign n357 = n139 & n1206;
  assign n358 = ~pi05 & ~n23;
  assign n359 = n192 & n358;
  assign n360 = ~n46 & n76;
  assign n361 = ~n359 & ~n360;
  assign n362 = ~n357 & ~n359;
  assign n363 = ~n360 & n362;
  assign n364 = ~n357 & n361;
  assign n365 = ~n356 & n1226;
  assign n366 = pi01 & ~n365;
  assign n367 = n1193 & n261;
  assign n368 = ~n150 & n367;
  assign n369 = ~pi11 & n24;
  assign n370 = ~n1200 & ~n369;
  assign n371 = ~n1193 & ~n370;
  assign n372 = ~n261 & n371;
  assign n373 = ~pi00 & ~pi01;
  assign n374 = n1206 & n373;
  assign n375 = n23 & n240;
  assign n376 = n192 & n375;
  assign n377 = ~n374 & ~n376;
  assign n378 = pi11 & ~n377;
  assign n379 = n23 & ~n224;
  assign n380 = ~n23 & ~n235;
  assign n381 = n192 & ~n380;
  assign n382 = ~n23 & n235;
  assign n383 = n23 & n224;
  assign n384 = ~n382 & ~n383;
  assign n385 = n192 & ~n384;
  assign n386 = ~n379 & n381;
  assign n387 = ~n378 & ~n1227;
  assign n388 = ~n372 & n387;
  assign n389 = ~n368 & n388;
  assign n390 = ~n366 & n389;
  assign n391 = ~n352 & n390;
  assign n392 = ~n346 & n391;
  assign n393 = ~n1222 & n392;
  assign n394 = ~n368 & ~n372;
  assign n395 = ~n1227 & n394;
  assign n396 = ~n352 & n395;
  assign n397 = ~n366 & n396;
  assign n398 = ~n1222 & n397;
  assign n399 = ~n378 & n398;
  assign n400 = ~n315 & n399;
  assign n401 = ~n346 & n400;
  assign n402 = ~n315 & n393;
  assign n403 = pi13 & ~n1228;
  assign n404 = n1210 & n403;
  assign n405 = n1210 & ~n1228;
  assign n406 = ~n88 & ~n235;
  assign n407 = n88 & ~n237;
  assign n408 = ~n235 & ~n407;
  assign n409 = ~n237 & ~n406;
  assign n410 = ~pi06 & n1230;
  assign n411 = pi09 & n1230;
  assign n412 = ~pi06 & n411;
  assign n413 = pi09 & n410;
  assign n414 = pi06 & ~n1230;
  assign n415 = n54 & ~n1230;
  assign n416 = pi06 & n415;
  assign n417 = n54 & n414;
  assign n418 = ~n1231 & ~n1232;
  assign n419 = pi02 & ~n418;
  assign n420 = ~pi02 & pi09;
  assign n421 = ~n414 & n420;
  assign n422 = ~n54 & n1230;
  assign n423 = ~n410 & ~n422;
  assign n424 = ~pi02 & ~n410;
  assign n425 = pi09 & ~n414;
  assign n426 = ~n422 & n425;
  assign n427 = n424 & n426;
  assign n428 = ~pi06 & ~n1230;
  assign n429 = n54 & n1230;
  assign n430 = pi06 & n429;
  assign n431 = ~n428 & ~n430;
  assign n432 = pi09 & ~n431;
  assign n433 = ~pi02 & n432;
  assign n434 = n421 & n423;
  assign n435 = pi01 & pi11;
  assign n436 = n233 & n435;
  assign n437 = ~n1233 & ~n436;
  assign n438 = ~n419 & ~n436;
  assign n439 = ~n1233 & n438;
  assign n440 = ~n419 & n437;
  assign n441 = ~pi08 & ~n1234;
  assign n442 = pi13 & n441;
  assign n443 = n28 & ~n1234;
  assign n444 = pi02 & pi06;
  assign n445 = ~n226 & n444;
  assign n446 = ~pi06 & ~n1189;
  assign n447 = ~pi02 & n1184;
  assign n448 = ~pi02 & ~pi06;
  assign n449 = n1190 & ~n448;
  assign n450 = ~n447 & ~n449;
  assign n451 = ~n446 & n450;
  assign n452 = ~n445 & ~n446;
  assign n453 = n450 & n452;
  assign n454 = ~n445 & n451;
  assign n455 = ~n1235 & n1236;
  assign n456 = n1182 & n444;
  assign n457 = ~pi02 & n455;
  assign n458 = n1181 & ~n457;
  assign n459 = ~pi06 & ~pi09;
  assign n460 = pi02 & pi08;
  assign n461 = ~n459 & n460;
  assign n462 = ~pi08 & n455;
  assign n463 = ~n461 & ~n462;
  assign n464 = pi09 & n455;
  assign n465 = n108 & ~n464;
  assign n466 = n45 & n455;
  assign n467 = pi09 & ~n455;
  assign n468 = pi06 & ~pi09;
  assign n469 = ~n467 & ~n468;
  assign n470 = pi08 & ~n469;
  assign n471 = pi02 & n470;
  assign n472 = ~n466 & ~n471;
  assign n473 = n108 & ~n472;
  assign n474 = ~n463 & n465;
  assign n475 = ~n458 & ~n1237;
  assign n476 = n1196 & n475;
  assign n477 = ~n456 & ~n476;
  assign n478 = n455 & n477;
  assign n479 = ~n455 & ~n477;
  assign n480 = ~n478 & ~n479;
  assign n481 = ~n261 & ~n287;
  assign n482 = ~n286 & ~n481;
  assign n483 = ~n480 & n482;
  assign n484 = n480 & ~n482;
  assign n485 = n60 & ~n484;
  assign n486 = ~n480 & ~n482;
  assign n487 = n480 & n482;
  assign n488 = ~n486 & ~n487;
  assign n489 = n60 & ~n488;
  assign n490 = n60 & ~n483;
  assign n491 = ~n484 & n490;
  assign n492 = ~n483 & n485;
  assign n493 = pi06 & n168;
  assign n494 = pi01 & ~n301;
  assign n495 = ~pi01 & ~n300;
  assign n496 = ~n282 & ~n495;
  assign n497 = pi01 & n300;
  assign n498 = ~n496 & ~n497;
  assign n499 = ~n303 & ~n494;
  assign n500 = ~n475 & ~n1239;
  assign n501 = n475 & n1239;
  assign n502 = ~n475 & n1239;
  assign n503 = n475 & ~n1239;
  assign n504 = ~n502 & ~n503;
  assign n505 = ~n500 & ~n501;
  assign n506 = pi02 & ~pi08;
  assign n507 = ~pi08 & n1240;
  assign n508 = pi02 & n507;
  assign n509 = n1240 & n506;
  assign n510 = ~n493 & ~n1241;
  assign n511 = ~n1238 & n510;
  assign n512 = n52 & ~n511;
  assign n513 = ~n282 & ~n317;
  assign n514 = n477 & ~n513;
  assign n515 = ~n477 & n513;
  assign n516 = ~n514 & ~n515;
  assign n517 = n475 & ~n516;
  assign n518 = ~n475 & n516;
  assign n519 = n1202 & ~n518;
  assign n520 = ~n475 & n513;
  assign n521 = n475 & ~n513;
  assign n522 = ~n475 & ~n513;
  assign n523 = n475 & n513;
  assign n524 = ~n522 & ~n523;
  assign n525 = ~n520 & ~n521;
  assign n526 = ~n477 & n1242;
  assign n527 = n477 & ~n1242;
  assign n528 = ~n526 & ~n527;
  assign n529 = n1202 & ~n528;
  assign n530 = n1202 & ~n517;
  assign n531 = ~n518 & n530;
  assign n532 = ~n517 & n519;
  assign n533 = n53 & ~n1240;
  assign n534 = n52 & n533;
  assign n535 = n1186 & ~n1240;
  assign n536 = ~pi01 & ~n335;
  assign n537 = ~pi01 & ~n1194;
  assign n538 = ~n261 & ~n537;
  assign n539 = pi01 & n1194;
  assign n540 = ~n538 & ~n539;
  assign n541 = pi01 & ~n336;
  assign n542 = ~n335 & ~n541;
  assign n543 = ~n336 & ~n536;
  assign n544 = n334 & ~n455;
  assign n545 = n334 & n1245;
  assign n546 = ~n455 & n545;
  assign n547 = n1245 & n544;
  assign n548 = ~n1244 & ~n1246;
  assign n549 = ~pi02 & ~n548;
  assign n550 = ~n347 & ~n475;
  assign n551 = n347 & n475;
  assign n552 = ~pi11 & ~n551;
  assign n553 = ~n550 & n552;
  assign n554 = ~pi02 & n373;
  assign n555 = pi02 & ~n373;
  assign n556 = pi11 & ~n555;
  assign n557 = ~n554 & n556;
  assign n558 = n1206 & ~n557;
  assign n559 = ~n550 & ~n551;
  assign n560 = ~pi11 & ~n559;
  assign n561 = pi11 & n554;
  assign n562 = pi02 & pi11;
  assign n563 = ~n373 & n562;
  assign n564 = ~n561 & ~n563;
  assign n565 = ~n560 & n564;
  assign n566 = n1206 & ~n565;
  assign n567 = ~n553 & n558;
  assign n568 = ~n455 & ~n1245;
  assign n569 = ~n1225 & ~n1245;
  assign n570 = n334 & ~n1245;
  assign n571 = ~n455 & n1248;
  assign n572 = ~n1225 & n568;
  assign n573 = ~n360 & ~n1249;
  assign n574 = pi02 & ~n573;
  assign n575 = ~pi02 & n334;
  assign n576 = ~n1225 & n1245;
  assign n577 = ~n575 & ~n576;
  assign n578 = ~pi02 & n1245;
  assign n579 = n455 & ~n578;
  assign n580 = ~pi02 & n1248;
  assign n581 = ~n1245 & n575;
  assign n582 = pi02 & n576;
  assign n583 = ~n1250 & ~n582;
  assign n584 = n455 & ~n583;
  assign n585 = ~n577 & n579;
  assign n586 = ~pi11 & n157;
  assign n587 = ~pi10 & n369;
  assign n588 = n367 & ~n1252;
  assign n589 = ~n370 & ~n455;
  assign n590 = ~n367 & ~n370;
  assign n591 = ~n1252 & ~n590;
  assign n592 = ~n455 & ~n591;
  assign n593 = ~n588 & n589;
  assign n594 = ~n23 & ~n224;
  assign n595 = n23 & ~n240;
  assign n596 = ~n224 & ~n595;
  assign n597 = ~n240 & ~n594;
  assign n598 = pi11 & n448;
  assign n599 = ~n444 & ~n598;
  assign n600 = ~n1254 & n599;
  assign n601 = ~pi02 & pi06;
  assign n602 = pi02 & ~pi06;
  assign n603 = ~n601 & ~n602;
  assign n604 = ~n444 & ~n448;
  assign n605 = n1254 & n1255;
  assign n606 = n192 & ~n605;
  assign n607 = ~n1254 & ~n599;
  assign n608 = n1254 & ~n1255;
  assign n609 = ~n607 & ~n608;
  assign n610 = n192 & ~n609;
  assign n611 = ~n600 & n606;
  assign n612 = n367 & n455;
  assign n613 = ~n150 & n612;
  assign n614 = n368 & n455;
  assign n615 = ~n1256 & ~n1257;
  assign n616 = ~n1253 & n615;
  assign n617 = ~n1251 & n616;
  assign n618 = n455 & n1245;
  assign n619 = ~n568 & ~n618;
  assign n620 = ~n1225 & ~n619;
  assign n621 = ~n360 & ~n620;
  assign n622 = pi02 & ~n621;
  assign n623 = ~n368 & ~n1250;
  assign n624 = n455 & ~n623;
  assign n625 = ~n1253 & ~n1256;
  assign n626 = ~n624 & n625;
  assign n627 = ~n622 & n626;
  assign n628 = ~n574 & n617;
  assign n629 = ~n1247 & n1258;
  assign n630 = ~n549 & n629;
  assign n631 = ~n1243 & n630;
  assign n632 = ~n1247 & ~n1257;
  assign n633 = ~n1253 & n632;
  assign n634 = ~n574 & n633;
  assign n635 = ~n512 & n634;
  assign n636 = ~n1243 & n635;
  assign n637 = ~n549 & n636;
  assign n638 = ~n1256 & n637;
  assign n639 = ~n1251 & n638;
  assign n640 = ~n512 & n631;
  assign n641 = pi13 & ~n1259;
  assign n642 = n1229 & n641;
  assign n643 = n1229 & ~n1259;
  assign n644 = n233 & n562;
  assign n645 = n1230 & ~n601;
  assign n646 = ~n414 & ~n424;
  assign n647 = pi02 & ~n414;
  assign n648 = ~n410 & ~n647;
  assign n649 = ~n602 & ~n645;
  assign n650 = ~pi03 & ~pi07;
  assign n651 = pi09 & n650;
  assign n652 = pi09 & ~n1261;
  assign n653 = n650 & n652;
  assign n654 = ~n1261 & n651;
  assign n655 = ~n644 & ~n1262;
  assign n656 = pi13 & ~n655;
  assign po5 = pi03 & pi07;
  assign n658 = n54 & ~n1261;
  assign n659 = pi13 & n658;
  assign n660 = n108 & ~n1261;
  assign n661 = ~n1197 & ~n1263;
  assign n662 = po5 & ~n661;
  assign n663 = pi07 & pi09;
  assign n664 = n108 & n663;
  assign n665 = pi07 & pi13;
  assign n666 = pi09 & n54;
  assign n667 = n1261 & n666;
  assign n668 = n665 & n667;
  assign n669 = n1261 & n664;
  assign n670 = ~n1183 & ~n1264;
  assign n671 = ~pi03 & ~n670;
  assign n672 = ~n662 & ~n671;
  assign n673 = ~n656 & ~n671;
  assign n674 = ~n662 & n673;
  assign n675 = ~n656 & n672;
  assign n676 = ~pi08 & ~n1265;
  assign n677 = pi03 & n25;
  assign n678 = pi09 & n1261;
  assign n679 = pi03 & n678;
  assign n680 = n28 & n679;
  assign n681 = n1261 & n677;
  assign n682 = n1189 & ~n1266;
  assign n683 = ~pi07 & ~n682;
  assign n684 = n1190 & ~n650;
  assign n685 = ~n1185 & ~n1197;
  assign n686 = pi13 & po5;
  assign n687 = pi13 & ~n685;
  assign n688 = po5 & n687;
  assign n689 = ~n685 & n686;
  assign n690 = ~n684 & ~n1267;
  assign n691 = ~n683 & n690;
  assign n692 = ~n676 & n690;
  assign n693 = ~n683 & n692;
  assign n694 = ~n676 & n691;
  assign n695 = ~pi03 & n1268;
  assign n696 = n1181 & ~n695;
  assign n697 = pi03 & ~n1268;
  assign n698 = n46 & n697;
  assign n699 = n45 & n1268;
  assign n700 = n79 & po5;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n698 & ~n700;
  assign n703 = ~n699 & n702;
  assign n704 = ~n698 & n701;
  assign n705 = n108 & ~n1269;
  assign n706 = ~n696 & ~n705;
  assign n707 = n1182 & po5;
  assign n708 = n1196 & n706;
  assign n709 = ~n707 & ~n708;
  assign n710 = ~n475 & ~n514;
  assign n711 = n709 & ~n710;
  assign n712 = ~n709 & n710;
  assign n713 = ~n711 & ~n712;
  assign n714 = ~n706 & n713;
  assign n715 = n706 & ~n713;
  assign n716 = n157 & ~n715;
  assign n717 = ~n706 & n710;
  assign n718 = n706 & ~n710;
  assign n719 = ~n706 & ~n710;
  assign n720 = n706 & n710;
  assign n721 = ~n719 & ~n720;
  assign n722 = ~n717 & ~n718;
  assign n723 = ~n709 & n1270;
  assign n724 = n709 & ~n1270;
  assign n725 = ~n723 & ~n724;
  assign n726 = n157 & ~n725;
  assign n727 = ~n714 & n716;
  assign n728 = ~pi03 & n192;
  assign n729 = ~n444 & n1254;
  assign n730 = ~n448 & ~n1254;
  assign n731 = ~n444 & ~n730;
  assign n732 = ~n448 & ~n729;
  assign n733 = ~pi07 & ~n1272;
  assign n734 = n650 & ~n1272;
  assign n735 = n192 & n734;
  assign n736 = n728 & n733;
  assign n737 = ~pi03 & n1206;
  assign n738 = ~pi03 & n554;
  assign n739 = n1206 & n738;
  assign n740 = n554 & n737;
  assign n741 = ~n1273 & ~n1274;
  assign n742 = ~n1271 & n741;
  assign n743 = pi11 & ~n742;
  assign n744 = ~pi02 & n475;
  assign n745 = ~n1239 & ~n744;
  assign n746 = pi02 & ~n475;
  assign n747 = pi02 & ~n501;
  assign n748 = ~n500 & ~n747;
  assign n749 = ~pi02 & n1239;
  assign n750 = ~n475 & ~n749;
  assign n751 = pi02 & ~n1239;
  assign n752 = ~n750 & ~n751;
  assign n753 = ~n745 & ~n746;
  assign n754 = ~n706 & ~n1275;
  assign n755 = ~pi03 & ~n754;
  assign n756 = n706 & n1275;
  assign n757 = ~pi08 & ~n756;
  assign n758 = n706 & ~n1275;
  assign n759 = ~n706 & n1275;
  assign n760 = ~n758 & ~n759;
  assign n761 = ~n754 & ~n756;
  assign n762 = ~pi08 & ~n1276;
  assign n763 = ~pi03 & n762;
  assign n764 = n755 & n757;
  assign n765 = ~n1268 & ~n709;
  assign n766 = n1268 & n709;
  assign n767 = ~n1268 & n709;
  assign n768 = n1268 & ~n709;
  assign n769 = ~n767 & ~n768;
  assign n770 = ~n765 & ~n766;
  assign n771 = n477 & n482;
  assign n772 = ~n455 & ~n771;
  assign n773 = ~n477 & ~n482;
  assign n774 = ~n772 & ~n773;
  assign n775 = ~n479 & n482;
  assign n776 = ~n1278 & ~n1279;
  assign n777 = n1278 & n1279;
  assign n778 = pi08 & ~n777;
  assign n779 = n1278 & ~n1279;
  assign n780 = ~n1278 & n1279;
  assign n781 = ~n779 & ~n780;
  assign n782 = pi08 & ~n781;
  assign n783 = ~n776 & n778;
  assign n784 = ~n1277 & ~n1280;
  assign n785 = n1197 & ~n784;
  assign n786 = pi03 & n45;
  assign n787 = n45 & n1276;
  assign n788 = pi03 & n787;
  assign n789 = n1276 & n786;
  assign n790 = pi07 & n192;
  assign n791 = n551 & n706;
  assign n792 = ~n551 & ~n706;
  assign n793 = ~n791 & ~n792;
  assign n794 = n1206 & ~n793;
  assign n795 = ~n790 & ~n794;
  assign n796 = ~n1281 & ~n790;
  assign n797 = ~n794 & n796;
  assign n798 = ~n1281 & n795;
  assign n799 = ~pi11 & ~n1282;
  assign n800 = ~pi02 & ~n568;
  assign n801 = ~n455 & ~n578;
  assign n802 = pi02 & ~n1245;
  assign n803 = ~n801 & ~n802;
  assign n804 = pi02 & ~n618;
  assign n805 = ~n568 & ~n804;
  assign n806 = ~n618 & ~n800;
  assign n807 = ~n1268 & ~n1283;
  assign n808 = n1268 & n1283;
  assign n809 = ~n1268 & n1283;
  assign n810 = n1268 & ~n1283;
  assign n811 = ~n809 & ~n810;
  assign n812 = ~n807 & ~n808;
  assign n813 = ~n1225 & n1284;
  assign n814 = ~n360 & ~n813;
  assign n815 = pi03 & ~n814;
  assign n816 = n334 & ~n1284;
  assign n817 = pi07 & n1272;
  assign n818 = n192 & n817;
  assign n819 = n1272 & n790;
  assign n820 = ~n816 & ~n1285;
  assign n821 = ~pi03 & ~n820;
  assign n822 = ~n1252 & n612;
  assign n823 = ~n370 & ~n1268;
  assign n824 = ~n370 & ~n612;
  assign n825 = ~n1252 & ~n824;
  assign n826 = ~n370 & ~n822;
  assign n827 = ~n1268 & ~n1286;
  assign n828 = ~n822 & n823;
  assign n829 = n612 & n1268;
  assign n830 = ~n150 & n829;
  assign n831 = n1257 & n1268;
  assign n832 = pi03 & n192;
  assign n833 = ~n733 & n832;
  assign n834 = ~pi07 & n1272;
  assign n835 = pi03 & n834;
  assign n836 = po5 & ~n1272;
  assign n837 = ~n835 & ~n836;
  assign n838 = n192 & ~n837;
  assign n839 = ~n817 & n833;
  assign n840 = pi03 & pi11;
  assign n841 = n1206 & n840;
  assign n842 = ~n554 & n840;
  assign n843 = n1206 & n842;
  assign n844 = ~n554 & n841;
  assign n845 = ~n1289 & ~n1290;
  assign n846 = ~n1288 & n845;
  assign n847 = ~n1287 & n845;
  assign n848 = ~n1288 & n847;
  assign n849 = ~n1287 & n846;
  assign n850 = ~n821 & n1291;
  assign n851 = ~n815 & n850;
  assign n852 = ~n799 & n851;
  assign n853 = ~n785 & n852;
  assign n854 = ~n1288 & ~n1290;
  assign n855 = ~n815 & n854;
  assign n856 = ~n1289 & n855;
  assign n857 = ~n799 & n856;
  assign n858 = ~n821 & n857;
  assign n859 = ~n743 & n858;
  assign n860 = ~n785 & n859;
  assign n861 = ~n1287 & n860;
  assign n862 = ~n743 & n853;
  assign n863 = pi13 & ~n1292;
  assign n864 = n1260 & n863;
  assign n865 = n1260 & ~n1292;
  assign n866 = ~n1260 & n1292;
  assign n867 = pi13 & ~n866;
  assign n868 = ~n1260 & n863;
  assign n869 = n1260 & ~n863;
  assign n870 = ~n868 & ~n869;
  assign n871 = ~n1293 & n867;
  assign n872 = ~pi11 & n46;
  assign n873 = n46 & n76;
  assign n874 = pi13 & n873;
  assign n875 = ~pi11 & pi13;
  assign n876 = n143 & n875;
  assign n877 = n78 & n872;
  assign n878 = ~pi13 & n29;
  assign n879 = n29 & n233;
  assign n880 = ~pi13 & n879;
  assign n881 = n233 & n878;
  assign n882 = ~n1295 & ~n1296;
  assign n883 = pi08 & n76;
  assign n884 = ~n53 & ~n883;
  assign n885 = n1268 & ~n884;
  assign n886 = ~pi07 & n120;
  assign n887 = ~pi09 & ~n886;
  assign n888 = ~n885 & n887;
  assign n889 = n60 & n697;
  assign n890 = n55 & n650;
  assign n891 = ~pi11 & ~n53;
  assign n892 = po5 & ~n891;
  assign n893 = pi09 & ~n892;
  assign n894 = ~n890 & n893;
  assign n895 = ~n889 & n894;
  assign n896 = ~n890 & ~n892;
  assign n897 = ~n889 & n896;
  assign n898 = pi09 & ~n897;
  assign n899 = ~n885 & ~n886;
  assign n900 = ~pi09 & ~n899;
  assign n901 = ~n898 & ~n900;
  assign n902 = ~n888 & ~n895;
  assign n903 = ~pi09 & ~n54;
  assign n904 = pi10 & pi11;
  assign n905 = ~n40 & ~n904;
  assign n906 = ~pi09 & ~n905;
  assign n907 = ~pi09 & ~n168;
  assign n908 = ~n54 & n907;
  assign n909 = ~n168 & n903;
  assign n910 = pi07 & n40;
  assign n911 = ~n1298 & ~n910;
  assign n912 = ~n1268 & ~n911;
  assign n913 = ~pi07 & ~pi09;
  assign n914 = n132 & ~n913;
  assign n915 = n840 & ~n914;
  assign n916 = ~n24 & ~n728;
  assign n917 = pi07 & pi11;
  assign n918 = pi09 & n29;
  assign n919 = ~pi03 & n168;
  assign n920 = pi11 & n168;
  assign n921 = ~pi03 & n920;
  assign n922 = ~pi09 & n921;
  assign n923 = n61 & n919;
  assign n924 = ~n918 & ~n1299;
  assign n925 = pi07 & ~n924;
  assign n926 = ~n916 & n917;
  assign n927 = ~n915 & ~n1300;
  assign n928 = ~n912 & n927;
  assign n929 = n1297 & ~n1300;
  assign n930 = ~n912 & n929;
  assign n931 = ~n915 & n930;
  assign n932 = ~n900 & n928;
  assign n933 = ~n898 & n932;
  assign n934 = n1297 & n928;
  assign n935 = ~pi13 & ~n1301;
  assign n936 = n882 & ~n935;
  assign n937 = n1294 & n936;
  assign n938 = ~pi03 & n1275;
  assign n939 = ~n706 & ~n938;
  assign n940 = pi03 & ~n1275;
  assign n941 = ~n939 & ~n940;
  assign n942 = ~pi08 & ~n941;
  assign n943 = ~n755 & n757;
  assign n944 = ~n709 & ~n1279;
  assign n945 = n1268 & ~n944;
  assign n946 = n1268 & n1279;
  assign n947 = ~n709 & ~n1303;
  assign n948 = ~n1268 & ~n1279;
  assign n949 = ~n947 & ~n948;
  assign n950 = n709 & n1279;
  assign n951 = pi08 & ~n950;
  assign n952 = ~n1303 & n951;
  assign n953 = ~n765 & n1279;
  assign n954 = ~n1302 & n1304;
  assign n955 = n233 & ~n954;
  assign n956 = pi10 & ~n791;
  assign n957 = n46 & ~n956;
  assign n958 = n46 & n791;
  assign n959 = ~n955 & ~n1305;
  assign n960 = ~pi11 & ~n959;
  assign n961 = n157 & ~n711;
  assign n962 = ~n706 & n961;
  assign n963 = ~n706 & ~n711;
  assign n964 = ~n697 & n1283;
  assign n965 = ~n333 & ~n695;
  assign n966 = ~n695 & ~n1283;
  assign n967 = ~n697 & ~n966;
  assign n968 = ~n333 & ~n967;
  assign n969 = ~n964 & n965;
  assign n970 = ~po5 & n1272;
  assign n971 = n192 & ~n650;
  assign n972 = ~n650 & ~n1272;
  assign n973 = ~po5 & ~n972;
  assign n974 = n192 & ~n973;
  assign n975 = ~n970 & n971;
  assign n976 = ~n1274 & ~n1308;
  assign n977 = ~n1274 & ~n1307;
  assign n978 = ~n1308 & n977;
  assign n979 = ~n1307 & n976;
  assign n980 = ~n1306 & n1309;
  assign n981 = pi11 & ~n980;
  assign n982 = ~n55 & ~n168;
  assign n983 = pi09 & ~n982;
  assign n984 = ~n143 & ~n1201;
  assign n985 = n612 & n1310;
  assign n986 = n829 & n1310;
  assign n987 = n1268 & n985;
  assign n988 = ~n981 & ~n1311;
  assign n989 = ~n960 & n988;
  assign n990 = ~n1293 & ~n960;
  assign n991 = ~n981 & n990;
  assign n992 = ~n1311 & n991;
  assign n993 = ~n1293 & n989;
  assign po6 = pi13 & ~n1312;
  assign n995 = ~n1229 & n1259;
  assign n996 = pi13 & ~n1260;
  assign n997 = ~n1229 & n641;
  assign n998 = n1229 & ~n641;
  assign n999 = ~n997 & ~n998;
  assign n1000 = pi13 & ~n995;
  assign n1001 = ~n1260 & n1000;
  assign n1002 = ~n995 & n996;
  assign n1003 = n455 & ~n884;
  assign n1004 = ~pi06 & n120;
  assign n1005 = ~n1003 & ~n1004;
  assign n1006 = ~pi09 & ~n1005;
  assign n1007 = pi02 & n60;
  assign n1008 = pi09 & n1007;
  assign n1009 = pi02 & n1206;
  assign n1010 = pi06 & n40;
  assign n1011 = ~n1298 & ~n1010;
  assign n1012 = ~n1298 & ~n1314;
  assign n1013 = ~n1010 & n1012;
  assign n1014 = ~n1314 & n1011;
  assign n1015 = ~n455 & ~n1315;
  assign n1016 = n444 & ~n891;
  assign n1017 = n55 & n448;
  assign n1018 = ~n1016 & ~n1017;
  assign n1019 = pi09 & ~n1018;
  assign n1020 = n132 & ~n459;
  assign n1021 = n562 & ~n1020;
  assign n1022 = ~pi02 & n168;
  assign n1023 = ~pi02 & n920;
  assign n1024 = ~pi09 & n1023;
  assign n1025 = n61 & n1022;
  assign n1026 = ~pi02 & n192;
  assign n1027 = ~n24 & ~n1026;
  assign n1028 = pi11 & ~n1027;
  assign n1029 = ~n918 & ~n1316;
  assign n1030 = pi06 & n1317;
  assign n1031 = ~n1021 & ~n1030;
  assign n1032 = ~n1019 & n1031;
  assign n1033 = ~n1015 & n1032;
  assign n1034 = n40 & ~n455;
  assign n1035 = ~n1317 & ~n1034;
  assign n1036 = pi06 & ~n1035;
  assign n1037 = ~n455 & ~n1012;
  assign n1038 = ~n1019 & ~n1021;
  assign n1039 = ~n1037 & n1038;
  assign n1040 = ~n1006 & n1039;
  assign n1041 = ~n1036 & n1040;
  assign n1042 = ~n1006 & ~n1019;
  assign n1043 = ~n1030 & n1042;
  assign n1044 = ~n1015 & n1043;
  assign n1045 = ~n1021 & n1044;
  assign n1046 = ~n1006 & n1033;
  assign n1047 = ~pi13 & ~n1318;
  assign n1048 = n882 & ~n1047;
  assign n1049 = n1313 & n1048;
  assign n1050 = ~n1210 & n1228;
  assign n1051 = pi13 & ~n1050;
  assign n1052 = ~n1210 & n403;
  assign n1053 = n1210 & ~n403;
  assign n1054 = ~n1052 & ~n1053;
  assign n1055 = ~n1229 & n1051;
  assign n1056 = n261 & ~n884;
  assign n1057 = ~pi01 & ~n168;
  assign n1058 = ~n224 & ~n240;
  assign n1059 = pi11 & n1058;
  assign n1060 = pi11 & n237;
  assign n1061 = n235 & n920;
  assign n1062 = ~n1060 & ~n1061;
  assign n1063 = ~pi01 & ~n312;
  assign n1064 = pi11 & ~n224;
  assign n1065 = ~n1063 & n1064;
  assign n1066 = ~n1057 & n1059;
  assign n1067 = ~pi05 & n120;
  assign n1068 = ~pi09 & ~n1067;
  assign n1069 = n1320 & n1068;
  assign n1070 = ~n1056 & n1069;
  assign n1071 = ~pi01 & ~n29;
  assign n1072 = pi05 & ~n891;
  assign n1073 = pi01 & ~n891;
  assign n1074 = ~n29 & ~n1073;
  assign n1075 = pi05 & ~n1074;
  assign n1076 = ~n1071 & n1072;
  assign n1077 = n55 & n240;
  assign n1078 = pi09 & ~n1077;
  assign n1079 = ~n1321 & n1078;
  assign n1080 = n1320 & ~n1067;
  assign n1081 = ~n1056 & ~n1067;
  assign n1082 = n1320 & n1081;
  assign n1083 = ~n1056 & n1080;
  assign n1084 = ~pi09 & ~n1322;
  assign n1085 = pi05 & n29;
  assign n1086 = n224 & ~n891;
  assign n1087 = ~n1077 & ~n1086;
  assign n1088 = ~n1085 & n1087;
  assign n1089 = ~n1321 & ~n1077;
  assign n1090 = pi09 & ~n1323;
  assign n1091 = ~n1084 & ~n1090;
  assign n1092 = ~n1070 & ~n1079;
  assign n1093 = pi05 & n40;
  assign n1094 = ~n1298 & ~n1093;
  assign n1095 = ~n261 & ~n1094;
  assign n1096 = pi11 & ~n132;
  assign n1097 = n1206 & ~n261;
  assign n1098 = ~n1096 & ~n1097;
  assign n1099 = pi01 & ~n1098;
  assign n1100 = ~n1095 & ~n1099;
  assign n1101 = n1324 & ~n1095;
  assign n1102 = ~n1099 & n1101;
  assign n1103 = ~n1090 & ~n1095;
  assign n1104 = ~n1099 & n1103;
  assign n1105 = ~n1084 & n1104;
  assign n1106 = n1324 & n1100;
  assign n1107 = ~pi13 & ~n1325;
  assign n1108 = n882 & ~n1107;
  assign n1109 = n1319 & n1108;
  assign n1110 = pi12 & n1209;
  assign n1111 = pi13 & ~n1210;
  assign n1112 = pi12 & n221;
  assign n1113 = ~pi12 & ~n221;
  assign n1114 = ~n1112 & ~n1113;
  assign n1115 = pi13 & ~n1114;
  assign n1116 = ~n1110 & n1111;
  assign n1117 = n60 & n1194;
  assign n1118 = ~pi00 & ~n29;
  assign n1119 = pi04 & ~n891;
  assign n1120 = ~n1118 & n1119;
  assign n1121 = n55 & n75;
  assign n1122 = pi09 & ~n1121;
  assign n1123 = ~n1120 & n1122;
  assign n1124 = ~n1117 & n1123;
  assign n1125 = n1193 & ~n884;
  assign n1126 = ~n120 & ~n139;
  assign n1127 = ~pi04 & ~n1126;
  assign n1128 = n88 & n920;
  assign n1129 = n133 & n169;
  assign n1130 = ~pi09 & ~n1327;
  assign n1131 = ~n1127 & n1130;
  assign n1132 = ~n1125 & n1131;
  assign n1133 = ~n1124 & ~n1132;
  assign n1134 = ~n132 & n139;
  assign n1135 = pi04 & n40;
  assign n1136 = ~n1298 & ~n1135;
  assign n1137 = ~n1193 & ~n1136;
  assign n1138 = ~n1134 & ~n1137;
  assign n1139 = n23 & ~n891;
  assign n1140 = pi04 & n29;
  assign n1141 = ~n1121 & ~n1140;
  assign n1142 = ~n1139 & n1141;
  assign n1143 = ~n1117 & ~n1139;
  assign n1144 = n1141 & n1143;
  assign n1145 = ~n1117 & n1142;
  assign n1146 = pi09 & ~n1328;
  assign n1147 = ~n1127 & ~n1327;
  assign n1148 = ~pi04 & n120;
  assign n1149 = ~n1125 & ~n1148;
  assign n1150 = pi11 & n89;
  assign n1151 = ~n1327 & ~n1150;
  assign n1152 = n1149 & n1151;
  assign n1153 = ~n1125 & n1147;
  assign n1154 = ~pi09 & ~n1329;
  assign n1155 = ~n1134 & ~n1154;
  assign n1156 = ~n1146 & n1155;
  assign n1157 = ~n1137 & n1156;
  assign n1158 = n1138 & ~n1154;
  assign n1159 = ~n1146 & n1158;
  assign n1160 = ~n1133 & n1138;
  assign n1161 = ~pi13 & ~n1330;
  assign n1162 = n882 & ~n1161;
  assign n1163 = ~n1326 & n1162;
  assign n1164 = n1191 & ~n1058;
  assign n1165 = ~n650 & ~po5;
  assign n1166 = n1255 & ~n1165;
  assign n1167 = n373 & n444;
  assign n1168 = ~pi06 & n554;
  assign n1169 = ~n1167 & ~n1168;
  assign n1170 = ~pi05 & ~n1169;
  assign n1171 = ~pi04 & n1170;
  assign n1172 = n1191 & n224;
  assign n1173 = ~n375 & ~n1172;
  assign n1174 = n1255 & ~n1173;
  assign n1175 = ~n1171 & ~n1174;
  assign n1176 = ~n1165 & ~n1175;
  assign n1177 = n1191 & n1255;
  assign n1178 = ~n1058 & ~n1165;
  assign n1179 = n1177 & n1178;
  assign n1180 = n1164 & n1166;
  assign n1181 = n31 | n32;
  assign n1182 = n33 | n34;
  assign n1183 = n38 | n39;
  assign n1184 = n42 | n43;
  assign n1185 = n49 | n50;
  assign n1186 = n56 | n57;
  assign n1187 = n64 | n65;
  assign n1188 = n67 | n68;
  assign n1189 = n72 | n73;
  assign n1190 = n84 | n85;
  assign n1191 = n90 | ~n91;
  assign n1192 = n96 | n97;
  assign n1193 = n104 | n105;
  assign n1194 = n109 | n110;
  assign n1195 = n116 | n117;
  assign n1196 = n122 | n123;
  assign n1197 = n127 | n128;
  assign n1198 = n130 | n131;
  assign n1199 = n135 | n136;
  assign n1200 = n144 | n145;
  assign n1201 = n149 | n147 | n148;
  assign n1202 = n155 | n156;
  assign n1203 = n159 | n160;
  assign n1204 = n162 | n163;
  assign n1205 = n186 | n183 | n185;
  assign n1206 = n187 | n188;
  assign n1207 = n190 | n191;
  assign n1208 = n194 | n195;
  assign n1209 = n219 | n214 | n218;
  assign n1210 = n222 | n223;
  assign n1211 = n228 | n229;
  assign n1212 = n247 | n248;
  assign n1213 = n251 | n252;
  assign n1214 = n259 | n260;
  assign n1215 = n263 | n264;
  assign n1216 = n280 | n281;
  assign n1217 = n290 | ~n291;
  assign n1218 = n298 | n299;
  assign n1219 = n306 | ~n307;
  assign n1220 = n310 | n311;
  assign n1221 = n320 | ~n321;
  assign n1222 = n331 | n328 | n330;
  assign n1223 = n339 | ~n340;
  assign n1224 = n343 | n344;
  assign n1225 = n354 | ~n355;
  assign n1226 = n363 | n364;
  assign n1227 = n385 | n386;
  assign n1228 = n401 | n402;
  assign n1229 = n404 | n405;
  assign n1230 = n408 | ~n409;
  assign n1231 = n412 | n413;
  assign n1232 = n416 | n417;
  assign n1233 = n434 | n427 | n433;
  assign n1234 = n439 | n440;
  assign n1235 = n442 | n443;
  assign n1236 = n453 | n454;
  assign n1237 = n473 | n474;
  assign n1238 = n492 | n489 | n491;
  assign n1239 = n498 | n499;
  assign n1240 = n504 | ~n505;
  assign n1241 = n508 | n509;
  assign n1242 = n524 | ~n525;
  assign n1243 = n532 | n529 | n531;
  assign n1244 = n534 | n535;
  assign n1245 = ~n543 | n540 | n542;
  assign n1246 = n546 | n547;
  assign n1247 = n566 | n567;
  assign n1248 = n569 | n570;
  assign n1249 = n571 | n572;
  assign n1250 = n580 | n581;
  assign n1251 = n584 | n585;
  assign n1252 = n586 | n587;
  assign n1253 = n592 | n593;
  assign n1254 = n596 | ~n597;
  assign n1255 = n603 | ~n604;
  assign n1256 = n610 | n611;
  assign n1257 = n613 | n614;
  assign n1258 = n627 | n628;
  assign n1259 = n639 | n640;
  assign n1260 = n642 | n643;
  assign n1261 = ~n649 | n646 | ~n648;
  assign n1262 = n653 | n654;
  assign n1263 = n659 | n660;
  assign n1264 = n668 | n669;
  assign n1265 = n674 | n675;
  assign n1266 = n680 | n681;
  assign n1267 = n688 | n689;
  assign n1268 = n693 | n694;
  assign n1269 = n703 | n704;
  assign n1270 = n721 | ~n722;
  assign n1271 = n726 | n727;
  assign n1272 = n731 | ~n732;
  assign n1273 = n735 | n736;
  assign n1274 = n739 | n740;
  assign n1275 = n753 | n748 | n752;
  assign n1276 = n760 | ~n761;
  assign n1277 = n763 | n764;
  assign n1278 = n769 | ~n770;
  assign n1279 = n774 | n775;
  assign n1280 = n782 | n783;
  assign n1281 = n788 | n789;
  assign n1282 = n797 | n798;
  assign n1283 = ~n806 | n803 | n805;
  assign n1284 = n811 | ~n812;
  assign n1285 = n818 | n819;
  assign n1286 = n825 | ~n826;
  assign n1287 = n827 | n828;
  assign n1288 = n830 | n831;
  assign n1289 = n838 | n839;
  assign n1290 = n843 | n844;
  assign n1291 = n848 | n849;
  assign n1292 = n861 | n862;
  assign n1293 = n864 | n865;
  assign n1294 = n870 | ~n871;
  assign n1295 = n877 | n874 | n876;
  assign n1296 = n880 | n881;
  assign n1297 = n901 | ~n902;
  assign n1298 = n909 | n906 | n908;
  assign n1299 = n922 | n923;
  assign n1300 = n925 | n926;
  assign n1301 = n934 | n931 | n933;
  assign n1302 = n942 | n943;
  assign n1303 = n945 | n946;
  assign n1304 = n953 | n949 | ~n952;
  assign n1305 = n957 | n958;
  assign n1306 = n962 | n963;
  assign n1307 = n968 | n969;
  assign n1308 = n974 | n975;
  assign n1309 = n978 | n979;
  assign n1310 = n983 | ~n984;
  assign n1311 = n986 | n987;
  assign n1312 = n992 | n993;
  assign n1313 = ~n1002 | n999 | ~n1001;
  assign n1314 = n1008 | n1009;
  assign n1315 = n1013 | n1014;
  assign n1316 = n1024 | n1025;
  assign n1317 = n1028 | ~n1029;
  assign n1318 = n1046 | n1041 | n1045;
  assign n1319 = n1054 | ~n1055;
  assign n1320 = ~n1066 | n1062 | ~n1065;
  assign n1321 = n1075 | n1076;
  assign n1322 = n1082 | n1083;
  assign n1323 = n1088 | n1089;
  assign n1324 = n1091 | ~n1092;
  assign n1325 = n1106 | n1102 | n1105;
  assign n1326 = n1115 | n1116;
  assign n1327 = n1128 | n1129;
  assign n1328 = n1144 | n1145;
  assign n1329 = n1152 | n1153;
  assign n1330 = n1160 | n1157 | n1159;
  assign po7 = n1180 | n1176 | n1179;
  assign po0 = ~n1163;
  assign po1 = ~n1109;
  assign po2 = ~n1049;
  assign po3 = ~n937;
  assign po4 = ~n1165;
endmodule
