module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n338, n339,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n417, n419, n420,
    n421, n422, n423, n424, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n439, n440, n441, n442, n443,
    n444, n445, n446, n448, n449, n450, n451,
    n452, n453, n454, n455, n456, n457, n458,
    n460, n461, n462, n463, n464, n465, n466,
    n468, n469, n470, n471, n472, n473, n475,
    n476, n477, n478, n479, n480, n481, n482,
    n484, n485, n486, n487, n488, n490, n491,
    n492, n493, n494, n496, n497, n498, n499,
    n500, n501, n502, n503, n505, n506, n507,
    n508, n509, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n527, n528, n529, n530,
    n531, n533, n534, n535, n536, n537, n539,
    n540, n541, n542, n543, n544, n546, n547,
    n548, n549, n551, n552, n553, n554, n555,
    n556, n557, n558, n559, n560, n562, n563,
    n564, n565, n567, n568, n569, n570, n571,
    n572, n573, n574, n576, n577, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602,
    n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n634, n635, n636, n637, n638,
    n639, n640, n642, n643, n644, n645, n646,
    n647, n648, n649, n650, n651, n653, n654,
    n655, n656, n657, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n717, n718, n719,
    n720, n721, n722, n724, n725, n726, n727,
    n728, n729, n731, n732, n733, n734, n735,
    n736, n738, n739, n740, n741, n742, n743,
    n745, n746, n747, n748, n749, n750, n752,
    n753, n754, n755, n756, n757, n759, n760,
    n761, n762, n763, n764, n766, n767, n768,
    n769, n770, n771, n773, n774, n775, n776,
    n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n796, n797, n798,
    n799, n800, n801, n802, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813,
    n814, n816, n817, n818, n819, n820, n821,
    n822, n823, n824, n825, n826, n827, n829,
    n830, n831, n832, n833, n834, n835, n836,
    n837, n838, n839, n840, n841, n842, n843,
    n844, n845, n846, n847, n848, n850, n851,
    n852, n853, n854, n855, n856, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881,
    n882, n883, n884, n885, n886, n888, n889,
    n890, n891, n892, n893, n894, n895, n896,
    n897, n898, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n910, n911, n912,
    n913, n914, n915, n916, n917, n918, n919,
    n920, n921, n923, n924, n925, n926, n927,
    n928, n929, n930, n931, n932, n933, n935,
    n936, n937, n938, n939, n940, n941, n943,
    n944, n945, n947, n948, n949, n951, n952,
    n953, n954, n958, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977,
    n978, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n997, n998, n999, n1000,
    n1001, n1002, n1004, n1005, n1006, n1007,
    n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1017, n1018, n1020,
    n1021, n1022, n1024, n1025, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1036, n1037, n1038, n1040, n1041, n1042,
    n1044, n1045, n1046, n1048, n1049, n1050,
    n1051, n1052, n1054, n1055, n1056, n1058,
    n1059, n1060, n1062, n1063, n1064, n1066,
    n1067, n1068, n1070, n1071, n1072, n1074,
    n1075, n1076, n1078, n1079, n1080, n1082,
    n1083, n1084, n1086, n1087, n1088, n1090,
    n1091, n1092, n1094, n1095, n1096, n1098,
    n1099, n1100, n1101, n1102, n1104, n1105,
    n1106, n1108, n1109, n1110, n1112, n1113,
    n1114, n1116, n1117, n1118, n1120, n1121,
    n1122, n1123, n1124, n1125, n1126, n1127,
    n1128, n1129, n1130, n1131, n1132, n1133,
    n1134, n1135, n1136, n1137, n1139, n1140,
    n1141, n1143, n1144, n1145, n1146, n1148,
    n1149, n1150, n1152, n1153, n1154, n1156,
    n1157, n1158, n1159, n1160, n1162, n1163,
    n1164, n1166, n1167, n1168, n1170, n1171,
    n1172, n1174, n1175, n1176, n1178, n1179,
    n1180, n1182, n1183, n1184, n1185, n1186,
    n1187, n1189, n1190, n1191, n1192, n1193,
    n1194, n1196, n1197, n1198, n1200, n1201,
    n1202, n1204, n1205, n1206, n1208, n1209,
    n1210, n1212, n1213, n1214, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223,
    n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1234, n1235, n1236,
    n1237, n1238, n1239, n1240, n1241, n1242,
    n1243, n1244, n1245, n1246, n1247, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255,
    n1256, n1257, n1258, n1259, n1260, n1261,
    n1262, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1297, n1298, n1299, n1301,
    n1302, n1303, n1304, n1305, n1306, n1307,
    n1308, n1309, n1310, n1311, n1312, n1313,
    n1314, n1315, n1316, n1317, n1319, n1320,
    n1321, n1322, n1323, n1324, n1325, n1326,
    n1327, n1328, n1329, n1330, n1331, n1332,
    n1333, n1334, n1335, n1337, n1338, n1340,
    n1341, n1343, n1344, n1345, n1346, n1348,
    n1349, n1350, n1351, n1353, n1354, n1355,
    n1356, n1358, n1359, n1360, n1361, n1363,
    n1364, n1365, n1368, n1369, n1372, n1373,
    n1375, n1380, n1381, n1383;
  assign n291 = ~pi8 & ~pi21;
  assign n292 = ~pi17 & n291;
  assign n293 = ~pi22 & n292;
  assign n294 = ~pi4 & ~pi19;
  assign n295 = ~pi18 & n294;
  assign n296 = ~pi16 & n295;
  assign n297 = ~pi9 & ~pi11;
  assign n298 = ~pi5 & ~pi7;
  assign n299 = ~pi6 & n298;
  assign n300 = ~pi13 & n299;
  assign n301 = ~pi12 & n300;
  assign n302 = ~pi14 & n301;
  assign n303 = n297 & n302;
  assign n304 = n296 & n303;
  assign n305 = n293 & n304;
  assign n306 = pi54 & ~n305;
  assign n307 = ~pi0 & ~n306;
  assign n308 = ~pi5 & ~pi22;
  assign n309 = pi56 & ~n308;
  assign n310 = ~pi7 & n291;
  assign n311 = ~pi13 & ~pi14;
  assign n312 = ~n310 & ~n311;
  assign n313 = ~pi13 & pi14;
  assign n314 = pi7 & ~n291;
  assign n315 = pi8 & pi21;
  assign n316 = ~n310 & ~n315;
  assign n317 = ~n314 & n316;
  assign n318 = ~pi13 & ~n317;
  assign n319 = ~pi14 & ~n318;
  assign n320 = ~n313 & ~n319;
  assign n321 = ~pi10 & ~n320;
  assign n322 = ~n312 & n321;
  assign n323 = pi10 & ~pi14;
  assign n324 = ~pi13 & n323;
  assign n325 = n310 & n324;
  assign n326 = ~n322 & ~n325;
  assign n327 = ~pi6 & ~pi12;
  assign n328 = ~pi17 & n296;
  assign n329 = n327 & n328;
  assign n330 = ~n326 & n329;
  assign n331 = n308 & ~n330;
  assign n332 = n297 & ~n331;
  assign n333 = ~n309 & n332;
  assign n334 = ~pi56 & ~n297;
  assign n335 = n308 & n334;
  assign n336 = ~n333 & ~n335;
  assign n337 = pi54 & ~n336;
  assign n338 = ~n307 & ~n337;
  assign n339 = ~pi3 & ~pi129;
  assign po15 = n338 | ~n339;
  assign n341 = ~pi10 & ~pi22;
  assign n342 = n311 & n341;
  assign n343 = ~pi11 & n291;
  assign n344 = ~pi12 & n296;
  assign n345 = n343 & n344;
  assign n346 = n299 & n345;
  assign n347 = n342 & n346;
  assign n348 = ~pi17 & ~n347;
  assign n349 = pi54 & n348;
  assign n350 = ~pi1 & ~n349;
  assign n351 = pi9 & ~n301;
  assign n352 = n341 & ~n351;
  assign n353 = ~pi14 & pi54;
  assign n354 = ~pi5 & n327;
  assign n355 = pi5 & ~n327;
  assign n356 = pi6 & pi12;
  assign n357 = ~n355 & ~n356;
  assign n358 = ~n354 & n357;
  assign n359 = ~pi7 & ~n358;
  assign n360 = pi7 & ~n354;
  assign n361 = ~pi13 & ~n360;
  assign n362 = ~n359 & n361;
  assign n363 = n298 & n327;
  assign n364 = pi13 & n363;
  assign n365 = ~pi9 & ~n364;
  assign n366 = ~n362 & n365;
  assign n367 = ~pi11 & n292;
  assign n368 = n296 & n367;
  assign n369 = ~n366 & n368;
  assign n370 = n353 & n369;
  assign n371 = n352 & n370;
  assign n372 = ~n350 & ~n371;
  assign po16 = ~n339 | n372;
  assign n374 = ~pi42 & ~pi44;
  assign n375 = ~pi40 & n374;
  assign n376 = ~pi46 & ~pi50;
  assign n377 = ~pi38 & n376;
  assign n378 = ~pi41 & ~pi43;
  assign n379 = n377 & n378;
  assign n380 = n375 & n379;
  assign n381 = pi82 & ~n380;
  assign n382 = pi122 & pi127;
  assign n383 = ~pi82 & n382;
  assign n384 = ~pi15 & ~pi20;
  assign n385 = ~pi24 & ~pi49;
  assign n386 = n384 & n385;
  assign n387 = ~pi45 & ~pi48;
  assign n388 = ~pi47 & n387;
  assign n389 = n386 & n388;
  assign n390 = pi82 & ~n389;
  assign n391 = ~n383 & ~n390;
  assign n392 = ~n381 & n391;
  assign n393 = pi2 & ~n392;
  assign n394 = n374 & n379;
  assign n395 = ~pi2 & n386;
  assign n396 = ~pi45 & n395;
  assign n397 = ~pi47 & n396;
  assign n398 = ~pi48 & n397;
  assign n399 = n394 & n398;
  assign n400 = pi82 & ~n399;
  assign n401 = ~n382 & ~n400;
  assign n402 = ~n381 & n401;
  assign n403 = ~pi65 & n402;
  assign n404 = ~n393 & ~n403;
  assign po17 = ~pi129 & ~n404;
  assign n406 = pi0 & ~pi123;
  assign n407 = ~pi113 & n406;
  assign n408 = ~pi17 & ~pi18;
  assign n409 = ~pi9 & ~pi22;
  assign n410 = ~pi10 & ~pi14;
  assign n411 = n409 & n410;
  assign n412 = n301 & n411;
  assign n413 = n345 & n412;
  assign n414 = n408 & n413;
  assign n415 = ~pi61 & ~n414;
  assign n416 = ~pi118 & n415;
  assign n417 = ~n407 & ~n416;
  assign po18 = ~pi129 & ~n417;
  assign n419 = pi4 & ~pi54;
  assign n420 = pi54 & n368;
  assign n421 = n323 & n409;
  assign n422 = n301 & n421;
  assign n423 = n420 & n422;
  assign n424 = ~n419 & ~n423;
  assign po19 = n339 & ~n424;
  assign n426 = pi5 & pi54;
  assign n427 = ~pi13 & n411;
  assign n428 = ~pi25 & n427;
  assign n429 = ~pi59 & n428;
  assign n430 = ~pi7 & ~pi12;
  assign n431 = ~pi6 & ~pi29;
  assign n432 = n430 & n431;
  assign n433 = pi28 & n432;
  assign n434 = n420 & n433;
  assign n435 = n429 & n434;
  assign n436 = ~pi5 & ~n435;
  assign n437 = n339 & ~n436;
  assign po20 = ~n426 & n437;
  assign n439 = pi6 & ~pi54;
  assign n440 = n420 & n427;
  assign n441 = pi25 & ~pi59;
  assign n442 = ~pi29 & n363;
  assign n443 = ~pi28 & n442;
  assign n444 = n441 & n443;
  assign n445 = n440 & n444;
  assign n446 = ~n439 & ~n445;
  assign po21 = n339 & ~n446;
  assign n448 = pi7 & ~pi54;
  assign n449 = ~pi11 & n408;
  assign n450 = n317 & n449;
  assign n451 = n354 & n450;
  assign n452 = ~pi16 & pi54;
  assign n453 = ~pi4 & n452;
  assign n454 = ~pi19 & n453;
  assign n455 = pi8 & n454;
  assign n456 = n427 & n455;
  assign n457 = n451 & n456;
  assign n458 = ~n448 & ~n457;
  assign po22 = n339 & ~n458;
  assign n460 = pi8 & ~pi54;
  assign n461 = ~pi8 & n449;
  assign n462 = n412 & n453;
  assign n463 = n461 & n462;
  assign n464 = ~pi19 & n463;
  assign n465 = pi21 & n464;
  assign n466 = ~n460 & ~n465;
  assign po23 = n339 & ~n466;
  assign n468 = pi9 & ~pi54;
  assign n469 = n295 & n452;
  assign n470 = pi11 & n412;
  assign n471 = n292 & n470;
  assign n472 = n469 & n471;
  assign n473 = ~n468 & ~n472;
  assign po24 = n339 & ~n473;
  assign n475 = pi10 & ~pi54;
  assign n476 = ~pi9 & ~pi10;
  assign n477 = ~pi11 & n476;
  assign n478 = n363 & n477;
  assign n479 = n293 & n478;
  assign n480 = n313 & n479;
  assign n481 = n469 & n480;
  assign n482 = ~n475 & ~n481;
  assign po25 = n339 & ~n482;
  assign n484 = pi11 & ~pi54;
  assign n485 = pi22 & n420;
  assign n486 = n302 & n485;
  assign n487 = n476 & n486;
  assign n488 = ~n484 & ~n487;
  assign po26 = n339 & ~n488;
  assign n490 = pi12 & ~pi54;
  assign n491 = pi18 & n412;
  assign n492 = n367 & n491;
  assign n493 = n454 & n492;
  assign n494 = ~n490 & ~n493;
  assign po27 = n339 & ~n494;
  assign n496 = pi13 & ~pi54;
  assign n497 = ~pi25 & ~pi28;
  assign n498 = pi29 & n497;
  assign n499 = pi54 & ~pi59;
  assign n500 = n498 & n499;
  assign n501 = n363 & n500;
  assign n502 = n440 & n501;
  assign n503 = ~n496 & ~n502;
  assign po28 = n339 & ~n503;
  assign n505 = pi14 & ~pi54;
  assign n506 = pi13 & n479;
  assign n507 = n296 & n506;
  assign n508 = n353 & n507;
  assign n509 = ~n505 & ~n508;
  assign po29 = n339 & ~n509;
  assign n511 = n380 & n388;
  assign n512 = n385 & n511;
  assign n513 = pi15 & ~n512;
  assign n514 = ~pi15 & n512;
  assign n515 = ~pi49 & n384;
  assign n516 = ~pi2 & n515;
  assign n517 = n514 & ~n516;
  assign n518 = ~n513 & ~n517;
  assign n519 = pi82 & ~n518;
  assign n520 = pi15 & n383;
  assign n521 = ~n519 & ~n520;
  assign n522 = pi82 & ~n514;
  assign n523 = ~pi70 & ~n522;
  assign n524 = ~n382 & n523;
  assign n525 = n521 & ~n524;
  assign po30 = ~pi129 & ~n525;
  assign n527 = pi16 & ~pi54;
  assign n528 = pi6 & n420;
  assign n529 = n362 & n528;
  assign n530 = n411 & n529;
  assign n531 = ~n527 & ~n530;
  assign po31 = n339 & ~n531;
  assign n533 = pi17 & ~pi54;
  assign n534 = pi59 & n443;
  assign n535 = n420 & n534;
  assign n536 = n428 & n535;
  assign n537 = ~n533 & ~n536;
  assign po32 = n339 & ~n537;
  assign n539 = pi18 & ~pi54;
  assign n540 = pi16 & n367;
  assign n541 = pi54 & n540;
  assign n542 = n295 & n541;
  assign n543 = n412 & n542;
  assign n544 = ~n539 & ~n543;
  assign po33 = n339 & ~n544;
  assign n546 = pi19 & ~pi54;
  assign n547 = pi17 & pi54;
  assign n548 = n413 & n547;
  assign n549 = ~n546 & ~n548;
  assign po34 = n339 & ~n549;
  assign n551 = n384 & n512;
  assign n552 = pi2 & n551;
  assign n553 = pi20 & ~n514;
  assign n554 = ~n552 & ~n553;
  assign n555 = pi82 & ~n554;
  assign n556 = pi20 & n383;
  assign n557 = ~n555 & ~n556;
  assign n558 = ~pi71 & ~n382;
  assign n559 = n392 & n558;
  assign n560 = n557 & ~n559;
  assign po35 = ~pi129 & ~n560;
  assign n562 = pi21 & ~pi54;
  assign n563 = ~pi21 & n463;
  assign n564 = pi19 & n563;
  assign n565 = ~n562 & ~n564;
  assign po36 = n339 & ~n565;
  assign n567 = pi22 & ~pi54;
  assign n568 = pi5 & ~pi7;
  assign n569 = n311 & n568;
  assign n570 = n293 & n569;
  assign n571 = n327 & n477;
  assign n572 = n469 & n571;
  assign n573 = n570 & n572;
  assign n574 = ~n567 & ~n573;
  assign po37 = n339 & ~n574;
  assign n576 = ~pi23 & pi55;
  assign n577 = pi61 & ~n576;
  assign po38 = ~pi129 & n577;
  assign n579 = pi82 & ~n511;
  assign n580 = pi82 & ~n516;
  assign n581 = n382 & ~n580;
  assign n582 = ~n579 & ~n581;
  assign n583 = pi63 & ~n580;
  assign n584 = n582 & n583;
  assign n585 = ~pi24 & ~n582;
  assign n586 = pi24 & pi82;
  assign n587 = n511 & n586;
  assign n588 = ~pi129 & ~n587;
  assign n589 = ~n585 & n588;
  assign po39 = ~n584 & n589;
  assign n591 = ~pi96 & ~pi110;
  assign n592 = ~pi85 & ~n591;
  assign n593 = pi85 & ~pi116;
  assign n594 = pi100 & ~n593;
  assign n595 = ~n592 & n594;
  assign n596 = pi25 & ~pi116;
  assign n597 = pi85 & n596;
  assign n598 = ~n595 & ~n597;
  assign n599 = ~pi26 & ~n598;
  assign n600 = ~pi95 & ~pi100;
  assign n601 = ~pi97 & n600;
  assign n602 = ~pi110 & ~n601;
  assign n603 = pi25 & ~n602;
  assign n604 = pi26 & pi116;
  assign n605 = ~n603 & ~n604;
  assign n606 = ~pi39 & ~pi52;
  assign n607 = ~pi51 & n606;
  assign n608 = ~n605 & ~n607;
  assign n609 = pi26 & n596;
  assign n610 = ~n608 & ~n609;
  assign n611 = ~pi85 & ~n610;
  assign n612 = ~n599 & ~n611;
  assign n613 = ~pi27 & ~n612;
  assign n614 = pi116 & n607;
  assign n615 = ~n596 & ~n614;
  assign n616 = pi27 & ~n615;
  assign n617 = n603 & n607;
  assign n618 = ~n616 & ~n617;
  assign n619 = ~pi26 & ~pi85;
  assign n620 = ~n618 & n619;
  assign n621 = ~n613 & ~n620;
  assign n622 = ~pi53 & ~n621;
  assign n623 = pi53 & ~pi85;
  assign n624 = ~pi26 & ~pi27;
  assign n625 = n596 & n624;
  assign n626 = n623 & n625;
  assign n627 = ~n622 & ~n626;
  assign n628 = ~pi58 & ~n627;
  assign n629 = ~pi53 & pi58;
  assign n630 = n619 & n629;
  assign n631 = n625 & n630;
  assign n632 = ~n628 & ~n631;
  assign po40 = n339 & ~n632;
  assign n634 = ~pi53 & ~pi58;
  assign n635 = ~pi27 & n634;
  assign n636 = ~pi85 & ~n614;
  assign n637 = pi26 & n636;
  assign n638 = n595 & ~n604;
  assign n639 = ~n637 & ~n638;
  assign n640 = n339 & ~n639;
  assign po41 = n635 & n640;
  assign n642 = pi27 & n636;
  assign n643 = pi95 & n591;
  assign n644 = ~pi85 & ~n643;
  assign n645 = ~pi100 & ~n644;
  assign n646 = pi27 & pi116;
  assign n647 = ~n593 & ~n646;
  assign n648 = n645 & n647;
  assign n649 = ~n642 & ~n648;
  assign n650 = n634 & ~n649;
  assign n651 = ~pi26 & n339;
  assign po42 = n650 & n651;
  assign n653 = ~pi26 & n643;
  assign n654 = ~pi100 & n653;
  assign n655 = n604 & n607;
  assign n656 = ~n654 & ~n655;
  assign n657 = ~pi27 & ~n656;
  assign n658 = ~pi26 & ~n607;
  assign n659 = ~pi27 & n607;
  assign n660 = ~n658 & ~n659;
  assign n661 = ~n602 & ~n660;
  assign n662 = pi26 & ~pi27;
  assign n663 = ~pi26 & pi27;
  assign n664 = ~n662 & ~n663;
  assign n665 = ~pi116 & ~n664;
  assign n666 = ~n661 & ~n665;
  assign n667 = pi28 & ~n666;
  assign n668 = n646 & n658;
  assign n669 = ~n667 & ~n668;
  assign n670 = ~n657 & n669;
  assign n671 = ~pi85 & ~n670;
  assign n672 = ~pi28 & ~pi116;
  assign n673 = pi85 & ~n672;
  assign n674 = pi100 & pi116;
  assign n675 = n624 & ~n674;
  assign n676 = n673 & n675;
  assign n677 = ~n671 & ~n676;
  assign n678 = ~pi53 & ~n677;
  assign n679 = ~pi27 & pi28;
  assign n680 = ~pi116 & n679;
  assign n681 = ~pi26 & n623;
  assign n682 = n680 & n681;
  assign n683 = ~n678 & ~n682;
  assign n684 = ~pi58 & ~n683;
  assign n685 = n630 & n680;
  assign n686 = ~n684 & ~n685;
  assign po43 = n339 & ~n686;
  assign n688 = pi53 & ~pi58;
  assign n689 = ~n629 & ~n688;
  assign n690 = ~pi116 & ~n689;
  assign n691 = ~n602 & n634;
  assign n692 = ~n690 & ~n691;
  assign n693 = pi29 & ~n692;
  assign n694 = pi58 & pi116;
  assign n695 = ~pi58 & n591;
  assign n696 = n600 & n695;
  assign n697 = ~n694 & ~n696;
  assign n698 = ~pi53 & pi97;
  assign n699 = ~n697 & n698;
  assign n700 = ~n693 & ~n699;
  assign n701 = ~pi27 & ~n700;
  assign n702 = pi29 & ~pi116;
  assign n703 = pi27 & n702;
  assign n704 = n634 & n703;
  assign n705 = ~n701 & ~n704;
  assign n706 = ~pi85 & ~n705;
  assign n707 = pi85 & n634;
  assign n708 = ~pi27 & n707;
  assign n709 = n702 & n708;
  assign n710 = ~n706 & ~n709;
  assign n711 = ~pi26 & ~n710;
  assign n712 = ~pi85 & n634;
  assign n713 = n662 & n712;
  assign n714 = n702 & n713;
  assign n715 = ~n711 & ~n714;
  assign po44 = n339 & ~n715;
  assign n717 = pi30 & ~pi109;
  assign n718 = pi60 & pi109;
  assign n719 = ~pi106 & ~n718;
  assign n720 = ~n717 & n719;
  assign n721 = ~pi88 & pi106;
  assign n722 = ~pi129 & ~n721;
  assign po45 = ~n720 & n722;
  assign n724 = pi31 & ~pi109;
  assign n725 = pi30 & pi109;
  assign n726 = ~pi106 & ~n725;
  assign n727 = ~n724 & n726;
  assign n728 = ~pi89 & pi106;
  assign n729 = ~pi129 & ~n728;
  assign po46 = ~n727 & n729;
  assign n731 = pi32 & ~pi109;
  assign n732 = pi31 & pi109;
  assign n733 = ~pi106 & ~n732;
  assign n734 = ~n731 & n733;
  assign n735 = ~pi99 & pi106;
  assign n736 = ~pi129 & ~n735;
  assign po47 = ~n734 & n736;
  assign n738 = pi33 & ~pi109;
  assign n739 = pi32 & pi109;
  assign n740 = ~pi106 & ~n739;
  assign n741 = ~n738 & n740;
  assign n742 = ~pi90 & pi106;
  assign n743 = ~pi129 & ~n742;
  assign po48 = ~n741 & n743;
  assign n745 = pi34 & ~pi109;
  assign n746 = pi33 & pi109;
  assign n747 = ~pi106 & ~n746;
  assign n748 = ~n745 & n747;
  assign n749 = ~pi91 & pi106;
  assign n750 = ~pi129 & ~n749;
  assign po49 = ~n748 & n750;
  assign n752 = pi35 & ~pi109;
  assign n753 = pi34 & pi109;
  assign n754 = ~pi106 & ~n753;
  assign n755 = ~n752 & n754;
  assign n756 = ~pi92 & pi106;
  assign n757 = ~pi129 & ~n756;
  assign po50 = ~n755 & n757;
  assign n759 = pi36 & ~pi109;
  assign n760 = pi35 & pi109;
  assign n761 = ~pi106 & ~n760;
  assign n762 = ~n759 & n761;
  assign n763 = ~pi98 & pi106;
  assign n764 = ~pi129 & ~n763;
  assign po51 = ~n762 & n764;
  assign n766 = pi37 & ~pi109;
  assign n767 = pi36 & pi109;
  assign n768 = ~pi106 & ~n767;
  assign n769 = ~n766 & n768;
  assign n770 = ~pi93 & pi106;
  assign n771 = ~pi129 & ~n770;
  assign po52 = ~n769 & n771;
  assign n773 = pi82 & ~n375;
  assign n774 = ~pi43 & ~pi47;
  assign n775 = ~pi48 & n396;
  assign n776 = n774 & n775;
  assign n777 = pi82 & ~n776;
  assign n778 = n382 & ~n777;
  assign n779 = ~pi41 & n376;
  assign n780 = n391 & ~n779;
  assign n781 = n778 & ~n780;
  assign n782 = ~n773 & ~n781;
  assign n783 = ~pi38 & ~n782;
  assign n784 = ~pi38 & n375;
  assign n785 = pi82 & ~n784;
  assign n786 = n375 & n785;
  assign n787 = ~pi129 & ~n786;
  assign n788 = n378 & n398;
  assign n789 = n375 & n788;
  assign n790 = n376 & n789;
  assign n791 = pi82 & ~n790;
  assign n792 = ~n382 & ~n791;
  assign n793 = pi74 & n792;
  assign n794 = n787 & ~n793;
  assign po53 = ~n783 & n794;
  assign n796 = ~pi51 & ~pi52;
  assign n797 = pi109 & n796;
  assign n798 = pi39 & ~n797;
  assign n799 = ~pi51 & pi109;
  assign n800 = n606 & n799;
  assign n801 = ~pi106 & ~n800;
  assign n802 = ~n798 & n801;
  assign po54 = ~pi129 & ~n802;
  assign n804 = n374 & n773;
  assign n805 = pi82 & ~n374;
  assign n806 = pi82 & ~n398;
  assign n807 = n382 & ~n806;
  assign n808 = ~n379 & n391;
  assign n809 = n807 & ~n808;
  assign n810 = ~n805 & ~n809;
  assign n811 = ~pi40 & ~n810;
  assign n812 = pi73 & n401;
  assign n813 = ~pi129 & ~n812;
  assign n814 = ~n811 & n813;
  assign po55 = ~n804 & n814;
  assign n816 = n375 & n377;
  assign n817 = n776 & n816;
  assign n818 = pi82 & ~n817;
  assign n819 = ~n382 & ~n818;
  assign n820 = pi76 & n819;
  assign n821 = ~pi41 & n816;
  assign n822 = pi82 & ~n821;
  assign n823 = n816 & n822;
  assign n824 = ~pi129 & ~n823;
  assign n825 = ~n820 & n824;
  assign n826 = ~n778 & ~n822;
  assign n827 = ~pi41 & ~n826;
  assign po56 = n825 & ~n827;
  assign n829 = pi44 & pi82;
  assign n830 = ~pi38 & ~pi40;
  assign n831 = ~pi50 & n830;
  assign n832 = ~pi44 & n831;
  assign n833 = ~pi47 & n378;
  assign n834 = ~pi46 & n833;
  assign n835 = ~pi48 & n834;
  assign n836 = n395 & n835;
  assign n837 = ~pi45 & n836;
  assign n838 = n832 & n837;
  assign n839 = pi82 & ~n838;
  assign n840 = n382 & ~n839;
  assign n841 = ~n829 & ~n840;
  assign n842 = ~pi42 & ~n841;
  assign n843 = ~pi44 & pi82;
  assign n844 = pi42 & n843;
  assign n845 = ~pi129 & ~n844;
  assign n846 = ~n382 & ~n839;
  assign n847 = pi72 & n846;
  assign n848 = n845 & ~n847;
  assign po57 = ~n842 & n848;
  assign n850 = ~n807 & ~n822;
  assign n851 = ~pi43 & ~n850;
  assign n852 = ~n806 & n850;
  assign n853 = pi77 & n852;
  assign n854 = n381 & n821;
  assign n855 = ~pi129 & ~n854;
  assign n856 = ~n853 & n855;
  assign po58 = ~n851 & n856;
  assign n858 = ~pi42 & n834;
  assign n859 = n775 & n831;
  assign n860 = n858 & n859;
  assign n861 = pi82 & ~n860;
  assign n862 = ~pi67 & ~n382;
  assign n863 = pi44 & n382;
  assign n864 = ~n862 & ~n863;
  assign n865 = ~n861 & n864;
  assign n866 = ~pi129 & ~n829;
  assign po59 = ~n865 & n866;
  assign n868 = pi82 & ~n395;
  assign n869 = n382 & ~n868;
  assign n870 = n774 & n779;
  assign n871 = n843 & n870;
  assign n872 = pi48 & n871;
  assign n873 = ~n869 & ~n872;
  assign n874 = pi47 & pi82;
  assign n875 = ~n381 & ~n874;
  assign n876 = n873 & n875;
  assign n877 = ~pi45 & ~n876;
  assign n878 = n374 & n831;
  assign n879 = n836 & n878;
  assign n880 = pi82 & ~n879;
  assign n881 = ~n382 & ~n880;
  assign n882 = pi68 & n881;
  assign n883 = n835 & n878;
  assign n884 = n579 & n883;
  assign n885 = ~pi129 & ~n884;
  assign n886 = ~n882 & n885;
  assign po60 = ~n877 & n886;
  assign n888 = pi82 & ~n878;
  assign n889 = pi82 & ~n788;
  assign n890 = n382 & ~n889;
  assign n891 = ~n888 & ~n890;
  assign n892 = pi75 & ~n889;
  assign n893 = n891 & n892;
  assign n894 = pi82 & n878;
  assign n895 = pi46 & n894;
  assign n896 = ~pi46 & ~n891;
  assign n897 = ~pi129 & ~n896;
  assign n898 = ~n895 & n897;
  assign po61 = ~n893 & n898;
  assign n900 = pi82 & ~n775;
  assign n901 = n382 & ~n900;
  assign n902 = ~n381 & ~n901;
  assign n903 = pi64 & ~n900;
  assign n904 = n902 & n903;
  assign n905 = ~pi47 & ~n902;
  assign n906 = ~pi129 & ~n905;
  assign n907 = ~n904 & n906;
  assign n908 = n380 & n874;
  assign po62 = n907 & ~n908;
  assign n910 = pi82 & ~n837;
  assign n911 = n382 & ~n910;
  assign n912 = n875 & ~n911;
  assign n913 = ~pi48 & ~n912;
  assign n914 = n380 & n397;
  assign n915 = pi82 & ~n914;
  assign n916 = ~n382 & ~n915;
  assign n917 = pi62 & n916;
  assign n918 = ~pi42 & n830;
  assign n919 = n872 & n918;
  assign n920 = ~pi129 & ~n919;
  assign n921 = ~n917 & n920;
  assign po63 = ~n913 & n921;
  assign n923 = ~pi24 & n511;
  assign n924 = pi49 & ~n923;
  assign n925 = n512 & ~n775;
  assign n926 = ~n924 & ~n925;
  assign n927 = pi82 & ~n926;
  assign n928 = pi49 & n383;
  assign n929 = ~n927 & ~n928;
  assign n930 = pi82 & ~n512;
  assign n931 = ~pi69 & ~n930;
  assign n932 = ~n382 & n931;
  assign n933 = n929 & ~n932;
  assign po64 = ~pi129 & ~n933;
  assign n935 = ~n785 & ~n911;
  assign n936 = ~pi50 & ~n935;
  assign n937 = ~n785 & n888;
  assign n938 = ~pi129 & ~n937;
  assign n939 = pi66 & ~n910;
  assign n940 = n935 & n939;
  assign n941 = n938 & ~n940;
  assign po65 = ~n936 & n941;
  assign n943 = pi51 & ~pi109;
  assign n944 = ~pi106 & ~n799;
  assign n945 = ~n943 & n944;
  assign po66 = ~pi129 & ~n945;
  assign n947 = pi52 & ~n799;
  assign n948 = ~pi106 & ~n797;
  assign n949 = ~n947 & n948;
  assign po67 = ~pi129 & ~n949;
  assign n951 = ~pi116 & n688;
  assign n952 = ~n699 & ~n951;
  assign n953 = n339 & ~n952;
  assign n954 = ~pi85 & n953;
  assign po68 = n624 & n954;
  assign po69 = pi129 | n402;
  assign po129 = pi123 | pi129;
  assign n958 = pi114 & ~pi122;
  assign po70 = ~po129 & n958;
  assign n960 = ~pi26 & pi58;
  assign n961 = n604 & ~n694;
  assign n962 = ~n960 & ~n961;
  assign n963 = pi94 & ~n962;
  assign n964 = pi58 & ~pi116;
  assign n965 = pi37 & ~pi116;
  assign n966 = ~n960 & ~n965;
  assign n967 = ~n964 & ~n966;
  assign n968 = ~n963 & ~n967;
  assign n969 = ~pi53 & ~n968;
  assign n970 = ~pi26 & pi37;
  assign n971 = ~pi58 & n970;
  assign n972 = ~n969 & ~n971;
  assign n973 = ~pi85 & ~n972;
  assign n974 = n634 & n970;
  assign n975 = ~n973 & ~n974;
  assign n976 = ~pi27 & ~n975;
  assign n977 = n712 & n970;
  assign n978 = ~n976 & ~n977;
  assign po71 = n339 & ~n978;
  assign n980 = ~pi26 & ~pi53;
  assign n981 = ~pi85 & n980;
  assign n982 = ~pi116 & n981;
  assign n983 = pi26 & pi53;
  assign n984 = pi85 & ~n980;
  assign n985 = ~pi58 & ~n984;
  assign n986 = ~n983 & n985;
  assign n987 = ~n982 & ~n986;
  assign n988 = pi57 & ~n987;
  assign n989 = pi60 & n630;
  assign n990 = pi116 & n989;
  assign n991 = ~n988 & ~n990;
  assign n992 = ~pi27 & ~n991;
  assign n993 = pi57 & ~pi58;
  assign n994 = n981 & n993;
  assign n995 = ~n992 & ~n994;
  assign po72 = n339 & ~n995;
  assign n997 = n624 & n964;
  assign n998 = ~pi58 & ~n664;
  assign n999 = n614 & n998;
  assign n1000 = ~n997 & ~n999;
  assign n1001 = ~pi53 & ~n1000;
  assign n1002 = ~pi85 & n339;
  assign po73 = n1001 & n1002;
  assign n1004 = pi59 & ~n692;
  assign n1005 = pi96 & n634;
  assign n1006 = n602 & n1005;
  assign n1007 = ~n1004 & ~n1006;
  assign n1008 = ~pi85 & ~n1007;
  assign n1009 = pi59 & ~pi116;
  assign n1010 = n707 & n1009;
  assign n1011 = ~n1008 & ~n1010;
  assign n1012 = ~pi27 & ~n1011;
  assign n1013 = pi27 & n712;
  assign n1014 = n1009 & n1013;
  assign n1015 = ~n1012 & ~n1014;
  assign n1016 = ~pi26 & ~n1015;
  assign n1017 = n713 & n1009;
  assign n1018 = ~n1016 & ~n1017;
  assign po74 = n339 & ~n1018;
  assign n1020 = ~pi117 & ~pi122;
  assign n1021 = pi60 & ~n1020;
  assign n1022 = pi123 & n1020;
  assign po75 = n1021 | n1022;
  assign n1024 = ~pi114 & ~pi129;
  assign n1025 = ~pi122 & pi123;
  assign po76 = n1024 & n1025;
  assign n1027 = pi136 & ~pi137;
  assign n1028 = pi132 & pi133;
  assign n1029 = pi131 & n1028;
  assign n1030 = ~pi138 & n1029;
  assign n1031 = n1027 & n1030;
  assign n1032 = ~pi62 & ~n1031;
  assign n1033 = pi140 & n1031;
  assign n1034 = ~pi129 & ~n1033;
  assign po77 = n1032 | ~n1034;
  assign n1036 = ~pi63 & ~n1031;
  assign n1037 = pi142 & n1031;
  assign n1038 = ~pi129 & ~n1037;
  assign po78 = n1036 | ~n1038;
  assign n1040 = ~pi64 & ~n1031;
  assign n1041 = pi139 & n1031;
  assign n1042 = ~pi129 & ~n1041;
  assign po79 = n1040 | ~n1042;
  assign n1044 = ~pi65 & ~n1031;
  assign n1045 = pi146 & n1031;
  assign n1046 = ~pi129 & ~n1045;
  assign po80 = n1044 | ~n1046;
  assign n1048 = ~pi136 & ~pi137;
  assign n1049 = n1030 & n1048;
  assign n1050 = ~pi66 & ~n1049;
  assign n1051 = pi143 & n1049;
  assign n1052 = ~pi129 & ~n1051;
  assign po81 = n1050 | ~n1052;
  assign n1054 = ~pi67 & ~n1049;
  assign n1055 = pi139 & n1049;
  assign n1056 = ~pi129 & ~n1055;
  assign po82 = n1054 | ~n1056;
  assign n1058 = ~pi68 & ~n1031;
  assign n1059 = pi141 & n1031;
  assign n1060 = ~pi129 & ~n1059;
  assign po83 = n1058 | ~n1060;
  assign n1062 = ~pi69 & ~n1031;
  assign n1063 = pi143 & n1031;
  assign n1064 = ~pi129 & ~n1063;
  assign po84 = n1062 | ~n1064;
  assign n1066 = ~pi70 & ~n1031;
  assign n1067 = pi144 & n1031;
  assign n1068 = ~pi129 & ~n1067;
  assign po85 = n1066 | ~n1068;
  assign n1070 = ~pi71 & ~n1031;
  assign n1071 = pi145 & n1031;
  assign n1072 = ~pi129 & ~n1071;
  assign po86 = n1070 | ~n1072;
  assign n1074 = ~pi72 & ~n1049;
  assign n1075 = pi140 & n1049;
  assign n1076 = ~pi129 & ~n1075;
  assign po87 = n1074 | ~n1076;
  assign n1078 = ~pi73 & ~n1049;
  assign n1079 = pi141 & n1049;
  assign n1080 = ~pi129 & ~n1079;
  assign po88 = n1078 | ~n1080;
  assign n1082 = ~pi74 & ~n1049;
  assign n1083 = pi142 & n1049;
  assign n1084 = ~pi129 & ~n1083;
  assign po89 = n1082 | ~n1084;
  assign n1086 = ~pi75 & ~n1049;
  assign n1087 = pi144 & n1049;
  assign n1088 = ~pi129 & ~n1087;
  assign po90 = n1086 | ~n1088;
  assign n1090 = ~pi76 & ~n1049;
  assign n1091 = pi145 & n1049;
  assign n1092 = ~pi129 & ~n1091;
  assign po91 = n1090 | ~n1092;
  assign n1094 = ~pi77 & ~n1049;
  assign n1095 = pi146 & n1049;
  assign n1096 = ~pi129 & ~n1095;
  assign po92 = n1094 | ~n1096;
  assign n1098 = ~pi136 & pi137;
  assign n1099 = n1030 & n1098;
  assign n1100 = ~pi78 & ~n1099;
  assign n1101 = ~pi142 & n1099;
  assign n1102 = ~pi129 & ~n1101;
  assign po93 = ~n1100 & n1102;
  assign n1104 = ~pi79 & ~n1099;
  assign n1105 = ~pi143 & n1099;
  assign n1106 = ~pi129 & ~n1105;
  assign po94 = ~n1104 & n1106;
  assign n1108 = ~pi80 & ~n1099;
  assign n1109 = ~pi144 & n1099;
  assign n1110 = ~pi129 & ~n1109;
  assign po95 = ~n1108 & n1110;
  assign n1112 = ~pi81 & ~n1099;
  assign n1113 = ~pi145 & n1099;
  assign n1114 = ~pi129 & ~n1113;
  assign po96 = ~n1112 & n1114;
  assign n1116 = ~pi82 & ~n1099;
  assign n1117 = ~pi146 & n1099;
  assign n1118 = ~pi129 & ~n1117;
  assign po97 = ~n1116 & n1118;
  assign n1120 = ~pi89 & pi138;
  assign n1121 = pi62 & ~pi138;
  assign n1122 = pi136 & ~n1121;
  assign n1123 = ~n1120 & n1122;
  assign n1124 = ~pi119 & pi138;
  assign n1125 = pi72 & ~pi138;
  assign n1126 = ~pi136 & ~n1125;
  assign n1127 = ~n1124 & n1126;
  assign n1128 = ~n1123 & ~n1127;
  assign n1129 = ~pi137 & ~n1128;
  assign n1130 = pi136 & ~pi138;
  assign n1131 = pi31 & n1130;
  assign n1132 = ~pi87 & ~pi138;
  assign n1133 = pi115 & pi138;
  assign n1134 = ~pi136 & ~n1133;
  assign n1135 = ~n1132 & n1134;
  assign n1136 = ~n1131 & ~n1135;
  assign n1137 = pi137 & ~n1136;
  assign po98 = n1129 | n1137;
  assign n1139 = ~pi84 & ~n1099;
  assign n1140 = ~pi141 & n1099;
  assign n1141 = ~pi129 & ~n1140;
  assign po99 = ~n1139 & n1141;
  assign n1143 = n592 & n602;
  assign n1144 = ~n593 & ~n1143;
  assign n1145 = n624 & n634;
  assign n1146 = n339 & n1145;
  assign po100 = ~n1144 & n1146;
  assign n1148 = ~pi86 & ~n1099;
  assign n1149 = ~pi139 & n1099;
  assign n1150 = ~pi129 & ~n1149;
  assign po101 = ~n1148 & n1150;
  assign n1152 = ~pi87 & ~n1099;
  assign n1153 = ~pi140 & n1099;
  assign n1154 = ~pi129 & ~n1153;
  assign po102 = ~n1152 & n1154;
  assign n1156 = pi137 & n1130;
  assign n1157 = n1029 & n1156;
  assign n1158 = ~pi88 & ~n1157;
  assign n1159 = ~pi139 & n1157;
  assign n1160 = ~pi129 & ~n1159;
  assign po103 = ~n1158 & n1160;
  assign n1162 = ~pi89 & ~n1157;
  assign n1163 = ~pi140 & n1157;
  assign n1164 = ~pi129 & ~n1163;
  assign po104 = ~n1162 & n1164;
  assign n1166 = ~pi90 & ~n1157;
  assign n1167 = ~pi142 & n1157;
  assign n1168 = ~pi129 & ~n1167;
  assign po105 = ~n1166 & n1168;
  assign n1170 = ~pi91 & ~n1157;
  assign n1171 = ~pi143 & n1157;
  assign n1172 = ~pi129 & ~n1171;
  assign po106 = ~n1170 & n1172;
  assign n1174 = ~pi92 & ~n1157;
  assign n1175 = ~pi144 & n1157;
  assign n1176 = ~pi129 & ~n1175;
  assign po107 = ~n1174 & n1176;
  assign n1178 = ~pi93 & ~n1157;
  assign n1179 = ~pi146 & n1157;
  assign n1180 = ~pi129 & ~n1179;
  assign po108 = ~n1178 & n1180;
  assign n1182 = pi82 & pi138;
  assign n1183 = n1048 & n1182;
  assign n1184 = n1029 & n1183;
  assign n1185 = ~pi94 & ~n1184;
  assign n1186 = ~pi142 & n1184;
  assign n1187 = ~pi129 & ~n1186;
  assign po109 = ~n1185 & n1187;
  assign n1189 = ~pi3 & ~pi110;
  assign n1190 = ~n1029 & ~n1189;
  assign n1191 = ~n1184 & ~n1190;
  assign n1192 = pi95 & n1191;
  assign n1193 = pi143 & n1184;
  assign n1194 = ~n1192 & ~n1193;
  assign po110 = ~pi129 & ~n1194;
  assign n1196 = pi96 & n1191;
  assign n1197 = pi146 & n1184;
  assign n1198 = ~n1196 & ~n1197;
  assign po111 = ~pi129 & ~n1198;
  assign n1200 = pi97 & n1191;
  assign n1201 = pi145 & n1184;
  assign n1202 = ~n1200 & ~n1201;
  assign po112 = ~pi129 & ~n1202;
  assign n1204 = ~pi98 & ~n1157;
  assign n1205 = ~pi145 & n1157;
  assign n1206 = ~pi129 & ~n1205;
  assign po113 = ~n1204 & n1206;
  assign n1208 = ~pi99 & ~n1157;
  assign n1209 = ~pi141 & n1157;
  assign n1210 = ~pi129 & ~n1209;
  assign po114 = ~n1208 & n1210;
  assign n1212 = pi100 & n1191;
  assign n1213 = pi144 & n1184;
  assign n1214 = ~n1212 & ~n1213;
  assign po115 = ~pi129 & ~n1214;
  assign n1216 = ~pi124 & pi138;
  assign n1217 = pi77 & ~pi138;
  assign n1218 = ~pi136 & ~n1217;
  assign n1219 = ~n1216 & n1218;
  assign n1220 = ~pi93 & pi138;
  assign n1221 = pi65 & ~pi138;
  assign n1222 = pi136 & ~n1221;
  assign n1223 = ~n1220 & n1222;
  assign n1224 = ~n1219 & ~n1223;
  assign n1225 = ~pi137 & ~n1224;
  assign n1226 = pi37 & n1130;
  assign n1227 = ~pi82 & ~pi138;
  assign n1228 = ~pi96 & pi138;
  assign n1229 = ~pi136 & ~n1228;
  assign n1230 = ~n1227 & n1229;
  assign n1231 = ~n1226 & ~n1230;
  assign n1232 = pi137 & ~n1231;
  assign po116 = n1225 | n1232;
  assign n1234 = pi91 & n1027;
  assign n1235 = pi95 & n1098;
  assign n1236 = ~n1234 & ~n1235;
  assign n1237 = pi138 & ~n1236;
  assign n1238 = ~pi79 & ~pi136;
  assign n1239 = ~pi34 & pi136;
  assign n1240 = pi137 & ~n1239;
  assign n1241 = ~n1238 & n1240;
  assign n1242 = pi66 & ~pi136;
  assign n1243 = pi69 & pi136;
  assign n1244 = ~pi137 & ~n1243;
  assign n1245 = ~n1242 & n1244;
  assign n1246 = ~n1241 & ~n1245;
  assign n1247 = ~pi138 & ~n1246;
  assign po117 = n1237 | n1247;
  assign n1249 = pi90 & n1027;
  assign n1250 = pi94 & n1098;
  assign n1251 = ~n1249 & ~n1250;
  assign n1252 = pi138 & ~n1251;
  assign n1253 = ~pi78 & ~pi136;
  assign n1254 = ~pi33 & pi136;
  assign n1255 = pi137 & ~n1254;
  assign n1256 = ~n1253 & n1255;
  assign n1257 = pi74 & ~pi136;
  assign n1258 = pi63 & pi136;
  assign n1259 = ~pi137 & ~n1258;
  assign n1260 = ~n1257 & n1259;
  assign n1261 = ~n1256 & ~n1260;
  assign n1262 = ~pi138 & ~n1261;
  assign po118 = n1252 | n1262;
  assign n1264 = pi99 & n1027;
  assign n1265 = ~pi112 & n1098;
  assign n1266 = ~n1264 & ~n1265;
  assign n1267 = pi138 & ~n1266;
  assign n1268 = pi73 & ~pi136;
  assign n1269 = pi68 & pi136;
  assign n1270 = ~pi137 & ~n1269;
  assign n1271 = ~n1268 & n1270;
  assign n1272 = ~pi84 & ~pi136;
  assign n1273 = ~pi32 & pi136;
  assign n1274 = pi137 & ~n1273;
  assign n1275 = ~n1272 & n1274;
  assign n1276 = ~n1271 & ~n1275;
  assign n1277 = ~pi138 & ~n1276;
  assign po119 = n1267 | n1277;
  assign n1279 = ~pi92 & pi138;
  assign n1280 = pi70 & ~pi138;
  assign n1281 = pi136 & ~n1280;
  assign n1282 = ~n1279 & n1281;
  assign n1283 = ~pi125 & pi138;
  assign n1284 = pi75 & ~pi138;
  assign n1285 = ~pi136 & ~n1284;
  assign n1286 = ~n1283 & n1285;
  assign n1287 = ~n1282 & ~n1286;
  assign n1288 = ~pi137 & ~n1287;
  assign n1289 = pi35 & n1130;
  assign n1290 = ~pi80 & ~pi138;
  assign n1291 = ~pi100 & pi138;
  assign n1292 = ~pi136 & ~n1291;
  assign n1293 = ~n1290 & n1292;
  assign n1294 = ~n1289 & ~n1293;
  assign n1295 = pi137 & ~n1294;
  assign po120 = n1288 | n1295;
  assign n1297 = n602 & n1145;
  assign n1298 = ~pi85 & ~n1297;
  assign n1299 = n339 & ~n593;
  assign po121 = ~n1298 & n1299;
  assign n1301 = ~pi98 & pi138;
  assign n1302 = pi71 & ~pi138;
  assign n1303 = pi136 & ~n1302;
  assign n1304 = ~n1301 & n1303;
  assign n1305 = ~pi23 & pi138;
  assign n1306 = pi76 & ~pi138;
  assign n1307 = ~pi136 & ~n1306;
  assign n1308 = ~n1305 & n1307;
  assign n1309 = ~n1304 & ~n1308;
  assign n1310 = ~pi137 & ~n1309;
  assign n1311 = pi36 & n1130;
  assign n1312 = ~pi81 & ~pi138;
  assign n1313 = ~pi97 & pi138;
  assign n1314 = ~pi136 & ~n1313;
  assign n1315 = ~n1312 & n1314;
  assign n1316 = ~n1311 & ~n1315;
  assign n1317 = pi137 & ~n1316;
  assign po122 = n1310 | n1317;
  assign n1319 = ~pi88 & pi138;
  assign n1320 = pi64 & ~pi138;
  assign n1321 = pi136 & ~n1320;
  assign n1322 = ~n1319 & n1321;
  assign n1323 = ~pi120 & pi138;
  assign n1324 = pi67 & ~pi138;
  assign n1325 = ~pi136 & ~n1324;
  assign n1326 = ~n1323 & n1325;
  assign n1327 = ~n1322 & ~n1326;
  assign n1328 = ~pi137 & ~n1327;
  assign n1329 = pi30 & n1130;
  assign n1330 = ~pi86 & ~pi138;
  assign n1331 = ~pi111 & pi138;
  assign n1332 = ~pi136 & ~n1331;
  assign n1333 = ~n1330 & n1332;
  assign n1334 = ~n1329 & ~n1333;
  assign n1335 = pi137 & ~n1334;
  assign po123 = n1328 | n1335;
  assign n1337 = pi116 & n339;
  assign n1338 = ~n662 & ~n668;
  assign po124 = n1337 & ~n1338;
  assign n1340 = ~pi97 & n629;
  assign n1341 = ~n688 & ~n1340;
  assign po125 = n1337 & ~n1341;
  assign n1343 = ~pi111 & ~n1183;
  assign n1344 = n1029 & ~n1343;
  assign n1345 = ~pi139 & n1183;
  assign n1346 = ~pi129 & ~n1345;
  assign po126 = n1344 & n1346;
  assign n1348 = pi112 & ~n1183;
  assign n1349 = ~pi141 & n1183;
  assign n1350 = n1029 & ~n1349;
  assign n1351 = ~pi129 & n1350;
  assign po127 = ~n1348 & n1351;
  assign n1353 = ~pi11 & pi54;
  assign n1354 = ~pi22 & n1353;
  assign n1355 = ~pi54 & pi113;
  assign n1356 = n339 & ~n1355;
  assign po128 = ~n1354 & n1356;
  assign n1358 = pi115 & ~n1183;
  assign n1359 = ~pi140 & n1183;
  assign n1360 = n1029 & ~n1359;
  assign n1361 = ~pi129 & n1360;
  assign po130 = ~n1358 & n1361;
  assign n1363 = pi54 & n339;
  assign n1364 = ~pi4 & n430;
  assign n1365 = ~pi9 & n1364;
  assign po131 = n1363 & ~n1365;
  assign po132 = ~pi122 | pi129;
  assign n1368 = ~pi54 & pi118;
  assign n1369 = ~n500 & ~n1368;
  assign po133 = ~pi129 & ~n1369;
  assign po134 = ~pi129 & ~n600;
  assign n1372 = ~pi120 & n1189;
  assign n1373 = ~pi111 & ~n1372;
  assign po135 = ~pi129 & n1373;
  assign n1375 = pi81 & pi120;
  assign po136 = ~pi129 & n1375;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi57 & ~pi129;
  assign n1380 = ~pi96 & pi125;
  assign n1381 = ~pi3 & ~n1380;
  assign po140 = ~pi129 & ~n1381;
  assign n1383 = ~pi126 & pi132;
  assign po141 = pi133 & n1383;
  assign po12 = 1'b1;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
endmodule
