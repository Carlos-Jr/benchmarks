module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 , pi30 , pi31 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 ;
  wire n65, n66, n67, n68, n69, n70, n71,
    n72, n73, n74, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87,
    n88, n89, n90, n91, n92, n93, n94, n95,
    n96, n97, n98, n99, n100, n101, n102,
    n103, n104, n105, n106, n107, n108, n109,
    n110, n111, n112, n113, n114, n115, n116,
    n117, n118, n119, n120, n121, n122, n123,
    n124, n125, n126, n127, n128, n129, n130,
    n131, n132, n133, n134, n135, n136, n137,
    n138, n139, n140, n141, n142, n143, n144,
    n145, n146, n147, n148, n149, n150, n151,
    n152, n153, n154, n155, n156, n157, n158,
    n159, n160, n161, n162, n163, n164, n165,
    n166, n167, n168, n169, n170, n171, n172,
    n173, n174, n175, n176, n177, n178, n179,
    n180, n181, n182, n183, n184, n185, n186,
    n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200,
    n201, n202, n203, n204, n205, n206, n207,
    n208, n209, n210, n211, n212, n213, n214,
    n215, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225, n226, n227, n228,
    n229, n230, n231, n232, n233, n234, n235,
    n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249,
    n250, n251, n252, n253, n254, n255, n256,
    n257, n258, n259, n260, n261, n262, n263,
    n264, n265, n266, n267, n268, n269, n270,
    n271, n272, n273, n274, n275, n276, n277,
    n278, n279, n280, n281, n282, n283, n284,
    n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298,
    n299, n300, n301, n302, n303, n304, n305,
    n306, n307, n308, n309, n310, n311, n312,
    n313, n314, n315, n316, n317, n318, n319,
    n320, n321, n322, n323, n324, n325, n326,
    n327, n328, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n485, n486, n487,
    n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501,
    n502, n503, n504, n505, n506, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n540, n541, n542, n543,
    n544, n545, n546, n547, n548, n549, n550,
    n551, n552, n553, n554, n555, n556, n557,
    n558, n559, n560, n561, n562, n563, n564,
    n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578,
    n579, n580, n581, n582, n583, n584, n585,
    n586, n587, n588, n589, n590, n591, n592,
    n593, n594, n595, n596, n597, n598, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n607, n608, n609, n610, n611, n612, n613,
    n614, n615, n616, n617, n618, n619, n620,
    n621, n622, n623, n624, n625, n626, n627,
    n628, n629, n630, n631, n632, n633, n634,
    n635, n636, n637, n638, n639, n640, n641,
    n642, n643, n644, n645, n646, n647, n648,
    n649, n650, n651, n652, n653, n654, n655,
    n656, n657, n658, n659, n660, n661, n662,
    n663, n664, n665, n666, n667, n668, n669,
    n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683,
    n684, n685, n686, n687, n688, n689, n690,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n718,
    n719, n720, n721, n722, n723, n724, n725,
    n726, n727, n728, n729, n730, n731, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767,
    n768, n769, n770, n771, n772, n773, n774,
    n775, n776, n777, n778, n779, n780, n781,
    n782, n783, n784, n785, n786, n787, n788,
    n789, n790, n791, n792, n793, n794, n795,
    n796, n797, n798, n799, n800, n801, n802,
    n803, n804, n805, n806, n807, n808, n809,
    n810, n811, n812, n813, n814, n815, n816,
    n817, n818, n819, n820, n821, n822, n823,
    n824, n825, n826, n827, n828, n829, n830,
    n831, n832, n833, n834, n835, n836, n837,
    n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851,
    n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865,
    n866, n867, n868, n869, n870, n871, n872,
    n873, n874, n875, n876, n877, n878, n879,
    n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893,
    n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n908, n909, n910, n911, n912, n913, n914,
    n915, n916, n917, n918, n919, n920, n921,
    n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n946, n947, n948, n949,
    n950, n951, n952, n953, n954, n955, n956,
    n957, n958, n959, n960, n961, n962, n963,
    n964, n965, n966, n967, n968, n969, n970,
    n971, n972, n973, n974, n975, n976, n977,
    n978, n979, n980, n981, n982, n983, n984,
    n985, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998,
    n999, n1000, n1001, n1002, n1003, n1004,
    n1005, n1006, n1007, n1008, n1009, n1010,
    n1011, n1012, n1013, n1014, n1015, n1016,
    n1017, n1018, n1019, n1020, n1021, n1022,
    n1023, n1024, n1025, n1026, n1027, n1028,
    n1029, n1030, n1031, n1032, n1033, n1034,
    n1035, n1036, n1037, n1038, n1039, n1040,
    n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052,
    n1053, n1054, n1055, n1056, n1057, n1058,
    n1059, n1060, n1061, n1062, n1063, n1064,
    n1065, n1066, n1067, n1068, n1069, n1070,
    n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082,
    n1083, n1084, n1085, n1086, n1087, n1088,
    n1089, n1090, n1091, n1092, n1093, n1094,
    n1095, n1096, n1097, n1098, n1099, n1100,
    n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1115, n1116, n1117, n1118,
    n1119, n1120, n1121, n1122, n1123, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130,
    n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142,
    n1143, n1144, n1145, n1146, n1147, n1148,
    n1149, n1150, n1151, n1152, n1153, n1154,
    n1155, n1156, n1157, n1158, n1159, n1160,
    n1161, n1162, n1163, n1164, n1165, n1166,
    n1167, n1168, n1169, n1170, n1171, n1172,
    n1173, n1174, n1175, n1176, n1177, n1178,
    n1179, n1180, n1181, n1182, n1183, n1184,
    n1185, n1186, n1187, n1188, n1189, n1190,
    n1191, n1192, n1193, n1194, n1195, n1196,
    n1197, n1198, n1199, n1200, n1201, n1202,
    n1203, n1204, n1205, n1206, n1207, n1208,
    n1209, n1210, n1211, n1212, n1213, n1214,
    n1215, n1216, n1217, n1218, n1219, n1220,
    n1221, n1222, n1223, n1224, n1225, n1226,
    n1227, n1228, n1229, n1230, n1231, n1232,
    n1233, n1234, n1235, n1236, n1237, n1238,
    n1239, n1240, n1241, n1242, n1243, n1244,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1262,
    n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274,
    n1275, n1276, n1277, n1278, n1279, n1280,
    n1281, n1282, n1283, n1284, n1285, n1286,
    n1287, n1288, n1289, n1290, n1291, n1292,
    n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304,
    n1305, n1306, n1307, n1308, n1309, n1310,
    n1311, n1312, n1313, n1314, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328,
    n1329, n1330, n1331, n1332, n1333, n1334,
    n1335, n1336, n1337, n1338, n1339, n1340,
    n1341, n1342, n1343, n1344, n1345, n1346,
    n1347, n1348, n1349, n1350, n1351, n1352,
    n1353, n1354, n1355, n1356, n1357, n1358,
    n1359, n1360, n1361, n1362, n1363, n1364,
    n1365, n1366, n1367, n1368, n1369, n1370,
    n1371, n1372, n1373, n1374, n1375, n1376,
    n1377, n1378, n1379, n1380, n1381, n1382,
    n1383, n1384, n1385, n1386, n1387, n1388,
    n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400,
    n1401, n1402, n1403, n1404, n1405, n1406,
    n1407, n1408, n1409, n1410, n1411, n1412,
    n1413, n1414, n1415, n1416, n1417, n1418,
    n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436,
    n1437, n1438, n1439, n1440, n1441, n1442,
    n1443, n1444, n1445, n1446, n1447, n1448,
    n1449, n1450, n1451, n1452, n1453, n1454,
    n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466,
    n1467, n1468, n1469, n1470, n1471, n1472,
    n1473, n1474, n1475, n1476, n1477, n1478,
    n1479, n1480, n1481, n1482, n1483, n1484,
    n1485, n1486, n1487, n1488, n1489, n1490,
    n1491, n1492, n1493, n1494, n1495, n1496,
    n1497, n1498, n1499, n1500, n1501, n1502,
    n1503, n1504, n1505, n1506, n1507, n1508,
    n1509, n1510, n1511, n1512, n1513, n1514,
    n1515, n1516, n1517, n1518, n1519, n1520,
    n1521, n1522, n1523, n1524, n1525, n1526,
    n1527, n1528, n1529, n1530, n1531, n1532,
    n1533, n1534, n1535, n1536, n1537, n1538,
    n1539, n1540, n1541, n1542, n1543, n1544,
    n1545, n1546, n1547, n1548, n1549, n1550,
    n1551, n1552, n1553, n1554, n1555, n1556,
    n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568,
    n1569, n1570, n1571, n1572, n1573, n1574,
    n1575, n1576, n1577, n1578, n1579, n1580,
    n1581, n1582, n1583, n1584, n1585, n1586,
    n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598,
    n1599, n1600, n1601, n1602, n1603, n1604,
    n1605, n1606, n1607, n1608, n1609, n1610,
    n1611, n1612, n1613, n1614, n1615, n1616,
    n1617, n1618, n1619, n1620, n1621, n1622,
    n1623, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634,
    n1635, n1636, n1637, n1638, n1639, n1640,
    n1641, n1642, n1643, n1644, n1645, n1646,
    n1647, n1648, n1649, n1650, n1651, n1652,
    n1653, n1654, n1655, n1656, n1657, n1658,
    n1659, n1660, n1661, n1662, n1663, n1664,
    n1665, n1666, n1667, n1668, n1669, n1670,
    n1671, n1672, n1673, n1674, n1675, n1676,
    n1677, n1678, n1679, n1680, n1681, n1682,
    n1683, n1684, n1685, n1686, n1687, n1688,
    n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700,
    n1701, n1702, n1703, n1704, n1705, n1706,
    n1707, n1708, n1709, n1710, n1711, n1712,
    n1713, n1714, n1715, n1716, n1717, n1718,
    n1719, n1720, n1721, n1722, n1723, n1724,
    n1725, n1726, n1727, n1728, n1729, n1730,
    n1731, n1732, n1733, n1734, n1735, n1736,
    n1737, n1738, n1739, n1740, n1741, n1742,
    n1743, n1744, n1745, n1746, n1747, n1748,
    n1749, n1750, n1751, n1752, n1753, n1754,
    n1755, n1756, n1757, n1758, n1759, n1760,
    n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772,
    n1773, n1774, n1775, n1776, n1777, n1778,
    n1779, n1780, n1781, n1782, n1783, n1784,
    n1785, n1786, n1787, n1788, n1789, n1790,
    n1791, n1792, n1793, n1794, n1795, n1796,
    n1797, n1798, n1799, n1800, n1801, n1802,
    n1803, n1804, n1805, n1806, n1807, n1808,
    n1809, n1810, n1811, n1812, n1813, n1814,
    n1815, n1816, n1817, n1818, n1819, n1820,
    n1821, n1822, n1823, n1824, n1825, n1826,
    n1827, n1828, n1829, n1830, n1831, n1832,
    n1833, n1834, n1835, n1836, n1837, n1838,
    n1839, n1840, n1841, n1842, n1843, n1844,
    n1845, n1846, n1847, n1848, n1849, n1850,
    n1851, n1852, n1853, n1854, n1855, n1856,
    n1857, n1858, n1859, n1860, n1861, n1862,
    n1863, n1864, n1865, n1866, n1867, n1868,
    n1869, n1870, n1871, n1872, n1873, n1874,
    n1875, n1876, n1877, n1878, n1879, n1880,
    n1881, n1882, n1883, n1884, n1885, n1886,
    n1887, n1888, n1889, n1890, n1891, n1892,
    n1893, n1894, n1895, n1896, n1897, n1898,
    n1899, n1900, n1901, n1902, n1903, n1904,
    n1905, n1906, n1907, n1908, n1909, n1910,
    n1911, n1912, n1913, n1914, n1915, n1916,
    n1917, n1918, n1919, n1920, n1921, n1922,
    n1923, n1924, n1925, n1926, n1927, n1928,
    n1929, n1930, n1931, n1932, n1933, n1934,
    n1935, n1936, n1937, n1938, n1939, n1940,
    n1941, n1942, n1943, n1944, n1945, n1946,
    n1947, n1948, n1949, n1950, n1951, n1952,
    n1953, n1954, n1955, n1956, n1957, n1958,
    n1959, n1960, n1961, n1962, n1963, n1964,
    n1965, n1966, n1967, n1968, n1969, n1970,
    n1971, n1972, n1973, n1974, n1975, n1976,
    n1977, n1978, n1979, n1980, n1981, n1982,
    n1983, n1984, n1985, n1986, n1987, n1988,
    n1989, n1990, n1991, n1992, n1993, n1994,
    n1995, n1996, n1997, n1998, n1999, n2000,
    n2001, n2002, n2003, n2004, n2005, n2006,
    n2007, n2008, n2009, n2010, n2011, n2012,
    n2013, n2014, n2015, n2016, n2017, n2018,
    n2019, n2020, n2021, n2022, n2023, n2024,
    n2025, n2026, n2027, n2028, n2029, n2030,
    n2031, n2032, n2033, n2034, n2035, n2036,
    n2037, n2038, n2039, n2040, n2041, n2042,
    n2043, n2044, n2045, n2046, n2047, n2048,
    n2049, n2050, n2051, n2052, n2053, n2054,
    n2055, n2056, n2057, n2058, n2059, n2060,
    n2061, n2062, n2063, n2064, n2065, n2066,
    n2067, n2068, n2069, n2070, n2071, n2072,
    n2073, n2074, n2075, n2076, n2077, n2078,
    n2079, n2080, n2081, n2082, n2083, n2084,
    n2085, n2086, n2087, n2088, n2089, n2090,
    n2091, n2092, n2093, n2094, n2095, n2096,
    n2097, n2098, n2099, n2100, n2101, n2102,
    n2103, n2104, n2105, n2106, n2107, n2108,
    n2109, n2110, n2111, n2112, n2113, n2114,
    n2115, n2116, n2117, n2118, n2119, n2120,
    n2121, n2122, n2123, n2124, n2125, n2126,
    n2127, n2128, n2129, n2130, n2131, n2132,
    n2133, n2134, n2135, n2136, n2137, n2138,
    n2139, n2140, n2141, n2142, n2143, n2144,
    n2145, n2146, n2147, n2148, n2149, n2150,
    n2151, n2152, n2153, n2154, n2155, n2156,
    n2157, n2158, n2159, n2160, n2161, n2162,
    n2163, n2164, n2165, n2166, n2167, n2168,
    n2169, n2170, n2171, n2172, n2173, n2174,
    n2175, n2176, n2177, n2178, n2179, n2180,
    n2181, n2182, n2183, n2184, n2185, n2186,
    n2187, n2188, n2189, n2190, n2191, n2192,
    n2193, n2194, n2195, n2196, n2197, n2198,
    n2199, n2200, n2201, n2202, n2203, n2204,
    n2205, n2206, n2207, n2208, n2209, n2210,
    n2211, n2212, n2213, n2214, n2215, n2216,
    n2217, n2218, n2219, n2220, n2221, n2222,
    n2223, n2224, n2225, n2226, n2227, n2228,
    n2229, n2230, n2231, n2232, n2233, n2234,
    n2235, n2236, n2237, n2238, n2239, n2240,
    n2241, n2242, n2243, n2244, n2245, n2246,
    n2247, n2248, n2249, n2250, n2251, n2252,
    n2253, n2254, n2255, n2256, n2257, n2258,
    n2259, n2260, n2261, n2262, n2263, n2264,
    n2265, n2266, n2267, n2268, n2269, n2270,
    n2271, n2272, n2273, n2274, n2275, n2276,
    n2277, n2278, n2279, n2280, n2281, n2282,
    n2283, n2284, n2285, n2286, n2287, n2288,
    n2289, n2290, n2291, n2292, n2293, n2294,
    n2295, n2296, n2297, n2298, n2299, n2300,
    n2301, n2302, n2303, n2304, n2305, n2306,
    n2307, n2308, n2309, n2310, n2311, n2312,
    n2313, n2314, n2315, n2316, n2317, n2318,
    n2319, n2320, n2321, n2322, n2323, n2324,
    n2325, n2326, n2327, n2328, n2329, n2330,
    n2331, n2332, n2333, n2334, n2335, n2336,
    n2337, n2338, n2339, n2340, n2341, n2342,
    n2343, n2344, n2345, n2346, n2347, n2348,
    n2349, n2350, n2351, n2352, n2353, n2354,
    n2355, n2356, n2357, n2358, n2359, n2360,
    n2361, n2362, n2363, n2364, n2365, n2366,
    n2367, n2368, n2369, n2370, n2371, n2372,
    n2373, n2374, n2375, n2376, n2377, n2378,
    n2379, n2380, n2381, n2382, n2383, n2384,
    n2385, n2386, n2387, n2388, n2389, n2390,
    n2391, n2392, n2393, n2394, n2395, n2396,
    n2397, n2398, n2399, n2400, n2401, n2402,
    n2403, n2404, n2405, n2406, n2407, n2408,
    n2409, n2410, n2411, n2412, n2413, n2414,
    n2415, n2416, n2417, n2418, n2419, n2420,
    n2421, n2422, n2423, n2424, n2425, n2426,
    n2427, n2428, n2429, n2430, n2431, n2432,
    n2433, n2434, n2435, n2436, n2437, n2438,
    n2439, n2440, n2441, n2442, n2443, n2444,
    n2445, n2446, n2447, n2448, n2449, n2450,
    n2451, n2452, n2453, n2454, n2455, n2456,
    n2457, n2458, n2459, n2460, n2461, n2462,
    n2463, n2464, n2465, n2466, n2467, n2468,
    n2469, n2470, n2471, n2472, n2473, n2474,
    n2475, n2476, n2477, n2478, n2479, n2480,
    n2481, n2482, n2483, n2484, n2485, n2486,
    n2487, n2488, n2489, n2490, n2491, n2492,
    n2493, n2494, n2495, n2496, n2497, n2498,
    n2499, n2500, n2501, n2502, n2503, n2504,
    n2505, n2506, n2507, n2508, n2509, n2510,
    n2511, n2512, n2513, n2514, n2515, n2516,
    n2517, n2518, n2519, n2520, n2521, n2522,
    n2523, n2524, n2525, n2526, n2527, n2528,
    n2529, n2530, n2531, n2532, n2533, n2534,
    n2535, n2536, n2537, n2538, n2539, n2540,
    n2541, n2542, n2543, n2544, n2545, n2546,
    n2547, n2548, n2549, n2550, n2551, n2552,
    n2553, n2554, n2555, n2556, n2557, n2558,
    n2559, n2560, n2561, n2562, n2563, n2564,
    n2565, n2566, n2567, n2568, n2569, n2570,
    n2571, n2572, n2573, n2574, n2575, n2576,
    n2577, n2578, n2579, n2580, n2581, n2582,
    n2583, n2584, n2585, n2586, n2587, n2588,
    n2589, n2590, n2591, n2592, n2593, n2594,
    n2595, n2596, n2597, n2598, n2599, n2600,
    n2601, n2602, n2603, n2604, n2605, n2606,
    n2607, n2608, n2609, n2610, n2611, n2612,
    n2613, n2614, n2615, n2616, n2617, n2618,
    n2619, n2620, n2621, n2622, n2623, n2624,
    n2625, n2626, n2627, n2628, n2629, n2630,
    n2631, n2632, n2633, n2634, n2635, n2636,
    n2637, n2638, n2639, n2640, n2641, n2642,
    n2643, n2644, n2645, n2646, n2647, n2648,
    n2649, n2650, n2651, n2652, n2653, n2654,
    n2655, n2656, n2657, n2658, n2659, n2660,
    n2661, n2662, n2663, n2664, n2665, n2666,
    n2667, n2668, n2669, n2670, n2671, n2672,
    n2673, n2674, n2675, n2676, n2677, n2678,
    n2679, n2680, n2681, n2682, n2683, n2684,
    n2685, n2686, n2687, n2688, n2689, n2690,
    n2691, n2692, n2693, n2694, n2695, n2696,
    n2697, n2698, n2699, n2700, n2701, n2702,
    n2703, n2704, n2705, n2706, n2707, n2708,
    n2709, n2710, n2711, n2712, n2713, n2714,
    n2715, n2716, n2717, n2718, n2719, n2720,
    n2721, n2722, n2723, n2724, n2725, n2726,
    n2727, n2728, n2729, n2730, n2731, n2732,
    n2733, n2734, n2735, n2736, n2737, n2738,
    n2739, n2740, n2741, n2742, n2743, n2744,
    n2745, n2746, n2747, n2748, n2749, n2750,
    n2751, n2752, n2753, n2754, n2755, n2756,
    n2757, n2758, n2759, n2760, n2761, n2762,
    n2763, n2764, n2765, n2766, n2767, n2768,
    n2769, n2770, n2771, n2772, n2773, n2774,
    n2775, n2776, n2777, n2778, n2779, n2780,
    n2781, n2782, n2783, n2784, n2785, n2786,
    n2787, n2788, n2789, n2790, n2791, n2792,
    n2793, n2794, n2795, n2796, n2797, n2798,
    n2799, n2800, n2801, n2802, n2803, n2804,
    n2805, n2806, n2807, n2808, n2809, n2810,
    n2811, n2812, n2813, n2814, n2815, n2816,
    n2817, n2818, n2819, n2820, n2821, n2822,
    n2823, n2824, n2825, n2826, n2827, n2828,
    n2829, n2830, n2831, n2832, n2833, n2834,
    n2835, n2836, n2837, n2838, n2839, n2840,
    n2841, n2842, n2843, n2844, n2845, n2846,
    n2847, n2848, n2849, n2850, n2851, n2852,
    n2853, n2854, n2855, n2856, n2857, n2858,
    n2859, n2860, n2861, n2862, n2863, n2864,
    n2865, n2866, n2867, n2868, n2869, n2870,
    n2871, n2872, n2873, n2874, n2875, n2876,
    n2877, n2878, n2879, n2880, n2881, n2882,
    n2883, n2884, n2885, n2886, n2887, n2888,
    n2889, n2890, n2891, n2892, n2893, n2894,
    n2895, n2896, n2897, n2898, n2899, n2900,
    n2901, n2902, n2903, n2904, n2905, n2906,
    n2907, n2908, n2909, n2910, n2911, n2912,
    n2913, n2914, n2915, n2916, n2917, n2918,
    n2919, n2920, n2921, n2922, n2923, n2924,
    n2925, n2926, n2927, n2928, n2929, n2930,
    n2931, n2932, n2933, n2934, n2935, n2936,
    n2937, n2938, n2939, n2940, n2941, n2942,
    n2943, n2944, n2945, n2946, n2947, n2948,
    n2949, n2950, n2951, n2952, n2953, n2954,
    n2955, n2956, n2957, n2958, n2959, n2960,
    n2961, n2962, n2963, n2964, n2965, n2966,
    n2967, n2968, n2969, n2970, n2971, n2972,
    n2973, n2974, n2975, n2976, n2977, n2978,
    n2979, n2980, n2981, n2982, n2983, n2984,
    n2985, n2986, n2987, n2988, n2989, n2990,
    n2991, n2992, n2993, n2994, n2995, n2996,
    n2997, n2998, n2999, n3000, n3001, n3002,
    n3003, n3004, n3005, n3006, n3007, n3008,
    n3009, n3010, n3011, n3012, n3013, n3014,
    n3015, n3016, n3017, n3018, n3019, n3020,
    n3021, n3022, n3023, n3024, n3025, n3026,
    n3027, n3028, n3029, n3030, n3031, n3032,
    n3033, n3034, n3035, n3036, n3037, n3038,
    n3039, n3040, n3041, n3042, n3043, n3044,
    n3045, n3046, n3047, n3048, n3049, n3050,
    n3051, n3052, n3053, n3054, n3055, n3056,
    n3057, n3058, n3059, n3060, n3061, n3062,
    n3063, n3064, n3065, n3066, n3067, n3068,
    n3069, n3070, n3071, n3072, n3073, n3074,
    n3075, n3076, n3077, n3078, n3079, n3080,
    n3081, n3082, n3083, n3084, n3085, n3086,
    n3087, n3088, n3089, n3090, n3091, n3092,
    n3093, n3094, n3095, n3096, n3097, n3098,
    n3099, n3100, n3101, n3102, n3103, n3104,
    n3105, n3106, n3107, n3108, n3109, n3110,
    n3111, n3112, n3113, n3114, n3115, n3116,
    n3117, n3118, n3119, n3120, n3121, n3122,
    n3123, n3124, n3125, n3126, n3127, n3128,
    n3129, n3130, n3131, n3132, n3133, n3134,
    n3135, n3136, n3137, n3138, n3139, n3140,
    n3141, n3142, n3143, n3144, n3145, n3146,
    n3147, n3148, n3149, n3150, n3151, n3152,
    n3153, n3154, n3155, n3156, n3157, n3158,
    n3159, n3160, n3161, n3162, n3163, n3164,
    n3165, n3166, n3167, n3168, n3169, n3170,
    n3171, n3172, n3173, n3174, n3175, n3176,
    n3177, n3178, n3179, n3180, n3181, n3182,
    n3183, n3184, n3185, n3186, n3187, n3188,
    n3189, n3190, n3191, n3192, n3193, n3194,
    n3195, n3196, n3197, n3198, n3199, n3200,
    n3201, n3202, n3203, n3204, n3205, n3206,
    n3207, n3208, n3209, n3210, n3211, n3212,
    n3213, n3214, n3215, n3216, n3217, n3218,
    n3219, n3220, n3221, n3222, n3223, n3224,
    n3225, n3226, n3227, n3228, n3229, n3230,
    n3231, n3232, n3233, n3234, n3235, n3236,
    n3237, n3238, n3239, n3240, n3241, n3242,
    n3243, n3244, n3245, n3246, n3247, n3248,
    n3249, n3250, n3251, n3252, n3253, n3254,
    n3255, n3256, n3257, n3258, n3259, n3260,
    n3261, n3262, n3263, n3264, n3265, n3266,
    n3267, n3268, n3269, n3270, n3271, n3272,
    n3273, n3274, n3275, n3276, n3277, n3278,
    n3279, n3280, n3281, n3282, n3283, n3284,
    n3285, n3286, n3287, n3288, n3289, n3290,
    n3291, n3292, n3293, n3294, n3295, n3296,
    n3297, n3298, n3299, n3300, n3301, n3302,
    n3303, n3304, n3305, n3306, n3307, n3308,
    n3309, n3310, n3311, n3312, n3313, n3314,
    n3315, n3316, n3317, n3318, n3319, n3320,
    n3321, n3322, n3323, n3324, n3325, n3326,
    n3327, n3328, n3329, n3330, n3331, n3332,
    n3333, n3334, n3335, n3336, n3337, n3338,
    n3339, n3340, n3341, n3342, n3343, n3344,
    n3345, n3346, n3347, n3348, n3349, n3350,
    n3351, n3352, n3353, n3354, n3355, n3356,
    n3357, n3358, n3359, n3360, n3361, n3362,
    n3363, n3364, n3365, n3366, n3367, n3368,
    n3369, n3370, n3371, n3372, n3373, n3374,
    n3375, n3376, n3377, n3378, n3379, n3380,
    n3381, n3382, n3383, n3384, n3385, n3386,
    n3387, n3388, n3389, n3390, n3391, n3392,
    n3393, n3394, n3395, n3396, n3397, n3398,
    n3399, n3400, n3401, n3402, n3403, n3404,
    n3405, n3406, n3407, n3408, n3409, n3410,
    n3411, n3412, n3413, n3414, n3415, n3416,
    n3417, n3418, n3419, n3420, n3421, n3422,
    n3423, n3424, n3425, n3426, n3427, n3428,
    n3429, n3430, n3431, n3432, n3433, n3434,
    n3435, n3436, n3437, n3438, n3439, n3440,
    n3441, n3442, n3443, n3444, n3445, n3446,
    n3447, n3448, n3449, n3450, n3451, n3452,
    n3453, n3454, n3455, n3456, n3457, n3458,
    n3459, n3460, n3461, n3462, n3463, n3464,
    n3465, n3466, n3467, n3468, n3469, n3470,
    n3471, n3472, n3473, n3474, n3475, n3476,
    n3477, n3478, n3479, n3480, n3481, n3482,
    n3483, n3484, n3485, n3486, n3487, n3488,
    n3489, n3490, n3491, n3492, n3493, n3494,
    n3495, n3496, n3497, n3498, n3499, n3500,
    n3501, n3502, n3503, n3504, n3505, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3678, n3679, n3680,
    n3681, n3682, n3683, n3684, n3685, n3686,
    n3687, n3688, n3689, n3690, n3691, n3692,
    n3693, n3694, n3695, n3696, n3697, n3698,
    n3699, n3700, n3701, n3702, n3703, n3704,
    n3705, n3706, n3707, n3708, n3709, n3710,
    n3711, n3712, n3713, n3714, n3715, n3716,
    n3717, n3718, n3719, n3720, n3721, n3722,
    n3723, n3724, n3725, n3726, n3727, n3728,
    n3729, n3730, n3731, n3732, n3733, n3734,
    n3735, n3736, n3737, n3738, n3739, n3740,
    n3741, n3742, n3743, n3744, n3745, n3746,
    n3747, n3748, n3749, n3750, n3751, n3752,
    n3753, n3754, n3755, n3756, n3757, n3758,
    n3759, n3760, n3761, n3762, n3763, n3764,
    n3765, n3766, n3767, n3768, n3769, n3770,
    n3771, n3772, n3773, n3774, n3775, n3776,
    n3777, n3778, n3779, n3780, n3781, n3782,
    n3783, n3784, n3785, n3786, n3787, n3788,
    n3789, n3790, n3791, n3792, n3793, n3794,
    n3795, n3796, n3797, n3798, n3799, n3800,
    n3801, n3802, n3803, n3804, n3805, n3806,
    n3807, n3808, n3809, n3810, n3811, n3812,
    n3813, n3814, n3815, n3816, n3817, n3818,
    n3819, n3820, n3821, n3822, n3823, n3824,
    n3825, n3826, n3827, n3828, n3829, n3830,
    n3831, n3832, n3833, n3834, n3835, n3836,
    n3837, n3838, n3839, n3840, n3841, n3842,
    n3843, n3844, n3845, n3846, n3847, n3848,
    n3849, n3850, n3851, n3852, n3853, n3854,
    n3855, n3856, n3857, n3858, n3859, n3860,
    n3861, n3862, n3863, n3864, n3865, n3866,
    n3867, n3868, n3869, n3870, n3871, n3872,
    n3873, n3874, n3875, n3876, n3877, n3878,
    n3879, n3880, n3881, n3882, n3883, n3884,
    n3885, n3886, n3887, n3888, n3889, n3890,
    n3891, n3892, n3893, n3894, n3895, n3896,
    n3897, n3898, n3899, n3900, n3901, n3902,
    n3903, n3904, n3905, n3906, n3907, n3908,
    n3909, n3910, n3911, n3912, n3913, n3914,
    n3915, n3916, n3917, n3918, n3919, n3920,
    n3921, n3922, n3923, n3924, n3925, n3926,
    n3927, n3928, n3929, n3930, n3931, n3932,
    n3933, n3934, n3935, n3936, n3937, n3938,
    n3939, n3940, n3941, n3942, n3943, n3944,
    n3945, n3946, n3947, n3948, n3949, n3950,
    n3951, n3952, n3953, n3954, n3955, n3956,
    n3957, n3958, n3959, n3960, n3961, n3962,
    n3963, n3964, n3965, n3966, n3967, n3968,
    n3969, n3970, n3971, n3972, n3973, n3974,
    n3975, n3976, n3977, n3978, n3979, n3980,
    n3981, n3982, n3983, n3984, n3985, n3986,
    n3987, n3988, n3989, n3990, n3991, n3992,
    n3993, n3994, n3995, n3996, n3997, n3998,
    n3999, n4000, n4001, n4002, n4003, n4004,
    n4005, n4006, n4007, n4008, n4009, n4010,
    n4011, n4012, n4013, n4014, n4015, n4016,
    n4017, n4018, n4019, n4020, n4021, n4022,
    n4023, n4024, n4025, n4026, n4027, n4028,
    n4029, n4030, n4031, n4032, n4033, n4034,
    n4035, n4036, n4037, n4038, n4039, n4040,
    n4041, n4042, n4043, n4044, n4045, n4046,
    n4047, n4048, n4049, n4050, n4051, n4052,
    n4053, n4054, n4055, n4056, n4057, n4058,
    n4059, n4060, n4061, n4062, n4063, n4064,
    n4065, n4066, n4067, n4068, n4069, n4070,
    n4071, n4072, n4073, n4074, n4075, n4076,
    n4077, n4078, n4079, n4080, n4081, n4082,
    n4083, n4084, n4085, n4086, n4087, n4088,
    n4089, n4090, n4091, n4092, n4093, n4094,
    n4095, n4096, n4097, n4098, n4099, n4100,
    n4101, n4102, n4103, n4104, n4105, n4106,
    n4107, n4108, n4109, n4110, n4111, n4112,
    n4113, n4114, n4115, n4116, n4117, n4118,
    n4119, n4120, n4121, n4122, n4123, n4124,
    n4125, n4126, n4127, n4128, n4129, n4130,
    n4131, n4132, n4133, n4134, n4135, n4136,
    n4137, n4138, n4139, n4140, n4141, n4142,
    n4143, n4144, n4145, n4146, n4147, n4148,
    n4149, n4150, n4151, n4152, n4153, n4154,
    n4155, n4156, n4157, n4158, n4159, n4160,
    n4161, n4162, n4163, n4164, n4165, n4166,
    n4167, n4168, n4169, n4170, n4171, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4276, n4277, n4278, n4279, n4280,
    n4281, n4282, n4283, n4284, n4285, n4286,
    n4287, n4288, n4289, n4290, n4291, n4292,
    n4293, n4294, n4295, n4296, n4297, n4298,
    n4299, n4300, n4301, n4302, n4303, n4304,
    n4305, n4306, n4307, n4308, n4309, n4310,
    n4311, n4312, n4313, n4314, n4315, n4316,
    n4317, n4318, n4319, n4320, n4321, n4322,
    n4323, n4324, n4325, n4326, n4327, n4328,
    n4329, n4330, n4331, n4332, n4333, n4334,
    n4335, n4336, n4337, n4338, n4339, n4340,
    n4341, n4342, n4343, n4344, n4345, n4346,
    n4347, n4348, n4349, n4350, n4351, n4352,
    n4353, n4354, n4355, n4356, n4357, n4358,
    n4359, n4360, n4361, n4362, n4363, n4364,
    n4365, n4366, n4367, n4368, n4369, n4370,
    n4371, n4372, n4373, n4374, n4375, n4376,
    n4377, n4378, n4379, n4380, n4381, n4382,
    n4383, n4384, n4385, n4386, n4387, n4388,
    n4389, n4390, n4391, n4392, n4393, n4394,
    n4395, n4396, n4397, n4398, n4399, n4400,
    n4401, n4402, n4403, n4404, n4405, n4406,
    n4407, n4408, n4409, n4410, n4411, n4412,
    n4413, n4414, n4415, n4416, n4417, n4418,
    n4419, n4420, n4421, n4422, n4423, n4424,
    n4425, n4426, n4427, n4428, n4429, n4430,
    n4431, n4432, n4433, n4434, n4435, n4436,
    n4437, n4438, n4439, n4440, n4441, n4442,
    n4443, n4444, n4445, n4446, n4447, n4448,
    n4449, n4450, n4451, n4452, n4453, n4454,
    n4455, n4456, n4457, n4458, n4459, n4460,
    n4461, n4462, n4463, n4464, n4465, n4466,
    n4467, n4468, n4469, n4470, n4471, n4472,
    n4473, n4474, n4475, n4476, n4477, n4478,
    n4479, n4480, n4481, n4482, n4483, n4484,
    n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496,
    n4497, n4498, n4499, n4500, n4501, n4502,
    n4503, n4504, n4505, n4506, n4507, n4508,
    n4509, n4510, n4511, n4512, n4513, n4514,
    n4515, n4516, n4517, n4518, n4519, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526,
    n4527, n4528, n4529, n4530, n4531, n4532,
    n4533, n4534, n4535, n4536, n4537, n4538,
    n4539, n4540, n4541, n4542, n4543, n4544,
    n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556,
    n4557, n4558, n4559, n4560, n4561, n4562,
    n4563, n4564, n4565, n4566, n4567, n4568,
    n4569, n4570, n4571, n4572, n4573, n4574,
    n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586,
    n4587, n4588, n4589, n4590, n4591, n4592,
    n4593, n4594, n4595, n4596, n4597, n4598,
    n4599, n4600, n4601, n4602, n4603, n4604,
    n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616,
    n4617, n4618, n4619, n4620, n4621, n4622,
    n4623, n4624, n4625, n4626, n4627, n4628,
    n4629, n4630, n4631, n4632, n4633, n4634,
    n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646,
    n4647, n4648, n4649, n4650, n4651, n4652,
    n4653, n4654, n4655, n4656, n4657, n4658,
    n4659, n4660, n4661, n4662, n4663, n4664,
    n4665, n4666, n4667, n4668, n4669, n4670,
    n4671, n4672, n4673, n4674, n4675, n4676,
    n4677, n4678, n4679, n4680, n4681, n4682,
    n4683, n4684, n4685, n4686, n4687, n4688,
    n4689, n4690, n4691, n4692, n4693, n4694,
    n4695, n4696, n4697, n4698, n4699, n4700,
    n4701, n4702, n4703, n4704, n4705, n4706,
    n4707, n4708, n4709, n4710, n4711, n4712,
    n4713, n4714, n4715, n4716, n4717, n4718,
    n4719, n4720, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4784,
    n4785, n4786, n4787, n4788, n4789, n4790,
    n4791, n4792, n4793, n4794, n4795, n4796,
    n4797, n4798, n4799, n4800, n4801, n4802,
    n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5023, n5024,
    n5025, n5026, n5027, n5028, n5029, n5030,
    n5031, n5032, n5033, n5034, n5035, n5036,
    n5037, n5038, n5039, n5040, n5041, n5042,
    n5043, n5044, n5045, n5046, n5047, n5048,
    n5049, n5050, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072,
    n5073, n5074, n5075, n5076, n5077, n5078,
    n5079, n5080, n5081, n5082, n5083, n5084,
    n5085, n5086, n5087, n5088, n5089, n5090,
    n5091, n5092, n5093, n5094, n5095, n5096,
    n5097, n5098, n5099, n5100, n5101, n5102,
    n5103, n5104, n5105, n5106, n5107, n5108,
    n5109, n5110, n5111, n5112, n5113, n5114,
    n5115, n5116, n5117, n5118, n5119, n5120,
    n5121, n5122, n5123, n5124, n5125, n5126,
    n5127, n5128, n5129, n5130, n5131, n5132,
    n5133, n5134, n5135, n5136, n5137, n5138,
    n5139, n5140, n5141, n5142, n5143, n5144,
    n5145, n5146, n5147, n5148, n5149, n5150,
    n5151, n5152, n5153, n5154, n5155, n5156,
    n5157, n5158, n5159, n5160, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5170, n5171, n5172, n5173, n5174,
    n5175, n5176, n5177, n5178, n5179, n5180,
    n5181, n5182, n5183, n5184, n5185, n5186,
    n5187, n5188, n5189, n5190, n5191, n5192,
    n5193, n5194, n5195, n5196, n5197, n5198,
    n5199, n5200, n5201, n5202, n5203, n5204,
    n5205, n5206, n5207, n5208, n5209, n5210,
    n5211, n5212, n5213, n5214, n5215, n5216,
    n5217, n5218, n5219, n5220, n5221, n5222,
    n5223, n5224, n5225, n5226, n5227, n5228,
    n5229, n5230, n5231, n5232, n5233, n5234,
    n5235, n5236, n5237, n5238, n5239, n5240,
    n5241, n5242, n5243, n5244, n5245, n5246,
    n5247, n5248, n5249, n5250, n5251, n5252,
    n5253, n5254, n5255, n5256, n5257, n5258,
    n5259, n5260, n5261, n5262, n5263, n5264,
    n5265, n5266, n5267, n5268, n5269, n5270,
    n5271, n5272, n5273, n5274, n5275, n5276,
    n5277, n5278, n5279, n5280, n5281, n5282,
    n5283, n5284, n5285, n5286, n5287, n5288,
    n5289, n5290, n5291, n5292, n5293, n5294,
    n5295, n5296, n5297, n5298, n5299, n5300,
    n5301, n5302, n5303, n5304, n5305, n5306,
    n5307, n5308, n5309, n5310, n5311, n5312,
    n5313, n5314, n5315, n5316, n5317, n5318,
    n5319, n5320, n5321, n5322, n5323, n5324,
    n5325, n5326, n5327, n5328, n5329, n5330,
    n5331, n5332, n5333, n5334, n5335, n5336,
    n5337, n5338, n5339, n5340, n5341, n5342,
    n5343, n5344, n5345, n5346, n5347, n5348,
    n5349, n5350, n5351, n5352, n5353, n5354,
    n5355, n5356, n5357, n5358, n5359, n5360,
    n5361, n5362, n5363, n5364, n5365, n5366,
    n5367, n5368, n5369, n5370, n5371, n5372,
    n5373, n5374, n5375, n5376, n5377, n5378,
    n5379, n5380, n5381, n5382, n5383, n5384,
    n5385, n5386, n5387, n5388, n5389, n5390,
    n5391, n5392, n5393, n5394, n5395, n5396,
    n5397, n5398, n5399, n5400, n5401, n5402,
    n5403, n5404, n5405, n5406, n5407, n5408,
    n5409, n5410, n5411, n5412, n5413, n5414,
    n5415, n5416, n5417, n5418, n5419, n5420,
    n5421, n5422, n5423, n5424, n5425, n5426,
    n5427, n5428, n5429, n5430, n5431, n5432,
    n5433, n5434, n5435, n5436, n5437, n5438,
    n5439, n5440, n5441, n5442, n5443, n5444,
    n5445, n5446, n5447, n5448, n5449, n5450,
    n5451, n5452, n5453, n5454, n5455, n5456,
    n5457, n5458, n5459, n5460, n5461, n5462,
    n5463, n5464, n5465, n5466, n5467, n5468,
    n5469, n5470, n5471, n5472, n5473, n5474,
    n5475, n5476, n5477, n5478, n5479, n5480,
    n5481, n5482, n5483, n5484, n5485, n5486,
    n5487, n5488, n5489, n5490, n5491, n5492,
    n5493, n5494, n5495, n5496, n5497, n5498,
    n5499, n5500, n5501, n5502, n5503, n5504,
    n5505, n5506, n5507, n5508, n5509, n5510,
    n5511, n5512, n5513, n5514, n5515, n5516,
    n5517, n5518, n5519, n5520, n5521, n5522,
    n5523, n5524, n5525, n5526, n5527, n5528,
    n5529, n5530, n5531, n5532, n5533, n5534,
    n5535, n5536, n5537, n5538, n5539, n5540,
    n5541, n5542, n5543, n5544, n5545, n5546,
    n5547, n5548, n5549, n5550, n5551, n5552,
    n5553, n5554, n5555, n5556, n5557, n5558,
    n5559, n5560, n5561, n5562, n5563, n5564,
    n5565, n5566, n5567, n5568, n5569, n5570,
    n5571, n5572, n5573, n5574, n5575, n5576,
    n5577, n5578, n5579, n5580, n5581, n5582,
    n5583, n5584, n5585, n5586, n5587, n5588,
    n5589, n5590, n5591, n5592, n5593, n5594,
    n5595, n5596, n5597, n5598, n5599, n5600,
    n5601, n5602, n5603, n5604, n5605, n5606,
    n5607, n5608, n5609, n5610, n5611, n5612,
    n5613, n5614, n5615, n5616, n5617, n5618,
    n5619, n5620, n5621, n5622, n5623, n5624,
    n5625, n5626, n5627, n5628, n5629, n5630,
    n5631, n5632, n5633, n5634, n5635, n5636,
    n5637, n5638, n5639, n5640, n5641, n5642,
    n5643, n5644, n5645, n5646, n5647, n5648,
    n5649, n5650, n5651, n5652, n5653, n5654,
    n5655, n5656, n5657, n5658, n5659, n5660,
    n5661, n5662, n5663, n5664, n5665, n5666,
    n5667, n5668, n5669, n5670, n5671, n5672,
    n5673, n5674, n5675, n5676, n5677, n5678,
    n5679, n5680, n5681, n5682, n5683, n5684,
    n5685, n5686, n5687, n5688, n5689, n5690,
    n5691, n5692, n5693, n5694, n5695, n5696,
    n5697, n5698, n5699, n5700, n5701, n5702,
    n5703, n5704, n5705, n5706, n5707, n5708,
    n5709, n5710, n5711, n5712, n5713, n5714,
    n5715, n5716, n5717, n5718, n5719, n5720,
    n5721, n5722, n5723, n5724, n5725, n5726,
    n5727, n5728, n5729, n5730, n5731, n5732,
    n5733, n5734, n5735, n5736, n5737, n5738,
    n5739, n5740, n5741, n5742, n5743, n5744,
    n5745, n5746, n5747, n5748, n5749, n5750,
    n5751, n5752, n5753, n5754, n5755, n5756,
    n5757, n5758, n5759, n5760, n5761, n5762,
    n5763, n5764, n5765, n5766, n5767, n5768,
    n5769, n5770, n5771, n5772, n5773, n5774,
    n5775, n5776, n5777, n5778, n5779, n5780,
    n5781, n5782, n5783, n5784, n5785, n5786,
    n5787, n5788, n5789, n5790, n5791, n5792,
    n5793, n5794, n5795, n5796, n5797, n5798,
    n5799, n5800, n5801, n5802, n5803, n5804,
    n5805, n5806, n5807, n5808, n5809, n5810,
    n5811, n5812, n5813, n5814, n5815, n5816,
    n5817, n5818, n5819, n5820, n5821, n5822,
    n5823, n5824, n5825, n5826, n5827, n5828,
    n5829, n5830, n5831, n5832, n5833, n5834,
    n5835, n5836, n5837, n5838, n5839, n5840,
    n5841, n5842, n5843, n5844, n5845, n5846,
    n5847, n5848, n5849, n5850, n5851, n5852,
    n5853, n5854, n5855, n5856, n5857, n5858,
    n5859, n5860, n5861, n5862, n5863, n5864,
    n5865, n5866, n5867, n5868, n5869, n5870,
    n5871, n5872, n5873, n5874, n5875, n5876,
    n5877, n5878, n5879, n5880, n5881, n5882,
    n5883, n5884, n5885, n5886, n5887, n5888,
    n5889, n5890, n5891, n5892, n5893, n5894,
    n5895, n5896, n5897, n5898, n5899, n5900,
    n5901, n5902, n5903, n5904, n5905, n5906,
    n5907, n5908, n5909, n5910, n5911, n5912,
    n5913, n5914, n5915, n5916, n5917, n5918,
    n5919, n5920, n5921, n5922, n5923, n5924,
    n5925, n5926, n5927, n5928, n5929, n5930,
    n5931, n5932, n5933, n5934, n5935, n5936,
    n5937, n5938, n5939, n5940, n5941, n5942,
    n5943, n5944, n5945, n5946, n5947, n5948,
    n5949, n5950, n5951, n5952, n5953, n5954,
    n5955, n5956, n5957, n5958, n5959, n5960,
    n5961, n5962, n5963, n5964, n5965, n5966,
    n5967, n5968, n5969, n5970, n5971, n5972,
    n5973, n5974, n5975, n5976, n5977, n5978,
    n5979, n5980, n5981, n5982, n5983, n5984,
    n5985, n5986, n5987, n5988, n5989, n5990,
    n5991, n5992, n5993, n5994, n5995, n5996,
    n5997, n5998, n5999, n6000, n6001, n6002,
    n6003, n6004, n6005, n6006, n6007, n6008,
    n6009, n6010, n6011, n6012, n6013, n6014,
    n6015, n6016, n6017, n6018, n6019, n6020,
    n6021, n6022, n6023, n6024, n6025, n6026,
    n6027, n6028, n6029, n6030, n6031, n6032,
    n6033, n6034, n6035, n6036, n6037, n6038,
    n6039, n6040, n6041, n6042, n6043, n6044,
    n6045, n6046, n6047, n6048, n6049, n6050,
    n6051, n6052, n6053, n6054, n6055, n6056,
    n6057, n6058, n6059, n6060, n6061, n6062,
    n6063, n6064, n6065, n6066, n6067, n6068,
    n6069, n6070, n6071, n6072, n6073, n6074,
    n6075, n6076, n6077, n6078, n6079, n6080,
    n6081, n6082, n6083, n6084, n6085, n6086,
    n6087, n6088, n6089, n6090, n6091, n6092,
    n6093, n6094, n6095, n6096, n6097, n6098,
    n6099, n6100, n6101, n6102, n6103, n6104,
    n6105, n6106, n6107, n6108, n6109, n6110,
    n6111, n6112, n6113, n6114, n6115, n6116,
    n6117, n6118, n6119, n6120, n6121, n6122,
    n6123, n6124, n6125, n6126, n6127, n6128,
    n6129, n6130, n6131, n6132, n6133, n6134,
    n6135, n6136, n6137, n6138, n6139, n6140,
    n6141, n6142, n6143, n6144, n6145, n6146,
    n6147, n6148, n6149, n6150, n6151, n6152,
    n6153, n6154, n6155, n6156, n6157, n6158,
    n6159, n6160, n6161, n6162, n6163, n6164,
    n6165, n6166, n6167, n6168, n6169, n6170,
    n6171, n6172, n6173, n6174, n6175, n6176,
    n6177, n6178, n6179, n6180, n6181, n6182,
    n6183, n6184, n6185, n6186, n6187, n6188,
    n6189, n6190, n6191, n6192, n6193, n6194,
    n6195, n6196, n6197, n6198, n6199, n6200,
    n6201, n6202, n6203, n6204, n6205, n6206,
    n6207, n6208, n6209, n6210, n6211, n6212,
    n6213, n6214, n6215, n6216, n6217, n6218,
    n6219, n6220, n6221, n6222, n6223, n6224,
    n6225, n6226, n6227, n6228, n6229, n6230,
    n6231, n6232, n6233, n6234, n6235, n6236,
    n6237, n6238, n6239, n6240, n6241, n6242,
    n6243, n6244, n6245, n6246, n6247, n6248,
    n6249, n6250, n6251, n6252, n6253, n6254,
    n6255, n6256, n6257, n6258, n6259, n6260,
    n6261, n6262, n6263, n6264, n6265, n6266,
    n6267, n6268, n6269, n6270, n6271, n6272,
    n6273, n6274, n6275, n6276, n6277, n6278,
    n6279, n6280, n6281, n6282, n6283, n6284,
    n6285, n6286, n6287, n6288, n6289, n6290,
    n6291, n6292, n6293, n6294, n6295, n6296,
    n6297, n6298, n6299, n6300, n6301, n6302,
    n6303, n6304, n6305, n6306, n6307, n6308,
    n6309, n6310, n6311, n6312, n6313, n6314,
    n6315, n6316, n6317, n6318, n6319, n6320,
    n6321, n6322, n6323, n6324, n6325, n6326,
    n6327, n6328, n6329, n6330, n6331, n6332,
    n6333, n6334, n6335, n6336, n6337, n6338,
    n6339, n6340, n6341, n6342, n6343, n6344,
    n6345, n6346, n6347, n6348, n6349, n6350,
    n6351, n6352, n6353, n6354, n6355, n6356,
    n6357, n6358, n6359, n6360, n6361, n6362,
    n6363, n6364, n6365, n6366, n6367, n6368,
    n6369, n6370, n6371, n6372, n6373, n6374,
    n6375, n6376, n6377, n6378, n6379, n6380,
    n6381, n6382, n6383, n6384, n6385, n6386,
    n6387, n6388, n6389, n6390, n6391, n6392,
    n6393, n6394, n6395, n6396, n6397, n6398,
    n6399, n6400, n6401, n6402, n6403, n6404,
    n6405, n6406, n6407, n6408, n6409, n6410,
    n6411, n6412, n6413, n6414, n6415, n6416,
    n6417, n6418, n6419, n6420, n6421, n6422,
    n6423, n6424, n6425, n6426, n6427, n6428,
    n6429, n6430, n6431, n6432, n6433, n6434,
    n6435, n6436, n6437, n6438, n6439, n6440,
    n6441, n6442, n6443, n6444, n6445, n6446,
    n6447, n6448, n6449, n6450, n6451, n6452,
    n6453, n6454, n6455, n6456, n6457, n6458,
    n6459, n6460, n6461, n6462, n6463, n6464,
    n6465, n6466, n6467, n6468, n6469, n6470,
    n6471, n6472, n6473, n6474, n6475, n6476,
    n6477, n6478, n6479, n6480, n6481, n6482,
    n6483, n6484, n6485, n6486, n6487, n6488,
    n6489, n6490, n6491, n6492, n6493, n6494,
    n6495, n6496, n6497, n6498, n6499, n6500,
    n6501, n6502, n6503, n6504, n6505, n6506,
    n6507, n6508, n6509, n6510, n6511, n6512,
    n6513, n6514, n6515, n6516, n6517, n6518,
    n6519, n6520, n6521, n6522, n6523, n6524,
    n6525, n6526, n6527, n6528, n6529, n6530,
    n6531, n6532, n6533, n6534, n6535, n6536,
    n6537, n6538, n6539, n6540, n6541, n6542,
    n6543, n6544, n6545, n6546, n6547, n6548,
    n6549, n6550, n6551, n6552, n6553, n6554,
    n6555, n6556, n6557, n6558, n6559, n6560,
    n6561, n6562, n6563, n6564, n6565, n6566,
    n6567, n6568, n6569, n6570, n6571, n6572,
    n6573, n6574, n6575, n6576, n6577, n6578,
    n6579, n6580, n6581, n6582, n6583, n6584,
    n6585, n6586, n6587, n6588, n6589, n6590,
    n6591, n6592, n6593, n6594, n6595, n6596,
    n6597, n6598, n6599, n6600, n6601, n6602,
    n6603, n6604, n6605, n6606, n6607, n6608,
    n6609, n6610, n6611, n6612, n6613, n6614,
    n6615, n6616, n6617, n6618, n6619, n6620,
    n6621, n6622, n6623, n6624, n6625, n6626,
    n6627, n6628, n6629, n6630, n6631, n6632,
    n6633, n6634, n6635, n6636, n6637, n6638,
    n6639, n6640, n6641, n6642, n6643, n6644,
    n6645, n6646, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6772, n6773, n6774, n6775, n6776,
    n6777, n6778, n6779, n6780, n6781, n6782,
    n6783, n6784, n6785, n6786, n6787, n6788,
    n6789, n6790, n6791, n6792, n6793, n6794,
    n6795, n6796, n6797, n6798, n6799, n6800,
    n6801, n6802, n6803, n6804, n6805, n6806,
    n6807, n6808, n6809, n6810, n6811, n6812,
    n6813, n6814, n6815, n6816, n6817, n6818,
    n6819, n6820, n6821, n6822, n6823, n6824,
    n6825, n6826, n6827, n6828, n6829, n6830,
    n6831, n6832, n6833, n6834, n6835, n6836,
    n6837, n6838, n6839, n6840, n6841, n6842,
    n6843, n6844, n6845, n6846, n6847, n6848,
    n6849, n6850, n6851, n6852, n6853, n6854,
    n6855, n6856, n6857, n6858, n6859, n6860,
    n6861, n6862, n6863, n6864, n6865, n6866,
    n6867, n6868, n6869, n6870, n6871, n6872,
    n6873, n6874, n6875, n6876, n6877, n6878,
    n6879, n6880, n6881, n6882, n6883, n6884,
    n6885, n6886, n6887, n6888, n6889, n6890,
    n6891, n6892, n6893, n6894, n6895, n6896,
    n6897, n6898, n6899, n6900, n6901, n6902,
    n6903, n6904, n6905, n6906, n6907, n6908,
    n6909, n6910, n6911, n6912, n6913, n6914,
    n6915, n6916, n6917, n6918, n6919, n6920,
    n6921, n6922, n6923, n6924, n6925, n6926,
    n6927, n6928, n6929, n6930, n6931, n6932,
    n6933, n6934, n6935, n6936, n6937, n6938,
    n6939, n6940, n6941, n6942, n6943, n6944,
    n6945, n6946, n6947, n6948, n6949, n6950,
    n6951, n6952, n6953, n6954, n6955, n6956,
    n6957, n6958, n6959, n6960, n6961, n6962,
    n6963, n6964, n6965, n6966, n6967, n6968,
    n6969, n6970, n6971, n6972, n6973, n6974,
    n6975, n6976, n6977, n6978, n6979, n6980,
    n6981, n6982, n6983, n6984, n6985, n6986,
    n6987, n6988, n6989, n6990, n6991, n6992,
    n6993, n6994, n6995, n6996, n6997, n6998,
    n6999, n7000, n7001, n7002, n7003, n7004,
    n7005, n7006, n7007, n7008, n7009, n7010,
    n7011, n7012, n7013, n7014, n7015, n7016,
    n7017, n7018, n7019, n7020, n7021, n7022,
    n7023, n7024, n7025, n7026, n7027, n7028,
    n7029, n7030, n7031, n7032, n7033, n7034,
    n7035, n7036, n7037, n7038, n7039, n7040,
    n7041, n7042, n7043, n7044, n7045, n7046,
    n7047, n7048, n7049, n7050, n7051, n7052,
    n7053, n7054, n7055, n7056, n7057, n7058,
    n7059, n7060, n7061, n7062, n7063, n7064,
    n7065, n7066, n7067, n7068, n7069, n7070,
    n7071, n7072, n7073, n7074, n7075, n7076,
    n7077, n7078, n7079, n7080, n7081, n7082,
    n7083, n7084, n7085, n7086, n7087, n7088,
    n7089, n7090, n7091, n7092, n7093, n7094,
    n7095, n7096, n7097, n7098, n7099, n7100,
    n7101, n7102, n7103, n7104, n7105, n7106,
    n7107, n7108, n7109, n7110, n7111, n7112,
    n7113, n7114, n7115, n7116, n7117, n7118,
    n7119, n7120, n7121, n7122, n7123, n7124,
    n7125, n7126, n7127, n7128, n7129, n7130,
    n7131, n7132, n7133, n7134, n7135, n7136,
    n7137, n7138, n7139, n7140, n7141, n7142,
    n7143, n7144, n7145, n7146, n7147, n7148,
    n7149, n7150, n7151, n7152, n7153, n7154,
    n7155, n7156, n7157, n7158, n7159, n7160,
    n7161, n7162, n7163, n7164, n7165, n7166,
    n7167, n7168, n7169, n7170, n7171, n7172,
    n7173, n7174, n7175, n7176, n7177, n7178,
    n7179, n7180, n7181, n7182, n7183, n7184,
    n7185, n7186, n7187, n7188, n7189, n7190,
    n7191, n7192, n7193, n7194, n7195, n7196,
    n7197, n7198, n7199, n7200, n7201, n7202,
    n7203, n7204, n7205, n7206, n7207, n7208,
    n7209, n7210, n7211, n7212, n7213, n7214,
    n7215, n7216, n7217, n7218, n7219, n7220,
    n7221, n7222, n7223, n7224, n7225, n7226,
    n7227, n7228, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7282, n7283, n7284, n7285, n7286,
    n7287, n7288, n7289, n7290, n7291, n7292,
    n7293, n7294, n7295, n7296, n7297, n7298,
    n7299, n7300, n7301, n7302, n7303, n7304,
    n7305, n7306, n7307, n7308, n7309, n7310,
    n7311, n7312, n7313, n7314, n7315, n7316,
    n7317, n7318, n7319, n7320, n7321, n7322,
    n7323, n7324, n7325, n7326, n7327, n7328,
    n7329, n7330, n7331, n7332, n7333, n7334,
    n7335, n7336, n7337, n7338, n7339, n7340,
    n7341, n7342, n7343, n7344, n7345, n7346,
    n7347, n7348, n7349, n7350, n7351, n7352,
    n7353, n7354, n7355, n7356, n7357, n7358,
    n7359, n7360, n7361, n7362, n7363, n7364,
    n7365, n7366, n7367, n7368, n7369, n7370,
    n7371, n7372, n7373, n7374, n7375, n7376,
    n7377, n7378, n7379, n7380, n7381, n7382,
    n7383, n7384, n7385, n7386, n7387, n7388,
    n7389, n7390, n7391, n7392, n7393, n7394,
    n7395, n7396, n7397, n7398, n7399, n7400,
    n7401, n7402, n7403, n7404, n7405, n7406,
    n7407, n7408, n7409, n7410, n7411, n7412,
    n7413, n7414, n7415, n7416, n7417, n7418,
    n7419, n7420, n7421, n7422, n7423, n7424,
    n7425, n7426, n7427, n7428, n7429, n7430,
    n7431, n7432, n7433, n7434, n7435, n7436,
    n7437, n7438, n7439, n7440, n7441, n7442,
    n7443, n7444, n7445, n7446, n7447, n7448,
    n7449, n7450, n7451, n7452, n7453, n7454,
    n7455, n7456, n7457, n7458, n7459, n7460,
    n7461, n7462, n7463, n7464, n7465, n7466,
    n7467, n7468, n7469, n7470, n7471, n7472,
    n7473, n7474, n7475, n7476, n7477, n7478,
    n7479, n7480, n7481, n7482, n7483, n7484,
    n7485, n7486, n7487, n7488, n7489, n7490,
    n7491, n7492, n7493, n7494, n7495, n7496,
    n7497, n7498, n7499, n7500, n7501, n7502,
    n7503, n7504, n7505, n7506, n7507, n7508,
    n7509, n7510, n7511, n7512, n7513, n7514,
    n7515, n7516, n7517, n7518, n7519, n7520,
    n7521, n7522, n7523, n7524, n7525, n7526,
    n7527, n7528, n7529, n7530, n7531, n7532,
    n7533, n7534, n7535, n7536, n7537, n7538,
    n7539, n7540, n7541, n7542, n7543, n7544,
    n7545, n7546, n7547, n7548, n7549, n7550,
    n7551, n7552, n7553, n7554, n7555, n7556,
    n7557, n7558, n7559, n7560, n7561, n7562,
    n7563, n7564, n7565, n7566, n7567, n7568,
    n7569, n7570, n7571, n7572, n7573, n7574,
    n7575, n7576, n7577, n7578, n7579, n7580,
    n7581, n7582, n7583, n7584, n7585, n7586,
    n7587, n7588, n7589, n7590, n7591, n7592,
    n7593, n7594, n7595, n7596, n7597, n7598,
    n7599, n7600, n7601, n7602, n7603, n7604,
    n7605, n7606, n7607, n7608, n7609, n7610,
    n7611, n7612, n7613, n7614, n7615, n7616,
    n7617, n7618, n7619, n7620, n7621, n7622,
    n7623, n7624, n7625, n7626, n7627, n7628,
    n7629, n7630, n7631, n7632, n7633, n7634,
    n7635, n7636, n7637, n7638, n7639, n7640,
    n7641, n7642, n7643, n7644, n7645, n7646,
    n7647, n7648, n7649, n7650, n7651, n7652,
    n7653, n7654, n7655, n7656, n7657, n7658,
    n7659, n7660, n7661, n7662, n7663, n7664,
    n7665, n7666, n7667, n7668, n7669, n7670,
    n7671, n7672, n7673, n7674, n7675, n7676,
    n7677, n7678, n7679, n7680, n7681, n7682,
    n7683, n7684, n7685, n7686, n7687, n7688,
    n7689, n7690, n7691, n7692, n7693, n7694,
    n7695, n7696, n7697, n7698, n7699, n7700,
    n7701, n7702, n7703, n7704, n7705, n7706,
    n7707, n7708, n7709, n7710, n7711, n7712,
    n7713, n7714, n7715, n7716, n7717, n7718,
    n7719, n7720, n7721, n7722, n7723, n7724,
    n7725, n7726, n7727, n7728, n7729, n7730,
    n7731, n7732, n7733, n7734, n7735, n7736,
    n7737, n7738, n7739, n7740, n7741, n7742,
    n7743, n7744, n7745, n7746, n7747, n7748,
    n7749, n7750, n7751, n7752, n7753, n7754,
    n7755, n7756, n7757, n7758, n7759, n7760,
    n7761, n7762, n7763, n7764, n7765, n7766,
    n7767, n7768, n7769, n7770, n7771, n7772,
    n7773, n7774, n7775, n7776, n7777, n7778,
    n7779, n7780, n7781, n7782, n7783, n7784,
    n7785, n7786, n7787, n7788, n7789, n7790,
    n7791, n7792, n7793, n7794, n7795, n7796,
    n7797, n7798, n7799, n7800, n7801, n7802,
    n7803, n7804, n7805, n7806, n7807, n7808,
    n7809, n7810, n7811, n7812, n7813, n7814,
    n7815, n7816, n7817, n7818, n7819, n7820,
    n7821, n7822, n7823, n7824, n7825, n7826,
    n7827, n7828, n7829, n7830, n7831, n7832,
    n7833, n7834, n7835, n7836, n7837, n7838,
    n7839, n7840, n7841, n7842, n7843, n7844,
    n7845, n7846, n7847, n7848, n7849, n7850,
    n7851, n7852, n7853, n7854, n7855, n7856,
    n7857, n7858, n7859, n7860, n7861, n7862,
    n7863, n7864, n7865, n7866, n7867, n7868,
    n7869, n7870, n7871, n7872, n7873, n7874,
    n7875, n7876, n7877, n7878, n7879, n7880,
    n7881, n7882, n7883, n7884, n7885, n7886,
    n7887, n7888, n7889, n7890, n7891, n7892,
    n7893, n7894, n7895, n7896, n7897, n7898,
    n7899, n7900, n7901, n7902, n7903, n7904,
    n7905, n7906, n7907, n7908, n7909, n7910,
    n7911, n7912, n7913, n7914, n7915, n7916,
    n7917, n7918, n7919, n7920, n7921, n7922,
    n7923, n7924, n7925, n7926, n7927, n7928,
    n7929, n7930, n7931, n7932, n7933, n7934,
    n7935, n7936, n7937, n7938, n7939, n7940,
    n7941, n7942, n7943, n7944, n7945, n7946,
    n7947, n7948, n7949, n7950, n7951, n7952,
    n7953, n7954, n7955, n7956, n7957, n7958,
    n7959, n7960, n7961, n7962, n7963, n7964,
    n7965, n7966, n7967, n7968, n7969, n7970,
    n7971, n7972, n7973, n7974, n7975, n7976,
    n7977, n7978, n7979, n7980, n7981, n7982,
    n7983, n7984, n7985, n7986, n7987, n7988,
    n7989, n7990, n7991, n7992, n7993, n7994,
    n7995, n7996, n7997, n7998, n7999, n8000,
    n8001, n8002, n8003, n8004, n8005, n8006,
    n8007, n8008, n8009, n8010, n8011, n8012,
    n8013, n8014, n8015, n8016, n8017, n8018,
    n8019, n8020, n8021, n8022, n8023, n8024,
    n8025, n8026, n8027, n8028, n8029, n8030,
    n8031, n8032, n8033, n8034, n8035, n8036,
    n8037, n8038, n8039, n8040, n8041, n8042,
    n8043, n8044, n8045, n8046, n8047, n8048,
    n8049, n8050, n8051, n8052, n8053, n8054,
    n8055, n8056, n8057, n8058, n8059, n8060,
    n8061, n8062, n8063, n8064, n8065, n8066,
    n8067, n8068, n8069, n8070, n8071, n8072,
    n8073, n8074, n8075, n8076, n8077, n8078,
    n8079, n8080, n8081, n8082, n8083, n8084,
    n8085, n8086, n8087, n8088, n8089, n8090,
    n8091, n8092, n8093, n8094, n8095, n8096,
    n8097, n8098, n8099, n8100, n8101, n8102,
    n8103, n8104, n8105, n8106, n8107, n8108,
    n8109, n8110, n8111, n8112, n8113, n8114,
    n8115, n8116, n8117, n8118, n8119, n8120,
    n8121, n8122, n8123, n8124, n8125, n8126,
    n8127, n8128, n8129, n8130, n8131, n8132,
    n8133, n8134, n8135, n8136, n8137, n8138,
    n8139, n8140, n8141, n8142, n8143, n8144,
    n8145, n8146, n8147, n8148, n8149, n8150,
    n8151, n8152, n8153, n8154, n8155, n8156,
    n8157, n8158, n8159, n8160, n8161, n8162,
    n8163, n8164, n8165, n8166, n8167, n8168,
    n8169, n8170, n8171, n8172, n8173, n8174,
    n8175, n8176, n8177, n8178, n8179, n8180,
    n8181, n8182, n8183, n8184, n8185, n8186,
    n8187, n8188, n8189, n8190, n8191, n8192,
    n8193, n8194, n8195, n8196, n8197, n8198,
    n8199, n8200, n8201, n8202, n8203, n8204,
    n8205, n8206, n8207, n8208, n8209, n8210,
    n8211, n8212, n8213, n8214, n8215, n8216,
    n8217, n8218, n8219, n8220, n8221, n8222,
    n8223, n8224, n8225, n8226, n8227, n8228,
    n8229, n8230, n8231, n8232, n8233, n8234,
    n8235, n8236, n8237, n8238, n8239, n8240,
    n8241, n8242, n8243, n8244, n8245, n8246,
    n8247, n8248, n8249, n8250, n8251, n8252,
    n8253, n8254, n8255, n8256, n8257, n8258,
    n8259, n8260, n8261, n8262, n8263, n8264,
    n8265, n8266, n8267, n8268, n8269, n8270,
    n8271, n8272, n8273, n8274, n8275, n8276,
    n8277, n8278, n8279, n8280, n8281, n8282,
    n8283, n8284, n8285, n8286, n8287, n8288,
    n8289, n8290, n8291, n8292, n8293, n8294,
    n8295, n8296, n8297, n8298, n8299, n8300,
    n8301, n8302, n8303, n8304, n8305, n8306,
    n8307, n8308, n8309, n8310, n8311, n8312,
    n8313, n8314, n8315, n8316, n8317, n8318,
    n8319, n8320, n8321, n8322, n8323, n8324,
    n8325, n8326, n8327, n8328, n8329, n8330,
    n8331, n8332, n8333, n8334, n8335, n8336,
    n8337, n8338, n8339, n8340, n8341, n8342,
    n8343, n8344, n8345, n8346, n8347, n8348,
    n8349, n8350, n8351, n8352, n8353, n8354,
    n8355, n8356, n8357, n8358, n8359, n8360,
    n8361, n8362, n8363, n8364, n8365, n8366,
    n8367, n8368, n8369, n8370, n8371, n8372,
    n8373, n8374, n8375, n8376, n8377, n8378,
    n8379, n8380, n8381, n8382, n8383, n8384,
    n8385, n8386, n8387, n8388, n8389, n8390,
    n8391, n8392, n8393, n8394, n8395, n8396,
    n8397, n8398, n8399, n8400, n8401, n8402,
    n8403, n8404, n8405, n8406, n8407, n8408,
    n8409, n8410, n8411, n8412, n8413, n8414,
    n8415, n8416, n8417, n8418, n8419, n8420,
    n8421, n8422, n8423, n8424, n8425, n8426,
    n8427, n8428, n8429, n8430, n8431, n8432,
    n8433, n8434, n8435, n8436, n8437, n8438,
    n8439, n8440, n8441, n8442, n8443, n8444,
    n8445, n8446, n8447, n8448, n8449, n8450,
    n8451, n8452, n8453, n8454, n8455, n8456,
    n8457, n8458, n8459, n8460, n8461, n8462,
    n8463, n8464, n8465, n8466, n8467, n8468,
    n8469, n8470, n8471, n8472, n8473, n8474,
    n8475, n8476, n8477, n8478, n8479, n8480,
    n8481, n8482, n8483, n8484, n8485, n8486,
    n8487, n8488, n8489, n8490, n8491, n8492,
    n8493, n8494, n8495, n8496, n8497, n8498,
    n8499, n8500, n8501, n8502, n8503, n8504,
    n8505, n8506, n8507, n8508, n8509, n8510,
    n8511, n8512, n8513, n8514, n8515, n8516,
    n8517, n8518, n8519, n8520, n8521, n8522,
    n8523, n8524, n8525, n8526, n8527, n8528,
    n8529, n8530, n8531, n8532, n8533, n8534,
    n8535, n8536, n8537, n8538, n8539, n8540,
    n8541, n8542, n8543, n8544, n8545, n8546,
    n8547, n8548, n8549, n8550, n8551, n8552,
    n8553, n8554, n8555, n8556, n8557, n8558,
    n8559, n8560, n8561, n8562, n8563, n8564,
    n8565, n8566, n8567, n8568, n8569, n8570,
    n8571, n8572, n8573, n8574, n8575, n8576,
    n8577, n8578, n8579, n8580, n8581, n8582,
    n8583, n8584, n8585, n8586, n8587, n8588,
    n8589, n8590, n8591, n8592, n8593, n8594,
    n8595, n8596, n8597, n8598, n8599, n8600,
    n8601, n8602, n8603, n8604, n8605, n8606,
    n8607, n8608, n8609, n8610, n8611, n8612,
    n8613, n8614, n8615, n8616, n8617, n8618,
    n8619, n8620, n8621, n8622, n8623, n8624,
    n8625, n8626, n8627, n8628, n8629, n8630,
    n8631, n8632, n8633, n8634, n8635, n8636,
    n8637, n8638, n8639, n8640, n8641, n8642,
    n8643, n8644, n8645, n8646, n8647, n8648,
    n8649, n8650, n8651, n8652, n8653, n8654,
    n8655, n8656, n8657, n8658, n8659, n8660,
    n8661, n8662, n8663, n8664, n8665, n8666,
    n8667, n8668, n8669, n8670, n8671, n8672,
    n8673, n8674, n8675, n8676, n8677, n8678,
    n8679, n8680, n8681, n8682, n8683, n8684,
    n8685, n8686, n8687, n8688, n8689, n8690,
    n8691, n8692, n8693, n8694, n8695, n8696,
    n8697, n8698, n8699, n8700, n8701, n8702,
    n8703, n8704, n8705, n8706, n8707, n8708,
    n8709, n8710, n8711, n8712, n8713, n8714,
    n8715, n8716, n8717, n8718, n8719, n8720,
    n8721, n8722, n8723, n8724, n8725, n8726,
    n8727, n8728, n8729, n8730, n8731, n8732,
    n8733, n8734, n8735, n8736, n8737, n8738,
    n8739, n8740, n8741, n8742, n8743, n8744,
    n8745, n8746, n8747, n8748, n8749, n8750,
    n8751, n8752, n8753, n8754, n8755, n8756,
    n8757, n8758, n8759, n8760, n8761, n8762,
    n8763, n8764, n8765, n8766, n8767, n8768,
    n8769, n8770, n8771, n8772, n8773, n8774,
    n8775, n8776, n8777, n8778, n8779, n8780,
    n8781, n8782, n8783, n8784, n8785, n8786,
    n8787, n8788, n8789, n8790, n8791, n8792,
    n8793, n8794, n8795, n8796, n8797, n8798,
    n8799, n8800, n8801, n8802, n8803, n8804,
    n8805, n8806, n8807, n8808, n8809, n8810,
    n8811, n8812, n8813, n8814, n8815, n8816,
    n8817, n8818, n8819, n8820, n8821, n8822,
    n8823, n8824, n8825, n8826, n8827, n8828,
    n8829, n8830, n8831, n8832, n8833, n8834,
    n8835, n8836, n8837, n8838, n8839, n8840,
    n8841, n8842, n8843, n8844, n8845, n8846,
    n8847, n8848, n8849, n8850, n8851, n8852,
    n8853, n8854, n8855, n8856, n8857, n8858,
    n8859, n8860, n8861, n8862, n8863, n8864,
    n8865, n8866, n8867, n8868, n8869, n8870,
    n8871, n8872, n8873, n8874, n8875, n8876,
    n8877, n8878, n8879, n8880, n8881, n8882,
    n8883, n8884, n8885, n8886, n8887, n8888,
    n8889, n8890, n8891, n8892, n8893, n8894,
    n8895, n8896, n8897, n8898, n8899, n8900,
    n8901, n8902, n8903, n8904, n8905, n8906,
    n8907, n8908, n8909, n8910, n8911, n8912,
    n8913, n8914, n8915, n8916, n8917, n8918,
    n8919, n8920, n8921, n8922, n8923, n8924,
    n8925, n8926, n8927, n8928, n8929, n8930,
    n8931, n8932, n8933, n8934, n8935, n8936,
    n8937, n8938, n8939, n8940, n8941, n8942,
    n8943, n8944, n8945, n8946, n8947, n8948,
    n8949, n8950, n8951, n8952, n8953, n8954,
    n8955, n8956, n8957, n8958, n8959, n8960,
    n8961, n8962, n8963, n8964, n8965, n8966,
    n8967, n8968, n8969, n8970, n8971, n8972,
    n8973, n8974, n8975, n8976, n8977, n8978,
    n8979, n8980, n8981, n8982, n8983, n8984,
    n8985, n8986, n8987, n8988, n8989, n8990,
    n8991, n8992, n8993, n8994, n8995, n8996,
    n8997, n8998, n8999, n9000, n9001, n9002,
    n9003, n9004, n9005, n9006, n9007, n9008,
    n9009, n9010, n9011, n9012, n9013, n9014,
    n9015, n9016, n9017, n9018, n9019, n9020,
    n9021, n9022, n9023, n9024, n9025, n9026,
    n9027, n9028, n9029, n9030, n9031, n9032,
    n9033, n9034, n9035, n9036, n9037, n9038,
    n9039, n9040, n9041, n9042, n9043, n9044,
    n9045, n9046, n9047, n9048, n9049, n9050,
    n9051, n9052, n9053, n9054, n9055, n9056,
    n9057, n9058, n9059, n9060, n9061, n9062,
    n9063, n9064, n9065, n9066, n9067, n9068,
    n9069, n9070, n9071, n9072, n9073, n9074,
    n9075, n9076, n9077, n9078, n9079, n9080,
    n9081, n9082, n9083, n9084, n9085, n9086,
    n9087, n9088, n9089, n9090, n9091, n9092,
    n9093, n9094, n9095, n9096, n9097, n9098,
    n9099, n9100, n9101, n9102, n9103, n9104,
    n9105, n9106, n9107, n9108, n9109, n9110,
    n9111, n9112, n9113, n9114, n9115, n9116,
    n9117, n9118, n9119, n9120, n9121, n9122,
    n9123, n9124, n9125, n9126, n9127, n9128,
    n9129, n9130, n9131, n9132, n9133, n9134,
    n9135, n9136, n9137, n9138, n9139, n9140,
    n9141, n9142, n9143, n9144, n9145, n9146,
    n9147, n9148, n9149, n9150, n9151, n9152,
    n9153, n9154, n9155, n9156, n9157, n9158,
    n9159, n9160, n9161, n9162, n9163, n9164,
    n9165, n9166, n9167, n9168, n9169, n9170,
    n9171, n9172, n9173, n9174, n9175, n9176,
    n9177, n9178, n9179, n9180, n9181, n9182,
    n9183, n9184, n9185, n9186, n9187, n9188,
    n9189, n9190, n9191, n9192, n9193, n9194,
    n9195, n9196, n9197, n9198, n9199, n9200,
    n9201, n9202, n9203, n9204, n9205, n9206,
    n9207, n9208, n9209, n9210, n9211, n9212,
    n9213, n9214, n9215, n9216, n9217, n9218,
    n9219, n9220, n9221, n9222, n9223, n9224,
    n9225, n9226, n9227, n9228, n9229, n9230,
    n9231, n9232, n9233, n9234, n9235, n9236,
    n9237, n9238, n9239, n9240, n9241, n9242,
    n9243, n9244, n9245, n9246, n9247, n9248,
    n9249, n9250, n9251, n9252, n9253, n9254,
    n9255, n9256, n9257, n9258, n9259, n9260,
    n9261, n9262, n9263, n9264, n9265, n9266,
    n9267, n9268, n9269, n9270, n9271, n9272,
    n9273, n9274, n9275, n9276, n9277, n9278,
    n9279, n9280, n9281, n9282, n9283, n9284,
    n9285, n9286, n9287, n9288, n9289, n9290,
    n9291, n9292, n9293, n9294, n9295, n9296,
    n9297, n9298, n9299, n9300, n9301, n9302,
    n9303, n9304, n9305, n9306, n9307, n9308,
    n9309, n9310, n9311, n9312, n9313, n9314,
    n9315, n9316, n9317, n9318, n9319, n9320,
    n9321, n9322, n9323, n9324, n9325, n9326,
    n9327, n9328, n9329, n9330, n9331, n9332,
    n9333, n9334, n9335, n9336, n9337, n9338,
    n9339, n9340, n9341, n9342, n9343, n9344,
    n9345, n9346, n9347, n9348, n9349, n9350,
    n9351, n9352, n9353, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386,
    n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416,
    n9417, n9418, n9419, n9420, n9421, n9422,
    n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446,
    n9447, n9448, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9703, n9704,
    n9705, n9706, n9707, n9708, n9709, n9710,
    n9711, n9712, n9713, n9714, n9715, n9716,
    n9717, n9718, n9719, n9720, n9721, n9722,
    n9723, n9724, n9725, n9726, n9727, n9728,
    n9729, n9730, n9731, n9732, n9733, n9734,
    n9735, n9736, n9737, n9738, n9739, n9740,
    n9741, n9742, n9743, n9744, n9745, n9746,
    n9747, n9748, n9749, n9750, n9751, n9752,
    n9753, n9754, n9755, n9756, n9757, n9758,
    n9759, n9760, n9761, n9762, n9763, n9764,
    n9765, n9766, n9767, n9768, n9769, n9770,
    n9771, n9772, n9773, n9774, n9775, n9776,
    n9777, n9778, n9779, n9780, n9781, n9782,
    n9783, n9784, n9785, n9786, n9787, n9788,
    n9789, n9790, n9791, n9792, n9793, n9794,
    n9795, n9796, n9797, n9798, n9799, n9800,
    n9801, n9802, n9803, n9804, n9805, n9806,
    n9807, n9808, n9809, n9810, n9811, n9812,
    n9813, n9814, n9815, n9816, n9817, n9818,
    n9819, n9820, n9821, n9822, n9823, n9824,
    n9825, n9826, n9827, n9828, n9829, n9830,
    n9831, n9832, n9833, n9834, n9835, n9836,
    n9837, n9838, n9839, n9840, n9841, n9842,
    n9843, n9844, n9845, n9846, n9847, n9848,
    n9849, n9850, n9851, n9852, n9853, n9854,
    n9855, n9856, n9857, n9858, n9859, n9860,
    n9861, n9862, n9863, n9864, n9865, n9866,
    n9867, n9868, n9869, n9870, n9871, n9872,
    n9873, n9874, n9875, n9876, n9877, n9878,
    n9879, n9880, n9881, n9882, n9883, n9884,
    n9885, n9886, n9887, n9888, n9889, n9890,
    n9891, n9892, n9893, n9894, n9895, n9896,
    n9897, n9898, n9899, n9900, n9901, n9902,
    n9903, n9904, n9905, n9906, n9907, n9908,
    n9909, n9910, n9911, n9912, n9913, n9914,
    n9915, n9916, n9917, n9918, n9919, n9920,
    n9921, n9922, n9923, n9924, n9925, n9926,
    n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052,
    n10053, n10054, n10055, n10056, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064,
    n10065, n10066, n10067, n10068, n10069, n10070,
    n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10082,
    n10083, n10084, n10085, n10086, n10087, n10088,
    n10089, n10090, n10091, n10092, n10093, n10094,
    n10095, n10096, n10097, n10098, n10099, n10100,
    n10101, n10102, n10103, n10104, n10105, n10106,
    n10107, n10108, n10109, n10110, n10111, n10112,
    n10113, n10114, n10115, n10116, n10117, n10118,
    n10119, n10120, n10121, n10122, n10123, n10124,
    n10125, n10126, n10127, n10128, n10129, n10130,
    n10131, n10132, n10133, n10134, n10135, n10136,
    n10137, n10138, n10139, n10140, n10141, n10142,
    n10143, n10144, n10145, n10146, n10147, n10148,
    n10149, n10150, n10151, n10152, n10153, n10154,
    n10155, n10156, n10157, n10158, n10159, n10160,
    n10161, n10162, n10163, n10164, n10165, n10166,
    n10167, n10168, n10169, n10170, n10171, n10172,
    n10173, n10174, n10175, n10176, n10177, n10178,
    n10179, n10180, n10181, n10182, n10183, n10184,
    n10185, n10186, n10187, n10188, n10189, n10190,
    n10191, n10192, n10193, n10194, n10195, n10196,
    n10197, n10198, n10199, n10200, n10201, n10202,
    n10203, n10204, n10205, n10206, n10207, n10208,
    n10209, n10210, n10211, n10212, n10213, n10214,
    n10215, n10216, n10217, n10218, n10219, n10220,
    n10221, n10222, n10223, n10224, n10225, n10226,
    n10227, n10228, n10229, n10230, n10231, n10232,
    n10233, n10234, n10235, n10236, n10237, n10238,
    n10239, n10240, n10241, n10242, n10243, n10244,
    n10245, n10246, n10247, n10248, n10249, n10250,
    n10251, n10252, n10253, n10254, n10255, n10256,
    n10257, n10258, n10259, n10260, n10261, n10262,
    n10263, n10264, n10265, n10266, n10267, n10268,
    n10269, n10270, n10271, n10272, n10273, n10274,
    n10275, n10276, n10277, n10278, n10279, n10280,
    n10281, n10282, n10283, n10284, n10285, n10286,
    n10287, n10288, n10289, n10290, n10291, n10292,
    n10293, n10294, n10295, n10296, n10297, n10298,
    n10299, n10300, n10301, n10302, n10303, n10304,
    n10305, n10306, n10307, n10308, n10309, n10310,
    n10311, n10312, n10313, n10314, n10315, n10316,
    n10317, n10318, n10319, n10320, n10321, n10322,
    n10323, n10324, n10325, n10326, n10327, n10328,
    n10329, n10330, n10331, n10332, n10333, n10334,
    n10335, n10336, n10337, n10338, n10339, n10340,
    n10341, n10342, n10343, n10344, n10345, n10346,
    n10347, n10348, n10349, n10350, n10351, n10352,
    n10353, n10354, n10355, n10356, n10357, n10358,
    n10359, n10360, n10361, n10362, n10363, n10364,
    n10365, n10366, n10367, n10368, n10369, n10370,
    n10371, n10372, n10373, n10374, n10375, n10376,
    n10377, n10378, n10379, n10380, n10381, n10382,
    n10383, n10384, n10385, n10386, n10387, n10388,
    n10389, n10390, n10391, n10392, n10393, n10394,
    n10395, n10396, n10397, n10398, n10399, n10400,
    n10401, n10402, n10403, n10404, n10405, n10406,
    n10407, n10408, n10409, n10410, n10411, n10412,
    n10413, n10414, n10415, n10416, n10417, n10418,
    n10419, n10420, n10421, n10422, n10423, n10424,
    n10425, n10426, n10427, n10428, n10429, n10430,
    n10431, n10432, n10433, n10434, n10435, n10436,
    n10437, n10438, n10439, n10440, n10441, n10442,
    n10443, n10444, n10445, n10446, n10447, n10448,
    n10449, n10450, n10451, n10452, n10453, n10454,
    n10455, n10456, n10457, n10458, n10459, n10460,
    n10461, n10462, n10463, n10464, n10465, n10466,
    n10467, n10468, n10469, n10470, n10471, n10472,
    n10473, n10474, n10475, n10476, n10477, n10478,
    n10479, n10480, n10481, n10482, n10483, n10484,
    n10485, n10486, n10487, n10488, n10489, n10490,
    n10491, n10492, n10493, n10494, n10495, n10496,
    n10497, n10498, n10499, n10500, n10501, n10502,
    n10503, n10504, n10505, n10506, n10507, n10508,
    n10509, n10510, n10511, n10512, n10513, n10514,
    n10515, n10516, n10517, n10518, n10519, n10520,
    n10521, n10522, n10523, n10524, n10525, n10526,
    n10527, n10528, n10529, n10530, n10531, n10532,
    n10533, n10534, n10535, n10536, n10537, n10538,
    n10539, n10540, n10541, n10542, n10543, n10544,
    n10545, n10546, n10547, n10548, n10549, n10550,
    n10551, n10552, n10553, n10554, n10555, n10556,
    n10557, n10558, n10559, n10560, n10561, n10562,
    n10563, n10564, n10565, n10566, n10567, n10568,
    n10569, n10570, n10571, n10572, n10573, n10574,
    n10575, n10576, n10577, n10578, n10579, n10580,
    n10581, n10582, n10583, n10584, n10585, n10586,
    n10587, n10588, n10589, n10590, n10591, n10592,
    n10593, n10594, n10595, n10596, n10597, n10598,
    n10599, n10600, n10601, n10602, n10603, n10604,
    n10605, n10606, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10651, n10652,
    n10653, n10654, n10655, n10656, n10657, n10658,
    n10659, n10660, n10661, n10662, n10663, n10664,
    n10665, n10666, n10667, n10668, n10669, n10670,
    n10671, n10672, n10673, n10674, n10675, n10676,
    n10677, n10678, n10679, n10680, n10681, n10682,
    n10683, n10684, n10685, n10686, n10687, n10688,
    n10689, n10690, n10691, n10692, n10693, n10694,
    n10695, n10696, n10697, n10698, n10699, n10700,
    n10701, n10702, n10703, n10704, n10705, n10706,
    n10707, n10708, n10709, n10710, n10711, n10712,
    n10713, n10714, n10715, n10716, n10717, n10718,
    n10719, n10720, n10721, n10722, n10723, n10724,
    n10725, n10726, n10727, n10728, n10729, n10730,
    n10731, n10732, n10733, n10734, n10735, n10736,
    n10737, n10738, n10739, n10740, n10741, n10742,
    n10743, n10744, n10745, n10746, n10747, n10748,
    n10749, n10750, n10751, n10752, n10753, n10754,
    n10755, n10756, n10757, n10758, n10759, n10760,
    n10761, n10762, n10763, n10764, n10765, n10766,
    n10767, n10768, n10769, n10770, n10771, n10772,
    n10773, n10774, n10775, n10776, n10777, n10778,
    n10779, n10780, n10781, n10782, n10783, n10784,
    n10785, n10786, n10787, n10788, n10789, n10790,
    n10791, n10792, n10793, n10794, n10795, n10796,
    n10797, n10798, n10799, n10800, n10801, n10802,
    n10803, n10804, n10805, n10806, n10807, n10808,
    n10809, n10810, n10811, n10812, n10813, n10814,
    n10815, n10816, n10817, n10818, n10819, n10820,
    n10821, n10822, n10823, n10824, n10825, n10826,
    n10827, n10828, n10829, n10830, n10831, n10832,
    n10833, n10834, n10835, n10836, n10837, n10838,
    n10839, n10840, n10841, n10842, n10843, n10844,
    n10845, n10846, n10847, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10859, n10860, n10861, n10862,
    n10863, n10864, n10865, n10866, n10867, n10868,
    n10869, n10870, n10871, n10872, n10873, n10874,
    n10875, n10876, n10877, n10878, n10879, n10880,
    n10881, n10882, n10883, n10884, n10885, n10886,
    n10887, n10888, n10889, n10890, n10891, n10892,
    n10893, n10894, n10895, n10896, n10897, n10898,
    n10899, n10900, n10901, n10902, n10903, n10904,
    n10905, n10906, n10907, n10908, n10909, n10910,
    n10911, n10912, n10913, n10914, n10915, n10916,
    n10917, n10918, n10919, n10920, n10921, n10922,
    n10923, n10924, n10925, n10926, n10927, n10928,
    n10929, n10930, n10931, n10932, n10933, n10934,
    n10935, n10936, n10937, n10938, n10939, n10940,
    n10941, n10942, n10943, n10944, n10945, n10946,
    n10947, n10948, n10949, n10950, n10951, n10952,
    n10953, n10954, n10955, n10956, n10957, n10958,
    n10959, n10960, n10961, n10962, n10963, n10964,
    n10965, n10966, n10967, n10968, n10969, n10970,
    n10971, n10972, n10973, n10974, n10975, n10976,
    n10977, n10978, n10979, n10980, n10981, n10982,
    n10983, n10984, n10985, n10986, n10987, n10988,
    n10989, n10990, n10991, n10992, n10993, n10994,
    n10995, n10996, n10997, n10998, n10999, n11000,
    n11001, n11002, n11003, n11004, n11005, n11006,
    n11007, n11008, n11009, n11010, n11011, n11012,
    n11013, n11014, n11015, n11016, n11017, n11018,
    n11019, n11020, n11021, n11022, n11023, n11024,
    n11025, n11026, n11027, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11048,
    n11049, n11050, n11051, n11052, n11053, n11054,
    n11055, n11056, n11057, n11058, n11059, n11060,
    n11061, n11062, n11063, n11064, n11065, n11066,
    n11067, n11068, n11069, n11070, n11071, n11072,
    n11073, n11074, n11075, n11076, n11077, n11078,
    n11079, n11080, n11081, n11082, n11083, n11084,
    n11085, n11086, n11087, n11088, n11089, n11090,
    n11091, n11092, n11093, n11094, n11095, n11096,
    n11097, n11098, n11099, n11100, n11101, n11102,
    n11103, n11104, n11105, n11106, n11107, n11108,
    n11109, n11110, n11111, n11112, n11113, n11114,
    n11115, n11116, n11117, n11118, n11119, n11120,
    n11121, n11122, n11123, n11124, n11125, n11126,
    n11127, n11128, n11129, n11130, n11131, n11132,
    n11133, n11134, n11135, n11136, n11137, n11138,
    n11139, n11140, n11141, n11142, n11143, n11144,
    n11145, n11146, n11147, n11148, n11149, n11150,
    n11151, n11152, n11153, n11154, n11155, n11156,
    n11157, n11158, n11159, n11160, n11161, n11162,
    n11163, n11164, n11165, n11166, n11167, n11168,
    n11169, n11170, n11171, n11172, n11173, n11174,
    n11175, n11176, n11177, n11178, n11179, n11180,
    n11181, n11182, n11183, n11184, n11185, n11186,
    n11187, n11188, n11189, n11190, n11191, n11192,
    n11193, n11194, n11195, n11196, n11197, n11198,
    n11199, n11200, n11201, n11202, n11203, n11204,
    n11205, n11206, n11207, n11208, n11209, n11210,
    n11211, n11212, n11213, n11214, n11215, n11216,
    n11217, n11218, n11219, n11220, n11221, n11222,
    n11223, n11224, n11225, n11226, n11227, n11228,
    n11229, n11230, n11231, n11232, n11233, n11234,
    n11235, n11236, n11237, n11238, n11239, n11240,
    n11241, n11242, n11243, n11244, n11245, n11246,
    n11247, n11248, n11249, n11250, n11251, n11252,
    n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11261, n11262, n11263, n11264,
    n11265, n11266, n11267, n11268, n11269, n11270,
    n11271, n11272, n11273, n11274, n11275, n11276,
    n11277, n11278, n11279, n11280, n11281, n11282,
    n11283, n11284, n11285, n11286, n11287, n11288,
    n11289, n11290, n11291, n11292, n11293, n11294,
    n11295, n11296, n11297, n11298, n11299, n11300,
    n11301, n11302, n11303, n11304, n11305, n11306,
    n11307, n11308, n11309, n11310, n11311, n11312,
    n11313, n11314, n11315, n11316, n11317, n11318,
    n11319, n11320, n11321, n11322, n11323, n11324,
    n11325, n11326, n11327, n11328, n11329, n11330,
    n11331, n11332, n11333, n11334, n11335, n11336,
    n11337, n11338, n11339, n11340, n11341, n11342,
    n11343, n11344, n11345, n11346, n11347, n11348,
    n11349, n11350, n11351, n11352, n11353, n11354,
    n11355, n11356, n11357, n11358, n11359, n11360,
    n11361, n11362, n11363, n11364, n11365, n11366,
    n11367, n11368, n11369, n11370, n11371, n11372,
    n11373, n11374, n11375, n11376, n11377, n11378,
    n11379, n11380, n11381, n11382, n11383, n11384,
    n11385, n11386, n11387, n11388, n11389, n11390,
    n11391, n11392, n11393, n11394, n11395, n11396,
    n11397, n11398, n11399, n11400, n11401, n11402,
    n11403, n11404, n11405, n11406, n11407, n11408,
    n11409, n11410, n11411, n11412, n11413, n11414,
    n11415, n11416, n11417, n11418, n11419, n11420,
    n11421, n11422, n11423, n11424, n11425, n11426,
    n11427, n11428, n11429, n11430, n11431, n11432,
    n11433, n11434, n11435, n11436, n11437, n11438,
    n11439, n11440, n11441, n11442, n11443, n11444,
    n11445, n11446, n11447, n11448, n11449, n11450,
    n11451, n11452, n11453, n11454, n11455, n11456,
    n11457, n11458, n11459, n11460, n11461, n11462,
    n11463, n11464, n11465, n11466, n11467, n11468,
    n11469, n11470, n11471, n11472, n11473, n11474,
    n11475, n11476, n11477, n11478, n11479, n11480,
    n11481, n11482, n11483, n11484, n11485, n11486,
    n11487, n11488, n11489, n11490, n11491, n11492,
    n11493, n11494, n11495, n11496, n11497, n11498,
    n11499, n11500, n11501, n11502, n11503, n11504,
    n11505, n11506, n11507, n11508, n11509, n11510,
    n11511, n11512, n11513, n11514, n11515, n11516,
    n11517, n11518, n11519, n11520, n11521, n11522,
    n11523, n11524, n11525, n11526, n11527, n11528,
    n11529, n11530, n11531, n11532, n11533, n11534,
    n11535, n11536, n11537, n11538, n11539, n11540,
    n11541, n11542, n11543, n11544, n11545, n11546,
    n11547, n11548, n11549, n11550, n11551, n11552,
    n11553, n11554, n11555, n11556, n11557, n11558,
    n11559, n11560, n11561, n11562, n11563, n11564,
    n11565, n11566, n11567, n11568, n11569, n11570,
    n11571, n11572, n11573, n11574, n11575, n11576,
    n11577, n11578, n11579, n11580, n11581, n11582,
    n11583, n11584, n11585, n11586, n11587, n11588,
    n11589, n11590, n11591, n11592, n11593, n11594,
    n11595, n11596, n11597, n11598, n11599, n11600,
    n11601, n11602, n11603, n11604, n11605, n11606,
    n11607, n11608, n11609, n11610, n11611, n11612,
    n11613, n11614, n11615, n11616, n11617, n11618,
    n11619, n11620, n11621, n11622, n11623, n11624,
    n11625, n11626, n11627, n11628, n11629, n11630,
    n11631, n11632, n11633, n11634, n11635, n11636,
    n11637, n11638, n11639, n11640, n11641, n11642,
    n11643, n11644, n11645, n11646, n11647, n11648,
    n11649, n11650, n11651, n11652, n11653, n11654,
    n11655, n11656, n11657, n11658, n11659, n11660,
    n11661, n11662, n11663, n11664, n11665, n11666,
    n11667, n11668, n11669, n11670, n11671, n11672,
    n11673, n11674, n11675, n11676, n11677, n11678,
    n11679, n11680, n11681, n11682, n11683, n11684,
    n11685, n11686, n11687, n11688, n11689, n11690,
    n11691, n11692, n11693, n11694, n11695, n11696,
    n11697, n11698, n11699, n11700, n11701, n11702,
    n11703, n11704, n11705, n11706, n11707, n11708,
    n11709, n11710, n11711, n11712, n11713, n11714,
    n11715, n11716, n11717, n11718, n11719, n11720,
    n11721, n11722, n11723, n11724, n11725, n11726,
    n11727, n11728, n11729, n11730, n11731, n11732,
    n11733, n11734, n11735, n11736, n11737, n11738,
    n11739, n11740, n11741, n11742, n11743, n11744,
    n11745, n11746, n11747, n11748, n11749, n11750,
    n11751, n11752, n11753, n11754, n11755, n11756,
    n11757, n11758, n11759, n11760, n11761, n11762,
    n11763, n11764, n11765, n11766, n11767, n11768,
    n11769, n11770, n11771, n11772, n11773, n11774,
    n11775, n11776, n11777, n11778, n11779, n11780,
    n11781, n11782, n11783, n11784, n11785, n11786,
    n11787, n11788, n11789, n11790, n11791, n11792,
    n11793, n11794, n11795, n11796, n11797, n11798,
    n11799, n11800, n11801, n11802, n11803, n11804,
    n11805, n11806, n11807, n11808, n11809, n11810,
    n11811, n11812, n11813, n11814, n11815, n11816,
    n11817, n11818, n11819, n11820, n11821, n11822,
    n11823, n11824, n11825, n11826, n11827, n11828,
    n11829, n11830, n11831, n11832, n11833, n11834,
    n11835, n11836, n11837, n11838, n11839, n11840,
    n11841, n11842, n11843, n11844, n11845, n11846,
    n11847, n11848, n11849, n11850, n11851, n11852,
    n11853, n11854, n11855, n11856, n11857, n11858,
    n11859, n11860, n11861, n11862, n11863, n11864,
    n11865, n11866, n11867, n11868, n11869, n11870,
    n11871, n11872, n11873, n11874, n11875, n11876,
    n11877, n11878, n11879, n11880, n11881, n11882,
    n11883, n11884, n11885, n11886, n11887, n11888,
    n11889, n11890, n11891, n11892, n11893, n11894,
    n11895, n11896, n11897, n11898, n11899, n11900,
    n11901, n11902, n11903, n11904, n11905, n11906,
    n11907, n11908, n11909, n11910, n11911, n11912,
    n11913, n11914, n11915, n11916, n11917, n11918,
    n11919, n11920, n11921, n11922, n11923, n11924,
    n11925, n11926, n11927, n11928, n11929, n11930,
    n11931, n11932, n11933, n11934, n11935, n11936,
    n11937, n11938, n11939, n11940, n11941, n11942,
    n11943, n11944, n11945, n11946, n11947, n11948,
    n11949, n11950, n11951, n11952, n11953, n11954,
    n11955, n11956, n11957, n11958, n11959, n11960,
    n11961, n11962, n11963, n11964, n11965, n11966,
    n11967, n11968, n11969, n11970, n11971, n11972,
    n11973, n11974, n11975, n11976, n11977, n11978,
    n11979, n11980, n11981, n11982, n11983, n11984,
    n11985, n11986, n11987, n11988, n11989, n11990,
    n11991, n11992, n11993, n11994, n11995, n11996,
    n11997, n11998, n11999, n12000, n12001, n12002,
    n12003, n12004, n12005, n12006, n12007, n12008,
    n12009, n12010, n12011, n12012, n12013, n12014,
    n12015, n12016, n12017, n12018, n12019, n12020,
    n12021, n12022, n12023, n12024, n12025, n12026,
    n12027, n12028, n12029, n12030, n12031, n12032,
    n12033, n12034, n12035, n12036, n12037, n12038,
    n12039, n12040, n12041, n12042, n12043, n12044,
    n12045, n12046, n12047, n12048, n12049, n12050,
    n12051, n12052, n12053, n12054, n12055, n12056,
    n12057, n12058, n12059, n12060, n12061, n12062,
    n12063, n12064, n12065, n12066, n12067, n12068,
    n12069, n12070, n12071, n12072, n12073, n12074,
    n12075, n12076, n12077, n12078, n12079, n12080,
    n12081, n12082, n12083, n12084, n12085, n12086,
    n12087, n12088, n12089, n12090, n12091, n12092,
    n12093, n12094, n12095, n12096, n12097, n12098,
    n12099, n12100, n12101, n12102, n12103, n12104,
    n12105, n12106, n12107, n12108, n12109, n12110,
    n12111, n12112, n12113, n12114, n12115, n12116,
    n12117, n12118, n12119, n12120, n12121, n12122,
    n12123, n12124, n12125, n12126, n12127, n12128,
    n12129, n12130, n12131, n12132, n12133, n12134,
    n12135, n12136, n12137, n12138, n12139, n12140,
    n12141, n12142, n12143, n12144, n12145, n12146,
    n12147, n12148, n12149, n12150, n12151, n12152,
    n12153, n12154, n12155, n12156, n12157, n12158,
    n12159, n12160, n12161, n12162, n12163, n12164,
    n12165, n12166, n12167, n12168, n12169, n12170,
    n12171, n12172, n12173, n12174, n12175, n12176,
    n12177, n12178, n12179, n12180, n12181, n12182,
    n12183, n12184, n12185, n12186, n12187, n12188,
    n12189, n12190, n12191, n12192, n12193, n12194,
    n12195, n12196, n12197, n12198, n12199, n12200,
    n12201, n12202, n12203, n12204, n12205, n12206,
    n12207, n12208, n12209, n12210, n12211, n12212,
    n12213, n12214, n12215, n12216, n12217, n12218,
    n12219, n12220, n12221, n12222, n12223, n12224,
    n12225, n12226, n12227, n12228, n12229, n12230,
    n12231, n12232, n12233, n12234, n12235, n12236,
    n12237, n12238, n12239, n12240, n12241, n12242,
    n12243, n12244, n12245, n12246, n12247, n12248,
    n12249, n12250, n12251, n12252, n12253, n12254,
    n12255, n12256, n12257, n12258, n12259, n12260,
    n12261, n12262, n12263, n12264, n12265, n12266,
    n12267, n12268, n12269, n12270, n12271, n12272,
    n12273, n12274, n12275, n12276, n12277, n12278,
    n12279, n12280, n12281, n12282, n12283, n12284,
    n12285, n12286, n12287, n12288, n12289, n12290,
    n12291, n12292, n12293, n12294, n12295, n12296,
    n12297, n12298, n12299, n12300, n12301, n12302,
    n12303, n12304, n12305, n12306, n12307, n12308,
    n12309, n12310, n12311, n12312, n12313, n12314,
    n12315, n12316, n12317, n12318, n12319, n12320,
    n12321, n12322, n12323, n12324, n12325, n12326,
    n12327, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12340, n12341, n12342, n12343, n12344,
    n12345, n12346, n12347, n12348, n12349, n12350,
    n12351, n12352, n12353, n12354, n12355, n12356,
    n12357, n12358, n12359, n12360, n12361, n12362,
    n12363, n12364, n12365, n12366, n12367, n12368,
    n12369, n12370, n12371, n12372, n12373, n12374,
    n12375, n12376, n12377, n12378, n12379, n12380,
    n12381, n12382, n12383, n12384, n12385, n12386,
    n12387, n12388, n12389, n12390, n12391, n12392,
    n12393, n12394, n12395, n12396, n12397, n12398,
    n12399, n12400, n12401, n12402, n12403, n12404,
    n12405, n12406, n12407, n12408, n12409, n12410,
    n12411, n12412, n12413, n12414, n12415, n12416,
    n12417, n12418, n12419, n12420, n12421, n12422,
    n12423, n12424, n12425, n12426, n12427, n12428,
    n12429, n12430, n12431, n12432, n12433, n12434,
    n12435, n12436, n12437, n12438, n12439, n12440,
    n12441, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12451, n12452,
    n12453, n12454, n12455, n12456, n12457, n12458,
    n12459, n12460, n12461, n12462, n12463, n12464,
    n12465, n12466, n12467, n12468, n12469, n12470,
    n12471, n12472, n12473, n12474, n12475, n12476,
    n12477, n12478, n12479, n12480, n12481, n12482,
    n12483, n12484, n12485, n12486, n12487, n12488,
    n12489, n12490, n12491, n12492, n12493, n12494,
    n12495, n12496, n12497, n12498, n12499, n12500,
    n12501, n12502, n12503, n12504, n12505, n12506,
    n12507, n12508, n12509, n12510, n12511, n12512,
    n12513, n12514, n12515, n12516, n12517, n12518,
    n12519, n12520, n12521, n12522, n12523, n12524,
    n12525, n12526, n12527, n12528, n12529, n12530,
    n12531, n12532, n12533, n12534, n12535, n12536,
    n12537, n12538, n12539, n12540, n12541, n12542,
    n12543, n12544, n12545, n12546, n12547, n12548,
    n12549, n12550, n12551, n12552, n12553, n12554,
    n12555, n12556, n12557, n12558, n12559, n12560,
    n12561, n12562, n12563, n12564, n12565, n12566,
    n12567, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578,
    n12579, n12580, n12581, n12582, n12583, n12584,
    n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596,
    n12597, n12598, n12599, n12600, n12601, n12602,
    n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614,
    n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632,
    n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12644,
    n12645, n12646, n12647, n12648, n12649, n12650,
    n12651, n12652, n12653, n12654, n12655, n12656,
    n12657, n12658, n12659, n12660, n12661, n12662,
    n12663, n12664, n12665, n12666, n12667, n12668,
    n12669, n12670, n12671, n12672, n12673, n12674,
    n12675, n12676, n12677, n12678, n12679, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12691, n12692,
    n12693, n12694, n12695, n12696, n12697, n12698,
    n12699, n12700, n12701, n12702, n12703, n12704,
    n12705, n12706, n12707, n12708, n12709, n12710,
    n12711, n12712, n12713, n12714, n12715, n12716,
    n12717, n12718, n12719, n12720, n12721, n12722,
    n12723, n12724, n12725, n12726, n12727, n12728,
    n12729, n12730, n12731, n12732, n12733, n12734,
    n12735, n12736, n12737, n12738, n12739, n12740,
    n12741, n12742, n12743, n12744, n12745, n12746,
    n12747, n12748, n12749, n12750, n12751, n12752,
    n12753, n12754, n12755, n12756, n12757, n12758,
    n12759, n12760, n12761, n12762, n12763, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776,
    n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794,
    n12795, n12796, n12797, n12798, n12799, n12800,
    n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12810, n12811, n12812,
    n12813, n12814, n12815, n12816, n12817, n12818,
    n12819, n12820, n12821, n12822, n12823, n12824,
    n12825, n12826, n12827, n12828, n12829, n12830,
    n12831, n12832, n12833, n12834, n12835, n12836,
    n12837, n12838, n12839, n12840, n12841, n12842,
    n12843, n12844, n12845, n12846, n12847, n12848,
    n12849, n12850, n12851, n12852, n12853, n12854,
    n12855, n12856, n12857, n12858, n12859, n12860,
    n12861, n12862, n12863, n12864, n12865, n12866,
    n12867, n12868, n12869, n12870, n12871, n12872,
    n12873, n12874, n12875, n12876, n12877, n12878,
    n12879, n12880, n12881, n12882, n12883, n12884,
    n12885, n12886, n12887, n12888, n12889, n12890,
    n12891, n12892, n12893, n12894, n12895, n12896,
    n12897, n12898, n12899, n12900, n12901, n12902,
    n12903, n12904, n12905, n12906, n12907, n12908,
    n12909, n12910, n12911, n12912, n12913, n12914,
    n12915, n12916, n12917, n12918, n12919, n12920,
    n12921, n12922, n12923, n12924, n12925, n12926,
    n12927, n12928, n12929, n12930, n12931, n12932,
    n12933, n12934, n12935, n12936, n12937, n12938,
    n12939, n12940, n12941, n12942, n12943, n12944,
    n12945, n12946, n12947, n12948, n12949, n12950,
    n12951, n12952, n12953, n12954, n12955, n12956,
    n12957, n12958, n12959, n12960, n12961, n12962,
    n12963, n12964, n12965, n12966, n12967, n12968,
    n12969, n12970, n12971, n12972, n12973, n12974,
    n12975, n12976, n12977, n12978, n12979, n12980,
    n12981, n12982, n12983, n12984, n12985, n12986,
    n12987, n12988, n12989, n12990, n12991, n12992,
    n12993, n12994, n12995, n12996, n12997, n12998,
    n12999, n13000, n13001, n13002, n13003, n13004,
    n13005, n13006, n13007, n13008, n13009, n13010,
    n13011, n13012, n13013, n13014, n13015, n13016,
    n13017, n13018, n13019, n13020, n13021, n13022,
    n13023, n13024, n13025, n13026, n13027, n13028,
    n13029, n13030, n13031, n13032, n13033, n13034,
    n13035, n13036, n13037, n13038, n13039, n13040,
    n13041, n13042, n13043, n13044, n13045, n13046,
    n13047, n13048, n13049, n13050, n13051, n13052,
    n13053, n13054, n13055, n13056, n13057, n13058,
    n13059, n13060, n13061, n13062, n13063, n13064,
    n13065, n13066, n13067, n13068, n13069, n13070,
    n13071, n13072, n13073, n13074, n13075, n13076,
    n13077, n13078, n13079, n13080, n13081, n13082,
    n13083, n13084, n13085, n13086, n13087, n13088,
    n13089, n13090, n13091, n13092, n13093, n13094,
    n13095, n13096, n13097, n13098, n13099, n13100,
    n13101, n13102, n13103, n13104, n13105, n13106,
    n13107, n13108, n13109, n13110, n13111, n13112,
    n13113, n13114, n13115, n13116, n13117, n13118,
    n13119, n13120, n13121, n13122, n13123, n13124,
    n13125, n13126, n13127, n13128, n13129, n13130,
    n13131, n13132, n13133, n13134, n13135, n13136,
    n13137, n13138, n13139, n13140, n13141, n13142,
    n13143, n13144, n13145, n13146, n13147, n13148,
    n13149, n13150, n13151, n13152, n13153, n13154,
    n13155, n13156, n13157, n13158, n13159, n13160,
    n13161, n13162, n13163, n13164, n13165, n13166,
    n13167, n13168, n13169, n13170, n13171, n13172,
    n13173, n13174, n13175, n13176, n13177, n13178,
    n13179, n13180, n13181, n13182, n13183, n13184,
    n13185, n13186, n13187, n13188, n13189, n13190,
    n13191, n13192, n13193, n13194, n13195, n13196,
    n13197, n13198, n13199, n13200, n13201, n13202,
    n13203, n13204, n13205, n13206, n13207, n13208,
    n13209, n13210, n13211, n13212, n13213, n13214,
    n13215, n13216, n13217, n13218, n13219, n13220,
    n13221, n13222, n13223, n13224, n13225, n13226,
    n13227, n13228, n13229, n13230, n13231, n13232,
    n13233, n13234, n13235, n13236, n13237, n13238,
    n13239, n13240, n13241, n13242, n13243, n13244,
    n13245, n13246, n13247, n13248, n13249, n13250,
    n13251, n13252, n13253, n13254, n13255, n13256,
    n13257, n13258, n13259, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322,
    n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13354, n13355, n13356, n13357, n13358,
    n13359, n13360, n13361, n13362, n13363, n13364,
    n13365, n13366, n13367, n13368, n13369, n13370,
    n13371, n13372, n13373, n13374, n13375, n13376,
    n13377, n13378, n13379, n13380, n13381, n13382,
    n13383, n13384, n13385, n13386, n13387, n13388,
    n13389, n13390, n13391, n13392, n13393, n13394,
    n13395, n13396, n13397, n13398, n13399, n13400,
    n13401, n13402, n13403, n13404, n13405, n13406,
    n13407, n13408, n13409, n13410, n13411, n13412,
    n13413, n13414, n13415, n13416, n13417, n13418,
    n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430,
    n13431, n13432, n13433, n13434, n13435, n13436,
    n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448,
    n13449, n13450, n13451, n13452, n13453, n13454,
    n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13464, n13465, n13466,
    n13467, n13468, n13469, n13470, n13471, n13472,
    n13473, n13474, n13475, n13476, n13477, n13478,
    n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13486, n13487, n13488, n13489, n13490,
    n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502,
    n13503, n13504, n13505, n13506, n13507, n13508,
    n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13516, n13517, n13518, n13519, n13520,
    n13521, n13522, n13523, n13524, n13525, n13526,
    n13527, n13528, n13529, n13530, n13531, n13532,
    n13533, n13534, n13535, n13536, n13537, n13538,
    n13539, n13540, n13541, n13542, n13543, n13544,
    n13545, n13546, n13547, n13548, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562,
    n13563, n13564, n13565, n13566, n13567, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580,
    n13581, n13582, n13583, n13584, n13585, n13586,
    n13587, n13588, n13589, n13590, n13591, n13592,
    n13593, n13594, n13595, n13596, n13597, n13598,
    n13599, n13600, n13601, n13602, n13603, n13604,
    n13605, n13606, n13607, n13608, n13609, n13610,
    n13611, n13612, n13613, n13614, n13615, n13616,
    n13617, n13618, n13619, n13620, n13621, n13622,
    n13623, n13624, n13625, n13626, n13627, n13628,
    n13629, n13630, n13631, n13632, n13633, n13634,
    n13635, n13636, n13637, n13638, n13639, n13640,
    n13641, n13642, n13643, n13644, n13645, n13646,
    n13647, n13648, n13649, n13650, n13651, n13652,
    n13653, n13654, n13655, n13656, n13657, n13658,
    n13659, n13660, n13661, n13662, n13663, n13664,
    n13665, n13666, n13667, n13668, n13669, n13670,
    n13671, n13672, n13673, n13674, n13675, n13676,
    n13677, n13678, n13679, n13680, n13681, n13682,
    n13683, n13684, n13685, n13686, n13687, n13688,
    n13689, n13690, n13691, n13692, n13693, n13694,
    n13695, n13696, n13697, n13698, n13699, n13700,
    n13701, n13702, n13703, n13704, n13705, n13706,
    n13707, n13708, n13709, n13710, n13711, n13712,
    n13713, n13714, n13715, n13716, n13717, n13718,
    n13719, n13720, n13721, n13722, n13723, n13724,
    n13725, n13726, n13727, n13728, n13729, n13730,
    n13731, n13732, n13733, n13734, n13735, n13736,
    n13737, n13738, n13739, n13740, n13741, n13742,
    n13743, n13744, n13745, n13746, n13747, n13748,
    n13749, n13750, n13751, n13752, n13753, n13754,
    n13755, n13756, n13757, n13758, n13759, n13760,
    n13761, n13762, n13763, n13764, n13765, n13766,
    n13767, n13768, n13769, n13770, n13771, n13772,
    n13773, n13774, n13775, n13776, n13777, n13778,
    n13779, n13780, n13781, n13782, n13783, n13784,
    n13785, n13786, n13787, n13788, n13789, n13790,
    n13791, n13792, n13793, n13794, n13795, n13796,
    n13797, n13798, n13799, n13800, n13801, n13802,
    n13803, n13804, n13805, n13806, n13807, n13808,
    n13809, n13810, n13811, n13812, n13813, n13814,
    n13815, n13816, n13817, n13818, n13819, n13820,
    n13821, n13822, n13823, n13824, n13825, n13826,
    n13827, n13828, n13829, n13830, n13831, n13832,
    n13833, n13834, n13835, n13836, n13837, n13838,
    n13839, n13840, n13841, n13842, n13843, n13844,
    n13845, n13846, n13847, n13848, n13849, n13850,
    n13851, n13852, n13853, n13854, n13855, n13856,
    n13857, n13858, n13859, n13860, n13861, n13862,
    n13863, n13864, n13865, n13866, n13867, n13868,
    n13869, n13870, n13871, n13872, n13873, n13874,
    n13875, n13876, n13877, n13878, n13879, n13880,
    n13881, n13882, n13883, n13884, n13885, n13886,
    n13887, n13888, n13889, n13890, n13891, n13892,
    n13893, n13894, n13895, n13896, n13897, n13898,
    n13899, n13900, n13901, n13902, n13903, n13904,
    n13905, n13906, n13907, n13908, n13909, n13910,
    n13911, n13912, n13913, n13914, n13915, n13916,
    n13917, n13918, n13919, n13920, n13921, n13922,
    n13923, n13924, n13925, n13926, n13927, n13928,
    n13929, n13930, n13931, n13932, n13933, n13934,
    n13935, n13936, n13937, n13938, n13939, n13940,
    n13941, n13942, n13943, n13944, n13945, n13946,
    n13947, n13948, n13949, n13950, n13951, n13952,
    n13953, n13954, n13955, n13956, n13957, n13958,
    n13959, n13960, n13961, n13962, n13963, n13964,
    n13965, n13966, n13967, n13968, n13969, n13970,
    n13971, n13972, n13973, n13974, n13975, n13976,
    n13977, n13978, n13979, n13980, n13981, n13982,
    n13983, n13984, n13985, n13986, n13987, n13988,
    n13989, n13990, n13991, n13992, n13993, n13994,
    n13995, n13996, n13997, n13998, n13999, n14000,
    n14001, n14002, n14003, n14004, n14005, n14006,
    n14007, n14008, n14009, n14010, n14011, n14012,
    n14013, n14014, n14015, n14016, n14017, n14018,
    n14019, n14020, n14021, n14022, n14023, n14024,
    n14025, n14026, n14027, n14028, n14029, n14030,
    n14031, n14032, n14033, n14034, n14035, n14036,
    n14037, n14038, n14039, n14040, n14041, n14042,
    n14043, n14044, n14045, n14046, n14047, n14048,
    n14049, n14050, n14051, n14052, n14053, n14054,
    n14055, n14056, n14057, n14058, n14059, n14060,
    n14061, n14062, n14063, n14064, n14065, n14066,
    n14067, n14068, n14069, n14070, n14071, n14072,
    n14073, n14074, n14075, n14076, n14077, n14078,
    n14079, n14080, n14081, n14082, n14083, n14084,
    n14085, n14086, n14087, n14088, n14089, n14090,
    n14091, n14092, n14093, n14094, n14095, n14096,
    n14097, n14098, n14099, n14100, n14101, n14102,
    n14103, n14104, n14105, n14106, n14107, n14108,
    n14109, n14110, n14111, n14112, n14113, n14114,
    n14115, n14116, n14117, n14118, n14119, n14120,
    n14121, n14122, n14123, n14124, n14125, n14126,
    n14127, n14128, n14129, n14130, n14131, n14132,
    n14133, n14134, n14135, n14136, n14137, n14138,
    n14139, n14140, n14141, n14142, n14143, n14144,
    n14145, n14146, n14147, n14148, n14149, n14150,
    n14151, n14152, n14153, n14154, n14155, n14156,
    n14157, n14158, n14159, n14160, n14161, n14162,
    n14163, n14164, n14165, n14166, n14167, n14168,
    n14169, n14170, n14171, n14172, n14173, n14174,
    n14175, n14176, n14177, n14178, n14179, n14180,
    n14181, n14182, n14183, n14184, n14185, n14186,
    n14187, n14188, n14189, n14190, n14191, n14192,
    n14193, n14194, n14195, n14196, n14197, n14198,
    n14199, n14200, n14201, n14202, n14203, n14204,
    n14205, n14206, n14207, n14208, n14209, n14210,
    n14211, n14212, n14213, n14214, n14215, n14216,
    n14217, n14218, n14219, n14220, n14221, n14222,
    n14223, n14224, n14225, n14226, n14227, n14228,
    n14229, n14230, n14231, n14232, n14233, n14234,
    n14235, n14236, n14237, n14238, n14239, n14240,
    n14241, n14242, n14243, n14244, n14245, n14246,
    n14247, n14248, n14249, n14250, n14251, n14252,
    n14253, n14254, n14255, n14256, n14257, n14258,
    n14259, n14260, n14261, n14262, n14263, n14264,
    n14265, n14266, n14267, n14268, n14269, n14270,
    n14271, n14272, n14273, n14274, n14275, n14276,
    n14277, n14278, n14279, n14280, n14281, n14282,
    n14283, n14284, n14285, n14286, n14287, n14288,
    n14289, n14290, n14291, n14292, n14293, n14294,
    n14295, n14296, n14297, n14298, n14299, n14300,
    n14301, n14302, n14303, n14304, n14305, n14306,
    n14307, n14308, n14309, n14310, n14311, n14312,
    n14313, n14314, n14315, n14316, n14317, n14318,
    n14319, n14320, n14321, n14322, n14323, n14324,
    n14325, n14326, n14327, n14328, n14329, n14330,
    n14331, n14332, n14333, n14334, n14335, n14336,
    n14337, n14338, n14339, n14340, n14341, n14342,
    n14343, n14344, n14345, n14346, n14347, n14348,
    n14349, n14350, n14351, n14352, n14353, n14354,
    n14355, n14356, n14357, n14358, n14359, n14360,
    n14361, n14362, n14363, n14364, n14365, n14366,
    n14367, n14368, n14369, n14370, n14371, n14372,
    n14373, n14374, n14375, n14376, n14377, n14378,
    n14379, n14380, n14381, n14382, n14383, n14384,
    n14385, n14386, n14387, n14388, n14389, n14390,
    n14391, n14392, n14393, n14394, n14395, n14396,
    n14397, n14398, n14399, n14400, n14401, n14402,
    n14403, n14404, n14405, n14406, n14407, n14408,
    n14409, n14410, n14411, n14412, n14413, n14414,
    n14415, n14416, n14417, n14418, n14419, n14420,
    n14421, n14422, n14423, n14424, n14425, n14426,
    n14427, n14428, n14429, n14430, n14431, n14432,
    n14433, n14434, n14435, n14436, n14437, n14438,
    n14439, n14440, n14441, n14442, n14443, n14444,
    n14445, n14446, n14447, n14448, n14449, n14450,
    n14451, n14452, n14453, n14454, n14455, n14456,
    n14457, n14458, n14459, n14460, n14461, n14462,
    n14463, n14464, n14465, n14466, n14467, n14468,
    n14469, n14470, n14471, n14472, n14473, n14474,
    n14475, n14476, n14477, n14478, n14479, n14480,
    n14481, n14482, n14483, n14484, n14485, n14486,
    n14487, n14488, n14489, n14490, n14491, n14492,
    n14493, n14494, n14495, n14496, n14497, n14498,
    n14499, n14500, n14501, n14502, n14503, n14504,
    n14505, n14506, n14507, n14508, n14509, n14510,
    n14511, n14512, n14513, n14514, n14515, n14516,
    n14517, n14518, n14519, n14520, n14521, n14522,
    n14523, n14524, n14525, n14526, n14527, n14528,
    n14529, n14530, n14531, n14532, n14533, n14534,
    n14535, n14536, n14537, n14538, n14539, n14540,
    n14541, n14542, n14543, n14544, n14545, n14546,
    n14547, n14548, n14549, n14550, n14551, n14552,
    n14553, n14554, n14555, n14556, n14557, n14558,
    n14559, n14560, n14561, n14562, n14563, n14564,
    n14565, n14566, n14567, n14568, n14569, n14570,
    n14571, n14572, n14573, n14574, n14575, n14576,
    n14577, n14578, n14579, n14580, n14581, n14582,
    n14583, n14584, n14585, n14586, n14587, n14588,
    n14589, n14590, n14591, n14592, n14593, n14594,
    n14595, n14596, n14597, n14598, n14599, n14600,
    n14601, n14602, n14603, n14604, n14605, n14606,
    n14607, n14608, n14609, n14610, n14611, n14612,
    n14613, n14614, n14615, n14616, n14617, n14618,
    n14619, n14620, n14621, n14622, n14623, n14624,
    n14625, n14626, n14627, n14628, n14629, n14630,
    n14631, n14632, n14633, n14634, n14635, n14636,
    n14637, n14638, n14639, n14640, n14641, n14642,
    n14643, n14644, n14645, n14646, n14647, n14648,
    n14649, n14650, n14651, n14652, n14653, n14654,
    n14655, n14656, n14657, n14658, n14659, n14660,
    n14661, n14662, n14663, n14664, n14665, n14666,
    n14667, n14668, n14669, n14670, n14671, n14672,
    n14673, n14674, n14675, n14676, n14677, n14678,
    n14679, n14680, n14681, n14682, n14683, n14684,
    n14685, n14686, n14687, n14688, n14689, n14690,
    n14691, n14692, n14693, n14694, n14695, n14696,
    n14697, n14698, n14699, n14700, n14701, n14702,
    n14703, n14704, n14705, n14706, n14707, n14708,
    n14709, n14710, n14711, n14712, n14713, n14714,
    n14715, n14716, n14717, n14718, n14719, n14720,
    n14721, n14722, n14723, n14724, n14725, n14726,
    n14727, n14728, n14729, n14730, n14731, n14732,
    n14733, n14734, n14735, n14736, n14737, n14738,
    n14739, n14740, n14741, n14742, n14743, n14744,
    n14745, n14746, n14747, n14748, n14749, n14750,
    n14751, n14752, n14753, n14754, n14755, n14756,
    n14757, n14758, n14759, n14760, n14761, n14762,
    n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816,
    n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14830, n14831, n14832, n14833, n14834,
    n14835, n14836, n14837, n14838, n14839, n14840,
    n14841, n14842, n14843, n14844, n14845, n14846,
    n14847, n14848, n14849, n14850, n14851, n14852,
    n14853, n14854, n14855, n14856, n14857, n14858,
    n14859, n14860, n14861, n14862, n14863, n14864,
    n14865, n14866, n14867, n14868, n14869, n14870,
    n14871, n14872, n14873, n14874, n14875, n14876,
    n14877, n14878, n14879, n14880, n14881, n14882,
    n14883, n14884, n14885, n14886, n14887, n14888,
    n14889, n14890, n14891, n14892, n14893, n14894,
    n14895, n14896, n14897, n14898, n14899, n14900,
    n14901, n14902, n14903, n14904, n14905, n14906,
    n14907, n14908, n14909, n14910, n14911, n14912,
    n14913, n14914, n14915, n14916, n14917, n14918,
    n14919, n14920, n14921, n14922, n14923, n14924,
    n14925, n14926, n14927, n14928, n14929, n14930,
    n14931, n14932, n14933, n14934, n14935, n14936,
    n14937, n14938, n14939, n14940, n14941, n14942,
    n14943, n14944, n14945, n14946, n14947, n14948,
    n14949, n14950, n14951, n14952, n14953, n14954,
    n14955, n14956, n14957, n14958, n14959, n14960,
    n14961, n14962, n14963, n14964, n14965, n14966,
    n14967, n14968, n14969, n14970, n14971, n14972,
    n14973, n14974, n14975, n14976, n14977, n14978,
    n14979, n14980, n14981, n14982, n14983, n14984,
    n14985, n14986, n14987, n14988, n14989, n14990,
    n14991, n14992, n14993, n14994, n14995, n14996,
    n14997, n14998, n14999, n15000, n15001, n15002,
    n15003, n15004, n15005, n15006, n15007, n15008,
    n15009, n15010, n15011, n15012, n15013, n15014,
    n15015, n15016, n15017, n15018, n15019, n15020,
    n15021, n15022, n15023, n15024, n15025, n15026,
    n15027, n15028, n15029, n15030, n15031, n15032,
    n15033, n15034, n15035, n15036, n15037, n15038,
    n15039, n15040, n15041, n15042, n15043, n15044,
    n15045, n15046, n15047, n15048, n15049, n15050,
    n15051, n15052, n15053, n15054, n15055, n15056,
    n15057, n15058, n15059, n15060, n15061, n15062,
    n15063, n15064, n15065, n15066, n15067, n15068,
    n15069, n15070, n15071, n15072, n15073, n15074,
    n15075, n15076, n15077, n15078, n15079, n15080,
    n15081, n15082, n15083, n15084, n15085, n15086,
    n15087, n15088, n15089, n15090, n15091, n15092,
    n15093, n15094, n15095, n15096, n15097, n15098,
    n15099, n15100, n15101, n15102, n15103, n15104,
    n15105, n15106, n15107, n15108, n15109, n15110,
    n15111, n15112, n15113, n15114, n15115, n15116,
    n15117, n15118, n15119, n15120, n15121, n15122,
    n15123, n15124, n15125, n15126, n15127, n15128,
    n15129, n15130, n15131, n15132, n15133, n15134,
    n15135, n15136, n15137, n15138, n15139, n15140,
    n15141, n15142, n15143, n15144, n15145, n15146,
    n15147, n15148, n15149, n15150, n15151, n15152,
    n15153, n15154, n15155, n15156, n15157, n15158,
    n15159, n15160, n15161, n15162, n15163, n15164,
    n15165, n15166, n15167, n15168, n15169, n15170,
    n15171, n15172, n15173, n15174, n15175, n15176,
    n15177, n15178, n15179, n15180, n15181, n15182,
    n15183, n15184, n15185, n15186, n15187, n15188,
    n15189, n15190, n15191, n15192, n15193, n15194,
    n15195, n15196, n15197, n15198, n15199, n15200,
    n15201, n15202, n15203, n15204, n15205, n15206,
    n15207, n15208, n15209, n15210, n15211, n15212,
    n15213, n15214, n15215, n15216, n15217, n15218,
    n15219, n15220, n15221, n15222, n15223, n15224,
    n15225, n15226, n15227, n15228, n15229, n15230,
    n15231, n15232, n15233, n15234, n15235, n15236,
    n15237, n15238, n15239, n15240, n15241, n15242,
    n15243, n15244, n15245, n15246, n15247, n15248,
    n15249, n15250, n15251, n15252, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15281, n15282, n15283, n15284,
    n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302,
    n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314,
    n15315, n15316, n15317, n15318, n15319, n15320,
    n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338,
    n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15355, n15356,
    n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15365, n15366, n15367, n15368,
    n15369, n15370, n15371, n15372, n15373, n15374,
    n15375, n15376, n15377, n15378, n15379, n15380,
    n15381, n15382, n15383, n15384, n15385, n15386,
    n15387, n15388, n15389, n15390, n15391, n15392,
    n15393, n15394, n15395, n15396, n15397, n15398,
    n15399, n15400, n15401, n15402, n15403, n15404,
    n15405, n15406, n15407, n15408, n15409, n15410,
    n15411, n15412, n15413, n15414, n15415, n15416,
    n15417, n15418, n15419, n15420, n15421, n15422,
    n15423, n15424, n15425, n15426, n15427, n15428,
    n15429, n15430, n15431, n15432, n15433, n15434,
    n15435, n15436, n15437, n15438, n15439, n15440,
    n15441, n15442, n15443, n15444, n15445, n15446,
    n15447, n15448, n15449, n15450, n15451, n15452,
    n15453, n15454, n15455, n15456, n15457, n15458,
    n15459, n15460, n15461, n15462, n15463, n15464,
    n15465, n15466, n15467, n15468, n15469, n15470,
    n15471, n15472, n15473, n15474, n15475, n15476,
    n15477, n15478, n15479, n15480, n15481, n15482,
    n15483, n15484, n15485, n15486, n15487, n15488,
    n15489, n15490, n15491, n15492, n15493, n15494,
    n15495, n15496, n15497, n15498, n15499, n15500,
    n15501, n15502, n15503, n15504, n15505, n15506,
    n15507, n15508, n15509, n15510, n15511, n15512,
    n15513, n15514, n15515, n15516, n15517, n15518,
    n15519, n15520, n15521, n15522, n15523, n15524,
    n15525, n15526, n15527, n15528, n15529, n15530,
    n15531, n15532, n15533, n15534, n15535, n15536,
    n15537, n15538, n15539, n15540, n15541, n15542,
    n15543, n15544, n15545, n15546, n15547, n15548,
    n15549, n15550, n15551, n15552, n15553, n15554,
    n15555, n15556, n15557, n15558, n15559, n15560,
    n15561, n15562, n15563, n15564, n15565, n15566,
    n15567, n15568, n15569, n15570, n15571, n15572,
    n15573, n15574, n15575, n15576, n15577, n15578,
    n15579, n15580, n15581, n15582, n15583, n15584,
    n15585, n15586, n15587, n15588, n15589, n15590,
    n15591, n15592, n15593, n15594, n15595, n15596,
    n15597, n15598, n15599, n15600, n15601, n15602,
    n15603, n15604, n15605, n15606, n15607, n15608,
    n15609, n15610, n15611, n15612, n15613, n15614,
    n15615, n15616, n15617, n15618, n15619, n15620,
    n15621, n15622, n15623, n15624, n15625, n15626,
    n15627, n15628, n15629, n15630, n15631, n15632,
    n15633, n15634, n15635, n15636, n15637, n15638,
    n15639, n15640, n15641, n15642, n15643, n15644,
    n15645, n15646, n15647, n15648, n15649, n15650,
    n15651, n15652, n15653, n15654, n15655, n15656,
    n15657, n15658, n15659, n15660, n15661, n15662,
    n15663, n15664, n15665, n15666, n15667, n15668,
    n15669, n15670, n15671, n15672, n15673, n15674,
    n15675, n15676, n15677, n15678, n15679, n15680,
    n15681, n15682, n15683, n15684, n15685, n15686,
    n15687, n15688, n15689, n15690, n15691, n15692,
    n15693, n15694, n15695, n15696, n15697, n15698,
    n15699, n15700, n15701, n15702, n15703, n15704,
    n15705, n15706, n15707, n15708, n15709, n15710,
    n15711, n15712, n15713, n15714, n15715, n15716,
    n15717, n15718, n15719, n15720, n15721, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15768, n15769, n15770,
    n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782,
    n15783, n15784, n15785, n15786, n15787, n15788,
    n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800,
    n15801, n15802, n15803, n15804, n15805, n15806,
    n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824,
    n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854,
    n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872,
    n15873, n15874, n15875, n15876, n15877, n15878,
    n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890,
    n15891, n15892, n15893, n15894, n15895, n15896,
    n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908,
    n15909, n15910, n15911, n15912, n15913, n15914,
    n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926,
    n15927, n15928, n15929, n15930, n15931, n15932,
    n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944,
    n15945, n15946, n15947, n15948, n15949, n15950,
    n15951, n15952, n15953, n15954, n15955, n15956,
    n15957, n15958, n15959, n15960, n15961, n15962,
    n15963, n15964, n15965, n15966, n15967, n15968,
    n15969, n15970, n15971, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980,
    n15981, n15982, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998,
    n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016,
    n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034,
    n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106,
    n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178,
    n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196,
    n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214,
    n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232,
    n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250,
    n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262,
    n16263, n16264, n16265, n16266, n16267, n16268,
    n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280,
    n16281, n16282, n16283, n16284, n16285, n16286,
    n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16302, n16303, n16304,
    n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316,
    n16317, n16318, n16319, n16320, n16321, n16322,
    n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334,
    n16335, n16336, n16337, n16338, n16339, n16340,
    n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352,
    n16353, n16354, n16355, n16356, n16357, n16358,
    n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370,
    n16371, n16372, n16373, n16374, n16375, n16376,
    n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388,
    n16389, n16390, n16391, n16392, n16393, n16394,
    n16395, n16396, n16397, n16398, n16399, n16400,
    n16401, n16402, n16403, n16404, n16405, n16406,
    n16407, n16408, n16409, n16410, n16411, n16412,
    n16413, n16414, n16415, n16416, n16417, n16418,
    n16419, n16420, n16421, n16422, n16423, n16424,
    n16425, n16426, n16427, n16428, n16429, n16430,
    n16431, n16432, n16433, n16434, n16435, n16436,
    n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448,
    n16449, n16450, n16451, n16452, n16453, n16454,
    n16455, n16456, n16457, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466,
    n16467, n16468, n16469, n16470, n16471, n16472,
    n16473, n16474, n16475, n16476, n16477, n16478,
    n16479, n16480, n16481, n16482, n16483, n16484,
    n16485, n16486, n16487, n16488, n16489, n16490,
    n16491, n16492, n16493, n16494, n16495, n16496,
    n16497, n16498, n16499, n16500, n16501, n16502,
    n16503, n16504, n16505, n16506, n16507, n16508,
    n16509, n16510, n16511, n16512, n16513, n16514,
    n16515, n16516, n16517, n16518, n16519, n16520,
    n16521, n16522, n16523, n16524, n16525, n16526,
    n16527, n16528, n16529, n16530, n16531, n16532,
    n16533, n16534, n16535, n16536, n16537, n16538,
    n16539, n16540, n16541, n16542, n16543, n16544,
    n16545, n16546, n16547, n16548, n16549, n16550,
    n16551, n16552, n16553, n16554, n16555, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562,
    n16563, n16564, n16565, n16566, n16567, n16568,
    n16569, n16570, n16571, n16572, n16573, n16574,
    n16575, n16576, n16577, n16578, n16579, n16580,
    n16581, n16582, n16583, n16584, n16585, n16586,
    n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598,
    n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652,
    n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670,
    n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16687, n16688,
    n16689, n16690, n16691, n16692, n16693, n16694,
    n16695, n16696, n16697, n16698, n16699, n16700,
    n16701, n16702, n16703, n16704, n16705, n16706,
    n16707, n16708, n16709, n16710, n16711, n16712,
    n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724,
    n16725, n16726, n16727, n16728, n16729, n16730,
    n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742,
    n16743, n16744, n16745, n16746, n16747, n16748,
    n16749, n16750, n16751, n16752, n16753, n16754,
    n16755, n16756, n16757, n16758, n16759, n16760,
    n16761, n16762, n16763, n16764, n16765, n16766,
    n16767, n16768, n16769, n16770, n16771, n16772,
    n16773, n16774, n16775, n16776, n16777, n16778,
    n16779, n16780, n16781, n16782, n16783, n16784,
    n16785, n16786, n16787, n16788, n16789, n16790,
    n16791, n16792, n16793, n16794, n16795, n16796,
    n16797, n16798, n16799, n16800, n16801, n16802,
    n16803, n16804, n16805, n16806, n16807, n16808,
    n16809, n16810, n16811, n16812, n16813, n16814,
    n16815, n16816, n16817, n16818, n16819, n16820,
    n16821, n16822, n16823, n16824, n16825, n16826,
    n16827, n16828, n16829, n16830, n16831, n16832,
    n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844,
    n16845, n16846, n16847, n16848, n16849, n16850,
    n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16868,
    n16869, n16870, n16871, n16872, n16873, n16874,
    n16875, n16876, n16877, n16878, n16879, n16880,
    n16881, n16882, n16883, n16884, n16885, n16886,
    n16887, n16888, n16889, n16890, n16891, n16892,
    n16893, n16894, n16895, n16896, n16897, n16898,
    n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16906, n16907, n16908, n16909, n16910,
    n16911, n16912, n16913, n16914, n16915, n16916,
    n16917, n16918, n16919, n16920, n16921, n16922,
    n16923, n16924, n16925, n16926, n16927, n16928,
    n16929, n16930, n16931, n16932, n16933, n16934,
    n16935, n16936, n16937, n16938, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16952,
    n16953, n16954, n16955, n16956, n16957, n16958,
    n16959, n16960, n16961, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976,
    n16977, n16978, n16979, n16980, n16981, n16982,
    n16983, n16984, n16985, n16986, n16987, n16988,
    n16989, n16990, n16991, n16992, n16993, n16994,
    n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17004, n17005, n17006,
    n17007, n17008, n17009, n17010, n17011, n17012,
    n17013, n17014, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024,
    n17025, n17026, n17027, n17028, n17029, n17030,
    n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042,
    n17043, n17044, n17045, n17046, n17047, n17048,
    n17049, n17050, n17051, n17052, n17053, n17054,
    n17055, n17056, n17057, n17058, n17059, n17060,
    n17061, n17062, n17063, n17064, n17065, n17066,
    n17067, n17068, n17069, n17070, n17071, n17072,
    n17073, n17074, n17075, n17076, n17077, n17078,
    n17079, n17080, n17081, n17082, n17083, n17084,
    n17085, n17086, n17087, n17088, n17089, n17090,
    n17091, n17092, n17093, n17094, n17095, n17096,
    n17097, n17098, n17099, n17100, n17101, n17102,
    n17103, n17104, n17105, n17106, n17107, n17108,
    n17109, n17110, n17111, n17112, n17113, n17114,
    n17115, n17116, n17117, n17118, n17119, n17120,
    n17121, n17122, n17123, n17124, n17125, n17126,
    n17127, n17128, n17129, n17130, n17131, n17132,
    n17133, n17134, n17135, n17136, n17137, n17138,
    n17139, n17140, n17141, n17142, n17143, n17144,
    n17145, n17146, n17147, n17148, n17149, n17150,
    n17151, n17152, n17153, n17154, n17155, n17156,
    n17157, n17158, n17159, n17160, n17161, n17162,
    n17163, n17164, n17165, n17166, n17167, n17168,
    n17169, n17170, n17171, n17172, n17173, n17174,
    n17175, n17176, n17177, n17178, n17179, n17180,
    n17181, n17182, n17183, n17184, n17185, n17186,
    n17187, n17188, n17189, n17190, n17191, n17192,
    n17193, n17194, n17195, n17196, n17197, n17198,
    n17199, n17200, n17201, n17202, n17203, n17204,
    n17205, n17206, n17207, n17208, n17209, n17210,
    n17211, n17212, n17213, n17214, n17215, n17216,
    n17217, n17218, n17219, n17220, n17221, n17222,
    n17223, n17224, n17225, n17226, n17227, n17228,
    n17229, n17230, n17231, n17232, n17233, n17234,
    n17235, n17236, n17237, n17238, n17239, n17240,
    n17241, n17242, n17243, n17244, n17245, n17246,
    n17247, n17248, n17249, n17250, n17251, n17252,
    n17253, n17254, n17255, n17256, n17257, n17258,
    n17259, n17260, n17261, n17262, n17263, n17264,
    n17265, n17266, n17267, n17268, n17269, n17270,
    n17271, n17272, n17273, n17274, n17275, n17276,
    n17277, n17278, n17279, n17280, n17281, n17282,
    n17283, n17284, n17285, n17286, n17287, n17288,
    n17289, n17290, n17291, n17292, n17293, n17294,
    n17295, n17296, n17297, n17298, n17299, n17300,
    n17301, n17302, n17303, n17304, n17305, n17306,
    n17307, n17308, n17309, n17310, n17311, n17312,
    n17313, n17314, n17315, n17316, n17317, n17318,
    n17319, n17320, n17321, n17322, n17323, n17324,
    n17325, n17326, n17327, n17328, n17329, n17330,
    n17331, n17332, n17333, n17334, n17335, n17336,
    n17337, n17338, n17339, n17340, n17341, n17342,
    n17343, n17344, n17345, n17346, n17347, n17348,
    n17349, n17350, n17351, n17352, n17353, n17354,
    n17355, n17356, n17357, n17358, n17359, n17360,
    n17361, n17362, n17363, n17364, n17365, n17366,
    n17367, n17368, n17369, n17370, n17371, n17372,
    n17373, n17374, n17375, n17376, n17377, n17378,
    n17379, n17380, n17381, n17382, n17383, n17384,
    n17385, n17386, n17387, n17388, n17389, n17390,
    n17391, n17392, n17393, n17394, n17395, n17396,
    n17397, n17398, n17399, n17400, n17401, n17402,
    n17403, n17404, n17405, n17406, n17407, n17408,
    n17409, n17410, n17411, n17412, n17413, n17414,
    n17415, n17416, n17417, n17418, n17419, n17420,
    n17421, n17422, n17423, n17424, n17425, n17426,
    n17427, n17428, n17429, n17430, n17431, n17432,
    n17433, n17434, n17435, n17436, n17437, n17438,
    n17439, n17440, n17441, n17442, n17443, n17444,
    n17445, n17446, n17447, n17448, n17449, n17450,
    n17451, n17452, n17453, n17454, n17455, n17456,
    n17457, n17458, n17459, n17460, n17461, n17462,
    n17463, n17464, n17465, n17466, n17467, n17468,
    n17469, n17470, n17471, n17472, n17473, n17474,
    n17475, n17476, n17477, n17478, n17479, n17480,
    n17481, n17482, n17483, n17484, n17485, n17486,
    n17487, n17488, n17489, n17490, n17491, n17492,
    n17493, n17494, n17495, n17496, n17497, n17498,
    n17499, n17500, n17501, n17502, n17503, n17504,
    n17505, n17506, n17507, n17508, n17509, n17510,
    n17511, n17512, n17513, n17514, n17515, n17516,
    n17517, n17518, n17519, n17520, n17521, n17522,
    n17523, n17524, n17525, n17526, n17527, n17528,
    n17529, n17530, n17531, n17532, n17533, n17534,
    n17535, n17536, n17537, n17538, n17539, n17540,
    n17541, n17542, n17543, n17544, n17545, n17546,
    n17547, n17548, n17549, n17550, n17551, n17552,
    n17553, n17554, n17555, n17556, n17557, n17558,
    n17559, n17560, n17561, n17562, n17563, n17564,
    n17565, n17566, n17567, n17568, n17569, n17570,
    n17571, n17572, n17573, n17574, n17575, n17576,
    n17577, n17578, n17579, n17580, n17581, n17582,
    n17583, n17584, n17585, n17586, n17587, n17588,
    n17589, n17590, n17591, n17592, n17593, n17594,
    n17595, n17596, n17597, n17598, n17599, n17600,
    n17601, n17602, n17603, n17604, n17605, n17606,
    n17607, n17608, n17609, n17610, n17611, n17612,
    n17613, n17614, n17615, n17616, n17617, n17618,
    n17619, n17620, n17621, n17622, n17623, n17624,
    n17625, n17626, n17627, n17628, n17629, n17630,
    n17631, n17632, n17633, n17634, n17635, n17636,
    n17637, n17638, n17639, n17640, n17641, n17642,
    n17643, n17644, n17645, n17646, n17647, n17648,
    n17649, n17650, n17651, n17652, n17653, n17654,
    n17655, n17656, n17657, n17658, n17659, n17660,
    n17661, n17662, n17663, n17664, n17665, n17666,
    n17667, n17668, n17669, n17670, n17671, n17672,
    n17673, n17674, n17675, n17676, n17677, n17678,
    n17679, n17680, n17681, n17682, n17683, n17684,
    n17685, n17686, n17687, n17688, n17689, n17690,
    n17691, n17692, n17693, n17694, n17695, n17696,
    n17697, n17698, n17699, n17700, n17701, n17702,
    n17703, n17704, n17705, n17706, n17707, n17708,
    n17709, n17710, n17711, n17712, n17713, n17714,
    n17715, n17716, n17717, n17718, n17719, n17720,
    n17721, n17722, n17723, n17724, n17725, n17726,
    n17727, n17728, n17729, n17730, n17731, n17732,
    n17733, n17734, n17735, n17736, n17737, n17738,
    n17739, n17740, n17741, n17742, n17743, n17744,
    n17745, n17746, n17747, n17748, n17749, n17750,
    n17751, n17752, n17753, n17754, n17755, n17756,
    n17757, n17758, n17759, n17760, n17761, n17762,
    n17763, n17764, n17765, n17766, n17767, n17768,
    n17769, n17770, n17771, n17772, n17773, n17774,
    n17775, n17776, n17777, n17778, n17779, n17780,
    n17781, n17782, n17783, n17784, n17785, n17786,
    n17787, n17788, n17789, n17790, n17791, n17792,
    n17793, n17794, n17795, n17796, n17797, n17798,
    n17799, n17800, n17801, n17802, n17803, n17804,
    n17805, n17806, n17807, n17808, n17809, n17810,
    n17811, n17812, n17813, n17814, n17815, n17816,
    n17817, n17818, n17819, n17820, n17821, n17822,
    n17823, n17824, n17825, n17826, n17827, n17828,
    n17829, n17830, n17831, n17832, n17833, n17834,
    n17835, n17836, n17837, n17838, n17839, n17840,
    n17841, n17842, n17843, n17844, n17845, n17846,
    n17847, n17848, n17849, n17850, n17851, n17852,
    n17853, n17854, n17855, n17856, n17857, n17858,
    n17859, n17860, n17861, n17862, n17863, n17864,
    n17865, n17866, n17867, n17868, n17869, n17870,
    n17871, n17872, n17873, n17874, n17875, n17876,
    n17877, n17878, n17879, n17880, n17881, n17882,
    n17883, n17884, n17885, n17886, n17887, n17888,
    n17889, n17890, n17891, n17892, n17893, n17894,
    n17895, n17896, n17897, n17898, n17899, n17900,
    n17901, n17902, n17903, n17904, n17905, n17906,
    n17907, n17908, n17909, n17910, n17911, n17912,
    n17913, n17914, n17915, n17916, n17917, n17918,
    n17919, n17920, n17921, n17922, n17923, n17924,
    n17925, n17926, n17927, n17928, n17929, n17930,
    n17931, n17932, n17933, n17934, n17935, n17936,
    n17937, n17938, n17939, n17940, n17941, n17942,
    n17943, n17944, n17945, n17946, n17947, n17948,
    n17949, n17950, n17951, n17952, n17953, n17954,
    n17955, n17956, n17957, n17958, n17959, n17960,
    n17961, n17962, n17963, n17964, n17965, n17966,
    n17967, n17968, n17969, n17970, n17971, n17972,
    n17973, n17974, n17975, n17976, n17977, n17978,
    n17979, n17980, n17981, n17982, n17983, n17984,
    n17985, n17986, n17987, n17988, n17989, n17990,
    n17991, n17992, n17993, n17994, n17995, n17996,
    n17997, n17998, n17999, n18000, n18001, n18002,
    n18003, n18004, n18005, n18006, n18007, n18008,
    n18009, n18010, n18011, n18012, n18013, n18014,
    n18015, n18016, n18017, n18018, n18019, n18020,
    n18021, n18022, n18023, n18024, n18025, n18026,
    n18027, n18028, n18029, n18030, n18031, n18032,
    n18033, n18034, n18035, n18036, n18037, n18038,
    n18039, n18040, n18041, n18042, n18043, n18044,
    n18045, n18046, n18047, n18048, n18049, n18050,
    n18051, n18052, n18053, n18054, n18055, n18056,
    n18057, n18058, n18059, n18060, n18061, n18062,
    n18063, n18064, n18065, n18066, n18067, n18068,
    n18069, n18070, n18071, n18072, n18073, n18074,
    n18075, n18076, n18077, n18078, n18079, n18080,
    n18081, n18082, n18083, n18084, n18085, n18086,
    n18087, n18088, n18089, n18090, n18091, n18092,
    n18093, n18094, n18095, n18096, n18097, n18098,
    n18099, n18100, n18101, n18102, n18103, n18104,
    n18105, n18106, n18107, n18108, n18109, n18110,
    n18111, n18112, n18113, n18114, n18115, n18116,
    n18117, n18118, n18119, n18120, n18121, n18122,
    n18123, n18124, n18125, n18126, n18127, n18128,
    n18129, n18130, n18131, n18132, n18133, n18134,
    n18135, n18136, n18137, n18138, n18139, n18140,
    n18141, n18142, n18143, n18144, n18145, n18146,
    n18147, n18148, n18149, n18150, n18151, n18152,
    n18153, n18154, n18155, n18156, n18157, n18158,
    n18159, n18160, n18161, n18162, n18163, n18164,
    n18165, n18166, n18167, n18168, n18169, n18170,
    n18171, n18172, n18173, n18174, n18175, n18176,
    n18177, n18178, n18179, n18180, n18181, n18182,
    n18183, n18184, n18185, n18186, n18187, n18188,
    n18189, n18190, n18191, n18192, n18193, n18194,
    n18195, n18196, n18197, n18198, n18199, n18200,
    n18201, n18202, n18203, n18204, n18205, n18206,
    n18207, n18208, n18209, n18210, n18211, n18212,
    n18213, n18214, n18215, n18216, n18217, n18218,
    n18219, n18220, n18221, n18222, n18223, n18224,
    n18225, n18226, n18227, n18228, n18229, n18230,
    n18231, n18232, n18233, n18234, n18235, n18236,
    n18237, n18238, n18239, n18240, n18241, n18242,
    n18243, n18244, n18245, n18246, n18247, n18248,
    n18249, n18250, n18251, n18252, n18253, n18254,
    n18255, n18256, n18257, n18258, n18259, n18260,
    n18261, n18262, n18263, n18264, n18265, n18266,
    n18267, n18268, n18269, n18270, n18271, n18272,
    n18273, n18274, n18275, n18276, n18277, n18278,
    n18279, n18280, n18281, n18282, n18283, n18284,
    n18285, n18286, n18287, n18288, n18289, n18290,
    n18291, n18292, n18293, n18294, n18295, n18296,
    n18297, n18298, n18299, n18300, n18301, n18302,
    n18303, n18304, n18305, n18306, n18307, n18308,
    n18309, n18310, n18311, n18312, n18313, n18314,
    n18315, n18316, n18317, n18318, n18319, n18320,
    n18321, n18322, n18323, n18324, n18325, n18326,
    n18327, n18328, n18329, n18330, n18331, n18332,
    n18333, n18334, n18335, n18336, n18337, n18338,
    n18339, n18340, n18341, n18342, n18343, n18344,
    n18345, n18346, n18347, n18348, n18349, n18350,
    n18351, n18352, n18353, n18354, n18355, n18356,
    n18357, n18358, n18359, n18360, n18361, n18362,
    n18363, n18364, n18365, n18366, n18367, n18368,
    n18369, n18370, n18371, n18372, n18373, n18374,
    n18375, n18376, n18377, n18378, n18379, n18380,
    n18381, n18382, n18383, n18384, n18385, n18386,
    n18387, n18388, n18389, n18390, n18391, n18392,
    n18393, n18394, n18395, n18396, n18397, n18398,
    n18399, n18400, n18401, n18402, n18403, n18404,
    n18405, n18406, n18407, n18408, n18409, n18410,
    n18411, n18412, n18413, n18414, n18415, n18416,
    n18417, n18418, n18419, n18420, n18421, n18422,
    n18423, n18424, n18425, n18426, n18427, n18428,
    n18429, n18430, n18431, n18432, n18433, n18434,
    n18435, n18436, n18437, n18438, n18439, n18440,
    n18441, n18442, n18443, n18444, n18445, n18446,
    n18447, n18448, n18449, n18450, n18451, n18452,
    n18453, n18454, n18455, n18456, n18457, n18458,
    n18459, n18460, n18461, n18462, n18463, n18464,
    n18465, n18466, n18467, n18468, n18469, n18470,
    n18471, n18472, n18473, n18474, n18475, n18476,
    n18477, n18478, n18479, n18480, n18481, n18482,
    n18483, n18484, n18485, n18486, n18487, n18488,
    n18489, n18490, n18491, n18492, n18493, n18494,
    n18495, n18496, n18497, n18498, n18499, n18500,
    n18501, n18502, n18503, n18504, n18505, n18506,
    n18507, n18508, n18509, n18510, n18511, n18512,
    n18513, n18514, n18515, n18516, n18517, n18518,
    n18519, n18520, n18521, n18522, n18523, n18524,
    n18525, n18526, n18527, n18528, n18529, n18530,
    n18531, n18532, n18533, n18534, n18535, n18536,
    n18537, n18538, n18539, n18540, n18541, n18542,
    n18543, n18544, n18545, n18546, n18547, n18548,
    n18549, n18550, n18551, n18552, n18553, n18554,
    n18555, n18556, n18557, n18558, n18559, n18560,
    n18561, n18562, n18563, n18564, n18565, n18566,
    n18567, n18568, n18569, n18570, n18571, n18572,
    n18573, n18574, n18575, n18576, n18577, n18578,
    n18579, n18580, n18581, n18582, n18583, n18584,
    n18585, n18586, n18587, n18588, n18589, n18590,
    n18591, n18592, n18593, n18594, n18595, n18596,
    n18597, n18598, n18599, n18600, n18601, n18602,
    n18603, n18604, n18605, n18606, n18607, n18608,
    n18609, n18610, n18611, n18612, n18613, n18614,
    n18615, n18616, n18617, n18618, n18619, n18620,
    n18621, n18622, n18623, n18624, n18625, n18626,
    n18627, n18628, n18629, n18630, n18631, n18632,
    n18633, n18634, n18635, n18636, n18637, n18638,
    n18639, n18640, n18641, n18642, n18643, n18644,
    n18645, n18646, n18647, n18648, n18649, n18650,
    n18651, n18652, n18653, n18654, n18655, n18656,
    n18657, n18658, n18659, n18660, n18661, n18662,
    n18663, n18664, n18665, n18666, n18667, n18668,
    n18669, n18670, n18671, n18672, n18673, n18674,
    n18675, n18676, n18677, n18678, n18679, n18680,
    n18681, n18682, n18683, n18684, n18685, n18686,
    n18687, n18688, n18689, n18690, n18691, n18692,
    n18693, n18694, n18695, n18696, n18697, n18698,
    n18699, n18700, n18701, n18702, n18703, n18704,
    n18705, n18706, n18707, n18708, n18709, n18710,
    n18711, n18712, n18713, n18714, n18715, n18716,
    n18717, n18718, n18719, n18720, n18721, n18722,
    n18723, n18724, n18725, n18726, n18727, n18728,
    n18729, n18730, n18731, n18732, n18733, n18734,
    n18735, n18736, n18737, n18738, n18739, n18740,
    n18741, n18742, n18743, n18744, n18745, n18746,
    n18747, n18748, n18749, n18750, n18751, n18752,
    n18753, n18754, n18755, n18756, n18757, n18758,
    n18759, n18760, n18761, n18762, n18763, n18764,
    n18765, n18766, n18767, n18768, n18769, n18770,
    n18771, n18772, n18773, n18774, n18775, n18776,
    n18777, n18778, n18779, n18780, n18781, n18782,
    n18783, n18784, n18785, n18786, n18787, n18788,
    n18789, n18790, n18791, n18792, n18793, n18794,
    n18795, n18796, n18797, n18798, n18799, n18800,
    n18801, n18802, n18803, n18804, n18805, n18806,
    n18807, n18808, n18809, n18810, n18811, n18812,
    n18813, n18814, n18815, n18816, n18817, n18818,
    n18819, n18820, n18821, n18822, n18823, n18824,
    n18825, n18826, n18827, n18828, n18829, n18830,
    n18831, n18832, n18833, n18834, n18835, n18836,
    n18837, n18838, n18839, n18840, n18841, n18842,
    n18843, n18844, n18845, n18846, n18847, n18848,
    n18849, n18850, n18851, n18852, n18853, n18854,
    n18855, n18856, n18857, n18858, n18859, n18860,
    n18861, n18862, n18863, n18864, n18865, n18866,
    n18867, n18868, n18869, n18870, n18871, n18872,
    n18873, n18874, n18875, n18876, n18877, n18878,
    n18879, n18880, n18881, n18882, n18883, n18884,
    n18885, n18886, n18887, n18888, n18889, n18890,
    n18891, n18892, n18893, n18894, n18895, n18896,
    n18897, n18898, n18899, n18900, n18901, n18902,
    n18903, n18904, n18905, n18906, n18907, n18908,
    n18909, n18910, n18911, n18912, n18913, n18914,
    n18915, n18916, n18917, n18918, n18919, n18920,
    n18921, n18922, n18923, n18924, n18925, n18926,
    n18927, n18928, n18929, n18930, n18931, n18932,
    n18933, n18934, n18935, n18936, n18937, n18938,
    n18939, n18940, n18941, n18942, n18943, n18944,
    n18945, n18946, n18947, n18948, n18949, n18950,
    n18951, n18952, n18953, n18954, n18955, n18956,
    n18957, n18958, n18959, n18960, n18961, n18962,
    n18963, n18964, n18965, n18966, n18967, n18968,
    n18969, n18970, n18971, n18972, n18973, n18974,
    n18975, n18976, n18977, n18978, n18979, n18980,
    n18981, n18982, n18983, n18984, n18985, n18986,
    n18987, n18988, n18989, n18990, n18991, n18992,
    n18993, n18994, n18995, n18996, n18997, n18998,
    n18999, n19000, n19001, n19002, n19003, n19004,
    n19005, n19006, n19007, n19008, n19009, n19010,
    n19011, n19012, n19013, n19014, n19015, n19016,
    n19017, n19018, n19019, n19020, n19021, n19022,
    n19023, n19024, n19025, n19026, n19027, n19028,
    n19029, n19030, n19031, n19032, n19033, n19034,
    n19035, n19036, n19037, n19038, n19039, n19040,
    n19041, n19042, n19043, n19044, n19045, n19046,
    n19047, n19048, n19049, n19050, n19051, n19052,
    n19053, n19054, n19055, n19056, n19057, n19058,
    n19059, n19060, n19061, n19062, n19063, n19064,
    n19065, n19066, n19067, n19068, n19069, n19070,
    n19071, n19072, n19073, n19074, n19075, n19076,
    n19077, n19078, n19079, n19080, n19081, n19082,
    n19083, n19084, n19085, n19086, n19087, n19088,
    n19089, n19090, n19091, n19092, n19093, n19094,
    n19095, n19096, n19097, n19098, n19099, n19100,
    n19101, n19102, n19103, n19104, n19105, n19106,
    n19107, n19108, n19109, n19110, n19111, n19112,
    n19113, n19114, n19115, n19116, n19117, n19118,
    n19119, n19120, n19121, n19122, n19123, n19124,
    n19125, n19126, n19127, n19128, n19129, n19130,
    n19131, n19132, n19133, n19134, n19135, n19136,
    n19137, n19138, n19139, n19140, n19141, n19142,
    n19143, n19144, n19145, n19146, n19147, n19148,
    n19149, n19150, n19151, n19152, n19153, n19154,
    n19155, n19156, n19157, n19158, n19159, n19160,
    n19161, n19162, n19163, n19164, n19165, n19166,
    n19167, n19168, n19169, n19170, n19171, n19172,
    n19173, n19174, n19175, n19176, n19177, n19178,
    n19179, n19180, n19181, n19182, n19183, n19184,
    n19185, n19186, n19187, n19188, n19189, n19190,
    n19191, n19192, n19193, n19194, n19195, n19196,
    n19197, n19198, n19199, n19200, n19201, n19202,
    n19203, n19204, n19205, n19206, n19207, n19208,
    n19209, n19210, n19211, n19212, n19213, n19214,
    n19215, n19216, n19217, n19218, n19219, n19220,
    n19221, n19222, n19223, n19224, n19225, n19226,
    n19227, n19228, n19229, n19230, n19231, n19232,
    n19233, n19234, n19235, n19236, n19237, n19238,
    n19239, n19240, n19241, n19242, n19243, n19244,
    n19245, n19246, n19247, n19248, n19249, n19250,
    n19251, n19252, n19253, n19254, n19255, n19256,
    n19257, n19258, n19259, n19260, n19261, n19262,
    n19263, n19264, n19265, n19266, n19267, n19268,
    n19269, n19270, n19271, n19272, n19273, n19274,
    n19275, n19276, n19277, n19278, n19279, n19280,
    n19281, n19282, n19283, n19284, n19285, n19286,
    n19287, n19288, n19289, n19290, n19291, n19292,
    n19293, n19294, n19295, n19296, n19297, n19298,
    n19299, n19300, n19301, n19302, n19303, n19304,
    n19305, n19306, n19307, n19308, n19309, n19310,
    n19311, n19312, n19313, n19314, n19315, n19316,
    n19317, n19318, n19319, n19320, n19321, n19322,
    n19323, n19324, n19325, n19326, n19327, n19328,
    n19329, n19330, n19331, n19332, n19333, n19334,
    n19335, n19336, n19337, n19338, n19339, n19340,
    n19341, n19342, n19343, n19344, n19345, n19346,
    n19347, n19348, n19349, n19350, n19351, n19352,
    n19353, n19354, n19355, n19356, n19357, n19358,
    n19359, n19360, n19361, n19362, n19363, n19364,
    n19365, n19366, n19367, n19368, n19369, n19370,
    n19371, n19372, n19373, n19374, n19375, n19376,
    n19377, n19378, n19379, n19380, n19381, n19382,
    n19383, n19384, n19385, n19386, n19387, n19388,
    n19389, n19390, n19391, n19392, n19393, n19394,
    n19395, n19396, n19397, n19398, n19399, n19400,
    n19401, n19402, n19403, n19404, n19405, n19406,
    n19407, n19408, n19409, n19410, n19411, n19412,
    n19413, n19414, n19415, n19416, n19417, n19418,
    n19419, n19420, n19421, n19422, n19423, n19424,
    n19425, n19426, n19427, n19428, n19429, n19430,
    n19431, n19432, n19433, n19434, n19435, n19436,
    n19437, n19438, n19439, n19440, n19441, n19442,
    n19443, n19444, n19445, n19446, n19447, n19448,
    n19449, n19450, n19451, n19452, n19453, n19454,
    n19455, n19456, n19457, n19458, n19459, n19460,
    n19461, n19462, n19463, n19464, n19465, n19466,
    n19467, n19468, n19469, n19470, n19471, n19472,
    n19473, n19474, n19475, n19476, n19477, n19478,
    n19479, n19480, n19481, n19482, n19483, n19484,
    n19485, n19486, n19487, n19488, n19489, n19490,
    n19491, n19492, n19493, n19494, n19495, n19496,
    n19497, n19498, n19499, n19500, n19501, n19502,
    n19503, n19504, n19505, n19506, n19507, n19508,
    n19509, n19510, n19511, n19512, n19513, n19514,
    n19515, n19516, n19517, n19518, n19519, n19520,
    n19521, n19522, n19523, n19524, n19525, n19526,
    n19527, n19528, n19529, n19530, n19531, n19532,
    n19533, n19534, n19535, n19536, n19537, n19538,
    n19539, n19540, n19541, n19542, n19543, n19544,
    n19545, n19546, n19547, n19548, n19549, n19550,
    n19551, n19552, n19553, n19554, n19555, n19556,
    n19557, n19558, n19559, n19560, n19561, n19562,
    n19563, n19564, n19565, n19566, n19567, n19568,
    n19569, n19570, n19571, n19572, n19573, n19574,
    n19575, n19576, n19577, n19578, n19579, n19580,
    n19581, n19582, n19583, n19584, n19585, n19586,
    n19587, n19588, n19589, n19590, n19591, n19592,
    n19593, n19594, n19595, n19596, n19597, n19598,
    n19599, n19600, n19601, n19602, n19603, n19604,
    n19605, n19606, n19607, n19608, n19609, n19610,
    n19611, n19612, n19613, n19614, n19615, n19616,
    n19617, n19618, n19619, n19620, n19621, n19622,
    n19623, n19624, n19625, n19626, n19627, n19628,
    n19629, n19630, n19631, n19632, n19633, n19634,
    n19635, n19636, n19637, n19638, n19639, n19640,
    n19641, n19642, n19643, n19644, n19645, n19646,
    n19647, n19648, n19649, n19650, n19651, n19652,
    n19653, n19654, n19655, n19656, n19657, n19658,
    n19659, n19660, n19661, n19662, n19663, n19664,
    n19665, n19666, n19667, n19668, n19669, n19670,
    n19671, n19672, n19673, n19674, n19675, n19676,
    n19677, n19678, n19679, n19680, n19681, n19682,
    n19683, n19684, n19685, n19686, n19687, n19688,
    n19689, n19690, n19691, n19692, n19693, n19694,
    n19695, n19696, n19697, n19698, n19699, n19700,
    n19701, n19702, n19703, n19704, n19705, n19706,
    n19707, n19708, n19709, n19710, n19711, n19712,
    n19713, n19714, n19715, n19716, n19717, n19718,
    n19719, n19720, n19721, n19722, n19723, n19724,
    n19725, n19726, n19727, n19728, n19729, n19730,
    n19731, n19732, n19733, n19734, n19735, n19736,
    n19737, n19738, n19739, n19740, n19741, n19742,
    n19743, n19744, n19745, n19746, n19747, n19748,
    n19749, n19750, n19751, n19752, n19753, n19754,
    n19755, n19756, n19757, n19758, n19759, n19760,
    n19761, n19762, n19763, n19764, n19765, n19766,
    n19767, n19768, n19769, n19770, n19771, n19772,
    n19773, n19774, n19775, n19776, n19777, n19778,
    n19779, n19780, n19781, n19782, n19783, n19784,
    n19785, n19786, n19787, n19788, n19789, n19790,
    n19791, n19792, n19793, n19794, n19795, n19796,
    n19797, n19798, n19799, n19800, n19801, n19802,
    n19803, n19804, n19805, n19806, n19807, n19808,
    n19809, n19810, n19811, n19812, n19813, n19814,
    n19815, n19816, n19817, n19818, n19819, n19820,
    n19821, n19822, n19823, n19824, n19825, n19826,
    n19827, n19828, n19829, n19830, n19831, n19832,
    n19833, n19834, n19835, n19836, n19837, n19838,
    n19839, n19840, n19841, n19842, n19843, n19844,
    n19845, n19846, n19847, n19848, n19849, n19850,
    n19851, n19852, n19853, n19854, n19855, n19856,
    n19857, n19858, n19859, n19860, n19861, n19862,
    n19863, n19864, n19865, n19866, n19867, n19868,
    n19869, n19870, n19871, n19872, n19873, n19874,
    n19875, n19876, n19877, n19878, n19879, n19880,
    n19881, n19882, n19883, n19884, n19885, n19886,
    n19887, n19888, n19889, n19890, n19891, n19892,
    n19893, n19894, n19895, n19896, n19897, n19898,
    n19899, n19900, n19901, n19902, n19903, n19904,
    n19905, n19906, n19907, n19908, n19909, n19910,
    n19911, n19912, n19913, n19914, n19915, n19916,
    n19917, n19918, n19919, n19920, n19921, n19922,
    n19923, n19924, n19925, n19926, n19927, n19928,
    n19929, n19930, n19931, n19932, n19933, n19934,
    n19935, n19936, n19937, n19938, n19939, n19940,
    n19941, n19942, n19943, n19944, n19945, n19946,
    n19947, n19948, n19949, n19950, n19951, n19952,
    n19953, n19954, n19955, n19956, n19957, n19958,
    n19959, n19960, n19961, n19962, n19963, n19964,
    n19965, n19966, n19967, n19968, n19969, n19970,
    n19971, n19972, n19973, n19974, n19975, n19976,
    n19977, n19978, n19979, n19980, n19981, n19982,
    n19983, n19984, n19985, n19986, n19987, n19988,
    n19989, n19990, n19991, n19992, n19993, n19994,
    n19995, n19996, n19997, n19998, n19999, n20000,
    n20001, n20002, n20003, n20004, n20005, n20006,
    n20007, n20008, n20009, n20010, n20011, n20012,
    n20013, n20014, n20015, n20016, n20017, n20018,
    n20019, n20020, n20021, n20022, n20023, n20024,
    n20025, n20026, n20027, n20028, n20029, n20030,
    n20031, n20032, n20033, n20034, n20035, n20036,
    n20037, n20038, n20039, n20040, n20041, n20042,
    n20043, n20044, n20045, n20046, n20047, n20048,
    n20049, n20050, n20051, n20052, n20053, n20054,
    n20055, n20056, n20057, n20058, n20059, n20060,
    n20061, n20062, n20063, n20064, n20065, n20066,
    n20067, n20068, n20069, n20070, n20071, n20072,
    n20073, n20074, n20075, n20076, n20077, n20078,
    n20079, n20080, n20081, n20082, n20083, n20084,
    n20085, n20086, n20087, n20088, n20089, n20090,
    n20091, n20092, n20093, n20094, n20095, n20096,
    n20097, n20098, n20099, n20100, n20101, n20102,
    n20103, n20104, n20105, n20106, n20107, n20108,
    n20109, n20110, n20111, n20112, n20113, n20114,
    n20115, n20116, n20117, n20118, n20119, n20120,
    n20121, n20122, n20123, n20124, n20125, n20126,
    n20127, n20128, n20129, n20130, n20131, n20132,
    n20133, n20134, n20135, n20136, n20137, n20138,
    n20139, n20140, n20141, n20142, n20143, n20144,
    n20145, n20146, n20147, n20148, n20149, n20150,
    n20151, n20152, n20153, n20154, n20155, n20156,
    n20157, n20158, n20159, n20160, n20161, n20162,
    n20163, n20164, n20165, n20166, n20167, n20168,
    n20169, n20170, n20171, n20172, n20173, n20174,
    n20175, n20176, n20177, n20178, n20179, n20180,
    n20181, n20182, n20183, n20184, n20185, n20186,
    n20187, n20188, n20189, n20190, n20191, n20192,
    n20193, n20194, n20195, n20196, n20197, n20198,
    n20199, n20200, n20201, n20202, n20203, n20204,
    n20205, n20206, n20207, n20208, n20209, n20210,
    n20211, n20212, n20213, n20214, n20215, n20216,
    n20217, n20218, n20219, n20220, n20221, n20222,
    n20223, n20224, n20225, n20226, n20227, n20228,
    n20229, n20230, n20231, n20232, n20233, n20234,
    n20235, n20236, n20237, n20238, n20239, n20240,
    n20241, n20242, n20243, n20244, n20245, n20246,
    n20247, n20248, n20249, n20250, n20251, n20252,
    n20253, n20254, n20255, n20256, n20257, n20258,
    n20259, n20260, n20261, n20262, n20263, n20264,
    n20265, n20266, n20267, n20268, n20269, n20270,
    n20271, n20272, n20273, n20274, n20275, n20276,
    n20277, n20278, n20279, n20280, n20281, n20282,
    n20283, n20284, n20285, n20286, n20287, n20288,
    n20289, n20290, n20291, n20292, n20293, n20294,
    n20295, n20296, n20297, n20298, n20299, n20300,
    n20301, n20302, n20303, n20304, n20305, n20306,
    n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318,
    n20319, n20320, n20321, n20322, n20323, n20324,
    n20325, n20326, n20327, n20328, n20329, n20330,
    n20331, n20332, n20333, n20334, n20335, n20336,
    n20337, n20338, n20339, n20340, n20341, n20342,
    n20343, n20344, n20345, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354,
    n20355, n20356, n20357, n20358, n20359, n20360,
    n20361, n20362, n20363, n20364, n20365, n20366,
    n20367, n20368, n20369, n20370, n20371, n20372,
    n20373, n20374, n20375, n20376, n20377, n20378,
    n20379, n20380, n20381, n20382, n20383, n20384,
    n20385, n20386, n20387, n20388, n20389, n20390,
    n20391, n20392, n20393, n20394, n20395, n20396,
    n20397, n20398, n20399, n20400, n20401, n20402,
    n20403, n20404, n20405, n20406, n20407, n20408,
    n20409, n20410, n20411, n20412, n20413, n20414,
    n20415, n20416, n20417, n20418, n20419, n20420,
    n20421, n20422, n20423, n20424, n20425, n20426,
    n20427, n20428, n20429, n20430, n20431, n20432,
    n20433, n20434, n20435, n20436, n20437, n20438,
    n20439, n20440, n20441, n20442, n20443, n20444,
    n20445, n20446, n20447, n20448, n20449, n20450,
    n20451, n20452, n20453, n20454, n20455, n20456,
    n20457, n20458, n20459, n20460, n20461, n20462,
    n20463, n20464, n20465, n20466, n20467, n20468,
    n20469, n20470, n20471, n20472, n20473, n20474,
    n20475, n20476, n20477, n20478, n20479, n20480,
    n20481, n20482, n20483, n20484, n20485, n20486,
    n20487, n20488, n20489, n20490, n20491, n20492,
    n20493, n20494, n20495, n20496, n20497, n20498,
    n20499, n20500, n20501, n20502, n20503, n20504,
    n20505, n20506, n20507, n20508, n20509, n20510,
    n20511, n20512, n20513, n20514, n20515, n20516,
    n20517, n20518, n20519, n20520, n20521, n20522,
    n20523, n20524, n20525, n20526, n20527, n20528,
    n20529, n20530, n20531, n20532, n20533, n20534,
    n20535, n20536, n20537, n20538, n20539, n20540,
    n20541, n20542, n20543, n20544, n20545, n20546,
    n20547, n20548, n20549, n20550, n20551, n20552,
    n20553, n20554, n20555, n20556, n20557, n20558,
    n20559, n20560, n20561, n20562, n20563, n20564,
    n20565, n20566, n20567, n20568, n20569, n20570,
    n20571, n20572, n20573, n20574, n20575, n20576,
    n20577, n20578, n20579, n20580, n20581, n20582,
    n20583, n20584, n20585, n20586, n20587, n20588,
    n20589, n20590, n20591, n20592, n20593, n20594,
    n20595, n20596, n20597, n20598, n20599, n20600,
    n20601, n20602, n20603, n20604, n20605, n20606,
    n20607, n20608, n20609, n20610, n20611, n20612,
    n20613, n20614, n20615, n20616, n20617, n20618,
    n20619, n20620, n20621, n20622, n20623, n20624,
    n20625, n20626, n20627, n20628, n20629, n20630,
    n20631, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20645, n20646, n20647, n20648,
    n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660,
    n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20675, n20676, n20677, n20678,
    n20679, n20680, n20681, n20682, n20683, n20684,
    n20685, n20686, n20687, n20688, n20689, n20690,
    n20691, n20692, n20693, n20694, n20695, n20696,
    n20697, n20698, n20699, n20700, n20701, n20702,
    n20703, n20704, n20705, n20706, n20707, n20708,
    n20709, n20710, n20711, n20712, n20713, n20714,
    n20715, n20716, n20717, n20718, n20719, n20720,
    n20721, n20722, n20723, n20724, n20725, n20726,
    n20727, n20728, n20729, n20730, n20731, n20732,
    n20733, n20734, n20735, n20736, n20737, n20738,
    n20739, n20740, n20741, n20742, n20743, n20744,
    n20745, n20746, n20747, n20748, n20749, n20750,
    n20751, n20752, n20753, n20754, n20755, n20756,
    n20757, n20758, n20759, n20760, n20761, n20762,
    n20763, n20764, n20765, n20766, n20767, n20768,
    n20769, n20770, n20771, n20772, n20773, n20774,
    n20775, n20776, n20777, n20778, n20779, n20780,
    n20781, n20782, n20783, n20784, n20785, n20786,
    n20787, n20788, n20789, n20790, n20791, n20792,
    n20793, n20794, n20795, n20796, n20797, n20798,
    n20799, n20800, n20801, n20802, n20803, n20804,
    n20805, n20806, n20807, n20808, n20809, n20810,
    n20811, n20812, n20813, n20814, n20815, n20816,
    n20817, n20818, n20819, n20820, n20821, n20822,
    n20823, n20824, n20825, n20826, n20827, n20828,
    n20829, n20830, n20831, n20832, n20833, n20834,
    n20835, n20836, n20837, n20838, n20839, n20840,
    n20841, n20842, n20843, n20844, n20845, n20846,
    n20847, n20848, n20849, n20850, n20851, n20852,
    n20853, n20854, n20855, n20856, n20857, n20858,
    n20859, n20860, n20861, n20862, n20863, n20864,
    n20865, n20866, n20867, n20868, n20869, n20870,
    n20871, n20872, n20873, n20874, n20875, n20876,
    n20877, n20878, n20879, n20880, n20881, n20882,
    n20883, n20884, n20885, n20886, n20887, n20888,
    n20889, n20890, n20891, n20892, n20893, n20894,
    n20895, n20896, n20897, n20898, n20899, n20900,
    n20901, n20902, n20903, n20904, n20905, n20906,
    n20907, n20908, n20909, n20910, n20911, n20912,
    n20913, n20914, n20915, n20916, n20917, n20918,
    n20919, n20920, n20921, n20922, n20923, n20924,
    n20925, n20926, n20927, n20928, n20929, n20930,
    n20931, n20932, n20933, n20934, n20935, n20936,
    n20937, n20938, n20939, n20940, n20941, n20942,
    n20943, n20944, n20945, n20946, n20947, n20948,
    n20949, n20950, n20951, n20952, n20953, n20954,
    n20955, n20956, n20957, n20958, n20959, n20960,
    n20961, n20962, n20963, n20964, n20965, n20966,
    n20967, n20968, n20969, n20970, n20971, n20972,
    n20973, n20974, n20975, n20976, n20977, n20978,
    n20979, n20980, n20981, n20982, n20983, n20984,
    n20985, n20986, n20987, n20988, n20989, n20990,
    n20991, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008,
    n21009, n21010, n21011, n21012, n21013, n21014,
    n21015, n21016, n21017, n21018, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026,
    n21027, n21028, n21029, n21030, n21031, n21032,
    n21033, n21034, n21035, n21036, n21037, n21038,
    n21039, n21040, n21041, n21042, n21043, n21044,
    n21045, n21046, n21047, n21048, n21049, n21050,
    n21051, n21052, n21053, n21054, n21055, n21056,
    n21057, n21058, n21059, n21060, n21061, n21062,
    n21063, n21064, n21065, n21066, n21067, n21068,
    n21069, n21070, n21071, n21072, n21073, n21074,
    n21075, n21076, n21077, n21078, n21079, n21080,
    n21081, n21082, n21083, n21084, n21085, n21086,
    n21087, n21088, n21089, n21090, n21091, n21092,
    n21093, n21094, n21095, n21096, n21097, n21098,
    n21099, n21100, n21101, n21102, n21103, n21104,
    n21105, n21106, n21107, n21108, n21109, n21110,
    n21111, n21112, n21113, n21114, n21115, n21116,
    n21117, n21118, n21119, n21120, n21121, n21122,
    n21123, n21124, n21125, n21126, n21127, n21128,
    n21129, n21130, n21131, n21132, n21133, n21134,
    n21135, n21136, n21137, n21138, n21139, n21140,
    n21141, n21142, n21143, n21144, n21145, n21146,
    n21147, n21148, n21149, n21150, n21151, n21152,
    n21153, n21154, n21155, n21156, n21157, n21158,
    n21159, n21160, n21161, n21162, n21163, n21164,
    n21165, n21166, n21167, n21168, n21169, n21170,
    n21171, n21172, n21173, n21174, n21175, n21176,
    n21177, n21178, n21179, n21180, n21181, n21182,
    n21183, n21184, n21185, n21186, n21187, n21188,
    n21189, n21190, n21191, n21192, n21193, n21194,
    n21195, n21196, n21197, n21198, n21199, n21200,
    n21201, n21202, n21203, n21204, n21205, n21206,
    n21207, n21208, n21209, n21210, n21211, n21212,
    n21213, n21214, n21215, n21216, n21217, n21218,
    n21219, n21220, n21221, n21222, n21223, n21224,
    n21225, n21226, n21227, n21228, n21229, n21230,
    n21231, n21232, n21233, n21234, n21235, n21236,
    n21237, n21238, n21239, n21240, n21241, n21242,
    n21243, n21244, n21245, n21246, n21247, n21248,
    n21249, n21250, n21251, n21252, n21253, n21254,
    n21255, n21256, n21257, n21258, n21259, n21260,
    n21261, n21262, n21263, n21264, n21265, n21266,
    n21267, n21268, n21269, n21270, n21271, n21272,
    n21273, n21274, n21275, n21276, n21277, n21278,
    n21279, n21280, n21281, n21282, n21283, n21284,
    n21285, n21286, n21287, n21288, n21289, n21290,
    n21291, n21292, n21293, n21294, n21295, n21296,
    n21297, n21298, n21299, n21300, n21301, n21302,
    n21303, n21304, n21305, n21306, n21307, n21308,
    n21309, n21310, n21311, n21312, n21313, n21314,
    n21315, n21316, n21317, n21318, n21319, n21320,
    n21321, n21322, n21323, n21324, n21325, n21326,
    n21327, n21328, n21329, n21330, n21331, n21332,
    n21333, n21334, n21335, n21336, n21337, n21338,
    n21339, n21340, n21341, n21342, n21343, n21344,
    n21345, n21346, n21347, n21348, n21349, n21350,
    n21351, n21352, n21353, n21354, n21355, n21356,
    n21357, n21358, n21359, n21360, n21361, n21362,
    n21363, n21364, n21365, n21366, n21367, n21368,
    n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428,
    n21429, n21430, n21431, n21432, n21433, n21434,
    n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21446,
    n21447, n21448, n21449, n21450, n21451, n21452,
    n21453, n21454, n21455, n21456, n21457, n21458,
    n21459, n21460, n21461, n21462, n21463, n21464,
    n21465, n21466, n21467, n21468, n21469, n21470,
    n21471, n21472, n21473, n21474, n21475, n21476,
    n21477, n21478, n21479, n21480, n21481, n21482,
    n21483, n21484, n21485, n21486, n21487, n21488,
    n21489, n21490, n21491, n21492, n21493, n21494,
    n21495, n21496, n21497, n21498, n21499, n21500,
    n21501, n21502, n21503, n21504, n21505, n21506,
    n21507, n21508, n21509, n21510, n21511, n21512,
    n21513, n21514, n21515, n21516, n21517, n21518,
    n21519, n21520, n21521, n21522, n21523, n21524,
    n21525, n21526, n21527, n21528, n21529, n21530,
    n21531, n21532, n21533, n21534, n21535, n21536,
    n21537, n21538, n21539, n21540, n21541, n21542,
    n21543, n21544, n21545, n21546, n21547, n21548,
    n21549, n21550, n21551, n21552, n21553, n21554,
    n21555, n21556, n21557, n21558, n21559, n21560,
    n21561, n21562, n21563, n21564, n21565, n21566,
    n21567, n21568, n21569, n21570, n21571, n21572,
    n21573, n21574, n21575, n21576, n21577, n21578,
    n21579, n21580, n21581, n21582, n21583, n21584,
    n21585, n21586, n21587, n21588, n21589, n21590,
    n21591, n21592, n21593, n21594, n21595, n21596,
    n21597, n21598, n21599, n21600, n21601, n21602,
    n21603, n21604, n21605, n21606, n21607, n21608,
    n21609, n21610, n21611, n21612, n21613, n21614,
    n21615, n21616, n21617, n21618, n21619, n21620,
    n21621, n21622, n21623, n21624, n21625, n21626,
    n21627, n21628, n21629, n21630, n21631, n21632,
    n21633, n21634, n21635, n21636, n21637, n21638,
    n21639, n21640, n21641, n21642, n21643, n21644,
    n21645, n21646, n21647, n21648, n21649, n21650,
    n21651, n21652, n21653, n21654, n21655, n21656,
    n21657, n21658, n21659, n21660, n21661, n21662,
    n21663, n21664, n21665, n21666, n21667, n21668,
    n21669, n21670, n21671, n21672, n21673, n21674,
    n21675, n21676, n21677, n21678, n21679, n21680,
    n21681, n21682, n21683, n21684, n21685, n21686,
    n21687, n21688, n21689, n21690, n21691, n21692,
    n21693, n21694, n21695, n21696, n21697, n21698,
    n21699, n21700, n21701, n21702, n21703, n21704,
    n21705, n21706, n21707, n21708, n21709, n21710,
    n21711, n21712, n21713, n21714, n21715, n21716,
    n21717, n21718, n21719, n21720, n21721, n21722,
    n21723, n21724, n21725, n21726, n21727, n21728,
    n21729, n21730, n21731, n21732, n21733, n21734,
    n21735, n21736, n21737, n21738, n21739, n21740,
    n21741, n21742, n21743, n21744, n21745, n21746,
    n21747, n21748, n21749, n21750, n21751, n21752,
    n21753, n21754, n21755, n21756, n21757, n21758,
    n21759, n21760, n21761, n21762, n21763, n21764,
    n21765, n21766, n21767, n21768, n21769, n21770,
    n21771, n21772, n21773, n21774, n21775, n21776,
    n21777, n21778, n21779, n21780, n21781, n21782,
    n21783, n21784, n21785, n21786, n21787, n21788,
    n21789, n21790, n21791, n21792, n21793, n21794,
    n21795, n21796, n21797, n21798, n21799, n21800,
    n21801, n21802, n21803, n21804, n21805, n21806,
    n21807, n21808, n21809, n21810, n21811, n21812,
    n21813, n21814, n21815, n21816, n21817, n21818,
    n21819, n21820, n21821, n21822, n21823, n21824,
    n21825, n21826, n21827, n21828, n21829, n21830,
    n21831, n21832, n21833, n21834, n21835, n21836,
    n21837, n21838, n21839, n21840, n21841, n21842,
    n21843, n21844, n21845, n21846, n21847, n21848,
    n21849, n21850, n21851, n21852, n21853, n21854,
    n21855, n21856, n21857, n21858, n21859, n21860,
    n21861, n21862, n21863, n21864, n21865, n21866,
    n21867, n21868, n21869, n21870, n21871, n21872,
    n21873, n21874, n21875, n21876, n21877, n21878,
    n21879, n21880, n21881, n21882, n21883, n21884,
    n21885, n21886, n21887, n21888, n21889, n21890,
    n21891, n21892, n21893, n21894, n21895, n21896,
    n21897, n21898, n21899, n21900, n21901, n21902,
    n21903, n21904, n21905, n21906, n21907, n21908,
    n21909, n21910, n21911, n21912, n21913, n21914,
    n21915, n21916, n21917, n21918, n21919, n21920,
    n21921, n21922, n21923, n21924, n21925, n21926,
    n21927, n21928, n21929, n21930, n21931, n21932,
    n21933, n21934, n21935, n21936, n21937, n21938,
    n21939, n21940, n21941, n21942, n21943, n21944,
    n21945, n21946, n21947, n21948, n21949, n21950,
    n21951, n21952, n21953, n21954, n21955, n21956,
    n21957, n21958, n21959, n21960, n21961, n21962,
    n21963, n21964, n21965, n21966, n21967, n21968,
    n21969, n21970, n21971, n21972, n21973, n21974,
    n21975, n21976, n21977, n21978, n21979, n21980,
    n21981, n21982, n21983, n21984, n21985, n21986,
    n21987, n21988, n21989, n21990, n21991, n21992,
    n21993, n21994, n21995, n21996, n21997, n21998,
    n21999, n22000, n22001, n22002, n22003, n22004,
    n22005, n22006, n22007, n22008, n22009, n22010,
    n22011, n22012, n22013, n22014, n22015, n22016,
    n22017, n22018, n22019, n22020, n22021, n22022,
    n22023, n22024, n22025, n22026, n22027, n22028,
    n22029, n22030, n22031, n22032, n22033, n22034,
    n22035, n22036, n22037, n22038, n22039, n22040,
    n22041, n22042, n22043, n22044, n22045, n22046,
    n22047, n22048, n22049, n22050, n22051, n22052,
    n22053, n22054, n22055, n22056, n22057, n22058,
    n22059, n22060, n22061, n22062, n22063, n22064,
    n22065, n22066, n22067, n22068, n22069, n22070,
    n22071, n22072, n22073, n22074, n22075, n22076,
    n22077, n22078, n22079, n22080, n22081, n22082,
    n22083, n22084, n22085, n22086, n22087, n22088,
    n22089, n22090, n22091, n22092, n22093, n22094,
    n22095, n22096, n22097, n22098, n22099, n22100,
    n22101, n22102, n22103, n22104, n22105, n22106,
    n22107, n22108, n22109, n22110, n22111, n22112,
    n22113, n22114, n22115, n22116, n22117, n22118,
    n22119, n22120, n22121, n22122, n22123, n22124,
    n22125, n22126, n22127, n22128, n22129, n22130,
    n22131, n22132, n22133, n22134, n22135, n22136,
    n22137, n22138, n22139, n22140, n22141, n22142,
    n22143, n22144, n22145, n22146, n22147, n22148,
    n22149, n22150, n22151, n22152, n22153, n22154,
    n22155, n22156, n22157, n22158, n22159, n22160,
    n22161, n22162, n22163, n22164, n22165, n22166,
    n22167, n22168, n22169, n22170, n22171, n22172,
    n22173, n22174, n22175, n22176, n22177, n22178,
    n22179, n22180, n22181, n22182, n22183, n22184,
    n22185, n22186, n22187, n22188, n22189, n22190,
    n22191, n22192, n22193, n22194, n22195, n22196,
    n22197, n22198, n22199, n22200, n22201, n22202,
    n22203, n22204, n22205, n22206, n22207, n22208,
    n22209, n22210, n22211, n22212, n22213, n22214,
    n22215, n22216, n22217, n22218, n22219, n22220,
    n22221, n22222, n22223, n22224, n22225, n22226,
    n22227, n22228, n22229, n22230, n22231, n22232,
    n22233, n22234, n22235, n22236, n22237, n22238,
    n22239, n22240, n22241, n22242, n22243, n22244,
    n22245, n22246, n22247, n22248, n22249, n22250,
    n22251, n22252, n22253, n22254, n22255, n22256,
    n22257, n22258, n22259, n22260, n22261, n22262,
    n22263, n22264, n22265, n22266, n22267, n22268,
    n22269, n22270, n22271, n22272, n22273, n22274,
    n22275, n22276, n22277, n22278, n22279, n22280,
    n22281, n22282, n22283, n22284, n22285, n22286,
    n22287, n22288, n22289, n22290, n22291, n22292,
    n22293, n22294, n22295, n22296, n22297, n22298,
    n22299, n22300, n22301, n22302, n22303, n22304,
    n22305, n22306, n22307, n22308, n22309, n22310,
    n22311, n22312, n22313, n22314, n22315, n22316,
    n22317, n22318, n22319, n22320, n22321, n22322,
    n22323, n22324, n22325, n22326, n22327, n22328,
    n22329, n22330, n22331, n22332, n22333, n22334,
    n22335, n22336, n22337, n22338, n22339, n22340,
    n22341, n22342, n22343, n22344, n22345, n22346,
    n22347, n22348, n22349, n22350, n22351, n22352,
    n22353, n22354, n22355, n22356, n22357, n22358,
    n22359, n22360, n22361, n22362, n22363, n22364,
    n22365, n22366, n22367, n22368, n22369, n22370,
    n22371, n22372, n22373, n22374, n22375, n22376,
    n22377, n22378, n22379, n22380, n22381, n22382,
    n22383, n22384, n22385, n22386, n22387, n22388,
    n22389, n22390, n22391, n22392, n22393, n22394,
    n22395, n22396, n22397, n22398, n22399, n22400,
    n22401, n22402, n22403, n22404, n22405, n22406,
    n22407, n22408, n22409, n22410, n22411, n22412,
    n22413, n22414, n22415, n22416, n22417, n22418,
    n22419, n22420, n22421, n22422, n22423, n22424,
    n22425, n22426, n22427, n22428, n22429, n22430,
    n22431, n22432, n22433, n22434, n22435, n22436,
    n22437, n22438, n22439, n22440, n22441, n22442,
    n22443, n22444, n22445, n22446, n22447, n22448,
    n22449, n22450, n22451, n22452, n22453, n22454,
    n22455, n22456, n22457, n22458, n22459, n22460,
    n22461, n22462, n22463, n22464, n22465, n22466,
    n22467, n22468, n22469, n22470, n22471, n22472,
    n22473, n22474, n22475, n22476, n22477, n22478,
    n22479, n22480, n22481, n22482, n22483, n22484,
    n22485, n22486, n22487, n22488, n22489, n22490,
    n22491, n22492, n22493, n22494, n22495, n22496,
    n22497, n22498, n22499, n22500, n22501, n22502,
    n22503, n22504, n22505, n22506, n22507, n22508,
    n22509, n22510, n22511, n22512, n22513, n22514,
    n22515, n22516, n22517, n22518, n22519, n22520,
    n22521, n22522, n22523, n22524, n22525, n22526,
    n22527, n22528, n22529, n22530, n22531, n22532,
    n22533, n22534, n22535, n22536, n22537, n22538,
    n22539, n22540, n22541, n22542, n22543, n22544,
    n22545, n22546, n22547, n22548, n22549, n22550,
    n22551, n22552, n22553, n22554, n22555, n22556,
    n22557, n22558, n22559, n22560, n22561, n22562,
    n22563, n22564, n22565, n22566, n22567, n22568,
    n22569, n22570, n22571, n22572, n22573, n22574,
    n22575, n22576, n22577, n22578, n22579, n22580,
    n22581, n22582, n22583, n22584, n22585, n22586,
    n22587, n22588, n22589, n22590, n22591, n22592,
    n22593, n22594, n22595, n22596, n22597, n22598,
    n22599, n22600, n22601, n22602, n22603, n22604,
    n22605, n22606, n22607, n22608, n22609, n22610,
    n22611, n22612, n22613, n22614, n22615, n22616,
    n22617, n22618, n22619, n22620, n22621, n22622,
    n22623, n22624, n22625, n22626, n22627, n22628,
    n22629, n22630, n22631, n22632, n22633, n22634,
    n22635, n22636, n22637, n22638, n22639, n22640,
    n22641, n22642, n22643, n22644, n22645, n22646,
    n22647, n22648, n22649, n22650, n22651, n22652,
    n22653, n22654, n22655, n22656, n22657, n22658,
    n22659, n22660, n22661, n22662, n22663, n22664,
    n22665, n22666, n22667, n22668, n22669, n22670,
    n22671, n22672, n22673, n22674, n22675, n22676,
    n22677, n22678, n22679, n22680, n22681, n22682,
    n22683, n22684, n22685, n22686, n22687, n22688,
    n22689, n22690, n22691, n22692, n22693, n22694,
    n22695, n22696, n22697, n22698, n22699, n22700,
    n22701, n22702, n22703, n22704, n22705, n22706,
    n22707, n22708, n22709, n22710, n22711, n22712,
    n22713, n22714, n22715, n22716, n22717, n22718,
    n22719, n22720, n22721, n22722, n22723, n22724,
    n22725, n22726, n22727, n22728, n22729, n22730,
    n22731, n22732, n22733, n22734, n22735, n22736,
    n22737, n22738, n22739, n22740, n22741, n22742,
    n22743, n22744, n22745, n22746, n22747, n22748,
    n22749, n22750, n22751, n22752, n22753, n22754,
    n22755, n22756, n22757, n22758, n22759, n22760,
    n22761, n22762, n22763, n22764, n22765, n22766,
    n22767, n22768, n22769, n22770, n22771, n22772,
    n22773, n22774, n22775, n22776, n22777, n22778,
    n22779, n22780, n22781, n22782, n22783, n22784,
    n22785, n22786, n22787, n22788, n22789, n22790,
    n22791, n22792, n22793, n22794, n22795, n22796,
    n22797, n22798, n22799, n22800, n22801, n22802,
    n22803, n22804, n22805, n22806, n22807, n22808,
    n22809, n22810, n22811, n22812, n22813, n22814,
    n22815, n22816, n22817, n22818, n22819, n22820,
    n22821, n22822, n22823, n22824, n22825, n22826,
    n22827, n22828, n22829, n22830, n22831, n22832,
    n22833, n22834, n22835, n22836, n22837, n22838,
    n22839, n22840, n22841, n22842, n22843, n22844,
    n22845, n22846, n22847, n22848, n22849, n22850,
    n22851, n22852, n22853, n22854, n22855, n22856,
    n22857, n22858, n22859, n22860, n22861, n22862,
    n22863, n22864, n22865, n22866, n22867, n22868,
    n22869, n22870, n22871, n22872, n22873, n22874,
    n22875, n22876, n22877, n22878, n22879, n22880,
    n22881, n22882, n22883, n22884, n22885, n22886,
    n22887, n22888, n22889, n22890, n22891, n22892,
    n22893, n22894, n22895, n22896, n22897, n22898,
    n22899, n22900, n22901, n22902, n22903, n22904,
    n22905, n22906, n22907, n22908, n22909, n22910,
    n22911, n22912, n22913, n22914, n22915, n22916,
    n22917, n22918, n22919, n22920, n22921, n22922,
    n22923, n22924, n22925, n22926, n22927, n22928,
    n22929, n22930, n22931, n22932, n22933, n22934,
    n22935, n22936, n22937, n22938, n22939, n22940,
    n22941, n22942, n22943, n22944, n22945, n22946,
    n22947, n22948, n22949, n22950, n22951, n22952,
    n22953, n22954, n22955, n22956, n22957, n22958,
    n22959, n22960, n22961, n22962, n22963, n22964,
    n22965, n22966, n22967, n22968, n22969, n22970,
    n22971, n22972, n22973, n22974, n22975, n22976,
    n22977, n22978, n22979, n22980, n22981, n22982,
    n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994,
    n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012,
    n23013, n23014, n23015, n23016, n23017, n23018,
    n23019, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n23028, n23029, n23030,
    n23031, n23032, n23033, n23034, n23035, n23036,
    n23037, n23038, n23039, n23040, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048,
    n23049, n23050, n23051, n23052, n23053, n23054,
    n23055, n23056, n23057, n23058, n23059, n23060,
    n23061, n23062, n23063, n23064, n23065, n23066,
    n23067, n23068, n23069, n23070, n23071, n23072,
    n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084,
    n23085, n23086, n23087, n23088, n23089, n23090,
    n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102,
    n23103, n23104, n23105, n23106, n23107, n23108,
    n23109, n23110, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120,
    n23121, n23122, n23123, n23124, n23125, n23126,
    n23127, n23128, n23129, n23130, n23131, n23132,
    n23133, n23134, n23135, n23136, n23137, n23138,
    n23139, n23140, n23141, n23142, n23143, n23144,
    n23145, n23146, n23147, n23148, n23149, n23150,
    n23151, n23152, n23153, n23154, n23155, n23156,
    n23157, n23158, n23159, n23160, n23161, n23162,
    n23163, n23164, n23165, n23166, n23167, n23168,
    n23169, n23170, n23171, n23172, n23173, n23174,
    n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186,
    n23187, n23188, n23189, n23190, n23191, n23192,
    n23193, n23194, n23195, n23196, n23197, n23198,
    n23199, n23200, n23201, n23202, n23203, n23204,
    n23205, n23206, n23207, n23208, n23209, n23210,
    n23211, n23212, n23213, n23214, n23215, n23216,
    n23217, n23218, n23219, n23220, n23221, n23222,
    n23223, n23224, n23225, n23226, n23227, n23228,
    n23229, n23230, n23231, n23232, n23233, n23234,
    n23235, n23236, n23237, n23238, n23239, n23240,
    n23241, n23242, n23243, n23244, n23245, n23246,
    n23247, n23248, n23249, n23250, n23251, n23252,
    n23253, n23254, n23255, n23256, n23257, n23258,
    n23259, n23260, n23261, n23262, n23263, n23264,
    n23265, n23266, n23267, n23268, n23269, n23270,
    n23271, n23272, n23273, n23274, n23275, n23276,
    n23277, n23278, n23279, n23280, n23281, n23282,
    n23283, n23284, n23285, n23286, n23287, n23288,
    n23289, n23290, n23291, n23292, n23293, n23294,
    n23295, n23296, n23297, n23298, n23299, n23300,
    n23301, n23302, n23303, n23304, n23305, n23306,
    n23307, n23308, n23309, n23310, n23311, n23312,
    n23313, n23314, n23315, n23316, n23317, n23318,
    n23319, n23320, n23321, n23322, n23323, n23324,
    n23325, n23326, n23327, n23328, n23329, n23330,
    n23331, n23332, n23333, n23334, n23335, n23336,
    n23337, n23338, n23339, n23340, n23341, n23342,
    n23343, n23344, n23345, n23346, n23347, n23348,
    n23349, n23350, n23351, n23352, n23353, n23354,
    n23355, n23356, n23357, n23358, n23359, n23360,
    n23361, n23362, n23363, n23364, n23365, n23366,
    n23367, n23368, n23369, n23370, n23371, n23372,
    n23373, n23374, n23375, n23376, n23377, n23378,
    n23379, n23380, n23381, n23382, n23383, n23384,
    n23385, n23386, n23387, n23388, n23389, n23390,
    n23391, n23392, n23393, n23394, n23395, n23396,
    n23397, n23398, n23399, n23400, n23401, n23402,
    n23403, n23404, n23405, n23406, n23407, n23408,
    n23409, n23410, n23411, n23412, n23413, n23414,
    n23415, n23416, n23417, n23418, n23419, n23420,
    n23421, n23422, n23423, n23424, n23425, n23426,
    n23427, n23428, n23429, n23430, n23431, n23432,
    n23433, n23434, n23435, n23436, n23437, n23438,
    n23439, n23440, n23441, n23442, n23443, n23444,
    n23445, n23446, n23447, n23448, n23449, n23450,
    n23451, n23452, n23453, n23454, n23455, n23456,
    n23457, n23458, n23459, n23460, n23461, n23462,
    n23463, n23464, n23465, n23466, n23467, n23468,
    n23469, n23470, n23471, n23472, n23473, n23474,
    n23475, n23476, n23477, n23478, n23479, n23480,
    n23481, n23482, n23483, n23484, n23485, n23486,
    n23487, n23488, n23489, n23490, n23491, n23492,
    n23493, n23494, n23495, n23496, n23497, n23498,
    n23499, n23500, n23501, n23502, n23503, n23504,
    n23505, n23506, n23507, n23508, n23509, n23510,
    n23511, n23512, n23513, n23514, n23515, n23516,
    n23517, n23518, n23519, n23520, n23521, n23522,
    n23523, n23524, n23525, n23526, n23527, n23528,
    n23529, n23530, n23531, n23532, n23533, n23534,
    n23535, n23536, n23537, n23538, n23539, n23540,
    n23541, n23542, n23543, n23544, n23545, n23546,
    n23547, n23548, n23549, n23550, n23551, n23552,
    n23553, n23554, n23555, n23556, n23557, n23558,
    n23559, n23560, n23561, n23562, n23563, n23564,
    n23565, n23566, n23567, n23568, n23569, n23570,
    n23571, n23572, n23573, n23574, n23575, n23576,
    n23577, n23578, n23579, n23580, n23581, n23582,
    n23583, n23584, n23585, n23586, n23587, n23588,
    n23589, n23590, n23591, n23592, n23593, n23594,
    n23595, n23596, n23597, n23598, n23599, n23600,
    n23601, n23602, n23603, n23604, n23605, n23606,
    n23607, n23608, n23609, n23610, n23611, n23612,
    n23613, n23614, n23615, n23616, n23617, n23618,
    n23619, n23620, n23621, n23622, n23623, n23624,
    n23625, n23626, n23627, n23628, n23629, n23630,
    n23631, n23632, n23633, n23634, n23635, n23636,
    n23637, n23638, n23639, n23640, n23641, n23642,
    n23643, n23644, n23645, n23646, n23647, n23648,
    n23649, n23650, n23651, n23652, n23653, n23654,
    n23655, n23656, n23657, n23658, n23659, n23660,
    n23661, n23662, n23663, n23664, n23665, n23666,
    n23667, n23668, n23669, n23670, n23671, n23672,
    n23673, n23674, n23675, n23676, n23677, n23678,
    n23679, n23680, n23681, n23682, n23683, n23684,
    n23685, n23686, n23687, n23688, n23689, n23690,
    n23691, n23692, n23693, n23694, n23695, n23696,
    n23697, n23698, n23699, n23700, n23701, n23702,
    n23703, n23704, n23705, n23706, n23707, n23708,
    n23709, n23710, n23711, n23712, n23713, n23714,
    n23715, n23716, n23717, n23718, n23719, n23720,
    n23721, n23722, n23723, n23724, n23725, n23726,
    n23727, n23728, n23729, n23730, n23731, n23732,
    n23733, n23734, n23735, n23736, n23737, n23738,
    n23739, n23740, n23741, n23742, n23743, n23744,
    n23745, n23746, n23747, n23748, n23749, n23750,
    n23751, n23752, n23753, n23754, n23755, n23756,
    n23757, n23758, n23759, n23760, n23761, n23762,
    n23763, n23764, n23765, n23766, n23767, n23768,
    n23769, n23770, n23771, n23772, n23773, n23774,
    n23775, n23776, n23777, n23778, n23779, n23780,
    n23781, n23782, n23783, n23784, n23785, n23786,
    n23787, n23788, n23789, n23790, n23791, n23792,
    n23793, n23794, n23795, n23796, n23797, n23798,
    n23799, n23800, n23801, n23802, n23803, n23804,
    n23805, n23806, n23807, n23808, n23809, n23810,
    n23811, n23812, n23813, n23814, n23815, n23816,
    n23817, n23818, n23819, n23820, n23821, n23822,
    n23823, n23824, n23825, n23826, n23827, n23828,
    n23829, n23830, n23831, n23832, n23833, n23834,
    n23835, n23836, n23837, n23838, n23839, n23840,
    n23841, n23842, n23843, n23844, n23845, n23846,
    n23847, n23848, n23849, n23850, n23851, n23852,
    n23853, n23854, n23855, n23856, n23857, n23858,
    n23859, n23860, n23861, n23862, n23863, n23864,
    n23865, n23866, n23867, n23868, n23869, n23870,
    n23871, n23872, n23873, n23874, n23875, n23876,
    n23877, n23878, n23879, n23880, n23881, n23882,
    n23883, n23884, n23885, n23886, n23887, n23888,
    n23889, n23890, n23891, n23892, n23893, n23894,
    n23895, n23896, n23897, n23898, n23899, n23900,
    n23901, n23902, n23903, n23904, n23905, n23906,
    n23907, n23908, n23909, n23910, n23911, n23912,
    n23913, n23914, n23915, n23916, n23917, n23918,
    n23919, n23920, n23921, n23922, n23923, n23924,
    n23925, n23926, n23927, n23928, n23929, n23930,
    n23931, n23932, n23933, n23934, n23935, n23936,
    n23937, n23938, n23939, n23940, n23941, n23942,
    n23943, n23944, n23945, n23946, n23947, n23948,
    n23949, n23950, n23951, n23952, n23953, n23954,
    n23955, n23956, n23957, n23958, n23959, n23960,
    n23961, n23962, n23963, n23964, n23965, n23966,
    n23967, n23968, n23969, n23970, n23971, n23972,
    n23973, n23974, n23975, n23976, n23977, n23978,
    n23979, n23980, n23981, n23982, n23983, n23984,
    n23985, n23986, n23987, n23988, n23989, n23990,
    n23991, n23992, n23993, n23994, n23995, n23996,
    n23997, n23998, n23999, n24000, n24001, n24002,
    n24003, n24004, n24005, n24006, n24007, n24008,
    n24009, n24010, n24011, n24012, n24013, n24014,
    n24015, n24016, n24017, n24018, n24019, n24020,
    n24021, n24022, n24023, n24024, n24025, n24026,
    n24027, n24028, n24029, n24030, n24031, n24032,
    n24033, n24034, n24035, n24036, n24037, n24038,
    n24039, n24040, n24041, n24042, n24043, n24044,
    n24045, n24046, n24047, n24048, n24049, n24050,
    n24051, n24052, n24053, n24054, n24055, n24056,
    n24057, n24058, n24059, n24060, n24061, n24062,
    n24063, n24064, n24065, n24066, n24067, n24068,
    n24069, n24070, n24071, n24072, n24073, n24074,
    n24075, n24076, n24077, n24078, n24079, n24080,
    n24081, n24082, n24083, n24084, n24085, n24086,
    n24087, n24088, n24089, n24090, n24091, n24092,
    n24093, n24094, n24095, n24096, n24097, n24098,
    n24099, n24100, n24101, n24102, n24103, n24104,
    n24105, n24106, n24107, n24108, n24109, n24110,
    n24111, n24112, n24113, n24114, n24115, n24116,
    n24117, n24118, n24119, n24120, n24121, n24122,
    n24123, n24124, n24125, n24126, n24127, n24128,
    n24129, n24130, n24131, n24132, n24133, n24134,
    n24135, n24136, n24137, n24138, n24139, n24140,
    n24141, n24142, n24143, n24144, n24145, n24146,
    n24147, n24148, n24149, n24150, n24151, n24152,
    n24153, n24154, n24155, n24156, n24157, n24158,
    n24159, n24160, n24161, n24162, n24163, n24164,
    n24165, n24166, n24167, n24168, n24169, n24170,
    n24171, n24172, n24173, n24174, n24175, n24176,
    n24177, n24178, n24179, n24180, n24181, n24182,
    n24183, n24184, n24185, n24186, n24187, n24188,
    n24189, n24190, n24191, n24192, n24193, n24194,
    n24195, n24196, n24197, n24198, n24199, n24200,
    n24201, n24202, n24203, n24204, n24205, n24206,
    n24207, n24208, n24209, n24210, n24211, n24212,
    n24213, n24214, n24215, n24216, n24217, n24218,
    n24219, n24220, n24221, n24222, n24223, n24224,
    n24225, n24226, n24227, n24228, n24229, n24230,
    n24231, n24232, n24233, n24234, n24235, n24236,
    n24237, n24238, n24239, n24240, n24241, n24242,
    n24243, n24244, n24245, n24246, n24247, n24248,
    n24249, n24250, n24251, n24252, n24253, n24254,
    n24255, n24256, n24257, n24258, n24259, n24260,
    n24261, n24262, n24263, n24264, n24265, n24266,
    n24267, n24268, n24269, n24270, n24271, n24272,
    n24273, n24274, n24275, n24276, n24277, n24278,
    n24279, n24280, n24281, n24282, n24283, n24284,
    n24285, n24286, n24287, n24288, n24289, n24290,
    n24291, n24292, n24293, n24294, n24295, n24296,
    n24297, n24298, n24299, n24300, n24301, n24302,
    n24303, n24304, n24305, n24306, n24307, n24308,
    n24309, n24310, n24311, n24312, n24313, n24314,
    n24315, n24316, n24317, n24318, n24319, n24320,
    n24321, n24322, n24323, n24324, n24325, n24326,
    n24327, n24328, n24329, n24330, n24331, n24332,
    n24333, n24334, n24335, n24336, n24337, n24338,
    n24339, n24340, n24341, n24342, n24343, n24344,
    n24345, n24346, n24347, n24348, n24349, n24350,
    n24351, n24352, n24353, n24354, n24355, n24356,
    n24357, n24358, n24359, n24360, n24361, n24362,
    n24363, n24364, n24365, n24366, n24367, n24368,
    n24369, n24370, n24371, n24372, n24373, n24374,
    n24375, n24376, n24377, n24378, n24379, n24380,
    n24381, n24382, n24383, n24384, n24385, n24386,
    n24387, n24388, n24389, n24390, n24391, n24392,
    n24393, n24394, n24395, n24396, n24397, n24398,
    n24399, n24400, n24401, n24402, n24403, n24404,
    n24405, n24406, n24407, n24408, n24409, n24410,
    n24411, n24412, n24413, n24414, n24415, n24416,
    n24417, n24418, n24419, n24420, n24421, n24422,
    n24423, n24424, n24425, n24426, n24427, n24428,
    n24429, n24430, n24431, n24432, n24433, n24434,
    n24435, n24436, n24437, n24438, n24439, n24440,
    n24441, n24442, n24443, n24444, n24445, n24446,
    n24447, n24448, n24449, n24450, n24451, n24452,
    n24453, n24454, n24455, n24456, n24457, n24458,
    n24459, n24460, n24461, n24462, n24463, n24464,
    n24465, n24466, n24467, n24468, n24469, n24470,
    n24471, n24472, n24473, n24474, n24475, n24476,
    n24477, n24478, n24479, n24480, n24481, n24482,
    n24483, n24484, n24485, n24486, n24487, n24488,
    n24489, n24490, n24491, n24492, n24493, n24494,
    n24495, n24496, n24497, n24498, n24499, n24500,
    n24501, n24502, n24503, n24504, n24505, n24506,
    n24507, n24508, n24509, n24510, n24511, n24512,
    n24513, n24514, n24515, n24516, n24517, n24518,
    n24519, n24520, n24521, n24522, n24523, n24524,
    n24525, n24526, n24527, n24528, n24529, n24530,
    n24531, n24532, n24533, n24534, n24535, n24536,
    n24537, n24538, n24539, n24540, n24541, n24542,
    n24543, n24544, n24545, n24546, n24547, n24548,
    n24549, n24550, n24551, n24552, n24553, n24554,
    n24555, n24556, n24557, n24558, n24559, n24560,
    n24561, n24562, n24563, n24564, n24565, n24566,
    n24567, n24568, n24569, n24570, n24571, n24572,
    n24573, n24574, n24575, n24576, n24577, n24578,
    n24579, n24580, n24581, n24582, n24583, n24584,
    n24585, n24586, n24587, n24588, n24589, n24590,
    n24591, n24592, n24593, n24594, n24595, n24596,
    n24597, n24598, n24599, n24600, n24601, n24602,
    n24603, n24604, n24605, n24606, n24607, n24608,
    n24609, n24610, n24611, n24612, n24613, n24614,
    n24615, n24616, n24617, n24618, n24619, n24620,
    n24621, n24622, n24623, n24624, n24625, n24626,
    n24627, n24628, n24629, n24630, n24631, n24632,
    n24633, n24634, n24635, n24636, n24637, n24638,
    n24639, n24640, n24641, n24642, n24643, n24644,
    n24645, n24646, n24647, n24648, n24649, n24650,
    n24651, n24652, n24653, n24654, n24655, n24656,
    n24657, n24658, n24659, n24660, n24661, n24662,
    n24663, n24664, n24665, n24666, n24667, n24668,
    n24669, n24670, n24671, n24672, n24673, n24674,
    n24675, n24676, n24677, n24678, n24679, n24680,
    n24681, n24682, n24683, n24684, n24685, n24686,
    n24687, n24688, n24689, n24690, n24691, n24692,
    n24693, n24694, n24695, n24696, n24697, n24698,
    n24699, n24700, n24701, n24702, n24703, n24704,
    n24705, n24706, n24707, n24708, n24709, n24710,
    n24711, n24712, n24713, n24714, n24715, n24716,
    n24717, n24718, n24719, n24720, n24721, n24722,
    n24723, n24724, n24725, n24726, n24727, n24728,
    n24729, n24730, n24731, n24732, n24733, n24734,
    n24735, n24736, n24737, n24738, n24739, n24740,
    n24741, n24742, n24743, n24744, n24745, n24746,
    n24747, n24748, n24749, n24750, n24751, n24752,
    n24753, n24754, n24755, n24756, n24757, n24758,
    n24759, n24760, n24761, n24762, n24763, n24764,
    n24765, n24766, n24767, n24768, n24769, n24770,
    n24771, n24772, n24773, n24774, n24775, n24776,
    n24777, n24778, n24779, n24780, n24781, n24782,
    n24783, n24784, n24785, n24786, n24787, n24788,
    n24789, n24790, n24791, n24792, n24793, n24794,
    n24795, n24796, n24797, n24798, n24799, n24800,
    n24801, n24802, n24803, n24804, n24805, n24806,
    n24807, n24808, n24809, n24810, n24811, n24812,
    n24813, n24814, n24815, n24816, n24817, n24818,
    n24819, n24820, n24821, n24822, n24823, n24824,
    n24825, n24826, n24827, n24828, n24829, n24830,
    n24831, n24832, n24833, n24834, n24835, n24836,
    n24837, n24838, n24839, n24840, n24841, n24842,
    n24843, n24844, n24845, n24846, n24847, n24848,
    n24849, n24850, n24851, n24852, n24853, n24854,
    n24855, n24856, n24857, n24858, n24859, n24860,
    n24861, n24862, n24863, n24864, n24865, n24866,
    n24867, n24868, n24869, n24870, n24871, n24872,
    n24873, n24874, n24875, n24876, n24877, n24878,
    n24879, n24880, n24881, n24882, n24883, n24884,
    n24885, n24886, n24887, n24888, n24889, n24890,
    n24891, n24892, n24893, n24894, n24895, n24896,
    n24897, n24898, n24899, n24900, n24901, n24902,
    n24903, n24904, n24905, n24906, n24907, n24908,
    n24909, n24910, n24911, n24912, n24913, n24914,
    n24915, n24916, n24917, n24918, n24919, n24920,
    n24921, n24922, n24923, n24924, n24925, n24926,
    n24927, n24928, n24929, n24930, n24931, n24932,
    n24933, n24934, n24935, n24936, n24937, n24938,
    n24939, n24940, n24941, n24942, n24943, n24944,
    n24945, n24946, n24947, n24948, n24949, n24950,
    n24951, n24952, n24953, n24954, n24955, n24956,
    n24957, n24958, n24959, n24960, n24961, n24962,
    n24963, n24964, n24965, n24966, n24967, n24968,
    n24969, n24970, n24971, n24972, n24973, n24974,
    n24975, n24976, n24977, n24978, n24979, n24980,
    n24981, n24982, n24983, n24984, n24985, n24986,
    n24987, n24988, n24989, n24990, n24991, n24992,
    n24993, n24994, n24995, n24996, n24997, n24998,
    n24999, n25000, n25001, n25002, n25003, n25004,
    n25005, n25006, n25007, n25008, n25009, n25010,
    n25011, n25012, n25013, n25014, n25015, n25016,
    n25017, n25018, n25019, n25020, n25021, n25022,
    n25023, n25024, n25025, n25026, n25027, n25028,
    n25029, n25030, n25031, n25032, n25033, n25034,
    n25035, n25036, n25037, n25038, n25039, n25040,
    n25041, n25042, n25043, n25044, n25045, n25046,
    n25047, n25048, n25049, n25050, n25051, n25052,
    n25053, n25054, n25055, n25056, n25057, n25058,
    n25059, n25060, n25061, n25062, n25063, n25064,
    n25065, n25066, n25067, n25068, n25069, n25070,
    n25071, n25072, n25073, n25074, n25075, n25076,
    n25077, n25078, n25079, n25080, n25081, n25082,
    n25083, n25084, n25085, n25086, n25087, n25088,
    n25089, n25090, n25091, n25092, n25093, n25094,
    n25095, n25096, n25097, n25098, n25099, n25100,
    n25101, n25102, n25103, n25104, n25105, n25106,
    n25107, n25108, n25109, n25110, n25111, n25112,
    n25113, n25114, n25115, n25116, n25117, n25118,
    n25119, n25120, n25121, n25122, n25123, n25124,
    n25125, n25126, n25127, n25128, n25129, n25130,
    n25131, n25132, n25133, n25134, n25135, n25136,
    n25137, n25138, n25139, n25140, n25141, n25142,
    n25143, n25144, n25145, n25146, n25147, n25148,
    n25149, n25150, n25151, n25152, n25153, n25154,
    n25155, n25156, n25157, n25158, n25159, n25160,
    n25161, n25162, n25163, n25164, n25165, n25166,
    n25167, n25168, n25169, n25170, n25171, n25172,
    n25173, n25174, n25175, n25176, n25177, n25178,
    n25179, n25180, n25181, n25182, n25183, n25184,
    n25185, n25186, n25187, n25188, n25189, n25190,
    n25191, n25192, n25193, n25194, n25195, n25196,
    n25197, n25198, n25199, n25200, n25201, n25202,
    n25203, n25204, n25205, n25206, n25207, n25208,
    n25209, n25210, n25211, n25212, n25213, n25214,
    n25215, n25216, n25217, n25218, n25219, n25220,
    n25221, n25222, n25223, n25224, n25225, n25226,
    n25227, n25228, n25229, n25230, n25231, n25232,
    n25233, n25234, n25235, n25236, n25237, n25238,
    n25239, n25240, n25241, n25242, n25243, n25244,
    n25245, n25246, n25247, n25248, n25249, n25250,
    n25251, n25252, n25253, n25254, n25255, n25256,
    n25257, n25258, n25259, n25260, n25261, n25262,
    n25263, n25264, n25265, n25266, n25267, n25268,
    n25269, n25270, n25271, n25272, n25273, n25274,
    n25275, n25276, n25277, n25278, n25279, n25280,
    n25281, n25282, n25283, n25284, n25285, n25286,
    n25287, n25288, n25289, n25290, n25291, n25292,
    n25293, n25294, n25295, n25296, n25297, n25298,
    n25299, n25300, n25301, n25302, n25303, n25304,
    n25305, n25306, n25307, n25308, n25309, n25310,
    n25311, n25312, n25313, n25314, n25315, n25316,
    n25317, n25318, n25319, n25320, n25321, n25322,
    n25323, n25324, n25325, n25326, n25327, n25328,
    n25329, n25330, n25331, n25332, n25333, n25334,
    n25335, n25336, n25337, n25338, n25339, n25340,
    n25341, n25342, n25343, n25344, n25345, n25346,
    n25347, n25348, n25349, n25350, n25351, n25352,
    n25353, n25354, n25355, n25356, n25357, n25358,
    n25359, n25360, n25361, n25362, n25363, n25364,
    n25365, n25366, n25367, n25368, n25369, n25370,
    n25371, n25372, n25373, n25374, n25375, n25376,
    n25377, n25378, n25379, n25380, n25381, n25382,
    n25383, n25384, n25385, n25386, n25387, n25388,
    n25389, n25390, n25391, n25392, n25393, n25394,
    n25395, n25396, n25397, n25398, n25399, n25400,
    n25401, n25402, n25403, n25404, n25405, n25406,
    n25407, n25408, n25409, n25410, n25411, n25412,
    n25413, n25414, n25415, n25416, n25417, n25418,
    n25419, n25420, n25421, n25422, n25423, n25424,
    n25425, n25426, n25427, n25428, n25429, n25430,
    n25431, n25432, n25433, n25434, n25435, n25436,
    n25437, n25438, n25439, n25440, n25441, n25442,
    n25443, n25444, n25445, n25446, n25447, n25448,
    n25449, n25450, n25451, n25452, n25453, n25454,
    n25455, n25456, n25457, n25458, n25459, n25460,
    n25461, n25462, n25463, n25464, n25465, n25466,
    n25467, n25468, n25469, n25470, n25471, n25472,
    n25473, n25474, n25475, n25476, n25477, n25478,
    n25479, n25480, n25481, n25482, n25483, n25484,
    n25485, n25486, n25487, n25488, n25489, n25490,
    n25491, n25492, n25493, n25494, n25495, n25496,
    n25497, n25498, n25499, n25500, n25501, n25502,
    n25503, n25504, n25505, n25506, n25507, n25508,
    n25509, n25510, n25511, n25512, n25513, n25514,
    n25515, n25516, n25517, n25518, n25519, n25520,
    n25521, n25522, n25523, n25524, n25525, n25526,
    n25527, n25528, n25529, n25530, n25531, n25532,
    n25533, n25534, n25535, n25536, n25537, n25538,
    n25539, n25540, n25541, n25542, n25543, n25544,
    n25545, n25546, n25547, n25548, n25549, n25550,
    n25551, n25552, n25553, n25554, n25555, n25556,
    n25557, n25558, n25559, n25560, n25561, n25562,
    n25563, n25564, n25565, n25566, n25567, n25568,
    n25569, n25570, n25571, n25572, n25573, n25574,
    n25575, n25576, n25577, n25578, n25579, n25580,
    n25581, n25582, n25583, n25584, n25585, n25586,
    n25587, n25588, n25589, n25590, n25591, n25592,
    n25593, n25594, n25595, n25596, n25597, n25598,
    n25599, n25600, n25601, n25602, n25603, n25604,
    n25605, n25606, n25607, n25608, n25609, n25610,
    n25611, n25612, n25613, n25614, n25615, n25616,
    n25617, n25618, n25619, n25620, n25621, n25622,
    n25623, n25624, n25625, n25626, n25627, n25628,
    n25629, n25630, n25631, n25632, n25633, n25634,
    n25635, n25636, n25637, n25638, n25639, n25640,
    n25641, n25642, n25643, n25644, n25645, n25646,
    n25647, n25648, n25649, n25650, n25651, n25652,
    n25653, n25654, n25655, n25656, n25657, n25658,
    n25659, n25660, n25661, n25662, n25663, n25664,
    n25665, n25666, n25667, n25668, n25669, n25670,
    n25671, n25672, n25673, n25674, n25675, n25676,
    n25677, n25678, n25679, n25680, n25681, n25682,
    n25683, n25684, n25685, n25686, n25687, n25688,
    n25689, n25690, n25691, n25692, n25693, n25694,
    n25695, n25696, n25697, n25698, n25699, n25700,
    n25701, n25702, n25703, n25704, n25705, n25706,
    n25707, n25708, n25709, n25710, n25711, n25712,
    n25713, n25714, n25715, n25716, n25717, n25718,
    n25719, n25720, n25721, n25722, n25723, n25724,
    n25725, n25726, n25727, n25728, n25729, n25730,
    n25731, n25732, n25733, n25734, n25735, n25736,
    n25737, n25738, n25739, n25740, n25741, n25742,
    n25743, n25744, n25745, n25746, n25747, n25748,
    n25749, n25750, n25751, n25752, n25753, n25754,
    n25755, n25756, n25757, n25758, n25759, n25760,
    n25761, n25762, n25763, n25764, n25765, n25766,
    n25767, n25768, n25769, n25770, n25771, n25772,
    n25773, n25774, n25775, n25776, n25777, n25778,
    n25779, n25780, n25781, n25782, n25783, n25784,
    n25785, n25786, n25787, n25788, n25789, n25790,
    n25791, n25792, n25793, n25794, n25795, n25796,
    n25797, n25798, n25799, n25800, n25801, n25802,
    n25803, n25804, n25805, n25806, n25807, n25808,
    n25809, n25810, n25811, n25812, n25813, n25814,
    n25815, n25816, n25817, n25818, n25819, n25820,
    n25821, n25822, n25823, n25824, n25825, n25826,
    n25827, n25828, n25829, n25830, n25831, n25832,
    n25833, n25834, n25835, n25836, n25837, n25838,
    n25839, n25840, n25841, n25842, n25843, n25844,
    n25845, n25846, n25847, n25848, n25849, n25850,
    n25851, n25852, n25853, n25854, n25855, n25856,
    n25857, n25858, n25859, n25860, n25861, n25862,
    n25863, n25864, n25865, n25866, n25867, n25868,
    n25869, n25870, n25871, n25872, n25873, n25874,
    n25875, n25876, n25877, n25878, n25879, n25880,
    n25881, n25882, n25883, n25884, n25885, n25886,
    n25887, n25888, n25889, n25890, n25891, n25892,
    n25893, n25894, n25895, n25896, n25897, n25898,
    n25899, n25900, n25901, n25902, n25903, n25904,
    n25905, n25906, n25907, n25908, n25909, n25910,
    n25911, n25912, n25913, n25914, n25915, n25916,
    n25917, n25918, n25919, n25920, n25921, n25922,
    n25923, n25924, n25925, n25926, n25927, n25928,
    n25929, n25930, n25931, n25932, n25933, n25934,
    n25935, n25936, n25937, n25938, n25939, n25940,
    n25941, n25942, n25943, n25944, n25945, n25946,
    n25947, n25948, n25949, n25950, n25951, n25952,
    n25953, n25954, n25955, n25956, n25957, n25958,
    n25959, n25960, n25961, n25962, n25963, n25964,
    n25965, n25966, n25967, n25968, n25969, n25970,
    n25971, n25972, n25973, n25974, n25975, n25976,
    n25977, n25978, n25979, n25980, n25981, n25982,
    n25983, n25984, n25985, n25986, n25987, n25988,
    n25989, n25990, n25991, n25992, n25993, n25994,
    n25995, n25996, n25997, n25998, n25999, n26000,
    n26001, n26002, n26003, n26004, n26005, n26006,
    n26007, n26008, n26009, n26010, n26011, n26012,
    n26013, n26014, n26015, n26016, n26017, n26018,
    n26019, n26020, n26021, n26022, n26023, n26024,
    n26025, n26026, n26027, n26028, n26029, n26030,
    n26031, n26032, n26033, n26034, n26035, n26036,
    n26037, n26038, n26039, n26040, n26041, n26042,
    n26043, n26044, n26045, n26046, n26047, n26048,
    n26049, n26050, n26051, n26052, n26053, n26054,
    n26055, n26056, n26057, n26058, n26059, n26060,
    n26061, n26062, n26063, n26064, n26065, n26066,
    n26067, n26068, n26069, n26070, n26071, n26072,
    n26073, n26074, n26075, n26076, n26077, n26078,
    n26079, n26080, n26081, n26082, n26083, n26084,
    n26085, n26086, n26087, n26088, n26089, n26090,
    n26091, n26092, n26093, n26094, n26095, n26096,
    n26097, n26098, n26099, n26100, n26101, n26102,
    n26103, n26104, n26105, n26106, n26107, n26108,
    n26109, n26110, n26111, n26112, n26113, n26114,
    n26115, n26116, n26117, n26118, n26119, n26120,
    n26121, n26122, n26123, n26124, n26125, n26126,
    n26127, n26128, n26129, n26130, n26131, n26132,
    n26133, n26134, n26135, n26136, n26137, n26138,
    n26139, n26140, n26141, n26142, n26143, n26144,
    n26145, n26146, n26147, n26148, n26149, n26150,
    n26151, n26152, n26153, n26154, n26155, n26156,
    n26157, n26158, n26159, n26160, n26161, n26162,
    n26163, n26164, n26165, n26166, n26167, n26168,
    n26169, n26170, n26171, n26172, n26173, n26174,
    n26175, n26176, n26177, n26178, n26179, n26180,
    n26181, n26182, n26183, n26184, n26185, n26186,
    n26187, n26188, n26189, n26190, n26191, n26192,
    n26193, n26194, n26195, n26196, n26197, n26198,
    n26199, n26200, n26201, n26202, n26203, n26204,
    n26205, n26206, n26207, n26208, n26209, n26210,
    n26211, n26212, n26213, n26214, n26215, n26216,
    n26217, n26218, n26219, n26220, n26221, n26222,
    n26223, n26224, n26225, n26226, n26227, n26228,
    n26229, n26230, n26231, n26232, n26233, n26234,
    n26235, n26236, n26237, n26238, n26239, n26240,
    n26241, n26242, n26243, n26244, n26245, n26246,
    n26247, n26248, n26249, n26250, n26251, n26252,
    n26253, n26254, n26255, n26256, n26257, n26258,
    n26259, n26260, n26261, n26262, n26263, n26264,
    n26265, n26266, n26267, n26268, n26269, n26270,
    n26271, n26272, n26273, n26274, n26275, n26276,
    n26277, n26278, n26279, n26280, n26281, n26282,
    n26283, n26284, n26285, n26286, n26287, n26288,
    n26289, n26290, n26291, n26292, n26293, n26294,
    n26295, n26296, n26297, n26298, n26299, n26300,
    n26301, n26302, n26303, n26304, n26305, n26306,
    n26307, n26308, n26309, n26310, n26311, n26312,
    n26313, n26314, n26315, n26316, n26317, n26318,
    n26319, n26320, n26321, n26322, n26323, n26324,
    n26325, n26326, n26327, n26328, n26329, n26330,
    n26331, n26332, n26333, n26334, n26335, n26336,
    n26337, n26338, n26339, n26340, n26341, n26342,
    n26343, n26344, n26345, n26346, n26347, n26348,
    n26349, n26350, n26351, n26352, n26353, n26354,
    n26355, n26356, n26357, n26358, n26359, n26360,
    n26361, n26362, n26363, n26364, n26365, n26366,
    n26367, n26368, n26369, n26370, n26371, n26372,
    n26373, n26374, n26375, n26376, n26377, n26378,
    n26379, n26380, n26381, n26382, n26383, n26384,
    n26385, n26386, n26387, n26388, n26389, n26390,
    n26391, n26392, n26393, n26394, n26395, n26396,
    n26397, n26398, n26399, n26400, n26401, n26402,
    n26403, n26404, n26405, n26406, n26407, n26408,
    n26409, n26410, n26411, n26412, n26413, n26414,
    n26415, n26416, n26417, n26418, n26419, n26420,
    n26421, n26422, n26423, n26424, n26425, n26426,
    n26427, n26428, n26429, n26430, n26431, n26432,
    n26433, n26434, n26435, n26436, n26437, n26438,
    n26439, n26440, n26441, n26442, n26443, n26444,
    n26445, n26446, n26447, n26448, n26449, n26450,
    n26451, n26452, n26453, n26454, n26455, n26456,
    n26457, n26458, n26459, n26460, n26461, n26462,
    n26463, n26464, n26465, n26466, n26467, n26468,
    n26469, n26470, n26471, n26472, n26473, n26474,
    n26475, n26476, n26477, n26478, n26479, n26480,
    n26481, n26482, n26483, n26484, n26485, n26486,
    n26487, n26488, n26489, n26490, n26491, n26492,
    n26493, n26494, n26495, n26496, n26497, n26498,
    n26499, n26500, n26501, n26502, n26503, n26504,
    n26505, n26506, n26507, n26508, n26509, n26510,
    n26511, n26512, n26513, n26514, n26515, n26516,
    n26517, n26518, n26519, n26520, n26521, n26522,
    n26523, n26524, n26525, n26526, n26527, n26528,
    n26529, n26530, n26531, n26532, n26533, n26534,
    n26535, n26536, n26537, n26538, n26539, n26540,
    n26541, n26542, n26543, n26544, n26545, n26546,
    n26547, n26548, n26549, n26550, n26551, n26552,
    n26553, n26554, n26555, n26556, n26557, n26558,
    n26559, n26560, n26561, n26562, n26563, n26564,
    n26565, n26566, n26567, n26568, n26569, n26570,
    n26571, n26572, n26573, n26574, n26575, n26576,
    n26577, n26578, n26579, n26580, n26581, n26582,
    n26583, n26584, n26585, n26586, n26587, n26588,
    n26589, n26590, n26591, n26592, n26593, n26594,
    n26595, n26596, n26597, n26598, n26599, n26600,
    n26601, n26602, n26603, n26604, n26605, n26606,
    n26607, n26608, n26609, n26610, n26611, n26612,
    n26613, n26614, n26615, n26616, n26617, n26618,
    n26619, n26620, n26621, n26622, n26623, n26624,
    n26625, n26626, n26627, n26628, n26629, n26630,
    n26631, n26632, n26633, n26634, n26635, n26636,
    n26637, n26638, n26639, n26640, n26641, n26642,
    n26643, n26644, n26645, n26646, n26647, n26648,
    n26649, n26650, n26651, n26652, n26653, n26654,
    n26655, n26656, n26657, n26658, n26659, n26660,
    n26661, n26662, n26663, n26664, n26665, n26666,
    n26667, n26668, n26669, n26670, n26671, n26672,
    n26673, n26674, n26675, n26676, n26677, n26678,
    n26679, n26680, n26681, n26682, n26683, n26684,
    n26685, n26686, n26687, n26688, n26689, n26690,
    n26691, n26692, n26693, n26694, n26695, n26696,
    n26697, n26698, n26699, n26700, n26701, n26702,
    n26703, n26704, n26705, n26706, n26707, n26708,
    n26709, n26710, n26711, n26712, n26713, n26714,
    n26715, n26716, n26717, n26718, n26719, n26720,
    n26721, n26722, n26723, n26724, n26725, n26726,
    n26727, n26728, n26729, n26730, n26731, n26732,
    n26733, n26734, n26735, n26736, n26737, n26738,
    n26739, n26740, n26741, n26742, n26743, n26744,
    n26745, n26746, n26747, n26748, n26749, n26750,
    n26751, n26752, n26753, n26754, n26755, n26756,
    n26757, n26758, n26759, n26760, n26761, n26762,
    n26763, n26764, n26765, n26766, n26767, n26768,
    n26769, n26770, n26771, n26772, n26773, n26774,
    n26775, n26776, n26777, n26778, n26779, n26780,
    n26781, n26782, n26783, n26784, n26785, n26786,
    n26787, n26788, n26789, n26790, n26791, n26792,
    n26793, n26794, n26795, n26796, n26797, n26798,
    n26799, n26800, n26801, n26802, n26803, n26804,
    n26805, n26806, n26807, n26808, n26809, n26810,
    n26811, n26812, n26813, n26814, n26815, n26816,
    n26817, n26818, n26819, n26820, n26821, n26822,
    n26823, n26824, n26825, n26826, n26827, n26828,
    n26829, n26830, n26831, n26832, n26833, n26834,
    n26835, n26836, n26837, n26838, n26839, n26840,
    n26841, n26842, n26843, n26844, n26845, n26846,
    n26847, n26848, n26849, n26850, n26851, n26852,
    n26853, n26854, n26855, n26856, n26857, n26858,
    n26859, n26860, n26861, n26862, n26863, n26864,
    n26865, n26866, n26867, n26868, n26869, n26870,
    n26871, n26872, n26873, n26874, n26875, n26876,
    n26877, n26878, n26879, n26880, n26881, n26882,
    n26883, n26884, n26885, n26886, n26887, n26888,
    n26889, n26890, n26891, n26892, n26893, n26894,
    n26895, n26896, n26897, n26898, n26899, n26900,
    n26901, n26902, n26903, n26904, n26905, n26906,
    n26907, n26908, n26909, n26910, n26911, n26912,
    n26913, n26914, n26915, n26916, n26917, n26918,
    n26919, n26920, n26921, n26922, n26923, n26924,
    n26925, n26926, n26927, n26928, n26929, n26930,
    n26931, n26932, n26933, n26934, n26935, n26936,
    n26937, n26938, n26939, n26940, n26941, n26942,
    n26943, n26944, n26945, n26946, n26947, n26948,
    n26949, n26950, n26951, n26952, n26953, n26954,
    n26955, n26956, n26957, n26958, n26959, n26960,
    n26961, n26962, n26963, n26964, n26965, n26966,
    n26967, n26968, n26969, n26970, n26971, n26972,
    n26973, n26974, n26975, n26976, n26977, n26978,
    n26979, n26980, n26981, n26982, n26983, n26984,
    n26985, n26986, n26987, n26988, n26989, n26990,
    n26991, n26992, n26993, n26994, n26995, n26996,
    n26997, n26998, n26999, n27000, n27001, n27002,
    n27003, n27004, n27005, n27006, n27007, n27008,
    n27009, n27010, n27011, n27012, n27013, n27014,
    n27015, n27016, n27017, n27018, n27019, n27020,
    n27021, n27022, n27023, n27024, n27025, n27026,
    n27027, n27028, n27029, n27030, n27031, n27032,
    n27033, n27034, n27035, n27036, n27037, n27038,
    n27039, n27040, n27041, n27042, n27043, n27044,
    n27045, n27046, n27047, n27048, n27049, n27050,
    n27051, n27052, n27053, n27054, n27055, n27056,
    n27057, n27058, n27059, n27060, n27061, n27062,
    n27063, n27064, n27065, n27066, n27067, n27068,
    n27069, n27070, n27071, n27072, n27073, n27074,
    n27075, n27076, n27077, n27078, n27079, n27080,
    n27081, n27082, n27083, n27084, n27085, n27086,
    n27087, n27088, n27089, n27090, n27091, n27092,
    n27093, n27094, n27095, n27096, n27097, n27098,
    n27099, n27100, n27101, n27102, n27103, n27104,
    n27105, n27106, n27107, n27108, n27109, n27110,
    n27111, n27112, n27113, n27114, n27115, n27116,
    n27117, n27118, n27119, n27120, n27121, n27122,
    n27123, n27124, n27125, n27126, n27127, n27128,
    n27129, n27130, n27131, n27132, n27133, n27134,
    n27135, n27136, n27137, n27138, n27139, n27140,
    n27141, n27142, n27143, n27144, n27145, n27146,
    n27147, n27148, n27149, n27150, n27151, n27152,
    n27153, n27154, n27155, n27156, n27157, n27158,
    n27159, n27160, n27161, n27162, n27163, n27164,
    n27165, n27166, n27167, n27168, n27169, n27170,
    n27171, n27172, n27173, n27174, n27175, n27176,
    n27177, n27178, n27179, n27180, n27181, n27182,
    n27183, n27184, n27185, n27186, n27187, n27188,
    n27189, n27190, n27191, n27192, n27193, n27194,
    n27195, n27196, n27197, n27198, n27199, n27200,
    n27201, n27202, n27203, n27204, n27205, n27206,
    n27207, n27208, n27209, n27210, n27211, n27212,
    n27213, n27214, n27215, n27216, n27217, n27218,
    n27219, n27220, n27221, n27222, n27223, n27224,
    n27225, n27226, n27227, n27228, n27229, n27230,
    n27231, n27232, n27233, n27234, n27235, n27236,
    n27237, n27238, n27239, n27240, n27241, n27242,
    n27243, n27244, n27245, n27246, n27247, n27248,
    n27249, n27250, n27251, n27252, n27253, n27254,
    n27255, n27256, n27257, n27258, n27259, n27260,
    n27261, n27262, n27263, n27264, n27265, n27266,
    n27267, n27268, n27269, n27270, n27271, n27272,
    n27273, n27274, n27275, n27276, n27277, n27278,
    n27279, n27280, n27281, n27282, n27283, n27284,
    n27285, n27286, n27287, n27288, n27289, n27290,
    n27291, n27292, n27293, n27294, n27295, n27296,
    n27297, n27298, n27299, n27300, n27301, n27302,
    n27303, n27304, n27305, n27306, n27307, n27308,
    n27309, n27310, n27311, n27312, n27313, n27314,
    n27315, n27316, n27317, n27318, n27319, n27320,
    n27321, n27322, n27323, n27324, n27325, n27326,
    n27327, n27328, n27329, n27330, n27331, n27332,
    n27333, n27334, n27335, n27336, n27337, n27338,
    n27339, n27340, n27341, n27342, n27343, n27344,
    n27345, n27346, n27347, n27348, n27349, n27350,
    n27351, n27352, n27353, n27354, n27355, n27356,
    n27357, n27358, n27359, n27360, n27361, n27362,
    n27363, n27364, n27365, n27366, n27367, n27368,
    n27369, n27370, n27371, n27372, n27373, n27374,
    n27375, n27376, n27377, n27378, n27379, n27380,
    n27381, n27382, n27383, n27384, n27385, n27386,
    n27387, n27388, n27389, n27390, n27391, n27392,
    n27393, n27394, n27395, n27396, n27397, n27398,
    n27399, n27400, n27401, n27402, n27403, n27404,
    n27405, n27406, n27407, n27408, n27409, n27410,
    n27411, n27412, n27413, n27414, n27415, n27416,
    n27417, n27418, n27419, n27420, n27421, n27422,
    n27423, n27424, n27425, n27426, n27427, n27428,
    n27429, n27430, n27431, n27432, n27433, n27434,
    n27435, n27436, n27437, n27438, n27439, n27440,
    n27441, n27442, n27443, n27444, n27445, n27446,
    n27447, n27448, n27449, n27450, n27451, n27452,
    n27453, n27454, n27455, n27456, n27457, n27458,
    n27459, n27460, n27461, n27462, n27463, n27464,
    n27465, n27466, n27467, n27468, n27469, n27470,
    n27471, n27472, n27473, n27474, n27475, n27476,
    n27477, n27478, n27479, n27480, n27481, n27482,
    n27483, n27484, n27485, n27486, n27487, n27488,
    n27489, n27490, n27491, n27492, n27493, n27494,
    n27495, n27496, n27497, n27498, n27499, n27500,
    n27501, n27502, n27503, n27504, n27505, n27506,
    n27507, n27508, n27509, n27510, n27511, n27512,
    n27513, n27514, n27515, n27516, n27517, n27518,
    n27519, n27520, n27521, n27522, n27523, n27524,
    n27525, n27526, n27527, n27528, n27529, n27530,
    n27531, n27532, n27533, n27534, n27535, n27536,
    n27537, n27538, n27539, n27540, n27541, n27542,
    n27543, n27544, n27545, n27546, n27547, n27548,
    n27549, n27550, n27551, n27552, n27553, n27554,
    n27555, n27556, n27557, n27558, n27559, n27560,
    n27561, n27562, n27563, n27564, n27565, n27566,
    n27567, n27568, n27569, n27570, n27571, n27572,
    n27573, n27574, n27575, n27576, n27577, n27578,
    n27579, n27580, n27581, n27582, n27583, n27584,
    n27585, n27586, n27587, n27588, n27589, n27590,
    n27591, n27592, n27593, n27594, n27595, n27596,
    n27597, n27598, n27599, n27600, n27601, n27602,
    n27603, n27604, n27605, n27606, n27607, n27608,
    n27609, n27610, n27611, n27612, n27613, n27614,
    n27615, n27616, n27617, n27618, n27619, n27620,
    n27621, n27622, n27623, n27624, n27625, n27626,
    n27627, n27628, n27629, n27630, n27631, n27632,
    n27633, n27634, n27635, n27636, n27637, n27638,
    n27639, n27640, n27641, n27642, n27643, n27644,
    n27645, n27646, n27647, n27648, n27649, n27650,
    n27651, n27652, n27653, n27654, n27655, n27656,
    n27657, n27658, n27659, n27660, n27661, n27662,
    n27663, n27664, n27665, n27666, n27667, n27668,
    n27669, n27670, n27671, n27672, n27673, n27674,
    n27675, n27676, n27677, n27678, n27679, n27680,
    n27681, n27682, n27683, n27684, n27685, n27686,
    n27687, n27688, n27689, n27690, n27691, n27692,
    n27693, n27694, n27695, n27696, n27697, n27698,
    n27699, n27700, n27701, n27702, n27703, n27704,
    n27705, n27706, n27707, n27708, n27709, n27710,
    n27711, n27712, n27713, n27714, n27715, n27716,
    n27717, n27718, n27719, n27720, n27721, n27722,
    n27723, n27724, n27725, n27726, n27727, n27728,
    n27729, n27730, n27731, n27732, n27733, n27734,
    n27735, n27736, n27737, n27738, n27739, n27740,
    n27741, n27742, n27743, n27744, n27745, n27746,
    n27747, n27748, n27749, n27750, n27751, n27752,
    n27753, n27754, n27755, n27756, n27757, n27758,
    n27759, n27760, n27761, n27762, n27763, n27764,
    n27765, n27766, n27767, n27768, n27769, n27770,
    n27771, n27772, n27773, n27774, n27775, n27776,
    n27777, n27778, n27779, n27780, n27781, n27782,
    n27783, n27784, n27785, n27786, n27787, n27788,
    n27789, n27790, n27791, n27792, n27793, n27794,
    n27795, n27796, n27797, n27798, n27799, n27800,
    n27801, n27802, n27803, n27804, n27805, n27806,
    n27807, n27808, n27809, n27810, n27811, n27812,
    n27813, n27814, n27815, n27816, n27817, n27818,
    n27819, n27820, n27821, n27822, n27823, n27824,
    n27825, n27826, n27827, n27828, n27829, n27830,
    n27831, n27832, n27833, n27834, n27835, n27836,
    n27837, n27838, n27839, n27840, n27841, n27842,
    n27843, n27844, n27845, n27846, n27847, n27848,
    n27849, n27850, n27851, n27852, n27853, n27854,
    n27855, n27856, n27857, n27858, n27859, n27860,
    n27861, n27862, n27863, n27864, n27865, n27866,
    n27867, n27868, n27869, n27870, n27871, n27872,
    n27873, n27874, n27875, n27876, n27877, n27878,
    n27879, n27880, n27881, n27882, n27883, n27884,
    n27885, n27886, n27887, n27888, n27889, n27890,
    n27891, n27892, n27893, n27894, n27895, n27896,
    n27897, n27898, n27899, n27900, n27901, n27902,
    n27903, n27904, n27905, n27906, n27907, n27908,
    n27909, n27910, n27911, n27912, n27913, n27914,
    n27915, n27916, n27917, n27918, n27919, n27920,
    n27921, n27922, n27923, n27924, n27925, n27926,
    n27927, n27928, n27929, n27930, n27931, n27932,
    n27933, n27934, n27935, n27936, n27937, n27938,
    n27939, n27940, n27941, n27942, n27943, n27944,
    n27945, n27946, n27947, n27948, n27949, n27950,
    n27951, n27952, n27953, n27954, n27955, n27956,
    n27957, n27958, n27959, n27960, n27961, n27962,
    n27963, n27964, n27965, n27966, n27967, n27968,
    n27969, n27970, n27971, n27972, n27973, n27974,
    n27975, n27976, n27977, n27978, n27979, n27980,
    n27981, n27982, n27983, n27984, n27985, n27986,
    n27987, n27988, n27989, n27990, n27991, n27992,
    n27993, n27994, n27995, n27996, n27997, n27998,
    n27999, n28000, n28001, n28002, n28003, n28004,
    n28005, n28006, n28007, n28008, n28009, n28010,
    n28011, n28012, n28013, n28014, n28015, n28016,
    n28017, n28018, n28019, n28020, n28021, n28022,
    n28023, n28024, n28025, n28026, n28027, n28028,
    n28029, n28030, n28031, n28032, n28033, n28034,
    n28035, n28036, n28037, n28038, n28039, n28040,
    n28041, n28042, n28043, n28044, n28045, n28046,
    n28047, n28048, n28049, n28050, n28051, n28052,
    n28053, n28054, n28055, n28056, n28057, n28058,
    n28059, n28060, n28061, n28062, n28063, n28064,
    n28065, n28066, n28067, n28068, n28069, n28070,
    n28071, n28072, n28073, n28074, n28075, n28076,
    n28077, n28078, n28079, n28080, n28081, n28082,
    n28083, n28084, n28085, n28086, n28087, n28088,
    n28089, n28090, n28091, n28092, n28093, n28094,
    n28095, n28096, n28097, n28098, n28099, n28100,
    n28101, n28102, n28103, n28104, n28105, n28106,
    n28107, n28108, n28109, n28110, n28111, n28112,
    n28113, n28114, n28115, n28116, n28117, n28118,
    n28119, n28120, n28121, n28122, n28123, n28124,
    n28125, n28126, n28127, n28128, n28129, n28130,
    n28131, n28132, n28133, n28134, n28135, n28136,
    n28137, n28138, n28139, n28140, n28141, n28142,
    n28143, n28144, n28145, n28146, n28147, n28148,
    n28149, n28150, n28151, n28152, n28153, n28154,
    n28155, n28156, n28157, n28158, n28159, n28160,
    n28161, n28162, n28163, n28164, n28165, n28166,
    n28167, n28168, n28169, n28170, n28171, n28172,
    n28173, n28174, n28175, n28176, n28177, n28178,
    n28179, n28180, n28181, n28182, n28183, n28184,
    n28185, n28186, n28187, n28188, n28189, n28190,
    n28191, n28192, n28193, n28194, n28195, n28196,
    n28197, n28198, n28199, n28200, n28201, n28202,
    n28203, n28204, n28205, n28206, n28207, n28208,
    n28209, n28210, n28211, n28212, n28213, n28214,
    n28215, n28216, n28217, n28218, n28219, n28220,
    n28221, n28222, n28223, n28224, n28225, n28226,
    n28227, n28228, n28229, n28230, n28231, n28232,
    n28233, n28234, n28235, n28236, n28237, n28238,
    n28239, n28240, n28241, n28242, n28243, n28244,
    n28245, n28246, n28247, n28248, n28249, n28250,
    n28251, n28252, n28253, n28254, n28255, n28256,
    n28257, n28258, n28259, n28260, n28261, n28262,
    n28263, n28264, n28265, n28266, n28267, n28268,
    n28269, n28270, n28271, n28272, n28273, n28274,
    n28275, n28276, n28277, n28278, n28279, n28280,
    n28281, n28282, n28283, n28284, n28285, n28286,
    n28287, n28288, n28289, n28290, n28291, n28292,
    n28293, n28294, n28295, n28296, n28297, n28298,
    n28299, n28300, n28301, n28302, n28303, n28304,
    n28305, n28306, n28307, n28308, n28309, n28310,
    n28311, n28312, n28313, n28314, n28315, n28316,
    n28317, n28318, n28319, n28320, n28321, n28322,
    n28323, n28324, n28325, n28326, n28327, n28328,
    n28329, n28330, n28331, n28332, n28333, n28334,
    n28335, n28336, n28337, n28338, n28339, n28340,
    n28341, n28342, n28343, n28344, n28345, n28346,
    n28347, n28348, n28349, n28350, n28351, n28352,
    n28353, n28354, n28355, n28356, n28357, n28358,
    n28359, n28360, n28361, n28362, n28363, n28364,
    n28365, n28366, n28367, n28368, n28369, n28370,
    n28371, n28372, n28373, n28374, n28375, n28376,
    n28377, n28378, n28379, n28380, n28381, n28382,
    n28383, n28384, n28385, n28386, n28387, n28388,
    n28389, n28390, n28391, n28392, n28393, n28394,
    n28395, n28396, n28397, n28398, n28399, n28400,
    n28401, n28402, n28403, n28404, n28405, n28406,
    n28407, n28408, n28409, n28410, n28411, n28412,
    n28413, n28414, n28415, n28416, n28417, n28418,
    n28419, n28420, n28421, n28422, n28423, n28424,
    n28425, n28426, n28427, n28428, n28429, n28430,
    n28431, n28432, n28433, n28434, n28435, n28436,
    n28437, n28438, n28439, n28440, n28441, n28442,
    n28443, n28444, n28445, n28446, n28447, n28448,
    n28449, n28450, n28451, n28452, n28453, n28454,
    n28455, n28456, n28457, n28458, n28459, n28460,
    n28461, n28462, n28463, n28464, n28465, n28466,
    n28467, n28468, n28469, n28470, n28471, n28472,
    n28473, n28474, n28475, n28476, n28477, n28478,
    n28479, n28480, n28481, n28482, n28483, n28484,
    n28485, n28486, n28487, n28488, n28489, n28490,
    n28491, n28492, n28493, n28494, n28495, n28496,
    n28497, n28498, n28499, n28500, n28501, n28502,
    n28503, n28504, n28505, n28506, n28507, n28508,
    n28509, n28510, n28511, n28512, n28513, n28514,
    n28515, n28516, n28517, n28518, n28519, n28520,
    n28521, n28522, n28523, n28524, n28525, n28526,
    n28527, n28528, n28529, n28530, n28531, n28532,
    n28533, n28534, n28535, n28536, n28537, n28538,
    n28539, n28540, n28541, n28542, n28543, n28544,
    n28545, n28546, n28547, n28548, n28549, n28550,
    n28551, n28552, n28553, n28554, n28555, n28556,
    n28557, n28558, n28559, n28560, n28561, n28562,
    n28563, n28564, n28565, n28566, n28567, n28568,
    n28569, n28570, n28571, n28572, n28573, n28574,
    n28575, n28576, n28577, n28578, n28579, n28580,
    n28581, n28582, n28583, n28584, n28585, n28586,
    n28587, n28588, n28589, n28590, n28591, n28592,
    n28593, n28594, n28595, n28596, n28597, n28598,
    n28599, n28600, n28601, n28602, n28603, n28604,
    n28605, n28606, n28607, n28608, n28609, n28610,
    n28611, n28612, n28613, n28614, n28615, n28616,
    n28617, n28618, n28619, n28620, n28621, n28622,
    n28623, n28624, n28625, n28626, n28627, n28628,
    n28629, n28630, n28631, n28632, n28633, n28634,
    n28635, n28636, n28637, n28638, n28639, n28640,
    n28641, n28642, n28643, n28644, n28645, n28646,
    n28647, n28648, n28649, n28650, n28651, n28652,
    n28653, n28654, n28655, n28656, n28657, n28658,
    n28659, n28660, n28661, n28662, n28663, n28664,
    n28665, n28666, n28667, n28668, n28669, n28670,
    n28671, n28672, n28673, n28674, n28675, n28676,
    n28677, n28678, n28679, n28680, n28681, n28682,
    n28683, n28684, n28685, n28686, n28687, n28688,
    n28689, n28690, n28691, n28692, n28693, n28694,
    n28695, n28696, n28697, n28698, n28699, n28700,
    n28701, n28702, n28703, n28704, n28705, n28706,
    n28707, n28708, n28709, n28710, n28711, n28712,
    n28713, n28714, n28715, n28716, n28717, n28718,
    n28719, n28720, n28721, n28722, n28723, n28724,
    n28725, n28726, n28727, n28728, n28729, n28730,
    n28731, n28732, n28733, n28734, n28735, n28736,
    n28737, n28738, n28739, n28740, n28741, n28742,
    n28743, n28744, n28745, n28746, n28747, n28748,
    n28749, n28750, n28751, n28752, n28753, n28754,
    n28755, n28756, n28757, n28758, n28759, n28760,
    n28761, n28762, n28763, n28764, n28765, n28766,
    n28767, n28768, n28769, n28770, n28771, n28772,
    n28773, n28774, n28775, n28776, n28777, n28778,
    n28779, n28780, n28781, n28782, n28783, n28784,
    n28785, n28786, n28787, n28788, n28789, n28790,
    n28791, n28792, n28793, n28794, n28795, n28796,
    n28797, n28798, n28799, n28800, n28801, n28802,
    n28803, n28804, n28805, n28806, n28807, n28808,
    n28809, n28810, n28811, n28812, n28813, n28814,
    n28815, n28816, n28817, n28818, n28819, n28820,
    n28821, n28822, n28823, n28824, n28825, n28826,
    n28827, n28828, n28829, n28830, n28831, n28832,
    n28833, n28834, n28835, n28836, n28837, n28838,
    n28839, n28840, n28841, n28842, n28843, n28844,
    n28845, n28846, n28847, n28848, n28849, n28850,
    n28851, n28852, n28853, n28854, n28855, n28856,
    n28857, n28858, n28859, n28860, n28861, n28862,
    n28863, n28864, n28865, n28866, n28867, n28868,
    n28869, n28870, n28871, n28872, n28873, n28874,
    n28875, n28876, n28877, n28878, n28879, n28880,
    n28881, n28882, n28883, n28884, n28885, n28886,
    n28887, n28888, n28889, n28890, n28891, n28892,
    n28893, n28894, n28895, n28896, n28897, n28898,
    n28899, n28900, n28901, n28902, n28903, n28904,
    n28905, n28906, n28907, n28908, n28909, n28910,
    n28911, n28912, n28913, n28914, n28915, n28916,
    n28917, n28918, n28919, n28920, n28921, n28922,
    n28923, n28924, n28925, n28926, n28927, n28928,
    n28929, n28930, n28931, n28932, n28933, n28934,
    n28935, n28936, n28937, n28938, n28939, n28940,
    n28941, n28942, n28943, n28944, n28945, n28946,
    n28947, n28948, n28949, n28950, n28951, n28952,
    n28953, n28954, n28955, n28956, n28957, n28958,
    n28959, n28960, n28961, n28962, n28963, n28964,
    n28965, n28966, n28967, n28968, n28969, n28970,
    n28971, n28972, n28973, n28974, n28975, n28976,
    n28977, n28978, n28979, n28980, n28981, n28982,
    n28983, n28984, n28985, n28986, n28987, n28988,
    n28989, n28990, n28991, n28992, n28993, n28994,
    n28995, n28996, n28997, n28998, n28999, n29000,
    n29001, n29002, n29003, n29004, n29005, n29006,
    n29007, n29008, n29009, n29010, n29011, n29012,
    n29013, n29014, n29015, n29016, n29017, n29018,
    n29019, n29020, n29021, n29022, n29023, n29024,
    n29025, n29026, n29027, n29028, n29029, n29030,
    n29031, n29032, n29033, n29034, n29035, n29036,
    n29037, n29038, n29039, n29040, n29041, n29042,
    n29043, n29044, n29045, n29046, n29047, n29048,
    n29049, n29050, n29051, n29052, n29053, n29054,
    n29055, n29056, n29057, n29058, n29059, n29060,
    n29061, n29062, n29063, n29064, n29065, n29066,
    n29067, n29068, n29069, n29070, n29071, n29072,
    n29073, n29074, n29075, n29076, n29077, n29078,
    n29079, n29080, n29081, n29082, n29083, n29084,
    n29085, n29086, n29087, n29088, n29089, n29090,
    n29091, n29092, n29093, n29094, n29095, n29096,
    n29097, n29098, n29099, n29100, n29101, n29102,
    n29103, n29104, n29105, n29106, n29107, n29108,
    n29109, n29110, n29111, n29112, n29113, n29114,
    n29115, n29116, n29117, n29118, n29119, n29120,
    n29121, n29122, n29123, n29124, n29125, n29126,
    n29127, n29128, n29129, n29130, n29131, n29132,
    n29133, n29134, n29135, n29136, n29137, n29138,
    n29139, n29140, n29141, n29142, n29143, n29144,
    n29145, n29146, n29147, n29148, n29149, n29150,
    n29151, n29152, n29153, n29154, n29155, n29156,
    n29157, n29158, n29159, n29160, n29161, n29162,
    n29163, n29164, n29165, n29166, n29167, n29168,
    n29169, n29170, n29171, n29172, n29173, n29174,
    n29175, n29176, n29177, n29178, n29179, n29180,
    n29181, n29182, n29183, n29184, n29185, n29186,
    n29187, n29188, n29189, n29190, n29191, n29192,
    n29193, n29194, n29195, n29196, n29197, n29198,
    n29199, n29200, n29201, n29202, n29203, n29204,
    n29205, n29206, n29207, n29208, n29209, n29210,
    n29211, n29212, n29213, n29214, n29215, n29216,
    n29217, n29218, n29219, n29220, n29221, n29222,
    n29223, n29224, n29225, n29226, n29227, n29228,
    n29229, n29230, n29231, n29232, n29233, n29234,
    n29235, n29236, n29237, n29238, n29239, n29240,
    n29241, n29242, n29243, n29244, n29245, n29246,
    n29247, n29248, n29249, n29250, n29251, n29252,
    n29253, n29254, n29255, n29256, n29257, n29258,
    n29259, n29260, n29261, n29262, n29263, n29264,
    n29265, n29266, n29267, n29268, n29269, n29270,
    n29271, n29272, n29273, n29274, n29275, n29276,
    n29277, n29278, n29279, n29280, n29281, n29282,
    n29283, n29284, n29285, n29286, n29287, n29288,
    n29289, n29290, n29291, n29292, n29293, n29294,
    n29295, n29296, n29297, n29298, n29299, n29300,
    n29301, n29302, n29303, n29304, n29305, n29306,
    n29307, n29308, n29309, n29310, n29311, n29312,
    n29313, n29314, n29315, n29316, n29317, n29318,
    n29319, n29320, n29321, n29322, n29323, n29324,
    n29325, n29326, n29327, n29328, n29329, n29330,
    n29331, n29332, n29333, n29334, n29335, n29336,
    n29337, n29338, n29339, n29340, n29341, n29342,
    n29343, n29344, n29345, n29346, n29347, n29348,
    n29349, n29350, n29351, n29352, n29353, n29354,
    n29355, n29356, n29357, n29358, n29359, n29360,
    n29361, n29362, n29363, n29364, n29365, n29366,
    n29367, n29368, n29369, n29370, n29371, n29372,
    n29373, n29374, n29375, n29376, n29377, n29378,
    n29379, n29380, n29381, n29382, n29383, n29384,
    n29385, n29386, n29387, n29388, n29389, n29390,
    n29391, n29392, n29393, n29394, n29395, n29396,
    n29397, n29398, n29399, n29400, n29401, n29402,
    n29403, n29404, n29405, n29406, n29407, n29408,
    n29409, n29410, n29411, n29412, n29413, n29414,
    n29415, n29416, n29417, n29418, n29419, n29420,
    n29421, n29422, n29423, n29424, n29425, n29426,
    n29427, n29428, n29429, n29430, n29431, n29432,
    n29433, n29434, n29435, n29436, n29437, n29438,
    n29439, n29440, n29441, n29442, n29443, n29444,
    n29445, n29446, n29447, n29448, n29449, n29450,
    n29451, n29452, n29453, n29454, n29455, n29456,
    n29457, n29458, n29459, n29460, n29461, n29462,
    n29463, n29464, n29465, n29466, n29467, n29468,
    n29469, n29470, n29471, n29472, n29473, n29474,
    n29475, n29476, n29477, n29478, n29479, n29480,
    n29481, n29482, n29483, n29484, n29485, n29486,
    n29487, n29488, n29489, n29490, n29491, n29492,
    n29493, n29494, n29495, n29496, n29497, n29498,
    n29499, n29500, n29501, n29502, n29503, n29504,
    n29505, n29506, n29507, n29508, n29509, n29510,
    n29511, n29512, n29513, n29514, n29515, n29516,
    n29517, n29518, n29519, n29520, n29521, n29522,
    n29523, n29524, n29525, n29526, n29527, n29528,
    n29529, n29530, n29531, n29532, n29533, n29534,
    n29535, n29536, n29537, n29538, n29539, n29540,
    n29541, n29542, n29543, n29544, n29545, n29546,
    n29547, n29548, n29549, n29550, n29551, n29552,
    n29553, n29554, n29555, n29556, n29557, n29558,
    n29559, n29560, n29561, n29562, n29563, n29564,
    n29565, n29566, n29567, n29568, n29569, n29570,
    n29571, n29572, n29573, n29574, n29575, n29576,
    n29577, n29578, n29579, n29580, n29581, n29582,
    n29583, n29584, n29585, n29586, n29587, n29588,
    n29589, n29590, n29591, n29592, n29593, n29594,
    n29595, n29596, n29597, n29598, n29599, n29600,
    n29601, n29602, n29603, n29604, n29605, n29606,
    n29607, n29608, n29609, n29610, n29611, n29612,
    n29613, n29614, n29615, n29616, n29617, n29618,
    n29619, n29620, n29621, n29622, n29623, n29624,
    n29625, n29626, n29627, n29628, n29629, n29630,
    n29631, n29632, n29633, n29634, n29635, n29636,
    n29637, n29638, n29639, n29640, n29641, n29642,
    n29643, n29644, n29645, n29646, n29647, n29648,
    n29649, n29650, n29651, n29652, n29653, n29654,
    n29655, n29656, n29657, n29658, n29659, n29660,
    n29661, n29662, n29663, n29664, n29665, n29666,
    n29667, n29668, n29669, n29670, n29671, n29672,
    n29673, n29674, n29675, n29676, n29677, n29678,
    n29679, n29680, n29681, n29682, n29683, n29684,
    n29685, n29686, n29687, n29688, n29689, n29690,
    n29691, n29692, n29693, n29694, n29695, n29696,
    n29697, n29698, n29699, n29700, n29701, n29702,
    n29703, n29704, n29705, n29706, n29707, n29708,
    n29709, n29710, n29711, n29712, n29713, n29714,
    n29715, n29716, n29717, n29718, n29719, n29720,
    n29721, n29722, n29723, n29724, n29725, n29726,
    n29727, n29728, n29729, n29730, n29731, n29732,
    n29733, n29734, n29735, n29736, n29737, n29738,
    n29739, n29740, n29741, n29742, n29743, n29744,
    n29745, n29746, n29747, n29748, n29749, n29750,
    n29751, n29752, n29753, n29754, n29755, n29756,
    n29757, n29758, n29759, n29760, n29761, n29762,
    n29763, n29764, n29765, n29766, n29767, n29768,
    n29769, n29770, n29771, n29772, n29773, n29774,
    n29775, n29776, n29777, n29778, n29779, n29780,
    n29781, n29782, n29783, n29784, n29785, n29786,
    n29787, n29788, n29789, n29790, n29791, n29792,
    n29793, n29794, n29795, n29796, n29797, n29798,
    n29799, n29800, n29801, n29802, n29803, n29804,
    n29805, n29806, n29807, n29808, n29809, n29810,
    n29811, n29812, n29813, n29814, n29815, n29816,
    n29817, n29818, n29819, n29820, n29821, n29822,
    n29823, n29824, n29825, n29826, n29827, n29828,
    n29829, n29830, n29831, n29832, n29833, n29834,
    n29835, n29836, n29837, n29838, n29839, n29840,
    n29841, n29842, n29843, n29844, n29845, n29846,
    n29847, n29848, n29849, n29850, n29851, n29852,
    n29853, n29854, n29855, n29856, n29857, n29858,
    n29859, n29860, n29861, n29862, n29863, n29864,
    n29865, n29866, n29867, n29868, n29869, n29870,
    n29871, n29872, n29873, n29874, n29875, n29876,
    n29877, n29878, n29879, n29880, n29881, n29882,
    n29883, n29884, n29885, n29886, n29887, n29888,
    n29889, n29890, n29891, n29892, n29893, n29894,
    n29895, n29896, n29897, n29898, n29899, n29900,
    n29901, n29902, n29903, n29904, n29905, n29906,
    n29907, n29908, n29909, n29910, n29911, n29912,
    n29913, n29914, n29915, n29916, n29917, n29918,
    n29919, n29920, n29921, n29922, n29923, n29924,
    n29925, n29926, n29927, n29928, n29929, n29930,
    n29931, n29932, n29933, n29934, n29935, n29936,
    n29937, n29938, n29939, n29940, n29941, n29942,
    n29943, n29944, n29945, n29946, n29947, n29948,
    n29949, n29950, n29951, n29952, n29953, n29954,
    n29955, n29956, n29957, n29958, n29959, n29960,
    n29961, n29962, n29963, n29964, n29965, n29966,
    n29967, n29968, n29969, n29970, n29971, n29972,
    n29973, n29974, n29975, n29976, n29977, n29978,
    n29979, n29980, n29981, n29982, n29983, n29984,
    n29985, n29986, n29987, n29988, n29989, n29990,
    n29991, n29992, n29993, n29994, n29995, n29996,
    n29997, n29998, n29999, n30000, n30001, n30002,
    n30003, n30004, n30005, n30006, n30007, n30008,
    n30009, n30010, n30011, n30012, n30013, n30014,
    n30015, n30016, n30017, n30018, n30019, n30020,
    n30021, n30022, n30023, n30024, n30025, n30026,
    n30027, n30028, n30029, n30030, n30031, n30032,
    n30033, n30034, n30035, n30036, n30037, n30038,
    n30039, n30040, n30041, n30042, n30043, n30044,
    n30045, n30046, n30047, n30048, n30049, n30050,
    n30051, n30052, n30053, n30054, n30055, n30056,
    n30057, n30058, n30059, n30060, n30061, n30062,
    n30063, n30064, n30065, n30066, n30067, n30068,
    n30069, n30070, n30071, n30072, n30073, n30074,
    n30075, n30076, n30077, n30078, n30079, n30080,
    n30081, n30082, n30083, n30084, n30085, n30086,
    n30087, n30088, n30089, n30090, n30091, n30092,
    n30093, n30094, n30095, n30096, n30097, n30098,
    n30099, n30100, n30101, n30102, n30103, n30104,
    n30105, n30106, n30107, n30108, n30109, n30110,
    n30111, n30112, n30113, n30114, n30115, n30116,
    n30117, n30118, n30119, n30120, n30121, n30122,
    n30123, n30124, n30125, n30126, n30127, n30128,
    n30129, n30130, n30131, n30132, n30133, n30134,
    n30135, n30136, n30137, n30138, n30139, n30140,
    n30141, n30142, n30143, n30144, n30145, n30146,
    n30147, n30148, n30149, n30150, n30151, n30152,
    n30153, n30154, n30155, n30156, n30157, n30158,
    n30159, n30160, n30161, n30162, n30163, n30164,
    n30165, n30166, n30167, n30168, n30169, n30170,
    n30171, n30172, n30173, n30174, n30175, n30176,
    n30177, n30178, n30179, n30180, n30181, n30182,
    n30183, n30184, n30185, n30186, n30187, n30188,
    n30189, n30190, n30191, n30192, n30193, n30194,
    n30195, n30196, n30197, n30198, n30199, n30200,
    n30201, n30202, n30203, n30204, n30205, n30206,
    n30207, n30208, n30209, n30210, n30211, n30212,
    n30213, n30214, n30215, n30216, n30217, n30218,
    n30219, n30220, n30221, n30222, n30223, n30224,
    n30225, n30226, n30227, n30228, n30229, n30230,
    n30231, n30232, n30233, n30234, n30235, n30236,
    n30237, n30238, n30239, n30240, n30241, n30242,
    n30243, n30244, n30245, n30246, n30247, n30248,
    n30249, n30250, n30251, n30252, n30253, n30254,
    n30255, n30256, n30257, n30258, n30259, n30260,
    n30261, n30262, n30263, n30264, n30265, n30266,
    n30267, n30268, n30269, n30270, n30271, n30272,
    n30273, n30274, n30275, n30276, n30277, n30278,
    n30279, n30280, n30281, n30282, n30283, n30284,
    n30285, n30286, n30287, n30288, n30289, n30290,
    n30291, n30292, n30293, n30294, n30295, n30296,
    n30297, n30298, n30299, n30300, n30301, n30302,
    n30303, n30304, n30305, n30306, n30307, n30308,
    n30309, n30310, n30311, n30312, n30313, n30314,
    n30315, n30316, n30317, n30318, n30319, n30320,
    n30321, n30322, n30323, n30324, n30325, n30326,
    n30327, n30328, n30329, n30330, n30331, n30332,
    n30333, n30334, n30335, n30336, n30337, n30338,
    n30339, n30340, n30341, n30342, n30343, n30344,
    n30345, n30346, n30347, n30348, n30349, n30350,
    n30351, n30352, n30353, n30354, n30355, n30356,
    n30357, n30358, n30359, n30360, n30361, n30362,
    n30363, n30364, n30365, n30366, n30367, n30368,
    n30369, n30370, n30371, n30372, n30373, n30374,
    n30375, n30376, n30377, n30378, n30379, n30380,
    n30381, n30382, n30383, n30384, n30385, n30386,
    n30387, n30388, n30389, n30390, n30391, n30392,
    n30393, n30394, n30395, n30396, n30397, n30398,
    n30399, n30400, n30401, n30402, n30403, n30404,
    n30405, n30406, n30407, n30408, n30409, n30410,
    n30411, n30412, n30413, n30414, n30415, n30416,
    n30417, n30418, n30419, n30420, n30421, n30422,
    n30423, n30424, n30425, n30426, n30427, n30428,
    n30429, n30430, n30431, n30432, n30433, n30434,
    n30435, n30436, n30437, n30438, n30439, n30440,
    n30441, n30442, n30443, n30444, n30445, n30446,
    n30447, n30448, n30449, n30450, n30451, n30452,
    n30453, n30454, n30455, n30456, n30457, n30458,
    n30459, n30460, n30461, n30462, n30463, n30464,
    n30465, n30466, n30467, n30468, n30469, n30470,
    n30471, n30472, n30473, n30474, n30475, n30476,
    n30477, n30478, n30479, n30480, n30481, n30482,
    n30483, n30484, n30485, n30486, n30487, n30488,
    n30489, n30490, n30491, n30492, n30493, n30494,
    n30495, n30496, n30497, n30498, n30499, n30500,
    n30501, n30502, n30503, n30504, n30505, n30506,
    n30507, n30508, n30509, n30510, n30511, n30512,
    n30513, n30514, n30515, n30516, n30517, n30518,
    n30519, n30520, n30521, n30522, n30523, n30524,
    n30525, n30526, n30527, n30528, n30529, n30530,
    n30531, n30532, n30533, n30534, n30535, n30536,
    n30537, n30538, n30539, n30540, n30541, n30542,
    n30543, n30544, n30545, n30546, n30547, n30548,
    n30549, n30550, n30551, n30552, n30553, n30554,
    n30555, n30556, n30557, n30558, n30559, n30560,
    n30561, n30562, n30563, n30564, n30565, n30566,
    n30567, n30568, n30569, n30570, n30571, n30572,
    n30573, n30574, n30575, n30576, n30577, n30578,
    n30579, n30580, n30581, n30582, n30583, n30584,
    n30585, n30586, n30587, n30588, n30589, n30590,
    n30591, n30592, n30593, n30594, n30595, n30596,
    n30597, n30598, n30599, n30600, n30601, n30602,
    n30603, n30604, n30605, n30606, n30607, n30608,
    n30609, n30610, n30611, n30612, n30613, n30614,
    n30615, n30616, n30617, n30618, n30619, n30620,
    n30621, n30622, n30623, n30624, n30625, n30626,
    n30627, n30628, n30629, n30630, n30631, n30632,
    n30633, n30634, n30635, n30636, n30637, n30638,
    n30639, n30640, n30641, n30642, n30643, n30644,
    n30645, n30646, n30647, n30648, n30649, n30650,
    n30651, n30652, n30653, n30654, n30655, n30656,
    n30657, n30658, n30659, n30660, n30661, n30662,
    n30663, n30664, n30665, n30666, n30667, n30668,
    n30669, n30670, n30671, n30672, n30673, n30674,
    n30675, n30676, n30677, n30678, n30679, n30680,
    n30681, n30682, n30683, n30684, n30685, n30686,
    n30687, n30688, n30689, n30690, n30691, n30692,
    n30693, n30694, n30695, n30696, n30697, n30698,
    n30699, n30700, n30701, n30702, n30703, n30704,
    n30705, n30706, n30707, n30708, n30709, n30710,
    n30711, n30712, n30713, n30714, n30715, n30716,
    n30717, n30718, n30719, n30720, n30721, n30722,
    n30723, n30724, n30725, n30726, n30727, n30728,
    n30729, n30730, n30731, n30732, n30733, n30734,
    n30735, n30736, n30737, n30738, n30739, n30740,
    n30741, n30742, n30743, n30744, n30745, n30746,
    n30747, n30748, n30749, n30750, n30751, n30752,
    n30753, n30754, n30755, n30756, n30757, n30758,
    n30759, n30760, n30761, n30762, n30763, n30764,
    n30765, n30766, n30767, n30768, n30769, n30770,
    n30771, n30772, n30773, n30774, n30775, n30776,
    n30777, n30778, n30779, n30780, n30781, n30782,
    n30783, n30784, n30785, n30786, n30787, n30788,
    n30789, n30790, n30791, n30792, n30793, n30794,
    n30795, n30796, n30797, n30798, n30799, n30800,
    n30801, n30802, n30803, n30804, n30805, n30806,
    n30807, n30808, n30809, n30810, n30811, n30812,
    n30813, n30814, n30815, n30816, n30817, n30818,
    n30819, n30820, n30821, n30822, n30823, n30824,
    n30825, n30826, n30827, n30828, n30829, n30830,
    n30831, n30832, n30833, n30834, n30835, n30836,
    n30837, n30838, n30839, n30840, n30841, n30842,
    n30843, n30844, n30845, n30846, n30847, n30848,
    n30849, n30850, n30851, n30852, n30853, n30854,
    n30855, n30856, n30857, n30858, n30859, n30860,
    n30861, n30862, n30863, n30864, n30865, n30866,
    n30867, n30868, n30869, n30870, n30871, n30872,
    n30873, n30874, n30875, n30876, n30877, n30878,
    n30879, n30880, n30881, n30882, n30883, n30884,
    n30885, n30886, n30887, n30888, n30889, n30890,
    n30891, n30892, n30893, n30894, n30895, n30896,
    n30897, n30898, n30899, n30900, n30901, n30902,
    n30903, n30904, n30905, n30906, n30907, n30908,
    n30909, n30910, n30911, n30912, n30913, n30914,
    n30915, n30916, n30917, n30918, n30919, n30920,
    n30921, n30922, n30923, n30924, n30925, n30926,
    n30927, n30928, n30929, n30930, n30931, n30932,
    n30933, n30934, n30935, n30936, n30937, n30938,
    n30939, n30940, n30941, n30942, n30943, n30944,
    n30945, n30946, n30947, n30948, n30949, n30950,
    n30951, n30952, n30953, n30954, n30955, n30956,
    n30957, n30958, n30959, n30960, n30961, n30962,
    n30963, n30964, n30965, n30966, n30967, n30968,
    n30969, n30970, n30971, n30972, n30973, n30974,
    n30975, n30976, n30977, n30978, n30979, n30980,
    n30981, n30982, n30983, n30984, n30985, n30986,
    n30987, n30988, n30989, n30990, n30991, n30992,
    n30993, n30994, n30995, n30996, n30997, n30998,
    n30999, n31000, n31001, n31002, n31003, n31004,
    n31005, n31006, n31007, n31008, n31009, n31010,
    n31011, n31012, n31013, n31014, n31015, n31016,
    n31017, n31018, n31019, n31020, n31021, n31022,
    n31023, n31024, n31025, n31026, n31027, n31028,
    n31029, n31030, n31031, n31032, n31033, n31034,
    n31035, n31036, n31037, n31038, n31039, n31040,
    n31041, n31042, n31043, n31044, n31045, n31046,
    n31047, n31048, n31049, n31050, n31051, n31052,
    n31053, n31054, n31055, n31056, n31057, n31058,
    n31059, n31060, n31061, n31062, n31063, n31064,
    n31065, n31066, n31067, n31068, n31069, n31070,
    n31071, n31072, n31073, n31074, n31075, n31076,
    n31077, n31078, n31079, n31080, n31081, n31082,
    n31083, n31084, n31085, n31086, n31087, n31088,
    n31089, n31090, n31091, n31092, n31093, n31094,
    n31095, n31096, n31097, n31098, n31099, n31100,
    n31101, n31102, n31103, n31104, n31105, n31106,
    n31107, n31108, n31109, n31110, n31111, n31112,
    n31113, n31114, n31115, n31116, n31117, n31118,
    n31119, n31120, n31121, n31122, n31123, n31124,
    n31125, n31126, n31127, n31128, n31129, n31130,
    n31131, n31132, n31133, n31134, n31135, n31136,
    n31137, n31138, n31139, n31140, n31141, n31142,
    n31143, n31144, n31145, n31146, n31147, n31148,
    n31149, n31150, n31151, n31152, n31153, n31154,
    n31155, n31156, n31157, n31158, n31159, n31160,
    n31161, n31162, n31163, n31164, n31165, n31166,
    n31167, n31168, n31169, n31170, n31171, n31172,
    n31173, n31174, n31175, n31176, n31177, n31178,
    n31179, n31180, n31181, n31182, n31183, n31184,
    n31185, n31186, n31187, n31188, n31189, n31190,
    n31191, n31192, n31193, n31194, n31195, n31196,
    n31197, n31198, n31199, n31200, n31201, n31202,
    n31203, n31204, n31205, n31206, n31207, n31208,
    n31209, n31210, n31211, n31212, n31213, n31214,
    n31215, n31216, n31217, n31218, n31219, n31220,
    n31221, n31222, n31223, n31224, n31225, n31226,
    n31227, n31228, n31229, n31230, n31231, n31232,
    n31233, n31234, n31235, n31236, n31237, n31238,
    n31239, n31240, n31241, n31242, n31243, n31244,
    n31245, n31246, n31247, n31248, n31249, n31250,
    n31251, n31252, n31253, n31254, n31255, n31256,
    n31257, n31258, n31259, n31260, n31261, n31262,
    n31263, n31264, n31265, n31266, n31267, n31268,
    n31269, n31270, n31271, n31272, n31273, n31274,
    n31275, n31276, n31277, n31278, n31279, n31280,
    n31281, n31282, n31283, n31284, n31285, n31286,
    n31287, n31288, n31289, n31290, n31291, n31292,
    n31293, n31294, n31295, n31296, n31297, n31298,
    n31299, n31300, n31301, n31302, n31303, n31304,
    n31305, n31306, n31307, n31308, n31309, n31310,
    n31311, n31312, n31313, n31314, n31315, n31316,
    n31317, n31318, n31319, n31320, n31321, n31322,
    n31323, n31324, n31325, n31326, n31327, n31328,
    n31329, n31330, n31331, n31332, n31333, n31334,
    n31335, n31336, n31337, n31338, n31339, n31340,
    n31341, n31342, n31343, n31344, n31345, n31346,
    n31347, n31348, n31349, n31350, n31351, n31352,
    n31353, n31354, n31355, n31356, n31357, n31358,
    n31359, n31360, n31361, n31362, n31363, n31364,
    n31365, n31366, n31367, n31368, n31369, n31370,
    n31371, n31372, n31373, n31374, n31375, n31376,
    n31377, n31378, n31379, n31380, n31381, n31382,
    n31383, n31384, n31385, n31386, n31387, n31388,
    n31389, n31390, n31391, n31392, n31393, n31394,
    n31395, n31396, n31397, n31398, n31399, n31400,
    n31401, n31402, n31403, n31404, n31405, n31406,
    n31407, n31408, n31409, n31410, n31411, n31412,
    n31413, n31414, n31415, n31416, n31417, n31418,
    n31419, n31420, n31421, n31422, n31423, n31424,
    n31425, n31426, n31427, n31428, n31429, n31430,
    n31431, n31432, n31433, n31434, n31435, n31436,
    n31437, n31438, n31439, n31440, n31441, n31442,
    n31443, n31444, n31445, n31446, n31447, n31448,
    n31449, n31450, n31451, n31452, n31453, n31454,
    n31455, n31456, n31457, n31458, n31459, n31460,
    n31461, n31462, n31463, n31464, n31465, n31466,
    n31467, n31468, n31469, n31470, n31471, n31472,
    n31473, n31474, n31475, n31476, n31477, n31478,
    n31479, n31480, n31481, n31482, n31483, n31484,
    n31485, n31486, n31487, n31488, n31489, n31490,
    n31491, n31492, n31493, n31494, n31495, n31496,
    n31497, n31498, n31499, n31500, n31501, n31502,
    n31503, n31504, n31505, n31506, n31507, n31508,
    n31509, n31510, n31511, n31512, n31513, n31514,
    n31515, n31516, n31517, n31518, n31519, n31520,
    n31521, n31522, n31523, n31524, n31525, n31526,
    n31527, n31528, n31529, n31530, n31531, n31532,
    n31533, n31534, n31535, n31536, n31537, n31538,
    n31539, n31540, n31541, n31542, n31543, n31544,
    n31545, n31546, n31547, n31548, n31549, n31550,
    n31551, n31552, n31553, n31554, n31555, n31556,
    n31557, n31558, n31559, n31560, n31561, n31562,
    n31563, n31564, n31565, n31566, n31567, n31568,
    n31569, n31570, n31571, n31572, n31573, n31574,
    n31575, n31576, n31577, n31578, n31579, n31580,
    n31581, n31582, n31583, n31584, n31585, n31586,
    n31587, n31588, n31589, n31590, n31591, n31592,
    n31593, n31594, n31595, n31596, n31597, n31598,
    n31599, n31600, n31601, n31602, n31603, n31604,
    n31605, n31606, n31607, n31608, n31609, n31610,
    n31611, n31612, n31613, n31614, n31615, n31616,
    n31617, n31618, n31619, n31620, n31621, n31622,
    n31623, n31624, n31625, n31626, n31627, n31628,
    n31629, n31630, n31631, n31632, n31633, n31634,
    n31635, n31636, n31637, n31638, n31639, n31640,
    n31641, n31642, n31643, n31644, n31645, n31646,
    n31647, n31648, n31649, n31650, n31651, n31652,
    n31653, n31654, n31655, n31656, n31657, n31658,
    n31659, n31660, n31661, n31662, n31663, n31664,
    n31665, n31666, n31667, n31668, n31669, n31670,
    n31671, n31672, n31673, n31674, n31675, n31676,
    n31677, n31678, n31679, n31680, n31681, n31682,
    n31683, n31684, n31685, n31686, n31687, n31688,
    n31689, n31690, n31691, n31692, n31693, n31694,
    n31695, n31696, n31697, n31698, n31699, n31700,
    n31701, n31702, n31703, n31704, n31705, n31706,
    n31707, n31708, n31709, n31710, n31711, n31712,
    n31713, n31714, n31715, n31716, n31717, n31718,
    n31719, n31720, n31721, n31722, n31723, n31724,
    n31725, n31726, n31727, n31728, n31729, n31730,
    n31731, n31732, n31733, n31734, n31735, n31736,
    n31737, n31738, n31739, n31740, n31741, n31742,
    n31743, n31744, n31745, n31746, n31747, n31748,
    n31749, n31750, n31751, n31752, n31753, n31754,
    n31755, n31756, n31757, n31758, n31759, n31760,
    n31761, n31762, n31763, n31764, n31765, n31766,
    n31767, n31768, n31769, n31770, n31771, n31772,
    n31773, n31774, n31775, n31776, n31777, n31778,
    n31779, n31780, n31781, n31782, n31783, n31784,
    n31785, n31786, n31787, n31788, n31789, n31790,
    n31791, n31792, n31793, n31794, n31795, n31796,
    n31797, n31798, n31799, n31800, n31801, n31802,
    n31803, n31804, n31805, n31806, n31807, n31808,
    n31809, n31810, n31811, n31812, n31813, n31814,
    n31815, n31816, n31817, n31818, n31819, n31820,
    n31821, n31822, n31823, n31824, n31825, n31826,
    n31827, n31828, n31829, n31830, n31831, n31832,
    n31833, n31834, n31835, n31836, n31837, n31838,
    n31839, n31840, n31841, n31842, n31843, n31844,
    n31845, n31846, n31847, n31848, n31849, n31850,
    n31851, n31852, n31853, n31854, n31855, n31856,
    n31857, n31858, n31859, n31860, n31861, n31862,
    n31863, n31864, n31865, n31866, n31867, n31868,
    n31869, n31870, n31871, n31872, n31873, n31874,
    n31875, n31876, n31877, n31878, n31879, n31880,
    n31881, n31882, n31883, n31884, n31885, n31886,
    n31887, n31888, n31889, n31890, n31891, n31892,
    n31893, n31894, n31895, n31896, n31897, n31898,
    n31899, n31900, n31901, n31902, n31903, n31904,
    n31905, n31906, n31907, n31908, n31909, n31910,
    n31911, n31912, n31913, n31914, n31915, n31916,
    n31917, n31918, n31919, n31920, n31921, n31922,
    n31923, n31924, n31925, n31926, n31927, n31928,
    n31929, n31930, n31931, n31932, n31933, n31934,
    n31935, n31936, n31937, n31938, n31939, n31940,
    n31941, n31942, n31943, n31944, n31945, n31946,
    n31947, n31948, n31949, n31950, n31951, n31952,
    n31953, n31954, n31955, n31956, n31957, n31958,
    n31959, n31960, n31961, n31962, n31963, n31964,
    n31965, n31966, n31967, n31968, n31969, n31970,
    n31971, n31972, n31973, n31974, n31975, n31976,
    n31977, n31978, n31979, n31980, n31981, n31982,
    n31983, n31984, n31985, n31986, n31987, n31988,
    n31989, n31990, n31991, n31992, n31993, n31994,
    n31995, n31996, n31997, n31998, n31999, n32000,
    n32001, n32002, n32003, n32004, n32005, n32006,
    n32007, n32008, n32009, n32010, n32011, n32012,
    n32013, n32014, n32015, n32016, n32017, n32018,
    n32019, n32020, n32021, n32022, n32023, n32024,
    n32025, n32026, n32027, n32028, n32029, n32030,
    n32031, n32032, n32033, n32034, n32035, n32036,
    n32037, n32038, n32039, n32040, n32041, n32042,
    n32043, n32044, n32045, n32046, n32047, n32048,
    n32049, n32050, n32051, n32052, n32053, n32054,
    n32055, n32056, n32057, n32058, n32059, n32060,
    n32061, n32062, n32063, n32064, n32065, n32066,
    n32067, n32068, n32069, n32070, n32071, n32072,
    n32073, n32074, n32075, n32076, n32077, n32078,
    n32079, n32080, n32081, n32082, n32083, n32084,
    n32085, n32086, n32087, n32088, n32089, n32090,
    n32091, n32092, n32093, n32094, n32095, n32096,
    n32097, n32098, n32099, n32100, n32101, n32102,
    n32103, n32104, n32105, n32106, n32107, n32108,
    n32109, n32110, n32111, n32112, n32113, n32114,
    n32115, n32116, n32117, n32118, n32119, n32120,
    n32121, n32122, n32123, n32124, n32125, n32126,
    n32127, n32128, n32129, n32130, n32131, n32132,
    n32133, n32134, n32135, n32136, n32137, n32138,
    n32139, n32140, n32141, n32142, n32143, n32144,
    n32145, n32146, n32147, n32148, n32149, n32150,
    n32151, n32152, n32153, n32154, n32155, n32156,
    n32157, n32158, n32159, n32160, n32161, n32162,
    n32163, n32164, n32165, n32166, n32167, n32168,
    n32169, n32170, n32171, n32172, n32173, n32174,
    n32175, n32176, n32177, n32178, n32179, n32180,
    n32181, n32182, n32183, n32184, n32185, n32186,
    n32187, n32188, n32189, n32190, n32191, n32192,
    n32193, n32194, n32195, n32196, n32197, n32198,
    n32199, n32200, n32201, n32202, n32203, n32204,
    n32205, n32206, n32207, n32208, n32209, n32210,
    n32211, n32212, n32213, n32214, n32215, n32216,
    n32217, n32218, n32219, n32220, n32221, n32222,
    n32223, n32224, n32225, n32226, n32227, n32228,
    n32229, n32230, n32231, n32232, n32233, n32234,
    n32235, n32236, n32237, n32238, n32239, n32240,
    n32241, n32242, n32243, n32244, n32245, n32246,
    n32247, n32248, n32249, n32250, n32251, n32252,
    n32253, n32254, n32255, n32256, n32257, n32258,
    n32259, n32260, n32261, n32262, n32263, n32264,
    n32265, n32266, n32267, n32268, n32269, n32270,
    n32271, n32272, n32273, n32274, n32275, n32276,
    n32277, n32278, n32279, n32280, n32281, n32282,
    n32283, n32284, n32285, n32286, n32287, n32288,
    n32289, n32290, n32291, n32292, n32293, n32294,
    n32295, n32296, n32297, n32298, n32299, n32300,
    n32301, n32302, n32303, n32304, n32305, n32306,
    n32307, n32308, n32309, n32310, n32311, n32312,
    n32313, n32314, n32315, n32316, n32317, n32318,
    n32319, n32320, n32321, n32322, n32323, n32324,
    n32325, n32326, n32327, n32328, n32329, n32330,
    n32331, n32332, n32333, n32334, n32335, n32336,
    n32337, n32338, n32339, n32340, n32341, n32342,
    n32343, n32344, n32345, n32346, n32347, n32348,
    n32349, n32350, n32351, n32352, n32353, n32354,
    n32355, n32356, n32357, n32358, n32359, n32360,
    n32361, n32362, n32363, n32364, n32365, n32366,
    n32367, n32368, n32369, n32370, n32371, n32372,
    n32373, n32374, n32375, n32376, n32377, n32378,
    n32379, n32380, n32381, n32382, n32383, n32384,
    n32385, n32386, n32387, n32388, n32389, n32390,
    n32391, n32392, n32393, n32394, n32395, n32396,
    n32397, n32398, n32399, n32400, n32401, n32402,
    n32403, n32404, n32405, n32406, n32407, n32408,
    n32409, n32410, n32411, n32412, n32413, n32414,
    n32415, n32416, n32417, n32418, n32419, n32420,
    n32421, n32422, n32423, n32424, n32425, n32426,
    n32427, n32428, n32429, n32430, n32431, n32432,
    n32433, n32434, n32435, n32436, n32437, n32438,
    n32439, n32440, n32441, n32442, n32443, n32444,
    n32445, n32446, n32447, n32448, n32449, n32450,
    n32451, n32452, n32453, n32454, n32455, n32456,
    n32457, n32458, n32459, n32460, n32461, n32462,
    n32463, n32464, n32465, n32466, n32467, n32468,
    n32469, n32470, n32471, n32472, n32473, n32474,
    n32475, n32476, n32477, n32478, n32479, n32480,
    n32481, n32482, n32483, n32484, n32485, n32486,
    n32487, n32488, n32489, n32490, n32491, n32492,
    n32493, n32494, n32495, n32496, n32497, n32498,
    n32499, n32500, n32501, n32502, n32503, n32504,
    n32505, n32506, n32507, n32508, n32509, n32510,
    n32511, n32512, n32513, n32514, n32515, n32516,
    n32517, n32518, n32519, n32520, n32521, n32522,
    n32523, n32524, n32525, n32526, n32527, n32528,
    n32529, n32530, n32531, n32532, n32533, n32534,
    n32535, n32536, n32537, n32538, n32539, n32540,
    n32541, n32542, n32543, n32544, n32545, n32546,
    n32547, n32548, n32549, n32550, n32551, n32552,
    n32553, n32554, n32555, n32556, n32557, n32558,
    n32559, n32560, n32561, n32562, n32563, n32564,
    n32565, n32566, n32567, n32568, n32569, n32570,
    n32571, n32572, n32573, n32574, n32575, n32576,
    n32577, n32578, n32579, n32580, n32581, n32582,
    n32583, n32584, n32585, n32586, n32587, n32588,
    n32589, n32590, n32591, n32592, n32593, n32594,
    n32595, n32596, n32597, n32598, n32599, n32600,
    n32601, n32602, n32603, n32604, n32605, n32606,
    n32607, n32608, n32609, n32610, n32611, n32612,
    n32613, n32614, n32615, n32616, n32617, n32618,
    n32619, n32620, n32621, n32622, n32623, n32624,
    n32625, n32626, n32627, n32628, n32629, n32630,
    n32631, n32632, n32633, n32634, n32635, n32636,
    n32637, n32638, n32639, n32640, n32641, n32642,
    n32643, n32644, n32645, n32646, n32647, n32648,
    n32649, n32650, n32651, n32652, n32653, n32654,
    n32655, n32656, n32657, n32658, n32659, n32660,
    n32661, n32662, n32663, n32664, n32665, n32666,
    n32667, n32668, n32669, n32670, n32671, n32672,
    n32673, n32674, n32675, n32676, n32677, n32678,
    n32679, n32680, n32681, n32682, n32683, n32684,
    n32685, n32686, n32687, n32688, n32689, n32690,
    n32691, n32692, n32693, n32694, n32695, n32696,
    n32697, n32698, n32699, n32700, n32701, n32702,
    n32703, n32704, n32705, n32706, n32707, n32708,
    n32709, n32710, n32711, n32712, n32713, n32714,
    n32715, n32716, n32717, n32718, n32719, n32720,
    n32721, n32722, n32723, n32724, n32725, n32726,
    n32727, n32728, n32729, n32730, n32731, n32732,
    n32733, n32734, n32735, n32736, n32737, n32738,
    n32739, n32740, n32741, n32742, n32743, n32744,
    n32745, n32746, n32747, n32748, n32749, n32750,
    n32751, n32752, n32753, n32754, n32755, n32756,
    n32757, n32758, n32759, n32760, n32761, n32762,
    n32763, n32764, n32765, n32766, n32767, n32768,
    n32769, n32770, n32771, n32772, n32773, n32774,
    n32775, n32776, n32777, n32778, n32779, n32780,
    n32781, n32782, n32783, n32784, n32785, n32786,
    n32787, n32788, n32789, n32790, n32791, n32792,
    n32793, n32794, n32795, n32796, n32797, n32798,
    n32799, n32800, n32801, n32802, n32803, n32804,
    n32805, n32806, n32807, n32808, n32809, n32810,
    n32811, n32812, n32813, n32814, n32815, n32816,
    n32817, n32818, n32819, n32820, n32821, n32822,
    n32823, n32824, n32825, n32826, n32827, n32828,
    n32829, n32830, n32831, n32832, n32833, n32834,
    n32835, n32836, n32837, n32838, n32839, n32840,
    n32841, n32842, n32843, n32844, n32845, n32846,
    n32847, n32848, n32849, n32850, n32851, n32852,
    n32853, n32854, n32855, n32856, n32857, n32858,
    n32859, n32860, n32861, n32862, n32863, n32864,
    n32865, n32866, n32867, n32868, n32869, n32870,
    n32871, n32872, n32873, n32874, n32875, n32876,
    n32877, n32878, n32879, n32880, n32881, n32882,
    n32883, n32884, n32885, n32886, n32887, n32888,
    n32889, n32890, n32891, n32892, n32893, n32894,
    n32895, n32896, n32897, n32898, n32899, n32900,
    n32901, n32902, n32903, n32904, n32905, n32906,
    n32907, n32908, n32909, n32910, n32911, n32912,
    n32913, n32914, n32915, n32916, n32917, n32918,
    n32919, n32920, n32921, n32922, n32923, n32924,
    n32925, n32926, n32927, n32928, n32929, n32930,
    n32931, n32932, n32933, n32934, n32935, n32936,
    n32937, n32938, n32939, n32940, n32941, n32942,
    n32943, n32944, n32945, n32946, n32947, n32948,
    n32949, n32950, n32951, n32952, n32953, n32954,
    n32955, n32956, n32957, n32958, n32959, n32960,
    n32961, n32962, n32963, n32964, n32965, n32966,
    n32967, n32968, n32969, n32970, n32971, n32972,
    n32973, n32974, n32975, n32976, n32977, n32978,
    n32979, n32980, n32981, n32982, n32983, n32984,
    n32985, n32986, n32987, n32988, n32989, n32990,
    n32991, n32992, n32993, n32994, n32995, n32996,
    n32997, n32998, n32999, n33000, n33001, n33002,
    n33003, n33004, n33005, n33006, n33007, n33008,
    n33009, n33010, n33011, n33012, n33013, n33014,
    n33015, n33016, n33017, n33018, n33019, n33020,
    n33021, n33022, n33023, n33024, n33025, n33026,
    n33027, n33028, n33029, n33030, n33031, n33032,
    n33033, n33034, n33035, n33036, n33037, n33038,
    n33039, n33040, n33041, n33042, n33043, n33044,
    n33045, n33046, n33047, n33048, n33049, n33050,
    n33051, n33052, n33053, n33054, n33055, n33056,
    n33057, n33058, n33059, n33060, n33061, n33062,
    n33063, n33064, n33065, n33066, n33067, n33068,
    n33069, n33070, n33071, n33072, n33073, n33074,
    n33075, n33076, n33077, n33078, n33079, n33080,
    n33081, n33082, n33083, n33084, n33085, n33086,
    n33087, n33088, n33089, n33090, n33091, n33092,
    n33093, n33094, n33095, n33096, n33097, n33098,
    n33099, n33100, n33101, n33102, n33103, n33104,
    n33105, n33106, n33107, n33108, n33109, n33110,
    n33111, n33112, n33113, n33114, n33115, n33116,
    n33117, n33118, n33119, n33120, n33121, n33122,
    n33123, n33124, n33125, n33126, n33127, n33128,
    n33129, n33130, n33131, n33132, n33133, n33134,
    n33135, n33136, n33137, n33138, n33139, n33140,
    n33141, n33142, n33143, n33144, n33145, n33146,
    n33147, n33148, n33149, n33150, n33151, n33152,
    n33153, n33154, n33155, n33156, n33157, n33158,
    n33159, n33160, n33161, n33162, n33163, n33164,
    n33165, n33166, n33167, n33168, n33169, n33170,
    n33171, n33172, n33173, n33174, n33175, n33176,
    n33177, n33178, n33179, n33180, n33181, n33182,
    n33183, n33184, n33185, n33186, n33187, n33188,
    n33189, n33190, n33191, n33192, n33193, n33194,
    n33195, n33196, n33197, n33198, n33199, n33200,
    n33201, n33202, n33203, n33204, n33205, n33206,
    n33207, n33208, n33209, n33210, n33211, n33212,
    n33213, n33214, n33215, n33216, n33217, n33218,
    n33219, n33220, n33221, n33222, n33223, n33224,
    n33225, n33226, n33227, n33228, n33229, n33230,
    n33231, n33232, n33233, n33234, n33235, n33236,
    n33237, n33238, n33239, n33240, n33241, n33242,
    n33243, n33244, n33245, n33246, n33247, n33248,
    n33249, n33250, n33251, n33252, n33253, n33254,
    n33255, n33256, n33257, n33258, n33259, n33260,
    n33261, n33262, n33263, n33264, n33265, n33266,
    n33267, n33268, n33269, n33270, n33271, n33272,
    n33273, n33274, n33275, n33276, n33277, n33278,
    n33279, n33280, n33281, n33282, n33283, n33284,
    n33285, n33286, n33287, n33288, n33289, n33290,
    n33291, n33292, n33293, n33294, n33295, n33296,
    n33297, n33298, n33299, n33300, n33301, n33302,
    n33303, n33304, n33305, n33306, n33307, n33308,
    n33309, n33310, n33311, n33312, n33313, n33314,
    n33315, n33316, n33317, n33318, n33319, n33320,
    n33321, n33322, n33323, n33324, n33325, n33326,
    n33327, n33328, n33329, n33330, n33331, n33332,
    n33333, n33334, n33335, n33336, n33337, n33338,
    n33339, n33340, n33341, n33342, n33343, n33344,
    n33345, n33346, n33347, n33348, n33349, n33350,
    n33351, n33352, n33353, n33354, n33355, n33356,
    n33357, n33358, n33359, n33360, n33361, n33362,
    n33363, n33364, n33365, n33366, n33367, n33368,
    n33369, n33370, n33371, n33372, n33373, n33374,
    n33375, n33376, n33377, n33378, n33379, n33380,
    n33381, n33382, n33383, n33384, n33385, n33386,
    n33387, n33388, n33389, n33390, n33391, n33392,
    n33393, n33394, n33395, n33396, n33397, n33398,
    n33399, n33400, n33401, n33402, n33403, n33404,
    n33405, n33406, n33407, n33408, n33409, n33410,
    n33411, n33412, n33413, n33414, n33415, n33416,
    n33417, n33418, n33419, n33420, n33421, n33422,
    n33423, n33424, n33425, n33426, n33427, n33428,
    n33429, n33430, n33431, n33432, n33433, n33434,
    n33435, n33436, n33437, n33438, n33439, n33440,
    n33441, n33442, n33443, n33444, n33445, n33446,
    n33447, n33448, n33449, n33450, n33451, n33452,
    n33453, n33454, n33455, n33456, n33457, n33458,
    n33459, n33460, n33461, n33462, n33463, n33464,
    n33465, n33466, n33467, n33468, n33469, n33470,
    n33471, n33472, n33473, n33474, n33475, n33476,
    n33477, n33478, n33479, n33480, n33481, n33482,
    n33483, n33484, n33485, n33486, n33487, n33488,
    n33489, n33490, n33491, n33492, n33493, n33494,
    n33495, n33496, n33497, n33498, n33499, n33500,
    n33501, n33502, n33503, n33504, n33505, n33506,
    n33507, n33508, n33509, n33510, n33511, n33512,
    n33513, n33514, n33515, n33516, n33517, n33518,
    n33519, n33520, n33521, n33522, n33523, n33524,
    n33525, n33526, n33527, n33528, n33529, n33530,
    n33531, n33532, n33533, n33534, n33535, n33536,
    n33537, n33538, n33539, n33540, n33541, n33542,
    n33543, n33544, n33545, n33546, n33547, n33548,
    n33549, n33550, n33551, n33552, n33553, n33554,
    n33555, n33556, n33557, n33558, n33559, n33560,
    n33561, n33562, n33563, n33564, n33565, n33566,
    n33567, n33568, n33569, n33570, n33571, n33572,
    n33573, n33574, n33575, n33576, n33577, n33578,
    n33579, n33580, n33581, n33582, n33583, n33584,
    n33585, n33586, n33587, n33588, n33589, n33590,
    n33591, n33592, n33593, n33594, n33595, n33596,
    n33597, n33598, n33599, n33600, n33601, n33602,
    n33603, n33604, n33605, n33606, n33607, n33608,
    n33609, n33610, n33611, n33612, n33613, n33614,
    n33615, n33616, n33617, n33618, n33619, n33620,
    n33621, n33622, n33623, n33624, n33625, n33626,
    n33627, n33628, n33629, n33630, n33631, n33632,
    n33633, n33634, n33635, n33636, n33637, n33638,
    n33639, n33640, n33641, n33642, n33643, n33644,
    n33645, n33646, n33647, n33648, n33649, n33650,
    n33651, n33652, n33653, n33654, n33655, n33656,
    n33657, n33658, n33659, n33660, n33661, n33662,
    n33663, n33664, n33665, n33666, n33667, n33668,
    n33669, n33670, n33671, n33672, n33673, n33674,
    n33675, n33676, n33677, n33678, n33679, n33680,
    n33681, n33682, n33683, n33684, n33685, n33686,
    n33687, n33688, n33689, n33690, n33691, n33692,
    n33693, n33694, n33695, n33696, n33697, n33698,
    n33699, n33700, n33701, n33702, n33703, n33704,
    n33705, n33706, n33707, n33708, n33709, n33710,
    n33711, n33712, n33713, n33714, n33715, n33716,
    n33717, n33718, n33719, n33720, n33721, n33722,
    n33723, n33724, n33725, n33726, n33727, n33728,
    n33729, n33730, n33731, n33732, n33733, n33734,
    n33735, n33736, n33737, n33738, n33739, n33740,
    n33741, n33742, n33743, n33744, n33745, n33746,
    n33747, n33748, n33749, n33750, n33751, n33752,
    n33753, n33754, n33755, n33756, n33757, n33758,
    n33759, n33760, n33761, n33762, n33763, n33764,
    n33765, n33766, n33767, n33768, n33769, n33770,
    n33771, n33772, n33773, n33774, n33775, n33776,
    n33777, n33778, n33779, n33780, n33781, n33782,
    n33783, n33784, n33785, n33786, n33787, n33788,
    n33789, n33790, n33791, n33792, n33793, n33794,
    n33795, n33796, n33797, n33798, n33799, n33800,
    n33801, n33802, n33803, n33804, n33805, n33806,
    n33807, n33808, n33809, n33810, n33811, n33812,
    n33813, n33814, n33815, n33816, n33817, n33818,
    n33819, n33820, n33821, n33822, n33823, n33824,
    n33825, n33826, n33827, n33828, n33829, n33830,
    n33831, n33832, n33833, n33834, n33835, n33836,
    n33837, n33838, n33839, n33840, n33841, n33842,
    n33843, n33844, n33845, n33846, n33847, n33848,
    n33849, n33850, n33851, n33852, n33853, n33854,
    n33855, n33856, n33857, n33858, n33859, n33860,
    n33861, n33862, n33863, n33864, n33865, n33866,
    n33867, n33868, n33869, n33870, n33871, n33872,
    n33873, n33874, n33875, n33876, n33877, n33878,
    n33879, n33880, n33881, n33882, n33883, n33884,
    n33885, n33886, n33887, n33888, n33889, n33890,
    n33891, n33892, n33893, n33894, n33895, n33896,
    n33897, n33898, n33899, n33900, n33901, n33902,
    n33903, n33904, n33905, n33906, n33907, n33908,
    n33909, n33910, n33911, n33912, n33913, n33914,
    n33915, n33916, n33917, n33918, n33919, n33920,
    n33921, n33922, n33923, n33924, n33925, n33926,
    n33927, n33928, n33929, n33930, n33931, n33932,
    n33933, n33934, n33935, n33936, n33937, n33938,
    n33939, n33940, n33941, n33942, n33943, n33944,
    n33945, n33946, n33947, n33948, n33949, n33950,
    n33951, n33952, n33953, n33954, n33955, n33956,
    n33957, n33958, n33959, n33960, n33961, n33962,
    n33963, n33964, n33965, n33966, n33967, n33968,
    n33969, n33970, n33971, n33972, n33973, n33974,
    n33975, n33976, n33977, n33978, n33979, n33980,
    n33981, n33982, n33983, n33984, n33985, n33986,
    n33987, n33988, n33989, n33990, n33991, n33992,
    n33993, n33994, n33995, n33996, n33997, n33998,
    n33999, n34000, n34001, n34002, n34003, n34004,
    n34005, n34006, n34007, n34008, n34009, n34010,
    n34011, n34012, n34013, n34014, n34015, n34016,
    n34017, n34018, n34019, n34020, n34021, n34022,
    n34023, n34024, n34025, n34026, n34027, n34028,
    n34029, n34030, n34031, n34032, n34033, n34034,
    n34035, n34036, n34037, n34038, n34039, n34040,
    n34041, n34042, n34043, n34044, n34045, n34046,
    n34047, n34048, n34049, n34050, n34051, n34052,
    n34053, n34054, n34055, n34056, n34057, n34058,
    n34059, n34060, n34061, n34062, n34063, n34064,
    n34065, n34066, n34067, n34068, n34069, n34070,
    n34071, n34072, n34073, n34074, n34075, n34076,
    n34077, n34078, n34079, n34080, n34081, n34082,
    n34083, n34084, n34085, n34086, n34087, n34088,
    n34089, n34090, n34091, n34092, n34093, n34094,
    n34095, n34096, n34097, n34098, n34099, n34100,
    n34101, n34102, n34103, n34104, n34105, n34106,
    n34107, n34108, n34109, n34110, n34111, n34112,
    n34113, n34114, n34115, n34116, n34117, n34118,
    n34119, n34120, n34121, n34122, n34123, n34124,
    n34125, n34126, n34127, n34128, n34129, n34130,
    n34131, n34132, n34133, n34134, n34135, n34136,
    n34137, n34138, n34139, n34140, n34141, n34142,
    n34143, n34144, n34145, n34146, n34147, n34148,
    n34149, n34150, n34151, n34152, n34153, n34154,
    n34155, n34156, n34157, n34158, n34159, n34160,
    n34161, n34162, n34163, n34164, n34165, n34166,
    n34167, n34168, n34169, n34170, n34171, n34172,
    n34173, n34174, n34175, n34176, n34177, n34178,
    n34179, n34180, n34181, n34182, n34183, n34184,
    n34185, n34186, n34187, n34188, n34189, n34190,
    n34191, n34192, n34193, n34194, n34195, n34196,
    n34197, n34198, n34199, n34200, n34201, n34202,
    n34203, n34204, n34205, n34206, n34207, n34208,
    n34209, n34210, n34211, n34212, n34213, n34214,
    n34215, n34216, n34217, n34218, n34219, n34220,
    n34221, n34222, n34223, n34224, n34225, n34226,
    n34227, n34228, n34229, n34230, n34231, n34232,
    n34233, n34234, n34235, n34236, n34237, n34238,
    n34239, n34240, n34241, n34242, n34243, n34244,
    n34245, n34246, n34247, n34248, n34249, n34250,
    n34251, n34252, n34253, n34254, n34255, n34256,
    n34257, n34258, n34259, n34260, n34261, n34262,
    n34263, n34264, n34265, n34266, n34267, n34268,
    n34269, n34270, n34271, n34272, n34273, n34274,
    n34275, n34276, n34277, n34278, n34279, n34280,
    n34281, n34282, n34283, n34284, n34285, n34286,
    n34287, n34288, n34289, n34290, n34291, n34292,
    n34293, n34294, n34295, n34296, n34297, n34298,
    n34299, n34300, n34301, n34302, n34303, n34304,
    n34305, n34306, n34307, n34308, n34309, n34310,
    n34311, n34312, n34313, n34314, n34315, n34316,
    n34317, n34318, n34319, n34320, n34321, n34322,
    n34323, n34324, n34325, n34326, n34327, n34328,
    n34329, n34330, n34331, n34332, n34333, n34334,
    n34335, n34336, n34337, n34338, n34339, n34340,
    n34341, n34342, n34343, n34344, n34345, n34346,
    n34347, n34348, n34349, n34350, n34351, n34352,
    n34353, n34354, n34355, n34356, n34357, n34358,
    n34359, n34360, n34361, n34362, n34363, n34364,
    n34365, n34366, n34367, n34368, n34369, n34370,
    n34371, n34372, n34373, n34374, n34375, n34376,
    n34377, n34378, n34379, n34380, n34381, n34382,
    n34383, n34384, n34385, n34386, n34387, n34388,
    n34389, n34390, n34391, n34392, n34393, n34394,
    n34395, n34396, n34397, n34398, n34399, n34400,
    n34401, n34402, n34403, n34404, n34405, n34406,
    n34407, n34408, n34409, n34410, n34411, n34412,
    n34413, n34414, n34415, n34416, n34417, n34418,
    n34419, n34420, n34421, n34422, n34423, n34424,
    n34425, n34426, n34427, n34428, n34429, n34430,
    n34431, n34432, n34433, n34434, n34435, n34436,
    n34437, n34438, n34439, n34440, n34441, n34442,
    n34443, n34444, n34445, n34446, n34447, n34448,
    n34449, n34450, n34451, n34452, n34453, n34454,
    n34455, n34456, n34457, n34458, n34459, n34460,
    n34461, n34462, n34463, n34464, n34465, n34466,
    n34467, n34468, n34469, n34470, n34471, n34472,
    n34473, n34474, n34475, n34476, n34477, n34478,
    n34479, n34480, n34481, n34482, n34483, n34484,
    n34485, n34486, n34487, n34488, n34489, n34490,
    n34491, n34492, n34493, n34494, n34495, n34496,
    n34497, n34498, n34499, n34500, n34501, n34502,
    n34503, n34504, n34505, n34506, n34507, n34508,
    n34509, n34510, n34511, n34512, n34513, n34514,
    n34515, n34516, n34517, n34518, n34519, n34520,
    n34521, n34522, n34523, n34524, n34525, n34526,
    n34527, n34528, n34529, n34530, n34531, n34532,
    n34533, n34534, n34535, n34536, n34537, n34538,
    n34539, n34540, n34541, n34542, n34543, n34544,
    n34545, n34546, n34547, n34548, n34549, n34550,
    n34551, n34552, n34553, n34554, n34555, n34556,
    n34557, n34558, n34559, n34560, n34561, n34562,
    n34563, n34564, n34565, n34566, n34567, n34568,
    n34569, n34570, n34571, n34572, n34573, n34574,
    n34575, n34576, n34577, n34578, n34579, n34580,
    n34581, n34582, n34583, n34584, n34585, n34586,
    n34587, n34588, n34589, n34590, n34591, n34592,
    n34593, n34594, n34595, n34596, n34597, n34598,
    n34599, n34600, n34601, n34602, n34603, n34604,
    n34605, n34606, n34607, n34608, n34609, n34610,
    n34611, n34612, n34613, n34614, n34615, n34616,
    n34617, n34618, n34619, n34620, n34621, n34622,
    n34623, n34624, n34625, n34626, n34627, n34628,
    n34629, n34630, n34631, n34632, n34633, n34634,
    n34635, n34636, n34637, n34638, n34639, n34640,
    n34641, n34642, n34643, n34644, n34645, n34646,
    n34647, n34648, n34649, n34650, n34651, n34652,
    n34653, n34654, n34655, n34656, n34657, n34658,
    n34659, n34660, n34661, n34662, n34663, n34664,
    n34665, n34666, n34667, n34668, n34669, n34670,
    n34671, n34672, n34673, n34674, n34675, n34676,
    n34677, n34678, n34679, n34680, n34681, n34682,
    n34683, n34684, n34685, n34686, n34687, n34688,
    n34689, n34690, n34691, n34692, n34693, n34694,
    n34695, n34696, n34697, n34698, n34699, n34700,
    n34701, n34702, n34703, n34704, n34705, n34706,
    n34707, n34708, n34709, n34710, n34711, n34712,
    n34713, n34714, n34715, n34716, n34717, n34718,
    n34719, n34720, n34721, n34722, n34723, n34724,
    n34725, n34726, n34727, n34728, n34729, n34730,
    n34731, n34732, n34733, n34734, n34735, n34736,
    n34737, n34738, n34739, n34740, n34741, n34742,
    n34743, n34744, n34745, n34746, n34747, n34748,
    n34749, n34750, n34751, n34752, n34753, n34754,
    n34755, n34756, n34757, n34758, n34759, n34760,
    n34761, n34762, n34763, n34764, n34765, n34766,
    n34767, n34768, n34769, n34770, n34771, n34772,
    n34773, n34774, n34775, n34776, n34777, n34778,
    n34779, n34780, n34781, n34782, n34783, n34784,
    n34785, n34786, n34787, n34788, n34789, n34790,
    n34791, n34792, n34793, n34794, n34795, n34796,
    n34797, n34798, n34799, n34800, n34801, n34802,
    n34803, n34804, n34805, n34806, n34807, n34808,
    n34809, n34810, n34811, n34812, n34813, n34814,
    n34815, n34816, n34817, n34818, n34819, n34820,
    n34821, n34822, n34823, n34824, n34825, n34826,
    n34827, n34828, n34829, n34830, n34831, n34832,
    n34833, n34834, n34835, n34836, n34837, n34838,
    n34839, n34840, n34841, n34842, n34843, n34844,
    n34845, n34846, n34847, n34848, n34849, n34850,
    n34851, n34852, n34853, n34854, n34855, n34856,
    n34857, n34858, n34859, n34860, n34861, n34862,
    n34863, n34864, n34865, n34866, n34867, n34868,
    n34869, n34870, n34871, n34872, n34873, n34874,
    n34875, n34876, n34877, n34878, n34879, n34880,
    n34881, n34882, n34883, n34884, n34885, n34886,
    n34887, n34888, n34889, n34890, n34891, n34892,
    n34893, n34894, n34895, n34896, n34897, n34898,
    n34899, n34900, n34901, n34902, n34903, n34904,
    n34905, n34906, n34907, n34908, n34909, n34910,
    n34911, n34912, n34913, n34914, n34915, n34916,
    n34917, n34918, n34919, n34920, n34921, n34922,
    n34923, n34924, n34925, n34926, n34927, n34928,
    n34929, n34930, n34931, n34932, n34933, n34934,
    n34935, n34936, n34937, n34938, n34939, n34940,
    n34941, n34942, n34943, n34944, n34945, n34946,
    n34947, n34948, n34949, n34950, n34951, n34952,
    n34953, n34954, n34955, n34956, n34957, n34958,
    n34959, n34960, n34961, n34962, n34963, n34964,
    n34965, n34966, n34967, n34968, n34969, n34970,
    n34971, n34972, n34973, n34974, n34975, n34976,
    n34977, n34978, n34979, n34980, n34981, n34982,
    n34983, n34984, n34985, n34986, n34987, n34988,
    n34989, n34990, n34991, n34992, n34993, n34994,
    n34995, n34996, n34997, n34998, n34999, n35000,
    n35001, n35002, n35003, n35004, n35005, n35006,
    n35007, n35008, n35009, n35010, n35011, n35012,
    n35013, n35014, n35015, n35016, n35017, n35018,
    n35019, n35020, n35021, n35022, n35023, n35024,
    n35025, n35026, n35027, n35028, n35029, n35030,
    n35031, n35032, n35033, n35034, n35035, n35036,
    n35037, n35038, n35039, n35040, n35041, n35042,
    n35043, n35044, n35045, n35046, n35047, n35048,
    n35049, n35050, n35051, n35052, n35053, n35054,
    n35055, n35056, n35057, n35058, n35059, n35060,
    n35061, n35062, n35063, n35064, n35065, n35066,
    n35067, n35068, n35069, n35070, n35071, n35072,
    n35073, n35074, n35075, n35076, n35077, n35078,
    n35079, n35080, n35081, n35082, n35083, n35084,
    n35085, n35086, n35087, n35088, n35089, n35090,
    n35091, n35092, n35093, n35094, n35095, n35096,
    n35097, n35098, n35099, n35100, n35101, n35102,
    n35103, n35104, n35105, n35106, n35107, n35108,
    n35109, n35110, n35111, n35112, n35113, n35114,
    n35115, n35116, n35117, n35118, n35119, n35120,
    n35121, n35122, n35123, n35124, n35125, n35126,
    n35127, n35128, n35129, n35130, n35131, n35132,
    n35133, n35134, n35135, n35136, n35137, n35138,
    n35139, n35140, n35141, n35142, n35143, n35144,
    n35145, n35146, n35147, n35148, n35149, n35150,
    n35151, n35152, n35153, n35154, n35155, n35156,
    n35157, n35158, n35159, n35160, n35161, n35162,
    n35163, n35164, n35165, n35166, n35167, n35168,
    n35169, n35170, n35171, n35172, n35173, n35174,
    n35175, n35176, n35177, n35178, n35179, n35180,
    n35181, n35182, n35183, n35184, n35185, n35186,
    n35187, n35188, n35189, n35190, n35191, n35192,
    n35193, n35194, n35195, n35196, n35197, n35198,
    n35199, n35200, n35201, n35202, n35203, n35204,
    n35205, n35206, n35207, n35208, n35209, n35210,
    n35211, n35212, n35213, n35214, n35215, n35216,
    n35217, n35218, n35219, n35220, n35221, n35222,
    n35223, n35224, n35225, n35226, n35227, n35228,
    n35229, n35230, n35231, n35232, n35233, n35234,
    n35235, n35236, n35237, n35238, n35239, n35240,
    n35241, n35242, n35243, n35244, n35245, n35246,
    n35247, n35248, n35249, n35250, n35251, n35252,
    n35253, n35254, n35255, n35256, n35257, n35258,
    n35259, n35260, n35261, n35262, n35263, n35264,
    n35265, n35266, n35267, n35268, n35269, n35270,
    n35271, n35272, n35273, n35274, n35275, n35276,
    n35277, n35278, n35279, n35280, n35281, n35282,
    n35283, n35284, n35285, n35286, n35287, n35288,
    n35289, n35290, n35291, n35292, n35293, n35294,
    n35295, n35296, n35297, n35298, n35299, n35300,
    n35301, n35302, n35303, n35304, n35305, n35306,
    n35307, n35308, n35309, n35310, n35311, n35312,
    n35313, n35314, n35315, n35316, n35317, n35318,
    n35319, n35320, n35321, n35322, n35323, n35324,
    n35325, n35326, n35327, n35328, n35329, n35330,
    n35331, n35332, n35333, n35334, n35335, n35336,
    n35337, n35338, n35339, n35340, n35341, n35342,
    n35343, n35344, n35345, n35346, n35347, n35348,
    n35349, n35350, n35351, n35352, n35353, n35354,
    n35355, n35356, n35357, n35358, n35359, n35360,
    n35361, n35362, n35363, n35364, n35365, n35366,
    n35367, n35368, n35369, n35370, n35371, n35372,
    n35373, n35374, n35375, n35376, n35377, n35378,
    n35379, n35380, n35381, n35382, n35383, n35384,
    n35385, n35386, n35387, n35388, n35389, n35390,
    n35391, n35392, n35393, n35394, n35395, n35396,
    n35397, n35398, n35399, n35400, n35401, n35402,
    n35403, n35404, n35405, n35406, n35407, n35408,
    n35409, n35410, n35411, n35412, n35413, n35414,
    n35415, n35416, n35417, n35418, n35419, n35420,
    n35421, n35422, n35423, n35424, n35425, n35426,
    n35427, n35428, n35429, n35430, n35431, n35432,
    n35433, n35434, n35435, n35436, n35437, n35438,
    n35439, n35440, n35441, n35442, n35443, n35444,
    n35445, n35446, n35447, n35448, n35449, n35450,
    n35451, n35452, n35453, n35454, n35455, n35456,
    n35457, n35458, n35459, n35460, n35461, n35462,
    n35463, n35464, n35465, n35466, n35467, n35468,
    n35469, n35470, n35471, n35472, n35473, n35474,
    n35475, n35476, n35477, n35478, n35479, n35480,
    n35481, n35482, n35483, n35484, n35485, n35486,
    n35487, n35488, n35489, n35490, n35491, n35492,
    n35493, n35494, n35495, n35496, n35497, n35498,
    n35499, n35500, n35501, n35502, n35503, n35504,
    n35505, n35506, n35507, n35508, n35509, n35510,
    n35511, n35512, n35513, n35514, n35515, n35516,
    n35517, n35518, n35519, n35520, n35521, n35522,
    n35523, n35524, n35525, n35526, n35527, n35528,
    n35529, n35530, n35531, n35532, n35533, n35534,
    n35535, n35536, n35537, n35538, n35539, n35540,
    n35541, n35542, n35543, n35544, n35545, n35546,
    n35547, n35548, n35549, n35550, n35551, n35552,
    n35553, n35554, n35555, n35556, n35557, n35558,
    n35559, n35560, n35561, n35562, n35563, n35564,
    n35565, n35566, n35567, n35568, n35569, n35570,
    n35571, n35572, n35573, n35574, n35575, n35576,
    n35577, n35578, n35579, n35580, n35581, n35582,
    n35583, n35584, n35585, n35586, n35587, n35588,
    n35589, n35590, n35591, n35592, n35593, n35594,
    n35595, n35596, n35597, n35598, n35599, n35600,
    n35601, n35602, n35603, n35604, n35605, n35606,
    n35607, n35608, n35609, n35610, n35611, n35612,
    n35613, n35614, n35615, n35616, n35617, n35618,
    n35619, n35620, n35621, n35622, n35623, n35624,
    n35625, n35626, n35627, n35628, n35629, n35630,
    n35631, n35632, n35633, n35634, n35635, n35636,
    n35637, n35638, n35639, n35640, n35641, n35642,
    n35643, n35644, n35645, n35646, n35647, n35648,
    n35649, n35650, n35651, n35652, n35653, n35654,
    n35655, n35656, n35657, n35658, n35659, n35660,
    n35661, n35662, n35663, n35664, n35665, n35666,
    n35667, n35668, n35669, n35670, n35671, n35672,
    n35673, n35674, n35675, n35676, n35677, n35678,
    n35679, n35680, n35681, n35682, n35683, n35684,
    n35685, n35686, n35687, n35688, n35689, n35690,
    n35691, n35692, n35693, n35694, n35695, n35696,
    n35697, n35698, n35699, n35700, n35701, n35702,
    n35703, n35704, n35705, n35706, n35707, n35708,
    n35709, n35710, n35711, n35712, n35713, n35714,
    n35715, n35716, n35717, n35718, n35719, n35720,
    n35721, n35722, n35723, n35724, n35725, n35726,
    n35727, n35728, n35729, n35730, n35731, n35732,
    n35733, n35734, n35735, n35736, n35737, n35738,
    n35739, n35740, n35741, n35742, n35743, n35744,
    n35745, n35746, n35747, n35748, n35749, n35750,
    n35751, n35752, n35753, n35754, n35755, n35756,
    n35757, n35758, n35759, n35760, n35761, n35762,
    n35763, n35764, n35765, n35766, n35767, n35768,
    n35769, n35770, n35771, n35772, n35773, n35774,
    n35775, n35776, n35777, n35778, n35779, n35780,
    n35781, n35782, n35783, n35784, n35785, n35786,
    n35787, n35788, n35789, n35790, n35791, n35792,
    n35793, n35794, n35795, n35796, n35797, n35798,
    n35799, n35800, n35801, n35802, n35803, n35804,
    n35805, n35806, n35807, n35808, n35809, n35810,
    n35811, n35812, n35813, n35814, n35815, n35816,
    n35817, n35818, n35819, n35820, n35821, n35822,
    n35823, n35824, n35825, n35826, n35827, n35828,
    n35829, n35830, n35831, n35832, n35833, n35834,
    n35835, n35836, n35837, n35838, n35839, n35840,
    n35841, n35842, n35843, n35844, n35845, n35846,
    n35847, n35848, n35849, n35850, n35851, n35852,
    n35853, n35854, n35855, n35856, n35857, n35858,
    n35859, n35860, n35861, n35862, n35863, n35864,
    n35865, n35866, n35867, n35868, n35869, n35870,
    n35871, n35872, n35873, n35874, n35875, n35876,
    n35877, n35878, n35879, n35880, n35881, n35882,
    n35883, n35884, n35885, n35886, n35887, n35888,
    n35889, n35890, n35891, n35892, n35893, n35894,
    n35895, n35896, n35897, n35898, n35899, n35900,
    n35901, n35902, n35903, n35904, n35905, n35906,
    n35907, n35908, n35909, n35910, n35911, n35912,
    n35913, n35914, n35915, n35916, n35917, n35918,
    n35919, n35920, n35921, n35922, n35923, n35924,
    n35925, n35926, n35927, n35928, n35929, n35930,
    n35931, n35932, n35933, n35934, n35935, n35936,
    n35937, n35938, n35939, n35940, n35941, n35942,
    n35943, n35944, n35945, n35946, n35947, n35948,
    n35949, n35950, n35951, n35952, n35953, n35954,
    n35955, n35956, n35957, n35958, n35959, n35960,
    n35961, n35962, n35963, n35964, n35965, n35966,
    n35967, n35968, n35969, n35970, n35971, n35972,
    n35973, n35974, n35975, n35976, n35977, n35978,
    n35979, n35980, n35981, n35982, n35983, n35984,
    n35985, n35986, n35987, n35988, n35989, n35990,
    n35991, n35992, n35993, n35994, n35995, n35996,
    n35997, n35998, n35999, n36000, n36001, n36002,
    n36003, n36004, n36005, n36006, n36007, n36008,
    n36009, n36010, n36011, n36012, n36013, n36014,
    n36015, n36016, n36017, n36018, n36019, n36020,
    n36021, n36022, n36023, n36024, n36025, n36026,
    n36027, n36028, n36029, n36030, n36031, n36032,
    n36033, n36034, n36035, n36036, n36037, n36038,
    n36039, n36040, n36041, n36042, n36043, n36044,
    n36045, n36046, n36047, n36048, n36049, n36050,
    n36051, n36052, n36053, n36054, n36055, n36056,
    n36057, n36058, n36059, n36060, n36061, n36062,
    n36063, n36064, n36065, n36066, n36067, n36068,
    n36069, n36070, n36071, n36072, n36073, n36074,
    n36075, n36076, n36077, n36078, n36079, n36080,
    n36081, n36082, n36083, n36084, n36085, n36086,
    n36087, n36088, n36089, n36090, n36091, n36092,
    n36093, n36094, n36095, n36096, n36097, n36098,
    n36099, n36100, n36101, n36102, n36103, n36104,
    n36105, n36106, n36107, n36108, n36109, n36110,
    n36111, n36112, n36113, n36114, n36115, n36116,
    n36117, n36118, n36119, n36120, n36121, n36122,
    n36123, n36124, n36125, n36126, n36127, n36128,
    n36129, n36130, n36131, n36132, n36133, n36134,
    n36135, n36136, n36137, n36138, n36139, n36140,
    n36141, n36142, n36143, n36144, n36145, n36146,
    n36147, n36148, n36149, n36150, n36151, n36152,
    n36153, n36154, n36155, n36156, n36157, n36158,
    n36159, n36160, n36161, n36162, n36163, n36164,
    n36165, n36166, n36167, n36168, n36169, n36170,
    n36171, n36172, n36173, n36174, n36175, n36176,
    n36177, n36178, n36179, n36180, n36181, n36182,
    n36183, n36184, n36185, n36186, n36187, n36188,
    n36189, n36190, n36191, n36192, n36193, n36194,
    n36195, n36196, n36197, n36198, n36199, n36200,
    n36201, n36202, n36203, n36204, n36205, n36206,
    n36207, n36208, n36209, n36210, n36211, n36212,
    n36213, n36214, n36215, n36216, n36217, n36218,
    n36219, n36220, n36221, n36222, n36223, n36224,
    n36225, n36226, n36227, n36228, n36229, n36230,
    n36231, n36232, n36233, n36234, n36235, n36236,
    n36237, n36238, n36239, n36240, n36241, n36242,
    n36243, n36244, n36245, n36246, n36247, n36248,
    n36249, n36250, n36251, n36252, n36253, n36254,
    n36255, n36256, n36257, n36258, n36259, n36260,
    n36261, n36262, n36263, n36264, n36265, n36266,
    n36267, n36268, n36269, n36270, n36271, n36272,
    n36273, n36274, n36275, n36276, n36277, n36278,
    n36279, n36280, n36281, n36282, n36283, n36284,
    n36285, n36286, n36287, n36288, n36289, n36290,
    n36291, n36292, n36293, n36294, n36295, n36296,
    n36297, n36298, n36299, n36300, n36301, n36302,
    n36303, n36304, n36305, n36306, n36307, n36308,
    n36309, n36310, n36311, n36312, n36313, n36314,
    n36315, n36316, n36317, n36318, n36319, n36320,
    n36321, n36322, n36323, n36324, n36325, n36326,
    n36327, n36328, n36329, n36330, n36331, n36332,
    n36333, n36334, n36335, n36336, n36337, n36338,
    n36339, n36340, n36341, n36342, n36343, n36344,
    n36345, n36346, n36347, n36348, n36349, n36350,
    n36351, n36352, n36353, n36354, n36355, n36356,
    n36357, n36358, n36359, n36360, n36361, n36362,
    n36363, n36364, n36365, n36366, n36367, n36368,
    n36369, n36370, n36371, n36372, n36373, n36374,
    n36375, n36376, n36377, n36378, n36379, n36380,
    n36381, n36382, n36383, n36384, n36385, n36386,
    n36387, n36388, n36389, n36390, n36391, n36392,
    n36393, n36394, n36395, n36396, n36397, n36398,
    n36399, n36400, n36401, n36402, n36403, n36404,
    n36405, n36406, n36407, n36408, n36409, n36410,
    n36411, n36412, n36413, n36414, n36415, n36416,
    n36417, n36418, n36419, n36420, n36421, n36422,
    n36423, n36424, n36425, n36426, n36427, n36428,
    n36429, n36430, n36431, n36432, n36433, n36434,
    n36435, n36436, n36437, n36438, n36439, n36440,
    n36441, n36442, n36443, n36444, n36445, n36446,
    n36447, n36448, n36449, n36450, n36451, n36452,
    n36453, n36454, n36455, n36456, n36457, n36458,
    n36459, n36460, n36461, n36462, n36463, n36464,
    n36465, n36466, n36467, n36468, n36469, n36470,
    n36471, n36472, n36473, n36474, n36475, n36476,
    n36477, n36478, n36479, n36480, n36481, n36482,
    n36483, n36484, n36485, n36486, n36487, n36488,
    n36489, n36490, n36491, n36492, n36493, n36494,
    n36495, n36496, n36497, n36498, n36499, n36500,
    n36501, n36502, n36503, n36504, n36505, n36506,
    n36507, n36508, n36509, n36510, n36511, n36512,
    n36513, n36514, n36515, n36516, n36517, n36518,
    n36519, n36520, n36521, n36522, n36523, n36524,
    n36525, n36526, n36527, n36528, n36529, n36530,
    n36531, n36532, n36533, n36534, n36535, n36536,
    n36537, n36538, n36539, n36540, n36541, n36542,
    n36543, n36544, n36545, n36546, n36547, n36548,
    n36549, n36550, n36551, n36552, n36553, n36554,
    n36555, n36556, n36557, n36558, n36559, n36560,
    n36561, n36562, n36563, n36564, n36565, n36566,
    n36567, n36568, n36569, n36570, n36571, n36572,
    n36573, n36574, n36575, n36576, n36577, n36578,
    n36579, n36580, n36581, n36582, n36583, n36584,
    n36585, n36586, n36587, n36588, n36589, n36590,
    n36591, n36592, n36593, n36594, n36595, n36596,
    n36597, n36598, n36599, n36600, n36601, n36602,
    n36603, n36604, n36605, n36606, n36607, n36608,
    n36609, n36610, n36611, n36612, n36613, n36614,
    n36615, n36616, n36617, n36618, n36619, n36620,
    n36621, n36622, n36623, n36624, n36625, n36626,
    n36627, n36628, n36629, n36630, n36631, n36632,
    n36633, n36634, n36635, n36636, n36637, n36638,
    n36639, n36640, n36641, n36642, n36643, n36644,
    n36645, n36646, n36647, n36648, n36649, n36650,
    n36651, n36652, n36653, n36654, n36655, n36656,
    n36657, n36658, n36659, n36660, n36661, n36662,
    n36663, n36664, n36665, n36666, n36667, n36668,
    n36669, n36670, n36671, n36672, n36673, n36674,
    n36675, n36676, n36677, n36678, n36679, n36680,
    n36681, n36682, n36683, n36684, n36685, n36686,
    n36687, n36688, n36689, n36690, n36691, n36692,
    n36693, n36694, n36695, n36696, n36697, n36698,
    n36699, n36700, n36701, n36702, n36703, n36704,
    n36705, n36706, n36707, n36708, n36709, n36710,
    n36711, n36712, n36713, n36714, n36715, n36716,
    n36717, n36718, n36719, n36720, n36721, n36722,
    n36723, n36724, n36725, n36726, n36727, n36728,
    n36729, n36730, n36731, n36732, n36733, n36734,
    n36735, n36736, n36737, n36738, n36739, n36740,
    n36741, n36742, n36743, n36744, n36745, n36746,
    n36747, n36748, n36749, n36750, n36751, n36752,
    n36753, n36754, n36755, n36756, n36757, n36758,
    n36759, n36760, n36761, n36762, n36763, n36764,
    n36765, n36766, n36767, n36768, n36769, n36770,
    n36771, n36772, n36773, n36774, n36775, n36776,
    n36777, n36778, n36779, n36780, n36781, n36782,
    n36783, n36784, n36785, n36786, n36787, n36788,
    n36789, n36790, n36791, n36792, n36793, n36794,
    n36795, n36796, n36797, n36798, n36799, n36800,
    n36801, n36802, n36803, n36804, n36805, n36806,
    n36807, n36808, n36809, n36810, n36811, n36812,
    n36813, n36814, n36815, n36816, n36817, n36818,
    n36819, n36820, n36821, n36822, n36823, n36824,
    n36825, n36826, n36827, n36828, n36829, n36830,
    n36831, n36832, n36833, n36834, n36835, n36836,
    n36837, n36838, n36839, n36840, n36841, n36842,
    n36843, n36844, n36845, n36846, n36847, n36848,
    n36849, n36850, n36851, n36852, n36853, n36854,
    n36855, n36856, n36857, n36858, n36859, n36860,
    n36861, n36862, n36863, n36864, n36865, n36866,
    n36867, n36868, n36869, n36870, n36871, n36872,
    n36873, n36874, n36875, n36876, n36877, n36878,
    n36879, n36880, n36881, n36882, n36883, n36884,
    n36885, n36886, n36887, n36888, n36889, n36890,
    n36891, n36892, n36893, n36894, n36895, n36896,
    n36897, n36898, n36899, n36900, n36901, n36902,
    n36903, n36904, n36905, n36906, n36907, n36908,
    n36909, n36910, n36911, n36912, n36913, n36914,
    n36915, n36916, n36917, n36918, n36919, n36920,
    n36921, n36922, n36923, n36924, n36925, n36926,
    n36927, n36928, n36929, n36930, n36931, n36932,
    n36933, n36934, n36935, n36936, n36937, n36938,
    n36939, n36940, n36941, n36942, n36943, n36944,
    n36945, n36946, n36947, n36948, n36949, n36950,
    n36951, n36952, n36953, n36954, n36955, n36956,
    n36957, n36958, n36959, n36960, n36961, n36962,
    n36963, n36964, n36965, n36966, n36967, n36968,
    n36969, n36970, n36971, n36972, n36973, n36974,
    n36975, n36976, n36977, n36978, n36979, n36980,
    n36981, n36982, n36983, n36984, n36985, n36986,
    n36987, n36988, n36989, n36990, n36991, n36992,
    n36993, n36994, n36995, n36996, n36997, n36998,
    n36999, n37000, n37001, n37002, n37003, n37004,
    n37005, n37006, n37007, n37008, n37009, n37010,
    n37011, n37012, n37013, n37014, n37015, n37016,
    n37017, n37018, n37019, n37020, n37021, n37022,
    n37023, n37024, n37025, n37026, n37027, n37028,
    n37029, n37030, n37031, n37032, n37033, n37034,
    n37035, n37036, n37037, n37038, n37039, n37040,
    n37041, n37042, n37043, n37044, n37045, n37046,
    n37047, n37048, n37049, n37050, n37051, n37052,
    n37053, n37054, n37055, n37056, n37057, n37058,
    n37059, n37060, n37061, n37062, n37063, n37064,
    n37065, n37066, n37067, n37068, n37069, n37070,
    n37071, n37072, n37073, n37074, n37075, n37076,
    n37077, n37078, n37079, n37080, n37081, n37082,
    n37083, n37084, n37085, n37086, n37087, n37088,
    n37089, n37090, n37091, n37092, n37093, n37094,
    n37095, n37096, n37097, n37098, n37099, n37100,
    n37101, n37102, n37103, n37104, n37105, n37106,
    n37107, n37108, n37109, n37110, n37111, n37112,
    n37113, n37114, n37115, n37116, n37117, n37118,
    n37119, n37120, n37121, n37122, n37123, n37124,
    n37125, n37126, n37127, n37128, n37129, n37130,
    n37131, n37132, n37133, n37134, n37135, n37136,
    n37137, n37138, n37139, n37140, n37141, n37142,
    n37143, n37144, n37145, n37146, n37147, n37148,
    n37149, n37150, n37151, n37152, n37153, n37154,
    n37155, n37156, n37157, n37158, n37159, n37160,
    n37161, n37162, n37163, n37164, n37165, n37166,
    n37167, n37168, n37169, n37170, n37171, n37172,
    n37173, n37174, n37175, n37176, n37177, n37178,
    n37179, n37180, n37181, n37182, n37183, n37184,
    n37185, n37186, n37187, n37188, n37189, n37190,
    n37191, n37192, n37193, n37194, n37195, n37196,
    n37197, n37198, n37199, n37200, n37201, n37202,
    n37203, n37204, n37205, n37206, n37207, n37208,
    n37209, n37210, n37211, n37212, n37213, n37214,
    n37215, n37216, n37217, n37218, n37219, n37220,
    n37221, n37222, n37223, n37224, n37225, n37226,
    n37227, n37228, n37229, n37230, n37231, n37232,
    n37233, n37234, n37235, n37236, n37237, n37238,
    n37239, n37240, n37241, n37242, n37243, n37244,
    n37245, n37246, n37247, n37248, n37249, n37250,
    n37251, n37252, n37253, n37254, n37255, n37256,
    n37257, n37258, n37259, n37260, n37261, n37262,
    n37263, n37264, n37265, n37266, n37267, n37268,
    n37269, n37270, n37271, n37272, n37273, n37274,
    n37275, n37276, n37277, n37278, n37279, n37280,
    n37281, n37282, n37283, n37284, n37285, n37286,
    n37287, n37288, n37289, n37290, n37291, n37292,
    n37293, n37294, n37295, n37296, n37297, n37298,
    n37299, n37300, n37301, n37302, n37303, n37304,
    n37305, n37306, n37307, n37308, n37309, n37310,
    n37311, n37312, n37313, n37314, n37315, n37316,
    n37317, n37318, n37319, n37320, n37321, n37322,
    n37323, n37324, n37325, n37326, n37327, n37328,
    n37329, n37330, n37331, n37332, n37333, n37334,
    n37335, n37336, n37337, n37338, n37339, n37340,
    n37341, n37342, n37343, n37344, n37345, n37346,
    n37347, n37348, n37349, n37350, n37351, n37352,
    n37353, n37354, n37355, n37356, n37357, n37358,
    n37359, n37360, n37361, n37362, n37363, n37364,
    n37365, n37366, n37367, n37368, n37369, n37370,
    n37371, n37372, n37373, n37374, n37375, n37376,
    n37377, n37378, n37379, n37380, n37381, n37382,
    n37383, n37384, n37385, n37386, n37387, n37388,
    n37389, n37390, n37391, n37392, n37393, n37394,
    n37395, n37396, n37397, n37398, n37399, n37400,
    n37401, n37402, n37403, n37404, n37405, n37406,
    n37407, n37408, n37409, n37410, n37411, n37412,
    n37413, n37414, n37415, n37416, n37417, n37418,
    n37419, n37420, n37421, n37422, n37423, n37424,
    n37425, n37426, n37427, n37428, n37429, n37430,
    n37431, n37432, n37433, n37434, n37435, n37436,
    n37437, n37438, n37439, n37440, n37441, n37442,
    n37443, n37444, n37445, n37446, n37447, n37448,
    n37449, n37450, n37451, n37452, n37453, n37454,
    n37455, n37456, n37457, n37458, n37459, n37460,
    n37461, n37462, n37463, n37464, n37465, n37466,
    n37467, n37468, n37469, n37470, n37471, n37472,
    n37473, n37474, n37475, n37476, n37477, n37478,
    n37479, n37480, n37481, n37482, n37483, n37484,
    n37485, n37486, n37487, n37488, n37489, n37490,
    n37491, n37492, n37493, n37494, n37495, n37496,
    n37497, n37498, n37499, n37500, n37501, n37502,
    n37503, n37504, n37505, n37506, n37507, n37508,
    n37509, n37510, n37511, n37512, n37513, n37514,
    n37515, n37516, n37517, n37518, n37519, n37520,
    n37521, n37522, n37523, n37524, n37525, n37526,
    n37527, n37528, n37529, n37530, n37531, n37532,
    n37533, n37534, n37535, n37536, n37537, n37538,
    n37539, n37540, n37541, n37542, n37543, n37544,
    n37545, n37546, n37547, n37548, n37549, n37550,
    n37551, n37552, n37553, n37554, n37555, n37556,
    n37557, n37558, n37559, n37560, n37561, n37562,
    n37563, n37564, n37565, n37566, n37567, n37568,
    n37569, n37570, n37571, n37572, n37573, n37574,
    n37575, n37576, n37577, n37578, n37579, n37580,
    n37581, n37582, n37583, n37584, n37585, n37586,
    n37587, n37588, n37589, n37590, n37591, n37592,
    n37593, n37594, n37595, n37596, n37597, n37598,
    n37599, n37600, n37601, n37602, n37603, n37604,
    n37605, n37606, n37607, n37608, n37609, n37610,
    n37611, n37612, n37613, n37614, n37615, n37616,
    n37617, n37618, n37619, n37620, n37621, n37622,
    n37623, n37624, n37625, n37626, n37627, n37628,
    n37629, n37630, n37631, n37632, n37633, n37634,
    n37635, n37636, n37637, n37638, n37639, n37640,
    n37641, n37642, n37643, n37644, n37645, n37646,
    n37647, n37648, n37649, n37650, n37651, n37652,
    n37653, n37654, n37655, n37656, n37657, n37658,
    n37659, n37660, n37661, n37662, n37663, n37664,
    n37665, n37666, n37667, n37668, n37669, n37670,
    n37671, n37672, n37673, n37674, n37675, n37676,
    n37677, n37678, n37679, n37680, n37681, n37682,
    n37683, n37684, n37685, n37686, n37687, n37688,
    n37689, n37690, n37691, n37692, n37693, n37694,
    n37695, n37696, n37697, n37698, n37699, n37700,
    n37701, n37702, n37703, n37704, n37705, n37706,
    n37707, n37708, n37709, n37710, n37711, n37712,
    n37713, n37714, n37715, n37716, n37717, n37718,
    n37719, n37720, n37721, n37722, n37723, n37724,
    n37725, n37726, n37727, n37728, n37729, n37730,
    n37731, n37732, n37733, n37734, n37735, n37736,
    n37737, n37738, n37739, n37740, n37741, n37742,
    n37743, n37744, n37745, n37746, n37747, n37748,
    n37749, n37750, n37751, n37752, n37753, n37754,
    n37755, n37756, n37757, n37758, n37759, n37760,
    n37761, n37762, n37763, n37764, n37765, n37766,
    n37767, n37768, n37769, n37770, n37771, n37772,
    n37773, n37774, n37775, n37776, n37777, n37778,
    n37779, n37780, n37781, n37782, n37783, n37784,
    n37785, n37786, n37787, n37788, n37789, n37790,
    n37791, n37792, n37793, n37794, n37795, n37796,
    n37797, n37798, n37799, n37800, n37801, n37802,
    n37803, n37804, n37805, n37806, n37807, n37808,
    n37809, n37810, n37811, n37812, n37813, n37814,
    n37815, n37816, n37817, n37818, n37819, n37820,
    n37821, n37822, n37823, n37824, n37825, n37826,
    n37827, n37828, n37829, n37830, n37831, n37832,
    n37833, n37834, n37835, n37836, n37837, n37838,
    n37839, n37840, n37841, n37842, n37843, n37844,
    n37845, n37846, n37847, n37848, n37849, n37850,
    n37851, n37852, n37853, n37854, n37855, n37856,
    n37857, n37858, n37859, n37860, n37861, n37862,
    n37863, n37864, n37865, n37866, n37867, n37868,
    n37869, n37870, n37871, n37872, n37873, n37874,
    n37875, n37876, n37877, n37878, n37879, n37880,
    n37881, n37882, n37883, n37884, n37885, n37886,
    n37887, n37888, n37889, n37890, n37891, n37892,
    n37893, n37894, n37895, n37896, n37897, n37898,
    n37899, n37900, n37901, n37902, n37903, n37904,
    n37905, n37906, n37907, n37908, n37909, n37910,
    n37911, n37912, n37913, n37914, n37915, n37916,
    n37917, n37918, n37919, n37920, n37921, n37922,
    n37923, n37924, n37925, n37926, n37927, n37928,
    n37929, n37930, n37931, n37932, n37933, n37934,
    n37935, n37936, n37937, n37938, n37939, n37940,
    n37941, n37942, n37943, n37944, n37945, n37946,
    n37947, n37948, n37949, n37950, n37951, n37952,
    n37953, n37954, n37955, n37956, n37957, n37958,
    n37959, n37960, n37961, n37962, n37963, n37964,
    n37965, n37966, n37967, n37968, n37969, n37970,
    n37971, n37972, n37973, n37974, n37975, n37976,
    n37977, n37978, n37979, n37980, n37981, n37982,
    n37983, n37984, n37985, n37986, n37987, n37988,
    n37989, n37990, n37991, n37992, n37993, n37994,
    n37995, n37996, n37997, n37998, n37999, n38000,
    n38001, n38002, n38003, n38004, n38005, n38006,
    n38007, n38008, n38009, n38010, n38011, n38012,
    n38013, n38014, n38015, n38016, n38017, n38018,
    n38019, n38020, n38021, n38022, n38023, n38024,
    n38025, n38026, n38027, n38028, n38029, n38030,
    n38031, n38032, n38033, n38034, n38035, n38036,
    n38037, n38038, n38039, n38040, n38041, n38042,
    n38043, n38044, n38045, n38046, n38047, n38048,
    n38049, n38050, n38051, n38052, n38053, n38054,
    n38055, n38056, n38057, n38058, n38059, n38060,
    n38061, n38062, n38063, n38064, n38065, n38066,
    n38067, n38068, n38069, n38070, n38071, n38072,
    n38073, n38074, n38075, n38076, n38077, n38078,
    n38079, n38080, n38081, n38082, n38083, n38084,
    n38085, n38086, n38087, n38088, n38089, n38090,
    n38091, n38092, n38093, n38094, n38095, n38096,
    n38097, n38098, n38099, n38100, n38101, n38102,
    n38103, n38104, n38105, n38106, n38107, n38108,
    n38109, n38110, n38111, n38112, n38113, n38114,
    n38115, n38116, n38117, n38118, n38119, n38120,
    n38121, n38122, n38123, n38124, n38125, n38126,
    n38127, n38128, n38129, n38130, n38131, n38132,
    n38133, n38134, n38135, n38136, n38137, n38138,
    n38139, n38140, n38141, n38142, n38143, n38144,
    n38145, n38146, n38147, n38148, n38149, n38150,
    n38151, n38152, n38153, n38154, n38155, n38156,
    n38157, n38158, n38159, n38160, n38161, n38162,
    n38163, n38164, n38165, n38166, n38167, n38168,
    n38169, n38170, n38171, n38172, n38173, n38174,
    n38175, n38176, n38177, n38178, n38179, n38180,
    n38181, n38182, n38183, n38184, n38185, n38186,
    n38187, n38188, n38189, n38190, n38191, n38192,
    n38193, n38194, n38195, n38196, n38197, n38198,
    n38199, n38200, n38201, n38202, n38203, n38204,
    n38205, n38206, n38207, n38208, n38209, n38210,
    n38211, n38212, n38213, n38214, n38215, n38216,
    n38217, n38218, n38219, n38220, n38221, n38222,
    n38223, n38224, n38225, n38226, n38227, n38228,
    n38229, n38230, n38231, n38232, n38233, n38234,
    n38235, n38236, n38237, n38238, n38239, n38240,
    n38241, n38242, n38243, n38244, n38245, n38246,
    n38247, n38248, n38249, n38250, n38251, n38252,
    n38253, n38254, n38255, n38256, n38257, n38258,
    n38259, n38260, n38261, n38262, n38263, n38264,
    n38265, n38266, n38267, n38268, n38269, n38270,
    n38271, n38272, n38273, n38274, n38275, n38276,
    n38277, n38278, n38279, n38280, n38281, n38282,
    n38283, n38284, n38285, n38286, n38287, n38288,
    n38289, n38290, n38291, n38292, n38293, n38294,
    n38295, n38296, n38297, n38298, n38299, n38300,
    n38301, n38302, n38303, n38304, n38305, n38306,
    n38307, n38308, n38309, n38310, n38311, n38312,
    n38313, n38314, n38315, n38316, n38317, n38318,
    n38319, n38320, n38321, n38322, n38323, n38324,
    n38325, n38326, n38327, n38328, n38329, n38330,
    n38331, n38332, n38333, n38334, n38335, n38336,
    n38337, n38338, n38339, n38340, n38341, n38342,
    n38343, n38344, n38345, n38346, n38347, n38348,
    n38349, n38350, n38351, n38352, n38353, n38354,
    n38355, n38356, n38357, n38358, n38359, n38360,
    n38361, n38362, n38363, n38364, n38365, n38366,
    n38367, n38368, n38369, n38370, n38371, n38372,
    n38373, n38374, n38375, n38376, n38377, n38378,
    n38379, n38380, n38381, n38382, n38383, n38384,
    n38385, n38386, n38387, n38388, n38389, n38390,
    n38391, n38392, n38393, n38394, n38395, n38396,
    n38397, n38398, n38399, n38400, n38401, n38402,
    n38403, n38404, n38405, n38406, n38407, n38408,
    n38409, n38410, n38411, n38412, n38413, n38414,
    n38415, n38416, n38417, n38418, n38419, n38420,
    n38421, n38422, n38423, n38424, n38425, n38426,
    n38427, n38428, n38429, n38430, n38431, n38432,
    n38433, n38434, n38435, n38436, n38437, n38438,
    n38439, n38440, n38441, n38442, n38443, n38444,
    n38445, n38446, n38447, n38448, n38449, n38450,
    n38451, n38452, n38453, n38454, n38455, n38456,
    n38457, n38458, n38459, n38460, n38461, n38462,
    n38463, n38464, n38465, n38466, n38467, n38468,
    n38469, n38470, n38471, n38472, n38473, n38474,
    n38475, n38476, n38477, n38478, n38479, n38480,
    n38481, n38482, n38483, n38484, n38485, n38486,
    n38487, n38488, n38489, n38490, n38491, n38492,
    n38493, n38494, n38495, n38496, n38497, n38498,
    n38499, n38500, n38501, n38502, n38503, n38504,
    n38505, n38506, n38507, n38508, n38509, n38510,
    n38511, n38512, n38513, n38514, n38515, n38516,
    n38517, n38518, n38519, n38520, n38521, n38522,
    n38523, n38524, n38525, n38526, n38527, n38528,
    n38529, n38530, n38531, n38532, n38533, n38534,
    n38535, n38536, n38537, n38538, n38539, n38540,
    n38541, n38542, n38543, n38544, n38545, n38546,
    n38547, n38548, n38549, n38550, n38551, n38552,
    n38553, n38554, n38555, n38556, n38557, n38558,
    n38559, n38560, n38561, n38562, n38563, n38564,
    n38565, n38566, n38567, n38568, n38569, n38570,
    n38571, n38572, n38573, n38574, n38575, n38576,
    n38577, n38578, n38579, n38580, n38581, n38582,
    n38583, n38584, n38585, n38586, n38587, n38588,
    n38589, n38590, n38591, n38592, n38593, n38594,
    n38595, n38596, n38597, n38598, n38599, n38600,
    n38601, n38602, n38603, n38604, n38605, n38606,
    n38607, n38608, n38609, n38610, n38611, n38612,
    n38613, n38614, n38615, n38616, n38617, n38618,
    n38619, n38620, n38621, n38622, n38623, n38624,
    n38625, n38626, n38627, n38628, n38629, n38630,
    n38631, n38632, n38633, n38634, n38635, n38636,
    n38637, n38638, n38639, n38640, n38641, n38642,
    n38643, n38644, n38645, n38646, n38647, n38648,
    n38649, n38650, n38651, n38652, n38653, n38654,
    n38655, n38656, n38657, n38658, n38659, n38660,
    n38661, n38662, n38663, n38664, n38665, n38666,
    n38667, n38668, n38669, n38670, n38671, n38672,
    n38673, n38674, n38675, n38676, n38677, n38678,
    n38679, n38680, n38681, n38682, n38683, n38684,
    n38685, n38686, n38687, n38688, n38689, n38690,
    n38691, n38692, n38693, n38694, n38695, n38696,
    n38697, n38698, n38699, n38700, n38701, n38702,
    n38703, n38704, n38705, n38706, n38707, n38708,
    n38709, n38710, n38711, n38712, n38713, n38714,
    n38715, n38716, n38717, n38718, n38719, n38720,
    n38721, n38722, n38723, n38724, n38725, n38726,
    n38727, n38728, n38729, n38730, n38731, n38732,
    n38733, n38734, n38735, n38736, n38737, n38738,
    n38739, n38740, n38741, n38742, n38743, n38744,
    n38745, n38746, n38747, n38748, n38749, n38750,
    n38751, n38752, n38753, n38754, n38755, n38756,
    n38757, n38758, n38759, n38760, n38761, n38762,
    n38763, n38764, n38765, n38766, n38767, n38768,
    n38769, n38770, n38771, n38772, n38773, n38774,
    n38775, n38776, n38777, n38778, n38779, n38780,
    n38781, n38782, n38783, n38784, n38785, n38786,
    n38787, n38788, n38789, n38790, n38791, n38792,
    n38793, n38794, n38795, n38796, n38797, n38798,
    n38799, n38800, n38801, n38802, n38803, n38804,
    n38805, n38806, n38807, n38808, n38809, n38810,
    n38811, n38812, n38813, n38814, n38815, n38816,
    n38817, n38818, n38819, n38820, n38821, n38822,
    n38823, n38824, n38825, n38826, n38827, n38828,
    n38829, n38830, n38831, n38832, n38833, n38834,
    n38835, n38836, n38837, n38838, n38839, n38840,
    n38841, n38842, n38843, n38844, n38845, n38846,
    n38847, n38848, n38849, n38850, n38851, n38852,
    n38853, n38854, n38855, n38856, n38857, n38858,
    n38859, n38860, n38861, n38862, n38863, n38864,
    n38865, n38866, n38867, n38868, n38869, n38870,
    n38871, n38872, n38873, n38874, n38875, n38876,
    n38877, n38878, n38879, n38880, n38881, n38882,
    n38883, n38884, n38885, n38886, n38887, n38888,
    n38889, n38890, n38891, n38892, n38893, n38894,
    n38895, n38896, n38897, n38898, n38899, n38900,
    n38901, n38902, n38903, n38904, n38905, n38906,
    n38907, n38908, n38909, n38910, n38911, n38912,
    n38913, n38914, n38915, n38916, n38917, n38918,
    n38919, n38920, n38921, n38922, n38923, n38924,
    n38925, n38926, n38927, n38928, n38929, n38930,
    n38931, n38932, n38933, n38934, n38935, n38936,
    n38937, n38938, n38939, n38940, n38941, n38942,
    n38943, n38944, n38945, n38946, n38947, n38948,
    n38949, n38950, n38951, n38952, n38953, n38954,
    n38955, n38956, n38957, n38958, n38959, n38960,
    n38961, n38962, n38963, n38964, n38965, n38966,
    n38967, n38968, n38969, n38970, n38971, n38972,
    n38973, n38974, n38975, n38976, n38977, n38978,
    n38979, n38980, n38981, n38982, n38983, n38984,
    n38985, n38986, n38987, n38988, n38989, n38990,
    n38991, n38992, n38993, n38994, n38995, n38996,
    n38997, n38998, n38999, n39000, n39001, n39002,
    n39003, n39004, n39005, n39006, n39007, n39008,
    n39009, n39010, n39011, n39012, n39013, n39014,
    n39015, n39016, n39017, n39018, n39019, n39020,
    n39021, n39022, n39023, n39024, n39025, n39026,
    n39027, n39028, n39029, n39030, n39031, n39032,
    n39033, n39034, n39035, n39036, n39037, n39038,
    n39039, n39040, n39041, n39042, n39043, n39044,
    n39045, n39046, n39047, n39048, n39049, n39050,
    n39051, n39052, n39053, n39054, n39055, n39056,
    n39057, n39058, n39059, n39060, n39061, n39062,
    n39063, n39064, n39065, n39066, n39067, n39068,
    n39069, n39070, n39071, n39072, n39073, n39074,
    n39075, n39076, n39077, n39078, n39079, n39080,
    n39081, n39082, n39083, n39084, n39085, n39086,
    n39087, n39088, n39089, n39090, n39091, n39092,
    n39093, n39094, n39095, n39096, n39097, n39098,
    n39099, n39100, n39101, n39102, n39103, n39104,
    n39105, n39106, n39107, n39108, n39109, n39110,
    n39111, n39112, n39113, n39114, n39115, n39116,
    n39117, n39118, n39119, n39120, n39121, n39122,
    n39123, n39124, n39125, n39126, n39127, n39128,
    n39129, n39130, n39131, n39132, n39133, n39134,
    n39135, n39136, n39137, n39138, n39139, n39140,
    n39141, n39142, n39143, n39144, n39145, n39146,
    n39147, n39148, n39149, n39150, n39151, n39152,
    n39153, n39154, n39155, n39156, n39157, n39158,
    n39159, n39160, n39161, n39162, n39163, n39164,
    n39165, n39166, n39167, n39168, n39169, n39170,
    n39171, n39172, n39173, n39174, n39175, n39176,
    n39177, n39178, n39179, n39180, n39181, n39182,
    n39183, n39184, n39185, n39186, n39187, n39188,
    n39189, n39190, n39191, n39192, n39193, n39194,
    n39195, n39196, n39197, n39198, n39199, n39200,
    n39201, n39202, n39203, n39204, n39205, n39206,
    n39207, n39208, n39209, n39210, n39211, n39212,
    n39213, n39214, n39215, n39216, n39217, n39218,
    n39219, n39220, n39221, n39222, n39223, n39224,
    n39225, n39226, n39227, n39228, n39229, n39230,
    n39231, n39232, n39233, n39234, n39235, n39236,
    n39237, n39238, n39239, n39240, n39241, n39242,
    n39243, n39244, n39245, n39246, n39247, n39248,
    n39249, n39250, n39251, n39252, n39253, n39254,
    n39255, n39256, n39257, n39258, n39259, n39260,
    n39261, n39262, n39263, n39264, n39265, n39266,
    n39267, n39268, n39269, n39270, n39271, n39272,
    n39273, n39274, n39275, n39276, n39277, n39278,
    n39279, n39280, n39281, n39282, n39283, n39284,
    n39285, n39286, n39287, n39288, n39289, n39290,
    n39291, n39292, n39293, n39294, n39295, n39296,
    n39297, n39298, n39299, n39300, n39301, n39302,
    n39303, n39304, n39305, n39306, n39307, n39308,
    n39309, n39310, n39311, n39312, n39313, n39314,
    n39315, n39316, n39317, n39318, n39319, n39320,
    n39321, n39322, n39323, n39324, n39325, n39326,
    n39327, n39328, n39329, n39330, n39331, n39332,
    n39333, n39334, n39335, n39336, n39337, n39338,
    n39339, n39340, n39341, n39342, n39343, n39344,
    n39345, n39346, n39347, n39348, n39349, n39350,
    n39351, n39352, n39353, n39354, n39355, n39356,
    n39357, n39358, n39359, n39360, n39361, n39362,
    n39363, n39364, n39365, n39366, n39367, n39368,
    n39369, n39370, n39371, n39372, n39373, n39374,
    n39375, n39376, n39377, n39378, n39379, n39380,
    n39381, n39382, n39383, n39384, n39385, n39386,
    n39387, n39388, n39389, n39390, n39391, n39392,
    n39393, n39394, n39395, n39396, n39397, n39398,
    n39399, n39400, n39401, n39402, n39403, n39404,
    n39405, n39406, n39407, n39408, n39409, n39410,
    n39411, n39412, n39413, n39414, n39415, n39416,
    n39417, n39418, n39419, n39420, n39421, n39422,
    n39423, n39424, n39425, n39426, n39427, n39428,
    n39429, n39430, n39431, n39432, n39433, n39434,
    n39435, n39436, n39437, n39438, n39439, n39440,
    n39441, n39442, n39443, n39444, n39445, n39446,
    n39447, n39448, n39449, n39450, n39451, n39452,
    n39453, n39454, n39455, n39456, n39457, n39458,
    n39459, n39460, n39461, n39462, n39463, n39464,
    n39465, n39466, n39467, n39468, n39469, n39470,
    n39471, n39472, n39473, n39474, n39475, n39476,
    n39477, n39478, n39479, n39480, n39481, n39482,
    n39483, n39484, n39485, n39486, n39487, n39488,
    n39489, n39490, n39491, n39492, n39493, n39494,
    n39495, n39496, n39497, n39498, n39499, n39500,
    n39501, n39502, n39503, n39504, n39505, n39506,
    n39507, n39508, n39509, n39510, n39511, n39512,
    n39513, n39514, n39515, n39516, n39517, n39518,
    n39519, n39520, n39521, n39522, n39523, n39524,
    n39525, n39526, n39527, n39528, n39529, n39530,
    n39531, n39532, n39533, n39534, n39535, n39536,
    n39537, n39538, n39539, n39540, n39541, n39542,
    n39543, n39544, n39545, n39546, n39547, n39548,
    n39549, n39550, n39551, n39552, n39553, n39554,
    n39555, n39556, n39557, n39558, n39559, n39560,
    n39561, n39562, n39563, n39564, n39565, n39566,
    n39567, n39568, n39569, n39570, n39571, n39572,
    n39573, n39574, n39575, n39576, n39577, n39578,
    n39579, n39580, n39581, n39582, n39583, n39584,
    n39585, n39586, n39587, n39588, n39589, n39590,
    n39591, n39592, n39593, n39594, n39595, n39596,
    n39597, n39598, n39599, n39600, n39601, n39602,
    n39603, n39604, n39605, n39606, n39607, n39608,
    n39609, n39610, n39611, n39612, n39613, n39614,
    n39615, n39616, n39617, n39618, n39619, n39620,
    n39621, n39622, n39623, n39624, n39625, n39626,
    n39627, n39628, n39629, n39630, n39631, n39632,
    n39633, n39634, n39635, n39636, n39637, n39638,
    n39639, n39640, n39641, n39642, n39643, n39644,
    n39645, n39646, n39647, n39648, n39649, n39650,
    n39651, n39652, n39653, n39654, n39655, n39656,
    n39657, n39658, n39659, n39660, n39661, n39662,
    n39663, n39664, n39665, n39666, n39667, n39668,
    n39669, n39670, n39671, n39672, n39673, n39674,
    n39675, n39676, n39677, n39678, n39679, n39680,
    n39681, n39682, n39683, n39684, n39685, n39686,
    n39687, n39688, n39689, n39690, n39691, n39692,
    n39693, n39694, n39695, n39696, n39697, n39698,
    n39699, n39700, n39701, n39702, n39703, n39704,
    n39705, n39706, n39707, n39708, n39709, n39710,
    n39711, n39712, n39713, n39714, n39715, n39716,
    n39717, n39718, n39719, n39720, n39721, n39722,
    n39723, n39724, n39725, n39726, n39727, n39728,
    n39729, n39730, n39731, n39732, n39733, n39734,
    n39735, n39736, n39737, n39738, n39739, n39740,
    n39741, n39742, n39743, n39744, n39745, n39746,
    n39747, n39748, n39749, n39750, n39751, n39752,
    n39753, n39754, n39755, n39756, n39757, n39758,
    n39759, n39760, n39761, n39762, n39763, n39764,
    n39765, n39766, n39767, n39768, n39769, n39770,
    n39771, n39772, n39773, n39774, n39775, n39776,
    n39777, n39778, n39779, n39780, n39781, n39782,
    n39783, n39784, n39785, n39786, n39787, n39788,
    n39789, n39790, n39791, n39792, n39793, n39794,
    n39795, n39796, n39797, n39798, n39799, n39800,
    n39801, n39802, n39803, n39804, n39805, n39806,
    n39807, n39808, n39809, n39810, n39811, n39812,
    n39813, n39814, n39815, n39816, n39817, n39818,
    n39819, n39820, n39821, n39822, n39823, n39824,
    n39825, n39826, n39827, n39828, n39829, n39830,
    n39831, n39832, n39833, n39834, n39835, n39836,
    n39837, n39838, n39839, n39840, n39841, n39842,
    n39843, n39844, n39845, n39846, n39847, n39848,
    n39849, n39850, n39851, n39852, n39853, n39854,
    n39855, n39856, n39857, n39858, n39859, n39860,
    n39861, n39862, n39863, n39864, n39865, n39866,
    n39867, n39868, n39869, n39870, n39871, n39872,
    n39873, n39874, n39875, n39876, n39877, n39878,
    n39879, n39880, n39881, n39882, n39883, n39884,
    n39885, n39886, n39887, n39888, n39889, n39890,
    n39891, n39892, n39893, n39894, n39895, n39896,
    n39897, n39898, n39899, n39900, n39901, n39902,
    n39903, n39904, n39905, n39906, n39907, n39908,
    n39909, n39910, n39911, n39912, n39913, n39914,
    n39915, n39916, n39917, n39918, n39919, n39920,
    n39921, n39922, n39923, n39924, n39925, n39926,
    n39927, n39928, n39929, n39930, n39931, n39932,
    n39933, n39934, n39935, n39936, n39937, n39938,
    n39939, n39940, n39941, n39942, n39943, n39944,
    n39945, n39946, n39947, n39948, n39949, n39950,
    n39951, n39952, n39953, n39954, n39955, n39956,
    n39957, n39958, n39959, n39960, n39961, n39962,
    n39963, n39964, n39965, n39966, n39967, n39968,
    n39969, n39970, n39971, n39972, n39973, n39974,
    n39975, n39976, n39977, n39978, n39979, n39980,
    n39981, n39982, n39983, n39984, n39985, n39986,
    n39987, n39988, n39989, n39990, n39991, n39992,
    n39993, n39994, n39995, n39996, n39997, n39998,
    n39999, n40000, n40001, n40002, n40003, n40004,
    n40005, n40006, n40007, n40008, n40009, n40010,
    n40011, n40012, n40013, n40014, n40015, n40016,
    n40017, n40018, n40019, n40020, n40021, n40022,
    n40023, n40024, n40025, n40026, n40027, n40028,
    n40029, n40030, n40031, n40032, n40033, n40034,
    n40035, n40036, n40037, n40038, n40039, n40040,
    n40041, n40042, n40043, n40044, n40045, n40046,
    n40047, n40048, n40049, n40050, n40051, n40052,
    n40053, n40054, n40055, n40056, n40057, n40058,
    n40059, n40060, n40061, n40062, n40063, n40064,
    n40065, n40066, n40067, n40068, n40069, n40070,
    n40071, n40072, n40073, n40074, n40075, n40076,
    n40077, n40078, n40079, n40080, n40081, n40082,
    n40083, n40084, n40085, n40086, n40087, n40088,
    n40089, n40090, n40091, n40092, n40093, n40094,
    n40095, n40096, n40097, n40098, n40099, n40100,
    n40101, n40102, n40103, n40104, n40105, n40106,
    n40107, n40108, n40109, n40110, n40111, n40112,
    n40113, n40114, n40115, n40116, n40117, n40118,
    n40119, n40120, n40121, n40122, n40123, n40124,
    n40125, n40126, n40127, n40128, n40129, n40130,
    n40131, n40132, n40133, n40134, n40135, n40136,
    n40137, n40138, n40139, n40140, n40141, n40142,
    n40143, n40144, n40145, n40146, n40147, n40148,
    n40149, n40150, n40151, n40152, n40153, n40154,
    n40155, n40156, n40157, n40158, n40159, n40160,
    n40161, n40162, n40163, n40164, n40165, n40166,
    n40167, n40168, n40169, n40170, n40171, n40172,
    n40173, n40174, n40175, n40176, n40177, n40178,
    n40179, n40180, n40181, n40182, n40183, n40184,
    n40185, n40186, n40187, n40188, n40189, n40190,
    n40191, n40192, n40193, n40194, n40195, n40196,
    n40197, n40198, n40199, n40200, n40201, n40202,
    n40203, n40204, n40205, n40206, n40207, n40208,
    n40209, n40210, n40211, n40212, n40213, n40214,
    n40215, n40216, n40217, n40218, n40219, n40220,
    n40221, n40222, n40223, n40224, n40225, n40226,
    n40227, n40228, n40229, n40230, n40231, n40232,
    n40233, n40234, n40235, n40236, n40237, n40238,
    n40239, n40240, n40241, n40242, n40243, n40244,
    n40245, n40246, n40247, n40248, n40249, n40250,
    n40251, n40252, n40253, n40254, n40255, n40256,
    n40257, n40258, n40259, n40260, n40261, n40262,
    n40263, n40264, n40265, n40266, n40267, n40268,
    n40269, n40270, n40271, n40272, n40273, n40274,
    n40275, n40276, n40277, n40278, n40279, n40280,
    n40281, n40282, n40283, n40284, n40285, n40286,
    n40287, n40288, n40289, n40290, n40291, n40292,
    n40293, n40294, n40295, n40296, n40297, n40298,
    n40299, n40300, n40301, n40302, n40303, n40304,
    n40305, n40306, n40307, n40308, n40309, n40310,
    n40311, n40312, n40313, n40314, n40315, n40316,
    n40317, n40318, n40319, n40320, n40321, n40322,
    n40323, n40324, n40325, n40326, n40327, n40328,
    n40329, n40330, n40331, n40332, n40333, n40334,
    n40335, n40336, n40337, n40338, n40339, n40340,
    n40341, n40342, n40343, n40344, n40345, n40346,
    n40347, n40348, n40349, n40350, n40351, n40352,
    n40353, n40354, n40355, n40356, n40357, n40358,
    n40359, n40360, n40361, n40362, n40363, n40364,
    n40365, n40366, n40367, n40368, n40369, n40370,
    n40371, n40372, n40373, n40374, n40375, n40376,
    n40377, n40378, n40379, n40380, n40381, n40382,
    n40383, n40384, n40385, n40386, n40387, n40388,
    n40389, n40390, n40391, n40392, n40393, n40394,
    n40395, n40396, n40397, n40398, n40399, n40400,
    n40401, n40402, n40403, n40404, n40405, n40406,
    n40407, n40408, n40409, n40410, n40411, n40412,
    n40413, n40414, n40415, n40416, n40417, n40418,
    n40419, n40420, n40421, n40422, n40423, n40424,
    n40425, n40426, n40427, n40428, n40429, n40430,
    n40431, n40432, n40433, n40434, n40435, n40436,
    n40437, n40438, n40439, n40440, n40441, n40442,
    n40443, n40444, n40445, n40446, n40447, n40448,
    n40449, n40450, n40451, n40452, n40453, n40454,
    n40455, n40456, n40457, n40458, n40459, n40460,
    n40461, n40462, n40463, n40464, n40465, n40466,
    n40467, n40468, n40469, n40470, n40471, n40472,
    n40473, n40474, n40475, n40476, n40477, n40478,
    n40479, n40480, n40481, n40482, n40483, n40484,
    n40485, n40486, n40487, n40488, n40489, n40490,
    n40491, n40492, n40493, n40494, n40495, n40496,
    n40497, n40498, n40499, n40500, n40501, n40502,
    n40503, n40504, n40505, n40506, n40507, n40508,
    n40509, n40510, n40511, n40512, n40513, n40514,
    n40515, n40516, n40517, n40518, n40519, n40520,
    n40521, n40522, n40523, n40524, n40525, n40526,
    n40527, n40528, n40529, n40530, n40531, n40532,
    n40533, n40534, n40535, n40536, n40537, n40538,
    n40539, n40540, n40541, n40542, n40543, n40544,
    n40545, n40546, n40547, n40548, n40549, n40550,
    n40551, n40552, n40553, n40554, n40555, n40556,
    n40557, n40558, n40559, n40560, n40561, n40562,
    n40563, n40564, n40565, n40566, n40567, n40568,
    n40569, n40570, n40571, n40572, n40573, n40574,
    n40575, n40576, n40577, n40578, n40579, n40580,
    n40581, n40582, n40583, n40584, n40585, n40586,
    n40587, n40588, n40589, n40590, n40591, n40592,
    n40593, n40594, n40595, n40596, n40597, n40598,
    n40599, n40600, n40601, n40602, n40603, n40604,
    n40605, n40606, n40607, n40608, n40609, n40610,
    n40611, n40612, n40613, n40614, n40615, n40616,
    n40617, n40618, n40619, n40620, n40621, n40622,
    n40623, n40624, n40625, n40626, n40627, n40628,
    n40629, n40630, n40631, n40632, n40633, n40634,
    n40635, n40636, n40637, n40638, n40639, n40640,
    n40641, n40642, n40643, n40644, n40645, n40646,
    n40647, n40648, n40649, n40650, n40651, n40652,
    n40653, n40654, n40655, n40656, n40657, n40658,
    n40659, n40660, n40661, n40662, n40663, n40664,
    n40665, n40666, n40667, n40668, n40669, n40670,
    n40671, n40672, n40673, n40674, n40675, n40676,
    n40677, n40678, n40679, n40680, n40681, n40682,
    n40683, n40684, n40685, n40686, n40687, n40688,
    n40689, n40690, n40691, n40692, n40693, n40694,
    n40695, n40696, n40697, n40698, n40699, n40700,
    n40701, n40702, n40703, n40704, n40705, n40706,
    n40707, n40708, n40709, n40710, n40711, n40712,
    n40713, n40714, n40715, n40716, n40717, n40718,
    n40719, n40720, n40721, n40722, n40723, n40724,
    n40725, n40726, n40727, n40728, n40729, n40730,
    n40731, n40732, n40733, n40734, n40735, n40736,
    n40737, n40738, n40739, n40740, n40741, n40742,
    n40743, n40744, n40745, n40746, n40747, n40748,
    n40749, n40750, n40751, n40752, n40753, n40754,
    n40755, n40756, n40757, n40758, n40759, n40760,
    n40761, n40762, n40763, n40764, n40765, n40766,
    n40767, n40768, n40769, n40770, n40771, n40772,
    n40773, n40774, n40775, n40776, n40777, n40778,
    n40779, n40780, n40781, n40782, n40783, n40784,
    n40785, n40786, n40787, n40788, n40789, n40790,
    n40791, n40792, n40793, n40794, n40795, n40796,
    n40797, n40798, n40799, n40800, n40801, n40802,
    n40803, n40804, n40805, n40806, n40807, n40808,
    n40809, n40810, n40811, n40812, n40813, n40814,
    n40815, n40816, n40817, n40818, n40819, n40820,
    n40821, n40822, n40823, n40824, n40825, n40826,
    n40827, n40828, n40829, n40830, n40831, n40832,
    n40833, n40834, n40835, n40836, n40837, n40838,
    n40839, n40840, n40841, n40842, n40843, n40844,
    n40845, n40846, n40847, n40848, n40849, n40850,
    n40851, n40852, n40853, n40854, n40855, n40856,
    n40857, n40858, n40859, n40860, n40861, n40862,
    n40863, n40864, n40865, n40866, n40867, n40868,
    n40869, n40870, n40871, n40872, n40873, n40874,
    n40875, n40876, n40877, n40878, n40879, n40880,
    n40881, n40882, n40883, n40884, n40885, n40886,
    n40887, n40888, n40889, n40890, n40891, n40892,
    n40893, n40894, n40895, n40896, n40897, n40898,
    n40899, n40900, n40901, n40902, n40903, n40904,
    n40905, n40906, n40907, n40908, n40909, n40910,
    n40911, n40912, n40913, n40914, n40915, n40916,
    n40917, n40918, n40919, n40920, n40921, n40922,
    n40923, n40924, n40925, n40926, n40927, n40928,
    n40929, n40930, n40931, n40932, n40933, n40934,
    n40935, n40936, n40937, n40938, n40939, n40940,
    n40941, n40942, n40943, n40944, n40945, n40946,
    n40947, n40948, n40949, n40950, n40951, n40952,
    n40953, n40954, n40955, n40956, n40957, n40958,
    n40959, n40960, n40961, n40962, n40963, n40964,
    n40965, n40966, n40967, n40968, n40969, n40970,
    n40971, n40972, n40973, n40974, n40975, n40976,
    n40977, n40978, n40979, n40980, n40981, n40982,
    n40983, n40984, n40985, n40986, n40987, n40988,
    n40989, n40990, n40991, n40992, n40993, n40994,
    n40995, n40996, n40997, n40998, n40999, n41000,
    n41001, n41002, n41003, n41004, n41005, n41006,
    n41007, n41008, n41009, n41010, n41011, n41012,
    n41013, n41014, n41015, n41016, n41017, n41018,
    n41019, n41020, n41021, n41022, n41023, n41024,
    n41025, n41026, n41027, n41028, n41029, n41030,
    n41031, n41032, n41033, n41034, n41035, n41036,
    n41037, n41038, n41039, n41040, n41041, n41042,
    n41043, n41044, n41045, n41046, n41047, n41048,
    n41049, n41050, n41051, n41052, n41053, n41054,
    n41055, n41056, n41057, n41058, n41059, n41060,
    n41061, n41062, n41063, n41064, n41065, n41066,
    n41067, n41068, n41069, n41070, n41071, n41072,
    n41073, n41074, n41075, n41076, n41077, n41078,
    n41079, n41080, n41081, n41082, n41083, n41084,
    n41085, n41086, n41087, n41088, n41089, n41090,
    n41091, n41092, n41093, n41094, n41095, n41096,
    n41097, n41098, n41099, n41100, n41101, n41102,
    n41103, n41104, n41105, n41106, n41107, n41108,
    n41109, n41110, n41111, n41112, n41113, n41114,
    n41115, n41116, n41117, n41118, n41119, n41120,
    n41121, n41122, n41123, n41124, n41125, n41126,
    n41127, n41128, n41129, n41130, n41131, n41132,
    n41133, n41134, n41135, n41136, n41137, n41138,
    n41139, n41140, n41141, n41142, n41143, n41144,
    n41145, n41146, n41147, n41148, n41149, n41150,
    n41151, n41152, n41153, n41154, n41155, n41156,
    n41157, n41158, n41159, n41160, n41161, n41162,
    n41163, n41164, n41165, n41166, n41167, n41168,
    n41169, n41170, n41171, n41172, n41173, n41174,
    n41175, n41176, n41177, n41178, n41179, n41180,
    n41181, n41182, n41183, n41184, n41185, n41186,
    n41187, n41188, n41189, n41190, n41191, n41192,
    n41193, n41194, n41195, n41196, n41197, n41198,
    n41199, n41200, n41201, n41202, n41203, n41204,
    n41205, n41206, n41207, n41208, n41209, n41210,
    n41211, n41212, n41213, n41214, n41215, n41216,
    n41217, n41218, n41219, n41220, n41221, n41222,
    n41223, n41224, n41225, n41226, n41227, n41228,
    n41229, n41230, n41231, n41232, n41233, n41234,
    n41235, n41236, n41237, n41238, n41239, n41240,
    n41241, n41242, n41243, n41244, n41245, n41246,
    n41247, n41248, n41249, n41250, n41251, n41252,
    n41253, n41254, n41255, n41256, n41257, n41258,
    n41259, n41260, n41261, n41262, n41263, n41264,
    n41265, n41266, n41267, n41268, n41269, n41270,
    n41271, n41272, n41273, n41274, n41275, n41276,
    n41277, n41278, n41279, n41280, n41281, n41282,
    n41283, n41284, n41285, n41286, n41287, n41288,
    n41289, n41290, n41291, n41292, n41293, n41294,
    n41295, n41296, n41297, n41298, n41299, n41300,
    n41301, n41302, n41303, n41304, n41305, n41306,
    n41307, n41308, n41309, n41310, n41311, n41312,
    n41313, n41314, n41315, n41316, n41317, n41318,
    n41319, n41320, n41321, n41322, n41323, n41324,
    n41325, n41326, n41327, n41328, n41329, n41330,
    n41331, n41332, n41333, n41334, n41335, n41336,
    n41337, n41338, n41339, n41340, n41341, n41342,
    n41343, n41344, n41345, n41346, n41347, n41348,
    n41349, n41350, n41351, n41352, n41353, n41354,
    n41355, n41356, n41357, n41358, n41359, n41360,
    n41361, n41362, n41363, n41364, n41365, n41366,
    n41367, n41368, n41369, n41370, n41371, n41372,
    n41373, n41374, n41375, n41376, n41377, n41378,
    n41379, n41380, n41381, n41382, n41383, n41384,
    n41385, n41386, n41387, n41388, n41389, n41390,
    n41391, n41392, n41393, n41394, n41395, n41396,
    n41397, n41398, n41399, n41400, n41401, n41402,
    n41403, n41404, n41405, n41406, n41407, n41408,
    n41409, n41410, n41411, n41412, n41413, n41414,
    n41415, n41416, n41417, n41418, n41419, n41420,
    n41421, n41422, n41423, n41424, n41425, n41426,
    n41427, n41428, n41429, n41430, n41431, n41432,
    n41433, n41434, n41435, n41436, n41437, n41438,
    n41439, n41440, n41441, n41442, n41443, n41444,
    n41445, n41446, n41447, n41448, n41449, n41450,
    n41451, n41452, n41453, n41454, n41455, n41456,
    n41457, n41458, n41459, n41460, n41461, n41462,
    n41463, n41464, n41465, n41466, n41467, n41468,
    n41469, n41470, n41471, n41472, n41473, n41474,
    n41475, n41476, n41477, n41478, n41479, n41480,
    n41481, n41482, n41483, n41484, n41485, n41486,
    n41487, n41488, n41489, n41490, n41491, n41492,
    n41493, n41494, n41495, n41496, n41497, n41498,
    n41499, n41500, n41501, n41502, n41503, n41504,
    n41505, n41506, n41507, n41508, n41509, n41510,
    n41511, n41512, n41513, n41514, n41515, n41516,
    n41517, n41518, n41519, n41520, n41521, n41522,
    n41523, n41524, n41525, n41526, n41527, n41528,
    n41529, n41530, n41531, n41532, n41533, n41534,
    n41535, n41536, n41537, n41538, n41539, n41540,
    n41541, n41542, n41543, n41544, n41545, n41546,
    n41547, n41548, n41549, n41550, n41551, n41552,
    n41553, n41554, n41555, n41556, n41557, n41558,
    n41559, n41560, n41561, n41562, n41563, n41564,
    n41565, n41566, n41567, n41568, n41569, n41570,
    n41571, n41572, n41573, n41574, n41575, n41576,
    n41577, n41578, n41579, n41580, n41581, n41582,
    n41583, n41584, n41585, n41586, n41587, n41588,
    n41589, n41590, n41591, n41592, n41593, n41594,
    n41595, n41596, n41597, n41598, n41599, n41600,
    n41601, n41602, n41603, n41604, n41605, n41606,
    n41607, n41608, n41609, n41610, n41611, n41612,
    n41613, n41614, n41615, n41616, n41617, n41618,
    n41619, n41620, n41621, n41622, n41623, n41624,
    n41625, n41626, n41627, n41628, n41629, n41630,
    n41631, n41632, n41633, n41634, n41635, n41636,
    n41637, n41638, n41639, n41640, n41641, n41642,
    n41643, n41644, n41645, n41646, n41647, n41648,
    n41649, n41650, n41651, n41652, n41653, n41654,
    n41655, n41656, n41657, n41658, n41659, n41660,
    n41661, n41662, n41663, n41664, n41665, n41666,
    n41667, n41668, n41669, n41670, n41671, n41672,
    n41673, n41674, n41675, n41676, n41677, n41678,
    n41679, n41680, n41681, n41682, n41683, n41684,
    n41685, n41686, n41687, n41688, n41689, n41690,
    n41691, n41692, n41693, n41694, n41695, n41696,
    n41697, n41698, n41699, n41700, n41701, n41702,
    n41703, n41704, n41705, n41706, n41707, n41708,
    n41709, n41710, n41711, n41712, n41713, n41714,
    n41715, n41716, n41717, n41718, n41719, n41720,
    n41721, n41722, n41723, n41724, n41725, n41726,
    n41727, n41728, n41729, n41730, n41731, n41732,
    n41733, n41734, n41735, n41736, n41737, n41738,
    n41739, n41740, n41741, n41742, n41743, n41744,
    n41745, n41746, n41747, n41748, n41749, n41750,
    n41751, n41752, n41753, n41754, n41755, n41756,
    n41757, n41758, n41759, n41760, n41761, n41762,
    n41763, n41764, n41765, n41766, n41767, n41768,
    n41769, n41770, n41771, n41772, n41773, n41774,
    n41775, n41776, n41777, n41778, n41779, n41780,
    n41781, n41782, n41783, n41784, n41785, n41786,
    n41787, n41788, n41789, n41790, n41791, n41792,
    n41793, n41794, n41795, n41796, n41797, n41798,
    n41799, n41800, n41801, n41802, n41803, n41804,
    n41805, n41806, n41807, n41808, n41809, n41810,
    n41811, n41812, n41813, n41814, n41815, n41816,
    n41817, n41818, n41819, n41820, n41821, n41822,
    n41823, n41824, n41825, n41826, n41827, n41828,
    n41829, n41830, n41831, n41832, n41833, n41834,
    n41835, n41836, n41837, n41838, n41839, n41840,
    n41841, n41842, n41843, n41844, n41845, n41846,
    n41847, n41848, n41849, n41850, n41851, n41852,
    n41853, n41854, n41855, n41856, n41857, n41858,
    n41859, n41860, n41861, n41862, n41863, n41864,
    n41865, n41866, n41867, n41868, n41869, n41870,
    n41871, n41872, n41873, n41874, n41875, n41876,
    n41877, n41878, n41879, n41880, n41881, n41882,
    n41883, n41884, n41885, n41886, n41887, n41888,
    n41889, n41890, n41891, n41892, n41893, n41894,
    n41895, n41896, n41897, n41898, n41899, n41900,
    n41901, n41902, n41903, n41904, n41905, n41906,
    n41907, n41908, n41909, n41910, n41911, n41912,
    n41913, n41914, n41915, n41916, n41917, n41918,
    n41919, n41920, n41921, n41922, n41923, n41924,
    n41925, n41926, n41927, n41928, n41929, n41930,
    n41931, n41932, n41933, n41934, n41935, n41936,
    n41937, n41938, n41939, n41940, n41941, n41942,
    n41943, n41944, n41945, n41946, n41947, n41948,
    n41949, n41950, n41951, n41952, n41953, n41954,
    n41955, n41956, n41957, n41958, n41959, n41960,
    n41961, n41962, n41963, n41964, n41965, n41966,
    n41967, n41968, n41969, n41970, n41971, n41972,
    n41973, n41974, n41975, n41976, n41977, n41978,
    n41979, n41980, n41981, n41982, n41983, n41984,
    n41985, n41986, n41987, n41988, n41989, n41990,
    n41991, n41992, n41993, n41994, n41995, n41996,
    n41997, n41998, n41999, n42000, n42001, n42002,
    n42003, n42004, n42005, n42006, n42007, n42008,
    n42009, n42010, n42011, n42012, n42013, n42014,
    n42015, n42016, n42017, n42018, n42019, n42020,
    n42021, n42022, n42023, n42024, n42025, n42026,
    n42027, n42028, n42029, n42030, n42031, n42032,
    n42033, n42034, n42035, n42036, n42037, n42038,
    n42039, n42040, n42041, n42042, n42043, n42044,
    n42045, n42046, n42047, n42048, n42049, n42050,
    n42051, n42052, n42053, n42054, n42055, n42056,
    n42057, n42058, n42059, n42060, n42061, n42062,
    n42063, n42064, n42065, n42066, n42067, n42068,
    n42069, n42070, n42071, n42072, n42073, n42074,
    n42075, n42076, n42077, n42078, n42079, n42080,
    n42081, n42082, n42083, n42084, n42085, n42086,
    n42087, n42088, n42089, n42090, n42091, n42092,
    n42093, n42094, n42095, n42096, n42097, n42098,
    n42099, n42100, n42101, n42102, n42103, n42104,
    n42105, n42106, n42107, n42108, n42109, n42110,
    n42111, n42112, n42113, n42114, n42115, n42116,
    n42117, n42118, n42119, n42120, n42121, n42122,
    n42123, n42124, n42125, n42126, n42127, n42128,
    n42129, n42130, n42131, n42132, n42133, n42134,
    n42135, n42136, n42137, n42138, n42139, n42140,
    n42141, n42142, n42143, n42144, n42145, n42146,
    n42147, n42148, n42149, n42150, n42151, n42152,
    n42153, n42154, n42155, n42156, n42157, n42158,
    n42159, n42160, n42161, n42162, n42163, n42164,
    n42165, n42166, n42167, n42168, n42169, n42170,
    n42171, n42172, n42173, n42174, n42175, n42176,
    n42177, n42178, n42179, n42180, n42181, n42182,
    n42183, n42184, n42185, n42186, n42187, n42188,
    n42189, n42190, n42191, n42192, n42193, n42194,
    n42195, n42196, n42197, n42198, n42199, n42200,
    n42201, n42202, n42203, n42204, n42205, n42206,
    n42207, n42208, n42209, n42210, n42211, n42212,
    n42213, n42214, n42215, n42216, n42217, n42218,
    n42219, n42220, n42221, n42222, n42223, n42224,
    n42225, n42226, n42227, n42228, n42229, n42230,
    n42231, n42232, n42233, n42234, n42235, n42236,
    n42237, n42238, n42239, n42240, n42241, n42242,
    n42243, n42244, n42245, n42246, n42247, n42248,
    n42249, n42250, n42251, n42252, n42253, n42254,
    n42255, n42256, n42257, n42258, n42259, n42260,
    n42261, n42262, n42263, n42264, n42265, n42266,
    n42267, n42268, n42269, n42270, n42271, n42272,
    n42273, n42274, n42275, n42276, n42277, n42278,
    n42279, n42280, n42281, n42282, n42283, n42284,
    n42285, n42286, n42287, n42288, n42289, n42290,
    n42291, n42292, n42293, n42294, n42295, n42296,
    n42297, n42298, n42299, n42300, n42301, n42302,
    n42303, n42304, n42305, n42306, n42307, n42308,
    n42309, n42310, n42311, n42312, n42313, n42314,
    n42315, n42316, n42317, n42318, n42319, n42320,
    n42321, n42322, n42323, n42324, n42325, n42326,
    n42327, n42328, n42329, n42330, n42331, n42332,
    n42333, n42334, n42335, n42336, n42337, n42338,
    n42339, n42340, n42341, n42342, n42343, n42344,
    n42345, n42346, n42347, n42348, n42349, n42350,
    n42351, n42352, n42353, n42354, n42355, n42356,
    n42357, n42358, n42359, n42360, n42361, n42362,
    n42363, n42364, n42365, n42366, n42367, n42368,
    n42369, n42370, n42371, n42372, n42373, n42374,
    n42375, n42376, n42377, n42378, n42379, n42380,
    n42381, n42382, n42383, n42384, n42385, n42386,
    n42387, n42388, n42389, n42390, n42391, n42392,
    n42393, n42394, n42395, n42396, n42397, n42398,
    n42399, n42400, n42401, n42402, n42403, n42404,
    n42405, n42406, n42407, n42408, n42409, n42410,
    n42411, n42412, n42413, n42414, n42415, n42416,
    n42417, n42418, n42419, n42420, n42421, n42422,
    n42423, n42424, n42425, n42426, n42427, n42428,
    n42429, n42430, n42431, n42432, n42433, n42434,
    n42435, n42436, n42437, n42438, n42439, n42440,
    n42441, n42442, n42443, n42444, n42445, n42446,
    n42447, n42448, n42449, n42450, n42451, n42452,
    n42453, n42454, n42455, n42456, n42457, n42458,
    n42459, n42460, n42461, n42462, n42463, n42464,
    n42465, n42466, n42467, n42468, n42469, n42470,
    n42471, n42472, n42473, n42474, n42475, n42476,
    n42477, n42478, n42479, n42480, n42481, n42482,
    n42483, n42484, n42485, n42486, n42487, n42488,
    n42489, n42490, n42491, n42492, n42493, n42494,
    n42495, n42496, n42497, n42498, n42499, n42500,
    n42501, n42502, n42503, n42504, n42505, n42506,
    n42507, n42508, n42509, n42510, n42511, n42512,
    n42513, n42514, n42515, n42516, n42517, n42518,
    n42519, n42520, n42521, n42522, n42523, n42524,
    n42525, n42526, n42527, n42528, n42529, n42530,
    n42531, n42532, n42533, n42534, n42535, n42536,
    n42537, n42538, n42539, n42540, n42541, n42542,
    n42543, n42544, n42545, n42546, n42547, n42548,
    n42549, n42550, n42551, n42552, n42553, n42554,
    n42555, n42556, n42557, n42558, n42559, n42560,
    n42561, n42562, n42563, n42564, n42565, n42566,
    n42567, n42568, n42569, n42570, n42571, n42572,
    n42573, n42574, n42575, n42576, n42577, n42578,
    n42579, n42580, n42581, n42582, n42583, n42584,
    n42585, n42586, n42587, n42588, n42589, n42590,
    n42591, n42592, n42593, n42594, n42595, n42596,
    n42597, n42598, n42599, n42600, n42601, n42602,
    n42603, n42604, n42605, n42606, n42607, n42608,
    n42609, n42610, n42611, n42612, n42613, n42614,
    n42615, n42616, n42617, n42618, n42619, n42620,
    n42621, n42622, n42623, n42624, n42625, n42626,
    n42627, n42628, n42629, n42630, n42631, n42632,
    n42633, n42634, n42635, n42636, n42637, n42638,
    n42639, n42640, n42641, n42642, n42643, n42644,
    n42645, n42646, n42647, n42648, n42649, n42650,
    n42651, n42652, n42653, n42654, n42655, n42656,
    n42657, n42658, n42659, n42660, n42661, n42662,
    n42663, n42664, n42665, n42666, n42667, n42668,
    n42669, n42670, n42671, n42672, n42673, n42674,
    n42675, n42676, n42677, n42678, n42679, n42680,
    n42681, n42682, n42683, n42684, n42685, n42686,
    n42687, n42688, n42689, n42690, n42691, n42692,
    n42693, n42694, n42695, n42696, n42697, n42698,
    n42699, n42700, n42701, n42702, n42703, n42704,
    n42705, n42706, n42707, n42708, n42709, n42710,
    n42711, n42712, n42713, n42714, n42715, n42716,
    n42717, n42718, n42719, n42720, n42721, n42722,
    n42723, n42724, n42725, n42726, n42727, n42728,
    n42729, n42730, n42731, n42732, n42733, n42734,
    n42735, n42736, n42737, n42738, n42739, n42740,
    n42741, n42742, n42743, n42744, n42745, n42746,
    n42747, n42748, n42749, n42750, n42751, n42752,
    n42753, n42754, n42755, n42756, n42757, n42758,
    n42759, n42760, n42761, n42762, n42763, n42764,
    n42765, n42766, n42767, n42768, n42769, n42770,
    n42771, n42772, n42773, n42774, n42775, n42776,
    n42777, n42778, n42779, n42780, n42781, n42782,
    n42783, n42784, n42785, n42786, n42787, n42788,
    n42789, n42790, n42791, n42792, n42793, n42794,
    n42795, n42796, n42797, n42798, n42799, n42800,
    n42801, n42802, n42803, n42804, n42805, n42806,
    n42807, n42808, n42809, n42810, n42811, n42812,
    n42813, n42814, n42815, n42816, n42817, n42818,
    n42819, n42820, n42821, n42822, n42823, n42824,
    n42825, n42826, n42827, n42828, n42829, n42830,
    n42831, n42832, n42833, n42834, n42835, n42836,
    n42837, n42838, n42839, n42840, n42841, n42842,
    n42843, n42844, n42845, n42846, n42847, n42848,
    n42849, n42850, n42851, n42852, n42853, n42854,
    n42855, n42856, n42857, n42858, n42859, n42860,
    n42861, n42862, n42863, n42864, n42865, n42866,
    n42867, n42868, n42869, n42870, n42871, n42872,
    n42873, n42874, n42875, n42876, n42877, n42878,
    n42879, n42880, n42881, n42882, n42883, n42884,
    n42885, n42886, n42887, n42888, n42889, n42890,
    n42891, n42892, n42893, n42894, n42895, n42896,
    n42897, n42898, n42899, n42900, n42901, n42902,
    n42903, n42904, n42905, n42906, n42907, n42908,
    n42909, n42910, n42911, n42912, n42913, n42914,
    n42915, n42916, n42917, n42918, n42919, n42920,
    n42921, n42922, n42923, n42924, n42925, n42926,
    n42927, n42928, n42929, n42930, n42931, n42932,
    n42933, n42934, n42935, n42936, n42937, n42938,
    n42939, n42940, n42941, n42942, n42943, n42944,
    n42945, n42946, n42947, n42948, n42949, n42950,
    n42951, n42952, n42953, n42954, n42955, n42956,
    n42957, n42958, n42959, n42960, n42961, n42962,
    n42963, n42964, n42965, n42966, n42967, n42968,
    n42969, n42970, n42971, n42972, n42973, n42974,
    n42975, n42976, n42977, n42978, n42979, n42980,
    n42981, n42982, n42983, n42984, n42985, n42986,
    n42987, n42988, n42989, n42990, n42991, n42992,
    n42993, n42994, n42995, n42996, n42997, n42998,
    n42999, n43000, n43001, n43002, n43003, n43004,
    n43005, n43006, n43007, n43008, n43009, n43010,
    n43011, n43012, n43013, n43014, n43015, n43016,
    n43017, n43018, n43019, n43020, n43021, n43022,
    n43023, n43024, n43025, n43026, n43027, n43028,
    n43029, n43030, n43031, n43032, n43033, n43034,
    n43035, n43036, n43037, n43038, n43039, n43040,
    n43041, n43042, n43043, n43044, n43045, n43046,
    n43047, n43048, n43049, n43050, n43051, n43052,
    n43053, n43054, n43055, n43056, n43057, n43058,
    n43059, n43060, n43061, n43062, n43063, n43064,
    n43065, n43066, n43067, n43068, n43069, n43070,
    n43071, n43072, n43073, n43074, n43075, n43076,
    n43077, n43078, n43079, n43080, n43081, n43082,
    n43083, n43084, n43085, n43086, n43087, n43088,
    n43089, n43090, n43091, n43092, n43093, n43094,
    n43095, n43096, n43097, n43098, n43099, n43100,
    n43101, n43102, n43103, n43104, n43105, n43106,
    n43107, n43108, n43109, n43110, n43111, n43112,
    n43113, n43114, n43115, n43116, n43117, n43118,
    n43119, n43120, n43121, n43122, n43123, n43124,
    n43125, n43126, n43127, n43128, n43129, n43130,
    n43131, n43132, n43133, n43134, n43135, n43136,
    n43137, n43138, n43139, n43140, n43141, n43142,
    n43143, n43144, n43145, n43146, n43147, n43148,
    n43149, n43150, n43151, n43152, n43153, n43154,
    n43155, n43156, n43157, n43158, n43159, n43160,
    n43161, n43162, n43163, n43164, n43165, n43166,
    n43167, n43168, n43169, n43170, n43171, n43172,
    n43173, n43174, n43175, n43176, n43177, n43178,
    n43179, n43180, n43181, n43182, n43183, n43184,
    n43185, n43186, n43187, n43188, n43189, n43190,
    n43191, n43192, n43193, n43194, n43195, n43196,
    n43197, n43198, n43199, n43200, n43201, n43202,
    n43203, n43204, n43205, n43206, n43207, n43208,
    n43209, n43210, n43211, n43212, n43213, n43214,
    n43215, n43216, n43217, n43218, n43219, n43220,
    n43221, n43222, n43223, n43224, n43225, n43226,
    n43227, n43228, n43229, n43230, n43231, n43232,
    n43233, n43234, n43235, n43236, n43237, n43238,
    n43239, n43240, n43241, n43242, n43243, n43244,
    n43245, n43246, n43247, n43248, n43249, n43250,
    n43251, n43252, n43253, n43254, n43255, n43256,
    n43257, n43258, n43259, n43260, n43261, n43262,
    n43263, n43264, n43265, n43266, n43267, n43268,
    n43269, n43270, n43271, n43272, n43273, n43274,
    n43275, n43276, n43277, n43278, n43279, n43280,
    n43281, n43282, n43283, n43284, n43285, n43286,
    n43287, n43288, n43289, n43290, n43291, n43292,
    n43293, n43294, n43295, n43296, n43297, n43298,
    n43299, n43300, n43301, n43302, n43303, n43304,
    n43305, n43306, n43307, n43308, n43309, n43310,
    n43311, n43312, n43313, n43314, n43315, n43316,
    n43317, n43318, n43319, n43320, n43321, n43322,
    n43323, n43324, n43325, n43326, n43327, n43328,
    n43329, n43330, n43331, n43332, n43333, n43334,
    n43335, n43336, n43337, n43338, n43339, n43340,
    n43341, n43342, n43343, n43344, n43345, n43346,
    n43347, n43348, n43349, n43350, n43351, n43352,
    n43353, n43354, n43355, n43356, n43357, n43358,
    n43359, n43360, n43361, n43362, n43363, n43364,
    n43365, n43366, n43367, n43368, n43369, n43370,
    n43371, n43372, n43373, n43374, n43375, n43376,
    n43377, n43378, n43379, n43380, n43381, n43382,
    n43383, n43384, n43385, n43386, n43387, n43388,
    n43389, n43390, n43391, n43392, n43393, n43394,
    n43395, n43396, n43397, n43398, n43399, n43400,
    n43401, n43402, n43403, n43404, n43405, n43406,
    n43407, n43408, n43409, n43410, n43411, n43412,
    n43413, n43414, n43415, n43416, n43417, n43418,
    n43419, n43420, n43421, n43422, n43423, n43424,
    n43425, n43426, n43427, n43428, n43429, n43430,
    n43431, n43432, n43433, n43434, n43435, n43436,
    n43437, n43438, n43439, n43440, n43441, n43442,
    n43443, n43444, n43445, n43446, n43447, n43448,
    n43449, n43450, n43451, n43452, n43453, n43454,
    n43455, n43456, n43457, n43458, n43459, n43460,
    n43461, n43462, n43463, n43464, n43465, n43466,
    n43467, n43468, n43469, n43470, n43471, n43472,
    n43473, n43474, n43475, n43476, n43477, n43478,
    n43479, n43480, n43481, n43482, n43483, n43484,
    n43485, n43486, n43487, n43488, n43489, n43490,
    n43491, n43492, n43493, n43494, n43495, n43496,
    n43497, n43498, n43499, n43500, n43501, n43502,
    n43503, n43504, n43505, n43506, n43507, n43508,
    n43509, n43510, n43511, n43512, n43513, n43514,
    n43515, n43516, n43517, n43518, n43519, n43520,
    n43521, n43522, n43523, n43524, n43525, n43526,
    n43527, n43528, n43529, n43530, n43531, n43532,
    n43533, n43534, n43535, n43536, n43537, n43538,
    n43539, n43540, n43541, n43542, n43543, n43544,
    n43545, n43546, n43547, n43548, n43549, n43550,
    n43551, n43552, n43553, n43554, n43555, n43556,
    n43557, n43558, n43559, n43560, n43561, n43562,
    n43563, n43564, n43565, n43566, n43567, n43568,
    n43569, n43570, n43571, n43572, n43573, n43574,
    n43575, n43576, n43577, n43578, n43579, n43580,
    n43581, n43582, n43583, n43584, n43585, n43586,
    n43587, n43588, n43589, n43590, n43591, n43592,
    n43593, n43594, n43595, n43596, n43597, n43598,
    n43599, n43600, n43601, n43602, n43603, n43604,
    n43605, n43606, n43607, n43608, n43609, n43610,
    n43611, n43612, n43613, n43614, n43615, n43616,
    n43617, n43618, n43619, n43620, n43621, n43622,
    n43623, n43624, n43625, n43626, n43627, n43628,
    n43629, n43630, n43631, n43632, n43633, n43634,
    n43635, n43636, n43637, n43638, n43639, n43640,
    n43641, n43642, n43643, n43644, n43645, n43646,
    n43647, n43648, n43649, n43650, n43651, n43652,
    n43653, n43654, n43655, n43656, n43657, n43658,
    n43659, n43660, n43661, n43662, n43663, n43664,
    n43665, n43666, n43667, n43668, n43669, n43670,
    n43671, n43672, n43673, n43674, n43675, n43676,
    n43677, n43678, n43679, n43680, n43681, n43682,
    n43683, n43684, n43685, n43686, n43687, n43688,
    n43689, n43690, n43691, n43692, n43693, n43694,
    n43695, n43696, n43697, n43698, n43699, n43700,
    n43701, n43702, n43703, n43704, n43705, n43706,
    n43707, n43708, n43709, n43710, n43711, n43712,
    n43713, n43714, n43715, n43716, n43717, n43718,
    n43719, n43720, n43721, n43722, n43723, n43724,
    n43725, n43726, n43727, n43728, n43729, n43730,
    n43731, n43732, n43733, n43734, n43735, n43736,
    n43737, n43738, n43739, n43740, n43741, n43742,
    n43743, n43744, n43745, n43746, n43747, n43748,
    n43749, n43750, n43751, n43752, n43753, n43754,
    n43755, n43756, n43757, n43758, n43759, n43760,
    n43761, n43762, n43763, n43764, n43765, n43766,
    n43767, n43768, n43769, n43770, n43771, n43772,
    n43773, n43774, n43775, n43776, n43777, n43778,
    n43779, n43780, n43781, n43782, n43783, n43784,
    n43785, n43786, n43787, n43788, n43789, n43790,
    n43791, n43792, n43793, n43794, n43795, n43796,
    n43797, n43798, n43799, n43800, n43801, n43802,
    n43803, n43804, n43805, n43806, n43807, n43808,
    n43809, n43810, n43811, n43812, n43813, n43814,
    n43815, n43816, n43817, n43818, n43819, n43820,
    n43821, n43822, n43823, n43824, n43825, n43826,
    n43827, n43828, n43829, n43830, n43831, n43832,
    n43833, n43834, n43835, n43836, n43837, n43838,
    n43839, n43840, n43841, n43842, n43843, n43844,
    n43845, n43846, n43847, n43848, n43849, n43850,
    n43851, n43852, n43853, n43854, n43855, n43856,
    n43857, n43858, n43859, n43860, n43861, n43862,
    n43863, n43864, n43865, n43866, n43867, n43868,
    n43869, n43870, n43871, n43872, n43873, n43874,
    n43875, n43876, n43877, n43878, n43879, n43880,
    n43881, n43882, n43883, n43884, n43885, n43886,
    n43887, n43888, n43889, n43890, n43891, n43892,
    n43893, n43894, n43895, n43896, n43897, n43898,
    n43899, n43900, n43901, n43902, n43903, n43904,
    n43905, n43906, n43907, n43908, n43909, n43910,
    n43911, n43912, n43913, n43914, n43915, n43916,
    n43917, n43918, n43919, n43920, n43921, n43922,
    n43923, n43924, n43925, n43926, n43927, n43928,
    n43929, n43930, n43931, n43932, n43933, n43934,
    n43935, n43936, n43937, n43938, n43939, n43940,
    n43941, n43942, n43943, n43944, n43945, n43946,
    n43947, n43948, n43949, n43950, n43951, n43952,
    n43953, n43954, n43955, n43956, n43957, n43958,
    n43959, n43960, n43961, n43962, n43963, n43964,
    n43965, n43966, n43967, n43968, n43969, n43970,
    n43971, n43972, n43973, n43974, n43975, n43976,
    n43977, n43978, n43979, n43980, n43981, n43982,
    n43983, n43984, n43985, n43986, n43987, n43988,
    n43989, n43990, n43991, n43992, n43993, n43994,
    n43995, n43996, n43997, n43998, n43999, n44000,
    n44001, n44002, n44003, n44004, n44005, n44006,
    n44007, n44008, n44009, n44010, n44011, n44012,
    n44013, n44014, n44015, n44016, n44017, n44018,
    n44019, n44020, n44021, n44022, n44023, n44024,
    n44025, n44026, n44027, n44028, n44029, n44030,
    n44031, n44032, n44033, n44034, n44035, n44036,
    n44037, n44038, n44039, n44040, n44041, n44042,
    n44043, n44044, n44045, n44046, n44047, n44048,
    n44049, n44050, n44051, n44052, n44053, n44054,
    n44055, n44056, n44057, n44058, n44059, n44060,
    n44061, n44062, n44063, n44064, n44065, n44066,
    n44067, n44068, n44069, n44070, n44071, n44072,
    n44073, n44074, n44075, n44076, n44077, n44078,
    n44079, n44080, n44081, n44082, n44083, n44084,
    n44085, n44086, n44087, n44088, n44089, n44090,
    n44091, n44092, n44093, n44094, n44095, n44096,
    n44097, n44098, n44099, n44100, n44101, n44102,
    n44103, n44104, n44105, n44106, n44107, n44108,
    n44109, n44110, n44111, n44112, n44113, n44114,
    n44115, n44116, n44117, n44118, n44119, n44120,
    n44121, n44122, n44123, n44124, n44125, n44126,
    n44127, n44128, n44129, n44130, n44131, n44132,
    n44133, n44134, n44135, n44136, n44137, n44138,
    n44139, n44140, n44141, n44142, n44143, n44144,
    n44145, n44146, n44147, n44148, n44149, n44150,
    n44151, n44152, n44153, n44154, n44155, n44156,
    n44157, n44158, n44159, n44160, n44161, n44162,
    n44163, n44164, n44165, n44166, n44167, n44168,
    n44169, n44170, n44171, n44172, n44173, n44174,
    n44175, n44176, n44177, n44178, n44179, n44180,
    n44181, n44182, n44183, n44184, n44185, n44186,
    n44187, n44188, n44189, n44190, n44191, n44192,
    n44193, n44194, n44195, n44196, n44197, n44198,
    n44199, n44200, n44201, n44202, n44203, n44204,
    n44205, n44206, n44207, n44208, n44209, n44210,
    n44211, n44212, n44213, n44214, n44215, n44216,
    n44217, n44218, n44219, n44220, n44221, n44222,
    n44223, n44224, n44225, n44226, n44227, n44228,
    n44229, n44230, n44231, n44232, n44233, n44234,
    n44235, n44236, n44237, n44238, n44239, n44240,
    n44241, n44242, n44243, n44244, n44245, n44246,
    n44247, n44248, n44249, n44250, n44251, n44252,
    n44253, n44254, n44255, n44256, n44257, n44258,
    n44259, n44260, n44261, n44262, n44263, n44264,
    n44265, n44266, n44267, n44268, n44269, n44270,
    n44271, n44272, n44273, n44274, n44275, n44276,
    n44277, n44278, n44279, n44280, n44281, n44282,
    n44283, n44284, n44285, n44286, n44287, n44288,
    n44289, n44290, n44291, n44292, n44293, n44294,
    n44295, n44296, n44297, n44298, n44299, n44300,
    n44301, n44302, n44303, n44304, n44305, n44306,
    n44307, n44308, n44309, n44310, n44311, n44312,
    n44313, n44314, n44315, n44316, n44317, n44318,
    n44319, n44320, n44321, n44322, n44323, n44324,
    n44325, n44326, n44327, n44328, n44329, n44330,
    n44331, n44332, n44333, n44334, n44335, n44336,
    n44337, n44338, n44339, n44340, n44341, n44342,
    n44343, n44344, n44345, n44346, n44347, n44348,
    n44349, n44350, n44351, n44352, n44353, n44354,
    n44355, n44356, n44357, n44358, n44359, n44360,
    n44361, n44362, n44363, n44364, n44365, n44366,
    n44367, n44368, n44369, n44370, n44371, n44372,
    n44373, n44374, n44375, n44376, n44377, n44378,
    n44379, n44380, n44381, n44382, n44383, n44384,
    n44385, n44386, n44387, n44388, n44389, n44390,
    n44391, n44392, n44393, n44394, n44395, n44396,
    n44397, n44398, n44399, n44400, n44401, n44402,
    n44403, n44404, n44405, n44406, n44407, n44408,
    n44409, n44410, n44411, n44412, n44413, n44414,
    n44415, n44416, n44417, n44418, n44419, n44420,
    n44421, n44422, n44423, n44424, n44425, n44426,
    n44427, n44428, n44429, n44430, n44431, n44432,
    n44433, n44434, n44435, n44436, n44437, n44438,
    n44439, n44440, n44441, n44442, n44443, n44444,
    n44445, n44446, n44447, n44448, n44449, n44450,
    n44451, n44452, n44453, n44454, n44455, n44456,
    n44457, n44458, n44459, n44460, n44461, n44462,
    n44463, n44464, n44465, n44466, n44467, n44468,
    n44469, n44470, n44471, n44472, n44473, n44474,
    n44475, n44476, n44477, n44478, n44479, n44480,
    n44481, n44482, n44483, n44484, n44485, n44486,
    n44487, n44488, n44489, n44490, n44491, n44492,
    n44493, n44494, n44495, n44496, n44497, n44498,
    n44499, n44500, n44501, n44502, n44503, n44504,
    n44505, n44506, n44507, n44508, n44509, n44510,
    n44511, n44512, n44513, n44514, n44515, n44516,
    n44517, n44518, n44519, n44520, n44521, n44522,
    n44523, n44524, n44525, n44526, n44527, n44528,
    n44529, n44530, n44531, n44532, n44533, n44534,
    n44535, n44536, n44537, n44538, n44539, n44540,
    n44541, n44542, n44543, n44544, n44545, n44546,
    n44547, n44548, n44549, n44550, n44551, n44552,
    n44553, n44554, n44555, n44556, n44557, n44558,
    n44559, n44560, n44561, n44562, n44563, n44564,
    n44565, n44566, n44567, n44568, n44569, n44570,
    n44571, n44572, n44573, n44574, n44575, n44576,
    n44577, n44578, n44579, n44580, n44581, n44582,
    n44583, n44584, n44585, n44586, n44587, n44588,
    n44589, n44590, n44591, n44592, n44593, n44594,
    n44595, n44596, n44597, n44598, n44599, n44600,
    n44601, n44602, n44603, n44604, n44605, n44606,
    n44607, n44608, n44609, n44610, n44611, n44612,
    n44613, n44614, n44615, n44616, n44617, n44618,
    n44619, n44620, n44621, n44622, n44623, n44624,
    n44625, n44626, n44627, n44628, n44629, n44630,
    n44631, n44632, n44633, n44634, n44635, n44636,
    n44637, n44638, n44639, n44640, n44641, n44642,
    n44643, n44644, n44645, n44646, n44647, n44648,
    n44649, n44650, n44651, n44652, n44653, n44654,
    n44655, n44656, n44657, n44658, n44659, n44660,
    n44661, n44662, n44663, n44664, n44665, n44666,
    n44667, n44668, n44669, n44670, n44671, n44672,
    n44673, n44674, n44675, n44676, n44677, n44678,
    n44679, n44680, n44681, n44682, n44683, n44684,
    n44685, n44686, n44687, n44688, n44689, n44690,
    n44691, n44692, n44693, n44694, n44695, n44696,
    n44697, n44698, n44699, n44700, n44701, n44702,
    n44703, n44704, n44705, n44706, n44707, n44708,
    n44709, n44710, n44711, n44712, n44713, n44714,
    n44715, n44716, n44717, n44718, n44719, n44720,
    n44721, n44722, n44723, n44724, n44725, n44726,
    n44727, n44728, n44729, n44730, n44731, n44732,
    n44733, n44734, n44735, n44736, n44737, n44738,
    n44739, n44740, n44741, n44742, n44743, n44744,
    n44745, n44746, n44747, n44748, n44749, n44750,
    n44751, n44752, n44753, n44754, n44755, n44756,
    n44757, n44758, n44759, n44760, n44761, n44762,
    n44763, n44764, n44765, n44766, n44767, n44768,
    n44769, n44770, n44771, n44772, n44773, n44774,
    n44775, n44776, n44777, n44778, n44779, n44780,
    n44781, n44782, n44783, n44784, n44785, n44786,
    n44787, n44788, n44789, n44790, n44791, n44792,
    n44793, n44794, n44795, n44796, n44797, n44798,
    n44799, n44800, n44801, n44802, n44803, n44804,
    n44805, n44806, n44807, n44808, n44809, n44810,
    n44811, n44812, n44813, n44814, n44815, n44816,
    n44817, n44818, n44819, n44820, n44821, n44822,
    n44823, n44824, n44825, n44826, n44827, n44828,
    n44829, n44830, n44831, n44832, n44833, n44834,
    n44835, n44836, n44837, n44838, n44839, n44840,
    n44841, n44842, n44843, n44844, n44845, n44846,
    n44847, n44848, n44849, n44850, n44851, n44852,
    n44853, n44854, n44855, n44856, n44857, n44858,
    n44859, n44860, n44861, n44862, n44863, n44864,
    n44865, n44866, n44867, n44868, n44869, n44870,
    n44871, n44872, n44873, n44874, n44875, n44876,
    n44877, n44878, n44879, n44880, n44881, n44882,
    n44883, n44884, n44885, n44886, n44887, n44888,
    n44889, n44890, n44891, n44892, n44893, n44894,
    n44895, n44896, n44897, n44898, n44899, n44900,
    n44901, n44902, n44903, n44904, n44905, n44906,
    n44907, n44908, n44909, n44910, n44911, n44912,
    n44913, n44914, n44915, n44916, n44917, n44918,
    n44919, n44920, n44921, n44922, n44923, n44924,
    n44925, n44926, n44927, n44928, n44929, n44930,
    n44931, n44932, n44933, n44934, n44935, n44936,
    n44937, n44938, n44939, n44940, n44941, n44942,
    n44943, n44944, n44945, n44946, n44947, n44948,
    n44949, n44950, n44951, n44952, n44953, n44954,
    n44955, n44956, n44957, n44958, n44959, n44960,
    n44961, n44962, n44963, n44964, n44965, n44966,
    n44967, n44968, n44969, n44970, n44971, n44972,
    n44973, n44974, n44975, n44976, n44977, n44978,
    n44979, n44980, n44981, n44982, n44983, n44984,
    n44985, n44986, n44987, n44988, n44989, n44990,
    n44991, n44992, n44993, n44994, n44995, n44996,
    n44997, n44998, n44999, n45000, n45001, n45002,
    n45003, n45004, n45005, n45006, n45007, n45008,
    n45009, n45010, n45011, n45012, n45013, n45014,
    n45015, n45016, n45017, n45018, n45019, n45020,
    n45021, n45022, n45023, n45024, n45025, n45026,
    n45027, n45028, n45029, n45030, n45031, n45032,
    n45033, n45034, n45035, n45036, n45037, n45038,
    n45039, n45040, n45041, n45042, n45043, n45044,
    n45045, n45046, n45047, n45048, n45049, n45050,
    n45051, n45052, n45053, n45054, n45055, n45056,
    n45057, n45058, n45059, n45060, n45061, n45062,
    n45063, n45064, n45065, n45066, n45067, n45068,
    n45069, n45070, n45071, n45072, n45073, n45074,
    n45075, n45076, n45077, n45078, n45079, n45080,
    n45081, n45082, n45083, n45084, n45085, n45086,
    n45087, n45088, n45089, n45090, n45091, n45092,
    n45093, n45094, n45095, n45096, n45097, n45098,
    n45099, n45100, n45101, n45102, n45103, n45104,
    n45105, n45106, n45107, n45108, n45109, n45110,
    n45111, n45112, n45113, n45114, n45115, n45116,
    n45117, n45118, n45119, n45120, n45121, n45122,
    n45123, n45124, n45125, n45126, n45127, n45128,
    n45129, n45130, n45131, n45132, n45133, n45134,
    n45135, n45136, n45137, n45138, n45139, n45140,
    n45141, n45142, n45143, n45144, n45145, n45146,
    n45147, n45148, n45149, n45150, n45151, n45152,
    n45153, n45154, n45155, n45156, n45157, n45158,
    n45159, n45160, n45161, n45162, n45163, n45164,
    n45165, n45166, n45167, n45168, n45169, n45170,
    n45171, n45172, n45173, n45174, n45175, n45176,
    n45177, n45178, n45179, n45180, n45181, n45182,
    n45183, n45184, n45185, n45186, n45187, n45188,
    n45189, n45190, n45191, n45192, n45193, n45194,
    n45195, n45196, n45197, n45198, n45199, n45200,
    n45201, n45202, n45203, n45204, n45205, n45206,
    n45207, n45208, n45209, n45210, n45211, n45212,
    n45213, n45214, n45215, n45216, n45217, n45218,
    n45219, n45220, n45221, n45222, n45223, n45224,
    n45225, n45226, n45227, n45228, n45229, n45230,
    n45231, n45232, n45233, n45234, n45235, n45236,
    n45237, n45238, n45239, n45240, n45241, n45242,
    n45243, n45244, n45245, n45246, n45247, n45248,
    n45249, n45250, n45251, n45252, n45253, n45254,
    n45255, n45256, n45257, n45258, n45259, n45260,
    n45261, n45262, n45263, n45264, n45265, n45266,
    n45267, n45268, n45269, n45270, n45271, n45272,
    n45273, n45274, n45275, n45276, n45277, n45278,
    n45279, n45280, n45281, n45282, n45283, n45284,
    n45285, n45286, n45287, n45288, n45289, n45290,
    n45291, n45292, n45293, n45294, n45295, n45296,
    n45297, n45298, n45299, n45300, n45301, n45302,
    n45303, n45304, n45305, n45306, n45307, n45308,
    n45309, n45310, n45311, n45312, n45313, n45314,
    n45315, n45316, n45317, n45318, n45319, n45320,
    n45321, n45322, n45323, n45324, n45325, n45326,
    n45327, n45328, n45329, n45330, n45331, n45332,
    n45333, n45334, n45335, n45336, n45337, n45338,
    n45339, n45340, n45341, n45342, n45343, n45344,
    n45345, n45346, n45347, n45348, n45349, n45350,
    n45351, n45352, n45353, n45354, n45355, n45356,
    n45357, n45358, n45359, n45360, n45361, n45362,
    n45363, n45364, n45365, n45366, n45367, n45368,
    n45369, n45370, n45371, n45372, n45373, n45374,
    n45375, n45376, n45377, n45378, n45379, n45380,
    n45381, n45382, n45383, n45384, n45385, n45386,
    n45387, n45388, n45389, n45390, n45391, n45392,
    n45393, n45394, n45395, n45396, n45397, n45398,
    n45399, n45400, n45401, n45402, n45403, n45404,
    n45405, n45406, n45407, n45408, n45409, n45410,
    n45411, n45412, n45413, n45414, n45415, n45416,
    n45417, n45418, n45419, n45420, n45421, n45422,
    n45423, n45424, n45425, n45426, n45427, n45428,
    n45429, n45430, n45431, n45432, n45433, n45434,
    n45435, n45436, n45437, n45438, n45439, n45440,
    n45441, n45442, n45443, n45444, n45445, n45446,
    n45447, n45448, n45449, n45450, n45451, n45452,
    n45453, n45454, n45455, n45456, n45457, n45458,
    n45459, n45460, n45461, n45462, n45463, n45464,
    n45465, n45466, n45467, n45468, n45469, n45470,
    n45471, n45472, n45473, n45474, n45475, n45476,
    n45477, n45478, n45479, n45480, n45481, n45482,
    n45483, n45484, n45485, n45486, n45487, n45488,
    n45489, n45490, n45491, n45492, n45493, n45494,
    n45495, n45496, n45497, n45498, n45499, n45500,
    n45501, n45502, n45503, n45504, n45505, n45506,
    n45507, n45508, n45509, n45510, n45511, n45512,
    n45513, n45514, n45515, n45516, n45517, n45518,
    n45519, n45520, n45521, n45522, n45523, n45524,
    n45525, n45526, n45527, n45528, n45529, n45530,
    n45531, n45532, n45533, n45534, n45535, n45536,
    n45537, n45538, n45539, n45540, n45541, n45542,
    n45543, n45544, n45545, n45546, n45547, n45548,
    n45549, n45550, n45551, n45552, n45553, n45554,
    n45555, n45556, n45557, n45558, n45559, n45560,
    n45561, n45562, n45563, n45564, n45565, n45566,
    n45567, n45568, n45569, n45570, n45571, n45572,
    n45573, n45574, n45575, n45576, n45577, n45578,
    n45579, n45580, n45581, n45582, n45583, n45584,
    n45585, n45586, n45587, n45588, n45589, n45590,
    n45591, n45592, n45593, n45594, n45595, n45596,
    n45597, n45598, n45599, n45600, n45601, n45602,
    n45603, n45604, n45605, n45606, n45607, n45608,
    n45609, n45610, n45611, n45612, n45613, n45614,
    n45615, n45616, n45617, n45618, n45619, n45620,
    n45621, n45622, n45623, n45624, n45625, n45626,
    n45627, n45628, n45629, n45630, n45631, n45632,
    n45633, n45634, n45635, n45636, n45637, n45638,
    n45639, n45640, n45641, n45642, n45643, n45644,
    n45645, n45646, n45647, n45648, n45649, n45650,
    n45651, n45652, n45653, n45654, n45655, n45656,
    n45657, n45658, n45659, n45660, n45661, n45662,
    n45663, n45664, n45665, n45666, n45667, n45668,
    n45669, n45670, n45671, n45672, n45673, n45674,
    n45675, n45676, n45677, n45678, n45679, n45680,
    n45681, n45682, n45683, n45684, n45685, n45686,
    n45687, n45688, n45689, n45690, n45691, n45692,
    n45693, n45694, n45695, n45696, n45697, n45698,
    n45699, n45700, n45701, n45702, n45703, n45704,
    n45705, n45706, n45707, n45708, n45709, n45710,
    n45711, n45712, n45713, n45714, n45715, n45716,
    n45717, n45718, n45719, n45720, n45721, n45722,
    n45723, n45724, n45725, n45726, n45727, n45728,
    n45729, n45730, n45731, n45732, n45733, n45734,
    n45735, n45736, n45737, n45738, n45739, n45740,
    n45741, n45742, n45743, n45744, n45745, n45746,
    n45747, n45748, n45749, n45750, n45751, n45752,
    n45753, n45754, n45755, n45756, n45757, n45758,
    n45759, n45760, n45761, n45762, n45763, n45764,
    n45765, n45766, n45767, n45768, n45769, n45770,
    n45771, n45772, n45773, n45774, n45775, n45776,
    n45777, n45778, n45779, n45780, n45781, n45782,
    n45783, n45784, n45785, n45786, n45787, n45788,
    n45789, n45790, n45791, n45792, n45793, n45794,
    n45795, n45796, n45797, n45798, n45799, n45800,
    n45801, n45802, n45803, n45804, n45805, n45806,
    n45807, n45808, n45809, n45810, n45811, n45812,
    n45813, n45814, n45815, n45816, n45817, n45818,
    n45819, n45820, n45821, n45822, n45823, n45824,
    n45825, n45826, n45827, n45828, n45829, n45830,
    n45831, n45832, n45833, n45834, n45835, n45836,
    n45837, n45838, n45839, n45840, n45841, n45842,
    n45843, n45844, n45845, n45846, n45847, n45848,
    n45849, n45850, n45851, n45852, n45853, n45854,
    n45855, n45856, n45857, n45858, n45859, n45860,
    n45861, n45862, n45863, n45864, n45865, n45866,
    n45867, n45868, n45869, n45870, n45871, n45872,
    n45873, n45874, n45875, n45876, n45877, n45878,
    n45879, n45880, n45881, n45882, n45883, n45884,
    n45885, n45886, n45887, n45888, n45889, n45890,
    n45891, n45892, n45893, n45894, n45895, n45896,
    n45897, n45898, n45899, n45900, n45901, n45902,
    n45903, n45904, n45905, n45906, n45907, n45908,
    n45909, n45910, n45911, n45912, n45913, n45914,
    n45915, n45916, n45917, n45918, n45919, n45920,
    n45921, n45922, n45923, n45924, n45925, n45926,
    n45927, n45928, n45929, n45930, n45931, n45932,
    n45933, n45934, n45935, n45936, n45937, n45938,
    n45939, n45940, n45941, n45942, n45943, n45944,
    n45945, n45946, n45947, n45948, n45949, n45950,
    n45951, n45952, n45953, n45954, n45955, n45956,
    n45957, n45958, n45959, n45960, n45961, n45962,
    n45963, n45964, n45965, n45966, n45967, n45968,
    n45969, n45970, n45971, n45972, n45973, n45974,
    n45975, n45976, n45977, n45978, n45979, n45980,
    n45981, n45982, n45983, n45984, n45985, n45986,
    n45987, n45988, n45989, n45990, n45991, n45992,
    n45993, n45994, n45995, n45996, n45997, n45998,
    n45999, n46000, n46001, n46002, n46003, n46004,
    n46005, n46006, n46007, n46008, n46009, n46010,
    n46011, n46012, n46013, n46014, n46015, n46016,
    n46017, n46018, n46019, n46020, n46021, n46022,
    n46023, n46024, n46025, n46026, n46027, n46028,
    n46029, n46030, n46031, n46032, n46033, n46034,
    n46035, n46036, n46037, n46038, n46039, n46040,
    n46041, n46042, n46043, n46044, n46045, n46046,
    n46047, n46048, n46049, n46050, n46051, n46052,
    n46053, n46054, n46055, n46056, n46057, n46058,
    n46059, n46060, n46061, n46062, n46063, n46064,
    n46065, n46066, n46067, n46068, n46069, n46070,
    n46071, n46072, n46073, n46074, n46075, n46076,
    n46077, n46078, n46079, n46080, n46081, n46082,
    n46083, n46084, n46085, n46086, n46087, n46088,
    n46089, n46090, n46091, n46092, n46093, n46094,
    n46095, n46096, n46097, n46098, n46099, n46100,
    n46101, n46102, n46103, n46104, n46105, n46106,
    n46107, n46108, n46109, n46110, n46111, n46112,
    n46113, n46114, n46115, n46116, n46117, n46118,
    n46119, n46120, n46121, n46122, n46123, n46124,
    n46125, n46126, n46127, n46128, n46129, n46130,
    n46131, n46132, n46133, n46134, n46135, n46136,
    n46137, n46138, n46139, n46140, n46141, n46142,
    n46143, n46144, n46145, n46146, n46147, n46148,
    n46149, n46150, n46151, n46152, n46153, n46154,
    n46155, n46156, n46157, n46158, n46159, n46160,
    n46161, n46162, n46163, n46164, n46165, n46166,
    n46167, n46168, n46169, n46170, n46171, n46172,
    n46173, n46174, n46175, n46176, n46177, n46178,
    n46179, n46180, n46181, n46182, n46183, n46184,
    n46185, n46186, n46187, n46188, n46189, n46190,
    n46191, n46192, n46193, n46194, n46195, n46196,
    n46197, n46198, n46199, n46200, n46201, n46202,
    n46203, n46204, n46205, n46206, n46207, n46208,
    n46209, n46210, n46211, n46212, n46213, n46214,
    n46215, n46216, n46217, n46218, n46219, n46220,
    n46221, n46222, n46223, n46224, n46225, n46226,
    n46227, n46228, n46229, n46230, n46231, n46232,
    n46233, n46234, n46235, n46236, n46237, n46238,
    n46239, n46240, n46241, n46242, n46243, n46244,
    n46245, n46246, n46247, n46248, n46249, n46250,
    n46251, n46252, n46253, n46254, n46255, n46256,
    n46257, n46258, n46259, n46260, n46261, n46262,
    n46263, n46264, n46265, n46266, n46267, n46268,
    n46269, n46270, n46271, n46272, n46273, n46274,
    n46275, n46276, n46277, n46278, n46279, n46280,
    n46281, n46282, n46283, n46284, n46285, n46286,
    n46287, n46288, n46289, n46290, n46291, n46292,
    n46293, n46294, n46295, n46296, n46297, n46298,
    n46299, n46300, n46301, n46302, n46303, n46304,
    n46305, n46306, n46307, n46308, n46309, n46310,
    n46311, n46312, n46313, n46314, n46315, n46316,
    n46317, n46318, n46319, n46320, n46321, n46322,
    n46323, n46324, n46325, n46326, n46327, n46328,
    n46329, n46330, n46331, n46332, n46333, n46334,
    n46335, n46336, n46337, n46338, n46339, n46340,
    n46341, n46342, n46343, n46344, n46345, n46346,
    n46347, n46348, n46349, n46350, n46351, n46352,
    n46353, n46354, n46355, n46356, n46357, n46358,
    n46359, n46360, n46361, n46362, n46363, n46364,
    n46365, n46366, n46367, n46368, n46369, n46370,
    n46371, n46372, n46373, n46374, n46375, n46376,
    n46377, n46378, n46379, n46380, n46381, n46382,
    n46383, n46384, n46385, n46386, n46387, n46388,
    n46389, n46390, n46391, n46392, n46393, n46394,
    n46395, n46396, n46397, n46398, n46399, n46400,
    n46401, n46402, n46403, n46404, n46405, n46406,
    n46407, n46408, n46409, n46410, n46411, n46412,
    n46413, n46414, n46415, n46416, n46417, n46418,
    n46419, n46420, n46421, n46422, n46423, n46424,
    n46425, n46426, n46427, n46428, n46429, n46430,
    n46431, n46432, n46433, n46434, n46435, n46436,
    n46437, n46438, n46439, n46440, n46441, n46442,
    n46443, n46444, n46445, n46446, n46447, n46449,
    n46450, n46451, n46452, n46453, n46454, n46455,
    n46456, n46457, n46458, n46459, n46460, n46461,
    n46462, n46463, n46464, n46465, n46466, n46467,
    n46468, n46469, n46470, n46471, n46472, n46473,
    n46474, n46475, n46476, n46477, n46478, n46479,
    n46480, n46481, n46482, n46483, n46484, n46485,
    n46486, n46487, n46488, n46489, n46490, n46491,
    n46492, n46493, n46494, n46495, n46496, n46497,
    n46498, n46499, n46500, n46501, n46502, n46503,
    n46504, n46505, n46506, n46507, n46508, n46509,
    n46510, n46511, n46512, n46513, n46514, n46515,
    n46516, n46517, n46518, n46519, n46520, n46521,
    n46522, n46523, n46524, n46525, n46526, n46527,
    n46528, n46529, n46530, n46531, n46532, n46533,
    n46534, n46535, n46536, n46537, n46538, n46539,
    n46540, n46541, n46542, n46543, n46544, n46545,
    n46546, n46547, n46548, n46549, n46550, n46551,
    n46552, n46553, n46554, n46555, n46556, n46557,
    n46558, n46559, n46560, n46561, n46562, n46563,
    n46564, n46565, n46566, n46567, n46568, n46569,
    n46570, n46571, n46572, n46573, n46574, n46575,
    n46576, n46577, n46578, n46579, n46580, n46581,
    n46582, n46583, n46584, n46585, n46586, n46587,
    n46588, n46589, n46590, n46591, n46592, n46593,
    n46594, n46595, n46596, n46597, n46598, n46599,
    n46600, n46601, n46602, n46603, n46604, n46605,
    n46606, n46607, n46608, n46609, n46610, n46611,
    n46612, n46613, n46614, n46615, n46616, n46617,
    n46618, n46619, n46620, n46621, n46622, n46623,
    n46624, n46625, n46626, n46627, n46628, n46629,
    n46630, n46631, n46632, n46633, n46634, n46635,
    n46636, n46637, n46638, n46639, n46640, n46641,
    n46642, n46643, n46644, n46645, n46646, n46647,
    n46648, n46649, n46650, n46651, n46652, n46653,
    n46654, n46655, n46656, n46657, n46658, n46659,
    n46660, n46661, n46662, n46663, n46664, n46665,
    n46666, n46667, n46668, n46669, n46670, n46671,
    n46672, n46673, n46674, n46675, n46676, n46677,
    n46678, n46679, n46680, n46681, n46682, n46683,
    n46684, n46685, n46686, n46687, n46688, n46689,
    n46690, n46691, n46692, n46693, n46694, n46695,
    n46696, n46697, n46698, n46699, n46700, n46701,
    n46702, n46703, n46704, n46705, n46706, n46707,
    n46708, n46709, n46710, n46711, n46712, n46713,
    n46714, n46715, n46716, n46717, n46718, n46719,
    n46720, n46721, n46722, n46723, n46724, n46725,
    n46726, n46727, n46728, n46729, n46730, n46731,
    n46732, n46733, n46734, n46735, n46736, n46737,
    n46738, n46739, n46740, n46741, n46742, n46743,
    n46744, n46745, n46746, n46747, n46748, n46749,
    n46750, n46751, n46752, n46753, n46754, n46755,
    n46756, n46757, n46758, n46759, n46760, n46761,
    n46762, n46763, n46764, n46765, n46766, n46767,
    n46768, n46769, n46770, n46771, n46772, n46773,
    n46774, n46775, n46776, n46777, n46778, n46779,
    n46780, n46781, n46782, n46783, n46784, n46785,
    n46786, n46787, n46788, n46789, n46790, n46791,
    n46792, n46793, n46794, n46795, n46796, n46797,
    n46798, n46799, n46800, n46801, n46802, n46803,
    n46804, n46805, n46806, n46807, n46808, n46809,
    n46810, n46811, n46812, n46813, n46814, n46815,
    n46816, n46817, n46818, n46819, n46820, n46821,
    n46822, n46823, n46824, n46825, n46826, n46828,
    n46829, n46830, n46831, n46832, n46833, n46834,
    n46835, n46836, n46837, n46838, n46839, n46840,
    n46841, n46842, n46843, n46844, n46845, n46846,
    n46847, n46848, n46849, n46850, n46851, n46852,
    n46853, n46854, n46855, n46856, n46857, n46858,
    n46859, n46860, n46861, n46862, n46863, n46864,
    n46865, n46866, n46867, n46868, n46869, n46870,
    n46871, n46872, n46873, n46874, n46875, n46876,
    n46877, n46878, n46879, n46880, n46881, n46882,
    n46883, n46884, n46885, n46886, n46887, n46888,
    n46889, n46890, n46891, n46892, n46893, n46894,
    n46895, n46896, n46897, n46898, n46899, n46900,
    n46901, n46902, n46903, n46904, n46905, n46906,
    n46907, n46908, n46909, n46910, n46911, n46912,
    n46913, n46914, n46915, n46916, n46917, n46918,
    n46919, n46920, n46921, n46922, n46923, n46924,
    n46925, n46926, n46927, n46928, n46929, n46930,
    n46931, n46932, n46933, n46934, n46935, n46936,
    n46937, n46938, n46939, n46940, n46941, n46942,
    n46943, n46944, n46945, n46946, n46947, n46948,
    n46949, n46950, n46951, n46952, n46953, n46954,
    n46955, n46956, n46957, n46958, n46959, n46960,
    n46961, n46962, n46963, n46964, n46965, n46966,
    n46967, n46968, n46969, n46970, n46971, n46972,
    n46973, n46974, n46975, n46976, n46977, n46978,
    n46979, n46980, n46981, n46982, n46983, n46984,
    n46985, n46986, n46987, n46988, n46989, n46990,
    n46991, n46992, n46993, n46994, n46995, n46996,
    n46997, n46998, n46999, n47000, n47001, n47002,
    n47003, n47004, n47005, n47006, n47007, n47008,
    n47009, n47010, n47011, n47012, n47013, n47014,
    n47015, n47016, n47017, n47018, n47019, n47020,
    n47021, n47022, n47023, n47024, n47025, n47026,
    n47027, n47028, n47029, n47030, n47031, n47032,
    n47033, n47034, n47035, n47036, n47037, n47038,
    n47039, n47040, n47041, n47042, n47043, n47044,
    n47045, n47046, n47047, n47048, n47049, n47050,
    n47051, n47052, n47053, n47054, n47055, n47056,
    n47057, n47058, n47059, n47060, n47061, n47062,
    n47063, n47064, n47065, n47066, n47067, n47068,
    n47069, n47070, n47071, n47072, n47073, n47074,
    n47075, n47076, n47077, n47078, n47079, n47080,
    n47081, n47082, n47083, n47084, n47085, n47086,
    n47087, n47088, n47089, n47090, n47091, n47092,
    n47093, n47094, n47095, n47096, n47097, n47098,
    n47099, n47100, n47101, n47102, n47103, n47104,
    n47105, n47106, n47107, n47108, n47109, n47110,
    n47111, n47112, n47113, n47114, n47115, n47116,
    n47117, n47118, n47119, n47120, n47121, n47122,
    n47123, n47124, n47125, n47126, n47127, n47128,
    n47129, n47130, n47131, n47132, n47133, n47134,
    n47135, n47136, n47137, n47138, n47139, n47140,
    n47141, n47142, n47143, n47144, n47145, n47146,
    n47147, n47148, n47149, n47150, n47151, n47152,
    n47153, n47154, n47155, n47156, n47157, n47158,
    n47159, n47161, n47162, n47163, n47164, n47165,
    n47166, n47167, n47168, n47169, n47170, n47171,
    n47172, n47173, n47174, n47175, n47176, n47177,
    n47178, n47179, n47180, n47181, n47182, n47183,
    n47184, n47185, n47186, n47187, n47188, n47189,
    n47190, n47191, n47192, n47193, n47194, n47195,
    n47196, n47197, n47198, n47199, n47200, n47201,
    n47202, n47203, n47204, n47205, n47206, n47207,
    n47208, n47209, n47210, n47211, n47212, n47213,
    n47214, n47215, n47216, n47217, n47218, n47219,
    n47220, n47221, n47222, n47223, n47224, n47225,
    n47226, n47227, n47228, n47229, n47230, n47231,
    n47232, n47233, n47234, n47235, n47236, n47237,
    n47238, n47239, n47240, n47241, n47242, n47243,
    n47244, n47245, n47246, n47247, n47248, n47249,
    n47250, n47251, n47252, n47253, n47254, n47255,
    n47256, n47257, n47258, n47259, n47260, n47261,
    n47262, n47263, n47264, n47265, n47266, n47267,
    n47268, n47269, n47270, n47271, n47272, n47273,
    n47274, n47275, n47276, n47277, n47278, n47279,
    n47280, n47281, n47282, n47283, n47284, n47285,
    n47286, n47287, n47288, n47289, n47290, n47291,
    n47292, n47293, n47294, n47295, n47296, n47297,
    n47298, n47299, n47300, n47301, n47302, n47303,
    n47304, n47305, n47306, n47307, n47308, n47309,
    n47310, n47311, n47312, n47313, n47314, n47315,
    n47316, n47317, n47318, n47319, n47320, n47321,
    n47322, n47323, n47324, n47325, n47326, n47327,
    n47328, n47329, n47330, n47331, n47332, n47333,
    n47334, n47335, n47336, n47337, n47338, n47339,
    n47340, n47341, n47342, n47343, n47344, n47345,
    n47346, n47347, n47348, n47349, n47350, n47351,
    n47352, n47353, n47354, n47355, n47356, n47357,
    n47358, n47359, n47360, n47361, n47362, n47363,
    n47364, n47365, n47366, n47367, n47368, n47369,
    n47370, n47371, n47372, n47373, n47374, n47375,
    n47376, n47377, n47378, n47379, n47380, n47381,
    n47382, n47383, n47384, n47385, n47386, n47387,
    n47388, n47389, n47390, n47391, n47392, n47393,
    n47394, n47395, n47396, n47397, n47398, n47399,
    n47400, n47401, n47402, n47403, n47404, n47405,
    n47406, n47407, n47408, n47409, n47410, n47411,
    n47412, n47413, n47414, n47415, n47416, n47417,
    n47418, n47419, n47420, n47421, n47422, n47423,
    n47424, n47425, n47426, n47427, n47428, n47429,
    n47430, n47431, n47432, n47433, n47434, n47435,
    n47436, n47437, n47438, n47439, n47440, n47441,
    n47442, n47443, n47444, n47445, n47446, n47447,
    n47448, n47449, n47450, n47451, n47452, n47453,
    n47454, n47455, n47456, n47457, n47458, n47459,
    n47460, n47461, n47462, n47463, n47464, n47465,
    n47466, n47467, n47468, n47469, n47470, n47471,
    n47472, n47473, n47474, n47475, n47476, n47477,
    n47478, n47479, n47480, n47481, n47482, n47483,
    n47484, n47485, n47486, n47487, n47488, n47489,
    n47490, n47491, n47492, n47493, n47494, n47495,
    n47496, n47497, n47498, n47499, n47500, n47501,
    n47502, n47503, n47504, n47505, n47506, n47507,
    n47508, n47509, n47510, n47511, n47512, n47513,
    n47514, n47515, n47516, n47517, n47518, n47519,
    n47520, n47521, n47522, n47523, n47524, n47525,
    n47526, n47527, n47528, n47529, n47530, n47531,
    n47532, n47533, n47534, n47535, n47536, n47537,
    n47538, n47539, n47540, n47541, n47542, n47543,
    n47544, n47545, n47547, n47548, n47549, n47550,
    n47551, n47552, n47553, n47554, n47555, n47556,
    n47557, n47558, n47559, n47560, n47561, n47562,
    n47563, n47564, n47565, n47566, n47567, n47568,
    n47569, n47570, n47571, n47572, n47573, n47574,
    n47575, n47576, n47577, n47578, n47579, n47580,
    n47581, n47582, n47583, n47584, n47585, n47586,
    n47587, n47588, n47589, n47590, n47591, n47592,
    n47593, n47594, n47595, n47596, n47597, n47598,
    n47599, n47600, n47601, n47602, n47603, n47604,
    n47605, n47606, n47607, n47608, n47609, n47610,
    n47611, n47612, n47613, n47614, n47615, n47616,
    n47617, n47618, n47619, n47620, n47621, n47622,
    n47623, n47624, n47625, n47626, n47627, n47628,
    n47629, n47630, n47631, n47632, n47633, n47634,
    n47635, n47636, n47637, n47638, n47639, n47640,
    n47641, n47642, n47643, n47644, n47645, n47646,
    n47647, n47648, n47649, n47650, n47651, n47652,
    n47653, n47654, n47655, n47656, n47657, n47658,
    n47659, n47660, n47661, n47662, n47663, n47664,
    n47665, n47666, n47667, n47668, n47669, n47670,
    n47671, n47672, n47673, n47674, n47675, n47676,
    n47677, n47678, n47679, n47680, n47681, n47682,
    n47683, n47684, n47685, n47686, n47687, n47688,
    n47689, n47690, n47691, n47692, n47693, n47694,
    n47695, n47696, n47697, n47698, n47699, n47700,
    n47701, n47702, n47703, n47704, n47705, n47706,
    n47707, n47708, n47709, n47710, n47711, n47712,
    n47713, n47714, n47715, n47716, n47717, n47718,
    n47719, n47720, n47721, n47722, n47723, n47724,
    n47725, n47726, n47727, n47728, n47729, n47730,
    n47731, n47732, n47733, n47734, n47735, n47736,
    n47737, n47738, n47739, n47740, n47741, n47742,
    n47743, n47744, n47745, n47746, n47747, n47748,
    n47749, n47750, n47751, n47752, n47753, n47754,
    n47755, n47756, n47757, n47758, n47759, n47760,
    n47761, n47762, n47763, n47764, n47765, n47766,
    n47767, n47768, n47769, n47770, n47771, n47772,
    n47773, n47774, n47775, n47776, n47777, n47778,
    n47779, n47780, n47781, n47782, n47783, n47784,
    n47785, n47786, n47787, n47788, n47789, n47790,
    n47791, n47792, n47793, n47794, n47795, n47796,
    n47797, n47798, n47799, n47800, n47801, n47802,
    n47803, n47804, n47805, n47806, n47807, n47808,
    n47809, n47810, n47811, n47812, n47813, n47814,
    n47815, n47816, n47817, n47818, n47819, n47820,
    n47821, n47822, n47823, n47824, n47825, n47826,
    n47827, n47828, n47829, n47830, n47831, n47832,
    n47833, n47834, n47835, n47836, n47837, n47838,
    n47839, n47840, n47841, n47842, n47843, n47844,
    n47845, n47846, n47847, n47848, n47849, n47850,
    n47851, n47852, n47853, n47854, n47855, n47856,
    n47857, n47858, n47859, n47860, n47861, n47862,
    n47863, n47864, n47865, n47866, n47867, n47868,
    n47869, n47870, n47871, n47872, n47873, n47874,
    n47875, n47876, n47877, n47878, n47879, n47880,
    n47881, n47882, n47883, n47884, n47886, n47887,
    n47888, n47889, n47890, n47891, n47892, n47893,
    n47894, n47895, n47896, n47897, n47898, n47899,
    n47900, n47901, n47902, n47903, n47904, n47905,
    n47906, n47907, n47908, n47909, n47910, n47911,
    n47912, n47913, n47914, n47915, n47916, n47917,
    n47918, n47919, n47920, n47921, n47922, n47923,
    n47924, n47925, n47926, n47927, n47928, n47929,
    n47930, n47931, n47932, n47933, n47934, n47935,
    n47936, n47937, n47938, n47939, n47940, n47941,
    n47942, n47943, n47944, n47945, n47946, n47947,
    n47948, n47949, n47950, n47951, n47952, n47953,
    n47954, n47955, n47956, n47957, n47958, n47959,
    n47960, n47961, n47962, n47963, n47964, n47965,
    n47966, n47967, n47968, n47969, n47970, n47971,
    n47972, n47973, n47974, n47975, n47976, n47977,
    n47978, n47979, n47980, n47981, n47982, n47983,
    n47984, n47985, n47986, n47987, n47988, n47989,
    n47990, n47991, n47992, n47993, n47994, n47995,
    n47996, n47997, n47998, n47999, n48000, n48001,
    n48002, n48003, n48004, n48005, n48006, n48007,
    n48008, n48009, n48010, n48011, n48012, n48013,
    n48014, n48015, n48016, n48017, n48018, n48019,
    n48020, n48021, n48022, n48023, n48024, n48025,
    n48026, n48027, n48028, n48029, n48030, n48031,
    n48032, n48033, n48034, n48035, n48036, n48037,
    n48038, n48039, n48040, n48041, n48042, n48043,
    n48044, n48045, n48046, n48047, n48048, n48049,
    n48050, n48051, n48052, n48053, n48054, n48055,
    n48056, n48057, n48058, n48059, n48060, n48061,
    n48062, n48063, n48064, n48065, n48066, n48067,
    n48068, n48069, n48070, n48071, n48072, n48073,
    n48074, n48075, n48076, n48077, n48078, n48079,
    n48080, n48081, n48082, n48083, n48084, n48085,
    n48086, n48087, n48088, n48089, n48090, n48091,
    n48092, n48093, n48094, n48095, n48096, n48097,
    n48098, n48099, n48100, n48101, n48102, n48103,
    n48104, n48105, n48106, n48107, n48108, n48109,
    n48110, n48111, n48112, n48113, n48114, n48115,
    n48116, n48117, n48118, n48119, n48120, n48121,
    n48122, n48123, n48124, n48125, n48126, n48127,
    n48128, n48129, n48130, n48131, n48132, n48133,
    n48134, n48135, n48136, n48137, n48138, n48139,
    n48140, n48141, n48142, n48143, n48144, n48145,
    n48146, n48147, n48148, n48149, n48150, n48151,
    n48152, n48153, n48154, n48155, n48156, n48157,
    n48158, n48159, n48160, n48161, n48162, n48163,
    n48164, n48165, n48166, n48167, n48168, n48169,
    n48170, n48171, n48172, n48173, n48174, n48175,
    n48176, n48177, n48178, n48179, n48180, n48181,
    n48182, n48183, n48184, n48185, n48186, n48187,
    n48188, n48189, n48190, n48191, n48192, n48193,
    n48194, n48195, n48196, n48197, n48198, n48199,
    n48200, n48201, n48202, n48203, n48204, n48205,
    n48206, n48207, n48208, n48209, n48210, n48211,
    n48212, n48213, n48214, n48215, n48216, n48217,
    n48218, n48220, n48221, n48222, n48223, n48224,
    n48225, n48226, n48227, n48228, n48229, n48230,
    n48231, n48232, n48233, n48234, n48235, n48236,
    n48237, n48238, n48239, n48240, n48241, n48242,
    n48243, n48244, n48245, n48246, n48247, n48248,
    n48249, n48250, n48251, n48252, n48253, n48254,
    n48255, n48256, n48257, n48258, n48259, n48260,
    n48261, n48262, n48263, n48264, n48265, n48266,
    n48267, n48268, n48269, n48270, n48271, n48272,
    n48273, n48274, n48275, n48276, n48277, n48278,
    n48279, n48280, n48281, n48282, n48283, n48284,
    n48285, n48286, n48287, n48288, n48289, n48290,
    n48291, n48292, n48293, n48294, n48295, n48296,
    n48297, n48298, n48299, n48300, n48301, n48302,
    n48303, n48304, n48305, n48306, n48307, n48308,
    n48309, n48310, n48311, n48312, n48313, n48314,
    n48315, n48316, n48317, n48318, n48319, n48320,
    n48321, n48322, n48323, n48324, n48325, n48326,
    n48327, n48328, n48329, n48330, n48331, n48332,
    n48333, n48334, n48335, n48336, n48337, n48338,
    n48339, n48340, n48341, n48342, n48343, n48344,
    n48345, n48346, n48347, n48348, n48349, n48350,
    n48351, n48352, n48353, n48354, n48355, n48356,
    n48357, n48358, n48359, n48360, n48361, n48362,
    n48363, n48364, n48365, n48366, n48367, n48368,
    n48369, n48370, n48371, n48372, n48373, n48374,
    n48375, n48376, n48377, n48378, n48379, n48380,
    n48381, n48382, n48383, n48384, n48385, n48386,
    n48387, n48388, n48389, n48390, n48391, n48392,
    n48393, n48394, n48395, n48396, n48397, n48398,
    n48399, n48400, n48401, n48402, n48403, n48404,
    n48405, n48406, n48407, n48408, n48409, n48410,
    n48411, n48412, n48413, n48414, n48415, n48416,
    n48417, n48418, n48419, n48420, n48421, n48422,
    n48423, n48424, n48425, n48426, n48427, n48428,
    n48429, n48430, n48431, n48432, n48433, n48434,
    n48435, n48436, n48437, n48438, n48439, n48440,
    n48441, n48442, n48443, n48444, n48445, n48446,
    n48447, n48448, n48449, n48450, n48451, n48452,
    n48453, n48454, n48455, n48456, n48457, n48458,
    n48459, n48460, n48461, n48462, n48463, n48464,
    n48465, n48466, n48467, n48468, n48469, n48470,
    n48471, n48472, n48473, n48474, n48475, n48476,
    n48477, n48478, n48479, n48480, n48481, n48482,
    n48483, n48484, n48485, n48486, n48487, n48488,
    n48489, n48490, n48491, n48492, n48493, n48494,
    n48495, n48496, n48497, n48498, n48499, n48500,
    n48501, n48502, n48503, n48504, n48505, n48506,
    n48508, n48509, n48510, n48511, n48512, n48513,
    n48514, n48515, n48516, n48517, n48518, n48519,
    n48520, n48521, n48522, n48523, n48524, n48525,
    n48526, n48527, n48528, n48529, n48530, n48531,
    n48532, n48533, n48534, n48535, n48536, n48537,
    n48538, n48539, n48540, n48541, n48542, n48543,
    n48544, n48545, n48546, n48547, n48548, n48549,
    n48550, n48551, n48552, n48553, n48554, n48555,
    n48556, n48557, n48558, n48559, n48560, n48561,
    n48562, n48563, n48564, n48565, n48566, n48567,
    n48568, n48569, n48570, n48571, n48572, n48573,
    n48574, n48575, n48576, n48577, n48578, n48579,
    n48580, n48581, n48582, n48583, n48584, n48585,
    n48586, n48587, n48588, n48589, n48590, n48591,
    n48592, n48593, n48594, n48595, n48596, n48597,
    n48598, n48599, n48600, n48601, n48602, n48603,
    n48604, n48605, n48606, n48607, n48608, n48609,
    n48610, n48611, n48612, n48613, n48614, n48615,
    n48616, n48617, n48618, n48619, n48620, n48621,
    n48622, n48623, n48624, n48625, n48626, n48627,
    n48628, n48629, n48630, n48631, n48632, n48633,
    n48634, n48635, n48636, n48637, n48638, n48639,
    n48640, n48641, n48642, n48643, n48644, n48645,
    n48646, n48647, n48648, n48649, n48650, n48651,
    n48652, n48653, n48654, n48655, n48656, n48657,
    n48658, n48659, n48660, n48661, n48662, n48663,
    n48664, n48665, n48666, n48667, n48668, n48669,
    n48670, n48671, n48672, n48673, n48674, n48675,
    n48676, n48677, n48678, n48679, n48680, n48681,
    n48682, n48683, n48684, n48685, n48686, n48687,
    n48688, n48689, n48690, n48691, n48692, n48693,
    n48694, n48695, n48696, n48697, n48698, n48699,
    n48700, n48701, n48702, n48703, n48704, n48705,
    n48706, n48707, n48708, n48709, n48710, n48711,
    n48712, n48713, n48714, n48715, n48716, n48717,
    n48718, n48719, n48720, n48721, n48722, n48723,
    n48724, n48725, n48726, n48727, n48728, n48729,
    n48730, n48731, n48732, n48733, n48734, n48735,
    n48736, n48737, n48738, n48739, n48740, n48741,
    n48742, n48743, n48744, n48745, n48746, n48747,
    n48748, n48749, n48750, n48751, n48752, n48753,
    n48754, n48755, n48756, n48757, n48758, n48759,
    n48760, n48761, n48762, n48763, n48764, n48765,
    n48766, n48767, n48768, n48769, n48770, n48771,
    n48772, n48773, n48774, n48775, n48776, n48777,
    n48778, n48779, n48780, n48781, n48782, n48783,
    n48784, n48785, n48786, n48787, n48788, n48789,
    n48790, n48791, n48792, n48793, n48794, n48795,
    n48796, n48797, n48798, n48799, n48800, n48801,
    n48802, n48803, n48804, n48805, n48806, n48807,
    n48808, n48809, n48810, n48811, n48812, n48813,
    n48814, n48815, n48816, n48817, n48818, n48819,
    n48820, n48821, n48822, n48823, n48824, n48825,
    n48826, n48827, n48829, n48830, n48831, n48832,
    n48833, n48834, n48835, n48836, n48837, n48838,
    n48839, n48840, n48841, n48842, n48843, n48844,
    n48845, n48846, n48847, n48848, n48849, n48850,
    n48851, n48852, n48853, n48854, n48855, n48856,
    n48857, n48858, n48859, n48860, n48861, n48862,
    n48863, n48864, n48865, n48866, n48867, n48868,
    n48869, n48870, n48871, n48872, n48873, n48874,
    n48875, n48876, n48877, n48878, n48879, n48880,
    n48881, n48882, n48883, n48884, n48885, n48886,
    n48887, n48888, n48889, n48890, n48891, n48892,
    n48893, n48894, n48895, n48896, n48897, n48898,
    n48899, n48900, n48901, n48902, n48903, n48904,
    n48905, n48906, n48907, n48908, n48909, n48910,
    n48911, n48912, n48913, n48914, n48915, n48916,
    n48917, n48918, n48919, n48920, n48921, n48922,
    n48923, n48924, n48925, n48926, n48927, n48928,
    n48929, n48930, n48931, n48932, n48933, n48934,
    n48935, n48936, n48937, n48938, n48939, n48940,
    n48941, n48942, n48943, n48944, n48945, n48946,
    n48947, n48948, n48949, n48950, n48951, n48952,
    n48953, n48954, n48955, n48956, n48957, n48958,
    n48959, n48960, n48961, n48962, n48963, n48964,
    n48965, n48966, n48967, n48968, n48969, n48970,
    n48971, n48972, n48973, n48974, n48975, n48976,
    n48977, n48978, n48979, n48980, n48981, n48982,
    n48983, n48984, n48985, n48986, n48987, n48988,
    n48989, n48990, n48991, n48992, n48993, n48994,
    n48995, n48996, n48997, n48998, n48999, n49000,
    n49001, n49002, n49003, n49004, n49005, n49006,
    n49007, n49008, n49009, n49010, n49011, n49012,
    n49013, n49014, n49015, n49016, n49017, n49018,
    n49019, n49020, n49021, n49022, n49023, n49024,
    n49025, n49026, n49027, n49028, n49029, n49030,
    n49031, n49032, n49033, n49034, n49035, n49036,
    n49037, n49038, n49039, n49040, n49041, n49042,
    n49043, n49044, n49045, n49046, n49047, n49048,
    n49049, n49050, n49051, n49052, n49053, n49054,
    n49055, n49056, n49057, n49058, n49059, n49060,
    n49061, n49062, n49063, n49064, n49065, n49066,
    n49067, n49068, n49069, n49070, n49071, n49072,
    n49073, n49074, n49075, n49076, n49077, n49078,
    n49079, n49080, n49081, n49082, n49083, n49084,
    n49085, n49086, n49087, n49088, n49089, n49090,
    n49091, n49092, n49093, n49094, n49095, n49096,
    n49097, n49098, n49099, n49100, n49101, n49102,
    n49103, n49104, n49105, n49106, n49107, n49108,
    n49109, n49110, n49111, n49112, n49113, n49114,
    n49115, n49116, n49117, n49119, n49120, n49121,
    n49122, n49123, n49124, n49125, n49126, n49127,
    n49128, n49129, n49130, n49131, n49132, n49133,
    n49134, n49135, n49136, n49137, n49138, n49139,
    n49140, n49141, n49142, n49143, n49144, n49145,
    n49146, n49147, n49148, n49149, n49150, n49151,
    n49152, n49153, n49154, n49155, n49156, n49157,
    n49158, n49159, n49160, n49161, n49162, n49163,
    n49164, n49165, n49166, n49167, n49168, n49169,
    n49170, n49171, n49172, n49173, n49174, n49175,
    n49176, n49177, n49178, n49179, n49180, n49181,
    n49182, n49183, n49184, n49185, n49186, n49187,
    n49188, n49189, n49190, n49191, n49192, n49193,
    n49194, n49195, n49196, n49197, n49198, n49199,
    n49200, n49201, n49202, n49203, n49204, n49205,
    n49206, n49207, n49208, n49209, n49210, n49211,
    n49212, n49213, n49214, n49215, n49216, n49217,
    n49218, n49219, n49220, n49221, n49222, n49223,
    n49224, n49225, n49226, n49227, n49228, n49229,
    n49230, n49231, n49232, n49233, n49234, n49235,
    n49236, n49237, n49238, n49239, n49240, n49241,
    n49242, n49243, n49244, n49245, n49246, n49247,
    n49248, n49249, n49250, n49251, n49252, n49253,
    n49254, n49255, n49256, n49257, n49258, n49259,
    n49260, n49261, n49262, n49263, n49264, n49265,
    n49266, n49267, n49268, n49269, n49270, n49271,
    n49272, n49273, n49274, n49275, n49276, n49277,
    n49278, n49279, n49280, n49281, n49282, n49283,
    n49284, n49285, n49286, n49287, n49288, n49289,
    n49290, n49291, n49292, n49293, n49294, n49295,
    n49296, n49297, n49298, n49299, n49300, n49301,
    n49302, n49303, n49304, n49305, n49306, n49307,
    n49308, n49309, n49310, n49311, n49312, n49313,
    n49314, n49315, n49316, n49317, n49318, n49319,
    n49320, n49321, n49322, n49323, n49324, n49325,
    n49326, n49327, n49328, n49329, n49330, n49331,
    n49332, n49333, n49334, n49335, n49336, n49337,
    n49338, n49339, n49340, n49341, n49342, n49343,
    n49344, n49345, n49346, n49347, n49348, n49349,
    n49350, n49351, n49352, n49353, n49354, n49355,
    n49356, n49357, n49358, n49359, n49360, n49361,
    n49362, n49363, n49364, n49365, n49366, n49367,
    n49368, n49369, n49370, n49371, n49372, n49373,
    n49374, n49375, n49376, n49377, n49378, n49379,
    n49380, n49381, n49382, n49383, n49384, n49385,
    n49386, n49387, n49388, n49389, n49390, n49391,
    n49392, n49393, n49394, n49395, n49396, n49397,
    n49398, n49399, n49400, n49401, n49402, n49404,
    n49405, n49406, n49407, n49408, n49409, n49410,
    n49411, n49412, n49413, n49414, n49415, n49416,
    n49417, n49418, n49419, n49420, n49421, n49422,
    n49423, n49424, n49425, n49426, n49427, n49428,
    n49429, n49430, n49431, n49432, n49433, n49434,
    n49435, n49436, n49437, n49438, n49439, n49440,
    n49441, n49442, n49443, n49444, n49445, n49446,
    n49447, n49448, n49449, n49450, n49451, n49452,
    n49453, n49454, n49455, n49456, n49457, n49458,
    n49459, n49460, n49461, n49462, n49463, n49464,
    n49465, n49466, n49467, n49468, n49469, n49470,
    n49471, n49472, n49473, n49474, n49475, n49476,
    n49477, n49478, n49479, n49480, n49481, n49482,
    n49483, n49484, n49485, n49486, n49487, n49488,
    n49489, n49490, n49491, n49492, n49493, n49494,
    n49495, n49496, n49497, n49498, n49499, n49500,
    n49501, n49502, n49503, n49504, n49505, n49506,
    n49507, n49508, n49509, n49510, n49511, n49512,
    n49513, n49514, n49515, n49516, n49517, n49518,
    n49519, n49520, n49521, n49522, n49523, n49524,
    n49525, n49526, n49527, n49528, n49529, n49530,
    n49531, n49532, n49533, n49534, n49535, n49536,
    n49537, n49538, n49539, n49540, n49541, n49542,
    n49543, n49544, n49545, n49546, n49547, n49548,
    n49549, n49550, n49551, n49552, n49553, n49554,
    n49555, n49556, n49557, n49558, n49559, n49560,
    n49561, n49562, n49563, n49564, n49565, n49566,
    n49567, n49568, n49569, n49570, n49571, n49572,
    n49573, n49574, n49575, n49576, n49577, n49578,
    n49579, n49580, n49581, n49582, n49583, n49584,
    n49585, n49586, n49587, n49588, n49589, n49590,
    n49591, n49592, n49593, n49594, n49595, n49596,
    n49597, n49598, n49599, n49600, n49601, n49602,
    n49603, n49604, n49605, n49606, n49607, n49608,
    n49609, n49610, n49611, n49612, n49613, n49614,
    n49615, n49616, n49617, n49618, n49619, n49620,
    n49621, n49622, n49623, n49624, n49625, n49626,
    n49627, n49628, n49629, n49630, n49631, n49632,
    n49633, n49634, n49635, n49636, n49637, n49638,
    n49639, n49640, n49641, n49642, n49643, n49644,
    n49645, n49646, n49647, n49648, n49649, n49650,
    n49651, n49652, n49653, n49654, n49655, n49656,
    n49657, n49658, n49659, n49660, n49661, n49662,
    n49663, n49664, n49665, n49666, n49667, n49668,
    n49669, n49670, n49671, n49672, n49673, n49674,
    n49675, n49676, n49677, n49678, n49679, n49680,
    n49681, n49682, n49683, n49684, n49685, n49686,
    n49687, n49688, n49689, n49690, n49691, n49692,
    n49693, n49694, n49695, n49696, n49697, n49698,
    n49699, n49700, n49701, n49702, n49703, n49704,
    n49705, n49706, n49707, n49708, n49709, n49710,
    n49711, n49712, n49713, n49714, n49715, n49716,
    n49717, n49718, n49720, n49721, n49722, n49723,
    n49724, n49725, n49726, n49727, n49728, n49729,
    n49730, n49731, n49732, n49733, n49734, n49735,
    n49736, n49737, n49738, n49739, n49740, n49741,
    n49742, n49743, n49744, n49745, n49746, n49747,
    n49748, n49749, n49750, n49751, n49752, n49753,
    n49754, n49755, n49756, n49757, n49758, n49759,
    n49760, n49761, n49762, n49763, n49764, n49765,
    n49766, n49767, n49768, n49769, n49770, n49771,
    n49772, n49773, n49774, n49775, n49776, n49777,
    n49778, n49779, n49780, n49781, n49782, n49783,
    n49784, n49785, n49786, n49787, n49788, n49789,
    n49790, n49791, n49792, n49793, n49794, n49795,
    n49796, n49797, n49798, n49799, n49800, n49801,
    n49802, n49803, n49804, n49805, n49806, n49807,
    n49808, n49809, n49810, n49811, n49812, n49813,
    n49814, n49815, n49816, n49817, n49818, n49819,
    n49820, n49821, n49822, n49823, n49824, n49825,
    n49826, n49827, n49828, n49829, n49830, n49831,
    n49832, n49833, n49834, n49835, n49836, n49837,
    n49838, n49839, n49840, n49841, n49842, n49843,
    n49844, n49845, n49846, n49847, n49848, n49849,
    n49850, n49851, n49852, n49853, n49854, n49855,
    n49856, n49857, n49858, n49859, n49860, n49861,
    n49862, n49863, n49864, n49865, n49866, n49867,
    n49868, n49869, n49870, n49871, n49872, n49873,
    n49874, n49875, n49876, n49877, n49878, n49879,
    n49880, n49881, n49882, n49883, n49884, n49885,
    n49886, n49887, n49888, n49889, n49890, n49891,
    n49892, n49893, n49894, n49895, n49896, n49897,
    n49898, n49899, n49900, n49901, n49902, n49903,
    n49904, n49905, n49906, n49907, n49908, n49909,
    n49910, n49911, n49912, n49913, n49914, n49915,
    n49916, n49917, n49918, n49919, n49920, n49921,
    n49922, n49923, n49924, n49925, n49926, n49927,
    n49928, n49929, n49930, n49931, n49932, n49933,
    n49934, n49935, n49936, n49937, n49938, n49939,
    n49940, n49941, n49942, n49943, n49944, n49945,
    n49946, n49947, n49948, n49949, n49950, n49951,
    n49952, n49953, n49954, n49955, n49956, n49957,
    n49958, n49959, n49960, n49961, n49962, n49963,
    n49964, n49965, n49966, n49967, n49968, n49969,
    n49970, n49971, n49972, n49973, n49974, n49975,
    n49976, n49977, n49978, n49979, n49980, n49981,
    n49982, n49983, n49984, n49985, n49986, n49987,
    n49988, n49989, n49990, n49991, n49992, n49993,
    n49994, n49995, n49996, n49997, n49998, n49999,
    n50000, n50001, n50002, n50003, n50004, n50005,
    n50006, n50007, n50008, n50009, n50010, n50011,
    n50012, n50013, n50014, n50015, n50016, n50017,
    n50018, n50019, n50020, n50021, n50022, n50023,
    n50024, n50025, n50026, n50027, n50028, n50029,
    n50030, n50031, n50032, n50033, n50034, n50035,
    n50036, n50037, n50038, n50039, n50040, n50041,
    n50042, n50043, n50044, n50045, n50046, n50047,
    n50048, n50049, n50050, n50051, n50052, n50053,
    n50054, n50055, n50056, n50057, n50059, n50060,
    n50061, n50062, n50063, n50064, n50065, n50066,
    n50067, n50068, n50069, n50070, n50071, n50072,
    n50073, n50074, n50075, n50076, n50077, n50078,
    n50079, n50080, n50081, n50082, n50083, n50084,
    n50085, n50086, n50087, n50088, n50089, n50090,
    n50091, n50092, n50093, n50094, n50095, n50096,
    n50097, n50098, n50099, n50100, n50101, n50102,
    n50103, n50104, n50105, n50106, n50107, n50108,
    n50109, n50110, n50111, n50112, n50113, n50114,
    n50115, n50116, n50117, n50118, n50119, n50120,
    n50121, n50122, n50123, n50124, n50125, n50126,
    n50127, n50128, n50129, n50130, n50131, n50132,
    n50133, n50134, n50135, n50136, n50137, n50138,
    n50139, n50140, n50141, n50142, n50143, n50144,
    n50145, n50146, n50147, n50148, n50149, n50150,
    n50151, n50152, n50153, n50154, n50155, n50156,
    n50157, n50158, n50159, n50160, n50161, n50162,
    n50163, n50164, n50165, n50166, n50167, n50168,
    n50169, n50170, n50171, n50172, n50173, n50174,
    n50175, n50176, n50177, n50178, n50179, n50180,
    n50181, n50182, n50183, n50184, n50185, n50186,
    n50187, n50188, n50189, n50190, n50191, n50192,
    n50193, n50194, n50195, n50196, n50197, n50198,
    n50199, n50200, n50201, n50202, n50203, n50204,
    n50205, n50206, n50207, n50208, n50209, n50210,
    n50211, n50212, n50213, n50214, n50215, n50216,
    n50217, n50218, n50219, n50220, n50221, n50222,
    n50223, n50224, n50225, n50226, n50227, n50228,
    n50229, n50230, n50231, n50232, n50233, n50234,
    n50235, n50236, n50237, n50238, n50239, n50240,
    n50241, n50242, n50243, n50244, n50245, n50246,
    n50247, n50248, n50249, n50250, n50251, n50252,
    n50253, n50254, n50255, n50256, n50257, n50258,
    n50259, n50260, n50261, n50262, n50263, n50264,
    n50265, n50266, n50267, n50268, n50269, n50270,
    n50271, n50272, n50273, n50274, n50275, n50276,
    n50277, n50278, n50279, n50280, n50281, n50282,
    n50283, n50284, n50285, n50286, n50287, n50288,
    n50289, n50290, n50291, n50292, n50293, n50294,
    n50295, n50296, n50297, n50298, n50299, n50300,
    n50301, n50302, n50303, n50304, n50305, n50306,
    n50307, n50308, n50309, n50310, n50311, n50313,
    n50314, n50315, n50316, n50317, n50318, n50319,
    n50320, n50321, n50322, n50323, n50324, n50325,
    n50326, n50327, n50328, n50329, n50330, n50331,
    n50332, n50333, n50334, n50335, n50336, n50337,
    n50338, n50339, n50340, n50341, n50342, n50343,
    n50344, n50345, n50346, n50347, n50348, n50349,
    n50350, n50351, n50352, n50353, n50354, n50355,
    n50356, n50357, n50358, n50359, n50360, n50361,
    n50362, n50363, n50364, n50365, n50366, n50367,
    n50368, n50369, n50370, n50371, n50372, n50373,
    n50374, n50375, n50376, n50377, n50378, n50379,
    n50380, n50381, n50382, n50383, n50384, n50385,
    n50386, n50387, n50388, n50389, n50390, n50391,
    n50392, n50393, n50394, n50395, n50396, n50397,
    n50398, n50399, n50400, n50401, n50402, n50403,
    n50404, n50405, n50406, n50407, n50408, n50409,
    n50410, n50411, n50412, n50413, n50414, n50415,
    n50416, n50417, n50418, n50419, n50420, n50421,
    n50422, n50423, n50424, n50425, n50426, n50427,
    n50428, n50429, n50430, n50431, n50432, n50433,
    n50434, n50435, n50436, n50437, n50438, n50439,
    n50440, n50441, n50442, n50443, n50444, n50445,
    n50446, n50447, n50448, n50449, n50450, n50451,
    n50452, n50453, n50454, n50455, n50456, n50457,
    n50458, n50459, n50460, n50461, n50462, n50463,
    n50464, n50465, n50466, n50467, n50468, n50469,
    n50470, n50471, n50472, n50473, n50474, n50475,
    n50476, n50477, n50478, n50479, n50480, n50481,
    n50482, n50483, n50484, n50485, n50486, n50487,
    n50488, n50489, n50490, n50491, n50492, n50493,
    n50494, n50495, n50496, n50497, n50498, n50499,
    n50500, n50501, n50502, n50503, n50504, n50505,
    n50506, n50507, n50508, n50509, n50510, n50511,
    n50512, n50513, n50514, n50515, n50516, n50517,
    n50518, n50519, n50520, n50521, n50522, n50523,
    n50524, n50525, n50526, n50527, n50528, n50529,
    n50530, n50531, n50532, n50533, n50534, n50535,
    n50536, n50537, n50538, n50539, n50540, n50541,
    n50542, n50543, n50545, n50546, n50547, n50548,
    n50549, n50550, n50551, n50552, n50553, n50554,
    n50555, n50556, n50557, n50558, n50559, n50560,
    n50561, n50562, n50563, n50564, n50565, n50566,
    n50567, n50568, n50569, n50570, n50571, n50572,
    n50573, n50574, n50575, n50576, n50577, n50578,
    n50579, n50580, n50581, n50582, n50583, n50584,
    n50585, n50586, n50587, n50588, n50589, n50590,
    n50591, n50592, n50593, n50594, n50595, n50596,
    n50597, n50598, n50599, n50600, n50601, n50602,
    n50603, n50604, n50605, n50606, n50607, n50608,
    n50609, n50610, n50611, n50612, n50613, n50614,
    n50615, n50616, n50617, n50618, n50619, n50620,
    n50621, n50622, n50623, n50624, n50625, n50626,
    n50627, n50628, n50629, n50630, n50631, n50632,
    n50633, n50634, n50635, n50636, n50637, n50638,
    n50639, n50640, n50641, n50642, n50643, n50644,
    n50645, n50646, n50647, n50648, n50649, n50650,
    n50651, n50652, n50653, n50654, n50655, n50656,
    n50657, n50658, n50659, n50660, n50661, n50662,
    n50663, n50664, n50665, n50666, n50667, n50668,
    n50669, n50670, n50671, n50672, n50673, n50674,
    n50675, n50676, n50677, n50678, n50679, n50680,
    n50681, n50682, n50683, n50684, n50685, n50686,
    n50687, n50688, n50689, n50690, n50691, n50692,
    n50693, n50694, n50695, n50696, n50697, n50698,
    n50699, n50700, n50701, n50702, n50703, n50704,
    n50705, n50706, n50707, n50708, n50709, n50710,
    n50711, n50712, n50713, n50714, n50715, n50716,
    n50717, n50718, n50719, n50720, n50721, n50722,
    n50723, n50724, n50725, n50726, n50727, n50728,
    n50729, n50730, n50731, n50732, n50733, n50734,
    n50735, n50736, n50737, n50738, n50739, n50740,
    n50741, n50742, n50743, n50744, n50745, n50746,
    n50747, n50748, n50749, n50750, n50751, n50752,
    n50753, n50754, n50755, n50756, n50757, n50758,
    n50759, n50760, n50761, n50762, n50763, n50764,
    n50765, n50766, n50767, n50768, n50769, n50770,
    n50771, n50772, n50773, n50774, n50775, n50776,
    n50777, n50778, n50779, n50780, n50781, n50782,
    n50783, n50784, n50785, n50786, n50787, n50788,
    n50789, n50790, n50792, n50793, n50794, n50795,
    n50796, n50797, n50798, n50799, n50800, n50801,
    n50802, n50803, n50804, n50805, n50806, n50807,
    n50808, n50809, n50810, n50811, n50812, n50813,
    n50814, n50815, n50816, n50817, n50818, n50819,
    n50820, n50821, n50822, n50823, n50824, n50825,
    n50826, n50827, n50828, n50829, n50830, n50831,
    n50832, n50833, n50834, n50835, n50836, n50837,
    n50838, n50839, n50840, n50841, n50842, n50843,
    n50844, n50845, n50846, n50847, n50848, n50849,
    n50850, n50851, n50852, n50853, n50854, n50855,
    n50856, n50857, n50858, n50859, n50860, n50861,
    n50862, n50863, n50864, n50865, n50866, n50867,
    n50868, n50869, n50870, n50871, n50872, n50873,
    n50874, n50875, n50876, n50877, n50878, n50879,
    n50880, n50881, n50882, n50883, n50884, n50885,
    n50886, n50887, n50888, n50889, n50890, n50891,
    n50892, n50893, n50894, n50895, n50896, n50897,
    n50898, n50899, n50900, n50901, n50902, n50903,
    n50904, n50905, n50906, n50907, n50908, n50909,
    n50910, n50911, n50912, n50913, n50914, n50915,
    n50916, n50917, n50918, n50919, n50920, n50921,
    n50922, n50923, n50924, n50925, n50926, n50927,
    n50928, n50929, n50930, n50931, n50932, n50933,
    n50934, n50935, n50936, n50937, n50938, n50939,
    n50940, n50941, n50942, n50943, n50944, n50945,
    n50946, n50947, n50948, n50949, n50950, n50951,
    n50952, n50953, n50954, n50955, n50956, n50957,
    n50958, n50959, n50960, n50961, n50962, n50963,
    n50964, n50965, n50966, n50967, n50968, n50969,
    n50970, n50971, n50972, n50973, n50974, n50975,
    n50976, n50977, n50978, n50979, n50980, n50981,
    n50982, n50983, n50984, n50985, n50986, n50987,
    n50988, n50989, n50990, n50991, n50992, n50993,
    n50994, n50995, n50996, n50997, n50998, n50999,
    n51000, n51001, n51002, n51003, n51004, n51005,
    n51006, n51007, n51008, n51009, n51010, n51011,
    n51012, n51013, n51014, n51015, n51016, n51017,
    n51018, n51019, n51020, n51021, n51022, n51023,
    n51024, n51025, n51026, n51027, n51028, n51029,
    n51030, n51031, n51032, n51033, n51034, n51035,
    n51036, n51037, n51039, n51040, n51041, n51042,
    n51043, n51044, n51045, n51046, n51047, n51048,
    n51049, n51050, n51051, n51052, n51053, n51054,
    n51055, n51056, n51057, n51058, n51059, n51060,
    n51061, n51062, n51063, n51064, n51065, n51066,
    n51067, n51068, n51069, n51070, n51071, n51072,
    n51073, n51074, n51075, n51076, n51077, n51078,
    n51079, n51080, n51081, n51082, n51083, n51084,
    n51085, n51086, n51087, n51088, n51089, n51090,
    n51091, n51092, n51093, n51094, n51095, n51096,
    n51097, n51098, n51099, n51100, n51101, n51102,
    n51103, n51104, n51105, n51106, n51107, n51108,
    n51109, n51110, n51111, n51112, n51113, n51114,
    n51115, n51116, n51117, n51118, n51119, n51120,
    n51121, n51122, n51123, n51124, n51125, n51126,
    n51127, n51128, n51129, n51130, n51131, n51132,
    n51133, n51134, n51135, n51136, n51137, n51138,
    n51139, n51140, n51141, n51142, n51143, n51144,
    n51145, n51146, n51147, n51148, n51149, n51150,
    n51151, n51152, n51153, n51154, n51155, n51156,
    n51157, n51158, n51159, n51160, n51161, n51162,
    n51163, n51164, n51165, n51166, n51167, n51168,
    n51169, n51170, n51171, n51172, n51173, n51174,
    n51175, n51176, n51177, n51178, n51179, n51180,
    n51181, n51182, n51183, n51184, n51185, n51186,
    n51187, n51188, n51189, n51190, n51191, n51192,
    n51193, n51194, n51195, n51196, n51197, n51198,
    n51199, n51200, n51201, n51202, n51203, n51204,
    n51205, n51206, n51207, n51208, n51209, n51210,
    n51211, n51212, n51213, n51214, n51215, n51216,
    n51217, n51218, n51219, n51220, n51221, n51222,
    n51223, n51224, n51225, n51226, n51227, n51228,
    n51229, n51230, n51231, n51232, n51233, n51234,
    n51235, n51236, n51237, n51238, n51239, n51240,
    n51241, n51242, n51243, n51244, n51245, n51246,
    n51247, n51248, n51249, n51250, n51252, n51253,
    n51254, n51255, n51256, n51257, n51258, n51259,
    n51260, n51261, n51262, n51263, n51264, n51265,
    n51266, n51267, n51268, n51269, n51270, n51271,
    n51272, n51273, n51274, n51275, n51276, n51277,
    n51278, n51279, n51280, n51281, n51282, n51283,
    n51284, n51285, n51286, n51287, n51288, n51289,
    n51290, n51291, n51292, n51293, n51294, n51295,
    n51296, n51297, n51298, n51299, n51300, n51301,
    n51302, n51303, n51304, n51305, n51306, n51307,
    n51308, n51309, n51310, n51311, n51312, n51313,
    n51314, n51315, n51316, n51317, n51318, n51319,
    n51320, n51321, n51322, n51323, n51324, n51325,
    n51326, n51327, n51328, n51329, n51330, n51331,
    n51332, n51333, n51334, n51335, n51336, n51337,
    n51338, n51339, n51340, n51341, n51342, n51343,
    n51344, n51345, n51346, n51347, n51348, n51349,
    n51350, n51351, n51352, n51353, n51354, n51355,
    n51356, n51357, n51358, n51359, n51360, n51361,
    n51362, n51363, n51364, n51365, n51366, n51367,
    n51368, n51369, n51370, n51371, n51372, n51373,
    n51374, n51375, n51376, n51377, n51378, n51379,
    n51380, n51381, n51382, n51383, n51384, n51385,
    n51386, n51387, n51388, n51389, n51390, n51391,
    n51392, n51393, n51394, n51395, n51396, n51397,
    n51398, n51399, n51400, n51401, n51402, n51403,
    n51404, n51405, n51406, n51407, n51408, n51409,
    n51410, n51411, n51412, n51413, n51414, n51415,
    n51416, n51417, n51418, n51419, n51420, n51421,
    n51422, n51423, n51424, n51425, n51426, n51427,
    n51428, n51429, n51430, n51431, n51432, n51433,
    n51434, n51435, n51436, n51437, n51438, n51439,
    n51440, n51441, n51442, n51443, n51444, n51445,
    n51446, n51447, n51448, n51449, n51450, n51451,
    n51452, n51453, n51454, n51455, n51456, n51457,
    n51458, n51459, n51460, n51461, n51462, n51463,
    n51464, n51465, n51466, n51467, n51468, n51469,
    n51470, n51471, n51472, n51473, n51474, n51475,
    n51476, n51478, n51479, n51480, n51481, n51482,
    n51483, n51484, n51485, n51486, n51487, n51488,
    n51489, n51490, n51491, n51492, n51493, n51494,
    n51495, n51496, n51497, n51498, n51499, n51500,
    n51501, n51502, n51503, n51504, n51505, n51506,
    n51507, n51508, n51509, n51510, n51511, n51512,
    n51513, n51514, n51515, n51516, n51517, n51518,
    n51519, n51520, n51521, n51522, n51523, n51524,
    n51525, n51526, n51527, n51528, n51529, n51530,
    n51531, n51532, n51533, n51534, n51535, n51536,
    n51537, n51538, n51539, n51540, n51541, n51542,
    n51543, n51544, n51545, n51546, n51547, n51548,
    n51549, n51550, n51551, n51552, n51553, n51554,
    n51555, n51556, n51557, n51558, n51559, n51560,
    n51561, n51562, n51563, n51564, n51565, n51566,
    n51567, n51568, n51569, n51570, n51571, n51572,
    n51573, n51574, n51575, n51576, n51577, n51578,
    n51579, n51580, n51581, n51582, n51583, n51584,
    n51585, n51586, n51587, n51588, n51589, n51590,
    n51591, n51592, n51593, n51594, n51595, n51596,
    n51597, n51598, n51599, n51600, n51601, n51602,
    n51603, n51604, n51605, n51606, n51607, n51608,
    n51609, n51610, n51611, n51612, n51613, n51614,
    n51615, n51616, n51617, n51618, n51619, n51620,
    n51621, n51622, n51623, n51624, n51625, n51626,
    n51627, n51628, n51629, n51630, n51631, n51632,
    n51633, n51634, n51635, n51636, n51637, n51638,
    n51639, n51640, n51641, n51642, n51643, n51644,
    n51645, n51646, n51647, n51648, n51649, n51650,
    n51651, n51652, n51653, n51654, n51655, n51656,
    n51657, n51658, n51659, n51660, n51661, n51662,
    n51663, n51665, n51666, n51667, n51668, n51669,
    n51670, n51671, n51672, n51673, n51674, n51675,
    n51676, n51677, n51678, n51679, n51680, n51681,
    n51682, n51683, n51684, n51685, n51686, n51687,
    n51688, n51689, n51690, n51691, n51692, n51693,
    n51694, n51695, n51696, n51697, n51698, n51699,
    n51700, n51701, n51702, n51703, n51704, n51705,
    n51706, n51707, n51708, n51709, n51710, n51711,
    n51712, n51713, n51714, n51715, n51716, n51717,
    n51718, n51719, n51720, n51721, n51722, n51723,
    n51724, n51725, n51726, n51727, n51728, n51729,
    n51730, n51731, n51732, n51733, n51734, n51735,
    n51736, n51737, n51738, n51739, n51740, n51741,
    n51742, n51743, n51744, n51745, n51746, n51747,
    n51748, n51749, n51750, n51751, n51752, n51753,
    n51754, n51755, n51756, n51757, n51758, n51759,
    n51760, n51761, n51762, n51763, n51764, n51765,
    n51766, n51767, n51768, n51769, n51770, n51771,
    n51772, n51773, n51774, n51775, n51776, n51777,
    n51778, n51779, n51780, n51781, n51782, n51783,
    n51784, n51785, n51786, n51787, n51788, n51789,
    n51790, n51791, n51792, n51793, n51794, n51795,
    n51796, n51797, n51798, n51799, n51800, n51801,
    n51802, n51803, n51804, n51805, n51806, n51807,
    n51808, n51809, n51810, n51811, n51812, n51813,
    n51814, n51815, n51816, n51817, n51818, n51819,
    n51820, n51821, n51822, n51823, n51824, n51825,
    n51826, n51827, n51828, n51829, n51830, n51831,
    n51832, n51833, n51834, n51835, n51836, n51837,
    n51838, n51839, n51840, n51841, n51842, n51843,
    n51844, n51845, n51846, n51847, n51848, n51849,
    n51850, n51851, n51852, n51853, n51854, n51855,
    n51857, n51858, n51859, n51860, n51861, n51862,
    n51863, n51864, n51865, n51866, n51867, n51868,
    n51869, n51870, n51871, n51872, n51873, n51874,
    n51875, n51876, n51877, n51878, n51879, n51880,
    n51881, n51882, n51883, n51884, n51885, n51886,
    n51887, n51888, n51889, n51890, n51891, n51892,
    n51893, n51894, n51895, n51896, n51897, n51898,
    n51899, n51900, n51901, n51902, n51903, n51904,
    n51905, n51906, n51907, n51908, n51909, n51910,
    n51911, n51912, n51913, n51914, n51915, n51916,
    n51917, n51918, n51919, n51920, n51921, n51922,
    n51923, n51924, n51925, n51926, n51927, n51928,
    n51929, n51930, n51931, n51932, n51933, n51934,
    n51935, n51936, n51937, n51938, n51939, n51940,
    n51941, n51942, n51943, n51944, n51945, n51946,
    n51947, n51948, n51949, n51950, n51951, n51952,
    n51953, n51954, n51955, n51956, n51957, n51958,
    n51959, n51960, n51961, n51962, n51963, n51964,
    n51965, n51966, n51967, n51968, n51969, n51970,
    n51971, n51972, n51973, n51974, n51975, n51976,
    n51977, n51978, n51979, n51980, n51981, n51982,
    n51983, n51984, n51985, n51986, n51987, n51988,
    n51989, n51990, n51991, n51992, n51993, n51994,
    n51995, n51996, n51997, n51998, n51999, n52000,
    n52001, n52002, n52003, n52004, n52005, n52006,
    n52007, n52008, n52009, n52010, n52011, n52012,
    n52013, n52014, n52015, n52016, n52017, n52018,
    n52019, n52020, n52021, n52022, n52023, n52024,
    n52025, n52026, n52027, n52028, n52029, n52030,
    n52031, n52032, n52033, n52034, n52035, n52036,
    n52037, n52038, n52039, n52040, n52041, n52042,
    n52043, n52044, n52046, n52047, n52048, n52049,
    n52050, n52051, n52052, n52053, n52054, n52055,
    n52056, n52057, n52058, n52059, n52060, n52061,
    n52062, n52063, n52064, n52065, n52066, n52067,
    n52068, n52069, n52070, n52071, n52072, n52073,
    n52074, n52075, n52076, n52077, n52078, n52079,
    n52080, n52081, n52082, n52083, n52084, n52085,
    n52086, n52087, n52088, n52089, n52090, n52091,
    n52092, n52093, n52094, n52095, n52096, n52097,
    n52098, n52099, n52100, n52101, n52102, n52103,
    n52104, n52105, n52106, n52107, n52108, n52109,
    n52110, n52111, n52112, n52113, n52114, n52115,
    n52116, n52117, n52118, n52119, n52120, n52121,
    n52122, n52123, n52124, n52125, n52126, n52127,
    n52128, n52129, n52130, n52131, n52132, n52133,
    n52134, n52135, n52136, n52137, n52138, n52139,
    n52140, n52141, n52142, n52143, n52144, n52145,
    n52146, n52147, n52148, n52149, n52150, n52151,
    n52152, n52153, n52154, n52155, n52156, n52157,
    n52158, n52159, n52160, n52161, n52162, n52163,
    n52164, n52165, n52166, n52167, n52168, n52169,
    n52170, n52171, n52172, n52173, n52174, n52175,
    n52176, n52177, n52178, n52179, n52180, n52181,
    n52182, n52183, n52184, n52185, n52186, n52187,
    n52188, n52189, n52190, n52191, n52192, n52193,
    n52194, n52195, n52196, n52197, n52198, n52199,
    n52200, n52201, n52202, n52203, n52204, n52205,
    n52206, n52207, n52208, n52209, n52210, n52211,
    n52212, n52213, n52214, n52215, n52216, n52217,
    n52218, n52219, n52220, n52222, n52223, n52224,
    n52225, n52226, n52227, n52228, n52229, n52230,
    n52231, n52232, n52233, n52234, n52235, n52236,
    n52237, n52238, n52239, n52240, n52241, n52242,
    n52243, n52244, n52245, n52246, n52247, n52248,
    n52249, n52250, n52251, n52252, n52253, n52254,
    n52255, n52256, n52257, n52258, n52259, n52260,
    n52261, n52262, n52263, n52264, n52265, n52266,
    n52267, n52268, n52269, n52270, n52271, n52272,
    n52273, n52274, n52275, n52276, n52277, n52278,
    n52279, n52280, n52281, n52282, n52283, n52284,
    n52285, n52286, n52287, n52288, n52289, n52290,
    n52291, n52292, n52293, n52294, n52295, n52296,
    n52297, n52298, n52299, n52300, n52301, n52302,
    n52303, n52304, n52305, n52306, n52307, n52308,
    n52309, n52310, n52311, n52312, n52313, n52314,
    n52315, n52316, n52317, n52318, n52319, n52320,
    n52321, n52322, n52323, n52324, n52325, n52326,
    n52327, n52328, n52329, n52330, n52331, n52332,
    n52333, n52334, n52335, n52336, n52337, n52338,
    n52339, n52340, n52341, n52342, n52343, n52344,
    n52345, n52346, n52347, n52348, n52349, n52350,
    n52351, n52352, n52353, n52354, n52355, n52356,
    n52357, n52358, n52359, n52360, n52361, n52362,
    n52363, n52364, n52365, n52366, n52367, n52368,
    n52369, n52370, n52371, n52372, n52373, n52374,
    n52375, n52376, n52377, n52378, n52379, n52380,
    n52381, n52382, n52384, n52385, n52386, n52387,
    n52388, n52389, n52390, n52391, n52392, n52393,
    n52394, n52395, n52396, n52397, n52398, n52399,
    n52400, n52401, n52402, n52403, n52404, n52405,
    n52406, n52407, n52408, n52409, n52410, n52411,
    n52412, n52413, n52414, n52415, n52416, n52417,
    n52418, n52419, n52420, n52421, n52422, n52423,
    n52424, n52425, n52426, n52427, n52428, n52429,
    n52430, n52431, n52432, n52433, n52434, n52435,
    n52436, n52437, n52438, n52439, n52440, n52441,
    n52442, n52443, n52444, n52445, n52446, n52447,
    n52448, n52449, n52450, n52451, n52452, n52453,
    n52454, n52455, n52456, n52457, n52458, n52459,
    n52460, n52461, n52462, n52463, n52464, n52465,
    n52466, n52467, n52468, n52469, n52470, n52471,
    n52472, n52473, n52474, n52475, n52476, n52477,
    n52478, n52479, n52480, n52481, n52482, n52483,
    n52484, n52485, n52486, n52487, n52488, n52489,
    n52490, n52491, n52492, n52493, n52494, n52495,
    n52496, n52497, n52498, n52499, n52500, n52501,
    n52502, n52503, n52504, n52505, n52506, n52507,
    n52508, n52509, n52510, n52511, n52512, n52513,
    n52514, n52515, n52516, n52517, n52518, n52519,
    n52520, n52521, n52522, n52523, n52524, n52525,
    n52526, n52527, n52528, n52529, n52530, n52531,
    n52533, n52534, n52535, n52536, n52537, n52538,
    n52539, n52540, n52541, n52542, n52543, n52544,
    n52545, n52546, n52547, n52548, n52549, n52550,
    n52551, n52552, n52553, n52554, n52555, n52556,
    n52557, n52558, n52559, n52560, n52561, n52562,
    n52563, n52564, n52565, n52566, n52567, n52568,
    n52569, n52570, n52571, n52572, n52573, n52574,
    n52575, n52576, n52577, n52578, n52579, n52580,
    n52581, n52582, n52583, n52584, n52585, n52586,
    n52587, n52588, n52589, n52590, n52591, n52592,
    n52593, n52594, n52595, n52596, n52597, n52598,
    n52599, n52600, n52601, n52602, n52603, n52604,
    n52605, n52606, n52607, n52608, n52609, n52610,
    n52611, n52612, n52613, n52614, n52615, n52616,
    n52617, n52618, n52619, n52620, n52621, n52622,
    n52623, n52624, n52625, n52626, n52627, n52628,
    n52629, n52630, n52631, n52632, n52633, n52634,
    n52635, n52636, n52637, n52638, n52639, n52640,
    n52641, n52642, n52643, n52644, n52645, n52646,
    n52647, n52648, n52649, n52650, n52651, n52652,
    n52653, n52654, n52655, n52656, n52657, n52658,
    n52659, n52660, n52661, n52662, n52663, n52664,
    n52665, n52666, n52667, n52668, n52669, n52670,
    n52671, n52672, n52673, n52674, n52675, n52676,
    n52677, n52678, n52679, n52680, n52681, n52682,
    n52683, n52684, n52685, n52686, n52687, n52688,
    n52689, n52690, n52692, n52693, n52694, n52695,
    n52696, n52697, n52698, n52699, n52700, n52701,
    n52702, n52703, n52704, n52705, n52706, n52707,
    n52708, n52709, n52710, n52711, n52712, n52713,
    n52714, n52715, n52716, n52717, n52718, n52719,
    n52720, n52721, n52722, n52723, n52724, n52725,
    n52726, n52727, n52728, n52729, n52730, n52731,
    n52732, n52733, n52734, n52735, n52736, n52737,
    n52738, n52739, n52740, n52741, n52742, n52743,
    n52744, n52745, n52746, n52747, n52748, n52749,
    n52750, n52751, n52752, n52753, n52754, n52755,
    n52756, n52757, n52758, n52759, n52760, n52761,
    n52762, n52763, n52764, n52765, n52766, n52767,
    n52768, n52769, n52770, n52771, n52772, n52773,
    n52774, n52775, n52776, n52777, n52778, n52779,
    n52780, n52781, n52782, n52783, n52784, n52785,
    n52786, n52787, n52788, n52789, n52790, n52791,
    n52792, n52793, n52794, n52795, n52796, n52797,
    n52798, n52799, n52800, n52801, n52802, n52803,
    n52804, n52805, n52806, n52807, n52808, n52809,
    n52810, n52811, n52812, n52813, n52814, n52815,
    n52816, n52817, n52818, n52819, n52820, n52821,
    n52822, n52823, n52824, n52825, n52826, n52828,
    n52829, n52830, n52831, n52832, n52833, n52834,
    n52835, n52836, n52837, n52838, n52839, n52840,
    n52841, n52842, n52843, n52844, n52845, n52846,
    n52847, n52848, n52849, n52850, n52851, n52852,
    n52853, n52854, n52855, n52856, n52857, n52858,
    n52859, n52860, n52861, n52862, n52863, n52864,
    n52865, n52866, n52867, n52868, n52869, n52870,
    n52871, n52872, n52873, n52874, n52875, n52876,
    n52877, n52878, n52879, n52880, n52881, n52882,
    n52883, n52884, n52885, n52886, n52887, n52888,
    n52889, n52890, n52891, n52892, n52893, n52894,
    n52895, n52896, n52897, n52898, n52899, n52900,
    n52901, n52902, n52903, n52904, n52905, n52906,
    n52907, n52908, n52909, n52910, n52911, n52912,
    n52913, n52914, n52915, n52916, n52917, n52918,
    n52919, n52920, n52921, n52922, n52923, n52924,
    n52925, n52926, n52927, n52928, n52929, n52930,
    n52931, n52932, n52933, n52934, n52935, n52936,
    n52937, n52938, n52939, n52940, n52941, n52942,
    n52943, n52944, n52945, n52946, n52947, n52948,
    n52949, n52950, n52951, n52952, n52953, n52954,
    n52955, n52956, n52957, n52958, n52959, n52960,
    n52961, n52962, n52963, n52964, n52965, n52966,
    n52967, n52968, n52969, n52970, n52971, n52972,
    n52973, n52974, n52976, n52977, n52978, n52979,
    n52980, n52981, n52982, n52983, n52984, n52985,
    n52986, n52987, n52988, n52989, n52990, n52991,
    n52992, n52993, n52994, n52995, n52996, n52997,
    n52998, n52999, n53000, n53001, n53002, n53003,
    n53004, n53005, n53006, n53007, n53008, n53009,
    n53010, n53011, n53012, n53013, n53014, n53015,
    n53016, n53017, n53018, n53019, n53020, n53021,
    n53022, n53023, n53024, n53025, n53026, n53027,
    n53028, n53029, n53030, n53031, n53032, n53033,
    n53034, n53035, n53036, n53037, n53038, n53039,
    n53040, n53041, n53042, n53043, n53044, n53045,
    n53046, n53047, n53048, n53049, n53050, n53051,
    n53052, n53053, n53054, n53055, n53056, n53057,
    n53058, n53059, n53060, n53061, n53062, n53063,
    n53064, n53065, n53066, n53067, n53068, n53069,
    n53070, n53071, n53072, n53073, n53074, n53075,
    n53076, n53077, n53078, n53079, n53080, n53081,
    n53082, n53083, n53084, n53085, n53086, n53087,
    n53088, n53089, n53090, n53091, n53092, n53093,
    n53094, n53095, n53096, n53097, n53098, n53099,
    n53100, n53101, n53102, n53103, n53104, n53105,
    n53106, n53107, n53108, n53109, n53110, n53112,
    n53113, n53114, n53115, n53116, n53117, n53118,
    n53119, n53120, n53121, n53122, n53123, n53124,
    n53125, n53126, n53127, n53128, n53129, n53130,
    n53131, n53132, n53133, n53134, n53135, n53136,
    n53137, n53138, n53139, n53140, n53141, n53142,
    n53143, n53144, n53145, n53146, n53147, n53148,
    n53149, n53150, n53151, n53152, n53153, n53154,
    n53155, n53156, n53157, n53158, n53159, n53160,
    n53161, n53162, n53163, n53164, n53165, n53166,
    n53167, n53168, n53169, n53170, n53171, n53172,
    n53173, n53174, n53175, n53176, n53177, n53178,
    n53179, n53180, n53181, n53182, n53183, n53184,
    n53185, n53186, n53187, n53188, n53189, n53190,
    n53191, n53192, n53193, n53194, n53195, n53196,
    n53197, n53198, n53199, n53200, n53201, n53202,
    n53203, n53204, n53205, n53206, n53207, n53208,
    n53209, n53210, n53211, n53212, n53213, n53214,
    n53215, n53216, n53217, n53218, n53219, n53220,
    n53221, n53222, n53223, n53224, n53225, n53226,
    n53227, n53228, n53229, n53230, n53231, n53232,
    n53233, n53234, n53236, n53237, n53238, n53239,
    n53240, n53241, n53242, n53243, n53244, n53245,
    n53246, n53247, n53248, n53249, n53250, n53251,
    n53252, n53253, n53254, n53255, n53256, n53257,
    n53258, n53259, n53260, n53261, n53262, n53263,
    n53264, n53265, n53266, n53267, n53268, n53269,
    n53270, n53271, n53272, n53273, n53274, n53275,
    n53276, n53277, n53278, n53279, n53280, n53281,
    n53282, n53283, n53284, n53285, n53286, n53287,
    n53288, n53289, n53290, n53291, n53292, n53293,
    n53294, n53295, n53296, n53297, n53298, n53299,
    n53300, n53301, n53302, n53303, n53304, n53305,
    n53306, n53307, n53308, n53309, n53310, n53311,
    n53312, n53313, n53314, n53315, n53316, n53317,
    n53318, n53319, n53320, n53321, n53322, n53323,
    n53324, n53325, n53326, n53327, n53328, n53329,
    n53330, n53331, n53333, n53334, n53335, n53336,
    n53337, n53338, n53339, n53340, n53341, n53342,
    n53343, n53344, n53345, n53346, n53347, n53348,
    n53349, n53350, n53351, n53352, n53353, n53354,
    n53355, n53356, n53357, n53358, n53359, n53360,
    n53361, n53362, n53363, n53364, n53365, n53366,
    n53367, n53368, n53369, n53370, n53371, n53372,
    n53373, n53374, n53375, n53376, n53377, n53378,
    n53379, n53380, n53381, n53382, n53383, n53384,
    n53385, n53386, n53387, n53388, n53389, n53390,
    n53391, n53392, n53393, n53394, n53395, n53396,
    n53397, n53398, n53399, n53400, n53401, n53402,
    n53403, n53404, n53405, n53406, n53407, n53408,
    n53409, n53410, n53411, n53412, n53413, n53414,
    n53415, n53416, n53417, n53418, n53419, n53420,
    n53421, n53422, n53423, n53424, n53425, n53426,
    n53427, n53428, n53429, n53430, n53431, n53432,
    n53433, n53434, n53435, n53436, n53437, n53438,
    n53439, n53440, n53441, n53442, n53443, n53444,
    n53445, n53446, n53447, n53448, n53449, n53450,
    n53451, n53452, n53453, n53454, n53455, n53456,
    n53457, n53458, n53459, n53460, n53461, n53462,
    n53463, n53464, n53465, n53466, n53467, n53468,
    n53469, n53470, n53471, n53472, n53473, n53474,
    n53475, n53476, n53477, n53478, n53479, n53480,
    n53481, n53482, n53483, n53484, n53485, n53486,
    n53487, n53488, n53489, n53490, n53491, n53492,
    n53493, n53494, n53495, n53496, n53497, n53498,
    n53499, n53500, n53501, n53502, n53503, n53504,
    n53505, n53506, n53507, n53508, n53509, n53510,
    n53511, n53512, n53513, n53514, n53515, n53516,
    n53517, n53518, n53519, n53520, n53521, n53522,
    n53523, n53524, n53525, n53526, n53527, n53528,
    n53529, n53530, n53531, n53532, n53533, n53534,
    n53535, n53536, n53537, n53538, n53539, n53540,
    n53541, n53542, n53543, n53544, n53545, n53546,
    n53547, n53548, n53549, n53550, n53551, n53552,
    n53553, n53554, n53555, n53556, n53557, n53558,
    n53559, n53560, n53561, n53562, n53563, n53564,
    n53565, n53566, n53567, n53568, n53569, n53570,
    n53571, n53572, n53573, n53574, n53575, n53576,
    n53577, n53578, n53579, n53580, n53581, n53582,
    n53583, n53584, n53585, n53586, n53587, n53588,
    n53589, n53590, n53591, n53592, n53593, n53594,
    n53595, n53596, n53597, n53598, n53599, n53600,
    n53601, n53602, n53603, n53604, n53605, n53606,
    n53607, n53608, n53609, n53610, n53611, n53612,
    n53613, n53614, n53615, n53616, n53617, n53618,
    n53619, n53620, n53621, n53622, n53623, n53624,
    n53625, n53626, n53627, n53628, n53629, n53630,
    n53631, n53632, n53633, n53634, n53635, n53636,
    n53637, n53638, n53639, n53640, n53641, n53642,
    n53643, n53644, n53645, n53646, n53647, n53648,
    n53649, n53650, n53651, n53652, n53653, n53654,
    n53655, n53656, n53657, n53658, n53659, n53660,
    n53661, n53662, n53663, n53664, n53665, n53666,
    n53667, n53668, n53669, n53670, n53671, n53672,
    n53673, n53674, n53675, n53676, n53677, n53678,
    n53679, n53680, n53681, n53682, n53683, n53684,
    n53685, n53686, n53687, n53688, n53689, n53690,
    n53691, n53692, n53693, n53694, n53695, n53696,
    n53697, n53698, n53699, n53700, n53701, n53702,
    n53703, n53704, n53705, n53706, n53707, n53708,
    n53709, n53710, n53711, n53712, n53713, n53714,
    n53715, n53716, n53717, n53718, n53719, n53720,
    n53721, n53722, n53723, n53724, n53725, n53726,
    n53727, n53728, n53729, n53730, n53731, n53732,
    n53733, n53734, n53735, n53736, n53737, n53738,
    n53739, n53740, n53741, n53742, n53743, n53744,
    n53745, n53746, n53747, n53748, n53749, n53750,
    n53751, n53752, n53753, n53754, n53755, n53756,
    n53757, n53758, n53759, n53760, n53761, n53762,
    n53763, n53764, n53765, n53766, n53767, n53768,
    n53769, n53770, n53771, n53772, n53773, n53774,
    n53775, n53776, n53777, n53778, n53779, n53780,
    n53781, n53782, n53783, n53784, n53785, n53786,
    n53787, n53788, n53789, n53790, n53791, n53792,
    n53793, n53794, n53795, n53796, n53797, n53798,
    n53799, n53800, n53801, n53802, n53803, n53804,
    n53805, n53806, n53807, n53808, n53809, n53810,
    n53811, n53812, n53813, n53814, n53815, n53816,
    n53817, n53818, n53819, n53820, n53821, n53822,
    n53823, n53824, n53825, n53826, n53827, n53828,
    n53829, n53830, n53831, n53832, n53833, n53834,
    n53835, n53836, n53837, n53838, n53839, n53840,
    n53841, n53842, n53843, n53844, n53845, n53846,
    n53847, n53848, n53849, n53850, n53851, n53852,
    n53853, n53854, n53855, n53856, n53857, n53858,
    n53859, n53860, n53861, n53862, n53863, n53864,
    n53865, n53866, n53867, n53868, n53869, n53870,
    n53871, n53872, n53873, n53874, n53875, n53876,
    n53877, n53878, n53879, n53880, n53881, n53882,
    n53883, n53884, n53885, n53886, n53887, n53888,
    n53889, n53890, n53891, n53892, n53893, n53894,
    n53895, n53896, n53897, n53898, n53899, n53900,
    n53901, n53902, n53903, n53904, n53905, n53906,
    n53907, n53908, n53909, n53910, n53911, n53912,
    n53913, n53914, n53915, n53916, n53917, n53918,
    n53919, n53920, n53921, n53922, n53923, n53924,
    n53925, n53926, n53927, n53928, n53929, n53930,
    n53931, n53932, n53933, n53934, n53935, n53936,
    n53937, n53938, n53939, n53940, n53941, n53942,
    n53943, n53944, n53945, n53946, n53947, n53948,
    n53949, n53950, n53951, n53952, n53953, n53954,
    n53955, n53956, n53957, n53958, n53959, n53960,
    n53961, n53962, n53963, n53964, n53965, n53966,
    n53967, n53968, n53969, n53970, n53971, n53972,
    n53973, n53974, n53975, n53976, n53977, n53978,
    n53979, n53980, n53981, n53982, n53983, n53984,
    n53985, n53986, n53987, n53988, n53989, n53990,
    n53991, n53992, n53993, n53994, n53995, n53996,
    n53997, n53998, n53999, n54000, n54001, n54002,
    n54003, n54004, n54005, n54006, n54007, n54008,
    n54009, n54010, n54011, n54012, n54013, n54014,
    n54015, n54016, n54017, n54018, n54019, n54020,
    n54021, n54022, n54023, n54024, n54025, n54026,
    n54027, n54028, n54029, n54030, n54031, n54032,
    n54033, n54034, n54035, n54036, n54037, n54038,
    n54039, n54040, n54041, n54042, n54043, n54044,
    n54045, n54046, n54047, n54048, n54049, n54050,
    n54051, n54052, n54053, n54054, n54055, n54056,
    n54057, n54058, n54059, n54060, n54061, n54062,
    n54063, n54064, n54065, n54066, n54067, n54068,
    n54069, n54070, n54071, n54072, n54073, n54074,
    n54075, n54076, n54077, n54078, n54079, n54080,
    n54081, n54082, n54083, n54084, n54085, n54086,
    n54087, n54088, n54089, n54090, n54091, n54092,
    n54093, n54094, n54095, n54096, n54097, n54098,
    n54099, n54100, n54101, n54102, n54103, n54104,
    n54105, n54106, n54107, n54108, n54109, n54110,
    n54111, n54112, n54113, n54114, n54115, n54116,
    n54117, n54118, n54119, n54120, n54121, n54122,
    n54123, n54124, n54125, n54126, n54127, n54128,
    n54129, n54130, n54131, n54132, n54133, n54134,
    n54135, n54136, n54137, n54138, n54139, n54140,
    n54141, n54142, n54143, n54144, n54145, n54146,
    n54147, n54148, n54149, n54150, n54151, n54152,
    n54153, n54154, n54155, n54156, n54157, n54158,
    n54159, n54160, n54161, n54162, n54163, n54164,
    n54165, n54166, n54167, n54168, n54169, n54170,
    n54171, n54172, n54173, n54174, n54175, n54176,
    n54177, n54178, n54179, n54180, n54181, n54182,
    n54183, n54184, n54185, n54186, n54187, n54188,
    n54189, n54190, n54191, n54192, n54193, n54194,
    n54195, n54196, n54197, n54198, n54199, n54200,
    n54201, n54202, n54203, n54204, n54205, n54206,
    n54207, n54208, n54209, n54210, n54211, n54212,
    n54213, n54214, n54215, n54216, n54217, n54218,
    n54219, n54220, n54221, n54222, n54223, n54224,
    n54225, n54226, n54227, n54228, n54229, n54230,
    n54231, n54232, n54233, n54234, n54235, n54236,
    n54237, n54238, n54239, n54240, n54241, n54242,
    n54243, n54244, n54245, n54246, n54247, n54248,
    n54249, n54250, n54251, n54252, n54253, n54254,
    n54255, n54256, n54257, n54258, n54259, n54260,
    n54261, n54262, n54263, n54264, n54265, n54266,
    n54267, n54268, n54269, n54270, n54271, n54272,
    n54273, n54274, n54275, n54276, n54277, n54278,
    n54279, n54280, n54281, n54282, n54283, n54284,
    n54285, n54286, n54287, n54288, n54289, n54290,
    n54291, n54292, n54293, n54294, n54295, n54296,
    n54297, n54298, n54299, n54300, n54301, n54302,
    n54303, n54304, n54305, n54306, n54307, n54308,
    n54309, n54310, n54311, n54312, n54313, n54314,
    n54315, n54316, n54317, n54318, n54319, n54320,
    n54321, n54322, n54323, n54324, n54325, n54326,
    n54327, n54328, n54329, n54330, n54331, n54332,
    n54333, n54334, n54335, n54336, n54337, n54338,
    n54339, n54340, n54341, n54342, n54343, n54344,
    n54345, n54346, n54347, n54348, n54349, n54350,
    n54351, n54352, n54353, n54354, n54355, n54356,
    n54357, n54358, n54359, n54360, n54361, n54362,
    n54363, n54364, n54365, n54366, n54367, n54368,
    n54369, n54370, n54371, n54372, n54373, n54374,
    n54375, n54376, n54377, n54378, n54379, n54380,
    n54381, n54382, n54383, n54384, n54385, n54386,
    n54387, n54388, n54389, n54390, n54391, n54392,
    n54393, n54394, n54395, n54396, n54397, n54398,
    n54399, n54400, n54401, n54402, n54403, n54404,
    n54405, n54406, n54407, n54408, n54409, n54410,
    n54411, n54412, n54413, n54414, n54415, n54416,
    n54417, n54418, n54419, n54420, n54421, n54422,
    n54423, n54424, n54425, n54426, n54427, n54428,
    n54429, n54430, n54431, n54432, n54433, n54434,
    n54435, n54436, n54437, n54438, n54439, n54440,
    n54441, n54442, n54443, n54444, n54445, n54446,
    n54447, n54448, n54449, n54450, n54451, n54452,
    n54453, n54454, n54455, n54456, n54457, n54458,
    n54459, n54460, n54461, n54462, n54463, n54464,
    n54465, n54466, n54467, n54468, n54469, n54470,
    n54471, n54472, n54473, n54474, n54475, n54476,
    n54477, n54478, n54479, n54480, n54481, n54482,
    n54483, n54484, n54485, n54486, n54487, n54488,
    n54489, n54490, n54491, n54492, n54493, n54494,
    n54495, n54496, n54497, n54498, n54499, n54500,
    n54501, n54502, n54503, n54504, n54505, n54506,
    n54507, n54508, n54509, n54510, n54511, n54512,
    n54513, n54514, n54515, n54516, n54517, n54518,
    n54519, n54520, n54521, n54522, n54523, n54524,
    n54525, n54526, n54527, n54528, n54529, n54530,
    n54531, n54532, n54533, n54534, n54535, n54536,
    n54537, n54538, n54539, n54540, n54541, n54542,
    n54543, n54544, n54545, n54546, n54547, n54548,
    n54549, n54550, n54551, n54552, n54553, n54554,
    n54555, n54556, n54557, n54558, n54559, n54560,
    n54561, n54562, n54563, n54564, n54565, n54566,
    n54567, n54568, n54569, n54570, n54571, n54572,
    n54573, n54574, n54575, n54576, n54577, n54578,
    n54579, n54580, n54581, n54582, n54583, n54584,
    n54585, n54586, n54587, n54588, n54589, n54590,
    n54591, n54592, n54593, n54594, n54595, n54596,
    n54597, n54598, n54599, n54600, n54601, n54602,
    n54603, n54604, n54605, n54606, n54607, n54608,
    n54609, n54610, n54611, n54612, n54613, n54614,
    n54615, n54616, n54617, n54618, n54619, n54620,
    n54621, n54622, n54623, n54624, n54625, n54626,
    n54627, n54628, n54629, n54630, n54631, n54632,
    n54633, n54634, n54635, n54636, n54637, n54638,
    n54639, n54640, n54641, n54642, n54643, n54644,
    n54645, n54646, n54647, n54648, n54649, n54650,
    n54651, n54652, n54653, n54654, n54655, n54656,
    n54657, n54658, n54659, n54660, n54661, n54662,
    n54663, n54664, n54665, n54666, n54667, n54668,
    n54669, n54670, n54671, n54672, n54673, n54674,
    n54675, n54676, n54677, n54678, n54679, n54680,
    n54681, n54682, n54683, n54684, n54685, n54686,
    n54687, n54688, n54689, n54690, n54691, n54692,
    n54693, n54694, n54695, n54696, n54697, n54698,
    n54699, n54700, n54701, n54702, n54703, n54704,
    n54705, n54706, n54707, n54708, n54709, n54710,
    n54711, n54712, n54713, n54714, n54715, n54716,
    n54717, n54718, n54719, n54720, n54721, n54722,
    n54723, n54724, n54725, n54726, n54727, n54728,
    n54729, n54730, n54731, n54732, n54733, n54734,
    n54735, n54736, n54737, n54738, n54739, n54740,
    n54741, n54742, n54743, n54744, n54745, n54746,
    n54747, n54748, n54749, n54750, n54751, n54752,
    n54753, n54754, n54755, n54756, n54757, n54758,
    n54759, n54760, n54761, n54762, n54763, n54764,
    n54765, n54766, n54767, n54768, n54769, n54770,
    n54771, n54772, n54773, n54774, n54775, n54776,
    n54777, n54778, n54779, n54780, n54781, n54782,
    n54783, n54784, n54785, n54786, n54787, n54788,
    n54789, n54790, n54791, n54792, n54793, n54794,
    n54795, n54796, n54797, n54798, n54799, n54800,
    n54801, n54802, n54803, n54804, n54805, n54806,
    n54807, n54808, n54809, n54810, n54811, n54812,
    n54813, n54814, n54815, n54816, n54817, n54818,
    n54819, n54820, n54821, n54822, n54823, n54824,
    n54825, n54826, n54827, n54828, n54829, n54830,
    n54831, n54832, n54833, n54834, n54835, n54836,
    n54837, n54838, n54839, n54840, n54841, n54842,
    n54843, n54844, n54845, n54846, n54847, n54848,
    n54849, n54850, n54851, n54852, n54853, n54854,
    n54855, n54856, n54857, n54858, n54859, n54860,
    n54861, n54862, n54863, n54864, n54865, n54866,
    n54867, n54868, n54869, n54870, n54871, n54872,
    n54873, n54874, n54875, n54876, n54877, n54878,
    n54879, n54880, n54881, n54882, n54883, n54884,
    n54885, n54886, n54887, n54888, n54889, n54890,
    n54891, n54892, n54893, n54894, n54895, n54896,
    n54897, n54898, n54899, n54900, n54901, n54902,
    n54903, n54904, n54905, n54906, n54907, n54908,
    n54909, n54910, n54911, n54912, n54913, n54914,
    n54915, n54916, n54917, n54918, n54919, n54920,
    n54921, n54922, n54923, n54924, n54925, n54926,
    n54927, n54928, n54929, n54930, n54931, n54932,
    n54933, n54934, n54935, n54936, n54937, n54938,
    n54939, n54940, n54941, n54942, n54943, n54944,
    n54945, n54946, n54947, n54948, n54949, n54950,
    n54951, n54952, n54953, n54954, n54955, n54956,
    n54957, n54958, n54959, n54960, n54961, n54962,
    n54963, n54964, n54965, n54966, n54967, n54968,
    n54969, n54970, n54971, n54972, n54973, n54974,
    n54975, n54976, n54977, n54978, n54979, n54980,
    n54981, n54982, n54983, n54984, n54985, n54986,
    n54987, n54988, n54989, n54990, n54991, n54992,
    n54993, n54994, n54995, n54996, n54997, n54998,
    n54999, n55000, n55001, n55002, n55003, n55004,
    n55005, n55006, n55007, n55008, n55009, n55010,
    n55011, n55012, n55013, n55014, n55015, n55016,
    n55017, n55018, n55019, n55020, n55021, n55022,
    n55023, n55024, n55025, n55026, n55027, n55028,
    n55029, n55030, n55031, n55032, n55033, n55034,
    n55035, n55036, n55037, n55038, n55039, n55040,
    n55041, n55042, n55043, n55044, n55045, n55046,
    n55047, n55048, n55049, n55050, n55051, n55052,
    n55053, n55054, n55055, n55056, n55057, n55058,
    n55059, n55060, n55061, n55062, n55063, n55064,
    n55065, n55066, n55067, n55068, n55069, n55070,
    n55071, n55072, n55073, n55074, n55075, n55076,
    n55077, n55078, n55079, n55080, n55081, n55082,
    n55083, n55084, n55085, n55086, n55087, n55088,
    n55089, n55090, n55091, n55092, n55093, n55094,
    n55095, n55096, n55097, n55098, n55099, n55100,
    n55101, n55102, n55103, n55104, n55105, n55106,
    n55107, n55108, n55109, n55110, n55111, n55112,
    n55113, n55114, n55115, n55116, n55117, n55118,
    n55119, n55120, n55121, n55122, n55123, n55124,
    n55125, n55126, n55127, n55128, n55129, n55130,
    n55131, n55132, n55133, n55134, n55135, n55136,
    n55137, n55138, n55139, n55140, n55141, n55142,
    n55143, n55144, n55145, n55146, n55147, n55148,
    n55149, n55150, n55151, n55152, n55153, n55154,
    n55155, n55156, n55157, n55158, n55159, n55160,
    n55161, n55162, n55163, n55164, n55165, n55166,
    n55167, n55168, n55169, n55170, n55171, n55172,
    n55173, n55174, n55175, n55176, n55177, n55178,
    n55179, n55180, n55181, n55182, n55183, n55184,
    n55185, n55186, n55187, n55188, n55189, n55190,
    n55191, n55192, n55193, n55194, n55195, n55196,
    n55197, n55198, n55199, n55200, n55201, n55202,
    n55203, n55204, n55205, n55206, n55207, n55208,
    n55209, n55210, n55211, n55212, n55213, n55214,
    n55215, n55216, n55217, n55218, n55219, n55220,
    n55221, n55222, n55223, n55224, n55225, n55226,
    n55227, n55228, n55229, n55230, n55231, n55232,
    n55233, n55234, n55235, n55236, n55237, n55238,
    n55239, n55240, n55241, n55242, n55243, n55244,
    n55245, n55246, n55247, n55248, n55249, n55250,
    n55251, n55252, n55253, n55254, n55255, n55256,
    n55257, n55258, n55259, n55260, n55261, n55262,
    n55263, n55264, n55265, n55266, n55267, n55268,
    n55269, n55270, n55271, n55272, n55273, n55274,
    n55275, n55276, n55277, n55278, n55279, n55280,
    n55281, n55282, n55283, n55284, n55285, n55286,
    n55287, n55288, n55289, n55290, n55291, n55292,
    n55293, n55294, n55295, n55296, n55297, n55298,
    n55299, n55300, n55301, n55302, n55303, n55304,
    n55305, n55306, n55307, n55308, n55309, n55310,
    n55311, n55312, n55313, n55314, n55315, n55316,
    n55317, n55318, n55319, n55320, n55321, n55322,
    n55323, n55324, n55325, n55326, n55327, n55328,
    n55329, n55330, n55331, n55332, n55333, n55334,
    n55335, n55336, n55337, n55338, n55339, n55340,
    n55341, n55342, n55343, n55344, n55345, n55346,
    n55347, n55348, n55349, n55350, n55351, n55352,
    n55353, n55354, n55355, n55356, n55357, n55358,
    n55359, n55360, n55361, n55362, n55363, n55364,
    n55365, n55366, n55367, n55368, n55369, n55370,
    n55371, n55372, n55373, n55374, n55375, n55376,
    n55377, n55378, n55379, n55380, n55381, n55382,
    n55383, n55384, n55385, n55386, n55387, n55388,
    n55389, n55390, n55391, n55392, n55393, n55394,
    n55395, n55396, n55397, n55398, n55399, n55400,
    n55401, n55402, n55403, n55404, n55405, n55406,
    n55407, n55408, n55409, n55410, n55411, n55412,
    n55413, n55414, n55415, n55416, n55417, n55418,
    n55419, n55420, n55421, n55422, n55423, n55424,
    n55425, n55426, n55427, n55428, n55429, n55430,
    n55431, n55432, n55433, n55434, n55435, n55436,
    n55437, n55438, n55439, n55440, n55441, n55442,
    n55443, n55444, n55445, n55446, n55447, n55448,
    n55449, n55450, n55451, n55452, n55453, n55454,
    n55455, n55456, n55457, n55458, n55459, n55460,
    n55461, n55462, n55463, n55464, n55465, n55466,
    n55467, n55468, n55469, n55470, n55471, n55472,
    n55473, n55474, n55475, n55476, n55477, n55478,
    n55479, n55480, n55481, n55482, n55483, n55484,
    n55485, n55486, n55487, n55488, n55489, n55490,
    n55491, n55492, n55493, n55494, n55495, n55496,
    n55497, n55498, n55499, n55500, n55501, n55502,
    n55503, n55504, n55505, n55506, n55507, n55508,
    n55509, n55510, n55511, n55512, n55513, n55514,
    n55515, n55516, n55517, n55518, n55519, n55520,
    n55521, n55522, n55523, n55524, n55525, n55526,
    n55527, n55528, n55529, n55530, n55531, n55532,
    n55533, n55534, n55535, n55536, n55537, n55538,
    n55539, n55540, n55541, n55542, n55543, n55544,
    n55545, n55546, n55547, n55548, n55549, n55550,
    n55551, n55552, n55553, n55554, n55555, n55556,
    n55557, n55558, n55559, n55560, n55561, n55562,
    n55563, n55564, n55565, n55566, n55567, n55568,
    n55569, n55570, n55571, n55572, n55573, n55574,
    n55575, n55576, n55577, n55578, n55579, n55580,
    n55581, n55582, n55583, n55584, n55585, n55586,
    n55587, n55588, n55589, n55590, n55591, n55592,
    n55593, n55594, n55595, n55596, n55597, n55598,
    n55599, n55600, n55601, n55602, n55603, n55604,
    n55605, n55606, n55607, n55608, n55609, n55610,
    n55611, n55612, n55613, n55614, n55615, n55616,
    n55617, n55618, n55619, n55620, n55621, n55622,
    n55623, n55624, n55625, n55626, n55627, n55628,
    n55629, n55630, n55631, n55632, n55633, n55634,
    n55635, n55636, n55637, n55638, n55639, n55640,
    n55641, n55642, n55643, n55644, n55645, n55646,
    n55647, n55648, n55649, n55650, n55651, n55652,
    n55653, n55654, n55655, n55656, n55657, n55658,
    n55659, n55660, n55661, n55662, n55663, n55664,
    n55665, n55666, n55667, n55668, n55669, n55670,
    n55671, n55672, n55673, n55674, n55675, n55676,
    n55677, n55678, n55679, n55680, n55681, n55682,
    n55683, n55684, n55685, n55686, n55687, n55688,
    n55689, n55690, n55691, n55692, n55693, n55694,
    n55695, n55696, n55697, n55698, n55699, n55700,
    n55701, n55702, n55703, n55704, n55705, n55706,
    n55707, n55708, n55709, n55710, n55711, n55712,
    n55713, n55714, n55715, n55716, n55717, n55718,
    n55719, n55720, n55721, n55722, n55723, n55724,
    n55725, n55726, n55727, n55728, n55729, n55730,
    n55731, n55732, n55733, n55734, n55735, n55736,
    n55737, n55738, n55739, n55740, n55741, n55742,
    n55743, n55744, n55745, n55746, n55747, n55748,
    n55749, n55750, n55751, n55752, n55753, n55754,
    n55755, n55756, n55757, n55758, n55759, n55760,
    n55761, n55762, n55763, n55764, n55765, n55766,
    n55767, n55768, n55769, n55770, n55771, n55772,
    n55773, n55774, n55775, n55776, n55777, n55778,
    n55779, n55780, n55781, n55782, n55783, n55784,
    n55785, n55786, n55787, n55788, n55789, n55790,
    n55791, n55792, n55793, n55794, n55795, n55796,
    n55797, n55798, n55799, n55800, n55801, n55802,
    n55803, n55804, n55805, n55806, n55807, n55808,
    n55809, n55810, n55811, n55812, n55813, n55814,
    n55815, n55816, n55817, n55818, n55819, n55820,
    n55821, n55822, n55823, n55824, n55825, n55826,
    n55827, n55828, n55829, n55830, n55831, n55832,
    n55833, n55834, n55835, n55836, n55837, n55838,
    n55839, n55840, n55841, n55842, n55843, n55844,
    n55845, n55846, n55847, n55848, n55849, n55850,
    n55851, n55852, n55853, n55854, n55855, n55856,
    n55857, n55858, n55859, n55860, n55861, n55862,
    n55863, n55864, n55865, n55866, n55867, n55868,
    n55869, n55870, n55871, n55872, n55873, n55874,
    n55875, n55876, n55877, n55878, n55879, n55880,
    n55881, n55882, n55883, n55884, n55885, n55886,
    n55887, n55888, n55889, n55890, n55891, n55892,
    n55893, n55894, n55895, n55896, n55897, n55898,
    n55899, n55900, n55901, n55902, n55903, n55904,
    n55905, n55906, n55907, n55908, n55909, n55910,
    n55911, n55912, n55913, n55914, n55915, n55916,
    n55917, n55918, n55919, n55920, n55921, n55922,
    n55923, n55924, n55925, n55926, n55927, n55928,
    n55929, n55930, n55931, n55932, n55933, n55934,
    n55935, n55936, n55937, n55938, n55939, n55940,
    n55941, n55942, n55943, n55944, n55945, n55946,
    n55947, n55948, n55949, n55950, n55951, n55952,
    n55953, n55954, n55955, n55956, n55957, n55958,
    n55959, n55960, n55961, n55962, n55963, n55964,
    n55965, n55966, n55967, n55968, n55969, n55970,
    n55971, n55972, n55973, n55974, n55975, n55976,
    n55977, n55978, n55979, n55980, n55981, n55982,
    n55983, n55984, n55985, n55986, n55987, n55988,
    n55989, n55990, n55991, n55992, n55993, n55994,
    n55995, n55996, n55997, n55998, n55999, n56000,
    n56001, n56002, n56003, n56004, n56005, n56006,
    n56007, n56008, n56009, n56010, n56011, n56012,
    n56013, n56014, n56015, n56016, n56017, n56018,
    n56019, n56020, n56021, n56022, n56023, n56024,
    n56025, n56026, n56027, n56028, n56029, n56030,
    n56031, n56032, n56033, n56034, n56035, n56036,
    n56037, n56038, n56039, n56040, n56041, n56042,
    n56043, n56044, n56045, n56046, n56047, n56048,
    n56049, n56050, n56051, n56052, n56053, n56054,
    n56055, n56056, n56057, n56058, n56059, n56060,
    n56061, n56062, n56063, n56064, n56065, n56066,
    n56067, n56068, n56069, n56070, n56071, n56072,
    n56073, n56074, n56075, n56076, n56077, n56078,
    n56079, n56080, n56081, n56082, n56083, n56084,
    n56085, n56086, n56087, n56088, n56089, n56090,
    n56091, n56092, n56093, n56094, n56095, n56096,
    n56097, n56098, n56099, n56100, n56101, n56102,
    n56103, n56104, n56105, n56106, n56107, n56108,
    n56109, n56110, n56111, n56112, n56113, n56114,
    n56115, n56116, n56117, n56118, n56119, n56120,
    n56121, n56122, n56123, n56124, n56125, n56126,
    n56127, n56128, n56129, n56130, n56131, n56132,
    n56133, n56134, n56135, n56136, n56137, n56138,
    n56139, n56140, n56141, n56142, n56143, n56144,
    n56145, n56146, n56147, n56148, n56149, n56150,
    n56151, n56152, n56153, n56154, n56155, n56156,
    n56157, n56158, n56159, n56160, n56161, n56162,
    n56163, n56164, n56165, n56166, n56167, n56168,
    n56169, n56170, n56171, n56172, n56173, n56174,
    n56175, n56176, n56177, n56178, n56179, n56180,
    n56181, n56182, n56183, n56184, n56185, n56186,
    n56187, n56188, n56189, n56190, n56191, n56192,
    n56193, n56194, n56195, n56196, n56197, n56198,
    n56199, n56200, n56201, n56202, n56203, n56204,
    n56205, n56206, n56207, n56208, n56209, n56210,
    n56211, n56212, n56213, n56214, n56215, n56216,
    n56217, n56218, n56219, n56220, n56221, n56222,
    n56223, n56224, n56225, n56226, n56227, n56228,
    n56229, n56230, n56231, n56232, n56233, n56234,
    n56235, n56236, n56237, n56238, n56239, n56240,
    n56241, n56242, n56243, n56244, n56245, n56246,
    n56247, n56248, n56249, n56250, n56251, n56252,
    n56253, n56254, n56255, n56256, n56257, n56258,
    n56259, n56260, n56261, n56262, n56263, n56264,
    n56265, n56266, n56267, n56268, n56269, n56270,
    n56271, n56272, n56273, n56274, n56275, n56276,
    n56277, n56278, n56279, n56280, n56281, n56282,
    n56283, n56284, n56285, n56286, n56287, n56288,
    n56289, n56290, n56291, n56292, n56293, n56294,
    n56295, n56296, n56297, n56298, n56299, n56300,
    n56301, n56302, n56303, n56304, n56305, n56306,
    n56307, n56308, n56309, n56310, n56311, n56312,
    n56313, n56314, n56315, n56316, n56317, n56318,
    n56319, n56320, n56321, n56322, n56323, n56324,
    n56325, n56326, n56327, n56328, n56329, n56330,
    n56331, n56332, n56333, n56334, n56335, n56336,
    n56337, n56338, n56339, n56340, n56341, n56342,
    n56343, n56344, n56345, n56346, n56347, n56348,
    n56349, n56350, n56351, n56352, n56353, n56354,
    n56355, n56356, n56357, n56358, n56359, n56360,
    n56361, n56362, n56363, n56364, n56365, n56366,
    n56367, n56368, n56369, n56370, n56371, n56372,
    n56373, n56374, n56375, n56376, n56377, n56378,
    n56379, n56380, n56381, n56382, n56383, n56384,
    n56385, n56386, n56387, n56388, n56389, n56390,
    n56391, n56392, n56393, n56394, n56395, n56396,
    n56397, n56398, n56399, n56400, n56401, n56402,
    n56403, n56404, n56405, n56406, n56407, n56408,
    n56409, n56410, n56411, n56412, n56413, n56414,
    n56415, n56416, n56417, n56418, n56419, n56420,
    n56421, n56422, n56423, n56424, n56425, n56426,
    n56427, n56428, n56429, n56430, n56431, n56432,
    n56433, n56434, n56435, n56436, n56437, n56438,
    n56439, n56440, n56441, n56442, n56443, n56444,
    n56445, n56446, n56447, n56448, n56449, n56450,
    n56451, n56452, n56453, n56454, n56455, n56456,
    n56457, n56458, n56459, n56460, n56461, n56462,
    n56463, n56464, n56465, n56466, n56467, n56468,
    n56469, n56470, n56471, n56472, n56473, n56474,
    n56475, n56476, n56477, n56478, n56479, n56480,
    n56481, n56482, n56483, n56484, n56485, n56486,
    n56487, n56488, n56489, n56490, n56491, n56492,
    n56493, n56494, n56495, n56496, n56497, n56498,
    n56499, n56500, n56501, n56502, n56503, n56504,
    n56505, n56506, n56507, n56508, n56509, n56510,
    n56511, n56512, n56513, n56514, n56515, n56516,
    n56517, n56518, n56519, n56520, n56521, n56522,
    n56523, n56524, n56525, n56526, n56527, n56528,
    n56529, n56530, n56531, n56532, n56533, n56534,
    n56535, n56536, n56537, n56538, n56539, n56540,
    n56541, n56542, n56543, n56544, n56545, n56546,
    n56547, n56548, n56549, n56550, n56551, n56552,
    n56553, n56554, n56555, n56556, n56557, n56558,
    n56559, n56560, n56561, n56562, n56563, n56564,
    n56565, n56566, n56567, n56568, n56569, n56570,
    n56571, n56572, n56573, n56574, n56575, n56576,
    n56577, n56578, n56579, n56580, n56581, n56582,
    n56583, n56584, n56585, n56586, n56587, n56588,
    n56589, n56590, n56591, n56592, n56593, n56594,
    n56595, n56596, n56597, n56598, n56599, n56600,
    n56601, n56602, n56603, n56604, n56605, n56606,
    n56607, n56608, n56609, n56610, n56611, n56612,
    n56613, n56614, n56615, n56616, n56617, n56618,
    n56619, n56620, n56621, n56622, n56623, n56624,
    n56625, n56626, n56627, n56628, n56629, n56630,
    n56631, n56632, n56633, n56634, n56635, n56636,
    n56637, n56638, n56639, n56640, n56641, n56642,
    n56643, n56644, n56645, n56646, n56647, n56648,
    n56649, n56650, n56651, n56652, n56653, n56654,
    n56655, n56656, n56657, n56658, n56659, n56660,
    n56661, n56662, n56663, n56664, n56665, n56666,
    n56667, n56668, n56669, n56670, n56671, n56672,
    n56673, n56674, n56675, n56676, n56677, n56678,
    n56679, n56680, n56681, n56682, n56683, n56684,
    n56685, n56686, n56687, n56688, n56689, n56690,
    n56691, n56692, n56693, n56694, n56695, n56696,
    n56697, n56698, n56699, n56700, n56701, n56702,
    n56703, n56704, n56705, n56706, n56707, n56708,
    n56709, n56710, n56711, n56712, n56713, n56714,
    n56715, n56716, n56717, n56718, n56719, n56720,
    n56721, n56722, n56723, n56724, n56725, n56726,
    n56727, n56728, n56729, n56730, n56731, n56732,
    n56733, n56734, n56735, n56736, n56737, n56738,
    n56739, n56740, n56741, n56742, n56743, n56744,
    n56745, n56746, n56747, n56748, n56749, n56750,
    n56751, n56752, n56753, n56754, n56755, n56756,
    n56757, n56758, n56759, n56760, n56761, n56762,
    n56763, n56764, n56765, n56766, n56767, n56768,
    n56769, n56770, n56771, n56772, n56773, n56774,
    n56775, n56776, n56777, n56778, n56779, n56780,
    n56781, n56782, n56783, n56784, n56785, n56786,
    n56787, n56788, n56789, n56790, n56791, n56792,
    n56793, n56794, n56795, n56796, n56797, n56798,
    n56799, n56800, n56801, n56802, n56803, n56804,
    n56805, n56806, n56807, n56808, n56809, n56810,
    n56811, n56812, n56813, n56814, n56815, n56816,
    n56817, n56818, n56819, n56820, n56821, n56822,
    n56823, n56824, n56825, n56826, n56827, n56828,
    n56829, n56830, n56831, n56832, n56833, n56834,
    n56835, n56836, n56837, n56838, n56839, n56840,
    n56841, n56842, n56843, n56844, n56845, n56846,
    n56847, n56848, n56849, n56850, n56851, n56852,
    n56853, n56854, n56855, n56856, n56857, n56858,
    n56859, n56860, n56861, n56862, n56863, n56864,
    n56865, n56866, n56867, n56868, n56869, n56870,
    n56871, n56872, n56873, n56874, n56875, n56876,
    n56877, n56878, n56879, n56880, n56881, n56882,
    n56883, n56884, n56885, n56886, n56887, n56888,
    n56889, n56890, n56891, n56892, n56893, n56894,
    n56895, n56896, n56897, n56898, n56899, n56900,
    n56901, n56902, n56903, n56904, n56905, n56906,
    n56907, n56908, n56909, n56910, n56911, n56912,
    n56913, n56914, n56915, n56916, n56917, n56918,
    n56919, n56920, n56921, n56922, n56923, n56924,
    n56925, n56926, n56927, n56928, n56929, n56930,
    n56931, n56932, n56933, n56934, n56935, n56936,
    n56937, n56938, n56939, n56940, n56941, n56942,
    n56943, n56944, n56945, n56946, n56947, n56948,
    n56949, n56950, n56951, n56952, n56953, n56954,
    n56955, n56956, n56957, n56958, n56959, n56960,
    n56961, n56962, n56963, n56964, n56965, n56966,
    n56967, n56968, n56969, n56970, n56971, n56972,
    n56973, n56974, n56975, n56976, n56977, n56978,
    n56979, n56980, n56981, n56982, n56983, n56984,
    n56985, n56986, n56987, n56988, n56989, n56990,
    n56991, n56992, n56993, n56994, n56995, n56996,
    n56997, n56998, n56999, n57000, n57001, n57002,
    n57003, n57004, n57005, n57006, n57007, n57008,
    n57009, n57010, n57011, n57012, n57013, n57014,
    n57015, n57016, n57017, n57018, n57019, n57020,
    n57021, n57022, n57023, n57024, n57025, n57026,
    n57027, n57028, n57029, n57030, n57031, n57032,
    n57033, n57034, n57035, n57036, n57037, n57038,
    n57039, n57040, n57041, n57042, n57043, n57044,
    n57045, n57046, n57047, n57048, n57049, n57050,
    n57051, n57052, n57053, n57054, n57055, n57056,
    n57057, n57058, n57059, n57060, n57061, n57062,
    n57063, n57064, n57065, n57066, n57067, n57068,
    n57069, n57070, n57071, n57072, n57073, n57074,
    n57075, n57076, n57077, n57078, n57079, n57080,
    n57081, n57082, n57083, n57084, n57085, n57086,
    n57087, n57088, n57089, n57090, n57091, n57092,
    n57093, n57094, n57095, n57096, n57097, n57098,
    n57099, n57100, n57101, n57102, n57103, n57104,
    n57105, n57106, n57107, n57108, n57109, n57110,
    n57111, n57112, n57113, n57114, n57115, n57116,
    n57117, n57118, n57119, n57120, n57121, n57122,
    n57123, n57124, n57125, n57126, n57127, n57128,
    n57129, n57130, n57131, n57132, n57133, n57134,
    n57135, n57136, n57137, n57138, n57139, n57140,
    n57141, n57142, n57143, n57144, n57145, n57146,
    n57147, n57148, n57149, n57150, n57151, n57152,
    n57153, n57154, n57155, n57156, n57157, n57158,
    n57159, n57160, n57161, n57162, n57163, n57164,
    n57165, n57166, n57167, n57168, n57169, n57170,
    n57171, n57172, n57173, n57174, n57175, n57176,
    n57177, n57178, n57179, n57180, n57181, n57182,
    n57183, n57184, n57185, n57186, n57187, n57188,
    n57189, n57190, n57191, n57192, n57193, n57194,
    n57195, n57196, n57197, n57198, n57199, n57200,
    n57201, n57202, n57203, n57204, n57205, n57206,
    n57207, n57208, n57209, n57210, n57211, n57212,
    n57213, n57214, n57215, n57216, n57217, n57218,
    n57219, n57220, n57221, n57222, n57223, n57224,
    n57225, n57226, n57227, n57228, n57229, n57230,
    n57231, n57232, n57233, n57234, n57235, n57236,
    n57237, n57238, n57239, n57240, n57241, n57242,
    n57243, n57244, n57245, n57246, n57247, n57248,
    n57249, n57250, n57251, n57252, n57253, n57254,
    n57255, n57256, n57257, n57258, n57259, n57260,
    n57261, n57262, n57263, n57264, n57265, n57266,
    n57267, n57268, n57269, n57270, n57271, n57272,
    n57273, n57274, n57275, n57276, n57277, n57278,
    n57279, n57280, n57281, n57282, n57283, n57284,
    n57285, n57286, n57287, n57288, n57289, n57290,
    n57291, n57292, n57293, n57294, n57295, n57296,
    n57297, n57298, n57299, n57300, n57301, n57302,
    n57303, n57304, n57305, n57306, n57307, n57308,
    n57309, n57310, n57311, n57312, n57313, n57314,
    n57315, n57316, n57317, n57318, n57319, n57320,
    n57321, n57322, n57323, n57324, n57325, n57326,
    n57327, n57328, n57329, n57330, n57331, n57332,
    n57333, n57334, n57335, n57336, n57337, n57338,
    n57339, n57340, n57341, n57342, n57343, n57344,
    n57345, n57346, n57347, n57348, n57349, n57350,
    n57351, n57352, n57353, n57354, n57355, n57356,
    n57357, n57358, n57359, n57360, n57361, n57362,
    n57363, n57364, n57365, n57366, n57367, n57368,
    n57369, n57370, n57371, n57372, n57373, n57374,
    n57375, n57376, n57377, n57378, n57379, n57380,
    n57381, n57382, n57383, n57384, n57385, n57386,
    n57387, n57388, n57389, n57390, n57391, n57392,
    n57393, n57394, n57395, n57396, n57397, n57398,
    n57399, n57400, n57401, n57402, n57403, n57404,
    n57405, n57406, n57407, n57408, n57409, n57410,
    n57411, n57412, n57413, n57414, n57415, n57416,
    n57417, n57418, n57419, n57420, n57421, n57422,
    n57423, n57424, n57425, n57426, n57427, n57428,
    n57429, n57430, n57431, n57432, n57433, n57434,
    n57435, n57436, n57437, n57438, n57439, n57440,
    n57441, n57442, n57443, n57444, n57445, n57446,
    n57447, n57448, n57449, n57450, n57451, n57452,
    n57453, n57454, n57455, n57456, n57457, n57458,
    n57459, n57460, n57461, n57462, n57463, n57464,
    n57465, n57466, n57467, n57468, n57469, n57470,
    n57471, n57472, n57473, n57474, n57475, n57476,
    n57477, n57478, n57479, n57480, n57481, n57482,
    n57483, n57484, n57485, n57486, n57487, n57488,
    n57489, n57490, n57491, n57492, n57493, n57494,
    n57495, n57496, n57497, n57498, n57499, n57500,
    n57501, n57502, n57503, n57504, n57505, n57506,
    n57507, n57508, n57509, n57510, n57511, n57512,
    n57513, n57514, n57515, n57516, n57517, n57518,
    n57519, n57520, n57521, n57522, n57523, n57524,
    n57525, n57526, n57527, n57528, n57529, n57530,
    n57531, n57532, n57533, n57534, n57535, n57536,
    n57537, n57538, n57539, n57540, n57541, n57542,
    n57543, n57544, n57545, n57546, n57547, n57548,
    n57549, n57550, n57551, n57552, n57553, n57554,
    n57555, n57556, n57557, n57558, n57559, n57560,
    n57561, n57562, n57563, n57564, n57565, n57566,
    n57567, n57568, n57569, n57570, n57571, n57572,
    n57573, n57574, n57575, n57576, n57577, n57578,
    n57579, n57580, n57581, n57582, n57583, n57584,
    n57585, n57586, n57587, n57588, n57589, n57590,
    n57591, n57592, n57593, n57594, n57595, n57596,
    n57597, n57598, n57599, n57600, n57601, n57602,
    n57603, n57604, n57605, n57606, n57607, n57608,
    n57609, n57610, n57611, n57612, n57613, n57614,
    n57615, n57616, n57617, n57618, n57619, n57620,
    n57621, n57622, n57623, n57624, n57625, n57626,
    n57627, n57628, n57629, n57630, n57631, n57632,
    n57633, n57634, n57635, n57636, n57637, n57638,
    n57639, n57640, n57641, n57642, n57643, n57644,
    n57645, n57646, n57647, n57648, n57649, n57650,
    n57651, n57652, n57653, n57654, n57655, n57656,
    n57657, n57658, n57659, n57660, n57661, n57662,
    n57663, n57664, n57665, n57666, n57667, n57668,
    n57669, n57670, n57671, n57672, n57673, n57674,
    n57675, n57676, n57677, n57678, n57679, n57680,
    n57681, n57682, n57683, n57684, n57685, n57686,
    n57687, n57688, n57689, n57690, n57691, n57692,
    n57693, n57694, n57695, n57696, n57697, n57698,
    n57699, n57700, n57701, n57702, n57703, n57704,
    n57705, n57706, n57707, n57708, n57709, n57710,
    n57711, n57712, n57713, n57714, n57715, n57716,
    n57717, n57718, n57719, n57720, n57721, n57722,
    n57723, n57724, n57725, n57726, n57727, n57728,
    n57729, n57730, n57731, n57732, n57733, n57734,
    n57735, n57736, n57737, n57738, n57739, n57740,
    n57741, n57742, n57743, n57744, n57745, n57746,
    n57747, n57748, n57749, n57750, n57751, n57752,
    n57753, n57754, n57755, n57756, n57757, n57758,
    n57759, n57760, n57761, n57762, n57763, n57764,
    n57765, n57766, n57767, n57768, n57769, n57770,
    n57771, n57772, n57773, n57774, n57775, n57776,
    n57777, n57778, n57779, n57780, n57781, n57782,
    n57783, n57784, n57785, n57786, n57787, n57788,
    n57789, n57790, n57791, n57792, n57793, n57794,
    n57795, n57796, n57797, n57798, n57799, n57800,
    n57801, n57802, n57803, n57804, n57805, n57806,
    n57807, n57808, n57809, n57810, n57811, n57812,
    n57813, n57814, n57815, n57816, n57817, n57818,
    n57819, n57820, n57821, n57822, n57823, n57824,
    n57825, n57826, n57827, n57828, n57829, n57830,
    n57831, n57832, n57833, n57834, n57835, n57836,
    n57837, n57838, n57839, n57840, n57841, n57842,
    n57843, n57844, n57845, n57846, n57847, n57848,
    n57849, n57850, n57851, n57852, n57853, n57854,
    n57855, n57856, n57857, n57858, n57859, n57860,
    n57861, n57862, n57863, n57864, n57865, n57866,
    n57867, n57868, n57869, n57870, n57871, n57872,
    n57873, n57874, n57875, n57876, n57877, n57878,
    n57879, n57880, n57881, n57882, n57883, n57884,
    n57885, n57886, n57887, n57888, n57889, n57890,
    n57891, n57892, n57893, n57894, n57895, n57896,
    n57897, n57898, n57899, n57900, n57901, n57902,
    n57903, n57904, n57905, n57906, n57907, n57908,
    n57909, n57910, n57911, n57912, n57913, n57914,
    n57915, n57916, n57917, n57918, n57919, n57920,
    n57921, n57922, n57923, n57924, n57925, n57926,
    n57927, n57928, n57929, n57930, n57931, n57932,
    n57933, n57934, n57935, n57936, n57937, n57938,
    n57939, n57940, n57941, n57942, n57943, n57944,
    n57945, n57946, n57947, n57948, n57949, n57950,
    n57951, n57952, n57953, n57954, n57955, n57956,
    n57957, n57958, n57959, n57960, n57961, n57962,
    n57963, n57964, n57965, n57966, n57967, n57968,
    n57969, n57970, n57971, n57972, n57973, n57974,
    n57975, n57976, n57977, n57978, n57979, n57980,
    n57981, n57982, n57983, n57984, n57985, n57986,
    n57987, n57988, n57989, n57990, n57991, n57992,
    n57993, n57994, n57995, n57996, n57997, n57998,
    n57999, n58000, n58001, n58002, n58003, n58004,
    n58005, n58006, n58007, n58008, n58009, n58010,
    n58011, n58012, n58013, n58014, n58015, n58016,
    n58017, n58018, n58019, n58020, n58021, n58022,
    n58023, n58024, n58025, n58026, n58027, n58028,
    n58029, n58030, n58031, n58032, n58033, n58034,
    n58035, n58036, n58037, n58038, n58039, n58040,
    n58041, n58042, n58043, n58044, n58045, n58046,
    n58047, n58048, n58049, n58050, n58051, n58052,
    n58053, n58054, n58055, n58056, n58057, n58058,
    n58059, n58060, n58061, n58062, n58063, n58064,
    n58065, n58066, n58067, n58068, n58069, n58070,
    n58071, n58072, n58073, n58074, n58075, n58076,
    n58077, n58078, n58079, n58080, n58081, n58082,
    n58083, n58084, n58085, n58086, n58087, n58088,
    n58089, n58090, n58091, n58092, n58093, n58094,
    n58095, n58096, n58097, n58098, n58099, n58100,
    n58101, n58102, n58103, n58104, n58105, n58106,
    n58107, n58108, n58109, n58110, n58111, n58112,
    n58113, n58114, n58115, n58116, n58117, n58118,
    n58119, n58120, n58121, n58122, n58123, n58124,
    n58125, n58126, n58127, n58128, n58129, n58130,
    n58131, n58132, n58133, n58134, n58135, n58136,
    n58137, n58138, n58139, n58140, n58141, n58142,
    n58143, n58144, n58145, n58146, n58147, n58148,
    n58149, n58150, n58151, n58152, n58153, n58154,
    n58155, n58156, n58157, n58158, n58159, n58160,
    n58161, n58162, n58163, n58164, n58165, n58166,
    n58167, n58168, n58169, n58170, n58171, n58172,
    n58173, n58174, n58175, n58176, n58177, n58178,
    n58179, n58180, n58181, n58182, n58183, n58184,
    n58185, n58186, n58187, n58188, n58189, n58190,
    n58191, n58192, n58193, n58194, n58195, n58196,
    n58197, n58198, n58199, n58200, n58201, n58202,
    n58203, n58204, n58205, n58206, n58207, n58208,
    n58209, n58210, n58211, n58212, n58213, n58214,
    n58215, n58216, n58217, n58218, n58219, n58220,
    n58221, n58222, n58223, n58224, n58225, n58226,
    n58227, n58228, n58229, n58230, n58231, n58232,
    n58233, n58234, n58235, n58236, n58237, n58238,
    n58239, n58240, n58241, n58242, n58243, n58244,
    n58245, n58246, n58247, n58248, n58249, n58250,
    n58251, n58252, n58253, n58254, n58255, n58256,
    n58257, n58258, n58259, n58260, n58261, n58262,
    n58263, n58264, n58265, n58266, n58267, n58268,
    n58269, n58270, n58271, n58272, n58273, n58274,
    n58275, n58276, n58277, n58278, n58279, n58280,
    n58281, n58282, n58283, n58284, n58285, n58286,
    n58287, n58288, n58289, n58290, n58291, n58292,
    n58293, n58294, n58295, n58296, n58297, n58298,
    n58299, n58300, n58301, n58302, n58303, n58304,
    n58305, n58306, n58307, n58308, n58309, n58310,
    n58311, n58312, n58313, n58314, n58315, n58316,
    n58317, n58318, n58319, n58320, n58321, n58322,
    n58323, n58324, n58325, n58326, n58327, n58328,
    n58329, n58330, n58331, n58332, n58333, n58334,
    n58335, n58336, n58337, n58338, n58339, n58340,
    n58341, n58342, n58343, n58344, n58345, n58346,
    n58347, n58348, n58349, n58350, n58351, n58352,
    n58353, n58354, n58355, n58356, n58357, n58358,
    n58359, n58360, n58361, n58362, n58363, n58364,
    n58365, n58366, n58367, n58368, n58369, n58370,
    n58371, n58372, n58373, n58374, n58375, n58376,
    n58377, n58378, n58379, n58380, n58381, n58382,
    n58383, n58384, n58385, n58386, n58387, n58388,
    n58389, n58390, n58391, n58392, n58393, n58394,
    n58395, n58396, n58397, n58398, n58399, n58400,
    n58401, n58402, n58403, n58404, n58405, n58406,
    n58407, n58408, n58409, n58410, n58411, n58412,
    n58413, n58414, n58415, n58416, n58417, n58418,
    n58419, n58420, n58421, n58422, n58423, n58424,
    n58425, n58426, n58427, n58428, n58429, n58430,
    n58431, n58432, n58433, n58434, n58435, n58436,
    n58437, n58438, n58439, n58440, n58441, n58442,
    n58443, n58444, n58445, n58446, n58447, n58448,
    n58449, n58450, n58451, n58452, n58453, n58454,
    n58455, n58456, n58457, n58458, n58459, n58460,
    n58461, n58462, n58463, n58464, n58465, n58466,
    n58467, n58468, n58469, n58470, n58471, n58472,
    n58473, n58474, n58475, n58476, n58477, n58478,
    n58479, n58480, n58481, n58482, n58483, n58484,
    n58485, n58486, n58487, n58488, n58489, n58490,
    n58491, n58492, n58493, n58494, n58495, n58496,
    n58497, n58498, n58499, n58500, n58501, n58502,
    n58503, n58504, n58505, n58506, n58507, n58508,
    n58509, n58510, n58511, n58512, n58513, n58514,
    n58515, n58516, n58517, n58518, n58519, n58520,
    n58521, n58522, n58523, n58524, n58525, n58526,
    n58527, n58528, n58529, n58530, n58531, n58532,
    n58533, n58534, n58535, n58536, n58537, n58538,
    n58539, n58540, n58541, n58542, n58543, n58544,
    n58545, n58546, n58547, n58548, n58549, n58550,
    n58551, n58552, n58553, n58554, n58555, n58556,
    n58557, n58558, n58559, n58560, n58561, n58562,
    n58563, n58564, n58565, n58566, n58567, n58568,
    n58569, n58570, n58571, n58572, n58573, n58574,
    n58575, n58576, n58577, n58578, n58579, n58580,
    n58581, n58582, n58583, n58584, n58585, n58586,
    n58587, n58588, n58589, n58590, n58591, n58592,
    n58593, n58594, n58595, n58596, n58597, n58598,
    n58599, n58600, n58601, n58602, n58603, n58604,
    n58605, n58606, n58607, n58608, n58609, n58610,
    n58611, n58612, n58613, n58614, n58615, n58616,
    n58617, n58618, n58619, n58620, n58621, n58622,
    n58623, n58624, n58625, n58626, n58627, n58628,
    n58629, n58630, n58631, n58632, n58633, n58634,
    n58635, n58636, n58637, n58638, n58639, n58640,
    n58641, n58642, n58643, n58644, n58645, n58646,
    n58647, n58648, n58649, n58650, n58651, n58652,
    n58653, n58654, n58655, n58656, n58657, n58658,
    n58659, n58660, n58661, n58662, n58663, n58664,
    n58665, n58666, n58667, n58668, n58669, n58670,
    n58671, n58672, n58673, n58674, n58675, n58676,
    n58677, n58678, n58679, n58680, n58681, n58682,
    n58683, n58684, n58685, n58686, n58687, n58688,
    n58689, n58690, n58691, n58692, n58693, n58694,
    n58695, n58696, n58697, n58698, n58699, n58700,
    n58701, n58702, n58703, n58704, n58705, n58706,
    n58707, n58708, n58709, n58710, n58711, n58712,
    n58713, n58714, n58715, n58716, n58717, n58718,
    n58719, n58720, n58721, n58722, n58723, n58724,
    n58725, n58726, n58727, n58728, n58729, n58730,
    n58731, n58732, n58733, n58734, n58735, n58736,
    n58737, n58738, n58739, n58740, n58741, n58742,
    n58743, n58744, n58745, n58746, n58747, n58748,
    n58749, n58750, n58751, n58752, n58753, n58754,
    n58755, n58756, n58757, n58758, n58759, n58760,
    n58761, n58762, n58763, n58764, n58765, n58766,
    n58767, n58768, n58769, n58770, n58771, n58772,
    n58773, n58774, n58775, n58776, n58777, n58778,
    n58779, n58780, n58781, n58782, n58783, n58784,
    n58785, n58786, n58787, n58788, n58789, n58790,
    n58791, n58792, n58793, n58794, n58795, n58796,
    n58797, n58798, n58799, n58800, n58801, n58802,
    n58803, n58804, n58805, n58806, n58807, n58808,
    n58809, n58810, n58811, n58812, n58813, n58814,
    n58815, n58816, n58817, n58818, n58819, n58820,
    n58821, n58822, n58823, n58824, n58825, n58826,
    n58827, n58828, n58829, n58830, n58831, n58832,
    n58833, n58834, n58835, n58836, n58837, n58838,
    n58839, n58840, n58841, n58842, n58843, n58844,
    n58845, n58846, n58847, n58848, n58849, n58850,
    n58851, n58852, n58853, n58854, n58855, n58856,
    n58857, n58858, n58859, n58860, n58861, n58862,
    n58863, n58864, n58865, n58866, n58867, n58868,
    n58869, n58870, n58871, n58872, n58873, n58874,
    n58875, n58876, n58877, n58878, n58879, n58880,
    n58881, n58882, n58883, n58884, n58885, n58886,
    n58887, n58888, n58889, n58890, n58891, n58892,
    n58893, n58894, n58895, n58896, n58897, n58898,
    n58899, n58900, n58901, n58902, n58903, n58904,
    n58905, n58906, n58907, n58908, n58909, n58910,
    n58911, n58912, n58913, n58914, n58915, n58916,
    n58917, n58918, n58919, n58920, n58921, n58922,
    n58923, n58924, n58925, n58926, n58927, n58928,
    n58929, n58930, n58931, n58932, n58933, n58934,
    n58935, n58936, n58937, n58938, n58939, n58940,
    n58941, n58942, n58943, n58944, n58945, n58946,
    n58947, n58948, n58949, n58950, n58951, n58952,
    n58953, n58954, n58955, n58956, n58957, n58958,
    n58959, n58960, n58961, n58962, n58963, n58964,
    n58965, n58966, n58967, n58968, n58969, n58970,
    n58971, n58972, n58973, n58974, n58975, n58976,
    n58977, n58978, n58979, n58980, n58981, n58982,
    n58983, n58984, n58985, n58986, n58987, n58988,
    n58989, n58990, n58991, n58992, n58993, n58994,
    n58995, n58996, n58997, n58998, n58999, n59000,
    n59001, n59002, n59003, n59004, n59005, n59006,
    n59007, n59008, n59009, n59010, n59011, n59012,
    n59013, n59014, n59015, n59016, n59017, n59018,
    n59019, n59020, n59021, n59022, n59023, n59024,
    n59025, n59026, n59027, n59028, n59029, n59030,
    n59031, n59032, n59033, n59034, n59035, n59036,
    n59037, n59038, n59039, n59040, n59041, n59042,
    n59043, n59044, n59045, n59046, n59047, n59048,
    n59049, n59050, n59051, n59052, n59053, n59054,
    n59055, n59056, n59057, n59058, n59059, n59060,
    n59061, n59062, n59063, n59064, n59065, n59066,
    n59067, n59068, n59069, n59070, n59071, n59072,
    n59073, n59074, n59075, n59076, n59077, n59078,
    n59079, n59080, n59081, n59082, n59083, n59084,
    n59085, n59086, n59087, n59088, n59089, n59090,
    n59091, n59092, n59093, n59094, n59095, n59096,
    n59097, n59098, n59099, n59100, n59101, n59102,
    n59103, n59104, n59105, n59106, n59107, n59108,
    n59109, n59110, n59111, n59112, n59113, n59114,
    n59115, n59116, n59117, n59118, n59119, n59120,
    n59121, n59122, n59123, n59124, n59125, n59126,
    n59127, n59128, n59129, n59130, n59131, n59132,
    n59133, n59134, n59135, n59136, n59137, n59138,
    n59139, n59140, n59141, n59142, n59143, n59144,
    n59145, n59146, n59147, n59148, n59149, n59150,
    n59151, n59152, n59153, n59154, n59155, n59156,
    n59157, n59158, n59159, n59160, n59161, n59162,
    n59163, n59164, n59165, n59166, n59167, n59168,
    n59169, n59170, n59171, n59172, n59173, n59174,
    n59175, n59176, n59177, n59178, n59179, n59180,
    n59181, n59182, n59183, n59184, n59185, n59186,
    n59187, n59188, n59189, n59190, n59191, n59192,
    n59193, n59194, n59195, n59196, n59197, n59198,
    n59199, n59200, n59201, n59202, n59203, n59204,
    n59205, n59206, n59207, n59208, n59209, n59210,
    n59211, n59212, n59213, n59214, n59215, n59216,
    n59217, n59218, n59219, n59220, n59221, n59222,
    n59223, n59224, n59225, n59226, n59227, n59228,
    n59229, n59230, n59231, n59232, n59233, n59234,
    n59235, n59236, n59237, n59238, n59239, n59240,
    n59241, n59242, n59243, n59244, n59245, n59246,
    n59247, n59248, n59249, n59250, n59251, n59252,
    n59253, n59254, n59255, n59256, n59257, n59258,
    n59259, n59260, n59261, n59262, n59263, n59264,
    n59265, n59266, n59267, n59268, n59269, n59270,
    n59271, n59272, n59273, n59274, n59275, n59276,
    n59277, n59278, n59279, n59280, n59281, n59282,
    n59283, n59284, n59285, n59286, n59287, n59288,
    n59289, n59290, n59291, n59292, n59293, n59294,
    n59295, n59296, n59297, n59298, n59299, n59300,
    n59301, n59302, n59303, n59304, n59305, n59306,
    n59307, n59308, n59309, n59310, n59311, n59312,
    n59313, n59314, n59315, n59316, n59317, n59318,
    n59319, n59320, n59321, n59322, n59323, n59324,
    n59325, n59326, n59327, n59328, n59329, n59330,
    n59331, n59332, n59333, n59334, n59335, n59336,
    n59337, n59338, n59339, n59340, n59341, n59342,
    n59343, n59344, n59345, n59346, n59347, n59348,
    n59349, n59350, n59351, n59352, n59353, n59354,
    n59355, n59356, n59357, n59358, n59359, n59360,
    n59361, n59362, n59363, n59364, n59365, n59366,
    n59367, n59368, n59369, n59370, n59371, n59372,
    n59373, n59374, n59375, n59376, n59377, n59378,
    n59379, n59380, n59381, n59382, n59383, n59384,
    n59385, n59386, n59387, n59388, n59389, n59390,
    n59391, n59392, n59393, n59394, n59395, n59396,
    n59397, n59398, n59399, n59400, n59401, n59402,
    n59403, n59404, n59405, n59406, n59407, n59408,
    n59409, n59410, n59411, n59412, n59413, n59414,
    n59415, n59416, n59417, n59418, n59419, n59420,
    n59421, n59422, n59423, n59424, n59425, n59426,
    n59427, n59428, n59429, n59430, n59431, n59432,
    n59433, n59434, n59435, n59436, n59437, n59438,
    n59439, n59440, n59441, n59442, n59443, n59444,
    n59445, n59446, n59447, n59448, n59449, n59450,
    n59451, n59452, n59453, n59454, n59455, n59456,
    n59457, n59458, n59459, n59460, n59461, n59462,
    n59463, n59464, n59465, n59466, n59467, n59468,
    n59469, n59470, n59471, n59472, n59473, n59474,
    n59475, n59476, n59477, n59478, n59479, n59480,
    n59481, n59482, n59483, n59484, n59485, n59486,
    n59487, n59488, n59489, n59490, n59491, n59492,
    n59493, n59494, n59495, n59496, n59497, n59498,
    n59499, n59500, n59501, n59502, n59503, n59504,
    n59505, n59506, n59507, n59508, n59509, n59510,
    n59511, n59512, n59513, n59514, n59515, n59516,
    n59517, n59518, n59519, n59520, n59521, n59522,
    n59523, n59524, n59525, n59526, n59527, n59528,
    n59529, n59530, n59531, n59532, n59533, n59534,
    n59535, n59536, n59537, n59538, n59539, n59540,
    n59541, n59542, n59543, n59544, n59545, n59546,
    n59547, n59548, n59549, n59550, n59551, n59552,
    n59553, n59554, n59555, n59556, n59557, n59558,
    n59559, n59560, n59561, n59562, n59563, n59564,
    n59565, n59566, n59567, n59568, n59569, n59570,
    n59571, n59572, n59573, n59574, n59575, n59576,
    n59577, n59578, n59579, n59580, n59581, n59582,
    n59583, n59584, n59585, n59586, n59587, n59588,
    n59589, n59590, n59591, n59592, n59593, n59594,
    n59595, n59596, n59597, n59598, n59599, n59600,
    n59601, n59602, n59603, n59604, n59605, n59606,
    n59607, n59608, n59609, n59610, n59611, n59612,
    n59613, n59614, n59615, n59616, n59617, n59618,
    n59619, n59620, n59621, n59622, n59623, n59624,
    n59625, n59626, n59627, n59628, n59629, n59630,
    n59631, n59632, n59633, n59634, n59635, n59636,
    n59637, n59638, n59639, n59640, n59641, n59642,
    n59643, n59644, n59645, n59646, n59647, n59648,
    n59649, n59650, n59651, n59652, n59653, n59654,
    n59655, n59656, n59657, n59658, n59659, n59660,
    n59661, n59662, n59663, n59664, n59665, n59666,
    n59667, n59668, n59669, n59670, n59671, n59672,
    n59673, n59674, n59675, n59676, n59677, n59678,
    n59679, n59680, n59681, n59682, n59683, n59684,
    n59685, n59686, n59687, n59688, n59689, n59690,
    n59691, n59692, n59693, n59694, n59695, n59696,
    n59697, n59698, n59699, n59700, n59701, n59702,
    n59703, n59704, n59705, n59706, n59707, n59708,
    n59709, n59710, n59711, n59712, n59713, n59714,
    n59715, n59716, n59717, n59718, n59719, n59720,
    n59721, n59722, n59723, n59724, n59725, n59726,
    n59727, n59728, n59729, n59730, n59731, n59732,
    n59733, n59734, n59735, n59736, n59737, n59738,
    n59739, n59740, n59741, n59742, n59743, n59744,
    n59745, n59746, n59747, n59748, n59749, n59750,
    n59751, n59752, n59753, n59754, n59755, n59756,
    n59757, n59758, n59759, n59760, n59761, n59762,
    n59763, n59764, n59765, n59766, n59767, n59768,
    n59769, n59770, n59771, n59772, n59773, n59774,
    n59775, n59776, n59777, n59778, n59779, n59780,
    n59781, n59782, n59783, n59784, n59785, n59786,
    n59787, n59788, n59789, n59790, n59791, n59792,
    n59793, n59794, n59795, n59796, n59797, n59798,
    n59799, n59800, n59801, n59802, n59803, n59804,
    n59805, n59806, n59807, n59808, n59809, n59810,
    n59811, n59812, n59813, n59814, n59815, n59816,
    n59817, n59818, n59819, n59820, n59821, n59822,
    n59823, n59824, n59825, n59826, n59827, n59828,
    n59829, n59830, n59831, n59832, n59833, n59834,
    n59835, n59836, n59837, n59838, n59839, n59840,
    n59841, n59842, n59843, n59844, n59845, n59846,
    n59847, n59848, n59849, n59850, n59851, n59852,
    n59853, n59854, n59855, n59856, n59857, n59858,
    n59859, n59860, n59861, n59862, n59863, n59864,
    n59865, n59866, n59867, n59868, n59869, n59870,
    n59871, n59872, n59873, n59874, n59875, n59876,
    n59877, n59878, n59879, n59880, n59881, n59882,
    n59883, n59884, n59885, n59886, n59887, n59888,
    n59889, n59890, n59891, n59892, n59893, n59894,
    n59895, n59896, n59897, n59898, n59899, n59900,
    n59901, n59902, n59903, n59904, n59905, n59906,
    n59907, n59908, n59909, n59910, n59911, n59912,
    n59913, n59914, n59915, n59916, n59917, n59918,
    n59919, n59920, n59921, n59922, n59923, n59924,
    n59925, n59926, n59927, n59928, n59929, n59930,
    n59931, n59932, n59933, n59934, n59935, n59936,
    n59937, n59938, n59939, n59940, n59941, n59942,
    n59943, n59944, n59945, n59946, n59947, n59948,
    n59949, n59950, n59951, n59952, n59953, n59954,
    n59955, n59956, n59957, n59958, n59959, n59960,
    n59961, n59962, n59963, n59964, n59965, n59966,
    n59967, n59968, n59969, n59970, n59971, n59972,
    n59973, n59974, n59975, n59976, n59977, n59978,
    n59979, n59980, n59981, n59982, n59983, n59984,
    n59985, n59986, n59987, n59988, n59989, n59990,
    n59991, n59992, n59993, n59994, n59995, n59996,
    n59997, n59998, n59999, n60000, n60001, n60002,
    n60003, n60004, n60005, n60006, n60007, n60008,
    n60009, n60010, n60011, n60012, n60013, n60014,
    n60015, n60016, n60017, n60018, n60019, n60020,
    n60021, n60022, n60023, n60024, n60025, n60026,
    n60027, n60028, n60029, n60030, n60031, n60032,
    n60033, n60034, n60035, n60036, n60037, n60038,
    n60039, n60040, n60041, n60042, n60043, n60044,
    n60045, n60046, n60047, n60048, n60049, n60050,
    n60051, n60052, n60053, n60054, n60055, n60056,
    n60057, n60058, n60059, n60060, n60061, n60062,
    n60063, n60064, n60065, n60066, n60067, n60068,
    n60069, n60070, n60071, n60072, n60073, n60074,
    n60075, n60076, n60077, n60078, n60079, n60080,
    n60081, n60082, n60083, n60084, n60085, n60086,
    n60087, n60088, n60089, n60090, n60091, n60092,
    n60093, n60094, n60095, n60096, n60097, n60098,
    n60099, n60100, n60101, n60102, n60103, n60104,
    n60105, n60106, n60107, n60108, n60109, n60110,
    n60111, n60112, n60113, n60114, n60115, n60116,
    n60117, n60118, n60119, n60120, n60121, n60122,
    n60123, n60124, n60125, n60126, n60127, n60128,
    n60129, n60130, n60131, n60132, n60133, n60134,
    n60135, n60136, n60137, n60138, n60139, n60140,
    n60141, n60142, n60143, n60144, n60145, n60146,
    n60147, n60148, n60149, n60150, n60151, n60152,
    n60153, n60154, n60155, n60156, n60157, n60158,
    n60159, n60160, n60161, n60162, n60163, n60164,
    n60165, n60166, n60167, n60168, n60169, n60170,
    n60171, n60172, n60173, n60174, n60175, n60176,
    n60177, n60178, n60179, n60180, n60181, n60182,
    n60183, n60184, n60185, n60186, n60187, n60188,
    n60189, n60190, n60191, n60192, n60193, n60194,
    n60195, n60196, n60197, n60198, n60199, n60200,
    n60201, n60202, n60203, n60204, n60205, n60206,
    n60207, n60208, n60209, n60210, n60211, n60212,
    n60213, n60214, n60215, n60216, n60217, n60218,
    n60219, n60220, n60221, n60222, n60223, n60224,
    n60225, n60226, n60227, n60228, n60229, n60230,
    n60231, n60232, n60233, n60234, n60235, n60236,
    n60237, n60238, n60239, n60240, n60241, n60242,
    n60243, n60244, n60245, n60246, n60247, n60248,
    n60249, n60250, n60251, n60252, n60253, n60254,
    n60255, n60256, n60257, n60258, n60259, n60260,
    n60261, n60262, n60263, n60264, n60265, n60266,
    n60267, n60268, n60269, n60270, n60271, n60272,
    n60273, n60274, n60275, n60276, n60277, n60278,
    n60279, n60280, n60281, n60282, n60283, n60284,
    n60285, n60286, n60287, n60288, n60289, n60290,
    n60291, n60292, n60293, n60294, n60295, n60296,
    n60297, n60298, n60299, n60300, n60301, n60302,
    n60303, n60304, n60305, n60306, n60307, n60308,
    n60309, n60310, n60311, n60312, n60313, n60314,
    n60315, n60316, n60317, n60318, n60319, n60320,
    n60321, n60322, n60323, n60324, n60325, n60326,
    n60327, n60328, n60329, n60330, n60331, n60332,
    n60333, n60334, n60335, n60336, n60337, n60338,
    n60339, n60340, n60341, n60342, n60343, n60344,
    n60345, n60346, n60347, n60348, n60349, n60350,
    n60351, n60352, n60353, n60354, n60355, n60356,
    n60357, n60358, n60359, n60360, n60361, n60362,
    n60363, n60364, n60365, n60366, n60367, n60368,
    n60369, n60370, n60371, n60372, n60373, n60374,
    n60375, n60376, n60377, n60378, n60379, n60380,
    n60381, n60382, n60383, n60384, n60385, n60386,
    n60387, n60388, n60389, n60390, n60391, n60392,
    n60393, n60394, n60395, n60396, n60397, n60398,
    n60399, n60400, n60401, n60402;
  assign n65 = pi2  & ~pi3 ;
  assign n66 = ~pi2  & pi3 ;
  assign n67 = ~pi2  & ~pi3 ;
  assign n68 = pi2  & pi3 ;
  assign n69 = ~n67 & ~n68;
  assign n70 = ~n65 & ~n66;
  assign n71 = pi4  & ~pi5 ;
  assign n72 = ~pi4  & pi5 ;
  assign n73 = ~pi4  & ~pi5 ;
  assign n74 = pi4  & pi5 ;
  assign n75 = ~n73 & ~n74;
  assign n76 = ~n71 & ~n72;
  assign n77 = n53439 & n53440;
  assign n78 = pi20  & ~pi21 ;
  assign n79 = ~pi20  & pi21 ;
  assign n80 = ~pi20  & ~pi21 ;
  assign n81 = pi20  & pi21 ;
  assign n82 = ~n80 & ~n81;
  assign n83 = ~n78 & ~n79;
  assign n84 = pi22  & ~pi23 ;
  assign n85 = ~pi22  & pi23 ;
  assign n86 = ~pi22  & ~pi23 ;
  assign n87 = pi22  & pi23 ;
  assign n88 = ~n86 & ~n87;
  assign n89 = ~n84 & ~n85;
  assign n90 = n53441 & n53442;
  assign n91 = ~pi27  & pi28 ;
  assign n92 = ~pi29  & pi30 ;
  assign n93 = pi29  & ~pi30 ;
  assign n94 = ~n92 & ~n93;
  assign n95 = pi30  & n94;
  assign n96 = pi29  & pi30 ;
  assign n97 = n91 & n53443;
  assign n98 = ~pi24  & ~pi25 ;
  assign n99 = pi23  & pi26 ;
  assign n100 = n98 & n99;
  assign n101 = n97 & n100;
  assign n102 = ~pi24  & pi25 ;
  assign n103 = ~pi23  & ~pi26 ;
  assign n104 = n102 & n103;
  assign n105 = n97 & n104;
  assign n106 = ~n101 & ~n105;
  assign n107 = n98 & n103;
  assign n108 = n97 & n107;
  assign n109 = pi23  & ~pi26 ;
  assign n110 = pi24  & ~pi25 ;
  assign n111 = n109 & n110;
  assign n112 = n97 & n111;
  assign n113 = ~n108 & ~n112;
  assign n114 = pi24  & pi25 ;
  assign n115 = ~pi25  & pi26 ;
  assign n116 = pi25  & ~pi26 ;
  assign n117 = ~n115 & ~n116;
  assign n118 = ~pi23  & pi24 ;
  assign n119 = pi23  & ~pi24 ;
  assign n120 = ~n118 & ~n119;
  assign n121 = ~n98 & ~n114;
  assign n122 = n120 & ~n121;
  assign n123 = ~n117 & ~n120;
  assign n124 = ~n117 & n120;
  assign n125 = ~n121 & n124;
  assign n126 = ~n117 & n122;
  assign n127 = n120 & n121;
  assign n128 = n117 & ~n120;
  assign n129 = ~n127 & ~n128;
  assign n130 = ~n53444 & n129;
  assign n131 = ~n123 & n130;
  assign n132 = ~n123 & ~n53444;
  assign n133 = n129 & n132;
  assign n134 = n117 & n122;
  assign n135 = pi26  & ~n53445;
  assign n136 = pi26  & ~n135;
  assign n137 = pi26  & n53445;
  assign n138 = n99 & n114;
  assign n139 = pi27  & ~pi28 ;
  assign n140 = n53443 & n139;
  assign n141 = n53446 & n140;
  assign n142 = ~pi23  & pi26 ;
  assign n143 = n98 & n142;
  assign n144 = n97 & n143;
  assign n145 = ~n141 & ~n144;
  assign n146 = ~n108 & ~n144;
  assign n147 = ~n112 & ~n141;
  assign n148 = n146 & n147;
  assign n149 = n113 & n145;
  assign n150 = ~n101 & n113;
  assign n151 = ~n105 & n150;
  assign n152 = ~n144 & n151;
  assign n153 = ~n141 & n152;
  assign n154 = ~n105 & ~n144;
  assign n155 = ~n101 & ~n112;
  assign n156 = ~n108 & ~n141;
  assign n157 = n155 & n156;
  assign n158 = n154 & n157;
  assign n159 = n106 & n53447;
  assign n160 = n114 & n142;
  assign n161 = n140 & n160;
  assign n162 = n99 & n110;
  assign n163 = n97 & n162;
  assign n164 = ~n161 & ~n163;
  assign n165 = n99 & n102;
  assign n166 = n140 & n165;
  assign n167 = n109 & n114;
  assign n168 = n97 & n167;
  assign n169 = ~n166 & ~n168;
  assign n170 = n164 & n169;
  assign n171 = n103 & n110;
  assign n172 = n97 & n171;
  assign n173 = n110 & n142;
  assign n174 = n97 & n173;
  assign n175 = ~n172 & ~n174;
  assign n176 = n102 & n109;
  assign n177 = n97 & n176;
  assign n178 = n103 & n114;
  assign n179 = n97 & n178;
  assign n180 = ~n177 & ~n179;
  assign n181 = n102 & n142;
  assign n182 = n140 & n181;
  assign n183 = n98 & n109;
  assign n184 = n97 & n183;
  assign n185 = ~n182 & ~n184;
  assign n186 = n180 & n185;
  assign n187 = n175 & n186;
  assign n188 = n169 & n180;
  assign n189 = n164 & n175;
  assign n190 = n175 & n185;
  assign n191 = n164 & n190;
  assign n192 = n185 & n189;
  assign n193 = n188 & n53449;
  assign n194 = n169 & n175;
  assign n195 = n164 & n185;
  assign n196 = n180 & n195;
  assign n197 = n194 & n196;
  assign n198 = n170 & n187;
  assign n199 = n53448 & n185;
  assign n200 = n180 & n199;
  assign n201 = n175 & n200;
  assign n202 = n164 & n201;
  assign n203 = ~n168 & n202;
  assign n204 = ~n166 & n203;
  assign n205 = n53448 & n53450;
  assign n206 = n140 & n178;
  assign n207 = n140 & n162;
  assign n208 = ~n206 & ~n207;
  assign n209 = ~pi27  & ~pi28 ;
  assign n210 = n53443 & n209;
  assign n211 = n162 & n210;
  assign n212 = n53446 & n210;
  assign n213 = ~n211 & ~n212;
  assign n214 = n208 & n213;
  assign n215 = n160 & n210;
  assign n216 = n140 & n171;
  assign n217 = ~n215 & ~n216;
  assign n218 = n104 & n140;
  assign n219 = n173 & n210;
  assign n220 = ~n218 & ~n219;
  assign n221 = n140 & n176;
  assign n222 = n100 & n140;
  assign n223 = ~n221 & ~n222;
  assign n224 = n220 & n223;
  assign n225 = n217 & n223;
  assign n226 = n220 & n225;
  assign n227 = n217 & n224;
  assign n228 = n208 & n217;
  assign n229 = ~n219 & n228;
  assign n230 = ~n211 & n229;
  assign n231 = ~n212 & n230;
  assign n232 = ~n218 & n231;
  assign n233 = ~n222 & n232;
  assign n234 = ~n221 & n233;
  assign n235 = n213 & n220;
  assign n236 = n208 & n223;
  assign n237 = n217 & n236;
  assign n238 = n235 & n237;
  assign n239 = ~n211 & ~n219;
  assign n240 = n223 & n239;
  assign n241 = ~n212 & ~n218;
  assign n242 = n208 & n241;
  assign n243 = n217 & n242;
  assign n244 = n240 & n243;
  assign n245 = n214 & n53452;
  assign n246 = n140 & n167;
  assign n247 = n165 & n210;
  assign n248 = ~n246 & ~n247;
  assign n249 = n140 & n173;
  assign n250 = n143 & n210;
  assign n251 = ~n249 & ~n250;
  assign n252 = n248 & ~n250;
  assign n253 = ~n249 & n252;
  assign n254 = n248 & n251;
  assign n255 = n111 & n140;
  assign n256 = n107 & n140;
  assign n257 = ~n255 & ~n256;
  assign n258 = n181 & n210;
  assign n259 = n140 & n143;
  assign n260 = ~n258 & ~n259;
  assign n261 = n257 & n260;
  assign n262 = n53454 & n257;
  assign n263 = ~n258 & n262;
  assign n264 = ~n259 & n263;
  assign n265 = n53454 & n261;
  assign n266 = ~pi29  & ~pi30 ;
  assign n267 = n209 & n266;
  assign n268 = n107 & n267;
  assign n269 = n183 & n267;
  assign n270 = ~n268 & ~n269;
  assign n271 = n100 & n210;
  assign n272 = n140 & n183;
  assign n273 = ~n271 & ~n272;
  assign n274 = n171 & n267;
  assign n275 = n111 & n267;
  assign n276 = ~n274 & ~n275;
  assign n277 = n273 & n276;
  assign n278 = n270 & n273;
  assign n279 = n276 & n278;
  assign n280 = n270 & n277;
  assign n281 = n53455 & n53456;
  assign n282 = n53453 & n53455;
  assign n283 = n276 & n282;
  assign n284 = ~n271 & n283;
  assign n285 = ~n272 & n284;
  assign n286 = ~n269 & n285;
  assign n287 = ~n268 & n286;
  assign n288 = n53453 & n281;
  assign n289 = pi27  & pi28 ;
  assign n290 = n92 & n289;
  assign n291 = n160 & n290;
  assign n292 = n104 & n210;
  assign n293 = ~n291 & ~n292;
  assign n294 = n176 & n210;
  assign n295 = n53446 & n290;
  assign n296 = n181 & n290;
  assign n297 = ~n295 & ~n296;
  assign n298 = ~n294 & ~n295;
  assign n299 = ~n296 & n298;
  assign n300 = ~n294 & n297;
  assign n301 = n293 & ~n295;
  assign n302 = ~n296 & n301;
  assign n303 = ~n294 & n302;
  assign n304 = n293 & ~n294;
  assign n305 = n297 & n304;
  assign n306 = n293 & n53458;
  assign n307 = n107 & n210;
  assign n308 = n178 & n210;
  assign n309 = ~n307 & ~n308;
  assign n310 = n111 & n210;
  assign n311 = n171 & n210;
  assign n312 = ~n310 & ~n311;
  assign n313 = n309 & ~n310;
  assign n314 = ~n311 & n313;
  assign n315 = n309 & n312;
  assign n316 = n165 & n290;
  assign n317 = n167 & n210;
  assign n318 = ~n316 & ~n317;
  assign n319 = n104 & n267;
  assign n320 = n162 & n290;
  assign n321 = n183 & n210;
  assign n322 = ~n320 & ~n321;
  assign n323 = ~n319 & n322;
  assign n324 = n318 & ~n319;
  assign n325 = n322 & n324;
  assign n326 = n318 & n323;
  assign n327 = n53460 & n318;
  assign n328 = n323 & n327;
  assign n329 = n53460 & n53461;
  assign n330 = n53459 & n53462;
  assign n331 = n53457 & n330;
  assign n332 = n53459 & n53460;
  assign n333 = n53451 & n332;
  assign n334 = n53457 & n333;
  assign n335 = n322 & n334;
  assign n336 = n318 & n335;
  assign n337 = ~n319 & n336;
  assign n338 = n53451 & n331;
  assign n339 = n93 & n139;
  assign n340 = n171 & n339;
  assign n341 = n91 & n93;
  assign n342 = n171 & n341;
  assign n343 = ~n340 & ~n342;
  assign n344 = n100 & n339;
  assign n345 = n93 & n289;
  assign n346 = n107 & n345;
  assign n347 = ~n344 & ~n346;
  assign n348 = n162 & n341;
  assign n349 = n100 & n341;
  assign n350 = ~n348 & ~n349;
  assign n351 = n347 & n350;
  assign n352 = n343 & n351;
  assign n353 = n143 & n341;
  assign n354 = n181 & n341;
  assign n355 = ~n353 & ~n354;
  assign n356 = n167 & n339;
  assign n357 = n176 & n339;
  assign n358 = ~n356 & ~n357;
  assign n359 = n355 & n358;
  assign n360 = n167 & n341;
  assign n361 = n181 & n339;
  assign n362 = ~n360 & ~n361;
  assign n363 = n165 & n339;
  assign n364 = n111 & n339;
  assign n365 = ~n363 & ~n364;
  assign n366 = n362 & n365;
  assign n367 = n359 & n366;
  assign n368 = n343 & n347;
  assign n369 = n358 & n368;
  assign n370 = n355 & n369;
  assign n371 = ~n364 & n370;
  assign n372 = ~n363 & n371;
  assign n373 = ~n361 & n372;
  assign n374 = ~n360 & n373;
  assign n375 = ~n349 & n374;
  assign n376 = ~n348 & n375;
  assign n377 = ~n349 & ~n364;
  assign n378 = n343 & n377;
  assign n379 = n347 & n378;
  assign n380 = ~n361 & ~n363;
  assign n381 = ~n348 & ~n360;
  assign n382 = n380 & n381;
  assign n383 = n359 & n382;
  assign n384 = n379 & n383;
  assign n385 = n343 & n362;
  assign n386 = n347 & n385;
  assign n387 = ~n348 & ~n364;
  assign n388 = ~n349 & ~n363;
  assign n389 = n387 & n388;
  assign n390 = n359 & n389;
  assign n391 = n386 & n390;
  assign n392 = n343 & n359;
  assign n393 = ~n349 & ~n361;
  assign n394 = ~n360 & ~n363;
  assign n395 = n393 & n394;
  assign n396 = n347 & n387;
  assign n397 = n395 & n396;
  assign n398 = n392 & n397;
  assign n399 = n352 & n367;
  assign n400 = n53443 & n289;
  assign n401 = n181 & n400;
  assign n402 = n173 & n400;
  assign n403 = ~n401 & ~n402;
  assign n404 = n162 & n400;
  assign n405 = n53446 & n400;
  assign n406 = ~n404 & ~n405;
  assign n407 = n403 & n406;
  assign n408 = n167 & n290;
  assign n409 = n176 & n341;
  assign n410 = n165 & n341;
  assign n411 = ~n409 & ~n410;
  assign n412 = ~n408 & n411;
  assign n413 = n407 & n412;
  assign n414 = n178 & n290;
  assign n415 = n100 & n290;
  assign n416 = n143 & n290;
  assign n417 = ~n415 & ~n416;
  assign n418 = ~n414 & n417;
  assign n419 = n162 & n339;
  assign n420 = n178 & n339;
  assign n421 = ~n419 & ~n420;
  assign n422 = n104 & n290;
  assign n423 = n53446 & n339;
  assign n424 = ~n422 & ~n423;
  assign n425 = n421 & n424;
  assign n426 = n418 & n425;
  assign n427 = ~n408 & ~n414;
  assign n428 = n424 & n427;
  assign n429 = ~n408 & n424;
  assign n430 = n418 & n429;
  assign n431 = n417 & n428;
  assign n432 = ~n409 & n421;
  assign n433 = ~n410 & n432;
  assign n434 = n411 & n421;
  assign n435 = n407 & n53466;
  assign n436 = n53465 & n435;
  assign n437 = n413 & n426;
  assign n438 = n53464 & n53467;
  assign n439 = n91 & n266;
  assign n440 = n111 & n439;
  assign n441 = n178 & n267;
  assign n442 = ~n440 & ~n441;
  assign n443 = n100 & n267;
  assign n444 = n178 & n341;
  assign n445 = ~n443 & ~n444;
  assign n446 = n442 & n445;
  assign n447 = n173 & n341;
  assign n448 = n143 & n345;
  assign n449 = ~n447 & ~n448;
  assign n450 = n183 & n341;
  assign n451 = n107 & n341;
  assign n452 = ~n450 & ~n451;
  assign n453 = n449 & n452;
  assign n454 = n445 & n452;
  assign n455 = n442 & n449;
  assign n456 = n454 & n455;
  assign n457 = n446 & n453;
  assign n458 = n266 & n289;
  assign n459 = n183 & n458;
  assign n460 = n173 & n439;
  assign n461 = n162 & n439;
  assign n462 = ~n460 & ~n461;
  assign n463 = ~n459 & n462;
  assign n464 = n176 & n290;
  assign n465 = n143 & n339;
  assign n466 = n104 & n339;
  assign n467 = ~n465 & ~n466;
  assign n468 = ~n464 & ~n465;
  assign n469 = ~n466 & n468;
  assign n470 = ~n464 & n467;
  assign n471 = n463 & n53469;
  assign n472 = ~n459 & ~n466;
  assign n473 = n445 & n472;
  assign n474 = n452 & n473;
  assign n475 = n462 & n474;
  assign n476 = ~n464 & n475;
  assign n477 = ~n441 & n476;
  assign n478 = ~n440 & n477;
  assign n479 = ~n465 & n478;
  assign n480 = ~n447 & n479;
  assign n481 = ~n448 & n480;
  assign n482 = n452 & n462;
  assign n483 = n445 & n482;
  assign n484 = ~n447 & ~n465;
  assign n485 = n442 & n484;
  assign n486 = ~n448 & ~n464;
  assign n487 = n472 & n486;
  assign n488 = n485 & n487;
  assign n489 = n483 & n488;
  assign n490 = n53468 & n471;
  assign n491 = n160 & n439;
  assign n492 = n139 & n266;
  assign n493 = n165 & n492;
  assign n494 = ~n491 & ~n493;
  assign n495 = n53446 & n492;
  assign n496 = n107 & n439;
  assign n497 = ~n495 & ~n496;
  assign n498 = n104 & n439;
  assign n499 = n178 & n439;
  assign n500 = ~n498 & ~n499;
  assign n501 = n497 & n500;
  assign n502 = n494 & n501;
  assign n503 = n181 & n439;
  assign n504 = n171 & n458;
  assign n505 = ~n503 & ~n504;
  assign n506 = n176 & n439;
  assign n507 = n143 & n439;
  assign n508 = ~n506 & ~n507;
  assign n509 = n505 & n508;
  assign n510 = n171 & n439;
  assign n511 = n53446 & n439;
  assign n512 = ~n510 & ~n511;
  assign n513 = n100 & n439;
  assign n514 = n107 & n458;
  assign n515 = ~n513 & ~n514;
  assign n516 = n512 & n515;
  assign n517 = n509 & n516;
  assign n518 = n497 & n512;
  assign n519 = n500 & n518;
  assign n520 = n494 & n519;
  assign n521 = ~n514 & n520;
  assign n522 = ~n504 & n521;
  assign n523 = ~n503 & n522;
  assign n524 = ~n513 & n523;
  assign n525 = ~n506 & n524;
  assign n526 = ~n507 & n525;
  assign n527 = ~n506 & ~n513;
  assign n528 = n494 & n512;
  assign n529 = n527 & n528;
  assign n530 = ~n504 & ~n507;
  assign n531 = ~n503 & ~n514;
  assign n532 = n530 & n531;
  assign n533 = n501 & n532;
  assign n534 = n529 & n533;
  assign n535 = n494 & n518;
  assign n536 = ~n504 & ~n506;
  assign n537 = ~n507 & ~n514;
  assign n538 = n536 & n537;
  assign n539 = ~n503 & ~n513;
  assign n540 = n500 & n539;
  assign n541 = n505 & n515;
  assign n542 = n500 & n508;
  assign n543 = n541 & n542;
  assign n544 = n538 & n540;
  assign n545 = n535 & n53472;
  assign n546 = n502 & n517;
  assign n547 = n53470 & n53471;
  assign n548 = n53467 & n53470;
  assign n549 = n53464 & n53471;
  assign n550 = n548 & n549;
  assign n551 = n438 & n547;
  assign n552 = n167 & n400;
  assign n553 = n111 & n400;
  assign n554 = n143 & n400;
  assign n555 = ~n553 & ~n554;
  assign n556 = ~n552 & ~n553;
  assign n557 = ~n554 & n556;
  assign n558 = ~n552 & n555;
  assign n559 = n97 & n165;
  assign n560 = n171 & n400;
  assign n561 = ~n559 & ~n560;
  assign n562 = n176 & n400;
  assign n563 = n561 & ~n562;
  assign n564 = n104 & n400;
  assign n565 = n183 & n400;
  assign n566 = ~n564 & ~n565;
  assign n567 = n97 & n53446;
  assign n568 = n107 & n400;
  assign n569 = ~n567 & ~n568;
  assign n570 = n566 & n569;
  assign n571 = ~n562 & ~n564;
  assign n572 = ~n562 & n566;
  assign n573 = ~n565 & n571;
  assign n574 = n561 & n569;
  assign n575 = n53475 & n574;
  assign n576 = n563 & n570;
  assign n577 = n53474 & n561;
  assign n578 = ~n567 & n577;
  assign n579 = ~n568 & n578;
  assign n580 = ~n565 & n579;
  assign n581 = ~n564 & n580;
  assign n582 = ~n562 & n581;
  assign n583 = n53474 & n53476;
  assign n584 = n178 & n400;
  assign n585 = n111 & n345;
  assign n586 = ~n584 & ~n585;
  assign n587 = n167 & n267;
  assign n588 = n183 & n345;
  assign n589 = ~n587 & ~n588;
  assign n590 = n171 & n345;
  assign n591 = n167 & n439;
  assign n592 = ~n590 & ~n591;
  assign n593 = n589 & n592;
  assign n594 = n586 & n593;
  assign n595 = ~n584 & ~n587;
  assign n596 = n53477 & ~n584;
  assign n597 = ~n587 & n596;
  assign n598 = n53477 & n595;
  assign n599 = ~n585 & ~n590;
  assign n600 = ~n588 & ~n591;
  assign n601 = n599 & n600;
  assign n602 = n53478 & n601;
  assign n603 = n586 & n589;
  assign n604 = n53477 & n603;
  assign n605 = ~n591 & n604;
  assign n606 = ~n590 & n605;
  assign n607 = ~n585 & n592;
  assign n608 = n589 & n607;
  assign n609 = n596 & n608;
  assign n610 = n53477 & n594;
  assign n611 = n165 & n439;
  assign n612 = n176 & n267;
  assign n613 = ~n611 & ~n612;
  assign n614 = n104 & n345;
  assign n615 = n160 & n339;
  assign n616 = ~n614 & ~n615;
  assign n617 = n183 & n439;
  assign n618 = n160 & n492;
  assign n619 = ~n617 & ~n618;
  assign n620 = n616 & n619;
  assign n621 = n613 & n620;
  assign n622 = n176 & n345;
  assign n623 = n167 & n345;
  assign n624 = ~n622 & ~n623;
  assign n625 = n178 & n345;
  assign n626 = n624 & ~n625;
  assign n627 = n111 & n341;
  assign n628 = n111 & n290;
  assign n629 = ~n627 & ~n628;
  assign n630 = n143 & n267;
  assign n631 = n173 & n290;
  assign n632 = ~n630 & ~n631;
  assign n633 = n629 & n632;
  assign n634 = n626 & n633;
  assign n635 = n616 & n629;
  assign n636 = n613 & n616;
  assign n637 = n629 & n636;
  assign n638 = n613 & n635;
  assign n639 = ~n617 & ~n630;
  assign n640 = ~n618 & ~n631;
  assign n641 = n619 & n632;
  assign n642 = n639 & n640;
  assign n643 = n626 & n53481;
  assign n644 = n53480 & n643;
  assign n645 = n621 & n634;
  assign n646 = n53446 & n341;
  assign n647 = n183 & n339;
  assign n648 = ~n646 & ~n647;
  assign n649 = n173 & n339;
  assign n650 = n160 & n341;
  assign n651 = n104 & n341;
  assign n652 = ~n650 & ~n651;
  assign n653 = ~n649 & n652;
  assign n654 = n648 & n652;
  assign n655 = ~n649 & n654;
  assign n656 = n648 & ~n649;
  assign n657 = n652 & n656;
  assign n658 = n648 & n653;
  assign n659 = n97 & n181;
  assign n660 = n100 & n400;
  assign n661 = ~n659 & ~n660;
  assign n662 = n97 & n160;
  assign n663 = n165 & n400;
  assign n664 = n160 & n400;
  assign n665 = ~n663 & ~n664;
  assign n666 = ~n662 & n665;
  assign n667 = ~n659 & ~n662;
  assign n668 = ~n660 & n667;
  assign n669 = ~n664 & n668;
  assign n670 = ~n663 & n669;
  assign n671 = ~n662 & ~n664;
  assign n672 = ~n660 & ~n663;
  assign n673 = ~n659 & n672;
  assign n674 = n671 & n673;
  assign n675 = ~n660 & ~n662;
  assign n676 = ~n659 & n665;
  assign n677 = n675 & n676;
  assign n678 = ~n660 & n665;
  assign n679 = n667 & n678;
  assign n680 = n661 & n666;
  assign n681 = n53483 & n53484;
  assign n682 = n626 & n53483;
  assign n683 = n629 & n682;
  assign n684 = n613 & n683;
  assign n685 = n53484 & n684;
  assign n686 = ~n631 & n685;
  assign n687 = ~n618 & n686;
  assign n688 = ~n630 & n687;
  assign n689 = ~n617 & n688;
  assign n690 = ~n615 & n689;
  assign n691 = ~n614 & n690;
  assign n692 = n53482 & n681;
  assign n693 = n53479 & n53485;
  assign n694 = n53473 & n53485;
  assign n695 = n53479 & n694;
  assign n696 = n53473 & n693;
  assign n697 = n435 & n53485;
  assign n698 = n53470 & n697;
  assign n699 = n53463 & n698;
  assign n700 = n53479 & n699;
  assign n701 = n53471 & n700;
  assign n702 = n53464 & n701;
  assign n703 = n417 & n702;
  assign n704 = n424 & n703;
  assign n705 = ~n414 & n704;
  assign n706 = ~n408 & n705;
  assign n707 = n53463 & n53486;
  assign n708 = ~n444 & ~n465;
  assign n709 = n421 & n708;
  assign n710 = n53466 & n708;
  assign n711 = n411 & n709;
  assign n712 = ~n447 & ~n627;
  assign n713 = ~n466 & ~n615;
  assign n714 = ~n466 & n712;
  assign n715 = ~n615 & n714;
  assign n716 = n712 & n713;
  assign n717 = ~n423 & n452;
  assign n718 = n53489 & n717;
  assign n719 = ~n423 & ~n465;
  assign n720 = ~n444 & n719;
  assign n721 = n708 & n717;
  assign n722 = n452 & n720;
  assign n723 = n53466 & n53489;
  assign n724 = n53490 & n723;
  assign n725 = n53488 & n718;
  assign n726 = n53466 & n53483;
  assign n727 = n53489 & n726;
  assign n728 = n452 & n727;
  assign n729 = ~n423 & n728;
  assign n730 = ~n465 & n729;
  assign n731 = ~n444 & n730;
  assign n732 = n53483 & n53491;
  assign n733 = n107 & n339;
  assign n734 = n93 & n209;
  assign n735 = n173 & n734;
  assign n736 = ~n733 & ~n735;
  assign n737 = n53492 & ~n733;
  assign n738 = ~n735 & n737;
  assign n739 = n53492 & n736;
  assign n740 = n107 & n734;
  assign n741 = n176 & n734;
  assign n742 = n53446 & n458;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~n740 & ~n741;
  assign n745 = ~n742 & n744;
  assign n746 = ~n740 & n743;
  assign n747 = n183 & n734;
  assign n748 = n160 & n458;
  assign n749 = ~n747 & ~n748;
  assign n750 = n100 & n734;
  assign n751 = n111 & n734;
  assign n752 = ~n750 & ~n751;
  assign n753 = n53446 & n734;
  assign n754 = n167 & n734;
  assign n755 = ~n753 & ~n754;
  assign n756 = n752 & n755;
  assign n757 = n749 & n755;
  assign n758 = n752 & n757;
  assign n759 = n749 & n756;
  assign n760 = ~n742 & n757;
  assign n761 = ~n740 & n760;
  assign n762 = ~n741 & n761;
  assign n763 = ~n751 & n762;
  assign n764 = ~n750 & n763;
  assign n765 = ~n740 & n752;
  assign n766 = n743 & n749;
  assign n767 = n755 & n766;
  assign n768 = n765 & n767;
  assign n769 = n53494 & n53495;
  assign n770 = n181 & n734;
  assign n771 = n162 & n734;
  assign n772 = ~n770 & ~n771;
  assign n773 = n143 & n734;
  assign n774 = n104 & n734;
  assign n775 = ~n773 & ~n774;
  assign n776 = n178 & n734;
  assign n777 = n165 & n734;
  assign n778 = ~n776 & ~n777;
  assign n779 = n775 & n778;
  assign n780 = n772 & n778;
  assign n781 = n775 & n780;
  assign n782 = n772 & n779;
  assign n783 = n53496 & n775;
  assign n784 = n772 & n783;
  assign n785 = ~n776 & n784;
  assign n786 = ~n777 & n785;
  assign n787 = n53496 & n53497;
  assign n788 = n160 & n734;
  assign n789 = n171 & n734;
  assign n790 = ~n788 & ~n789;
  assign n791 = n53464 & n790;
  assign n792 = n53498 & n791;
  assign n793 = n53493 & n53498;
  assign n794 = n53464 & n793;
  assign n795 = ~n788 & n794;
  assign n796 = ~n789 & n795;
  assign n797 = n53493 & n792;
  assign n798 = ~n441 & ~n612;
  assign n799 = ~n448 & ~n614;
  assign n800 = ~n319 & n799;
  assign n801 = n798 & n800;
  assign n802 = n276 & ~n630;
  assign n803 = n626 & n802;
  assign n804 = ~n630 & n798;
  assign n805 = n276 & n804;
  assign n806 = n626 & n799;
  assign n807 = ~n319 & n806;
  assign n808 = n805 & n807;
  assign n809 = n626 & n798;
  assign n810 = n802 & n809;
  assign n811 = n799 & n810;
  assign n812 = ~n319 & n811;
  assign n813 = n801 & n803;
  assign n814 = ~n585 & ~n588;
  assign n815 = ~n268 & ~n590;
  assign n816 = ~n590 & n814;
  assign n817 = ~n588 & n599;
  assign n818 = ~n268 & n53501;
  assign n819 = ~n268 & n814;
  assign n820 = ~n590 & n819;
  assign n821 = n814 & n815;
  assign n822 = n176 & n458;
  assign n823 = n162 & n458;
  assign n824 = n143 & n458;
  assign n825 = ~n823 & ~n824;
  assign n826 = ~n822 & ~n823;
  assign n827 = ~n824 & n826;
  assign n828 = ~n822 & n825;
  assign n829 = n173 & n458;
  assign n830 = n181 & n458;
  assign n831 = ~n829 & ~n830;
  assign n832 = n167 & n458;
  assign n833 = n178 & n458;
  assign n834 = ~n832 & ~n833;
  assign n835 = n831 & n834;
  assign n836 = ~n823 & n831;
  assign n837 = ~n833 & n836;
  assign n838 = ~n824 & n837;
  assign n839 = ~n832 & n838;
  assign n840 = ~n822 & n839;
  assign n841 = ~n823 & n834;
  assign n842 = ~n822 & ~n824;
  assign n843 = n831 & n842;
  assign n844 = n841 & n843;
  assign n845 = n53503 & n835;
  assign n846 = ~n269 & ~n443;
  assign n847 = ~n587 & n846;
  assign n848 = n104 & n458;
  assign n849 = n111 & n458;
  assign n850 = ~n848 & ~n849;
  assign n851 = n100 & n458;
  assign n852 = n165 & n458;
  assign n853 = ~n851 & ~n852;
  assign n854 = n850 & n853;
  assign n855 = ~n587 & ~n852;
  assign n856 = ~n851 & n855;
  assign n857 = ~n587 & n853;
  assign n858 = n846 & n850;
  assign n859 = n53505 & n858;
  assign n860 = n847 & n854;
  assign n861 = n53504 & n53506;
  assign n862 = n53502 & n53506;
  assign n863 = n53504 & n862;
  assign n864 = n53502 & n861;
  assign n865 = n53500 & n53507;
  assign n866 = n53500 & n53502;
  assign n867 = n53499 & n866;
  assign n868 = n53504 & n867;
  assign n869 = n846 & n868;
  assign n870 = n850 & n869;
  assign n871 = ~n852 & n870;
  assign n872 = ~n851 & n871;
  assign n873 = ~n587 & n872;
  assign n874 = n53499 & n865;
  assign n875 = n53487 & ~n53508;
  assign n876 = ~n53487 & n53508;
  assign n877 = ~n875 & ~n876;
  assign n878 = n92 & n209;
  assign n879 = n178 & n878;
  assign n880 = n91 & n92;
  assign n881 = n181 & n880;
  assign n882 = ~n879 & ~n881;
  assign n883 = n165 & n880;
  assign n884 = ~n511 & ~n590;
  assign n885 = ~n590 & ~n883;
  assign n886 = ~n511 & n885;
  assign n887 = ~n511 & ~n883;
  assign n888 = ~n590 & n887;
  assign n889 = ~n883 & n884;
  assign n890 = n882 & ~n883;
  assign n891 = ~n511 & n890;
  assign n892 = ~n590 & n891;
  assign n893 = n882 & n53509;
  assign n894 = n107 & n290;
  assign n895 = ~n255 & ~n894;
  assign n896 = n183 & n290;
  assign n897 = ~n211 & ~n896;
  assign n898 = ~n272 & ~n459;
  assign n899 = n897 & n898;
  assign n900 = n895 & n899;
  assign n901 = n165 & n878;
  assign n902 = n100 & n880;
  assign n903 = ~n901 & ~n902;
  assign n904 = n406 & n903;
  assign n905 = ~n650 & ~n742;
  assign n906 = ~n733 & ~n852;
  assign n907 = n905 & n906;
  assign n908 = n904 & n907;
  assign n909 = n900 & n908;
  assign n910 = n53510 & n909;
  assign n911 = n162 & n492;
  assign n912 = ~n222 & ~n911;
  assign n913 = n217 & n912;
  assign n914 = n173 & n492;
  assign n915 = ~n259 & ~n914;
  assign n916 = ~n256 & ~n510;
  assign n917 = n915 & n916;
  assign n918 = n217 & n915;
  assign n919 = n912 & n916;
  assign n920 = n918 & n919;
  assign n921 = n913 & n917;
  assign n922 = n143 & n880;
  assign n923 = ~n269 & ~n588;
  assign n924 = ~n269 & ~n922;
  assign n925 = ~n588 & n924;
  assign n926 = ~n922 & n923;
  assign n927 = ~n249 & ~n342;
  assign n928 = ~n753 & ~n770;
  assign n929 = n927 & n928;
  assign n930 = n53512 & n929;
  assign n931 = n916 & n53512;
  assign n932 = n915 & n931;
  assign n933 = n217 & n932;
  assign n934 = ~n222 & n933;
  assign n935 = ~n249 & n934;
  assign n936 = ~n911 & n935;
  assign n937 = ~n342 & n936;
  assign n938 = ~n770 & n937;
  assign n939 = ~n753 & n938;
  assign n940 = ~n249 & ~n753;
  assign n941 = n217 & n940;
  assign n942 = n917 & n941;
  assign n943 = ~n342 & ~n770;
  assign n944 = n912 & n943;
  assign n945 = n53512 & n944;
  assign n946 = n942 & n945;
  assign n947 = n53511 & n930;
  assign n948 = n176 & n880;
  assign n949 = ~n258 & ~n552;
  assign n950 = ~n258 & ~n948;
  assign n951 = ~n552 & n950;
  assign n952 = ~n552 & ~n948;
  assign n953 = ~n258 & n952;
  assign n954 = ~n948 & n949;
  assign n955 = ~n207 & ~n491;
  assign n956 = n183 & n492;
  assign n957 = n100 & n878;
  assign n958 = ~n956 & ~n957;
  assign n959 = ~n491 & ~n957;
  assign n960 = ~n207 & ~n956;
  assign n961 = n959 & n960;
  assign n962 = n955 & n958;
  assign n963 = ~n443 & ~n615;
  assign n964 = ~n206 & ~n250;
  assign n965 = n963 & n964;
  assign n966 = n53515 & n965;
  assign n967 = n53514 & n964;
  assign n968 = ~n957 & n967;
  assign n969 = ~n207 & n968;
  assign n970 = ~n956 & n969;
  assign n971 = ~n443 & n970;
  assign n972 = ~n491 & n971;
  assign n973 = ~n615 & n972;
  assign n974 = n53514 & n966;
  assign n975 = n53446 & n267;
  assign n976 = ~n611 & ~n975;
  assign n977 = n167 & n878;
  assign n978 = ~n823 & ~n977;
  assign n979 = n976 & ~n977;
  assign n980 = ~n823 & n979;
  assign n981 = n976 & n978;
  assign n982 = ~n410 & ~n646;
  assign n983 = n173 & n878;
  assign n984 = n171 & n880;
  assign n985 = ~n983 & ~n984;
  assign n986 = n982 & n985;
  assign n987 = n53517 & n986;
  assign n988 = ~n308 & ~n363;
  assign n989 = ~n308 & ~n419;
  assign n990 = ~n363 & n989;
  assign n991 = ~n363 & ~n419;
  assign n992 = ~n308 & n991;
  assign n993 = ~n419 & n988;
  assign n994 = ~n499 & ~n584;
  assign n995 = ~n441 & ~n584;
  assign n996 = ~n440 & n995;
  assign n997 = ~n499 & n996;
  assign n998 = ~n440 & ~n499;
  assign n999 = n995 & n998;
  assign n1000 = n442 & n994;
  assign n1001 = n53518 & n53519;
  assign n1002 = n987 & n1001;
  assign n1003 = n53516 & n1002;
  assign n1004 = n53513 & n1003;
  assign n1005 = n903 & n906;
  assign n1006 = n897 & n1005;
  assign n1007 = ~n646 & ~n894;
  assign n1008 = n898 & n1007;
  assign n1009 = n406 & n905;
  assign n1010 = n1008 & n1009;
  assign n1011 = n903 & n905;
  assign n1012 = n898 & n1011;
  assign n1013 = n897 & n1007;
  assign n1014 = n406 & n906;
  assign n1015 = n1013 & n1014;
  assign n1016 = n1012 & n1015;
  assign n1017 = n1006 & n1010;
  assign n1018 = n53510 & n53520;
  assign n1019 = ~n255 & ~n984;
  assign n1020 = ~n410 & ~n983;
  assign n1021 = ~n255 & ~n983;
  assign n1022 = ~n410 & ~n984;
  assign n1023 = n1021 & n1022;
  assign n1024 = n1019 & n1020;
  assign n1025 = n53517 & n53521;
  assign n1026 = n1001 & n1025;
  assign n1027 = n53516 & n1026;
  assign n1028 = n53513 & n1027;
  assign n1029 = n1018 & n1028;
  assign n1030 = n910 & n1004;
  assign n1031 = n160 & n880;
  assign n1032 = ~n649 & ~n1031;
  assign n1033 = n111 & n880;
  assign n1034 = n107 & n492;
  assign n1035 = ~n777 & ~n1034;
  assign n1036 = ~n1033 & n1035;
  assign n1037 = n1032 & n1035;
  assign n1038 = ~n1033 & n1037;
  assign n1039 = n1032 & ~n1033;
  assign n1040 = n1035 & n1039;
  assign n1041 = n1032 & n1036;
  assign n1042 = n100 & n492;
  assign n1043 = ~n587 & ~n1042;
  assign n1044 = n104 & n880;
  assign n1045 = ~n361 & ~n1044;
  assign n1046 = n403 & n1045;
  assign n1047 = n403 & ~n1044;
  assign n1048 = ~n1042 & n1047;
  assign n1049 = ~n587 & n1048;
  assign n1050 = ~n361 & n1049;
  assign n1051 = ~n361 & ~n587;
  assign n1052 = ~n1042 & ~n1044;
  assign n1053 = ~n361 & ~n1042;
  assign n1054 = ~n587 & ~n1044;
  assign n1055 = n1053 & n1054;
  assign n1056 = n1051 & n1052;
  assign n1057 = n403 & n53525;
  assign n1058 = n1043 & n1046;
  assign n1059 = n171 & n492;
  assign n1060 = ~n504 & ~n1059;
  assign n1061 = n160 & n878;
  assign n1062 = n181 & n878;
  assign n1063 = ~n1061 & ~n1062;
  assign n1064 = n1060 & n1063;
  assign n1065 = n167 & n880;
  assign n1066 = ~n247 & ~n1065;
  assign n1067 = ~n271 & ~n317;
  assign n1068 = n1066 & n1067;
  assign n1069 = n1060 & n1066;
  assign n1070 = n1063 & n1067;
  assign n1071 = n1069 & n1070;
  assign n1072 = n1064 & n1068;
  assign n1073 = n53524 & n53526;
  assign n1074 = n53523 & n1073;
  assign n1075 = ~n660 & ~n740;
  assign n1076 = ~n614 & ~n664;
  assign n1077 = n1075 & n1076;
  assign n1078 = ~n218 & ~n750;
  assign n1079 = n53446 & n878;
  assign n1080 = n92 & n139;
  assign n1081 = n107 & n1080;
  assign n1082 = ~n1079 & ~n1081;
  assign n1083 = n1078 & n1082;
  assign n1084 = n1077 & n1083;
  assign n1085 = n53446 & n880;
  assign n1086 = ~n246 & ~n554;
  assign n1087 = ~n1085 & n1086;
  assign n1088 = n173 & n880;
  assign n1089 = ~n268 & ~n1088;
  assign n1090 = n171 & n290;
  assign n1091 = ~n829 & ~n1090;
  assign n1092 = n1089 & n1091;
  assign n1093 = n1087 & n1092;
  assign n1094 = ~n1085 & ~n1088;
  assign n1095 = n1078 & n1094;
  assign n1096 = n1076 & n1082;
  assign n1097 = n1094 & n1096;
  assign n1098 = n1078 & n1097;
  assign n1099 = n1095 & n1096;
  assign n1100 = n1091 & n53527;
  assign n1101 = ~n246 & n1100;
  assign n1102 = ~n660 & n1101;
  assign n1103 = ~n554 & n1102;
  assign n1104 = ~n268 & n1103;
  assign n1105 = ~n740 & n1104;
  assign n1106 = n1075 & n1078;
  assign n1107 = n1082 & n1091;
  assign n1108 = n1106 & n1107;
  assign n1109 = ~n246 & ~n268;
  assign n1110 = ~n554 & n1109;
  assign n1111 = ~n268 & n1086;
  assign n1112 = n1076 & n1094;
  assign n1113 = n53529 & n1112;
  assign n1114 = n1108 & n1113;
  assign n1115 = ~n554 & n1075;
  assign n1116 = n1091 & n1109;
  assign n1117 = n1115 & n1116;
  assign n1118 = n53527 & n1117;
  assign n1119 = n1084 & n1093;
  assign n1120 = ~n498 & ~n514;
  assign n1121 = ~n748 & n1120;
  assign n1122 = ~n585 & ~n630;
  assign n1123 = n452 & n1122;
  assign n1124 = n178 & n880;
  assign n1125 = n162 & n880;
  assign n1126 = ~n1124 & ~n1125;
  assign n1127 = n143 & n878;
  assign n1128 = ~n448 & ~n1127;
  assign n1129 = n1126 & n1128;
  assign n1130 = n1123 & n1129;
  assign n1131 = ~n748 & n1122;
  assign n1132 = n452 & n1120;
  assign n1133 = n1129 & n1132;
  assign n1134 = n1131 & n1133;
  assign n1135 = n1121 & n1130;
  assign n1136 = n53528 & n53530;
  assign n1137 = n53523 & n1060;
  assign n1138 = n53524 & n1137;
  assign n1139 = n452 & n1138;
  assign n1140 = n53528 & n1139;
  assign n1141 = n1067 & n1140;
  assign n1142 = n1128 & n1141;
  assign n1143 = ~n1124 & n1142;
  assign n1144 = ~n1125 & n1143;
  assign n1145 = ~n1065 & n1144;
  assign n1146 = ~n1062 & n1145;
  assign n1147 = ~n1061 & n1146;
  assign n1148 = ~n247 & n1147;
  assign n1149 = ~n514 & n1148;
  assign n1150 = ~n748 & n1149;
  assign n1151 = ~n630 & n1150;
  assign n1152 = ~n498 & n1151;
  assign n1153 = ~n585 & n1152;
  assign n1154 = n1060 & n1128;
  assign n1155 = n1068 & n1154;
  assign n1156 = n53524 & n1155;
  assign n1157 = n53523 & n1156;
  assign n1158 = ~n514 & ~n585;
  assign n1159 = ~n748 & n1158;
  assign n1160 = ~n498 & ~n630;
  assign n1161 = n1063 & n1160;
  assign n1162 = n452 & n1126;
  assign n1163 = n1161 & n1162;
  assign n1164 = n1159 & n1163;
  assign n1165 = n53528 & n1164;
  assign n1166 = n1157 & n1165;
  assign n1167 = n1060 & n1067;
  assign n1168 = n452 & n1128;
  assign n1169 = n1167 & n1168;
  assign n1170 = n53524 & n1169;
  assign n1171 = n53523 & n1170;
  assign n1172 = ~n498 & ~n585;
  assign n1173 = ~n247 & n1172;
  assign n1174 = ~n1061 & ~n1065;
  assign n1175 = ~n514 & ~n748;
  assign n1176 = n1174 & n1175;
  assign n1177 = ~n630 & ~n1062;
  assign n1178 = n1126 & n1177;
  assign n1179 = n1176 & n1178;
  assign n1180 = n1173 & n1179;
  assign n1181 = n53528 & n1180;
  assign n1182 = n1171 & n1181;
  assign n1183 = n1074 & n1136;
  assign n1184 = ~n423 & ~n788;
  assign n1185 = ~n219 & ~n663;
  assign n1186 = ~n212 & ~n771;
  assign n1187 = n1185 & n1186;
  assign n1188 = n1184 & n1187;
  assign n1189 = n143 & n492;
  assign n1190 = ~n506 & ~n1189;
  assign n1191 = n176 & n878;
  assign n1192 = n162 & n878;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = n1190 & n1193;
  assign n1195 = n171 & n1080;
  assign n1196 = n183 & n1080;
  assign n1197 = ~n1195 & ~n1196;
  assign n1198 = ~n221 & ~n346;
  assign n1199 = n1197 & n1198;
  assign n1200 = ~n221 & ~n1192;
  assign n1201 = ~n1189 & ~n1191;
  assign n1202 = ~n221 & ~n1189;
  assign n1203 = n1193 & n1202;
  assign n1204 = n1200 & n1201;
  assign n1205 = ~n346 & ~n506;
  assign n1206 = n1197 & n1205;
  assign n1207 = n53532 & n1206;
  assign n1208 = n1201 & n1205;
  assign n1209 = n1197 & n1200;
  assign n1210 = n1208 & n1209;
  assign n1211 = n1194 & n1199;
  assign n1212 = n626 & n53533;
  assign n1213 = n626 & n1186;
  assign n1214 = n1197 & n1213;
  assign n1215 = ~n1192 & n1214;
  assign n1216 = ~n1191 & n1215;
  assign n1217 = ~n219 & n1216;
  assign n1218 = ~n221 & n1217;
  assign n1219 = ~n663 & n1218;
  assign n1220 = ~n1189 & n1219;
  assign n1221 = ~n506 & n1220;
  assign n1222 = ~n423 & n1221;
  assign n1223 = ~n788 & n1222;
  assign n1224 = ~n346 & n1223;
  assign n1225 = n1184 & n1186;
  assign n1226 = n1197 & n1225;
  assign n1227 = ~n219 & ~n506;
  assign n1228 = ~n346 & ~n663;
  assign n1229 = n1227 & n1228;
  assign n1230 = n53532 & n1229;
  assign n1231 = n626 & n1230;
  assign n1232 = n1226 & n1231;
  assign n1233 = n1188 & n1212;
  assign n1234 = n181 & n492;
  assign n1235 = ~n830 & ~n1234;
  assign n1236 = ~n735 & ~n1234;
  assign n1237 = ~n830 & n1236;
  assign n1238 = ~n735 & n1235;
  assign n1239 = n53534 & ~n1234;
  assign n1240 = ~n830 & n1239;
  assign n1241 = ~n735 & n1240;
  assign n1242 = n53534 & n53535;
  assign n1243 = n53531 & n53536;
  assign n1244 = n897 & n53517;
  assign n1245 = n53536 & n1244;
  assign n1246 = n53510 & n1245;
  assign n1247 = n53531 & n1246;
  assign n1248 = n53513 & n1247;
  assign n1249 = n53519 & n1248;
  assign n1250 = n53518 & n1249;
  assign n1251 = n906 & n1250;
  assign n1252 = n53516 & n1251;
  assign n1253 = n905 & n1252;
  assign n1254 = n903 & n1253;
  assign n1255 = n406 & n1254;
  assign n1256 = ~n984 & n1255;
  assign n1257 = ~n894 & n1256;
  assign n1258 = ~n983 & n1257;
  assign n1259 = ~n255 & n1258;
  assign n1260 = ~n272 & n1259;
  assign n1261 = ~n459 & n1260;
  assign n1262 = ~n646 & n1261;
  assign n1263 = ~n410 & n1262;
  assign n1264 = n53522 & n1243;
  assign n1265 = ~n491 & ~n984;
  assign n1266 = ~n348 & ~n774;
  assign n1267 = ~n353 & ~n514;
  assign n1268 = n1266 & n1267;
  assign n1269 = n1265 & n1268;
  assign n1270 = ~n444 & ~n627;
  assign n1271 = ~n410 & ~n511;
  assign n1272 = n1270 & n1271;
  assign n1273 = ~n1044 & ~n1189;
  assign n1274 = ~n460 & ~n664;
  assign n1275 = n1273 & n1274;
  assign n1276 = n1272 & n1275;
  assign n1277 = ~n735 & ~n770;
  assign n1278 = ~n360 & ~n771;
  assign n1279 = n1277 & n1278;
  assign n1280 = n178 & n492;
  assign n1281 = ~n750 & ~n1280;
  assign n1282 = ~n894 & ~n1090;
  assign n1283 = n1281 & n1282;
  assign n1284 = n1279 & n1283;
  assign n1285 = n1276 & n1284;
  assign n1286 = n1269 & n1273;
  assign n1287 = n1277 & n1286;
  assign n1288 = n1278 & n1287;
  assign n1289 = ~n1090 & n1288;
  assign n1290 = ~n894 & n1289;
  assign n1291 = ~n664 & n1290;
  assign n1292 = ~n1280 & n1291;
  assign n1293 = ~n511 & n1292;
  assign n1294 = ~n460 & n1293;
  assign n1295 = ~n627 & n1294;
  assign n1296 = ~n410 & n1295;
  assign n1297 = ~n444 & n1296;
  assign n1298 = ~n750 & n1297;
  assign n1299 = n1265 & n1273;
  assign n1300 = n1266 & n1299;
  assign n1301 = ~n410 & ~n627;
  assign n1302 = ~n511 & ~n664;
  assign n1303 = n1301 & n1302;
  assign n1304 = ~n444 & ~n460;
  assign n1305 = n1267 & n1304;
  assign n1306 = n1303 & n1305;
  assign n1307 = n1284 & n1306;
  assign n1308 = n1300 & n1307;
  assign n1309 = n1267 & n1273;
  assign n1310 = n1265 & n1309;
  assign n1311 = ~n444 & ~n1090;
  assign n1312 = ~n511 & ~n1280;
  assign n1313 = n1311 & n1312;
  assign n1314 = ~n750 & ~n894;
  assign n1315 = n1266 & n1314;
  assign n1316 = n1313 & n1315;
  assign n1317 = n1274 & n1301;
  assign n1318 = n1279 & n1317;
  assign n1319 = n1316 & n1318;
  assign n1320 = n1310 & n1319;
  assign n1321 = n1268 & n1278;
  assign n1322 = ~n1090 & ~n1280;
  assign n1323 = n1265 & n1322;
  assign n1324 = n1273 & n1277;
  assign n1325 = n1323 & n1324;
  assign n1326 = ~n460 & ~n511;
  assign n1327 = ~n410 & ~n444;
  assign n1328 = n1326 & n1327;
  assign n1329 = ~n627 & ~n894;
  assign n1330 = ~n664 & ~n750;
  assign n1331 = n1329 & n1330;
  assign n1332 = n1328 & n1331;
  assign n1333 = n1325 & n1332;
  assign n1334 = n1321 & n1333;
  assign n1335 = n1269 & n1285;
  assign n1336 = ~n503 & ~n773;
  assign n1337 = n167 & n492;
  assign n1338 = ~n507 & ~n1337;
  assign n1339 = ~n1065 & ~n1337;
  assign n1340 = ~n507 & n1339;
  assign n1341 = ~n1065 & n1338;
  assign n1342 = ~n503 & n1339;
  assign n1343 = ~n507 & n1342;
  assign n1344 = ~n773 & n1343;
  assign n1345 = n1336 & n53539;
  assign n1346 = ~n741 & ~n754;
  assign n1347 = ~n459 & ~n776;
  assign n1348 = ~n914 & ~n1033;
  assign n1349 = ~n776 & ~n914;
  assign n1350 = ~n459 & ~n1033;
  assign n1351 = n1349 & n1350;
  assign n1352 = n1347 & n1348;
  assign n1353 = ~n1033 & n1346;
  assign n1354 = ~n914 & n1353;
  assign n1355 = ~n459 & n1354;
  assign n1356 = ~n776 & n1355;
  assign n1357 = n1346 & n53541;
  assign n1358 = ~n354 & ~n663;
  assign n1359 = n652 & n1358;
  assign n1360 = ~n447 & ~n902;
  assign n1361 = ~n611 & ~n789;
  assign n1362 = n1360 & n1361;
  assign n1363 = n1359 & n1362;
  assign n1364 = n53542 & n1363;
  assign n1365 = n53540 & n1364;
  assign n1366 = ~n922 & ~n1031;
  assign n1367 = ~n948 & n1366;
  assign n1368 = ~n883 & ~n896;
  assign n1369 = n1126 & n1368;
  assign n1370 = ~n1031 & ~n1124;
  assign n1371 = ~n1125 & n1370;
  assign n1372 = ~n948 & n1371;
  assign n1373 = ~n922 & n1372;
  assign n1374 = ~n883 & n1373;
  assign n1375 = ~n896 & n1374;
  assign n1376 = ~n883 & ~n948;
  assign n1377 = ~n948 & n1368;
  assign n1378 = ~n896 & n1376;
  assign n1379 = n1126 & n1366;
  assign n1380 = n53544 & n1379;
  assign n1381 = ~n883 & ~n1031;
  assign n1382 = ~n922 & n1381;
  assign n1383 = ~n896 & ~n948;
  assign n1384 = n1126 & n1383;
  assign n1385 = n1382 & n1384;
  assign n1386 = n1367 & n1369;
  assign n1387 = ~n881 & n1094;
  assign n1388 = n1094 & n53543;
  assign n1389 = ~n881 & n1388;
  assign n1390 = n53543 & n1387;
  assign n1391 = ~n513 & ~n660;
  assign n1392 = ~n349 & ~n409;
  assign n1393 = ~n409 & n1391;
  assign n1394 = ~n349 & n1393;
  assign n1395 = n1391 & n1392;
  assign n1396 = ~n461 & ~n751;
  assign n1397 = ~n1042 & n1396;
  assign n1398 = n407 & n1397;
  assign n1399 = n53546 & n1398;
  assign n1400 = n53545 & n1399;
  assign n1401 = ~n354 & ~n461;
  assign n1402 = n652 & n1401;
  assign n1403 = n1362 & n1402;
  assign n1404 = n53540 & n1403;
  assign n1405 = n53542 & n1404;
  assign n1406 = ~n663 & ~n751;
  assign n1407 = ~n1042 & n1406;
  assign n1408 = n407 & n1407;
  assign n1409 = n53546 & n1408;
  assign n1410 = n53545 & n1409;
  assign n1411 = n1405 & n1410;
  assign n1412 = ~n663 & ~n1042;
  assign n1413 = n1396 & n1412;
  assign n1414 = n652 & n1360;
  assign n1415 = n1413 & n1414;
  assign n1416 = n53542 & n1415;
  assign n1417 = n53540 & n1416;
  assign n1418 = ~n354 & ~n789;
  assign n1419 = ~n611 & n1418;
  assign n1420 = n53546 & n1419;
  assign n1421 = n407 & n1420;
  assign n1422 = n53545 & n1421;
  assign n1423 = n1417 & n1422;
  assign n1424 = ~n751 & ~n902;
  assign n1425 = ~n789 & ~n1042;
  assign n1426 = n1424 & n1425;
  assign n1427 = ~n447 & ~n611;
  assign n1428 = n652 & n1427;
  assign n1429 = n1426 & n1428;
  assign n1430 = n53542 & n1429;
  assign n1431 = n53540 & n1430;
  assign n1432 = ~n461 & ~n663;
  assign n1433 = ~n354 & n1432;
  assign n1434 = n53546 & n1433;
  assign n1435 = n407 & n1434;
  assign n1436 = n53545 & n1435;
  assign n1437 = n1431 & n1436;
  assign n1438 = n1365 & n1400;
  assign n1439 = n53545 & n53546;
  assign n1440 = n407 & n1439;
  assign n1441 = n652 & n1440;
  assign n1442 = n53540 & n1441;
  assign n1443 = n53538 & n1442;
  assign n1444 = n53542 & n1443;
  assign n1445 = ~n902 & n1444;
  assign n1446 = ~n663 & n1445;
  assign n1447 = ~n1042 & n1446;
  assign n1448 = ~n611 & n1447;
  assign n1449 = ~n461 & n1448;
  assign n1450 = ~n354 & n1449;
  assign n1451 = ~n447 & n1450;
  assign n1452 = ~n751 & n1451;
  assign n1453 = ~n789 & n1452;
  assign n1454 = n53538 & n53547;
  assign n1455 = n111 & n492;
  assign n1456 = ~n733 & ~n1455;
  assign n1457 = n176 & n492;
  assign n1458 = ~n788 & ~n1457;
  assign n1459 = ~n504 & n1458;
  assign n1460 = n1456 & n1459;
  assign n1461 = n53548 & n1456;
  assign n1462 = n1458 & n1461;
  assign n1463 = ~n504 & n1462;
  assign n1464 = n53548 & n1460;
  assign n1465 = n176 & n1080;
  assign n1466 = n178 & n1080;
  assign n1467 = ~n1465 & ~n1466;
  assign n1468 = n100 & n1080;
  assign n1469 = n173 & n1080;
  assign n1470 = ~n1468 & ~n1469;
  assign n1471 = n183 & n880;
  assign n1472 = n162 & n1080;
  assign n1473 = ~n1471 & ~n1472;
  assign n1474 = n1470 & n1473;
  assign n1475 = n1467 & n1474;
  assign n1476 = n165 & n1080;
  assign n1477 = n111 & n1080;
  assign n1478 = n104 & n1080;
  assign n1479 = ~n1477 & ~n1478;
  assign n1480 = ~n1476 & ~n1478;
  assign n1481 = ~n1477 & n1480;
  assign n1482 = ~n1476 & ~n1477;
  assign n1483 = ~n1478 & n1482;
  assign n1484 = ~n1476 & n1479;
  assign n1485 = n160 & n1080;
  assign n1486 = n107 & n880;
  assign n1487 = n167 & n1080;
  assign n1488 = ~n1486 & ~n1487;
  assign n1489 = ~n1485 & n1488;
  assign n1490 = n53446 & n1080;
  assign n1491 = n143 & n1080;
  assign n1492 = n181 & n1080;
  assign n1493 = ~n1491 & ~n1492;
  assign n1494 = ~n1490 & ~n1491;
  assign n1495 = ~n1492 & n1494;
  assign n1496 = ~n1490 & n1493;
  assign n1497 = n1489 & n53551;
  assign n1498 = n53550 & n1497;
  assign n1499 = n53550 & n53551;
  assign n1500 = n1467 & n1499;
  assign n1501 = n1488 & n1500;
  assign n1502 = ~n1471 & n1501;
  assign n1503 = ~n1472 & n1502;
  assign n1504 = ~n1469 & n1503;
  assign n1505 = ~n1485 & n1504;
  assign n1506 = ~n1468 & n1505;
  assign n1507 = ~n1468 & ~n1471;
  assign n1508 = n1488 & n1507;
  assign n1509 = n1467 & n1508;
  assign n1510 = ~n1472 & ~n1485;
  assign n1511 = ~n1469 & n1510;
  assign n1512 = n53550 & n1511;
  assign n1513 = n53551 & n1512;
  assign n1514 = n1509 & n1513;
  assign n1515 = ~n1469 & ~n1471;
  assign n1516 = n1488 & n1515;
  assign n1517 = n1467 & n1515;
  assign n1518 = n1488 & n1517;
  assign n1519 = n1467 & n1516;
  assign n1520 = ~n1468 & ~n1472;
  assign n1521 = ~n1485 & n1520;
  assign n1522 = ~n1468 & n1510;
  assign n1523 = n53551 & n53554;
  assign n1524 = n53550 & n53554;
  assign n1525 = n53551 & n1524;
  assign n1526 = n53550 & n1523;
  assign n1527 = n53553 & n53555;
  assign n1528 = n1475 & n1498;
  assign n1529 = ~n747 & ~n1234;
  assign n1530 = ~n646 & n1529;
  assign n1531 = ~n346 & ~n659;
  assign n1532 = ~n662 & ~n777;
  assign n1533 = n1531 & n1532;
  assign n1534 = ~n443 & ~n753;
  assign n1535 = n104 & n492;
  assign n1536 = ~n911 & ~n1535;
  assign n1537 = n1534 & n1536;
  assign n1538 = n1533 & n1537;
  assign n1539 = ~n646 & ~n753;
  assign n1540 = ~n443 & n1539;
  assign n1541 = ~n911 & ~n1234;
  assign n1542 = ~n747 & ~n1535;
  assign n1543 = n1529 & n1536;
  assign n1544 = n1541 & n1542;
  assign n1545 = n1533 & n53556;
  assign n1546 = n1540 & n1545;
  assign n1547 = n1530 & n1538;
  assign n1548 = n53500 & n53557;
  assign n1549 = n53552 & n1548;
  assign n1550 = n53451 & n53479;
  assign n1551 = n53451 & n53557;
  assign n1552 = n53500 & n53552;
  assign n1553 = n1551 & n1552;
  assign n1554 = n53479 & n1553;
  assign n1555 = n1549 & n1550;
  assign n1556 = n1533 & n1542;
  assign n1557 = n53549 & n1556;
  assign n1558 = n53500 & n1557;
  assign n1559 = n53552 & n1558;
  assign n1560 = n53479 & n1559;
  assign n1561 = n53451 & n1560;
  assign n1562 = n1541 & n1561;
  assign n1563 = ~n443 & n1562;
  assign n1564 = ~n646 & n1563;
  assign n1565 = ~n753 & n1564;
  assign n1566 = n53549 & n53558;
  assign n1567 = ~n53537 & ~n53559;
  assign n1568 = n53537 & n53559;
  assign n1569 = ~pi29  & ~n1567;
  assign n1570 = ~n1567 & ~n1568;
  assign n1571 = ~pi29  & n1570;
  assign n1572 = ~n1568 & n1569;
  assign n1573 = ~n1567 & ~n53560;
  assign n1574 = n53487 & ~n1573;
  assign n1575 = ~n53487 & n1573;
  assign n1576 = pi31  & ~n94;
  assign n1577 = ~n440 & ~n617;
  assign n1578 = ~n618 & ~n851;
  assign n1579 = n1577 & n1578;
  assign n1580 = n1541 & n1578;
  assign n1581 = n1577 & n1580;
  assign n1582 = n1541 & n1579;
  assign n1583 = ~n591 & ~n611;
  assign n1584 = n850 & n1583;
  assign n1585 = n463 & n1584;
  assign n1586 = n1541 & n1577;
  assign n1587 = n1583 & n1586;
  assign n1588 = n850 & n1578;
  assign n1589 = n463 & n1588;
  assign n1590 = n1587 & n1589;
  assign n1591 = n462 & n850;
  assign n1592 = n1578 & n1591;
  assign n1593 = ~n459 & ~n611;
  assign n1594 = ~n591 & n1593;
  assign n1595 = n1586 & n1594;
  assign n1596 = n1592 & n1595;
  assign n1597 = n53561 & n1585;
  assign n1598 = n53504 & n53562;
  assign n1599 = n53471 & n1577;
  assign n1600 = n53504 & n1599;
  assign n1601 = n1578 & n1600;
  assign n1602 = n1541 & n1601;
  assign n1603 = n850 & n1602;
  assign n1604 = n462 & n1603;
  assign n1605 = ~n459 & n1604;
  assign n1606 = ~n591 & n1605;
  assign n1607 = ~n611 & n1606;
  assign n1608 = n53471 & n1598;
  assign n1609 = ~n914 & ~n1280;
  assign n1610 = ~n1042 & ~n1337;
  assign n1611 = ~n1189 & n1610;
  assign n1612 = ~n1189 & ~n1280;
  assign n1613 = ~n914 & n1612;
  assign n1614 = ~n1337 & n1613;
  assign n1615 = ~n1042 & n1614;
  assign n1616 = ~n1042 & ~n1280;
  assign n1617 = ~n914 & ~n1189;
  assign n1618 = ~n1337 & n1617;
  assign n1619 = n1616 & n1618;
  assign n1620 = ~n1280 & ~n1337;
  assign n1621 = ~n914 & ~n1042;
  assign n1622 = ~n1189 & n1621;
  assign n1623 = n1620 & n1622;
  assign n1624 = n1609 & n1611;
  assign n1625 = ~n852 & ~n1457;
  assign n1626 = n53564 & n1625;
  assign n1627 = ~n1457 & n53564;
  assign n1628 = ~n852 & n53563;
  assign n1629 = n1627 & n1628;
  assign n1630 = n53563 & n53564;
  assign n1631 = ~n1457 & n1630;
  assign n1632 = ~n852 & n1631;
  assign n1633 = n53563 & n1626;
  assign n1634 = n162 & n267;
  assign n1635 = ~n1059 & ~n1455;
  assign n1636 = ~n1455 & ~n1634;
  assign n1637 = ~n1059 & n1636;
  assign n1638 = ~n1059 & ~n1634;
  assign n1639 = ~n1455 & n1638;
  assign n1640 = ~n1634 & n1635;
  assign n1641 = n173 & n267;
  assign n1642 = ~n975 & ~n1535;
  assign n1643 = ~n1641 & n1642;
  assign n1644 = n165 & n267;
  assign n1645 = ~n1034 & ~n1644;
  assign n1646 = n181 & n267;
  assign n1647 = ~n956 & ~n1646;
  assign n1648 = n1645 & n1647;
  assign n1649 = ~n1641 & ~n1646;
  assign n1650 = ~n1644 & ~n1646;
  assign n1651 = ~n1641 & n1650;
  assign n1652 = ~n1644 & n1649;
  assign n1653 = ~n956 & ~n1034;
  assign n1654 = n1642 & n1653;
  assign n1655 = n53567 & n1654;
  assign n1656 = n1643 & n1648;
  assign n1657 = n53566 & n53568;
  assign n1658 = n160 & n267;
  assign n1659 = ~n319 & ~n1658;
  assign n1660 = ~n268 & n1659;
  assign n1661 = n847 & n1660;
  assign n1662 = n846 & n1659;
  assign n1663 = n798 & n1662;
  assign n1664 = ~n268 & ~n587;
  assign n1665 = n1642 & n1664;
  assign n1666 = n802 & n1665;
  assign n1667 = n1663 & n1666;
  assign n1668 = n1642 & ~n1667;
  assign n1669 = n805 & n1661;
  assign n1670 = ~n105 & ~n627;
  assign n1671 = ~n316 & ~n911;
  assign n1672 = ~n272 & ~n822;
  assign n1673 = ~n246 & ~n1191;
  assign n1674 = ~n504 & ~n914;
  assign n1675 = ~n1487 & n1674;
  assign n1676 = ~n447 & ~n1492;
  assign n1677 = ~n447 & ~n1465;
  assign n1678 = ~n1492 & n1677;
  assign n1679 = ~n1465 & n1676;
  assign n1680 = n111 & n878;
  assign n1681 = n104 & n878;
  assign n1682 = ~n1680 & ~n1681;
  assign n1683 = ~n141 & ~n748;
  assign n1684 = n1682 & n1683;
  assign n1685 = n1184 & n1682;
  assign n1686 = n1683 & n1685;
  assign n1687 = n1184 & n1684;
  assign n1688 = ~n1465 & n1682;
  assign n1689 = ~n1492 & n1688;
  assign n1690 = ~n141 & n1689;
  assign n1691 = ~n748 & n1690;
  assign n1692 = ~n423 & n1691;
  assign n1693 = ~n447 & n1692;
  assign n1694 = ~n788 & n1693;
  assign n1695 = ~n1492 & n1683;
  assign n1696 = ~n423 & ~n447;
  assign n1697 = ~n788 & ~n1465;
  assign n1698 = n1696 & n1697;
  assign n1699 = n1682 & n1698;
  assign n1700 = n1695 & n1699;
  assign n1701 = n53570 & n53571;
  assign n1702 = ~n108 & ~n292;
  assign n1703 = n183 & n878;
  assign n1704 = ~n659 & ~n1703;
  assign n1705 = ~n414 & ~n564;
  assign n1706 = n1704 & n1705;
  assign n1707 = n1702 & n1706;
  assign n1708 = ~n902 & ~n1196;
  assign n1709 = ~n1280 & ~n1491;
  assign n1710 = n1708 & n1709;
  assign n1711 = ~n404 & ~n1337;
  assign n1712 = ~n559 & ~n646;
  assign n1713 = n1711 & n1712;
  assign n1714 = n1710 & n1713;
  assign n1715 = n162 & n345;
  assign n1716 = ~n848 & ~n1715;
  assign n1717 = ~n256 & ~n320;
  assign n1718 = ~n320 & n1716;
  assign n1719 = ~n256 & n1718;
  assign n1720 = n1716 & n1717;
  assign n1721 = ~n212 & ~n219;
  assign n1722 = ~n212 & ~n896;
  assign n1723 = ~n219 & n1722;
  assign n1724 = ~n896 & n1721;
  assign n1725 = n53573 & n53574;
  assign n1726 = n1714 & n1725;
  assign n1727 = n1704 & n1712;
  assign n1728 = n1702 & n1727;
  assign n1729 = n1705 & n1711;
  assign n1730 = n1710 & n1729;
  assign n1731 = n1725 & n1730;
  assign n1732 = n1728 & n1731;
  assign n1733 = n1705 & n1712;
  assign n1734 = n1708 & n1733;
  assign n1735 = n1702 & n1711;
  assign n1736 = n1704 & n1709;
  assign n1737 = n1735 & n1736;
  assign n1738 = n1725 & n1737;
  assign n1739 = n1734 & n1738;
  assign n1740 = n1709 & n1733;
  assign n1741 = n1704 & n1708;
  assign n1742 = n1735 & n1741;
  assign n1743 = n1725 & n1742;
  assign n1744 = n1740 & n1743;
  assign n1745 = n1707 & n1726;
  assign n1746 = n1709 & n1711;
  assign n1747 = n1702 & n1746;
  assign n1748 = n53573 & n1747;
  assign n1749 = n1705 & n1748;
  assign n1750 = n53572 & n1749;
  assign n1751 = n1712 & n1750;
  assign n1752 = n1704 & n1751;
  assign n1753 = n1708 & n1752;
  assign n1754 = ~n896 & n1753;
  assign n1755 = ~n219 & n1754;
  assign n1756 = ~n212 & n1755;
  assign n1757 = n53572 & n53575;
  assign n1758 = ~n206 & ~n496;
  assign n1759 = n624 & n1758;
  assign n1760 = ~n461 & ~n465;
  assign n1761 = n775 & n1760;
  assign n1762 = n1759 & n1761;
  assign n1763 = ~n222 & ~n823;
  assign n1764 = ~n823 & ~n1061;
  assign n1765 = ~n222 & n1764;
  assign n1766 = ~n222 & ~n1061;
  assign n1767 = ~n823 & n1766;
  assign n1768 = ~n1061 & n1763;
  assign n1769 = n165 & n345;
  assign n1770 = ~n733 & ~n1769;
  assign n1771 = ~n1471 & n1770;
  assign n1772 = n53577 & n1771;
  assign n1773 = ~n206 & ~n1471;
  assign n1774 = n775 & n1773;
  assign n1775 = n624 & n1760;
  assign n1776 = n1774 & n1775;
  assign n1777 = ~n496 & ~n733;
  assign n1778 = ~n1769 & n1777;
  assign n1779 = n53577 & n1778;
  assign n1780 = n1776 & n1779;
  assign n1781 = ~n733 & ~n1471;
  assign n1782 = ~n206 & ~n465;
  assign n1783 = n1781 & n1782;
  assign n1784 = n624 & n775;
  assign n1785 = n1783 & n1784;
  assign n1786 = ~n461 & ~n1769;
  assign n1787 = ~n496 & n1786;
  assign n1788 = n53577 & n1787;
  assign n1789 = n1785 & n1788;
  assign n1790 = n1762 & n1772;
  assign n1791 = n53576 & n53577;
  assign n1792 = n775 & n1791;
  assign n1793 = n624 & n1792;
  assign n1794 = ~n1471 & n1793;
  assign n1795 = ~n206 & n1794;
  assign n1796 = ~n496 & n1795;
  assign n1797 = ~n461 & n1796;
  assign n1798 = ~n733 & n1797;
  assign n1799 = ~n465 & n1798;
  assign n1800 = ~n1769 & n1799;
  assign n1801 = n53576 & n53578;
  assign n1802 = ~n1062 & ~n1457;
  assign n1803 = ~n651 & ~n1127;
  assign n1804 = ~n416 & ~n591;
  assign n1805 = n1803 & n1804;
  assign n1806 = ~n416 & n1803;
  assign n1807 = ~n1062 & n1806;
  assign n1808 = ~n1457 & n1807;
  assign n1809 = ~n591 & n1808;
  assign n1810 = ~n416 & ~n1062;
  assign n1811 = ~n591 & ~n1457;
  assign n1812 = n1802 & n1804;
  assign n1813 = n1810 & n1811;
  assign n1814 = n1803 & n53581;
  assign n1815 = n1802 & n1805;
  assign n1816 = ~n363 & ~n747;
  assign n1817 = ~n503 & n1816;
  assign n1818 = ~n450 & ~n617;
  assign n1819 = ~n565 & ~n735;
  assign n1820 = ~n357 & ~n983;
  assign n1821 = n1819 & n1820;
  assign n1822 = n1818 & n1820;
  assign n1823 = n1819 & n1822;
  assign n1824 = n1818 & n1821;
  assign n1825 = ~n503 & ~n983;
  assign n1826 = ~n357 & n1825;
  assign n1827 = n1816 & n1818;
  assign n1828 = n1819 & n1827;
  assign n1829 = n1826 & n1828;
  assign n1830 = ~n735 & ~n983;
  assign n1831 = ~n565 & n1830;
  assign n1832 = ~n357 & ~n503;
  assign n1833 = n1818 & n1832;
  assign n1834 = n1816 & n1833;
  assign n1835 = n1831 & n1834;
  assign n1836 = n1817 & n53582;
  assign n1837 = n53580 & n1816;
  assign n1838 = ~n983 & n1837;
  assign n1839 = ~n565 & n1838;
  assign n1840 = ~n503 & n1839;
  assign n1841 = ~n617 & n1840;
  assign n1842 = ~n357 & n1841;
  assign n1843 = ~n450 & n1842;
  assign n1844 = ~n735 & n1843;
  assign n1845 = n53580 & n53583;
  assign n1846 = ~n166 & ~n628;
  assign n1847 = ~n460 & ~n628;
  assign n1848 = ~n166 & n1847;
  assign n1849 = ~n460 & n1846;
  assign n1850 = ~n354 & ~n771;
  assign n1851 = ~n247 & ~n495;
  assign n1852 = ~n271 & ~n506;
  assign n1853 = n1851 & n1852;
  assign n1854 = ~n495 & ~n771;
  assign n1855 = ~n247 & ~n354;
  assign n1856 = n1854 & n1855;
  assign n1857 = n1852 & n1856;
  assign n1858 = n1850 & n1853;
  assign n1859 = ~n271 & n53585;
  assign n1860 = ~n247 & n1859;
  assign n1861 = ~n495 & n1860;
  assign n1862 = ~n506 & n1861;
  assign n1863 = ~n354 & n1862;
  assign n1864 = ~n771 & n1863;
  assign n1865 = n53585 & n53586;
  assign n1866 = ~n112 & ~n258;
  assign n1867 = n814 & n1866;
  assign n1868 = ~n514 & ~n1490;
  assign n1869 = ~n179 & ~n789;
  assign n1870 = ~n789 & ~n1490;
  assign n1871 = ~n179 & ~n514;
  assign n1872 = n1870 & n1871;
  assign n1873 = n1868 & n1869;
  assign n1874 = n1867 & n53588;
  assign n1875 = ~n182 & ~n296;
  assign n1876 = ~n296 & ~n1042;
  assign n1877 = ~n182 & n1876;
  assign n1878 = ~n182 & ~n1042;
  assign n1879 = ~n296 & n1878;
  assign n1880 = ~n1042 & n1875;
  assign n1881 = n100 & n345;
  assign n1882 = ~n364 & ~n1881;
  assign n1883 = n1273 & n1882;
  assign n1884 = n53474 & n1883;
  assign n1885 = n53589 & n1884;
  assign n1886 = n1273 & n1869;
  assign n1887 = n1866 & n1868;
  assign n1888 = n1886 & n1887;
  assign n1889 = n814 & n1882;
  assign n1890 = n53474 & n1889;
  assign n1891 = n53589 & n1890;
  assign n1892 = n1888 & n1891;
  assign n1893 = n1867 & n1883;
  assign n1894 = n53474 & n53588;
  assign n1895 = n53589 & n1894;
  assign n1896 = n1893 & n1895;
  assign n1897 = n1874 & n1885;
  assign n1898 = n53587 & n53590;
  assign n1899 = n1866 & n53589;
  assign n1900 = n53587 & n1899;
  assign n1901 = n53584 & n1900;
  assign n1902 = n814 & n1901;
  assign n1903 = n1273 & n1902;
  assign n1904 = n53474 & n1903;
  assign n1905 = ~n1490 & n1904;
  assign n1906 = ~n179 & n1905;
  assign n1907 = ~n514 & n1906;
  assign n1908 = ~n364 & n1907;
  assign n1909 = ~n789 & n1908;
  assign n1910 = ~n1881 & n1909;
  assign n1911 = n53584 & n1898;
  assign n1912 = n53446 & n345;
  assign n1913 = ~n353 & ~n618;
  assign n1914 = ~n618 & ~n1912;
  assign n1915 = ~n353 & n1914;
  assign n1916 = ~n353 & ~n1912;
  assign n1917 = ~n618 & n1916;
  assign n1918 = ~n1912 & n1913;
  assign n1919 = ~n255 & ~n1469;
  assign n1920 = ~n824 & n1346;
  assign n1921 = ~n824 & ~n1469;
  assign n1922 = ~n255 & n1921;
  assign n1923 = n1346 & n1922;
  assign n1924 = n1919 & n1920;
  assign n1925 = n1346 & n53592;
  assign n1926 = ~n1469 & n1925;
  assign n1927 = ~n255 & n1926;
  assign n1928 = ~n824 & n1927;
  assign n1929 = n53592 & n53593;
  assign n1930 = ~n444 & ~n742;
  assign n1931 = ~n1079 & ~n1477;
  assign n1932 = ~n444 & ~n1477;
  assign n1933 = ~n742 & ~n1079;
  assign n1934 = n1932 & n1933;
  assign n1935 = n1930 & n1931;
  assign n1936 = ~n568 & ~n1124;
  assign n1937 = n175 & n1936;
  assign n1938 = n53595 & n1937;
  assign n1939 = ~n879 & ~n894;
  assign n1940 = ~n405 & n1939;
  assign n1941 = ~n317 & ~n499;
  assign n1942 = ~n317 & ~n849;
  assign n1943 = ~n499 & n1942;
  assign n1944 = ~n849 & n1941;
  assign n1945 = n1940 & n53596;
  assign n1946 = n1938 & n1945;
  assign n1947 = ~n101 & ~n291;
  assign n1948 = ~n291 & ~n777;
  assign n1949 = ~n101 & n1948;
  assign n1950 = ~n777 & n1947;
  assign n1951 = ~n291 & n1032;
  assign n1952 = ~n101 & n1951;
  assign n1953 = ~n777 & n1952;
  assign n1954 = n1032 & n53597;
  assign n1955 = ~n415 & ~n511;
  assign n1956 = ~n321 & ~n1125;
  assign n1957 = ~n664 & ~n832;
  assign n1958 = n1956 & n1957;
  assign n1959 = n1955 & n1958;
  assign n1960 = n53598 & n1959;
  assign n1961 = n175 & n1955;
  assign n1962 = n53595 & n1961;
  assign n1963 = n1945 & n1962;
  assign n1964 = n1936 & n1956;
  assign n1965 = n1957 & n1964;
  assign n1966 = n53598 & n1965;
  assign n1967 = n1963 & n1966;
  assign n1968 = ~n742 & ~n1124;
  assign n1969 = ~n444 & ~n1079;
  assign n1970 = n1968 & n1969;
  assign n1971 = ~n568 & ~n1477;
  assign n1972 = n1957 & n1971;
  assign n1973 = n1970 & n1972;
  assign n1974 = n1945 & n1973;
  assign n1975 = n175 & n1956;
  assign n1976 = n1955 & n1975;
  assign n1977 = n53598 & n1976;
  assign n1978 = n1974 & n1977;
  assign n1979 = n1946 & n1960;
  assign n1980 = n53594 & n53599;
  assign n1981 = n53591 & n1980;
  assign n1982 = n1945 & n1956;
  assign n1983 = n53598 & n1982;
  assign n1984 = n53579 & n1983;
  assign n1985 = n53591 & n1984;
  assign n1986 = n53594 & n1985;
  assign n1987 = n1955 & n1986;
  assign n1988 = n1957 & n1987;
  assign n1989 = n175 & n1988;
  assign n1990 = ~n1124 & n1989;
  assign n1991 = ~n1079 & n1990;
  assign n1992 = ~n1477 & n1991;
  assign n1993 = ~n568 & n1992;
  assign n1994 = ~n742 & n1993;
  assign n1995 = ~n444 & n1994;
  assign n1996 = n53579 & n1981;
  assign n1997 = n171 & n878;
  assign n1998 = ~n346 & ~n1997;
  assign n1999 = ~n984 & ~n1085;
  assign n2000 = n1998 & n1999;
  assign n2001 = ~n310 & ~n647;
  assign n2002 = ~n308 & ~n567;
  assign n2003 = n2001 & n2002;
  assign n2004 = ~n1065 & ~n1466;
  assign n2005 = ~n584 & ~n829;
  assign n2006 = n2004 & n2005;
  assign n2007 = n2003 & n2006;
  assign n2008 = ~n1085 & n2004;
  assign n2009 = ~n984 & n2008;
  assign n2010 = ~n1997 & n2009;
  assign n2011 = ~n567 & n2010;
  assign n2012 = ~n308 & n2011;
  assign n2013 = ~n310 & n2012;
  assign n2014 = ~n584 & n2013;
  assign n2015 = ~n829 & n2014;
  assign n2016 = ~n647 & n2015;
  assign n2017 = ~n346 & n2016;
  assign n2018 = ~n308 & ~n984;
  assign n2019 = n2005 & n2018;
  assign n2020 = ~n346 & ~n1085;
  assign n2021 = ~n567 & ~n1997;
  assign n2022 = n2020 & n2021;
  assign n2023 = n2001 & n2004;
  assign n2024 = n2022 & n2023;
  assign n2025 = n2019 & n2024;
  assign n2026 = ~n346 & ~n984;
  assign n2027 = ~n308 & ~n310;
  assign n2028 = n2026 & n2027;
  assign n2029 = ~n829 & ~n1997;
  assign n2030 = ~n567 & ~n584;
  assign n2031 = n2029 & n2030;
  assign n2032 = ~n647 & ~n1085;
  assign n2033 = n2004 & n2032;
  assign n2034 = n2031 & n2033;
  assign n2035 = n2028 & n2034;
  assign n2036 = n2000 & n2007;
  assign n2037 = ~n663 & ~n830;
  assign n2038 = ~n615 & ~n1088;
  assign n2039 = ~n177 & ~n311;
  assign n2040 = n2038 & n2039;
  assign n2041 = n2037 & n2040;
  assign n2042 = n181 & n345;
  assign n2043 = ~n751 & ~n2042;
  assign n2044 = ~n510 & ~n1472;
  assign n2045 = ~n751 & n2044;
  assign n2046 = ~n2042 & n2045;
  assign n2047 = ~n1472 & ~n2042;
  assign n2048 = ~n510 & ~n751;
  assign n2049 = n2047 & n2048;
  assign n2050 = n2043 & n2044;
  assign n2051 = ~n410 & ~n753;
  assign n2052 = ~n1033 & n2051;
  assign n2053 = ~n356 & ~n440;
  assign n2054 = ~n211 & ~n216;
  assign n2055 = n2053 & n2054;
  assign n2056 = n2052 & n2055;
  assign n2057 = n53602 & n2056;
  assign n2058 = ~n663 & ~n1033;
  assign n2059 = n53602 & n2053;
  assign n2060 = n2038 & n2059;
  assign n2061 = n2058 & n2060;
  assign n2062 = ~n177 & n2061;
  assign n2063 = ~n211 & n2062;
  assign n2064 = ~n311 & n2063;
  assign n2065 = ~n216 & n2064;
  assign n2066 = ~n830 & n2065;
  assign n2067 = ~n410 & n2066;
  assign n2068 = ~n753 & n2067;
  assign n2069 = n2038 & n2053;
  assign n2070 = n2039 & n2069;
  assign n2071 = ~n211 & ~n830;
  assign n2072 = ~n410 & n2071;
  assign n2073 = ~n216 & ~n753;
  assign n2074 = n2058 & n2073;
  assign n2075 = ~n410 & ~n830;
  assign n2076 = ~n753 & n2075;
  assign n2077 = n2054 & n2058;
  assign n2078 = n2076 & n2077;
  assign n2079 = n2072 & n2074;
  assign n2080 = n53602 & n53604;
  assign n2081 = n2070 & n2080;
  assign n2082 = n2038 & n2058;
  assign n2083 = n2053 & n2082;
  assign n2084 = ~n216 & ~n830;
  assign n2085 = ~n410 & n2084;
  assign n2086 = ~n211 & ~n753;
  assign n2087 = n2039 & n2086;
  assign n2088 = n2085 & n2087;
  assign n2089 = n53602 & n2088;
  assign n2090 = n2083 & n2089;
  assign n2091 = n2041 & n2057;
  assign n2092 = ~n349 & ~n1192;
  assign n2093 = ~n977 & ~n1478;
  assign n2094 = ~n459 & ~n948;
  assign n2095 = n2093 & n2094;
  assign n2096 = n2092 & n2095;
  assign n2097 = ~n402 & ~n851;
  assign n2098 = n494 & n2097;
  assign n2099 = ~n340 & ~n466;
  assign n2100 = n799 & n2099;
  assign n2101 = n2098 & n2100;
  assign n2102 = ~n360 & ~n1486;
  assign n2103 = n107 & n878;
  assign n2104 = ~n221 & ~n2103;
  assign n2105 = ~n1486 & ~n2103;
  assign n2106 = ~n221 & n2105;
  assign n2107 = ~n360 & n2106;
  assign n2108 = n2102 & n2104;
  assign n2109 = n160 & n345;
  assign n2110 = ~n464 & ~n590;
  assign n2111 = ~n590 & ~n2109;
  assign n2112 = ~n464 & n2111;
  assign n2113 = ~n464 & ~n2109;
  assign n2114 = ~n590 & n2113;
  assign n2115 = ~n2109 & n2110;
  assign n2116 = n53605 & n53606;
  assign n2117 = n2101 & n2116;
  assign n2118 = n2092 & n2116;
  assign n2119 = n799 & n2118;
  assign n2120 = n494 & n2119;
  assign n2121 = n2093 & n2120;
  assign n2122 = n2094 & n2121;
  assign n2123 = ~n402 & n2122;
  assign n2124 = ~n851 & n2123;
  assign n2125 = ~n466 & n2124;
  assign n2126 = ~n340 & n2125;
  assign n2127 = n2092 & n2094;
  assign n2128 = n494 & n2127;
  assign n2129 = ~n340 & ~n851;
  assign n2130 = ~n402 & ~n466;
  assign n2131 = n2129 & n2130;
  assign n2132 = n799 & n2093;
  assign n2133 = n799 & n2097;
  assign n2134 = n2093 & n2099;
  assign n2135 = n2133 & n2134;
  assign n2136 = n2131 & n2132;
  assign n2137 = n2116 & n53608;
  assign n2138 = n2128 & n2137;
  assign n2139 = n2096 & n2117;
  assign n2140 = ~n184 & ~n770;
  assign n2141 = ~n631 & ~n1195;
  assign n2142 = ~n295 & ~n344;
  assign n2143 = n2141 & n2142;
  assign n2144 = ~n295 & ~n631;
  assign n2145 = ~n1195 & n2144;
  assign n2146 = ~n184 & n2145;
  assign n2147 = ~n344 & n2146;
  assign n2148 = ~n770 & n2147;
  assign n2149 = n2140 & n2141;
  assign n2150 = n2142 & n2149;
  assign n2151 = n2140 & n2143;
  assign n2152 = ~n207 & ~n662;
  assign n2153 = ~n498 & ~n776;
  assign n2154 = ~n776 & ~n1234;
  assign n2155 = ~n498 & n2154;
  assign n2156 = ~n1234 & n2153;
  assign n2157 = ~n1234 & n2152;
  assign n2158 = ~n498 & n2157;
  assign n2159 = ~n776 & n2158;
  assign n2160 = n2152 & n53610;
  assign n2161 = ~n342 & ~n833;
  assign n2162 = ~n307 & ~n1090;
  assign n2163 = ~n562 & ~n901;
  assign n2164 = n2162 & n2163;
  assign n2165 = n2161 & n2164;
  assign n2166 = n53611 & n2165;
  assign n2167 = n53609 & n2166;
  assign n2168 = ~n451 & ~n507;
  assign n2169 = ~n507 & ~n1468;
  assign n2170 = ~n451 & n2169;
  assign n2171 = ~n1468 & n2168;
  assign n2172 = ~n294 & ~n881;
  assign n2173 = ~n144 & n2172;
  assign n2174 = ~n883 & ~n1476;
  assign n2175 = ~n409 & ~n922;
  assign n2176 = n2174 & n2175;
  assign n2177 = ~n144 & ~n883;
  assign n2178 = ~n1476 & n2177;
  assign n2179 = n2172 & n2175;
  assign n2180 = n2178 & n2179;
  assign n2181 = ~n922 & n2177;
  assign n2182 = ~n409 & ~n1476;
  assign n2183 = n2172 & n2182;
  assign n2184 = n2181 & n2183;
  assign n2185 = n2173 & n2176;
  assign n2186 = n53612 & n2172;
  assign n2187 = ~n922 & n2186;
  assign n2188 = ~n883 & n2187;
  assign n2189 = ~n1476 & n2188;
  assign n2190 = ~n144 & n2189;
  assign n2191 = ~n409 & n2190;
  assign n2192 = n53612 & n53613;
  assign n2193 = ~n168 & ~n852;
  assign n2194 = ~n168 & ~n249;
  assign n2195 = ~n852 & n2194;
  assign n2196 = ~n249 & ~n852;
  assign n2197 = ~n168 & n2196;
  assign n2198 = ~n249 & n2193;
  assign n2199 = ~n218 & ~n401;
  assign n2200 = ~n740 & n2199;
  assign n2201 = n173 & n345;
  assign n2202 = ~n215 & ~n2201;
  assign n2203 = n421 & n2202;
  assign n2204 = n2200 & n2203;
  assign n2205 = n53615 & n2204;
  assign n2206 = n53614 & n2205;
  assign n2207 = n421 & n2163;
  assign n2208 = n2161 & n2207;
  assign n2209 = n53611 & n2208;
  assign n2210 = n53609 & n2209;
  assign n2211 = ~n218 & n2202;
  assign n2212 = ~n401 & ~n740;
  assign n2213 = n2162 & n2212;
  assign n2214 = n2211 & n2213;
  assign n2215 = n53615 & n2214;
  assign n2216 = n53614 & n2215;
  assign n2217 = n2210 & n2216;
  assign n2218 = ~n218 & ~n2201;
  assign n2219 = n2162 & n2218;
  assign n2220 = n421 & n2219;
  assign n2221 = n53611 & n2220;
  assign n2222 = n53609 & n2221;
  assign n2223 = ~n740 & n2161;
  assign n2224 = ~n215 & ~n401;
  assign n2225 = n2163 & n2224;
  assign n2226 = n2223 & n2225;
  assign n2227 = n53615 & n2226;
  assign n2228 = n53614 & n2227;
  assign n2229 = n2222 & n2228;
  assign n2230 = n2167 & n2206;
  assign n2231 = n53611 & n53615;
  assign n2232 = n53609 & n2231;
  assign n2233 = n53607 & n2232;
  assign n2234 = n53614 & n2233;
  assign n2235 = n421 & n2234;
  assign n2236 = ~n1090 & n2235;
  assign n2237 = ~n901 & n2236;
  assign n2238 = ~n215 & n2237;
  assign n2239 = ~n307 & n2238;
  assign n2240 = ~n218 & n2239;
  assign n2241 = ~n562 & n2240;
  assign n2242 = ~n401 & n2241;
  assign n2243 = ~n833 & n2242;
  assign n2244 = ~n342 & n2243;
  assign n2245 = ~n740 & n2244;
  assign n2246 = ~n2201 & n2245;
  assign n2247 = n53607 & n53616;
  assign n2248 = ~n259 & ~n611;
  assign n2249 = ~n259 & ~n1081;
  assign n2250 = ~n611 & n2249;
  assign n2251 = ~n1081 & n2248;
  assign n2252 = ~n1081 & n1391;
  assign n2253 = ~n259 & n2252;
  assign n2254 = ~n611 & n2253;
  assign n2255 = n1391 & n53618;
  assign n2256 = ~n361 & ~n560;
  assign n2257 = ~n250 & ~n422;
  assign n2258 = ~n650 & ~n957;
  assign n2259 = ~n422 & ~n957;
  assign n2260 = ~n250 & n2259;
  assign n2261 = ~n650 & n2260;
  assign n2262 = n2257 & n2258;
  assign n2263 = ~n408 & ~n625;
  assign n2264 = ~n408 & ~n750;
  assign n2265 = ~n625 & n2264;
  assign n2266 = ~n625 & ~n750;
  assign n2267 = ~n408 & n2266;
  assign n2268 = ~n750 & n2263;
  assign n2269 = n53620 & n53621;
  assign n2270 = n2256 & n2269;
  assign n2271 = n53619 & n2270;
  assign n2272 = n53617 & n2271;
  assign n2273 = n53603 & n2272;
  assign n2274 = n53601 & n2273;
  assign n2275 = n53600 & n2274;
  assign n2276 = n1675 & n2275;
  assign n2277 = n1673 & n2276;
  assign n2278 = n1672 & n2277;
  assign n2279 = n1671 & n2278;
  assign n2280 = n164 & n2279;
  assign n2281 = n1670 & n2280;
  assign n2282 = ~n1485 & n2281;
  assign n2283 = ~n348 & n2282;
  assign n2284 = n53567 & n1653;
  assign n2285 = n53566 & n1653;
  assign n2286 = ~n1646 & n2285;
  assign n2287 = ~n1644 & n2286;
  assign n2288 = ~n1641 & n2287;
  assign n2289 = n53566 & n2284;
  assign n2290 = n798 & n53623;
  assign n2291 = n846 & n2290;
  assign n2292 = n802 & n2291;
  assign n2293 = n1659 & n2292;
  assign n2294 = n1642 & n2293;
  assign n2295 = ~n587 & n2294;
  assign n2296 = ~n268 & n2295;
  assign n2297 = n1667 & n53623;
  assign n2298 = n1670 & n1671;
  assign n2299 = n1672 & n2298;
  assign n2300 = ~n348 & ~n1485;
  assign n2301 = n164 & n2300;
  assign n2302 = n1673 & n2256;
  assign n2303 = n2301 & n2302;
  assign n2304 = n164 & n1670;
  assign n2305 = n1672 & n2304;
  assign n2306 = n1671 & n2300;
  assign n2307 = n2302 & n2306;
  assign n2308 = n2305 & n2307;
  assign n2309 = n1671 & n1672;
  assign n2310 = n164 & n2309;
  assign n2311 = n2256 & n2300;
  assign n2312 = n1670 & n1673;
  assign n2313 = n2311 & n2312;
  assign n2314 = n2310 & n2313;
  assign n2315 = n2299 & n2303;
  assign n2316 = n53619 & n53624;
  assign n2317 = n1675 & n53620;
  assign n2318 = n53621 & n2317;
  assign n2319 = n53601 & n2318;
  assign n2320 = n2316 & n2319;
  assign n2321 = n53603 & n2320;
  assign n2322 = n53617 & n2321;
  assign n2323 = n53600 & n2322;
  assign n2324 = n1657 & ~n53569;
  assign n2325 = n53565 & ~n53622;
  assign n2326 = ~n879 & ~n1703;
  assign n2327 = ~n1191 & ~n2103;
  assign n2328 = ~n1061 & ~n1127;
  assign n2329 = n2327 & n2328;
  assign n2330 = n2326 & n2327;
  assign n2331 = n2328 & n2330;
  assign n2332 = n2326 & n2329;
  assign n2333 = ~n1079 & ~n1192;
  assign n2334 = ~n977 & ~n1997;
  assign n2335 = ~n1997 & n2333;
  assign n2336 = ~n977 & n2335;
  assign n2337 = n2333 & n2334;
  assign n2338 = ~n901 & ~n1912;
  assign n2339 = n1682 & n2338;
  assign n2340 = ~n957 & ~n1062;
  assign n2341 = ~n983 & n2340;
  assign n2342 = n2339 & n2341;
  assign n2343 = n53626 & n2342;
  assign n2344 = n1682 & n2328;
  assign n2345 = n53626 & n2344;
  assign n2346 = n2338 & n2345;
  assign n2347 = n2326 & n2346;
  assign n2348 = n2340 & n2347;
  assign n2349 = ~n1191 & n2348;
  assign n2350 = ~n983 & n2349;
  assign n2351 = ~n2103 & n2350;
  assign n2352 = n2326 & n2340;
  assign n2353 = n2328 & n2352;
  assign n2354 = ~n983 & ~n2103;
  assign n2355 = ~n983 & n2327;
  assign n2356 = ~n1191 & n2354;
  assign n2357 = n2339 & n53628;
  assign n2358 = n53626 & n2357;
  assign n2359 = n2353 & n2358;
  assign n2360 = n1682 & n2340;
  assign n2361 = n2328 & n2360;
  assign n2362 = n2326 & n2338;
  assign n2363 = n53628 & n2362;
  assign n2364 = n53626 & n2363;
  assign n2365 = n2361 & n2364;
  assign n2366 = n53625 & n2343;
  assign n2367 = ~n2042 & ~n2109;
  assign n2368 = ~n1769 & ~n2201;
  assign n2369 = ~n2201 & n2367;
  assign n2370 = ~n1769 & n2369;
  assign n2371 = n2367 & n2368;
  assign n2372 = ~n1715 & ~n1881;
  assign n2373 = n53629 & n2372;
  assign n2374 = n53627 & n53629;
  assign n2375 = ~n1715 & n2374;
  assign n2376 = ~n1881 & n2375;
  assign n2377 = n53627 & n2373;
  assign n2378 = ~n590 & n799;
  assign n2379 = n799 & n53501;
  assign n2380 = n814 & n2378;
  assign n2381 = n626 & n53631;
  assign n2382 = n806 & n53501;
  assign n2383 = n626 & n53630;
  assign n2384 = n814 & n2383;
  assign n2385 = n799 & n2384;
  assign n2386 = ~n590 & n2385;
  assign n2387 = n53630 & n53632;
  assign n2388 = n53499 & n53633;
  assign n2389 = ~n1081 & ~n1457;
  assign n2390 = ~n53622 & n2389;
  assign n2391 = ~n53622 & n2388;
  assign n2392 = ~n1081 & n2391;
  assign n2393 = ~n1457 & n2392;
  assign n2394 = n2388 & n2390;
  assign n2395 = ~n414 & ~n464;
  assign n2396 = n418 & ~n464;
  assign n2397 = n417 & ~n464;
  assign n2398 = ~n414 & n2397;
  assign n2399 = n417 & n2395;
  assign n2400 = ~n1033 & ~n1044;
  assign n2401 = ~n422 & ~n628;
  assign n2402 = n2141 & n2401;
  assign n2403 = n2400 & n2402;
  assign n2404 = ~n894 & n1708;
  assign n2405 = ~n408 & ~n984;
  assign n2406 = ~n1065 & ~n1090;
  assign n2407 = n2405 & n2406;
  assign n2408 = n2404 & n2407;
  assign n2409 = n2141 & n2400;
  assign n2410 = n2141 & n2405;
  assign n2411 = n2400 & n2410;
  assign n2412 = n2405 & n2409;
  assign n2413 = ~n422 & ~n1090;
  assign n2414 = ~n628 & ~n1065;
  assign n2415 = n2401 & n2406;
  assign n2416 = n2413 & n2414;
  assign n2417 = n2404 & n53637;
  assign n2418 = n53636 & n2417;
  assign n2419 = n2403 & n2408;
  assign n2420 = ~n984 & ~n1065;
  assign n2421 = ~n408 & ~n628;
  assign n2422 = n2420 & n2421;
  assign n2423 = n2413 & n2422;
  assign n2424 = n2404 & n2409;
  assign n2425 = n53635 & n2424;
  assign n2426 = n2423 & n2425;
  assign n2427 = n53635 & n53638;
  assign n2428 = n53545 & n53639;
  assign n2429 = n53545 & n53635;
  assign n2430 = n2404 & n2429;
  assign n2431 = n53552 & n2430;
  assign n2432 = ~n984 & n2431;
  assign n2433 = ~n1033 & n2432;
  assign n2434 = ~n1065 & n2433;
  assign n2435 = ~n1044 & n2434;
  assign n2436 = ~n631 & n2435;
  assign n2437 = ~n422 & n2436;
  assign n2438 = ~n628 & n2437;
  assign n2439 = ~n1090 & n2438;
  assign n2440 = ~n408 & n2439;
  assign n2441 = ~n1195 & n2440;
  assign n2442 = n53552 & n2428;
  assign n2443 = n53463 & n53478;
  assign n2444 = n53463 & n53640;
  assign n2445 = n53477 & n2444;
  assign n2446 = ~n584 & n2445;
  assign n2447 = ~n587 & n2446;
  assign n2448 = n53640 & n2443;
  assign n2449 = ~n364 & ~n788;
  assign n2450 = ~n733 & ~n788;
  assign n2451 = ~n364 & n2450;
  assign n2452 = ~n733 & n2449;
  assign n2453 = n497 & n619;
  assign n2454 = ~n510 & ~n647;
  assign n2455 = n2099 & n2454;
  assign n2456 = n497 & n2454;
  assign n2457 = n619 & n2099;
  assign n2458 = n2456 & n2457;
  assign n2459 = n2453 & n2455;
  assign n2460 = ~n618 & n2456;
  assign n2461 = ~n617 & n2460;
  assign n2462 = ~n733 & n2461;
  assign n2463 = ~n466 & n2462;
  assign n2464 = ~n364 & n2463;
  assign n2465 = ~n340 & n2464;
  assign n2466 = ~n788 & n2465;
  assign n2467 = ~n466 & ~n788;
  assign n2468 = ~n618 & n2467;
  assign n2469 = ~n340 & ~n617;
  assign n2470 = ~n364 & ~n733;
  assign n2471 = n2469 & n2470;
  assign n2472 = n2456 & n2471;
  assign n2473 = n2468 & n2472;
  assign n2474 = n53642 & n53643;
  assign n2475 = ~n440 & n500;
  assign n2476 = ~n506 & ~n735;
  assign n2477 = ~n493 & ~n789;
  assign n2478 = n1541 & n2477;
  assign n2479 = n2476 & n2478;
  assign n2480 = ~n440 & n1541;
  assign n2481 = n500 & n2476;
  assign n2482 = n2477 & n2481;
  assign n2483 = n2480 & n2482;
  assign n2484 = ~n440 & n2476;
  assign n2485 = n500 & n1541;
  assign n2486 = n2477 & n2485;
  assign n2487 = n2484 & n2486;
  assign n2488 = n2475 & n2479;
  assign n2489 = n53644 & n53645;
  assign n2490 = n53498 & n2477;
  assign n2491 = n53644 & n2490;
  assign n2492 = n500 & n2491;
  assign n2493 = n1541 & n2492;
  assign n2494 = n2476 & n2493;
  assign n2495 = ~n440 & n2494;
  assign n2496 = n53498 & n2489;
  assign n2497 = ~n363 & ~n662;
  assign n2498 = n421 & ~n662;
  assign n2499 = ~n363 & n2498;
  assign n2500 = n421 & n2497;
  assign n2501 = ~n344 & ~n361;
  assign n2502 = ~n465 & n2501;
  assign n2503 = ~n649 & ~n659;
  assign n2504 = n798 & n2503;
  assign n2505 = ~n361 & ~n659;
  assign n2506 = ~n649 & n2505;
  assign n2507 = ~n344 & ~n465;
  assign n2508 = n798 & n2507;
  assign n2509 = n2506 & n2508;
  assign n2510 = ~n659 & n2507;
  assign n2511 = ~n361 & ~n649;
  assign n2512 = n798 & n2511;
  assign n2513 = n2510 & n2512;
  assign n2514 = ~n649 & n2501;
  assign n2515 = ~n465 & ~n659;
  assign n2516 = n798 & n2515;
  assign n2517 = n2514 & n2516;
  assign n2518 = n2502 & n2504;
  assign n2519 = n798 & n53647;
  assign n2520 = ~n659 & n2519;
  assign n2521 = ~n649 & n2520;
  assign n2522 = ~n465 & n2521;
  assign n2523 = ~n344 & n2522;
  assign n2524 = ~n361 & n2523;
  assign n2525 = n53647 & n53648;
  assign n2526 = n358 & ~n591;
  assign n2527 = n53564 & n2526;
  assign n2528 = n53649 & n2527;
  assign n2529 = n53646 & n2528;
  assign n2530 = n53641 & n53646;
  assign n2531 = n53649 & n2530;
  assign n2532 = n53564 & n2531;
  assign n2533 = n358 & n2532;
  assign n2534 = ~n591 & n2533;
  assign n2535 = n53641 & n2529;
  assign n2536 = ~n53634 & ~n53650;
  assign n2537 = ~n646 & ~n1641;
  assign n2538 = ~n1634 & ~n1646;
  assign n2539 = ~n742 & ~n1644;
  assign n2540 = n2538 & n2539;
  assign n2541 = n2537 & n2540;
  assign n2542 = ~n346 & ~n443;
  assign n2543 = ~n740 & n2542;
  assign n2544 = n53635 & n2543;
  assign n2545 = ~n740 & ~n742;
  assign n2546 = ~n1644 & n2545;
  assign n2547 = n2537 & n2542;
  assign n2548 = n2538 & n2547;
  assign n2549 = ~n346 & ~n740;
  assign n2550 = ~n742 & n2549;
  assign n2551 = ~n443 & ~n1644;
  assign n2552 = n2538 & n2551;
  assign n2553 = n2537 & n2552;
  assign n2554 = n2550 & n2553;
  assign n2555 = n2546 & n2548;
  assign n2556 = n53635 & n53651;
  assign n2557 = n53635 & n2537;
  assign n2558 = ~n742 & n2557;
  assign n2559 = ~n1646 & n2558;
  assign n2560 = ~n1634 & n2559;
  assign n2561 = ~n1644 & n2560;
  assign n2562 = ~n443 & n2561;
  assign n2563 = ~n740 & n2562;
  assign n2564 = ~n346 & n2563;
  assign n2565 = n2541 & n2544;
  assign n2566 = ~n748 & n1541;
  assign n2567 = ~n615 & ~n630;
  assign n2568 = ~n493 & ~n747;
  assign n2569 = n2567 & n2568;
  assign n2570 = n717 & n2569;
  assign n2571 = ~n493 & ~n615;
  assign n2572 = ~n630 & n2571;
  assign n2573 = n749 & n1541;
  assign n2574 = n2572 & n2573;
  assign n2575 = n717 & n2574;
  assign n2576 = n2566 & n2570;
  assign n2577 = ~n342 & ~n408;
  assign n2578 = n2401 & n2577;
  assign n2579 = ~n269 & ~n1658;
  assign n2580 = n1197 & n2579;
  assign n2581 = n1197 & n2401;
  assign n2582 = n2577 & n2579;
  assign n2583 = n2581 & n2582;
  assign n2584 = n2578 & n2580;
  assign n2585 = n53502 & n53654;
  assign n2586 = ~n628 & n2571;
  assign n2587 = ~n422 & ~n630;
  assign n2588 = n1197 & n2587;
  assign n2589 = n2586 & n2588;
  assign n2590 = n717 & n2589;
  assign n2591 = n749 & n2577;
  assign n2592 = n1541 & n2579;
  assign n2593 = n2591 & n2592;
  assign n2594 = n53502 & n2593;
  assign n2595 = n2590 & n2594;
  assign n2596 = n452 & n1541;
  assign n2597 = n1197 & n2596;
  assign n2598 = n424 & n2567;
  assign n2599 = n2591 & n2598;
  assign n2600 = ~n493 & ~n628;
  assign n2601 = n2579 & n2600;
  assign n2602 = n53502 & n2601;
  assign n2603 = n2599 & n2602;
  assign n2604 = n2597 & n2603;
  assign n2605 = n53653 & n2585;
  assign n2606 = n53552 & n53655;
  assign n2607 = n53652 & n53655;
  assign n2608 = n53552 & n2607;
  assign n2609 = n53652 & n2606;
  assign n2610 = n452 & n53502;
  assign n2611 = n53552 & n2610;
  assign n2612 = n1197 & n2611;
  assign n2613 = n53652 & n2612;
  assign n2614 = n53548 & n2613;
  assign n2615 = n1541 & n2614;
  assign n2616 = n2577 & n2615;
  assign n2617 = n424 & n2616;
  assign n2618 = n749 & n2617;
  assign n2619 = ~n628 & n2618;
  assign n2620 = ~n493 & n2619;
  assign n2621 = ~n1658 & n2620;
  assign n2622 = ~n630 & n2621;
  assign n2623 = ~n269 & n2622;
  assign n2624 = ~n615 & n2623;
  assign n2625 = n53548 & n53656;
  assign n2626 = ~n53650 & ~n53657;
  assign n2627 = ~n292 & ~n405;
  assign n2628 = ~n1189 & n2627;
  assign n2629 = ~n311 & ~n317;
  assign n2630 = ~n311 & ~n751;
  assign n2631 = ~n317 & n2630;
  assign n2632 = ~n317 & ~n751;
  assign n2633 = ~n311 & n2632;
  assign n2634 = ~n751 & n2629;
  assign n2635 = ~n1469 & ~n1912;
  assign n2636 = ~n211 & ~n2201;
  assign n2637 = n2635 & n2636;
  assign n2638 = n53658 & n2637;
  assign n2639 = n2628 & n2635;
  assign n2640 = ~n211 & n2639;
  assign n2641 = ~n317 & n2640;
  assign n2642 = ~n311 & n2641;
  assign n2643 = ~n751 & n2642;
  assign n2644 = ~n2201 & n2643;
  assign n2645 = n2628 & n2638;
  assign n2646 = ~n984 & ~n1769;
  assign n2647 = ~n984 & ~n1492;
  assign n2648 = ~n1769 & n2647;
  assign n2649 = ~n1492 & n2646;
  assign n2650 = ~n1492 & n1711;
  assign n2651 = n2646 & n2650;
  assign n2652 = n1711 & n53660;
  assign n2653 = n1711 & n53659;
  assign n2654 = ~n984 & n2653;
  assign n2655 = ~n1492 & n2654;
  assign n2656 = ~n1769 & n2655;
  assign n2657 = n53659 & n53661;
  assign n2658 = ~n308 & ~n1042;
  assign n2659 = ~n1042 & ~n1487;
  assign n2660 = ~n308 & n2659;
  assign n2661 = ~n1487 & n2658;
  assign n2662 = n462 & n624;
  assign n2663 = n749 & n1391;
  assign n2664 = n2662 & n2663;
  assign n2665 = n53663 & n2664;
  assign n2666 = ~n291 & ~n443;
  assign n2667 = n1185 & n2666;
  assign n2668 = ~n291 & n53550;
  assign n2669 = ~n219 & n2668;
  assign n2670 = ~n663 & n2669;
  assign n2671 = ~n443 & n2670;
  assign n2672 = n53550 & n2667;
  assign n2673 = n297 & n2105;
  assign n2674 = ~n212 & ~n423;
  assign n2675 = ~n307 & ~n630;
  assign n2676 = n2674 & n2675;
  assign n2677 = ~n1486 & n2675;
  assign n2678 = ~n295 & n2677;
  assign n2679 = ~n296 & n2678;
  assign n2680 = ~n2103 & n2679;
  assign n2681 = ~n212 & n2680;
  assign n2682 = ~n423 & n2681;
  assign n2683 = ~n212 & ~n2103;
  assign n2684 = ~n296 & ~n1486;
  assign n2685 = n2683 & n2684;
  assign n2686 = ~n295 & ~n423;
  assign n2687 = n2675 & n2686;
  assign n2688 = n2685 & n2687;
  assign n2689 = n2673 & n2676;
  assign n2690 = ~n256 & ~n1465;
  assign n2691 = ~n215 & ~n1715;
  assign n2692 = n2690 & n2691;
  assign n2693 = ~n615 & ~n1881;
  assign n2694 = ~n250 & ~n1468;
  assign n2695 = n2693 & n2694;
  assign n2696 = n2690 & n2694;
  assign n2697 = n2691 & n2693;
  assign n2698 = n2696 & n2697;
  assign n2699 = n2692 & n2695;
  assign n2700 = n53665 & n53666;
  assign n2701 = n53664 & n2700;
  assign n2702 = n462 & n1391;
  assign n2703 = n624 & n2693;
  assign n2704 = n2702 & n2703;
  assign n2705 = n53663 & n2704;
  assign n2706 = n2691 & n2694;
  assign n2707 = n749 & n2690;
  assign n2708 = n2706 & n2707;
  assign n2709 = n53665 & n2708;
  assign n2710 = n53664 & n2709;
  assign n2711 = n2705 & n2710;
  assign n2712 = ~n308 & ~n1468;
  assign n2713 = ~n1487 & n2712;
  assign n2714 = ~n250 & ~n1042;
  assign n2715 = n624 & n2714;
  assign n2716 = n1391 & n2690;
  assign n2717 = n2715 & n2716;
  assign n2718 = n2713 & n2717;
  assign n2719 = n749 & n2693;
  assign n2720 = n462 & n2691;
  assign n2721 = n2719 & n2720;
  assign n2722 = n53664 & n2721;
  assign n2723 = n53665 & n2722;
  assign n2724 = n2718 & n2723;
  assign n2725 = n2665 & n2701;
  assign n2726 = n53662 & n2692;
  assign n2727 = n53665 & n2726;
  assign n2728 = n53664 & n2727;
  assign n2729 = n624 & n2728;
  assign n2730 = n749 & n2729;
  assign n2731 = n2693 & n2730;
  assign n2732 = n1391 & n2731;
  assign n2733 = n462 & n2732;
  assign n2734 = ~n1487 & n2733;
  assign n2735 = ~n1468 & n2734;
  assign n2736 = ~n308 & n2735;
  assign n2737 = ~n250 & n2736;
  assign n2738 = ~n1042 & n2737;
  assign n2739 = n53662 & n53667;
  assign n2740 = n799 & ~n1472;
  assign n2741 = ~n310 & ~n507;
  assign n2742 = ~n216 & ~n294;
  assign n2743 = n2367 & n2742;
  assign n2744 = n2741 & n2743;
  assign n2745 = n2740 & n2741;
  assign n2746 = n2367 & n2745;
  assign n2747 = ~n294 & n2746;
  assign n2748 = ~n216 & n2747;
  assign n2749 = n2740 & n2744;
  assign n2750 = ~n503 & ~n740;
  assign n2751 = ~n774 & n2750;
  assign n2752 = ~n1471 & ~n1490;
  assign n2753 = ~n247 & ~n625;
  assign n2754 = n2752 & n2753;
  assign n2755 = ~n247 & ~n503;
  assign n2756 = ~n740 & n2755;
  assign n2757 = ~n625 & ~n774;
  assign n2758 = n2752 & n2757;
  assign n2759 = n2756 & n2758;
  assign n2760 = ~n247 & ~n740;
  assign n2761 = ~n247 & ~n774;
  assign n2762 = ~n740 & n2761;
  assign n2763 = ~n774 & n2760;
  assign n2764 = ~n625 & ~n1471;
  assign n2765 = ~n503 & ~n1490;
  assign n2766 = ~n503 & ~n625;
  assign n2767 = n2752 & n2766;
  assign n2768 = n2764 & n2765;
  assign n2769 = n53671 & n53672;
  assign n2770 = n2751 & n2754;
  assign n2771 = n322 & ~n1485;
  assign n2772 = ~n451 & ~n664;
  assign n2773 = ~n258 & ~n1466;
  assign n2774 = ~n664 & n2773;
  assign n2775 = ~n451 & n2774;
  assign n2776 = ~n451 & ~n1466;
  assign n2777 = ~n258 & ~n664;
  assign n2778 = n2776 & n2777;
  assign n2779 = n2772 & n2773;
  assign n2780 = n2771 & n53673;
  assign n2781 = n53670 & n2780;
  assign n2782 = n273 & ~n342;
  assign n2783 = ~n316 & ~n742;
  assign n2784 = n1709 & n2783;
  assign n2785 = ~n271 & n2784;
  assign n2786 = ~n272 & n2785;
  assign n2787 = ~n342 & n2786;
  assign n2788 = ~n342 & n2783;
  assign n2789 = n273 & n1709;
  assign n2790 = n2788 & n2789;
  assign n2791 = n2782 & n2784;
  assign n2792 = ~n450 & ~n789;
  assign n2793 = ~n450 & ~n1641;
  assign n2794 = ~n789 & n2793;
  assign n2795 = ~n1641 & n2792;
  assign n2796 = n403 & ~n1641;
  assign n2797 = ~n450 & n2796;
  assign n2798 = ~n789 & n2797;
  assign n2799 = n403 & n53675;
  assign n2800 = n53674 & n53676;
  assign n2801 = n2781 & n2800;
  assign n2802 = n2771 & n53676;
  assign n2803 = n53669 & n2802;
  assign n2804 = n53674 & n2803;
  assign n2805 = n53673 & n2804;
  assign n2806 = ~n1471 & n2805;
  assign n2807 = ~n1490 & n2806;
  assign n2808 = ~n247 & n2807;
  assign n2809 = ~n503 & n2808;
  assign n2810 = ~n774 & n2809;
  assign n2811 = ~n740 & n2810;
  assign n2812 = ~n625 & n2811;
  assign n2813 = n53669 & n2801;
  assign n2814 = ~n319 & ~n956;
  assign n2815 = ~n218 & ~n360;
  assign n2816 = n1035 & n2815;
  assign n2817 = n2814 & n2815;
  assign n2818 = n1035 & n2817;
  assign n2819 = n2814 & n2816;
  assign n2820 = ~n504 & ~n832;
  assign n2821 = ~n832 & ~n975;
  assign n2822 = ~n504 & n2821;
  assign n2823 = ~n504 & ~n975;
  assign n2824 = ~n832 & n2823;
  assign n2825 = ~n975 & n2820;
  assign n2826 = ~n631 & ~n753;
  assign n2827 = n276 & n2826;
  assign n2828 = n850 & n1197;
  assign n2829 = n2827 & n2828;
  assign n2830 = n53679 & n2829;
  assign n2831 = n276 & n2814;
  assign n2832 = n850 & n2831;
  assign n2833 = ~n218 & ~n753;
  assign n2834 = ~n360 & ~n631;
  assign n2835 = ~n360 & ~n753;
  assign n2836 = ~n218 & ~n631;
  assign n2837 = n2835 & n2836;
  assign n2838 = n2833 & n2834;
  assign n2839 = n1035 & n1197;
  assign n2840 = n53680 & n2839;
  assign n2841 = n53679 & n2840;
  assign n2842 = n2832 & n2841;
  assign n2843 = n2814 & n2828;
  assign n2844 = n276 & n1035;
  assign n2845 = n53680 & n2844;
  assign n2846 = n53679 & n2845;
  assign n2847 = n2843 & n2846;
  assign n2848 = n53678 & n2830;
  assign n2849 = ~n353 & ~n444;
  assign n2850 = ~n627 & n2849;
  assign n2851 = ~n353 & n1270;
  assign n2852 = ~n409 & ~n822;
  assign n2853 = ~n651 & ~n1703;
  assign n2854 = ~n255 & ~n833;
  assign n2855 = n2853 & n2854;
  assign n2856 = ~n1703 & n2854;
  assign n2857 = ~n822 & n2856;
  assign n2858 = ~n409 & n2857;
  assign n2859 = ~n651 & n2858;
  assign n2860 = n2852 & n2855;
  assign n2861 = ~n627 & n53683;
  assign n2862 = ~n444 & n2861;
  assign n2863 = ~n353 & n2862;
  assign n2864 = ~n353 & ~n651;
  assign n2865 = ~n444 & n2864;
  assign n2866 = ~n409 & ~n627;
  assign n2867 = ~n822 & ~n1703;
  assign n2868 = n2866 & n2867;
  assign n2869 = n2854 & n2868;
  assign n2870 = n2865 & n2869;
  assign n2871 = n53682 & n53683;
  assign n2872 = n53644 & n53684;
  assign n2873 = n53681 & n2872;
  assign n2874 = n53677 & n2873;
  assign n2875 = n53668 & n53677;
  assign n2876 = n2873 & n2875;
  assign n2877 = n2814 & n53679;
  assign n2878 = n53644 & n2877;
  assign n2879 = n53677 & n2878;
  assign n2880 = n53684 & n2879;
  assign n2881 = n1197 & n2880;
  assign n2882 = n1035 & n2881;
  assign n2883 = n53668 & n2882;
  assign n2884 = n850 & n2883;
  assign n2885 = n276 & n2884;
  assign n2886 = ~n631 & n2885;
  assign n2887 = ~n218 & n2886;
  assign n2888 = ~n360 & n2887;
  assign n2889 = ~n753 & n2888;
  assign n2890 = n53668 & n2874;
  assign n2891 = ~n53657 & ~n53685;
  assign n2892 = ~n625 & ~n630;
  assign n2893 = ~n207 & ~n630;
  assign n2894 = ~n625 & n2893;
  assign n2895 = ~n207 & n2892;
  assign n2896 = ~n420 & ~n849;
  assign n2897 = ~n161 & ~n618;
  assign n2898 = ~n1124 & ~n1468;
  assign n2899 = n2897 & n2898;
  assign n2900 = ~n161 & ~n1124;
  assign n2901 = ~n849 & ~n1468;
  assign n2902 = ~n420 & ~n618;
  assign n2903 = n2901 & n2902;
  assign n2904 = n2900 & n2903;
  assign n2905 = n2896 & n2899;
  assign n2906 = ~n1124 & n53686;
  assign n2907 = ~n1468 & n2906;
  assign n2908 = ~n161 & n2907;
  assign n2909 = ~n618 & n2908;
  assign n2910 = ~n849 & n2909;
  assign n2911 = ~n420 & n2910;
  assign n2912 = n53686 & n53687;
  assign n2913 = ~n344 & ~n1191;
  assign n2914 = ~n623 & ~n1680;
  assign n2915 = n2913 & n2914;
  assign n2916 = ~n166 & ~n773;
  assign n2917 = ~n206 & ~n902;
  assign n2918 = n2916 & n2917;
  assign n2919 = n2915 & n2918;
  assign n2920 = ~n349 & ~n1088;
  assign n2921 = ~n268 & n2920;
  assign n2922 = ~n268 & ~n349;
  assign n2923 = ~n1088 & n2922;
  assign n2924 = ~n349 & n1089;
  assign n2925 = ~n246 & ~n614;
  assign n2926 = n2741 & n2925;
  assign n2927 = n53689 & n2926;
  assign n2928 = n2914 & n2925;
  assign n2929 = n2918 & n2928;
  assign n2930 = n2741 & n2913;
  assign n2931 = n53689 & n2930;
  assign n2932 = n2929 & n2931;
  assign n2933 = n1673 & n2917;
  assign n2934 = n2914 & n2916;
  assign n2935 = n2933 & n2934;
  assign n2936 = ~n344 & ~n614;
  assign n2937 = n2741 & n2936;
  assign n2938 = n53689 & n2937;
  assign n2939 = n2935 & n2938;
  assign n2940 = ~n614 & ~n623;
  assign n2941 = n1673 & n2940;
  assign n2942 = n2741 & n2916;
  assign n2943 = n2941 & n2942;
  assign n2944 = ~n344 & ~n1680;
  assign n2945 = n2917 & n2944;
  assign n2946 = n53689 & n2945;
  assign n2947 = n2943 & n2946;
  assign n2948 = n2919 & n2927;
  assign n2949 = ~n1337 & ~n1681;
  assign n2950 = n1035 & ~n1491;
  assign n2951 = n1035 & n2949;
  assign n2952 = ~n1491 & n2951;
  assign n2953 = n2949 & n2950;
  assign n2954 = ~n311 & ~n320;
  assign n2955 = ~n922 & n2954;
  assign n2956 = ~n922 & n2783;
  assign n2957 = ~n320 & n2956;
  assign n2958 = ~n311 & n2957;
  assign n2959 = n2783 & n2955;
  assign n2960 = n53691 & n53692;
  assign n2961 = n53690 & n2960;
  assign n2962 = n2942 & n53691;
  assign n2963 = n53689 & n2962;
  assign n2964 = n53692 & n2963;
  assign n2965 = n53688 & n2964;
  assign n2966 = n1673 & n2965;
  assign n2967 = ~n902 & n2966;
  assign n2968 = ~n1680 & n2967;
  assign n2969 = ~n206 & n2968;
  assign n2970 = ~n344 & n2969;
  assign n2971 = ~n614 & n2970;
  assign n2972 = ~n623 & n2971;
  assign n2973 = n53688 & n2961;
  assign n2974 = ~n259 & ~n879;
  assign n2975 = ~n504 & ~n1997;
  assign n2976 = ~n307 & ~n402;
  assign n2977 = n2975 & n2976;
  assign n2978 = n2974 & n2977;
  assign n2979 = n749 & n1128;
  assign n2980 = ~n249 & ~n1280;
  assign n2981 = ~n848 & ~n1487;
  assign n2982 = n2980 & n2981;
  assign n2983 = n749 & n2980;
  assign n2984 = n1128 & n2981;
  assign n2985 = n2983 & n2984;
  assign n2986 = n2979 & n2982;
  assign n2987 = n2975 & n2984;
  assign n2988 = n749 & n2974;
  assign n2989 = n2976 & n2980;
  assign n2990 = n2988 & n2989;
  assign n2991 = n2987 & n2990;
  assign n2992 = n2978 & n53694;
  assign n2993 = n53459 & n53695;
  assign n2994 = ~n182 & ~n465;
  assign n2995 = ~n881 & ~n975;
  assign n2996 = ~n465 & ~n975;
  assign n2997 = ~n182 & ~n881;
  assign n2998 = n2996 & n2997;
  assign n2999 = n2994 & n2995;
  assign n3000 = ~n612 & ~n883;
  assign n3001 = ~n321 & ~n441;
  assign n3002 = n1467 & n3001;
  assign n3003 = n3000 & n3001;
  assign n3004 = n1467 & n3003;
  assign n3005 = n3000 & n3002;
  assign n3006 = ~n881 & n53697;
  assign n3007 = ~n182 & n3006;
  assign n3008 = ~n975 & n3007;
  assign n3009 = ~n465 & n3008;
  assign n3010 = n53696 & n53697;
  assign n3011 = ~n1125 & n2093;
  assign n3012 = n223 & n497;
  assign n3013 = n3011 & n3012;
  assign n3014 = ~n1065 & ~n1477;
  assign n3015 = n1391 & n3014;
  assign n3016 = ~n622 & ~n740;
  assign n3017 = n358 & ~n740;
  assign n3018 = ~n622 & n3017;
  assign n3019 = n358 & n3016;
  assign n3020 = n3015 & n53699;
  assign n3021 = n3013 & n3020;
  assign n3022 = n53698 & n3021;
  assign n3023 = n3011 & n3015;
  assign n3024 = n53699 & n3023;
  assign n3025 = n497 & n3024;
  assign n3026 = n2981 & n3025;
  assign n3027 = n53698 & n3026;
  assign n3028 = n53459 & n3027;
  assign n3029 = n2974 & n3028;
  assign n3030 = n2975 & n3029;
  assign n3031 = n1128 & n3030;
  assign n3032 = n749 & n3031;
  assign n3033 = ~n307 & n3032;
  assign n3034 = ~n222 & n3033;
  assign n3035 = ~n221 & n3034;
  assign n3036 = ~n249 & n3035;
  assign n3037 = ~n402 & n3036;
  assign n3038 = ~n1280 & n3037;
  assign n3039 = n223 & n2976;
  assign n3040 = n2975 & n3039;
  assign n3041 = n53694 & n3040;
  assign n3042 = n53459 & n3041;
  assign n3043 = n497 & n2974;
  assign n3044 = n3011 & n3043;
  assign n3045 = n3020 & n3044;
  assign n3046 = n53698 & n3045;
  assign n3047 = n3042 & n3046;
  assign n3048 = n497 & n1128;
  assign n3049 = n2974 & n3048;
  assign n3050 = n2975 & n2980;
  assign n3051 = n749 & n2981;
  assign n3052 = n3050 & n3051;
  assign n3053 = n3049 & n3052;
  assign n3054 = n53459 & n3053;
  assign n3055 = n3011 & n3039;
  assign n3056 = n3020 & n3055;
  assign n3057 = n53698 & n3056;
  assign n3058 = n3054 & n3057;
  assign n3059 = n2993 & n3022;
  assign n3060 = n53693 & n53700;
  assign n3061 = n406 & n1197;
  assign n3062 = ~n112 & ~n914;
  assign n3063 = n2772 & n3062;
  assign n3064 = n3061 & n3063;
  assign n3065 = ~n354 & ~n631;
  assign n3066 = ~n342 & ~n733;
  assign n3067 = ~n631 & ~n733;
  assign n3068 = ~n342 & ~n354;
  assign n3069 = n3067 & n3068;
  assign n3070 = n3065 & n3066;
  assign n3071 = n53566 & n53701;
  assign n3072 = n3064 & n3071;
  assign n3073 = ~n172 & ~n498;
  assign n3074 = ~n274 & n2693;
  assign n3075 = ~n172 & n2693;
  assign n3076 = ~n274 & n3075;
  assign n3077 = ~n498 & n3076;
  assign n3078 = ~n172 & ~n274;
  assign n3079 = ~n498 & n3078;
  assign n3080 = n2693 & n3079;
  assign n3081 = n3073 & n3074;
  assign n3082 = ~n663 & ~n776;
  assign n3083 = ~n788 & ~n829;
  assign n3084 = n3082 & n3083;
  assign n3085 = ~n911 & ~n1646;
  assign n3086 = ~n108 & ~n423;
  assign n3087 = n3085 & n3086;
  assign n3088 = n3084 & n3087;
  assign n3089 = n53702 & n3088;
  assign n3090 = n2772 & n3085;
  assign n3091 = n3061 & n3090;
  assign n3092 = n3071 & n3091;
  assign n3093 = n3062 & n3083;
  assign n3094 = n3082 & n3086;
  assign n3095 = n3093 & n3094;
  assign n3096 = n53702 & n3095;
  assign n3097 = n3092 & n3096;
  assign n3098 = ~n342 & ~n451;
  assign n3099 = n1197 & n3098;
  assign n3100 = n406 & n3086;
  assign n3101 = n3099 & n3100;
  assign n3102 = ~n354 & ~n664;
  assign n3103 = n3067 & n3102;
  assign n3104 = n53566 & n3103;
  assign n3105 = n3101 & n3104;
  assign n3106 = n3062 & n3085;
  assign n3107 = n3084 & n3106;
  assign n3108 = n53702 & n3107;
  assign n3109 = n3105 & n3108;
  assign n3110 = ~n664 & ~n733;
  assign n3111 = n3083 & n3110;
  assign n3112 = n3082 & n3085;
  assign n3113 = n3111 & n3112;
  assign n3114 = ~n354 & ~n451;
  assign n3115 = ~n342 & ~n631;
  assign n3116 = n3114 & n3115;
  assign n3117 = n53566 & n3116;
  assign n3118 = n3113 & n3117;
  assign n3119 = n406 & n3062;
  assign n3120 = n1197 & n3086;
  assign n3121 = n3119 & n3120;
  assign n3122 = n53702 & n3121;
  assign n3123 = n3118 & n3122;
  assign n3124 = n3072 & n3089;
  assign n3125 = ~n105 & ~n443;
  assign n3126 = ~n491 & ~n824;
  assign n3127 = ~n443 & ~n491;
  assign n3128 = ~n105 & ~n824;
  assign n3129 = n3127 & n3128;
  assign n3130 = ~n105 & ~n491;
  assign n3131 = ~n443 & ~n824;
  assign n3132 = n3130 & n3131;
  assign n3133 = n3125 & n3126;
  assign n3134 = ~n401 & ~n447;
  assign n3135 = n2400 & n3134;
  assign n3136 = n2400 & n3126;
  assign n3137 = n3125 & n3134;
  assign n3138 = n3136 & n3137;
  assign n3139 = n53704 & n3135;
  assign n3140 = ~n177 & ~n450;
  assign n3141 = ~n177 & ~n948;
  assign n3142 = ~n450 & n3141;
  assign n3143 = ~n450 & ~n948;
  assign n3144 = ~n177 & n3143;
  assign n3145 = ~n948 & n3140;
  assign n3146 = ~n141 & ~n275;
  assign n3147 = ~n141 & ~n184;
  assign n3148 = ~n275 & n3147;
  assign n3149 = ~n184 & ~n275;
  assign n3150 = ~n141 & n3149;
  assign n3151 = ~n184 & n3146;
  assign n3152 = n53706 & n53707;
  assign n3153 = n3134 & n3152;
  assign n3154 = ~n1033 & n3153;
  assign n3155 = ~n1044 & n3154;
  assign n3156 = ~n105 & n3155;
  assign n3157 = ~n824 & n3156;
  assign n3158 = ~n443 & n3157;
  assign n3159 = ~n491 & n3158;
  assign n3160 = n53705 & n3152;
  assign n3161 = ~n440 & ~n741;
  assign n3162 = ~n741 & ~n2201;
  assign n3163 = ~n440 & n3162;
  assign n3164 = ~n2201 & n3161;
  assign n3165 = ~n410 & ~n851;
  assign n3166 = ~n348 & ~n611;
  assign n3167 = n755 & n3166;
  assign n3168 = n3165 & n3166;
  assign n3169 = n755 & n3168;
  assign n3170 = n3165 & n3167;
  assign n3171 = n755 & n3165;
  assign n3172 = ~n440 & n3171;
  assign n3173 = ~n611 & n3172;
  assign n3174 = ~n348 & n3173;
  assign n3175 = ~n741 & n3174;
  assign n3176 = ~n2201 & n3175;
  assign n3177 = ~n611 & ~n741;
  assign n3178 = ~n2201 & n3177;
  assign n3179 = ~n348 & ~n440;
  assign n3180 = n755 & n3179;
  assign n3181 = n3165 & n3180;
  assign n3182 = n3178 & n3181;
  assign n3183 = ~n440 & ~n2201;
  assign n3184 = ~n611 & n3183;
  assign n3185 = ~n348 & ~n741;
  assign n3186 = n755 & n3185;
  assign n3187 = n3165 & n3186;
  assign n3188 = n3184 & n3187;
  assign n3189 = n53709 & n53710;
  assign n3190 = n53708 & n53711;
  assign n3191 = n53703 & n3190;
  assign n3192 = n53566 & n3083;
  assign n3193 = n53702 & n3192;
  assign n3194 = n53711 & n3193;
  assign n3195 = n53700 & n3194;
  assign n3196 = n53693 & n3195;
  assign n3197 = n1197 & n3196;
  assign n3198 = n53708 & n3197;
  assign n3199 = n3085 & n3198;
  assign n3200 = n3086 & n3199;
  assign n3201 = n3082 & n3200;
  assign n3202 = n406 & n3201;
  assign n3203 = n3062 & n3202;
  assign n3204 = ~n631 & n3203;
  assign n3205 = ~n664 & n3204;
  assign n3206 = ~n733 & n3205;
  assign n3207 = ~n451 & n3206;
  assign n3208 = ~n354 & n3207;
  assign n3209 = ~n342 & n3208;
  assign n3210 = n53693 & n3191;
  assign n3211 = n53700 & n3210;
  assign n3212 = n3060 & n3191;
  assign n3213 = ~n53685 & ~n53712;
  assign n3214 = ~n751 & ~n894;
  assign n3215 = ~n750 & n3214;
  assign n3216 = n752 & ~n894;
  assign n3217 = ~n742 & ~n1769;
  assign n3218 = ~n741 & ~n896;
  assign n3219 = n3217 & n3218;
  assign n3220 = n3214 & n3217;
  assign n3221 = ~n896 & n3220;
  assign n3222 = ~n741 & n3221;
  assign n3223 = ~n750 & n3222;
  assign n3224 = ~n750 & n3218;
  assign n3225 = n3220 & n3224;
  assign n3226 = n53713 & n3219;
  assign n3227 = ~n914 & ~n1641;
  assign n3228 = ~n922 & ~n1059;
  assign n3229 = ~n922 & ~n1641;
  assign n3230 = ~n914 & ~n1059;
  assign n3231 = n3229 & n3230;
  assign n3232 = n3227 & n3228;
  assign n3233 = ~n168 & ~n405;
  assign n3234 = n3014 & n3233;
  assign n3235 = ~n922 & n3014;
  assign n3236 = ~n168 & n3235;
  assign n3237 = ~n405 & n3236;
  assign n3238 = ~n1059 & n3237;
  assign n3239 = ~n914 & n3238;
  assign n3240 = ~n1641 & n3239;
  assign n3241 = ~n168 & ~n1059;
  assign n3242 = n3229 & n3241;
  assign n3243 = ~n405 & ~n914;
  assign n3244 = n3014 & n3243;
  assign n3245 = n3242 & n3244;
  assign n3246 = ~n914 & ~n922;
  assign n3247 = n3233 & n3246;
  assign n3248 = ~n1059 & ~n1641;
  assign n3249 = n3014 & n3248;
  assign n3250 = n3247 & n3249;
  assign n3251 = n53715 & n3234;
  assign n3252 = ~n174 & ~n788;
  assign n3253 = ~n101 & ~n222;
  assign n3254 = n3252 & n3253;
  assign n3255 = ~n849 & ~n1680;
  assign n3256 = ~n776 & ~n1031;
  assign n3257 = n3255 & n3256;
  assign n3258 = n3254 & n3257;
  assign n3259 = n53716 & n3258;
  assign n3260 = n53714 & n3259;
  assign n3261 = ~n340 & ~n823;
  assign n3262 = ~n1715 & n3261;
  assign n3263 = ~n211 & ~n271;
  assign n3264 = ~n246 & ~n1085;
  assign n3265 = ~n211 & ~n1085;
  assign n3266 = ~n246 & ~n271;
  assign n3267 = n3265 & n3266;
  assign n3268 = ~n271 & ~n1085;
  assign n3269 = ~n211 & ~n246;
  assign n3270 = n3268 & n3269;
  assign n3271 = n3263 & n3264;
  assign n3272 = ~n401 & ~n1124;
  assign n3273 = ~n182 & ~n249;
  assign n3274 = n3272 & n3273;
  assign n3275 = n53717 & n3274;
  assign n3276 = n3262 & n3272;
  assign n3277 = n3273 & n3276;
  assign n3278 = ~n1085 & n3277;
  assign n3279 = ~n211 & n3278;
  assign n3280 = ~n271 & n3279;
  assign n3281 = ~n246 & n3280;
  assign n3282 = n3262 & n3275;
  assign n3283 = ~n957 & ~n1469;
  assign n3284 = ~n259 & ~n357;
  assign n3285 = ~n259 & n3283;
  assign n3286 = ~n357 & n3285;
  assign n3287 = n3283 & n3284;
  assign n3288 = ~n296 & ~n851;
  assign n3289 = ~n1192 & ~n1485;
  assign n3290 = ~n296 & ~n1192;
  assign n3291 = ~n1485 & n3290;
  assign n3292 = ~n851 & n3291;
  assign n3293 = ~n851 & ~n1485;
  assign n3294 = n3290 & n3293;
  assign n3295 = n3288 & n3289;
  assign n3296 = ~n346 & ~n451;
  assign n3297 = ~n1478 & n3296;
  assign n3298 = n53720 & n3297;
  assign n3299 = n53719 & n3298;
  assign n3300 = n53718 & n3299;
  assign n3301 = ~n346 & ~n1031;
  assign n3302 = n3252 & n3301;
  assign n3303 = ~n451 & ~n776;
  assign n3304 = n3255 & n3303;
  assign n3305 = n3255 & n3296;
  assign n3306 = n3252 & n3256;
  assign n3307 = n3305 & n3306;
  assign n3308 = n3302 & n3304;
  assign n3309 = n53714 & n53721;
  assign n3310 = n53716 & n53721;
  assign n3311 = n53714 & n3310;
  assign n3312 = n53716 & n3309;
  assign n3313 = ~n1478 & n3253;
  assign n3314 = n53720 & n3313;
  assign n3315 = n53719 & n3314;
  assign n3316 = n53718 & n3315;
  assign n3317 = n53722 & n3316;
  assign n3318 = ~n849 & ~n1031;
  assign n3319 = n3303 & n3318;
  assign n3320 = ~n101 & ~n174;
  assign n3321 = ~n788 & ~n1680;
  assign n3322 = n3320 & n3321;
  assign n3323 = n3319 & n3322;
  assign n3324 = n53716 & n3323;
  assign n3325 = n53714 & n3324;
  assign n3326 = ~n346 & ~n1478;
  assign n3327 = ~n222 & n3326;
  assign n3328 = n53720 & n3327;
  assign n3329 = n53719 & n3328;
  assign n3330 = n53718 & n3329;
  assign n3331 = n3325 & n3330;
  assign n3332 = n3260 & n3300;
  assign n3333 = n53485 & n53723;
  assign n3334 = ~n460 & ~n1196;
  assign n3335 = ~n291 & ~n409;
  assign n3336 = n1235 & n3335;
  assign n3337 = n1235 & n3334;
  assign n3338 = n3335 & n3337;
  assign n3339 = n3334 & n3336;
  assign n3340 = ~n308 & ~n559;
  assign n3341 = ~n308 & ~n514;
  assign n3342 = ~n559 & n3341;
  assign n3343 = ~n514 & ~n559;
  assign n3344 = ~n308 & n3343;
  assign n3345 = ~n514 & n3340;
  assign n3346 = ~n511 & ~n748;
  assign n3347 = ~n1472 & n3346;
  assign n3348 = n53725 & n3347;
  assign n3349 = n3334 & n53725;
  assign n3350 = ~n291 & n3349;
  assign n3351 = ~n1472 & n3350;
  assign n3352 = ~n1234 & n3351;
  assign n3353 = ~n830 & n3352;
  assign n3354 = ~n748 & n3353;
  assign n3355 = ~n511 & n3354;
  assign n3356 = ~n409 & n3355;
  assign n3357 = ~n409 & ~n1472;
  assign n3358 = ~n291 & ~n1234;
  assign n3359 = ~n1234 & ~n1472;
  assign n3360 = n3335 & n3359;
  assign n3361 = n3357 & n3358;
  assign n3362 = n3334 & n53727;
  assign n3363 = ~n511 & ~n830;
  assign n3364 = ~n748 & n3363;
  assign n3365 = ~n830 & n3346;
  assign n3366 = n53725 & n53728;
  assign n3367 = n3362 & n3366;
  assign n3368 = n53724 & n3348;
  assign n3369 = ~n402 & ~n822;
  assign n3370 = n2476 & n3369;
  assign n3371 = ~n163 & n421;
  assign n3372 = ~n1492 & ~n1681;
  assign n3373 = ~n1195 & n3372;
  assign n3374 = n3371 & n3373;
  assign n3375 = n3370 & n3373;
  assign n3376 = n3371 & n3375;
  assign n3377 = n3370 & n3374;
  assign n3378 = ~n1090 & ~n2042;
  assign n3379 = ~n1033 & ~n1476;
  assign n3380 = n3378 & n3379;
  assign n3381 = ~n1033 & n1642;
  assign n3382 = ~n1090 & n3381;
  assign n3383 = ~n1476 & n3382;
  assign n3384 = ~n2042 & n3383;
  assign n3385 = n1642 & n3380;
  assign n3386 = ~n250 & ~n504;
  assign n3387 = ~n824 & ~n1634;
  assign n3388 = n3386 & n3387;
  assign n3389 = ~n258 & ~n320;
  assign n3390 = ~n207 & ~n219;
  assign n3391 = n3389 & n3390;
  assign n3392 = ~n207 & ~n250;
  assign n3393 = n3387 & n3392;
  assign n3394 = ~n219 & ~n504;
  assign n3395 = n3389 & n3394;
  assign n3396 = n3393 & n3395;
  assign n3397 = n3388 & n3391;
  assign n3398 = n53730 & n53731;
  assign n3399 = ~n1492 & n3387;
  assign n3400 = n3371 & n3399;
  assign n3401 = n3370 & n3400;
  assign n3402 = ~n250 & ~n1681;
  assign n3403 = ~n504 & ~n1195;
  assign n3404 = n3402 & n3403;
  assign n3405 = n3391 & n3404;
  assign n3406 = n53730 & n3405;
  assign n3407 = n3401 & n3406;
  assign n3408 = ~n207 & ~n1195;
  assign n3409 = ~n1681 & n3408;
  assign n3410 = ~n250 & ~n824;
  assign n3411 = ~n219 & ~n1492;
  assign n3412 = n3410 & n3411;
  assign n3413 = n3409 & n3412;
  assign n3414 = n3371 & n3413;
  assign n3415 = ~n504 & ~n1634;
  assign n3416 = n3389 & n3415;
  assign n3417 = n3370 & n3416;
  assign n3418 = n53730 & n3417;
  assign n3419 = n3414 & n3418;
  assign n3420 = n53729 & n3398;
  assign n3421 = n3369 & n3371;
  assign n3422 = n53730 & n3421;
  assign n3423 = n53726 & n3422;
  assign n3424 = n2476 & n3423;
  assign n3425 = n3389 & n3424;
  assign n3426 = ~n1681 & n3425;
  assign n3427 = ~n1195 & n3426;
  assign n3428 = ~n1492 & n3427;
  assign n3429 = ~n219 & n3428;
  assign n3430 = ~n250 & n3429;
  assign n3431 = ~n207 & n3430;
  assign n3432 = ~n824 & n3431;
  assign n3433 = ~n504 & n3432;
  assign n3434 = ~n1634 & n3433;
  assign n3435 = n53726 & n53732;
  assign n3436 = ~n404 & ~n777;
  assign n3437 = ~n404 & ~n948;
  assign n3438 = ~n777 & n3437;
  assign n3439 = ~n948 & n3436;
  assign n3440 = ~n179 & ~n423;
  assign n3441 = ~n179 & ~n1062;
  assign n3442 = ~n423 & n3441;
  assign n3443 = ~n423 & ~n1062;
  assign n3444 = ~n179 & n3443;
  assign n3445 = ~n1062 & n3440;
  assign n3446 = n318 & n1273;
  assign n3447 = n53735 & n3446;
  assign n3448 = n53734 & n3447;
  assign n3449 = ~n349 & ~n507;
  assign n3450 = ~n789 & ~n1644;
  assign n3451 = ~n1997 & n3450;
  assign n3452 = ~n1644 & ~n1997;
  assign n3453 = ~n507 & n3452;
  assign n3454 = ~n349 & n3453;
  assign n3455 = ~n789 & n3454;
  assign n3456 = ~n507 & ~n1644;
  assign n3457 = ~n349 & ~n1997;
  assign n3458 = ~n789 & n3457;
  assign n3459 = n3456 & n3458;
  assign n3460 = ~n789 & n3449;
  assign n3461 = n3452 & n3460;
  assign n3462 = n3449 & n3451;
  assign n3463 = ~n274 & ~n1280;
  assign n3464 = ~n206 & ~n295;
  assign n3465 = ~n295 & ~n440;
  assign n3466 = ~n206 & n3465;
  assign n3467 = ~n206 & ~n440;
  assign n3468 = ~n295 & n3467;
  assign n3469 = ~n440 & n3464;
  assign n3470 = ~n295 & n3463;
  assign n3471 = ~n206 & n3470;
  assign n3472 = ~n440 & n3471;
  assign n3473 = n3463 & n53737;
  assign n3474 = ~n221 & ~n348;
  assign n3475 = ~n447 & ~n983;
  assign n3476 = ~n144 & ~n247;
  assign n3477 = n3475 & n3476;
  assign n3478 = n3474 & n3475;
  assign n3479 = n3476 & n3478;
  assign n3480 = n3474 & n3477;
  assign n3481 = n53738 & n53739;
  assign n3482 = n53736 & n3481;
  assign n3483 = n53734 & n3474;
  assign n3484 = n53736 & n3483;
  assign n3485 = n53738 & n3484;
  assign n3486 = n1273 & n3485;
  assign n3487 = n3476 & n3486;
  assign n3488 = n3475 & n3487;
  assign n3489 = n318 & n3488;
  assign n3490 = ~n1062 & n3489;
  assign n3491 = ~n179 & n3490;
  assign n3492 = ~n423 & n3491;
  assign n3493 = n1273 & n3476;
  assign n3494 = n53735 & n3493;
  assign n3495 = n53734 & n3494;
  assign n3496 = n318 & n3478;
  assign n3497 = n53738 & n3496;
  assign n3498 = n53736 & n3497;
  assign n3499 = n3495 & n3498;
  assign n3500 = n3448 & n3482;
  assign n3501 = n53733 & n53740;
  assign n3502 = n53714 & n53719;
  assign n3503 = n53485 & n3502;
  assign n3504 = n53720 & n3503;
  assign n3505 = n53716 & n3504;
  assign n3506 = n53733 & n3505;
  assign n3507 = n53718 & n3506;
  assign n3508 = n53740 & n3507;
  assign n3509 = ~n1031 & n3508;
  assign n3510 = ~n1680 & n3509;
  assign n3511 = ~n1478 & n3510;
  assign n3512 = ~n174 & n3511;
  assign n3513 = ~n101 & n3512;
  assign n3514 = ~n222 & n3513;
  assign n3515 = ~n849 & n3514;
  assign n3516 = ~n451 & n3515;
  assign n3517 = ~n788 & n3516;
  assign n3518 = ~n776 & n3517;
  assign n3519 = ~n346 & n3518;
  assign n3520 = n3333 & n3501;
  assign n3521 = ~n53712 & ~n53741;
  assign n3522 = ~n168 & ~n461;
  assign n3523 = ~n250 & ~n354;
  assign n3524 = n3522 & n3523;
  assign n3525 = ~n108 & ~n506;
  assign n3526 = n589 & n3525;
  assign n3527 = n3524 & n3526;
  assign n3528 = n1673 & n3463;
  assign n3529 = ~n317 & ~n356;
  assign n3530 = ~n902 & ~n1061;
  assign n3531 = ~n356 & ~n1061;
  assign n3532 = ~n317 & ~n902;
  assign n3533 = n3531 & n3532;
  assign n3534 = n3529 & n3530;
  assign n3535 = ~n511 & ~n1455;
  assign n3536 = ~n590 & ~n1088;
  assign n3537 = n3535 & n3536;
  assign n3538 = n53742 & n3537;
  assign n3539 = n3528 & n3538;
  assign n3540 = n3524 & n3537;
  assign n3541 = n3526 & n53742;
  assign n3542 = n3528 & n3541;
  assign n3543 = n3540 & n3542;
  assign n3544 = n3523 & n3535;
  assign n3545 = n589 & n3522;
  assign n3546 = n3544 & n3545;
  assign n3547 = n3525 & n3536;
  assign n3548 = n3528 & n3547;
  assign n3549 = n53742 & n3548;
  assign n3550 = n3546 & n3549;
  assign n3551 = n3463 & n3535;
  assign n3552 = n3522 & n3525;
  assign n3553 = n3551 & n3552;
  assign n3554 = n1673 & n3523;
  assign n3555 = n589 & n3536;
  assign n3556 = n3554 & n3555;
  assign n3557 = n53742 & n3556;
  assign n3558 = n3553 & n3557;
  assign n3559 = n3527 & n3539;
  assign n3560 = ~n166 & ~n1490;
  assign n3561 = ~n660 & ~n750;
  assign n3562 = ~n491 & ~n833;
  assign n3563 = n3561 & n3562;
  assign n3564 = n3560 & n3563;
  assign n3565 = ~n321 & ~n357;
  assign n3566 = ~n852 & n3565;
  assign n3567 = ~n627 & ~n647;
  assign n3568 = n500 & n3567;
  assign n3569 = ~n321 & ~n647;
  assign n3570 = ~n852 & n3569;
  assign n3571 = ~n357 & ~n627;
  assign n3572 = n500 & n3571;
  assign n3573 = n3570 & n3572;
  assign n3574 = n3566 & n3568;
  assign n3575 = n500 & n3561;
  assign n3576 = ~n1490 & n3575;
  assign n3577 = ~n321 & n3576;
  assign n3578 = ~n166 & n3577;
  assign n3579 = ~n833 & n3578;
  assign n3580 = ~n852 & n3579;
  assign n3581 = ~n491 & n3580;
  assign n3582 = ~n357 & n3581;
  assign n3583 = ~n647 & n3582;
  assign n3584 = ~n627 & n3583;
  assign n3585 = n500 & n3560;
  assign n3586 = n3562 & n3585;
  assign n3587 = ~n627 & n3565;
  assign n3588 = ~n647 & ~n852;
  assign n3589 = n3561 & n3588;
  assign n3590 = n3587 & n3589;
  assign n3591 = n3586 & n3590;
  assign n3592 = n3561 & n3567;
  assign n3593 = n500 & n3592;
  assign n3594 = ~n166 & ~n357;
  assign n3595 = ~n321 & n3594;
  assign n3596 = ~n852 & ~n1490;
  assign n3597 = n3562 & n3596;
  assign n3598 = n3595 & n3597;
  assign n3599 = n3593 & n3598;
  assign n3600 = n3564 & n53744;
  assign n3601 = ~n402 & ~n664;
  assign n3602 = ~n664 & ~n983;
  assign n3603 = ~n402 & n3602;
  assign n3604 = ~n983 & n3601;
  assign n3605 = n755 & n2690;
  assign n3606 = ~n649 & ~n957;
  assign n3607 = ~n221 & ~n422;
  assign n3608 = n3606 & n3607;
  assign n3609 = n2690 & n3606;
  assign n3610 = n755 & n3607;
  assign n3611 = n3609 & n3610;
  assign n3612 = n3605 & n3608;
  assign n3613 = n2690 & n3607;
  assign n3614 = n755 & n3613;
  assign n3615 = ~n957 & n3614;
  assign n3616 = ~n983 & n3615;
  assign n3617 = ~n664 & n3616;
  assign n3618 = ~n402 & n3617;
  assign n3619 = ~n649 & n3618;
  assign n3620 = n53746 & n53747;
  assign n3621 = n53745 & n53748;
  assign n3622 = n589 & n3523;
  assign n3623 = n3522 & n3622;
  assign n3624 = n3463 & n3623;
  assign n3625 = n53748 & n3624;
  assign n3626 = n53745 & n3625;
  assign n3627 = n3535 & n3626;
  assign n3628 = n1673 & n3627;
  assign n3629 = n3536 & n3628;
  assign n3630 = ~n902 & n3629;
  assign n3631 = ~n1061 & n3630;
  assign n3632 = ~n317 & n3631;
  assign n3633 = n3525 & n3632;
  assign n3634 = ~n356 & n3633;
  assign n3635 = n53743 & n3621;
  assign n3636 = ~n460 & ~n612;
  assign n3637 = ~n1646 & n3636;
  assign n3638 = ~n894 & ~n1196;
  assign n3639 = ~n741 & ~n1044;
  assign n3640 = n3638 & n3639;
  assign n3641 = ~n894 & ~n1646;
  assign n3642 = ~n612 & ~n1646;
  assign n3643 = ~n894 & n3642;
  assign n3644 = ~n612 & ~n894;
  assign n3645 = ~n1646 & n3644;
  assign n3646 = ~n612 & n3641;
  assign n3647 = n3334 & n3639;
  assign n3648 = n53750 & n3647;
  assign n3649 = n3637 & n3640;
  assign n3650 = ~n184 & ~n1042;
  assign n3651 = ~n184 & n799;
  assign n3652 = ~n1042 & n3651;
  assign n3653 = n799 & n3650;
  assign n3654 = ~n141 & ~n565;
  assign n3655 = ~n565 & ~n1469;
  assign n3656 = ~n141 & n3655;
  assign n3657 = ~n141 & ~n1469;
  assign n3658 = ~n565 & n3657;
  assign n3659 = ~n1469 & n3654;
  assign n3660 = n53752 & n53753;
  assign n3661 = n53751 & n3660;
  assign n3662 = n3334 & n53752;
  assign n3663 = n53753 & n3662;
  assign n3664 = n3639 & n3663;
  assign n3665 = n53749 & n3664;
  assign n3666 = ~n894 & n3665;
  assign n3667 = ~n612 & n3666;
  assign n3668 = ~n1646 & n3667;
  assign n3669 = n53749 & n3661;
  assign n3670 = ~n823 & ~n1634;
  assign n3671 = ~n308 & ~n1031;
  assign n3672 = ~n789 & ~n1059;
  assign n3673 = n3671 & n3672;
  assign n3674 = n3670 & n3673;
  assign n3675 = ~n567 & ~n1195;
  assign n3676 = ~n144 & ~n553;
  assign n3677 = n3675 & n3676;
  assign n3678 = ~n271 & ~n444;
  assign n3679 = n2256 & n3678;
  assign n3680 = n3677 & n3679;
  assign n3681 = ~n401 & ~n464;
  assign n3682 = n2691 & n3681;
  assign n3683 = ~n401 & ~n748;
  assign n3684 = ~n464 & n3683;
  assign n3685 = ~n748 & n3681;
  assign n3686 = n1541 & n2691;
  assign n3687 = n53755 & n3686;
  assign n3688 = n2566 & n3682;
  assign n3689 = n3680 & n53756;
  assign n3690 = n3672 & n3676;
  assign n3691 = n3671 & n3690;
  assign n3692 = n3675 & n3678;
  assign n3693 = n2256 & n3670;
  assign n3694 = n3692 & n3693;
  assign n3695 = n53756 & n3694;
  assign n3696 = n3691 & n3695;
  assign n3697 = n3676 & n3679;
  assign n3698 = n3672 & n3675;
  assign n3699 = n3670 & n3671;
  assign n3700 = n3698 & n3699;
  assign n3701 = n53756 & n3700;
  assign n3702 = n3697 & n3701;
  assign n3703 = n2691 & n3671;
  assign n3704 = n3676 & n3703;
  assign n3705 = n1541 & n3670;
  assign n3706 = n3698 & n3705;
  assign n3707 = n3679 & n53755;
  assign n3708 = n3706 & n3707;
  assign n3709 = n3704 & n3708;
  assign n3710 = n3674 & n3689;
  assign n3711 = ~n423 & ~n493;
  assign n3712 = ~n423 & ~n1457;
  assign n3713 = ~n493 & n3712;
  assign n3714 = ~n1457 & n3711;
  assign n3715 = ~n622 & ~n1486;
  assign n3716 = ~n1472 & ~n1644;
  assign n3717 = ~n174 & ~n646;
  assign n3718 = n3716 & n3717;
  assign n3719 = n3715 & n3718;
  assign n3720 = n3715 & n3716;
  assign n3721 = ~n174 & n3720;
  assign n3722 = ~n1457 & n3721;
  assign n3723 = ~n493 & n3722;
  assign n3724 = ~n423 & n3723;
  assign n3725 = ~n646 & n3724;
  assign n3726 = ~n174 & ~n423;
  assign n3727 = ~n1457 & n3726;
  assign n3728 = ~n493 & ~n646;
  assign n3729 = n3715 & n3728;
  assign n3730 = n3716 & n3729;
  assign n3731 = n3727 & n3730;
  assign n3732 = ~n1457 & n3728;
  assign n3733 = n3716 & n3726;
  assign n3734 = n3715 & n3733;
  assign n3735 = n3732 & n3734;
  assign n3736 = n53758 & n3719;
  assign n3737 = ~n101 & ~n1997;
  assign n3738 = ~n319 & ~n495;
  assign n3739 = ~n495 & n3737;
  assign n3740 = ~n319 & n3739;
  assign n3741 = n3737 & n3738;
  assign n3742 = ~n311 & ~n1085;
  assign n3743 = ~n651 & ~n948;
  assign n3744 = ~n948 & n3742;
  assign n3745 = ~n651 & n3744;
  assign n3746 = n3742 & n3743;
  assign n3747 = ~n296 & ~n618;
  assign n3748 = ~n296 & ~n320;
  assign n3749 = ~n618 & n3748;
  assign n3750 = ~n320 & ~n618;
  assign n3751 = ~n296 & n3750;
  assign n3752 = ~n320 & n3747;
  assign n3753 = n53761 & n53762;
  assign n3754 = n53760 & n53761;
  assign n3755 = n53762 & n3754;
  assign n3756 = n53760 & n53762;
  assign n3757 = n53761 & n3756;
  assign n3758 = n53760 & n3753;
  assign n3759 = n53759 & n53763;
  assign n3760 = n3676 & n53762;
  assign n3761 = n53761 & n3760;
  assign n3762 = n2691 & n3761;
  assign n3763 = n2256 & n3762;
  assign n3764 = n3678 & n3763;
  assign n3765 = n3671 & n3764;
  assign n3766 = n53760 & n3765;
  assign n3767 = n3675 & n3766;
  assign n3768 = n1541 & n3767;
  assign n3769 = n53759 & n3768;
  assign n3770 = n3670 & n3769;
  assign n3771 = n3672 & n3770;
  assign n3772 = ~n464 & n3771;
  assign n3773 = ~n401 & n3772;
  assign n3774 = ~n748 & n3773;
  assign n3775 = n53757 & n3759;
  assign n3776 = ~n212 & ~n1912;
  assign n3777 = ~n212 & n2338;
  assign n3778 = ~n901 & n3776;
  assign n3779 = n1675 & n53765;
  assign n3780 = ~n568 & ~n1337;
  assign n3781 = ~n822 & ~n2109;
  assign n3782 = ~n822 & n3780;
  assign n3783 = ~n2109 & n3782;
  assign n3784 = n3780 & n3781;
  assign n3785 = ~n206 & ~n631;
  assign n3786 = ~n161 & ~n269;
  assign n3787 = ~n161 & ~n631;
  assign n3788 = ~n206 & n3787;
  assign n3789 = ~n269 & n3788;
  assign n3790 = ~n161 & ~n206;
  assign n3791 = ~n269 & ~n631;
  assign n3792 = n3790 & n3791;
  assign n3793 = n3785 & n3786;
  assign n3794 = n53766 & n53767;
  assign n3795 = n1675 & n53767;
  assign n3796 = n53765 & n53766;
  assign n3797 = n3795 & n3796;
  assign n3798 = n3779 & n3794;
  assign n3799 = ~n450 & ~n630;
  assign n3800 = ~n1466 & n3799;
  assign n3801 = ~n740 & ~n777;
  assign n3802 = ~n465 & ~n1189;
  assign n3803 = n3801 & n3802;
  assign n3804 = ~n1466 & n3801;
  assign n3805 = ~n1189 & n3804;
  assign n3806 = ~n630 & n3805;
  assign n3807 = ~n465 & n3806;
  assign n3808 = ~n450 & n3807;
  assign n3809 = ~n465 & ~n1466;
  assign n3810 = ~n1189 & n3809;
  assign n3811 = n3799 & n3801;
  assign n3812 = n3810 & n3811;
  assign n3813 = ~n465 & ~n630;
  assign n3814 = ~n1189 & n3813;
  assign n3815 = ~n450 & ~n1466;
  assign n3816 = n3801 & n3815;
  assign n3817 = n3814 & n3816;
  assign n3818 = n3800 & n3803;
  assign n3819 = ~n364 & ~n404;
  assign n3820 = n2974 & n3819;
  assign n3821 = ~n349 & ~n956;
  assign n3822 = n2058 & n3821;
  assign n3823 = n2974 & n3821;
  assign n3824 = n2058 & n3819;
  assign n3825 = n3823 & n3824;
  assign n3826 = n2058 & n2974;
  assign n3827 = n3819 & n3821;
  assign n3828 = n3826 & n3827;
  assign n3829 = n3820 & n3822;
  assign n3830 = ~n307 & ~n615;
  assign n3831 = ~n307 & ~n824;
  assign n3832 = ~n615 & n3831;
  assign n3833 = ~n824 & n3830;
  assign n3834 = ~n179 & ~n650;
  assign n3835 = ~n771 & ~n1535;
  assign n3836 = ~n650 & ~n1535;
  assign n3837 = ~n179 & ~n771;
  assign n3838 = n3836 & n3837;
  assign n3839 = n3834 & n3835;
  assign n3840 = n53771 & n53772;
  assign n3841 = n53770 & n3840;
  assign n3842 = n53769 & n3841;
  assign n3843 = n53765 & n53771;
  assign n3844 = n1675 & n53766;
  assign n3845 = n3843 & n3844;
  assign n3846 = n53767 & n53772;
  assign n3847 = n53770 & n3846;
  assign n3848 = n53769 & n3847;
  assign n3849 = n3845 & n3848;
  assign n3850 = n53766 & n53771;
  assign n3851 = n3795 & n3850;
  assign n3852 = ~n179 & n3836;
  assign n3853 = n1186 & n2338;
  assign n3854 = n3852 & n3853;
  assign n3855 = n53770 & n3854;
  assign n3856 = n53769 & n3855;
  assign n3857 = n3851 & n3856;
  assign n3858 = n53768 & n3842;
  assign n3859 = n53764 & n53773;
  assign n3860 = n53766 & n3821;
  assign n3861 = n53771 & n3860;
  assign n3862 = n1186 & n3861;
  assign n3863 = n3819 & n3862;
  assign n3864 = n53767 & n3863;
  assign n3865 = n53754 & n3864;
  assign n3866 = n53764 & n3865;
  assign n3867 = n53769 & n3866;
  assign n3868 = n1675 & n3867;
  assign n3869 = n2974 & n3868;
  assign n3870 = n2338 & n3869;
  assign n3871 = n2058 & n3870;
  assign n3872 = ~n179 & n3871;
  assign n3873 = ~n1535 & n3872;
  assign n3874 = ~n650 & n3873;
  assign n3875 = n53754 & n3859;
  assign n3876 = ~n53741 & ~n53774;
  assign n3877 = ~n881 & ~n2103;
  assign n3878 = ~n1491 & ~n1634;
  assign n3879 = ~n292 & ~n614;
  assign n3880 = n3878 & n3879;
  assign n3881 = n3877 & n3880;
  assign n3882 = ~n402 & ~n585;
  assign n3883 = ~n567 & ~n611;
  assign n3884 = ~n402 & ~n567;
  assign n3885 = ~n611 & n3884;
  assign n3886 = ~n585 & n3885;
  assign n3887 = n3882 & n3883;
  assign n3888 = ~n346 & ~n410;
  assign n3889 = ~n513 & ~n1469;
  assign n3890 = n3888 & n3889;
  assign n3891 = n53775 & n3890;
  assign n3892 = n3878 & n53775;
  assign n3893 = ~n881 & n3892;
  assign n3894 = ~n2103 & n3893;
  assign n3895 = ~n1469 & n3894;
  assign n3896 = ~n292 & n3895;
  assign n3897 = ~n513 & n3896;
  assign n3898 = ~n410 & n3897;
  assign n3899 = ~n614 & n3898;
  assign n3900 = ~n346 & n3899;
  assign n3901 = ~n346 & ~n513;
  assign n3902 = n3877 & n3901;
  assign n3903 = n3878 & n3902;
  assign n3904 = ~n410 & ~n1469;
  assign n3905 = n3879 & n3904;
  assign n3906 = n53775 & n3905;
  assign n3907 = n3903 & n3906;
  assign n3908 = ~n292 & ~n2103;
  assign n3909 = n3901 & n3908;
  assign n3910 = n3878 & n3909;
  assign n3911 = ~n881 & ~n1469;
  assign n3912 = ~n410 & ~n614;
  assign n3913 = n3911 & n3912;
  assign n3914 = n53775 & n3913;
  assign n3915 = n3910 & n3914;
  assign n3916 = ~n513 & ~n614;
  assign n3917 = n3911 & n3916;
  assign n3918 = n3878 & n3917;
  assign n3919 = ~n292 & ~n346;
  assign n3920 = ~n410 & ~n2103;
  assign n3921 = n3919 & n3920;
  assign n3922 = n53775 & n3921;
  assign n3923 = n3918 & n3922;
  assign n3924 = n3881 & n3891;
  assign n3925 = ~n584 & ~n659;
  assign n3926 = ~n659 & ~n1033;
  assign n3927 = ~n584 & n3926;
  assign n3928 = ~n1033 & n3925;
  assign n3929 = ~n404 & ~n823;
  assign n3930 = ~n1124 & ~n1465;
  assign n3931 = n3929 & n3930;
  assign n3932 = ~n166 & ~n565;
  assign n3933 = ~n360 & ~n774;
  assign n3934 = n3932 & n3933;
  assign n3935 = n3931 & n3934;
  assign n3936 = n53777 & n3935;
  assign n3937 = ~n219 & ~n587;
  assign n3938 = ~n1059 & n2053;
  assign n3939 = ~n219 & n2053;
  assign n3940 = ~n1059 & n3939;
  assign n3941 = ~n587 & n3940;
  assign n3942 = ~n587 & ~n1059;
  assign n3943 = ~n1059 & n3937;
  assign n3944 = ~n219 & n3942;
  assign n3945 = n2053 & n53779;
  assign n3946 = n3937 & n3938;
  assign n3947 = ~n499 & ~n832;
  assign n3948 = ~n459 & ~n1471;
  assign n3949 = n3947 & n3948;
  assign n3950 = ~n364 & ~n1680;
  assign n3951 = ~n829 & ~n957;
  assign n3952 = n3950 & n3951;
  assign n3953 = n3949 & n3952;
  assign n3954 = n53778 & n3953;
  assign n3955 = n3947 & n3951;
  assign n3956 = n3931 & n3955;
  assign n3957 = n53777 & n3956;
  assign n3958 = n3948 & n3950;
  assign n3959 = n3934 & n3958;
  assign n3960 = n53778 & n3959;
  assign n3961 = n3957 & n3960;
  assign n3962 = ~n360 & ~n957;
  assign n3963 = ~n774 & ~n823;
  assign n3964 = n3962 & n3963;
  assign n3965 = ~n829 & ~n1465;
  assign n3966 = ~n404 & ~n1124;
  assign n3967 = n3965 & n3966;
  assign n3968 = ~n957 & ~n1465;
  assign n3969 = ~n829 & ~n1124;
  assign n3970 = n3968 & n3969;
  assign n3971 = n3929 & n3933;
  assign n3972 = n3970 & n3971;
  assign n3973 = n3964 & n3967;
  assign n3974 = n53777 & n53781;
  assign n3975 = n3932 & n3947;
  assign n3976 = n3958 & n3975;
  assign n3977 = n53778 & n3976;
  assign n3978 = n3974 & n3977;
  assign n3979 = n3936 & n3954;
  assign n3980 = n53778 & n3975;
  assign n3981 = n53776 & n3980;
  assign n3982 = n53777 & n3981;
  assign n3983 = n3950 & n3982;
  assign n3984 = ~n1124 & n3983;
  assign n3985 = ~n1471 & n3984;
  assign n3986 = ~n957 & n3985;
  assign n3987 = ~n1465 & n3986;
  assign n3988 = ~n404 & n3987;
  assign n3989 = ~n823 & n3988;
  assign n3990 = ~n459 & n3989;
  assign n3991 = ~n829 & n3990;
  assign n3992 = ~n360 & n3991;
  assign n3993 = ~n774 & n3992;
  assign n3994 = n53776 & n53780;
  assign n3995 = ~n357 & ~n588;
  assign n3996 = ~n754 & ~n776;
  assign n3997 = ~n357 & ~n776;
  assign n3998 = ~n588 & ~n754;
  assign n3999 = n3997 & n3998;
  assign n4000 = n3995 & n3996;
  assign n4001 = n53626 & n53783;
  assign n4002 = ~n562 & ~n956;
  assign n4003 = n903 & n4002;
  assign n4004 = ~n408 & ~n742;
  assign n4005 = ~n408 & ~n1881;
  assign n4006 = ~n742 & n4005;
  assign n4007 = ~n742 & ~n1881;
  assign n4008 = ~n408 & n4007;
  assign n4009 = ~n1881 & n4004;
  assign n4010 = n4003 & n53784;
  assign n4011 = n4001 & n4010;
  assign n4012 = ~n493 & ~n631;
  assign n4013 = ~n112 & ~n1044;
  assign n4014 = n445 & n4013;
  assign n4015 = ~n631 & n4014;
  assign n4016 = ~n493 & n4015;
  assign n4017 = n4012 & n4013;
  assign n4018 = n445 & n4017;
  assign n4019 = n4012 & n4014;
  assign n4020 = ~n206 & ~n1031;
  assign n4021 = ~n568 & ~n748;
  assign n4022 = ~n211 & ~n361;
  assign n4023 = n4021 & n4022;
  assign n4024 = n4020 & n4023;
  assign n4025 = n217 & n712;
  assign n4026 = ~n249 & ~n1490;
  assign n4027 = n3535 & n4026;
  assign n4028 = n4025 & n4027;
  assign n4029 = n4022 & n4026;
  assign n4030 = n4020 & n4029;
  assign n4031 = n3535 & n4021;
  assign n4032 = n4025 & n4031;
  assign n4033 = n4030 & n4032;
  assign n4034 = n712 & n4023;
  assign n4035 = n217 & n4020;
  assign n4036 = n4027 & n4035;
  assign n4037 = n4034 & n4036;
  assign n4038 = n4024 & n4028;
  assign n4039 = n53785 & n53786;
  assign n4040 = n53784 & n4021;
  assign n4041 = n4020 & n4040;
  assign n4042 = n53626 & n4041;
  assign n4043 = n53785 & n4042;
  assign n4044 = n217 & n4043;
  assign n4045 = n3535 & n4044;
  assign n4046 = n4002 & n4045;
  assign n4047 = n712 & n4046;
  assign n4048 = n4026 & n4047;
  assign n4049 = n903 & n4048;
  assign n4050 = ~n211 & n4049;
  assign n4051 = ~n357 & n4050;
  assign n4052 = ~n361 & n4051;
  assign n4053 = ~n754 & n4052;
  assign n4054 = ~n776 & n4053;
  assign n4055 = ~n588 & n4054;
  assign n4056 = n4020 & n4022;
  assign n4057 = n53783 & n4056;
  assign n4058 = n53626 & n53784;
  assign n4059 = n4057 & n4058;
  assign n4060 = n217 & n3535;
  assign n4061 = n903 & n4060;
  assign n4062 = n4002 & n4026;
  assign n4063 = n712 & n4021;
  assign n4064 = n4062 & n4063;
  assign n4065 = n4061 & n4064;
  assign n4066 = n53785 & n4065;
  assign n4067 = n4059 & n4066;
  assign n4068 = n4011 & n4039;
  assign n4069 = ~n618 & n1659;
  assign n4070 = ~n179 & ~n310;
  assign n4071 = ~n340 & ~n741;
  assign n4072 = n4070 & n4071;
  assign n4073 = n1659 & n4070;
  assign n4074 = ~n618 & n4073;
  assign n4075 = ~n340 & n4074;
  assign n4076 = ~n741 & n4075;
  assign n4077 = ~n618 & n4070;
  assign n4078 = n1659 & n4071;
  assign n4079 = n4077 & n4078;
  assign n4080 = ~n618 & n4071;
  assign n4081 = n4073 & n4080;
  assign n4082 = n4069 & n4072;
  assign n4083 = ~n363 & ~n1492;
  assign n4084 = ~n466 & ~n1191;
  assign n4085 = n1716 & n4084;
  assign n4086 = n1716 & n4083;
  assign n4087 = ~n1191 & n4086;
  assign n4088 = ~n466 & n4087;
  assign n4089 = n4083 & n4084;
  assign n4090 = n1716 & n4089;
  assign n4091 = n4083 & n4085;
  assign n4092 = ~n420 & ~n650;
  assign n4093 = n3607 & n4092;
  assign n4094 = ~n414 & ~n833;
  assign n4095 = ~n405 & ~n660;
  assign n4096 = n4094 & n4095;
  assign n4097 = n4092 & n4094;
  assign n4098 = n3607 & n4095;
  assign n4099 = n4097 & n4098;
  assign n4100 = n4093 & n4096;
  assign n4101 = n53789 & n53790;
  assign n4102 = n53788 & n4101;
  assign n4103 = ~n625 & ~n773;
  assign n4104 = ~n272 & ~n461;
  assign n4105 = ~n773 & n4104;
  assign n4106 = ~n625 & n4105;
  assign n4107 = ~n272 & ~n625;
  assign n4108 = ~n461 & ~n773;
  assign n4109 = n4107 & n4108;
  assign n4110 = n4103 & n4104;
  assign n4111 = ~n222 & ~n342;
  assign n4112 = ~n450 & ~n1196;
  assign n4113 = ~n342 & ~n450;
  assign n4114 = ~n222 & ~n1196;
  assign n4115 = n4113 & n4114;
  assign n4116 = n4111 & n4112;
  assign n4117 = ~n495 & ~n564;
  assign n4118 = n270 & n4117;
  assign n4119 = n4111 & n4117;
  assign n4120 = ~n268 & ~n450;
  assign n4121 = ~n269 & ~n1196;
  assign n4122 = n4120 & n4121;
  assign n4123 = n4119 & n4122;
  assign n4124 = n53792 & n4118;
  assign n4125 = ~n1196 & n53791;
  assign n4126 = ~n222 & n4125;
  assign n4127 = ~n564 & n4126;
  assign n4128 = ~n495 & n4127;
  assign n4129 = ~n269 & n4128;
  assign n4130 = ~n268 & n4129;
  assign n4131 = ~n450 & n4130;
  assign n4132 = ~n342 & n4131;
  assign n4133 = n53791 & n53793;
  assign n4134 = ~n168 & ~n510;
  assign n4135 = ~n168 & ~n1125;
  assign n4136 = ~n510 & n4135;
  assign n4137 = ~n1125 & n4134;
  assign n4138 = n164 & n2367;
  assign n4139 = n53795 & n4138;
  assign n4140 = ~n172 & ~n615;
  assign n4141 = ~n172 & n318;
  assign n4142 = ~n615 & n4141;
  assign n4143 = n318 & n4140;
  assign n4144 = ~n896 & ~n1477;
  assign n4145 = n309 & ~n896;
  assign n4146 = ~n1477 & n4145;
  assign n4147 = n309 & n4144;
  assign n4148 = n53796 & n53797;
  assign n4149 = n4139 & n4148;
  assign n4150 = n53794 & n4149;
  assign n4151 = n164 & n4095;
  assign n4152 = n4097 & n4151;
  assign n4153 = n53788 & n4152;
  assign n4154 = n53789 & n4153;
  assign n4155 = n2367 & n3607;
  assign n4156 = n53795 & n4155;
  assign n4157 = n4148 & n4156;
  assign n4158 = n53794 & n4157;
  assign n4159 = n4154 & n4158;
  assign n4160 = n2367 & n4094;
  assign n4161 = n164 & n3607;
  assign n4162 = n4160 & n4161;
  assign n4163 = n53788 & n4162;
  assign n4164 = n53789 & n4163;
  assign n4165 = ~n405 & ~n420;
  assign n4166 = ~n660 & n4165;
  assign n4167 = ~n510 & ~n1125;
  assign n4168 = ~n168 & ~n650;
  assign n4169 = n4167 & n4168;
  assign n4170 = n4166 & n4169;
  assign n4171 = n4148 & n4170;
  assign n4172 = n53794 & n4171;
  assign n4173 = n4164 & n4172;
  assign n4174 = n4102 & n4150;
  assign n4175 = n53787 & n53798;
  assign n4176 = n3607 & n53797;
  assign n4177 = n53796 & n4176;
  assign n4178 = n53789 & n4177;
  assign n4179 = n53788 & n4178;
  assign n4180 = n53794 & n4179;
  assign n4181 = n53787 & n4180;
  assign n4182 = n4094 & n4181;
  assign n4183 = n53782 & n4182;
  assign n4184 = n2367 & n4183;
  assign n4185 = n164 & n4184;
  assign n4186 = ~n1125 & n4185;
  assign n4187 = ~n168 & n4186;
  assign n4188 = ~n660 & n4187;
  assign n4189 = ~n405 & n4188;
  assign n4190 = ~n510 & n4189;
  assign n4191 = ~n420 & n4190;
  assign n4192 = ~n650 & n4191;
  assign n4193 = n53782 & n53798;
  assign n4194 = n53787 & n4193;
  assign n4195 = n53782 & n4175;
  assign n4196 = ~n53774 & ~n53799;
  assign n4197 = ~n172 & ~n879;
  assign n4198 = n2340 & n3561;
  assign n4199 = ~n879 & n4198;
  assign n4200 = ~n172 & n4199;
  assign n4201 = n2340 & n4197;
  assign n4202 = n3561 & n4201;
  assign n4203 = n4197 & n4198;
  assign n4204 = ~n307 & ~n984;
  assign n4205 = n772 & n4204;
  assign n4206 = ~n1125 & ~n1680;
  assign n4207 = n1577 & n4206;
  assign n4208 = n772 & n4207;
  assign n4209 = ~n984 & n4208;
  assign n4210 = ~n307 & n4209;
  assign n4211 = n4205 & n4207;
  assign n4212 = ~n507 & ~n552;
  assign n4213 = ~n448 & ~n568;
  assign n4214 = ~n587 & ~n741;
  assign n4215 = n4213 & n4214;
  assign n4216 = n4212 & n4214;
  assign n4217 = n4213 & n4216;
  assign n4218 = n4212 & n4215;
  assign n4219 = n53801 & n53802;
  assign n4220 = n53800 & n53802;
  assign n4221 = n53801 & n4220;
  assign n4222 = n53800 & n4219;
  assign n4223 = ~n349 & ~n495;
  assign n4224 = ~n179 & ~n1465;
  assign n4225 = ~n464 & ~n1127;
  assign n4226 = n4224 & n4225;
  assign n4227 = n4223 & n4226;
  assign n4228 = ~n615 & n1670;
  assign n4229 = ~n614 & n4228;
  assign n4230 = n616 & n1670;
  assign n4231 = ~n405 & ~n567;
  assign n4232 = ~n774 & ~n1081;
  assign n4233 = n4231 & n4232;
  assign n4234 = n53804 & n4233;
  assign n4235 = n4224 & n53804;
  assign n4236 = n4223 & n4235;
  assign n4237 = ~n464 & n4236;
  assign n4238 = ~n1127 & n4237;
  assign n4239 = ~n1081 & n4238;
  assign n4240 = ~n567 & n4239;
  assign n4241 = ~n405 & n4240;
  assign n4242 = ~n774 & n4241;
  assign n4243 = ~n405 & ~n774;
  assign n4244 = n4224 & n4243;
  assign n4245 = n4223 & n4244;
  assign n4246 = ~n567 & ~n1081;
  assign n4247 = n4225 & n4246;
  assign n4248 = n53804 & n4247;
  assign n4249 = n4245 & n4248;
  assign n4250 = ~n464 & ~n567;
  assign n4251 = n4223 & n4250;
  assign n4252 = n4224 & n4251;
  assign n4253 = ~n405 & ~n1127;
  assign n4254 = n4232 & n4253;
  assign n4255 = n53804 & n4254;
  assign n4256 = n4252 & n4255;
  assign n4257 = n4227 & n4234;
  assign n4258 = ~n166 & ~n564;
  assign n4259 = ~n622 & ~n1085;
  assign n4260 = n4258 & n4259;
  assign n4261 = ~n294 & ~n777;
  assign n4262 = ~n268 & ~n650;
  assign n4263 = n4261 & n4262;
  assign n4264 = n4259 & n4262;
  assign n4265 = n4258 & n4261;
  assign n4266 = n4264 & n4265;
  assign n4267 = n4260 & n4263;
  assign n4268 = ~n255 & ~n275;
  assign n4269 = ~n275 & ~n356;
  assign n4270 = ~n255 & n4269;
  assign n4271 = ~n255 & ~n356;
  assign n4272 = ~n275 & n4271;
  assign n4273 = ~n356 & n4268;
  assign n4274 = ~n788 & n3014;
  assign n4275 = n53807 & n4274;
  assign n4276 = n53806 & n4275;
  assign n4277 = n53805 & n4276;
  assign n4278 = n4213 & n4258;
  assign n4279 = n4212 & n4278;
  assign n4280 = n53800 & n4279;
  assign n4281 = n53801 & n4280;
  assign n4282 = n3014 & n4261;
  assign n4283 = n4264 & n4282;
  assign n4284 = ~n788 & n4214;
  assign n4285 = n53807 & n4284;
  assign n4286 = n4283 & n4285;
  assign n4287 = n53805 & n4286;
  assign n4288 = n4281 & n4287;
  assign n4289 = n4259 & n4261;
  assign n4290 = n4212 & n4289;
  assign n4291 = n53801 & n4290;
  assign n4292 = n53800 & n4291;
  assign n4293 = n4214 & n4262;
  assign n4294 = n3014 & n4258;
  assign n4295 = n4293 & n4294;
  assign n4296 = ~n788 & n4213;
  assign n4297 = n53807 & n4296;
  assign n4298 = n4295 & n4297;
  assign n4299 = n53805 & n4298;
  assign n4300 = n4292 & n4299;
  assign n4301 = n53803 & n4277;
  assign n4302 = ~n144 & ~n1769;
  assign n4303 = ~n144 & ~n1192;
  assign n4304 = ~n1769 & n4303;
  assign n4305 = ~n1192 & n4302;
  assign n4306 = ~n212 & ~n2109;
  assign n4307 = ~n212 & ~n1061;
  assign n4308 = ~n2109 & n4307;
  assign n4309 = ~n1061 & n4306;
  assign n4310 = n3085 & n4094;
  assign n4311 = n53810 & n4310;
  assign n4312 = n53809 & n4311;
  assign n4313 = ~n215 & ~n829;
  assign n4314 = ~n141 & ~n588;
  assign n4315 = n1032 & n4314;
  assign n4316 = n4313 & n4315;
  assign n4317 = ~n416 & ~n560;
  assign n4318 = n1816 & n4317;
  assign n4319 = ~n221 & ~n733;
  assign n4320 = ~n901 & ~n1466;
  assign n4321 = n4319 & n4320;
  assign n4322 = n4318 & n4321;
  assign n4323 = n4313 & n4319;
  assign n4324 = n4320 & n4323;
  assign n4325 = n1816 & n4314;
  assign n4326 = n1032 & n4317;
  assign n4327 = n4325 & n4326;
  assign n4328 = n4324 & n4327;
  assign n4329 = n4316 & n4322;
  assign n4330 = n1816 & n4320;
  assign n4331 = n4314 & n4330;
  assign n4332 = n4320 & n4325;
  assign n4333 = n1032 & n4313;
  assign n4334 = n4310 & n4333;
  assign n4335 = n3085 & n53812;
  assign n4336 = n4094 & n4335;
  assign n4337 = n4313 & n4336;
  assign n4338 = n1032 & n4337;
  assign n4339 = n53812 & n4334;
  assign n4340 = n53809 & n53813;
  assign n4341 = n4317 & n4340;
  assign n4342 = n4319 & n4341;
  assign n4343 = ~n1061 & n4342;
  assign n4344 = ~n212 & n4343;
  assign n4345 = ~n2109 & n4344;
  assign n4346 = n3085 & n4319;
  assign n4347 = n53810 & n4346;
  assign n4348 = n53809 & n4347;
  assign n4349 = n1816 & n4313;
  assign n4350 = n1032 & n4349;
  assign n4351 = n4094 & n4314;
  assign n4352 = n4317 & n4320;
  assign n4353 = n4351 & n4352;
  assign n4354 = n4350 & n4353;
  assign n4355 = n4348 & n4354;
  assign n4356 = n4317 & n4319;
  assign n4357 = n53810 & n4356;
  assign n4358 = n53809 & n4357;
  assign n4359 = n53813 & n4358;
  assign n4360 = n4312 & n53811;
  assign n4361 = n3001 & n3272;
  assign n4362 = n1673 & n4002;
  assign n4363 = n4361 & n4362;
  assign n4364 = ~n451 & ~n513;
  assign n4365 = ~n222 & ~n513;
  assign n4366 = ~n451 & n4365;
  assign n4367 = ~n222 & n4364;
  assign n4368 = ~n740 & n2093;
  assign n4369 = n53815 & n4368;
  assign n4370 = n2093 & n3272;
  assign n4371 = n4362 & n4370;
  assign n4372 = ~n740 & n3001;
  assign n4373 = n53815 & n4372;
  assign n4374 = n4371 & n4373;
  assign n4375 = n4363 & n4369;
  assign n4376 = ~n272 & ~n753;
  assign n4377 = ~n461 & ~n1881;
  assign n4378 = ~n269 & ~n983;
  assign n4379 = n4377 & n4378;
  assign n4380 = n4376 & n4379;
  assign n4381 = ~n360 & ~n1079;
  assign n4382 = n3948 & n4381;
  assign n4383 = ~n354 & ~n1457;
  assign n4384 = n2001 & n4383;
  assign n4385 = n4382 & n4384;
  assign n4386 = n4376 & n4381;
  assign n4387 = n4383 & n4386;
  assign n4388 = n3948 & n4377;
  assign n4389 = n2001 & n4378;
  assign n4390 = n4388 & n4389;
  assign n4391 = n4387 & n4390;
  assign n4392 = n4380 & n4385;
  assign n4393 = n3272 & n53815;
  assign n4394 = n3001 & n4393;
  assign n4395 = n4383 & n4394;
  assign n4396 = n4376 & n4395;
  assign n4397 = n1673 & n4396;
  assign n4398 = n4002 & n4397;
  assign n4399 = n4378 & n4398;
  assign n4400 = n2093 & n4399;
  assign n4401 = n4381 & n4400;
  assign n4402 = ~n1471 & n4401;
  assign n4403 = ~n310 & n4402;
  assign n4404 = ~n459 & n4403;
  assign n4405 = ~n461 & n4404;
  assign n4406 = ~n647 & n4405;
  assign n4407 = ~n740 & n4406;
  assign n4408 = ~n1881 & n4407;
  assign n4409 = n4002 & n4381;
  assign n4410 = n4379 & n4409;
  assign n4411 = ~n740 & n2001;
  assign n4412 = n53815 & n4411;
  assign n4413 = n4410 & n4412;
  assign n4414 = n3948 & n4376;
  assign n4415 = n4383 & n4414;
  assign n4416 = n1673 & n3001;
  assign n4417 = n4370 & n4416;
  assign n4418 = n4415 & n4417;
  assign n4419 = n4413 & n4418;
  assign n4420 = ~n647 & ~n1471;
  assign n4421 = ~n459 & ~n1881;
  assign n4422 = n4420 & n4421;
  assign n4423 = n2093 & n4381;
  assign n4424 = n4422 & n4423;
  assign n4425 = ~n461 & ~n740;
  assign n4426 = ~n310 & n4425;
  assign n4427 = n53815 & n4426;
  assign n4428 = n4424 & n4427;
  assign n4429 = n3001 & n4383;
  assign n4430 = n3272 & n4429;
  assign n4431 = n4002 & n4378;
  assign n4432 = n1673 & n4376;
  assign n4433 = n4431 & n4432;
  assign n4434 = n4430 & n4433;
  assign n4435 = n4428 & n4434;
  assign n4436 = n53816 & n53817;
  assign n4437 = n53814 & n53818;
  assign n4438 = n53808 & n4437;
  assign n4439 = n4212 & n4262;
  assign n4440 = n53807 & n4439;
  assign n4441 = n4259 & n4440;
  assign n4442 = n53800 & n4441;
  assign n4443 = n53805 & n4442;
  assign n4444 = n53818 & n4443;
  assign n4445 = n53814 & n4444;
  assign n4446 = n53733 & n4445;
  assign n4447 = n53801 & n4446;
  assign n4448 = n4261 & n4447;
  assign n4449 = n3014 & n4448;
  assign n4450 = n4258 & n4449;
  assign n4451 = n4214 & n4450;
  assign n4452 = ~n568 & n4451;
  assign n4453 = ~n788 & n4452;
  assign n4454 = ~n448 & n4453;
  assign n4455 = n53733 & n4438;
  assign n4456 = ~n53799 & ~n53819;
  assign n4457 = ~n419 & ~n2201;
  assign n4458 = ~n625 & n1674;
  assign n4459 = ~n419 & n1674;
  assign n4460 = ~n2201 & n4459;
  assign n4461 = ~n625 & n4460;
  assign n4462 = ~n625 & ~n2201;
  assign n4463 = ~n419 & ~n625;
  assign n4464 = ~n2201 & n4463;
  assign n4465 = ~n419 & n4462;
  assign n4466 = n1674 & n53821;
  assign n4467 = n4457 & n4458;
  assign n4468 = ~n1042 & ~n1088;
  assign n4469 = ~n1033 & n4468;
  assign n4470 = ~n650 & ~n1034;
  assign n4471 = n3678 & n4470;
  assign n4472 = ~n848 & ~n1478;
  assign n4473 = n1919 & n4472;
  assign n4474 = n1919 & n3678;
  assign n4475 = n4470 & n4472;
  assign n4476 = n4474 & n4475;
  assign n4477 = n4471 & n4473;
  assign n4478 = ~n1088 & ~n1478;
  assign n4479 = ~n848 & n4478;
  assign n4480 = ~n1033 & ~n1042;
  assign n4481 = n4470 & n4480;
  assign n4482 = n4474 & n4481;
  assign n4483 = n4479 & n4482;
  assign n4484 = ~n1033 & ~n1478;
  assign n4485 = ~n1088 & n4484;
  assign n4486 = ~n848 & ~n1469;
  assign n4487 = ~n255 & ~n1042;
  assign n4488 = n4486 & n4487;
  assign n4489 = n4471 & n4488;
  assign n4490 = n4485 & n4489;
  assign n4491 = n4469 & n53822;
  assign n4492 = n53820 & n4471;
  assign n4493 = ~n1088 & n4492;
  assign n4494 = ~n1033 & n4493;
  assign n4495 = ~n1469 & n4494;
  assign n4496 = ~n1478 & n4495;
  assign n4497 = ~n255 & n4496;
  assign n4498 = ~n1042 & n4497;
  assign n4499 = ~n848 & n4498;
  assign n4500 = n53820 & n53823;
  assign n4501 = ~n144 & ~n832;
  assign n4502 = ~n316 & n4501;
  assign n4503 = ~n590 & n3742;
  assign n4504 = ~n611 & ~n948;
  assign n4505 = n358 & ~n948;
  assign n4506 = ~n611 & n4505;
  assign n4507 = n358 & n4504;
  assign n4508 = n4503 & n53825;
  assign n4509 = n4502 & n4508;
  assign n4510 = ~n956 & n1659;
  assign n4511 = ~n1658 & n2814;
  assign n4512 = ~n272 & ~n733;
  assign n4513 = n2913 & n4512;
  assign n4514 = ~n1191 & n1659;
  assign n4515 = ~n272 & n4514;
  assign n4516 = ~n956 & n4515;
  assign n4517 = ~n733 & n4516;
  assign n4518 = ~n344 & n4517;
  assign n4519 = ~n344 & ~n956;
  assign n4520 = ~n1191 & n4519;
  assign n4521 = n1659 & n4512;
  assign n4522 = n4520 & n4521;
  assign n4523 = n53826 & n4513;
  assign n4524 = ~n554 & ~n740;
  assign n4525 = ~n1466 & n4524;
  assign n4526 = ~n317 & ~n614;
  assign n4527 = n2476 & n4526;
  assign n4528 = n4525 & n4527;
  assign n4529 = ~n651 & ~n2042;
  assign n4530 = ~n207 & ~n1641;
  assign n4531 = n4529 & n4530;
  assign n4532 = n53767 & n4531;
  assign n4533 = n4528 & n4532;
  assign n4534 = n53827 & n4533;
  assign n4535 = n53767 & n53825;
  assign n4536 = n53825 & n4532;
  assign n4537 = n4531 & n4535;
  assign n4538 = ~n590 & ~n740;
  assign n4539 = n318 & n2476;
  assign n4540 = n4538 & n4539;
  assign n4541 = ~n614 & ~n1466;
  assign n4542 = ~n554 & ~n614;
  assign n4543 = ~n1466 & n4542;
  assign n4544 = ~n554 & ~n1466;
  assign n4545 = ~n614 & n4544;
  assign n4546 = ~n554 & n4541;
  assign n4547 = n3742 & n4501;
  assign n4548 = n53829 & n4547;
  assign n4549 = n4538 & n4547;
  assign n4550 = n4539 & n53829;
  assign n4551 = n4549 & n4550;
  assign n4552 = n4540 & n4548;
  assign n4553 = n53827 & n53830;
  assign n4554 = n53828 & n4553;
  assign n4555 = n53767 & n53829;
  assign n4556 = n53825 & n4555;
  assign n4557 = n4501 & n4538;
  assign n4558 = n4529 & n4557;
  assign n4559 = n2476 & n3742;
  assign n4560 = n318 & n4530;
  assign n4561 = n4559 & n4560;
  assign n4562 = n4558 & n4561;
  assign n4563 = n53827 & n4562;
  assign n4564 = n4556 & n4563;
  assign n4565 = n4509 & n4534;
  assign n4566 = n53825 & n4529;
  assign n4567 = n4501 & n4566;
  assign n4568 = n53767 & n4567;
  assign n4569 = n53827 & n4568;
  assign n4570 = n4538 & n4569;
  assign n4571 = n53824 & n4570;
  assign n4572 = n2476 & n4571;
  assign n4573 = n4530 & n4572;
  assign n4574 = n318 & n4573;
  assign n4575 = n3742 & n4574;
  assign n4576 = ~n1466 & n4575;
  assign n4577 = ~n554 & n4576;
  assign n4578 = ~n614 & n4577;
  assign n4579 = n53824 & n53831;
  assign n4580 = ~n441 & ~n750;
  assign n4581 = ~n441 & n802;
  assign n4582 = ~n750 & n4581;
  assign n4583 = n802 & n4580;
  assign n4584 = ~n422 & ~n1680;
  assign n4585 = ~n141 & ~n1468;
  assign n4586 = n4584 & n4585;
  assign n4587 = ~n168 & ~n448;
  assign n4588 = n1186 & n4587;
  assign n4589 = n4586 & n4588;
  assign n4590 = ~n250 & ~n291;
  assign n4591 = n648 & n4590;
  assign n4592 = n4070 & n4258;
  assign n4593 = n4591 & n4592;
  assign n4594 = n4589 & n4593;
  assign n4595 = n53833 & n4594;
  assign n4596 = ~n101 & ~n182;
  assign n4597 = ~n101 & ~n459;
  assign n4598 = ~n182 & n4597;
  assign n4599 = ~n459 & n4596;
  assign n4600 = n2577 & n53834;
  assign n4601 = n53546 & n2577;
  assign n4602 = ~n101 & n4601;
  assign n4603 = ~n182 & n4602;
  assign n4604 = ~n459 & n4603;
  assign n4605 = n53546 & n4600;
  assign n4606 = ~n216 & ~n222;
  assign n4607 = ~n216 & ~n1477;
  assign n4608 = ~n222 & n4607;
  assign n4609 = ~n222 & ~n1477;
  assign n4610 = ~n216 & n4609;
  assign n4611 = ~n1477 & n4606;
  assign n4612 = ~n742 & ~n1337;
  assign n4613 = ~n1646 & n4612;
  assign n4614 = n53489 & n4613;
  assign n4615 = n53836 & n4614;
  assign n4616 = n53835 & n4615;
  assign n4617 = n53489 & n53833;
  assign n4618 = n1186 & n4617;
  assign n4619 = n53836 & n4618;
  assign n4620 = n648 & n4619;
  assign n4621 = n53835 & n4620;
  assign n4622 = n4585 & n4621;
  assign n4623 = n4584 & n4622;
  assign n4624 = n4070 & n4623;
  assign n4625 = n4587 & n4624;
  assign n4626 = n4258 & n4625;
  assign n4627 = ~n291 & n4626;
  assign n4628 = ~n250 & n4627;
  assign n4629 = ~n1337 & n4628;
  assign n4630 = ~n742 & n4629;
  assign n4631 = ~n1646 & n4630;
  assign n4632 = n4258 & n4584;
  assign n4633 = n1186 & n4585;
  assign n4634 = n4632 & n4633;
  assign n4635 = ~n250 & ~n1337;
  assign n4636 = n4587 & n4635;
  assign n4637 = n648 & n4070;
  assign n4638 = n4636 & n4637;
  assign n4639 = n4634 & n4638;
  assign n4640 = n53833 & n4639;
  assign n4641 = ~n291 & ~n742;
  assign n4642 = ~n1646 & n4641;
  assign n4643 = n53836 & n4642;
  assign n4644 = n53489 & n4643;
  assign n4645 = n53835 & n4644;
  assign n4646 = n4640 & n4645;
  assign n4647 = n4070 & n4587;
  assign n4648 = n648 & n4584;
  assign n4649 = n4647 & n4648;
  assign n4650 = ~n291 & ~n1646;
  assign n4651 = n1186 & n4650;
  assign n4652 = n4258 & n4585;
  assign n4653 = n4651 & n4652;
  assign n4654 = n4649 & n4653;
  assign n4655 = n53833 & n4654;
  assign n4656 = ~n250 & ~n742;
  assign n4657 = ~n1337 & n4656;
  assign n4658 = n53836 & n4657;
  assign n4659 = n53489 & n4658;
  assign n4660 = n53835 & n4659;
  assign n4661 = n4655 & n4660;
  assign n4662 = n4595 & n4616;
  assign n4663 = ~n663 & n1642;
  assign n4664 = n53592 & n53605;
  assign n4665 = n4663 & n4664;
  assign n4666 = ~n108 & n3672;
  assign n4667 = ~n443 & n4666;
  assign n4668 = ~n503 & ~n776;
  assign n4669 = ~n1681 & n4668;
  assign n4670 = ~n401 & ~n588;
  assign n4671 = n3562 & n4670;
  assign n4672 = n4669 & n4671;
  assign n4673 = n4667 & n4672;
  assign n4674 = ~n401 & ~n1681;
  assign n4675 = ~n503 & ~n588;
  assign n4676 = ~n588 & ~n1681;
  assign n4677 = ~n401 & ~n503;
  assign n4678 = n4676 & n4677;
  assign n4679 = n4674 & n4675;
  assign n4680 = n53592 & n53838;
  assign n4681 = n53605 & n53838;
  assign n4682 = n53592 & n4681;
  assign n4683 = n53605 & n4680;
  assign n4684 = n1642 & n3082;
  assign n4685 = n3562 & n4684;
  assign n4686 = n4667 & n4685;
  assign n4687 = n53839 & n4686;
  assign n4688 = n3562 & n4676;
  assign n4689 = n53605 & n4688;
  assign n4690 = n53592 & n4689;
  assign n4691 = n1642 & n4677;
  assign n4692 = n3082 & n4691;
  assign n4693 = n4667 & n4692;
  assign n4694 = n4690 & n4693;
  assign n4695 = n4665 & n4673;
  assign n4696 = n1368 & n2690;
  assign n4697 = ~n753 & ~n1065;
  assign n4698 = n2002 & n4697;
  assign n4699 = n4696 & n4698;
  assign n4700 = ~n218 & ~n249;
  assign n4701 = ~n218 & ~n507;
  assign n4702 = ~n249 & n4701;
  assign n4703 = ~n249 & ~n507;
  assign n4704 = ~n218 & n4703;
  assign n4705 = ~n507 & n4700;
  assign n4706 = ~n259 & ~n553;
  assign n4707 = ~n321 & ~n774;
  assign n4708 = n4706 & n4707;
  assign n4709 = n53841 & n4708;
  assign n4710 = ~n567 & ~n896;
  assign n4711 = n2690 & n53841;
  assign n4712 = n4710 & n4711;
  assign n4713 = ~n1065 & n4712;
  assign n4714 = ~n883 & n4713;
  assign n4715 = ~n308 & n4714;
  assign n4716 = ~n321 & n4715;
  assign n4717 = ~n259 & n4716;
  assign n4718 = ~n553 & n4717;
  assign n4719 = ~n774 & n4718;
  assign n4720 = ~n753 & n4719;
  assign n4721 = ~n259 & ~n321;
  assign n4722 = n2690 & n4721;
  assign n4723 = n4698 & n4722;
  assign n4724 = ~n553 & ~n774;
  assign n4725 = n1368 & n4724;
  assign n4726 = n53841 & n4725;
  assign n4727 = n4723 & n4726;
  assign n4728 = ~n259 & ~n774;
  assign n4729 = n4710 & n4728;
  assign n4730 = n2690 & n4697;
  assign n4731 = n4729 & n4730;
  assign n4732 = ~n321 & ~n883;
  assign n4733 = ~n308 & ~n553;
  assign n4734 = n4732 & n4733;
  assign n4735 = n53841 & n4734;
  assign n4736 = n4731 & n4735;
  assign n4737 = ~n259 & ~n753;
  assign n4738 = ~n553 & ~n1065;
  assign n4739 = n4737 & n4738;
  assign n4740 = n2690 & n4710;
  assign n4741 = n4739 & n4740;
  assign n4742 = ~n308 & ~n883;
  assign n4743 = n4707 & n4742;
  assign n4744 = n53841 & n4743;
  assign n4745 = n4741 & n4744;
  assign n4746 = n4699 & n4709;
  assign n4747 = ~n246 & ~n414;
  assign n4748 = ~n414 & ~n1280;
  assign n4749 = ~n246 & n4748;
  assign n4750 = ~n1280 & n4747;
  assign n4751 = ~n662 & ~n1189;
  assign n4752 = ~n1476 & ~n1769;
  assign n4753 = ~n499 & ~n1234;
  assign n4754 = n4752 & n4753;
  assign n4755 = n4751 & n4754;
  assign n4756 = n4751 & n4753;
  assign n4757 = ~n414 & n4756;
  assign n4758 = ~n1476 & n4757;
  assign n4759 = ~n246 & n4758;
  assign n4760 = ~n1280 & n4759;
  assign n4761 = ~n1769 & n4760;
  assign n4762 = ~n246 & n4752;
  assign n4763 = n4748 & n4753;
  assign n4764 = n4751 & n4763;
  assign n4765 = n4762 & n4764;
  assign n4766 = n53843 & n4755;
  assign n4767 = n53842 & n53844;
  assign n4768 = n53840 & n4767;
  assign n4769 = n53837 & n4768;
  assign n4770 = n53592 & n4667;
  assign n4771 = n53605 & n4770;
  assign n4772 = n53837 & n4771;
  assign n4773 = n53844 & n4772;
  assign n4774 = n3082 & n4773;
  assign n4775 = n53832 & n4774;
  assign n4776 = n53842 & n4775;
  assign n4777 = n1642 & n4776;
  assign n4778 = ~n1681 & n4777;
  assign n4779 = ~n401 & n4778;
  assign n4780 = ~n833 & n4779;
  assign n4781 = ~n503 & n4780;
  assign n4782 = ~n491 & n4781;
  assign n4783 = ~n588 & n4782;
  assign n4784 = n53832 & n4769;
  assign n4785 = ~n53819 & ~n53845;
  assign n4786 = ~n216 & ~n464;
  assign n4787 = ~n216 & ~n1641;
  assign n4788 = ~n464 & n4787;
  assign n4789 = ~n1641 & n4786;
  assign n4790 = n846 & n3165;
  assign n4791 = ~n161 & ~n1912;
  assign n4792 = n4538 & n4791;
  assign n4793 = n4790 & n4792;
  assign n4794 = n53846 & n4793;
  assign n4795 = ~n272 & ~n1469;
  assign n4796 = ~n177 & ~n585;
  assign n4797 = n4795 & n4796;
  assign n4798 = ~n879 & ~n1088;
  assign n4799 = ~n364 & ~n1658;
  assign n4800 = ~n1088 & n4799;
  assign n4801 = ~n879 & n4800;
  assign n4802 = n4798 & n4799;
  assign n4803 = ~n1469 & n53847;
  assign n4804 = ~n177 & n4803;
  assign n4805 = ~n272 & n4804;
  assign n4806 = ~n585 & n4805;
  assign n4807 = ~n585 & ~n879;
  assign n4808 = ~n177 & ~n1088;
  assign n4809 = n4796 & n4798;
  assign n4810 = ~n177 & ~n879;
  assign n4811 = ~n585 & ~n1088;
  assign n4812 = n4810 & n4811;
  assign n4813 = n4807 & n4808;
  assign n4814 = n4795 & n4799;
  assign n4815 = n53849 & n4814;
  assign n4816 = n4797 & n53847;
  assign n4817 = ~n295 & ~n342;
  assign n4818 = ~n754 & ~n914;
  assign n4819 = ~n977 & n4818;
  assign n4820 = ~n914 & ~n977;
  assign n4821 = ~n295 & ~n977;
  assign n4822 = ~n914 & n4821;
  assign n4823 = ~n295 & n4820;
  assign n4824 = ~n342 & n53850;
  assign n4825 = ~n754 & n4824;
  assign n4826 = ~n342 & ~n754;
  assign n4827 = n53850 & n4826;
  assign n4828 = ~n342 & ~n914;
  assign n4829 = ~n754 & n4828;
  assign n4830 = n4821 & n4829;
  assign n4831 = n4817 & n4819;
  assign n4832 = ~n317 & ~n460;
  assign n4833 = ~n770 & ~n984;
  assign n4834 = n1060 & n4833;
  assign n4835 = n4832 & n4834;
  assign n4836 = n53851 & n4835;
  assign n4837 = n53848 & n4836;
  assign n4838 = n1060 & n4790;
  assign n4839 = n53848 & n4838;
  assign n4840 = n1060 & n3165;
  assign n4841 = n53851 & n4840;
  assign n4842 = n846 & n4841;
  assign n4843 = n53848 & n4842;
  assign n4844 = n53851 & n4839;
  assign n4845 = n4833 & n53852;
  assign n4846 = n4538 & n4845;
  assign n4847 = ~n464 & n4846;
  assign n4848 = ~n317 & n4847;
  assign n4849 = ~n161 & n4848;
  assign n4850 = ~n216 & n4849;
  assign n4851 = ~n1641 & n4850;
  assign n4852 = ~n460 & n4851;
  assign n4853 = ~n1912 & n4852;
  assign n4854 = n4538 & n4832;
  assign n4855 = n4790 & n4854;
  assign n4856 = n53846 & n4855;
  assign n4857 = n4791 & n4834;
  assign n4858 = n53848 & n4857;
  assign n4859 = n53851 & n4858;
  assign n4860 = n4856 & n4859;
  assign n4861 = n3165 & n4538;
  assign n4862 = n4791 & n4832;
  assign n4863 = n4861 & n4862;
  assign n4864 = n53846 & n4863;
  assign n4865 = n846 & n1060;
  assign n4866 = n4833 & n4865;
  assign n4867 = n53851 & n4866;
  assign n4868 = n53848 & n4867;
  assign n4869 = n4864 & n4868;
  assign n4870 = ~n216 & n4832;
  assign n4871 = ~n464 & ~n1641;
  assign n4872 = n4791 & n4871;
  assign n4873 = n4538 & n4833;
  assign n4874 = n4872 & n4873;
  assign n4875 = n4870 & n4874;
  assign n4876 = n53852 & n4875;
  assign n4877 = n4794 & n4837;
  assign n4878 = ~n308 & ~n503;
  assign n4879 = ~n777 & ~n1125;
  assign n4880 = ~n503 & ~n1125;
  assign n4881 = ~n308 & ~n777;
  assign n4882 = n4880 & n4881;
  assign n4883 = n4878 & n4879;
  assign n4884 = ~n211 & ~n822;
  assign n4885 = n2256 & n4884;
  assign n4886 = ~n1125 & n4885;
  assign n4887 = ~n308 & n4886;
  assign n4888 = ~n503 & n4887;
  assign n4889 = ~n777 & n4888;
  assign n4890 = n53854 & n4885;
  assign n4891 = n2058 & n4223;
  assign n4892 = ~n849 & ~n1090;
  assign n4893 = ~n105 & ~n1127;
  assign n4894 = n4892 & n4893;
  assign n4895 = n4891 & n4894;
  assign n4896 = ~n101 & ~n591;
  assign n4897 = ~n101 & ~n405;
  assign n4898 = ~n591 & n4897;
  assign n4899 = ~n405 & n4896;
  assign n4900 = n421 & n3675;
  assign n4901 = n53856 & n4900;
  assign n4902 = n2058 & n3675;
  assign n4903 = n4223 & n4892;
  assign n4904 = n4902 & n4903;
  assign n4905 = n421 & n4893;
  assign n4906 = n53856 & n4905;
  assign n4907 = n4904 & n4906;
  assign n4908 = n4895 & n4901;
  assign n4909 = n53855 & n53857;
  assign n4910 = ~n611 & ~n630;
  assign n4911 = ~n316 & ~n630;
  assign n4912 = ~n611 & n4911;
  assign n4913 = ~n316 & n4910;
  assign n4914 = ~n824 & ~n1466;
  assign n4915 = n2367 & n4914;
  assign n4916 = ~n416 & n4212;
  assign n4917 = n4915 & n4916;
  assign n4918 = n53858 & n4917;
  assign n4919 = n53745 & n4918;
  assign n4920 = n3675 & n4892;
  assign n4921 = n4893 & n4914;
  assign n4922 = n4920 & n4921;
  assign n4923 = n421 & n4223;
  assign n4924 = n2058 & n2367;
  assign n4925 = n4923 & n4924;
  assign n4926 = n4922 & n4925;
  assign n4927 = n53855 & n4926;
  assign n4928 = n53856 & n4916;
  assign n4929 = n53858 & n4928;
  assign n4930 = n53745 & n4929;
  assign n4931 = n4927 & n4930;
  assign n4932 = n4909 & n4919;
  assign n4933 = n53576 & n53859;
  assign n4934 = n53858 & n4914;
  assign n4935 = n4893 & n4934;
  assign n4936 = n4892 & n4935;
  assign n4937 = n53853 & n4936;
  assign n4938 = n53576 & n4937;
  assign n4939 = n4916 & n4938;
  assign n4940 = n4223 & n4939;
  assign n4941 = n3675 & n4940;
  assign n4942 = n53745 & n4941;
  assign n4943 = n53855 & n4942;
  assign n4944 = n2058 & n4943;
  assign n4945 = n421 & n4944;
  assign n4946 = n2367 & n4945;
  assign n4947 = ~n101 & n4946;
  assign n4948 = ~n405 & n4947;
  assign n4949 = ~n591 & n4948;
  assign n4950 = n53853 & n4933;
  assign n4951 = ~n53845 & ~n53860;
  assign n4952 = ~n255 & ~n631;
  assign n4953 = ~n255 & ~n1455;
  assign n4954 = ~n631 & n4953;
  assign n4955 = ~n1455 & n4952;
  assign n4956 = ~n631 & n4206;
  assign n4957 = ~n255 & n4956;
  assign n4958 = ~n1455 & n4957;
  assign n4959 = n4206 & n53861;
  assign n4960 = ~n451 & ~n649;
  assign n4961 = ~n649 & n4663;
  assign n4962 = ~n451 & n4961;
  assign n4963 = ~n451 & ~n663;
  assign n4964 = ~n649 & n4963;
  assign n4965 = ~n663 & n4960;
  assign n4966 = n1642 & n53864;
  assign n4967 = n4663 & n4960;
  assign n4968 = n53524 & n53863;
  assign n4969 = n53524 & n53862;
  assign n4970 = n53863 & n4969;
  assign n4971 = n53862 & n4968;
  assign n4972 = ~n319 & ~n503;
  assign n4973 = n652 & n4972;
  assign n4974 = ~n177 & ~n630;
  assign n4975 = ~n622 & ~n741;
  assign n4976 = n4974 & n4975;
  assign n4977 = n652 & n4975;
  assign n4978 = n4972 & n4974;
  assign n4979 = n4977 & n4978;
  assign n4980 = ~n319 & ~n622;
  assign n4981 = ~n503 & ~n741;
  assign n4982 = n4980 & n4981;
  assign n4983 = n652 & n4974;
  assign n4984 = n4982 & n4983;
  assign n4985 = n4973 & n4976;
  assign n4986 = ~n342 & ~n514;
  assign n4987 = ~n342 & ~n735;
  assign n4988 = ~n514 & n4987;
  assign n4989 = ~n514 & ~n735;
  assign n4990 = ~n342 & n4989;
  assign n4991 = ~n735 & n4986;
  assign n4992 = ~n141 & ~n222;
  assign n4993 = ~n414 & ~n1191;
  assign n4994 = ~n141 & ~n414;
  assign n4995 = ~n222 & ~n1191;
  assign n4996 = n4994 & n4995;
  assign n4997 = n4992 & n4993;
  assign n4998 = n53867 & n53868;
  assign n4999 = n4974 & n53867;
  assign n5000 = n652 & n4999;
  assign n5001 = ~n414 & n5000;
  assign n5002 = ~n1191 & n5001;
  assign n5003 = ~n222 & n5002;
  assign n5004 = ~n141 & n5003;
  assign n5005 = ~n319 & n5004;
  assign n5006 = ~n503 & n5005;
  assign n5007 = ~n741 & n5006;
  assign n5008 = ~n622 & n5007;
  assign n5009 = ~n414 & ~n503;
  assign n5010 = n4974 & n5009;
  assign n5011 = n4977 & n5010;
  assign n5012 = ~n222 & ~n319;
  assign n5013 = ~n141 & ~n1191;
  assign n5014 = n5012 & n5013;
  assign n5015 = n53867 & n5014;
  assign n5016 = n5011 & n5015;
  assign n5017 = n53866 & n4998;
  assign n5018 = ~n565 & ~n823;
  assign n5019 = ~n830 & ~n2201;
  assign n5020 = n5018 & n5019;
  assign n5021 = ~n108 & ~n824;
  assign n5022 = n4319 & n5021;
  assign n5023 = n5020 & n5022;
  assign n5024 = ~n163 & n749;
  assign n5025 = n53762 & n5024;
  assign n5026 = n749 & n5021;
  assign n5027 = n4319 & n5018;
  assign n5028 = n5026 & n5027;
  assign n5029 = ~n163 & ~n830;
  assign n5030 = ~n2201 & n5029;
  assign n5031 = n53762 & n5030;
  assign n5032 = n5028 & n5031;
  assign n5033 = n4319 & n5019;
  assign n5034 = n5026 & n5033;
  assign n5035 = ~n163 & ~n823;
  assign n5036 = ~n565 & n5035;
  assign n5037 = n53762 & n5036;
  assign n5038 = n5034 & n5037;
  assign n5039 = n5023 & n5025;
  assign n5040 = n53869 & n53870;
  assign n5041 = n53516 & n53870;
  assign n5042 = n53869 & n5041;
  assign n5043 = n53516 & n5040;
  assign n5044 = n53762 & n53863;
  assign n5045 = n53524 & n5044;
  assign n5046 = n53869 & n5045;
  assign n5047 = n5021 & n5046;
  assign n5048 = n53516 & n5047;
  assign n5049 = n749 & n5048;
  assign n5050 = n53862 & n5049;
  assign n5051 = n4319 & n5050;
  assign n5052 = ~n163 & n5051;
  assign n5053 = ~n565 & n5052;
  assign n5054 = ~n823 & n5053;
  assign n5055 = ~n830 & n5054;
  assign n5056 = ~n2201 & n5055;
  assign n5057 = n53865 & n53871;
  assign n5058 = ~n219 & ~n311;
  assign n5059 = ~n356 & ~n560;
  assign n5060 = ~n983 & ~n1492;
  assign n5061 = n5059 & n5060;
  assign n5062 = n5058 & n5059;
  assign n5063 = n5060 & n5062;
  assign n5064 = n5058 & n5061;
  assign n5065 = ~n291 & ~n410;
  assign n5066 = ~n291 & ~n1703;
  assign n5067 = ~n410 & n5066;
  assign n5068 = ~n1703 & n5065;
  assign n5069 = ~n423 & ~n1491;
  assign n5070 = ~n754 & ~n1491;
  assign n5071 = ~n423 & n5070;
  assign n5072 = ~n754 & n5069;
  assign n5073 = ~n833 & ~n1912;
  assign n5074 = n3062 & n5073;
  assign n5075 = n53875 & n5074;
  assign n5076 = n53874 & n5075;
  assign n5077 = n53874 & n53875;
  assign n5078 = n5058 & n5077;
  assign n5079 = n5060 & n5078;
  assign n5080 = n3062 & n5079;
  assign n5081 = ~n560 & n5080;
  assign n5082 = ~n833 & n5081;
  assign n5083 = ~n356 & n5082;
  assign n5084 = ~n1912 & n5083;
  assign n5085 = n3062 & n5060;
  assign n5086 = n5058 & n5085;
  assign n5087 = n5059 & n5073;
  assign n5088 = n53875 & n5087;
  assign n5089 = n53874 & n5088;
  assign n5090 = n5086 & n5089;
  assign n5091 = n53873 & n5076;
  assign n5092 = ~n1457 & ~n1641;
  assign n5093 = ~n507 & ~n1280;
  assign n5094 = ~n1280 & ~n1457;
  assign n5095 = ~n1641 & n5094;
  assign n5096 = ~n507 & n5095;
  assign n5097 = ~n1280 & ~n1641;
  assign n5098 = ~n507 & ~n1457;
  assign n5099 = n5097 & n5098;
  assign n5100 = n5092 & n5093;
  assign n5101 = ~n422 & ~n447;
  assign n5102 = ~n1478 & ~n2103;
  assign n5103 = n5101 & n5102;
  assign n5104 = n53784 & n5103;
  assign n5105 = n53877 & n5104;
  assign n5106 = ~n307 & ~n584;
  assign n5107 = n355 & n1671;
  assign n5108 = ~n307 & n5107;
  assign n5109 = ~n584 & n5108;
  assign n5110 = n1671 & n5106;
  assign n5111 = n355 & n5110;
  assign n5112 = n5106 & n5107;
  assign n5113 = ~n405 & ~n1468;
  assign n5114 = n4501 & n5113;
  assign n5115 = ~n1466 & ~n1487;
  assign n5116 = ~n101 & ~n662;
  assign n5117 = n5115 & n5116;
  assign n5118 = n5114 & n5117;
  assign n5119 = n53878 & n5118;
  assign n5120 = n5102 & n5115;
  assign n5121 = n53784 & n5120;
  assign n5122 = n53877 & n5121;
  assign n5123 = n5113 & n5116;
  assign n5124 = n4501 & n5101;
  assign n5125 = n5123 & n5124;
  assign n5126 = n53878 & n5125;
  assign n5127 = n5122 & n5126;
  assign n5128 = ~n447 & ~n2103;
  assign n5129 = ~n1478 & ~n1487;
  assign n5130 = n5128 & n5129;
  assign n5131 = n53877 & n5130;
  assign n5132 = n53784 & n5131;
  assign n5133 = ~n422 & ~n1466;
  assign n5134 = n4501 & n5133;
  assign n5135 = n5123 & n5134;
  assign n5136 = n53878 & n5135;
  assign n5137 = n5132 & n5136;
  assign n5138 = n5105 & n5119;
  assign n5139 = n53784 & n4501;
  assign n5140 = n53878 & n5139;
  assign n5141 = n53876 & n5140;
  assign n5142 = n53877 & n5141;
  assign n5143 = n5116 & n5142;
  assign n5144 = n5113 & n5143;
  assign n5145 = ~n422 & n5144;
  assign n5146 = ~n2103 & n5145;
  assign n5147 = ~n1466 & n5146;
  assign n5148 = ~n1487 & n5147;
  assign n5149 = ~n1478 & n5148;
  assign n5150 = ~n447 & n5149;
  assign n5151 = n53876 & n53879;
  assign n5152 = ~n1634 & ~n2042;
  assign n5153 = n347 & n5152;
  assign n5154 = ~n1195 & ~n1997;
  assign n5155 = n3802 & n5154;
  assign n5156 = ~n321 & ~n404;
  assign n5157 = ~n611 & ~n776;
  assign n5158 = n5156 & n5157;
  assign n5159 = n3802 & n5156;
  assign n5160 = n5154 & n5157;
  assign n5161 = n5159 & n5160;
  assign n5162 = n5155 & n5158;
  assign n5163 = ~n465 & ~n1634;
  assign n5164 = ~n611 & ~n1189;
  assign n5165 = n5163 & n5164;
  assign n5166 = ~n776 & ~n2042;
  assign n5167 = n5154 & n5166;
  assign n5168 = n347 & n5156;
  assign n5169 = n5167 & n5168;
  assign n5170 = n5165 & n5169;
  assign n5171 = ~n776 & ~n1195;
  assign n5172 = ~n321 & ~n1189;
  assign n5173 = n5171 & n5172;
  assign n5174 = ~n611 & ~n1997;
  assign n5175 = ~n404 & ~n465;
  assign n5176 = n5174 & n5175;
  assign n5177 = n5153 & n5176;
  assign n5178 = n5173 & n5177;
  assign n5179 = n5153 & n53881;
  assign n5180 = ~n212 & ~n1486;
  assign n5181 = ~n902 & n1939;
  assign n5182 = ~n212 & ~n894;
  assign n5183 = ~n894 & ~n1486;
  assign n5184 = ~n212 & n5183;
  assign n5185 = ~n1486 & n5182;
  assign n5186 = ~n902 & n53883;
  assign n5187 = ~n879 & n5186;
  assign n5188 = ~n879 & ~n902;
  assign n5189 = n53883 & n5188;
  assign n5190 = n5180 & n5181;
  assign n5191 = ~n1476 & n4261;
  assign n5192 = n4261 & n4833;
  assign n5193 = ~n1476 & n5192;
  assign n5194 = n4833 & n5191;
  assign n5195 = n53884 & n53885;
  assign n5196 = n53882 & n5195;
  assign n5197 = n1712 & n3716;
  assign n5198 = ~n409 & ~n1646;
  assign n5199 = ~n295 & ~n357;
  assign n5200 = n5198 & n5199;
  assign n5201 = n5197 & n5200;
  assign n5202 = ~n308 & ~n360;
  assign n5203 = ~n499 & ~n788;
  assign n5204 = n5202 & n5203;
  assign n5205 = ~n259 & ~n590;
  assign n5206 = n3273 & n5205;
  assign n5207 = ~n259 & ~n308;
  assign n5208 = ~n590 & ~n788;
  assign n5209 = n5207 & n5208;
  assign n5210 = ~n360 & ~n499;
  assign n5211 = n3273 & n5210;
  assign n5212 = n5209 & n5211;
  assign n5213 = n5204 & n5206;
  assign n5214 = n3716 & n5198;
  assign n5215 = n3273 & n5214;
  assign n5216 = n5199 & n5215;
  assign n5217 = n1712 & n5216;
  assign n5218 = ~n308 & n5217;
  assign n5219 = ~n259 & n5218;
  assign n5220 = ~n360 & n5219;
  assign n5221 = n5203 & n5220;
  assign n5222 = ~n590 & n5221;
  assign n5223 = n1712 & n5199;
  assign n5224 = n5198 & n5203;
  assign n5225 = n5223 & n5224;
  assign n5226 = n5202 & n5205;
  assign n5227 = n3273 & n3716;
  assign n5228 = n5226 & n5227;
  assign n5229 = n5225 & n5228;
  assign n5230 = n1712 & n5203;
  assign n5231 = n5214 & n5230;
  assign n5232 = n3273 & n5199;
  assign n5233 = n5226 & n5232;
  assign n5234 = n5231 & n5233;
  assign n5235 = n5201 & n53886;
  assign n5236 = n53528 & n53887;
  assign n5237 = n5196 & n5236;
  assign n5238 = n53880 & n5237;
  assign n5239 = n53880 & n5195;
  assign n5240 = n53887 & n5239;
  assign n5241 = n53528 & n5240;
  assign n5242 = n347 & n5241;
  assign n5243 = n53872 & n5242;
  assign n5244 = ~n1997 & n5243;
  assign n5245 = ~n1195 & n5244;
  assign n5246 = ~n321 & n5245;
  assign n5247 = ~n404 & n5246;
  assign n5248 = ~n1189 & n5247;
  assign n5249 = ~n1634 & n5248;
  assign n5250 = ~n611 & n5249;
  assign n5251 = ~n465 & n5250;
  assign n5252 = ~n776 & n5251;
  assign n5253 = ~n2042 & n5252;
  assign n5254 = n53872 & n5238;
  assign n5255 = ~n53860 & ~n53888;
  assign n5256 = n4587 & n4710;
  assign n5257 = n1851 & n2038;
  assign n5258 = n1851 & n4587;
  assign n5259 = n2038 & n4710;
  assign n5260 = n5258 & n5259;
  assign n5261 = n5256 & n5257;
  assign n5262 = ~n416 & n772;
  assign n5263 = n3925 & n4103;
  assign n5264 = n5262 & n5263;
  assign n5265 = n772 & n3925;
  assign n5266 = n5257 & n5265;
  assign n5267 = ~n416 & n4587;
  assign n5268 = n4103 & n4710;
  assign n5269 = n5267 & n5268;
  assign n5270 = n5266 & n5269;
  assign n5271 = n53889 & n5264;
  assign n5272 = n53884 & n53890;
  assign n5273 = ~n491 & ~n1062;
  assign n5274 = ~n1062 & n53862;
  assign n5275 = ~n491 & n5274;
  assign n5276 = n53862 & n5273;
  assign n5277 = ~n776 & ~n1042;
  assign n5278 = n1458 & n5277;
  assign n5279 = n802 & n4666;
  assign n5280 = n5278 & n5279;
  assign n5281 = n53659 & n5280;
  assign n5282 = n53891 & n5281;
  assign n5283 = n2038 & n53891;
  assign n5284 = n53884 & n5283;
  assign n5285 = n802 & n5284;
  assign n5286 = n772 & n5285;
  assign n5287 = n5277 & n5286;
  assign n5288 = n4710 & n5287;
  assign n5289 = n53659 & n5288;
  assign n5290 = n4587 & n5289;
  assign n5291 = n1458 & n5290;
  assign n5292 = ~n416 & n5291;
  assign n5293 = n4666 & n5292;
  assign n5294 = ~n659 & n5293;
  assign n5295 = ~n247 & n5294;
  assign n5296 = ~n584 & n5295;
  assign n5297 = ~n495 & n5296;
  assign n5298 = ~n773 & n5297;
  assign n5299 = ~n625 & n5298;
  assign n5300 = n1458 & n2038;
  assign n5301 = n5256 & n5300;
  assign n5302 = ~n416 & ~n659;
  assign n5303 = n4103 & n5302;
  assign n5304 = n772 & n5277;
  assign n5305 = n5303 & n5304;
  assign n5306 = n5301 & n5305;
  assign n5307 = n53884 & n5306;
  assign n5308 = ~n495 & ~n584;
  assign n5309 = ~n247 & n5308;
  assign n5310 = n802 & n5309;
  assign n5311 = n4666 & n5310;
  assign n5312 = n53659 & n5311;
  assign n5313 = n53891 & n5312;
  assign n5314 = n5307 & n5313;
  assign n5315 = n5272 & n5282;
  assign n5316 = ~n747 & ~n1081;
  assign n5317 = ~n901 & ~n1476;
  assign n5318 = ~n1081 & ~n1476;
  assign n5319 = ~n747 & ~n901;
  assign n5320 = n5318 & n5319;
  assign n5321 = n5316 & n5317;
  assign n5322 = ~n112 & ~n824;
  assign n5323 = ~n161 & ~n553;
  assign n5324 = n5322 & n5323;
  assign n5325 = ~n824 & ~n901;
  assign n5326 = ~n112 & ~n1081;
  assign n5327 = n5325 & n5326;
  assign n5328 = ~n747 & ~n1476;
  assign n5329 = n5323 & n5328;
  assign n5330 = n5327 & n5329;
  assign n5331 = n53893 & n5324;
  assign n5332 = ~n1033 & ~n1715;
  assign n5333 = ~n440 & ~n591;
  assign n5334 = ~n591 & ~n1033;
  assign n5335 = ~n440 & n5334;
  assign n5336 = ~n1715 & n5335;
  assign n5337 = ~n591 & ~n1715;
  assign n5338 = ~n440 & ~n1033;
  assign n5339 = n5337 & n5338;
  assign n5340 = n5332 & n5333;
  assign n5341 = ~n346 & ~n1465;
  assign n5342 = ~n414 & ~n1465;
  assign n5343 = ~n346 & n5342;
  assign n5344 = ~n414 & n5341;
  assign n5345 = n53725 & n53896;
  assign n5346 = n53725 & n53895;
  assign n5347 = n53896 & n5346;
  assign n5348 = n53895 & n5345;
  assign n5349 = ~n901 & n53897;
  assign n5350 = ~n1476 & n5349;
  assign n5351 = ~n1081 & n5350;
  assign n5352 = ~n112 & n5351;
  assign n5353 = ~n161 & n5352;
  assign n5354 = ~n553 & n5353;
  assign n5355 = ~n824 & n5354;
  assign n5356 = ~n747 & n5355;
  assign n5357 = n53894 & n53897;
  assign n5358 = ~n623 & ~n822;
  assign n5359 = ~n774 & ~n1490;
  assign n5360 = n5358 & n5359;
  assign n5361 = ~n182 & ~n1124;
  assign n5362 = ~n464 & ~n565;
  assign n5363 = n5361 & n5362;
  assign n5364 = ~n1490 & n5363;
  assign n5365 = ~n822 & n5364;
  assign n5366 = ~n774 & n5365;
  assign n5367 = ~n623 & n5366;
  assign n5368 = n5360 & n5363;
  assign n5369 = ~n172 & ~n423;
  assign n5370 = ~n172 & ~n977;
  assign n5371 = ~n423 & n5370;
  assign n5372 = ~n977 & n5369;
  assign n5373 = ~n977 & n1035;
  assign n5374 = ~n172 & n5373;
  assign n5375 = ~n423 & n5374;
  assign n5376 = n1035 & n53900;
  assign n5377 = ~n833 & ~n1061;
  assign n5378 = ~n647 & ~n1031;
  assign n5379 = n3523 & n5378;
  assign n5380 = n5377 & n5378;
  assign n5381 = n3523 & n5380;
  assign n5382 = n5377 & n5379;
  assign n5383 = n53901 & n53902;
  assign n5384 = n53899 & n53902;
  assign n5385 = n53901 & n5384;
  assign n5386 = n53899 & n5383;
  assign n5387 = ~n444 & n1659;
  assign n5388 = ~n496 & ~n1634;
  assign n5389 = n53809 & n5388;
  assign n5390 = ~n444 & ~n496;
  assign n5391 = n53809 & n5390;
  assign n5392 = n1659 & n5391;
  assign n5393 = ~n1634 & n5392;
  assign n5394 = ~n1634 & n1659;
  assign n5395 = n5390 & n5394;
  assign n5396 = n53809 & n5395;
  assign n5397 = n5387 & n5389;
  assign n5398 = ~n735 & ~n1280;
  assign n5399 = ~n957 & ~n1044;
  assign n5400 = n5398 & n5399;
  assign n5401 = ~n256 & ~n552;
  assign n5402 = n2975 & n5401;
  assign n5403 = ~n735 & ~n957;
  assign n5404 = ~n552 & ~n1044;
  assign n5405 = n5403 & n5404;
  assign n5406 = ~n256 & ~n1280;
  assign n5407 = n2975 & n5406;
  assign n5408 = n5405 & n5407;
  assign n5409 = n5400 & n5402;
  assign n5410 = n53673 & n4531;
  assign n5411 = ~n552 & ~n1280;
  assign n5412 = n2975 & n5411;
  assign n5413 = n4531 & n5412;
  assign n5414 = ~n256 & ~n735;
  assign n5415 = n5399 & n5414;
  assign n5416 = n53673 & n5415;
  assign n5417 = n5413 & n5416;
  assign n5418 = n53905 & n5410;
  assign n5419 = n53904 & n53906;
  assign n5420 = n53903 & n5419;
  assign n5421 = n53898 & n5420;
  assign n5422 = n3523 & n4529;
  assign n5423 = n53901 & n5422;
  assign n5424 = n53904 & n5423;
  assign n5425 = n53898 & n5424;
  assign n5426 = n53892 & n5425;
  assign n5427 = n53899 & n5426;
  assign n5428 = n5378 & n5427;
  assign n5429 = n2975 & n5428;
  assign n5430 = n53673 & n5429;
  assign n5431 = n4530 & n5430;
  assign n5432 = n5377 & n5431;
  assign n5433 = ~n1044 & n5432;
  assign n5434 = ~n957 & n5433;
  assign n5435 = ~n256 & n5434;
  assign n5436 = ~n552 & n5435;
  assign n5437 = ~n1280 & n5436;
  assign n5438 = ~n735 & n5437;
  assign n5439 = n53892 & n5421;
  assign n5440 = ~n53888 & ~n53907;
  assign n5441 = ~n163 & ~n356;
  assign n5442 = ~n163 & ~n956;
  assign n5443 = ~n356 & n5442;
  assign n5444 = ~n956 & n5441;
  assign n5445 = ~n105 & n1391;
  assign n5446 = ~n294 & ~n514;
  assign n5447 = ~n493 & ~n1535;
  assign n5448 = ~n294 & ~n1535;
  assign n5449 = ~n493 & ~n514;
  assign n5450 = n5448 & n5449;
  assign n5451 = n5446 & n5447;
  assign n5452 = ~n514 & n5447;
  assign n5453 = ~n105 & ~n294;
  assign n5454 = n1391 & n5453;
  assign n5455 = n5452 & n5454;
  assign n5456 = n5445 & n53909;
  assign n5457 = n1391 & n53908;
  assign n5458 = ~n105 & n5457;
  assign n5459 = ~n294 & n5458;
  assign n5460 = ~n493 & n5459;
  assign n5461 = ~n1535 & n5460;
  assign n5462 = ~n514 & n5461;
  assign n5463 = n53908 & n53910;
  assign n5464 = ~n849 & ~n1085;
  assign n5465 = ~n1044 & n5464;
  assign n5466 = ~n308 & ~n615;
  assign n5467 = ~n748 & ~n770;
  assign n5468 = n5466 & n5467;
  assign n5469 = ~n308 & ~n849;
  assign n5470 = ~n1044 & n5469;
  assign n5471 = ~n770 & ~n1085;
  assign n5472 = ~n615 & ~n748;
  assign n5473 = n5471 & n5472;
  assign n5474 = n5470 & n5473;
  assign n5475 = n5465 & n5468;
  assign n5476 = ~n584 & ~n902;
  assign n5477 = ~n219 & ~n902;
  assign n5478 = ~n584 & n5477;
  assign n5479 = ~n219 & ~n584;
  assign n5480 = ~n902 & n5479;
  assign n5481 = ~n219 & n5476;
  assign n5482 = ~n311 & n4376;
  assign n5483 = n53913 & n5482;
  assign n5484 = n53912 & n5483;
  assign n5485 = ~n444 & ~n591;
  assign n5486 = n1032 & n4584;
  assign n5487 = n5485 & n5486;
  assign n5488 = n406 & n2326;
  assign n5489 = n3947 & n4319;
  assign n5490 = n5488 & n5489;
  assign n5491 = n4319 & n4584;
  assign n5492 = n5485 & n5491;
  assign n5493 = n1032 & n3947;
  assign n5494 = n5488 & n5493;
  assign n5495 = n5492 & n5494;
  assign n5496 = n4584 & n5485;
  assign n5497 = n2326 & n5496;
  assign n5498 = n406 & n4319;
  assign n5499 = n5493 & n5498;
  assign n5500 = n5497 & n5499;
  assign n5501 = n5487 & n5490;
  assign n5502 = ~n748 & ~n1044;
  assign n5503 = ~n308 & ~n770;
  assign n5504 = n5502 & n5503;
  assign n5505 = ~n615 & ~n849;
  assign n5506 = n2326 & n5505;
  assign n5507 = n5504 & n5506;
  assign n5508 = n53913 & n5507;
  assign n5509 = n406 & n4584;
  assign n5510 = n3947 & n5485;
  assign n5511 = n5509 & n5510;
  assign n5512 = n1032 & n4319;
  assign n5513 = n3742 & n4376;
  assign n5514 = n5512 & n5513;
  assign n5515 = n5511 & n5514;
  assign n5516 = n5508 & n5515;
  assign n5517 = n5484 & n53914;
  assign n5518 = n3947 & n53913;
  assign n5519 = n5485 & n5518;
  assign n5520 = n53911 & n5519;
  assign n5521 = n4584 & n5520;
  assign n5522 = n4376 & n5521;
  assign n5523 = n1032 & n5522;
  assign n5524 = n2326 & n5523;
  assign n5525 = n406 & n5524;
  assign n5526 = n4319 & n5525;
  assign n5527 = n3742 & n5526;
  assign n5528 = ~n1044 & n5527;
  assign n5529 = ~n308 & n5528;
  assign n5530 = ~n849 & n5529;
  assign n5531 = ~n748 & n5530;
  assign n5532 = ~n615 & n5531;
  assign n5533 = ~n770 & n5532;
  assign n5534 = n53911 & n53915;
  assign n5535 = ~n353 & ~n423;
  assign n5536 = ~n496 & ~n1088;
  assign n5537 = n5535 & n5536;
  assign n5538 = ~n256 & ~n410;
  assign n5539 = ~n440 & ~n450;
  assign n5540 = ~n271 & ~n628;
  assign n5541 = n5539 & n5540;
  assign n5542 = n5538 & n5541;
  assign n5543 = ~n1088 & n5538;
  assign n5544 = ~n628 & n5543;
  assign n5545 = ~n271 & n5544;
  assign n5546 = ~n496 & n5545;
  assign n5547 = ~n440 & n5546;
  assign n5548 = ~n423 & n5547;
  assign n5549 = ~n450 & n5548;
  assign n5550 = ~n353 & n5549;
  assign n5551 = ~n423 & ~n1088;
  assign n5552 = n5540 & n5551;
  assign n5553 = ~n353 & ~n496;
  assign n5554 = n5539 & n5553;
  assign n5555 = n5538 & n5554;
  assign n5556 = n5552 & n5555;
  assign n5557 = n5535 & n5540;
  assign n5558 = ~n450 & ~n496;
  assign n5559 = ~n440 & ~n1088;
  assign n5560 = n5558 & n5559;
  assign n5561 = n5538 & n5560;
  assign n5562 = n5557 & n5561;
  assign n5563 = ~n440 & ~n628;
  assign n5564 = n5536 & n5563;
  assign n5565 = ~n423 & ~n450;
  assign n5566 = ~n271 & ~n353;
  assign n5567 = n5565 & n5566;
  assign n5568 = n5538 & n5567;
  assign n5569 = n5564 & n5568;
  assign n5570 = n5537 & n5542;
  assign n5571 = ~n554 & ~n747;
  assign n5572 = ~n984 & ~n1469;
  assign n5573 = n5571 & n5572;
  assign n5574 = n403 & n4083;
  assign n5575 = n5573 & n5574;
  assign n5576 = n1675 & n53841;
  assign n5577 = n5575 & n5576;
  assign n5578 = ~n1061 & ~n1090;
  assign n5579 = ~n588 & ~n663;
  assign n5580 = ~n144 & ~n663;
  assign n5581 = ~n588 & n5580;
  assign n5582 = ~n144 & n5579;
  assign n5583 = ~n144 & n5578;
  assign n5584 = ~n663 & n5583;
  assign n5585 = ~n588 & n5584;
  assign n5586 = n5578 & n53918;
  assign n5587 = ~n1634 & ~n1641;
  assign n5588 = ~n320 & ~n461;
  assign n5589 = n4094 & n5588;
  assign n5590 = n5587 & n5589;
  assign n5591 = n53919 & n5590;
  assign n5592 = ~n1469 & ~n1641;
  assign n5593 = ~n747 & ~n984;
  assign n5594 = n5592 & n5593;
  assign n5595 = ~n554 & ~n1634;
  assign n5596 = n403 & n5595;
  assign n5597 = n5594 & n5596;
  assign n5598 = n5576 & n5597;
  assign n5599 = n4083 & n4094;
  assign n5600 = n5588 & n5599;
  assign n5601 = n53919 & n5600;
  assign n5602 = n5598 & n5601;
  assign n5603 = ~n984 & ~n1634;
  assign n5604 = n5571 & n5603;
  assign n5605 = n4094 & n5592;
  assign n5606 = n5604 & n5605;
  assign n5607 = n5576 & n5606;
  assign n5608 = n5574 & n5588;
  assign n5609 = n53919 & n5608;
  assign n5610 = n5607 & n5609;
  assign n5611 = n5577 & n5591;
  assign n5612 = n53841 & n5588;
  assign n5613 = n53919 & n5612;
  assign n5614 = n53917 & n5613;
  assign n5615 = n1675 & n5614;
  assign n5616 = n4094 & n5615;
  assign n5617 = n4083 & n5616;
  assign n5618 = n403 & n5617;
  assign n5619 = ~n984 & n5618;
  assign n5620 = ~n1469 & n5619;
  assign n5621 = ~n554 & n5620;
  assign n5622 = ~n1634 & n5621;
  assign n5623 = ~n1641 & n5622;
  assign n5624 = ~n747 & n5623;
  assign n5625 = n53917 & n53920;
  assign n5626 = ~n247 & ~n564;
  assign n5627 = ~n172 & ~n829;
  assign n5628 = ~n172 & ~n247;
  assign n5629 = ~n564 & ~n829;
  assign n5630 = n5628 & n5629;
  assign n5631 = n5626 & n5627;
  assign n5632 = n2004 & n3000;
  assign n5633 = ~n172 & n5632;
  assign n5634 = ~n247 & n5633;
  assign n5635 = ~n564 & n5634;
  assign n5636 = ~n829 & n5635;
  assign n5637 = n53922 & n5632;
  assign n5638 = ~n1681 & n3672;
  assign n5639 = ~n451 & ~n2103;
  assign n5640 = n3638 & n5639;
  assign n5641 = n3672 & n5639;
  assign n5642 = ~n894 & n5641;
  assign n5643 = ~n1681 & n5642;
  assign n5644 = ~n1196 & n5643;
  assign n5645 = ~n1681 & n5639;
  assign n5646 = n3638 & n3672;
  assign n5647 = n5645 & n5646;
  assign n5648 = ~n1681 & n3638;
  assign n5649 = n5641 & n5648;
  assign n5650 = n5638 & n5640;
  assign n5651 = ~n506 & ~n1042;
  assign n5652 = ~n503 & ~n2201;
  assign n5653 = n1458 & n5652;
  assign n5654 = n5651 & n5653;
  assign n5655 = n53924 & n5654;
  assign n5656 = n53923 & n5655;
  assign n5657 = ~n182 & ~n466;
  assign n5658 = ~n776 & ~n1644;
  assign n5659 = n5657 & n5658;
  assign n5660 = ~n321 & ~n830;
  assign n5661 = ~n773 & ~n1471;
  assign n5662 = n799 & n5661;
  assign n5663 = n5660 & n5662;
  assign n5664 = n799 & ~n1471;
  assign n5665 = ~n321 & n5664;
  assign n5666 = ~n182 & n5665;
  assign n5667 = ~n830 & n5666;
  assign n5668 = ~n1644 & n5667;
  assign n5669 = ~n466 & n5668;
  assign n5670 = ~n776 & n5669;
  assign n5671 = ~n773 & n5670;
  assign n5672 = ~n182 & ~n830;
  assign n5673 = n5658 & n5672;
  assign n5674 = ~n321 & ~n466;
  assign n5675 = n799 & n5674;
  assign n5676 = n5661 & n5675;
  assign n5677 = n5673 & n5676;
  assign n5678 = ~n321 & ~n1644;
  assign n5679 = n5657 & n5678;
  assign n5680 = ~n776 & ~n830;
  assign n5681 = n799 & n5680;
  assign n5682 = n5661 & n5681;
  assign n5683 = n5679 & n5682;
  assign n5684 = n5674 & n5680;
  assign n5685 = ~n182 & ~n1644;
  assign n5686 = n5661 & n5685;
  assign n5687 = n799 & n5686;
  assign n5688 = n5684 & n5687;
  assign n5689 = n5659 & n5663;
  assign n5690 = ~n511 & n1541;
  assign n5691 = ~n168 & ~n1490;
  assign n5692 = n1712 & n5691;
  assign n5693 = n3011 & n5692;
  assign n5694 = n5690 & n5693;
  assign n5695 = n53925 & n5694;
  assign n5696 = n1712 & n5652;
  assign n5697 = n1458 & n1712;
  assign n5698 = n5652 & n5697;
  assign n5699 = n1458 & n5696;
  assign n5700 = n53923 & n53926;
  assign n5701 = n53924 & n53926;
  assign n5702 = n53923 & n5701;
  assign n5703 = n53924 & n5700;
  assign n5704 = ~n168 & ~n506;
  assign n5705 = ~n1042 & ~n1490;
  assign n5706 = ~n168 & ~n1042;
  assign n5707 = ~n506 & ~n1490;
  assign n5708 = n5706 & n5707;
  assign n5709 = n5704 & n5705;
  assign n5710 = n3011 & n53928;
  assign n5711 = n5690 & n5710;
  assign n5712 = n53925 & n5711;
  assign n5713 = n53927 & n5712;
  assign n5714 = n5656 & n5695;
  assign n5715 = n53921 & n53929;
  assign n5716 = n3011 & n5690;
  assign n5717 = n53924 & n5716;
  assign n5718 = n53921 & n5717;
  assign n5719 = n53916 & n5718;
  assign n5720 = n5652 & n5719;
  assign n5721 = n1712 & n5720;
  assign n5722 = n53925 & n5721;
  assign n5723 = n53923 & n5722;
  assign n5724 = n1458 & n5723;
  assign n5725 = ~n1490 & n5724;
  assign n5726 = ~n168 & n5725;
  assign n5727 = ~n1042 & n5726;
  assign n5728 = ~n506 & n5727;
  assign n5729 = n53916 & n53929;
  assign n5730 = n53921 & n5729;
  assign n5731 = n53916 & n5715;
  assign n5732 = ~n53907 & ~n53930;
  assign n5733 = ~n832 & ~n1485;
  assign n5734 = ~n553 & ~n631;
  assign n5735 = ~n174 & ~n271;
  assign n5736 = ~n271 & ~n631;
  assign n5737 = ~n174 & ~n553;
  assign n5738 = n5736 & n5737;
  assign n5739 = ~n174 & ~n631;
  assign n5740 = ~n271 & ~n553;
  assign n5741 = n5739 & n5740;
  assign n5742 = n5734 & n5735;
  assign n5743 = n5733 & n53931;
  assign n5744 = ~n346 & ~n498;
  assign n5745 = n343 & ~n498;
  assign n5746 = ~n346 & n5745;
  assign n5747 = n343 & n5744;
  assign n5748 = ~n296 & ~n1196;
  assign n5749 = ~n465 & n5748;
  assign n5750 = ~n771 & ~n1125;
  assign n5751 = ~n883 & ~n894;
  assign n5752 = ~n894 & ~n1125;
  assign n5753 = ~n771 & ~n883;
  assign n5754 = n5752 & n5753;
  assign n5755 = n5750 & n5751;
  assign n5756 = n5749 & n53933;
  assign n5757 = n53932 & n5756;
  assign n5758 = n53932 & n5749;
  assign n5759 = n5733 & n5758;
  assign n5760 = ~n1125 & n5759;
  assign n5761 = ~n883 & n5760;
  assign n5762 = ~n631 & n5761;
  assign n5763 = ~n894 & n5762;
  assign n5764 = ~n174 & n5763;
  assign n5765 = ~n271 & n5764;
  assign n5766 = ~n553 & n5765;
  assign n5767 = ~n771 & n5766;
  assign n5768 = n5733 & n53933;
  assign n5769 = n53931 & n5749;
  assign n5770 = n53932 & n5769;
  assign n5771 = n5768 & n5770;
  assign n5772 = ~n174 & ~n894;
  assign n5773 = ~n271 & ~n1125;
  assign n5774 = n5772 & n5773;
  assign n5775 = n5733 & n5774;
  assign n5776 = ~n553 & ~n883;
  assign n5777 = ~n631 & ~n771;
  assign n5778 = n5776 & n5777;
  assign n5779 = n53932 & n5778;
  assign n5780 = n5749 & n5779;
  assign n5781 = n5775 & n5780;
  assign n5782 = n5743 & n5757;
  assign n5783 = ~n215 & ~n461;
  assign n5784 = ~n461 & ~n911;
  assign n5785 = ~n215 & n5784;
  assign n5786 = ~n215 & ~n911;
  assign n5787 = ~n461 & n5786;
  assign n5788 = ~n911 & n5783;
  assign n5789 = ~n419 & ~n1455;
  assign n5790 = ~n218 & ~n349;
  assign n5791 = ~n349 & ~n504;
  assign n5792 = ~n218 & n5791;
  assign n5793 = ~n504 & n5790;
  assign n5794 = ~n218 & ~n504;
  assign n5795 = ~n349 & ~n1455;
  assign n5796 = ~n419 & n5795;
  assign n5797 = n5794 & n5796;
  assign n5798 = n5789 & n53936;
  assign n5799 = ~n218 & n53935;
  assign n5800 = ~n1455 & n5799;
  assign n5801 = ~n504 & n5800;
  assign n5802 = ~n419 & n5801;
  assign n5803 = ~n349 & n5802;
  assign n5804 = n53935 & n53937;
  assign n5805 = ~n662 & ~n1912;
  assign n5806 = n452 & n5805;
  assign n5807 = n846 & n1035;
  assign n5808 = n5806 & n5807;
  assign n5809 = ~n222 & ~n587;
  assign n5810 = ~n587 & ~n753;
  assign n5811 = ~n222 & n5810;
  assign n5812 = ~n753 & n5809;
  assign n5813 = n53517 & n53939;
  assign n5814 = n5808 & n5813;
  assign n5815 = ~n585 & ~n617;
  assign n5816 = n1091 & n2326;
  assign n5817 = ~n617 & n5816;
  assign n5818 = ~n585 & n5817;
  assign n5819 = n1091 & n5815;
  assign n5820 = n2326 & n5819;
  assign n5821 = n2326 & n5815;
  assign n5822 = n1091 & n5821;
  assign n5823 = n5815 & n5816;
  assign n5824 = n1082 & n2917;
  assign n5825 = n5277 & n5824;
  assign n5826 = n53940 & n5825;
  assign n5827 = n1035 & n5805;
  assign n5828 = n452 & n2917;
  assign n5829 = n5827 & n5828;
  assign n5830 = n5813 & n5829;
  assign n5831 = n846 & n1082;
  assign n5832 = n5277 & n5831;
  assign n5833 = n53940 & n5832;
  assign n5834 = n5830 & n5833;
  assign n5835 = ~n206 & ~n662;
  assign n5836 = ~n902 & ~n1912;
  assign n5837 = n5835 & n5836;
  assign n5838 = n846 & n5277;
  assign n5839 = n5837 & n5838;
  assign n5840 = n5813 & n5839;
  assign n5841 = n1035 & n1082;
  assign n5842 = n452 & n5841;
  assign n5843 = n53940 & n5842;
  assign n5844 = n5840 & n5843;
  assign n5845 = n5814 & n5826;
  assign n5846 = n53938 & n53941;
  assign n5847 = n53934 & n5846;
  assign n5848 = ~n353 & n1672;
  assign n5849 = ~n307 & ~n754;
  assign n5850 = ~n663 & ~n1471;
  assign n5851 = ~n307 & ~n1471;
  assign n5852 = ~n663 & n5851;
  assign n5853 = ~n754 & n5852;
  assign n5854 = ~n754 & ~n1471;
  assign n5855 = ~n307 & ~n663;
  assign n5856 = n5854 & n5855;
  assign n5857 = ~n663 & ~n754;
  assign n5858 = n5851 & n5857;
  assign n5859 = n5849 & n5850;
  assign n5860 = n5848 & n53942;
  assign n5861 = ~n310 & ~n511;
  assign n5862 = ~n310 & n2693;
  assign n5863 = ~n511 & n5862;
  assign n5864 = n2693 & n5861;
  assign n5865 = ~n168 & ~n2103;
  assign n5866 = ~n1195 & ~n2103;
  assign n5867 = ~n168 & n5866;
  assign n5868 = ~n168 & ~n1195;
  assign n5869 = ~n2103 & n5868;
  assign n5870 = ~n1195 & n5865;
  assign n5871 = n53943 & n53944;
  assign n5872 = n5860 & n5871;
  assign n5873 = ~n348 & ~n773;
  assign n5874 = ~n625 & ~n948;
  assign n5875 = n4833 & n5874;
  assign n5876 = n4833 & n5873;
  assign n5877 = n5874 & n5876;
  assign n5878 = n5873 & n5875;
  assign n5879 = ~n321 & ~n503;
  assign n5880 = ~n851 & ~n1469;
  assign n5881 = ~n321 & ~n1469;
  assign n5882 = ~n851 & n5881;
  assign n5883 = ~n503 & n5882;
  assign n5884 = n5879 & n5880;
  assign n5885 = ~n255 & ~n292;
  assign n5886 = n2981 & n5885;
  assign n5887 = n53946 & n5886;
  assign n5888 = n2981 & n5873;
  assign n5889 = n4833 & n5888;
  assign n5890 = n2981 & n5876;
  assign n5891 = n5874 & n5885;
  assign n5892 = n53946 & n5891;
  assign n5893 = n53947 & n5892;
  assign n5894 = n53945 & n5887;
  assign n5895 = n53942 & n53946;
  assign n5896 = n5848 & n53943;
  assign n5897 = n53946 & n5896;
  assign n5898 = n53942 & n5897;
  assign n5899 = n5895 & n5896;
  assign n5900 = n53944 & n5891;
  assign n5901 = n53947 & n5900;
  assign n5902 = n53949 & n5901;
  assign n5903 = n5872 & n53948;
  assign n5904 = n2981 & n53949;
  assign n5905 = n53904 & n5904;
  assign n5906 = n53944 & n5905;
  assign n5907 = n5874 & n5906;
  assign n5908 = n4833 & n5907;
  assign n5909 = n5873 & n5908;
  assign n5910 = ~n292 & n5909;
  assign n5911 = ~n255 & n5910;
  assign n5912 = n53904 & n53950;
  assign n5913 = ~n317 & ~n628;
  assign n5914 = ~n614 & n5913;
  assign n5915 = ~n614 & ~n628;
  assign n5916 = ~n317 & n5915;
  assign n5917 = ~n628 & n4526;
  assign n5918 = ~n256 & ~n623;
  assign n5919 = ~n896 & ~n1234;
  assign n5920 = ~n623 & ~n896;
  assign n5921 = ~n256 & ~n1234;
  assign n5922 = n5920 & n5921;
  assign n5923 = n5918 & n5919;
  assign n5924 = ~n896 & n53952;
  assign n5925 = ~n256 & n5924;
  assign n5926 = ~n1234 & n5925;
  assign n5927 = ~n623 & n5926;
  assign n5928 = n53952 & n53953;
  assign n5929 = ~n274 & ~n344;
  assign n5930 = ~n1476 & n5929;
  assign n5931 = ~n1457 & ~n1476;
  assign n5932 = ~n274 & n5931;
  assign n5933 = ~n1641 & n5932;
  assign n5934 = ~n344 & n5933;
  assign n5935 = ~n344 & ~n1476;
  assign n5936 = ~n274 & n5092;
  assign n5937 = n5935 & n5936;
  assign n5938 = ~n274 & ~n1641;
  assign n5939 = ~n1457 & n5935;
  assign n5940 = n5938 & n5939;
  assign n5941 = n5092 & n5930;
  assign n5942 = ~n184 & ~n441;
  assign n5943 = ~n308 & ~n554;
  assign n5944 = n472 & n5943;
  assign n5945 = n5942 & n5943;
  assign n5946 = n472 & n5945;
  assign n5947 = n5942 & n5944;
  assign n5948 = n53955 & n53956;
  assign n5949 = n53954 & n5948;
  assign n5950 = ~n514 & ~n1124;
  assign n5951 = ~n1491 & n5950;
  assign n5952 = ~n258 & ~n881;
  assign n5953 = ~n166 & ~n219;
  assign n5954 = n5952 & n5953;
  assign n5955 = ~n363 & ~n422;
  assign n5956 = ~n649 & ~n830;
  assign n5957 = n5955 & n5956;
  assign n5958 = n5954 & n5957;
  assign n5959 = ~n1124 & ~n1491;
  assign n5960 = n5955 & n5959;
  assign n5961 = n5952 & n5956;
  assign n5962 = n5955 & n5961;
  assign n5963 = ~n1124 & n5962;
  assign n5964 = ~n1491 & n5963;
  assign n5965 = n5960 & n5961;
  assign n5966 = ~n219 & n53957;
  assign n5967 = ~n166 & n5966;
  assign n5968 = ~n514 & n5967;
  assign n5969 = ~n166 & ~n1124;
  assign n5970 = ~n1491 & n5969;
  assign n5971 = ~n219 & ~n514;
  assign n5972 = n5952 & n5971;
  assign n5973 = n5957 & n5972;
  assign n5974 = n5970 & n5973;
  assign n5975 = ~n514 & ~n1491;
  assign n5976 = ~n166 & n5975;
  assign n5977 = ~n219 & ~n1124;
  assign n5978 = n5952 & n5977;
  assign n5979 = n5957 & n5978;
  assign n5980 = n5976 & n5979;
  assign n5981 = ~n166 & n5971;
  assign n5982 = n53957 & n5981;
  assign n5983 = n5951 & n5958;
  assign n5984 = n2476 & n3672;
  assign n5985 = ~n356 & ~n591;
  assign n5986 = ~n740 & ~n1477;
  assign n5987 = n5985 & n5986;
  assign n5988 = ~n627 & ~n650;
  assign n5989 = n4320 & n5988;
  assign n5990 = ~n591 & ~n650;
  assign n5991 = n5986 & n5990;
  assign n5992 = ~n356 & ~n627;
  assign n5993 = n4320 & n5992;
  assign n5994 = n5991 & n5993;
  assign n5995 = n5987 & n5989;
  assign n5996 = ~n356 & ~n740;
  assign n5997 = ~n591 & ~n627;
  assign n5998 = n5996 & n5997;
  assign n5999 = ~n650 & ~n1477;
  assign n6000 = n2476 & n5999;
  assign n6001 = n3672 & n4320;
  assign n6002 = n6000 & n6001;
  assign n6003 = n5998 & n6002;
  assign n6004 = n5984 & n53959;
  assign n6005 = n53958 & n53960;
  assign n6006 = n472 & n4320;
  assign n6007 = n53955 & n6006;
  assign n6008 = n53958 & n6007;
  assign n6009 = n53954 & n6008;
  assign n6010 = n5943 & n6009;
  assign n6011 = n2476 & n6010;
  assign n6012 = n3672 & n6011;
  assign n6013 = ~n1477 & n6012;
  assign n6014 = ~n184 & n6013;
  assign n6015 = ~n441 & n6014;
  assign n6016 = ~n591 & n6015;
  assign n6017 = ~n356 & n6016;
  assign n6018 = ~n627 & n6017;
  assign n6019 = ~n650 & n6018;
  assign n6020 = ~n740 & n6019;
  assign n6021 = n3672 & n5943;
  assign n6022 = n472 & n6021;
  assign n6023 = n53954 & n6022;
  assign n6024 = n53955 & n6023;
  assign n6025 = ~n356 & ~n441;
  assign n6026 = ~n184 & ~n740;
  assign n6027 = n6025 & n6026;
  assign n6028 = ~n627 & ~n1477;
  assign n6029 = n5990 & n6028;
  assign n6030 = n2476 & n4320;
  assign n6031 = n6029 & n6030;
  assign n6032 = n6027 & n6031;
  assign n6033 = n53958 & n6032;
  assign n6034 = n6024 & n6033;
  assign n6035 = n5949 & n6005;
  assign n6036 = n53951 & n53961;
  assign n6037 = n1082 & n5813;
  assign n6038 = n53940 & n6037;
  assign n6039 = n452 & n6038;
  assign n6040 = n53951 & n6039;
  assign n6041 = n53938 & n6040;
  assign n6042 = n53934 & n6041;
  assign n6043 = n846 & n6042;
  assign n6044 = n53961 & n6043;
  assign n6045 = n5277 & n6044;
  assign n6046 = n1035 & n6045;
  assign n6047 = ~n902 & n6046;
  assign n6048 = ~n662 & n6047;
  assign n6049 = ~n206 & n6048;
  assign n6050 = ~n1912 & n6049;
  assign n6051 = n5847 & n6036;
  assign n6052 = ~n53930 & ~n53962;
  assign n6053 = ~n354 & ~n420;
  assign n6054 = ~n852 & n6053;
  assign n6055 = n53908 & n6054;
  assign n6056 = ~n513 & ~n618;
  assign n6057 = ~n618 & ~n1234;
  assign n6058 = ~n513 & n6057;
  assign n6059 = ~n747 & n6058;
  assign n6060 = ~n513 & ~n1234;
  assign n6061 = ~n618 & ~n747;
  assign n6062 = n6060 & n6061;
  assign n6063 = n1529 & n6056;
  assign n6064 = ~n177 & ~n1641;
  assign n6065 = ~n177 & ~n2109;
  assign n6066 = ~n1641 & n6065;
  assign n6067 = ~n1641 & ~n2109;
  assign n6068 = ~n177 & n6067;
  assign n6069 = ~n2109 & n6064;
  assign n6070 = n53963 & n53964;
  assign n6071 = n6055 & n6070;
  assign n6072 = ~n591 & ~n1466;
  assign n6073 = n4117 & n6072;
  assign n6074 = ~n320 & ~n1466;
  assign n6075 = ~n256 & n6074;
  assign n6076 = ~n564 & n6075;
  assign n6077 = ~n495 & n6076;
  assign n6078 = ~n591 & n6077;
  assign n6079 = n1717 & n4117;
  assign n6080 = n6072 & n6079;
  assign n6081 = n1717 & n6073;
  assign n6082 = ~n408 & ~n552;
  assign n6083 = n2949 & n6082;
  assign n6084 = n3950 & n6083;
  assign n6085 = n53965 & n6084;
  assign n6086 = ~n852 & n6082;
  assign n6087 = n53908 & n6086;
  assign n6088 = n6070 & n6087;
  assign n6089 = n2949 & n6053;
  assign n6090 = n3950 & n6089;
  assign n6091 = n53965 & n6090;
  assign n6092 = n6088 & n6091;
  assign n6093 = ~n552 & n6053;
  assign n6094 = n53908 & n6093;
  assign n6095 = n6070 & n6094;
  assign n6096 = ~n408 & ~n852;
  assign n6097 = n2949 & n6096;
  assign n6098 = n3950 & n6097;
  assign n6099 = n53965 & n6098;
  assign n6100 = n6095 & n6099;
  assign n6101 = ~n408 & ~n420;
  assign n6102 = ~n354 & n6101;
  assign n6103 = n53908 & n6102;
  assign n6104 = n6070 & n6103;
  assign n6105 = ~n552 & ~n852;
  assign n6106 = n3950 & n6105;
  assign n6107 = n2949 & n6106;
  assign n6108 = n53965 & n6107;
  assign n6109 = n6104 & n6108;
  assign n6110 = n6071 & n6085;
  assign n6111 = ~n623 & ~n627;
  assign n6112 = ~n216 & ~n627;
  assign n6113 = ~n623 & n6112;
  assign n6114 = ~n216 & ~n623;
  assign n6115 = ~n627 & n6114;
  assign n6116 = ~n216 & n6111;
  assign n6117 = ~n510 & ~n567;
  assign n6118 = ~n560 & ~n774;
  assign n6119 = n2477 & n6118;
  assign n6120 = ~n510 & ~n560;
  assign n6121 = ~n567 & ~n774;
  assign n6122 = n6120 & n6121;
  assign n6123 = n2477 & n6122;
  assign n6124 = n6117 & n6119;
  assign n6125 = n2477 & n53967;
  assign n6126 = ~n567 & n6125;
  assign n6127 = ~n560 & n6126;
  assign n6128 = ~n510 & n6127;
  assign n6129 = ~n774 & n6128;
  assign n6130 = n53967 & n53968;
  assign n6131 = n53887 & n53969;
  assign n6132 = n53966 & n6131;
  assign n6133 = n53951 & n6132;
  assign n6134 = n53908 & n53964;
  assign n6135 = n53963 & n6134;
  assign n6136 = n53965 & n6135;
  assign n6137 = n53951 & n6136;
  assign n6138 = n53887 & n6137;
  assign n6139 = n53969 & n6138;
  assign n6140 = n53531 & n6139;
  assign n6141 = n2949 & n6140;
  assign n6142 = n3950 & n6141;
  assign n6143 = ~n408 & n6142;
  assign n6144 = ~n552 & n6143;
  assign n6145 = ~n852 & n6144;
  assign n6146 = ~n420 & n6145;
  assign n6147 = ~n354 & n6146;
  assign n6148 = n53531 & n6133;
  assign n6149 = ~n53962 & ~n53970;
  assign n6150 = ~n275 & ~n346;
  assign n6151 = n589 & n6150;
  assign n6152 = ~n662 & ~n1457;
  assign n6153 = n905 & n6152;
  assign n6154 = n6151 & n6153;
  assign n6155 = ~n443 & ~n612;
  assign n6156 = n2338 & n6155;
  assign n6157 = n53875 & n6156;
  assign n6158 = n53867 & n6157;
  assign n6159 = n589 & n53875;
  assign n6160 = n53867 & n6159;
  assign n6161 = n2338 & n6160;
  assign n6162 = n6150 & n6161;
  assign n6163 = n905 & n6162;
  assign n6164 = ~n662 & n6163;
  assign n6165 = ~n1457 & n6164;
  assign n6166 = ~n612 & n6165;
  assign n6167 = ~n443 & n6166;
  assign n6168 = n905 & n2338;
  assign n6169 = n589 & n2338;
  assign n6170 = n905 & n6150;
  assign n6171 = n6169 & n6170;
  assign n6172 = n2338 & n6150;
  assign n6173 = n589 & n905;
  assign n6174 = n6172 & n6173;
  assign n6175 = n6151 & n6168;
  assign n6176 = ~n443 & ~n662;
  assign n6177 = ~n612 & ~n1457;
  assign n6178 = n6152 & n6155;
  assign n6179 = ~n612 & ~n662;
  assign n6180 = ~n443 & ~n1457;
  assign n6181 = n6179 & n6180;
  assign n6182 = n6176 & n6177;
  assign n6183 = n53867 & n53973;
  assign n6184 = n53875 & n53973;
  assign n6185 = n53867 & n6184;
  assign n6186 = n53875 & n6183;
  assign n6187 = n53972 & n53974;
  assign n6188 = n6154 & n6158;
  assign n6189 = ~n415 & ~n789;
  assign n6190 = ~n415 & ~n1476;
  assign n6191 = ~n789 & n6190;
  assign n6192 = ~n1476 & n6189;
  assign n6193 = n53809 & n53975;
  assign n6194 = ~n896 & ~n902;
  assign n6195 = n712 & ~n902;
  assign n6196 = ~n896 & n6195;
  assign n6197 = n712 & n6194;
  assign n6198 = ~n247 & ~n1127;
  assign n6199 = ~n1127 & n3536;
  assign n6200 = ~n247 & n6199;
  assign n6201 = n3536 & n6198;
  assign n6202 = n53976 & n53977;
  assign n6203 = n6193 & n6202;
  assign n6204 = ~n496 & ~n1469;
  assign n6205 = ~n101 & ~n320;
  assign n6206 = n2094 & n6205;
  assign n6207 = n6204 & n6205;
  assign n6208 = n2094 & n6207;
  assign n6209 = n6204 & n6206;
  assign n6210 = ~n206 & ~n562;
  assign n6211 = n175 & n6210;
  assign n6212 = n4378 & n5733;
  assign n6213 = n6211 & n6212;
  assign n6214 = n175 & n2094;
  assign n6215 = n175 & n6205;
  assign n6216 = n2094 & n6215;
  assign n6217 = n6205 & n6214;
  assign n6218 = n4378 & n6210;
  assign n6219 = n5733 & n6204;
  assign n6220 = n6218 & n6219;
  assign n6221 = n53979 & n6220;
  assign n6222 = n53978 & n6213;
  assign n6223 = ~n414 & ~n788;
  assign n6224 = ~n274 & ~n460;
  assign n6225 = ~n493 & ~n833;
  assign n6226 = ~n460 & ~n493;
  assign n6227 = ~n274 & ~n833;
  assign n6228 = n6226 & n6227;
  assign n6229 = n6224 & n6225;
  assign n6230 = ~n493 & n4094;
  assign n6231 = ~n274 & n6230;
  assign n6232 = ~n460 & n6231;
  assign n6233 = ~n788 & n6232;
  assign n6234 = ~n274 & ~n788;
  assign n6235 = ~n460 & ~n788;
  assign n6236 = ~n274 & ~n493;
  assign n6237 = n6235 & n6236;
  assign n6238 = n6226 & n6234;
  assign n6239 = n4094 & n53983;
  assign n6240 = n6223 & n53981;
  assign n6241 = ~n851 & n3272;
  assign n6242 = n1542 & n3272;
  assign n6243 = ~n851 & n6242;
  assign n6244 = ~n851 & n1542;
  assign n6245 = n3272 & n6244;
  assign n6246 = n1542 & n6241;
  assign n6247 = n53982 & n53984;
  assign n6248 = n53980 & n6247;
  assign n6249 = ~n562 & ~n789;
  assign n6250 = ~n1476 & n6249;
  assign n6251 = n53809 & n6250;
  assign n6252 = n6202 & n6251;
  assign n6253 = ~n206 & ~n415;
  assign n6254 = n175 & n6253;
  assign n6255 = n6212 & n6254;
  assign n6256 = n53978 & n6255;
  assign n6257 = n6247 & n6256;
  assign n6258 = n6252 & n6257;
  assign n6259 = ~n496 & n6249;
  assign n6260 = n53809 & n6259;
  assign n6261 = n6202 & n6260;
  assign n6262 = ~n415 & ~n1469;
  assign n6263 = ~n206 & ~n1476;
  assign n6264 = n6262 & n6263;
  assign n6265 = n6212 & n6264;
  assign n6266 = n53979 & n6265;
  assign n6267 = n6247 & n6266;
  assign n6268 = n6261 & n6267;
  assign n6269 = n6203 & n6248;
  assign n6270 = n53976 & n6205;
  assign n6271 = n53977 & n6270;
  assign n6272 = n5733 & n6271;
  assign n6273 = n53982 & n6272;
  assign n6274 = n53971 & n6273;
  assign n6275 = n53984 & n6274;
  assign n6276 = n53809 & n6275;
  assign n6277 = n4378 & n6276;
  assign n6278 = n175 & n6277;
  assign n6279 = n2094 & n6278;
  assign n6280 = ~n415 & n6279;
  assign n6281 = ~n1469 & n6280;
  assign n6282 = ~n1476 & n6281;
  assign n6283 = ~n206 & n6282;
  assign n6284 = ~n562 & n6283;
  assign n6285 = ~n496 & n6284;
  assign n6286 = ~n789 & n6285;
  assign n6287 = n53971 & n53985;
  assign n6288 = ~n649 & n3214;
  assign n6289 = ~n409 & ~n420;
  assign n6290 = ~n321 & ~n420;
  assign n6291 = ~n409 & n6290;
  assign n6292 = ~n321 & n6289;
  assign n6293 = ~n221 & ~n977;
  assign n6294 = ~n1465 & ~n1477;
  assign n6295 = n6293 & n6294;
  assign n6296 = n53987 & n6295;
  assign n6297 = n6288 & n6295;
  assign n6298 = n53987 & n6297;
  assign n6299 = n6288 & n6296;
  assign n6300 = ~n408 & ~n1059;
  assign n6301 = ~n364 & ~n625;
  assign n6302 = ~n357 & ~n506;
  assign n6303 = n6301 & n6302;
  assign n6304 = ~n506 & n6300;
  assign n6305 = ~n357 & n6304;
  assign n6306 = ~n364 & n6305;
  assign n6307 = ~n625 & n6306;
  assign n6308 = n6300 & n6303;
  assign n6309 = ~n219 & ~n1490;
  assign n6310 = ~n215 & ~n1044;
  assign n6311 = n5021 & n6310;
  assign n6312 = n6309 & n6311;
  assign n6313 = n53989 & n6312;
  assign n6314 = n6293 & n6310;
  assign n6315 = n6288 & n6314;
  assign n6316 = n53987 & n6315;
  assign n6317 = n5021 & n6294;
  assign n6318 = n6309 & n6317;
  assign n6319 = n53989 & n6318;
  assign n6320 = n6316 & n6319;
  assign n6321 = n53988 & n6313;
  assign n6322 = ~n451 & ~n823;
  assign n6323 = ~n105 & ~n614;
  assign n6324 = n1672 & n6323;
  assign n6325 = n6322 & n6324;
  assign n6326 = ~n259 & ~n503;
  assign n6327 = ~n344 & n6326;
  assign n6328 = ~n207 & ~n464;
  assign n6329 = ~n1280 & n6328;
  assign n6330 = n6327 & n6329;
  assign n6331 = n1672 & n6327;
  assign n6332 = ~n464 & n6331;
  assign n6333 = ~n105 & n6332;
  assign n6334 = ~n207 & n6333;
  assign n6335 = ~n1280 & n6334;
  assign n6336 = ~n823 & n6335;
  assign n6337 = ~n451 & n6336;
  assign n6338 = ~n614 & n6337;
  assign n6339 = ~n105 & ~n207;
  assign n6340 = ~n451 & ~n1280;
  assign n6341 = n6339 & n6340;
  assign n6342 = n1672 & n6341;
  assign n6343 = ~n614 & ~n823;
  assign n6344 = ~n464 & n6343;
  assign n6345 = n6327 & n6344;
  assign n6346 = n6342 & n6345;
  assign n6347 = ~n105 & ~n464;
  assign n6348 = ~n614 & ~n1280;
  assign n6349 = n6347 & n6348;
  assign n6350 = n1672 & n6349;
  assign n6351 = ~n207 & ~n451;
  assign n6352 = ~n823 & n6351;
  assign n6353 = n6327 & n6352;
  assign n6354 = n6350 & n6353;
  assign n6355 = n6325 & n6330;
  assign n6356 = ~n319 & ~n553;
  assign n6357 = ~n553 & ~n849;
  assign n6358 = ~n319 & n6357;
  assign n6359 = ~n849 & n6356;
  assign n6360 = ~n246 & ~n659;
  assign n6361 = ~n495 & ~n1881;
  assign n6362 = ~n922 & n6361;
  assign n6363 = ~n495 & ~n659;
  assign n6364 = ~n246 & ~n1881;
  assign n6365 = ~n922 & n6364;
  assign n6366 = n6363 & n6365;
  assign n6367 = ~n922 & ~n1881;
  assign n6368 = ~n246 & ~n495;
  assign n6369 = ~n659 & n6368;
  assign n6370 = n6367 & n6369;
  assign n6371 = ~n659 & ~n1881;
  assign n6372 = ~n922 & n6368;
  assign n6373 = n6371 & n6372;
  assign n6374 = n6360 & n6362;
  assign n6375 = ~n922 & n53992;
  assign n6376 = ~n659 & n6375;
  assign n6377 = ~n246 & n6376;
  assign n6378 = ~n495 & n6377;
  assign n6379 = ~n1881 & n6378;
  assign n6380 = n53992 & n53993;
  assign n6381 = n53991 & n53994;
  assign n6382 = n6288 & n53987;
  assign n6383 = n6309 & n6382;
  assign n6384 = n53989 & n6383;
  assign n6385 = n53991 & n6384;
  assign n6386 = n5021 & n6385;
  assign n6387 = n53994 & n6386;
  assign n6388 = ~n1044 & n6387;
  assign n6389 = ~n977 & n6388;
  assign n6390 = ~n1465 & n6389;
  assign n6391 = ~n1477 & n6390;
  assign n6392 = ~n215 & n6391;
  assign n6393 = ~n221 & n6392;
  assign n6394 = n53990 & n6381;
  assign n6395 = ~n422 & ~n448;
  assign n6396 = ~n444 & ~n975;
  assign n6397 = n4974 & n6396;
  assign n6398 = n4974 & n6395;
  assign n6399 = n6396 & n6398;
  assign n6400 = n6395 & n6397;
  assign n6401 = ~n404 & ~n461;
  assign n6402 = ~n461 & ~n507;
  assign n6403 = ~n404 & n6402;
  assign n6404 = ~n404 & ~n507;
  assign n6405 = ~n461 & n6404;
  assign n6406 = ~n507 & n6401;
  assign n6407 = ~n852 & ~n1715;
  assign n6408 = ~n1090 & n6407;
  assign n6409 = ~n161 & ~n770;
  assign n6410 = n3561 & n6409;
  assign n6411 = n6408 & n6410;
  assign n6412 = n53997 & n6411;
  assign n6413 = n4974 & n53997;
  assign n6414 = n3561 & n6413;
  assign n6415 = ~n422 & n6414;
  assign n6416 = ~n1090 & n6415;
  assign n6417 = ~n161 & n6416;
  assign n6418 = ~n852 & n6417;
  assign n6419 = ~n975 & n6418;
  assign n6420 = ~n444 & n6419;
  assign n6421 = ~n770 & n6420;
  assign n6422 = ~n448 & n6421;
  assign n6423 = ~n1715 & n6422;
  assign n6424 = n3561 & n6396;
  assign n6425 = n6395 & n6424;
  assign n6426 = ~n161 & ~n1090;
  assign n6427 = ~n770 & n6426;
  assign n6428 = n4974 & n6407;
  assign n6429 = n6427 & n6428;
  assign n6430 = n53997 & n6429;
  assign n6431 = n6425 & n6430;
  assign n6432 = ~n1090 & ~n1715;
  assign n6433 = n3561 & n6432;
  assign n6434 = n4974 & n6433;
  assign n6435 = ~n770 & ~n975;
  assign n6436 = ~n444 & n6435;
  assign n6437 = ~n161 & ~n852;
  assign n6438 = n6395 & n6437;
  assign n6439 = n6436 & n6438;
  assign n6440 = n53997 & n6439;
  assign n6441 = n6434 & n6440;
  assign n6442 = n53996 & n6412;
  assign n6443 = ~n222 & ~n552;
  assign n6444 = ~n311 & ~n1492;
  assign n6445 = ~n222 & n6444;
  assign n6446 = ~n552 & n6445;
  assign n6447 = ~n222 & ~n311;
  assign n6448 = ~n552 & ~n1492;
  assign n6449 = n6447 & n6448;
  assign n6450 = ~n311 & ~n552;
  assign n6451 = ~n222 & ~n1492;
  assign n6452 = n6450 & n6451;
  assign n6453 = n6443 & n6444;
  assign n6454 = ~n848 & ~n1189;
  assign n6455 = n2367 & n6454;
  assign n6456 = ~n218 & ~n848;
  assign n6457 = ~n360 & ~n1189;
  assign n6458 = n2815 & n6454;
  assign n6459 = n6456 & n6457;
  assign n6460 = n2367 & n54000;
  assign n6461 = n2815 & n6455;
  assign n6462 = n2367 & n53999;
  assign n6463 = ~n218 & n6462;
  assign n6464 = ~n1189 & n6463;
  assign n6465 = ~n848 & n6464;
  assign n6466 = ~n360 & n6465;
  assign n6467 = n53999 & n54001;
  assign n6468 = ~n292 & ~n356;
  assign n6469 = ~n1641 & n6468;
  assign n6470 = ~n559 & ~n611;
  assign n6471 = n257 & n6470;
  assign n6472 = ~n292 & ~n559;
  assign n6473 = ~n1641 & n6472;
  assign n6474 = ~n356 & ~n611;
  assign n6475 = n257 & n6474;
  assign n6476 = n6473 & n6475;
  assign n6477 = n6469 & n6471;
  assign n6478 = n1036 & n54003;
  assign n6479 = ~n466 & ~n1081;
  assign n6480 = n1488 & n6479;
  assign n6481 = ~n294 & ~n1062;
  assign n6482 = ~n883 & ~n1061;
  assign n6483 = n6481 & n6482;
  assign n6484 = n6480 & n6483;
  assign n6485 = n53878 & n6484;
  assign n6486 = ~n611 & ~n1641;
  assign n6487 = n6472 & n6486;
  assign n6488 = ~n356 & ~n1033;
  assign n6489 = n6482 & n6488;
  assign n6490 = n6480 & n6489;
  assign n6491 = n6487 & n6490;
  assign n6492 = n1035 & n6481;
  assign n6493 = n257 & n6492;
  assign n6494 = n53878 & n6493;
  assign n6495 = n6491 & n6494;
  assign n6496 = ~n292 & ~n1033;
  assign n6497 = n6479 & n6496;
  assign n6498 = ~n559 & ~n1641;
  assign n6499 = n6474 & n6498;
  assign n6500 = n1035 & n6482;
  assign n6501 = n6499 & n6500;
  assign n6502 = n6497 & n6501;
  assign n6503 = n1488 & n6481;
  assign n6504 = n257 & n6503;
  assign n6505 = n53878 & n6504;
  assign n6506 = n6502 & n6505;
  assign n6507 = n6478 & n6485;
  assign n6508 = n54002 & n54004;
  assign n6509 = n53998 & n6508;
  assign n6510 = n53995 & n6509;
  assign n6511 = n257 & n6481;
  assign n6512 = n53878 & n6511;
  assign n6513 = n53995 & n6512;
  assign n6514 = n53998 & n6513;
  assign n6515 = n1488 & n6514;
  assign n6516 = n53986 & n6515;
  assign n6517 = n54002 & n6516;
  assign n6518 = n1035 & n6517;
  assign n6519 = n6482 & n6518;
  assign n6520 = ~n1033 & n6519;
  assign n6521 = ~n1081 & n6520;
  assign n6522 = ~n559 & n6521;
  assign n6523 = ~n292 & n6522;
  assign n6524 = ~n1641 & n6523;
  assign n6525 = ~n611 & n6524;
  assign n6526 = ~n466 & n6525;
  assign n6527 = ~n356 & n6526;
  assign n6528 = n53986 & n6510;
  assign n6529 = ~n53970 & ~n54005;
  assign n6530 = ~n662 & ~n830;
  assign n6531 = n1531 & n5943;
  assign n6532 = n5943 & n6530;
  assign n6533 = n1531 & n6532;
  assign n6534 = n6530 & n6531;
  assign n6535 = ~n361 & ~n1471;
  assign n6536 = ~n849 & ~n2201;
  assign n6537 = ~n849 & n6535;
  assign n6538 = ~n2201 & n6537;
  assign n6539 = n6535 & n6536;
  assign n6540 = ~n216 & ~n564;
  assign n6541 = ~n564 & ~n1769;
  assign n6542 = ~n216 & n6541;
  assign n6543 = ~n1769 & n6540;
  assign n6544 = n53963 & n54008;
  assign n6545 = n54007 & n6544;
  assign n6546 = n1531 & n54007;
  assign n6547 = n53963 & n6546;
  assign n6548 = n6530 & n6547;
  assign n6549 = n5943 & n6548;
  assign n6550 = ~n216 & n6549;
  assign n6551 = ~n564 & n6550;
  assign n6552 = ~n1769 & n6551;
  assign n6553 = n54006 & n6545;
  assign n6554 = n53551 & n5848;
  assign n6555 = ~n553 & ~n584;
  assign n6556 = ~n108 & ~n584;
  assign n6557 = ~n553 & n6556;
  assign n6558 = ~n108 & ~n553;
  assign n6559 = ~n584 & n6558;
  assign n6560 = ~n108 & n6555;
  assign n6561 = n53952 & n54010;
  assign n6562 = n6554 & n6561;
  assign n6563 = ~n311 & ~n894;
  assign n6564 = ~n776 & ~n1191;
  assign n6565 = n6482 & n6564;
  assign n6566 = n6482 & n6563;
  assign n6567 = n6564 & n6566;
  assign n6568 = n6563 & n6565;
  assign n6569 = ~n354 & ~n560;
  assign n6570 = ~n514 & ~n741;
  assign n6571 = ~n560 & ~n741;
  assign n6572 = ~n354 & ~n514;
  assign n6573 = n6571 & n6572;
  assign n6574 = n6569 & n6570;
  assign n6575 = n500 & n3650;
  assign n6576 = n54012 & n6575;
  assign n6577 = ~n184 & ~n1191;
  assign n6578 = n500 & n5277;
  assign n6579 = n6577 & n6578;
  assign n6580 = n6566 & n54012;
  assign n6581 = n6579 & n6580;
  assign n6582 = n54011 & n6576;
  assign n6583 = ~n311 & n6570;
  assign n6584 = n53952 & n6583;
  assign n6585 = n53551 & n54010;
  assign n6586 = n6584 & n6585;
  assign n6587 = n355 & n1672;
  assign n6588 = n6577 & n6587;
  assign n6589 = ~n560 & ~n894;
  assign n6590 = n6482 & n6589;
  assign n6591 = n6578 & n6590;
  assign n6592 = n6588 & n6591;
  assign n6593 = n6586 & n6592;
  assign n6594 = n6562 & n54013;
  assign n6595 = n53551 & n53952;
  assign n6596 = n6577 & n6595;
  assign n6597 = n54010 & n6596;
  assign n6598 = n500 & n6597;
  assign n6599 = n54009 & n6598;
  assign n6600 = n1672 & n6599;
  assign n6601 = n5277 & n6600;
  assign n6602 = n355 & n6601;
  assign n6603 = n6482 & n6602;
  assign n6604 = ~n894 & n6603;
  assign n6605 = ~n311 & n6604;
  assign n6606 = ~n560 & n6605;
  assign n6607 = ~n514 & n6606;
  assign n6608 = ~n741 & n6607;
  assign n6609 = n54009 & n54014;
  assign n6610 = ~n404 & n1659;
  assign n6611 = n1659 & n54015;
  assign n6612 = ~n404 & n6611;
  assign n6613 = n54015 & n6610;
  assign n6614 = ~n466 & ~n922;
  assign n6615 = n5873 & n6614;
  assign n6616 = ~n342 & ~n1703;
  assign n6617 = n164 & ~n1703;
  assign n6618 = ~n342 & n6617;
  assign n6619 = n164 & n6616;
  assign n6620 = ~n249 & ~n1485;
  assign n6621 = ~n420 & n6620;
  assign n6622 = n54017 & n6621;
  assign n6623 = n6615 & n6622;
  assign n6624 = n2674 & n2741;
  assign n6625 = n3950 & n6624;
  assign n6626 = ~n268 & ~n464;
  assign n6627 = ~n1487 & ~n1644;
  assign n6628 = ~n464 & ~n1487;
  assign n6629 = ~n1644 & n6628;
  assign n6630 = ~n268 & n6629;
  assign n6631 = ~n464 & ~n1644;
  assign n6632 = ~n268 & ~n1487;
  assign n6633 = n6631 & n6632;
  assign n6634 = n6626 & n6627;
  assign n6635 = ~n631 & ~n1192;
  assign n6636 = n497 & n6635;
  assign n6637 = n54018 & n6636;
  assign n6638 = n6625 & n6637;
  assign n6639 = n53580 & n53885;
  assign n6640 = n6638 & n6639;
  assign n6641 = n2741 & n6621;
  assign n6642 = n53885 & n6641;
  assign n6643 = n54017 & n6642;
  assign n6644 = n497 & n6643;
  assign n6645 = n54018 & n6644;
  assign n6646 = n53580 & n6645;
  assign n6647 = n6614 & n6646;
  assign n6648 = n3950 & n6647;
  assign n6649 = n5873 & n6648;
  assign n6650 = ~n631 & n6649;
  assign n6651 = ~n1192 & n6650;
  assign n6652 = ~n212 & n6651;
  assign n6653 = ~n423 & n6652;
  assign n6654 = n6615 & n54018;
  assign n6655 = n6621 & n6654;
  assign n6656 = n54017 & n6636;
  assign n6657 = n6625 & n6656;
  assign n6658 = n6639 & n6657;
  assign n6659 = n6655 & n6658;
  assign n6660 = n54017 & n54018;
  assign n6661 = n6621 & n6660;
  assign n6662 = n497 & n6614;
  assign n6663 = n2741 & n6662;
  assign n6664 = n2674 & n6635;
  assign n6665 = n3950 & n5873;
  assign n6666 = n6664 & n6665;
  assign n6667 = n6663 & n6666;
  assign n6668 = n6639 & n6667;
  assign n6669 = n6661 & n6668;
  assign n6670 = n6623 & n6640;
  assign n6671 = n220 & n3536;
  assign n6672 = n906 & n4021;
  assign n6673 = n906 & n3536;
  assign n6674 = n220 & n4021;
  assign n6675 = n6673 & n6674;
  assign n6676 = n6671 & n6672;
  assign n6677 = ~n409 & ~n443;
  assign n6678 = ~n443 & ~n1681;
  assign n6679 = ~n409 & n6678;
  assign n6680 = ~n409 & ~n1681;
  assign n6681 = ~n443 & n6680;
  assign n6682 = ~n1681 & n6677;
  assign n6683 = ~n255 & ~n788;
  assign n6684 = ~n851 & ~n1189;
  assign n6685 = ~n255 & ~n1189;
  assign n6686 = ~n851 & n6685;
  assign n6687 = ~n788 & n6686;
  assign n6688 = ~n788 & ~n851;
  assign n6689 = n6685 & n6688;
  assign n6690 = n6683 & n6684;
  assign n6691 = ~n617 & ~n664;
  assign n6692 = ~n422 & ~n1486;
  assign n6693 = ~n664 & ~n1486;
  assign n6694 = ~n422 & ~n617;
  assign n6695 = n6693 & n6694;
  assign n6696 = n6691 & n6692;
  assign n6697 = n54022 & n54023;
  assign n6698 = n54021 & n6697;
  assign n6699 = ~n218 & ~n617;
  assign n6700 = n3536 & n6699;
  assign n6701 = n6672 & n6700;
  assign n6702 = ~n219 & ~n422;
  assign n6703 = n6693 & n6702;
  assign n6704 = n54022 & n6703;
  assign n6705 = n54021 & n6704;
  assign n6706 = n6701 & n6705;
  assign n6707 = n54020 & n6698;
  assign n6708 = ~n250 & ~n401;
  assign n6709 = n462 & n6708;
  assign n6710 = ~n250 & ~n1065;
  assign n6711 = ~n247 & ~n401;
  assign n6712 = n6710 & n6711;
  assign n6713 = n462 & n6712;
  assign n6714 = n1066 & n6709;
  assign n6715 = ~n172 & ~n647;
  assign n6716 = ~n172 & ~n975;
  assign n6717 = ~n647 & n6716;
  assign n6718 = ~n647 & ~n975;
  assign n6719 = ~n172 & n6718;
  assign n6720 = ~n975 & n6715;
  assign n6721 = ~n168 & ~n465;
  assign n6722 = ~n168 & ~n222;
  assign n6723 = ~n911 & n6722;
  assign n6724 = ~n465 & n6723;
  assign n6725 = n912 & n6721;
  assign n6726 = n54026 & n54027;
  assign n6727 = n462 & n6726;
  assign n6728 = ~n1065 & n6727;
  assign n6729 = ~n250 & n6728;
  assign n6730 = ~n247 & n6729;
  assign n6731 = ~n401 & n6730;
  assign n6732 = n54025 & n6726;
  assign n6733 = ~n612 & ~n1715;
  assign n6734 = ~n405 & ~n740;
  assign n6735 = n5199 & n6734;
  assign n6736 = n5199 & n6733;
  assign n6737 = n6734 & n6736;
  assign n6738 = n6733 & n6735;
  assign n6739 = ~n296 & ~n410;
  assign n6740 = ~n824 & ~n1079;
  assign n6741 = n6739 & n6740;
  assign n6742 = ~n587 & ~n663;
  assign n6743 = n3932 & n6742;
  assign n6744 = ~n410 & ~n587;
  assign n6745 = n6740 & n6744;
  assign n6746 = ~n296 & ~n663;
  assign n6747 = n3932 & n6746;
  assign n6748 = n6745 & n6747;
  assign n6749 = n6741 & n6743;
  assign n6750 = n3932 & n5199;
  assign n6751 = n3932 & n6733;
  assign n6752 = n5199 & n6751;
  assign n6753 = n6733 & n6750;
  assign n6754 = ~n296 & n54031;
  assign n6755 = ~n1079 & n6754;
  assign n6756 = ~n405 & n6755;
  assign n6757 = ~n663 & n6756;
  assign n6758 = ~n824 & n6757;
  assign n6759 = ~n587 & n6758;
  assign n6760 = ~n410 & n6759;
  assign n6761 = ~n740 & n6760;
  assign n6762 = ~n740 & ~n1079;
  assign n6763 = n6739 & n6762;
  assign n6764 = ~n587 & ~n824;
  assign n6765 = ~n405 & ~n663;
  assign n6766 = n6764 & n6765;
  assign n6767 = ~n663 & ~n1079;
  assign n6768 = n6739 & n6767;
  assign n6769 = ~n405 & ~n587;
  assign n6770 = ~n740 & ~n824;
  assign n6771 = n6769 & n6770;
  assign n6772 = n6768 & n6771;
  assign n6773 = n6763 & n6766;
  assign n6774 = n54031 & n54033;
  assign n6775 = n54029 & n54030;
  assign n6776 = n54028 & n54032;
  assign n6777 = n54024 & n6776;
  assign n6778 = n54019 & n6777;
  assign n6779 = n54016 & n54021;
  assign n6780 = n4021 & n6779;
  assign n6781 = n54022 & n6780;
  assign n6782 = n54032 & n6781;
  assign n6783 = n54019 & n6782;
  assign n6784 = n54028 & n6783;
  assign n6785 = n906 & n6784;
  assign n6786 = n3536 & n6785;
  assign n6787 = ~n1486 & n6786;
  assign n6788 = ~n422 & n6787;
  assign n6789 = ~n219 & n6788;
  assign n6790 = ~n218 & n6789;
  assign n6791 = ~n664 & n6790;
  assign n6792 = ~n617 & n6791;
  assign n6793 = n54016 & n6778;
  assign n6794 = ~n54005 & ~n54034;
  assign n6795 = ~n405 & ~n590;
  assign n6796 = ~n405 & n2974;
  assign n6797 = ~n590 & n6796;
  assign n6798 = n2974 & n6795;
  assign n6799 = ~n105 & ~n646;
  assign n6800 = ~n1337 & n6799;
  assign n6801 = n6288 & n6800;
  assign n6802 = n54035 & n6800;
  assign n6803 = n6288 & n6802;
  assign n6804 = n54035 & n6801;
  assign n6805 = n964 & n4470;
  assign n6806 = ~n219 & ~n441;
  assign n6807 = n6535 & n6806;
  assign n6808 = n6805 & n6807;
  assign n6809 = n343 & n2367;
  assign n6810 = n3776 & n4364;
  assign n6811 = n6809 & n6810;
  assign n6812 = n3776 & n6806;
  assign n6813 = n6805 & n6812;
  assign n6814 = n2367 & n4364;
  assign n6815 = n343 & n6535;
  assign n6816 = n6814 & n6815;
  assign n6817 = n6813 & n6816;
  assign n6818 = n6808 & n6811;
  assign n6819 = n755 & ~n1455;
  assign n6820 = n755 & n5874;
  assign n6821 = ~n1455 & n6820;
  assign n6822 = ~n1455 & n5874;
  assign n6823 = n755 & n6822;
  assign n6824 = n5874 & n6819;
  assign n6825 = n53611 & n54038;
  assign n6826 = n54037 & n6825;
  assign n6827 = ~n646 & ~n1337;
  assign n6828 = ~n451 & n6827;
  assign n6829 = n6288 & n6828;
  assign n6830 = n54035 & n6829;
  assign n6831 = n343 & n964;
  assign n6832 = n3776 & n6535;
  assign n6833 = n6831 & n6832;
  assign n6834 = ~n105 & ~n513;
  assign n6835 = n6806 & n6834;
  assign n6836 = n2367 & n4470;
  assign n6837 = n6835 & n6836;
  assign n6838 = n6833 & n6837;
  assign n6839 = n6825 & n6838;
  assign n6840 = n6830 & n6839;
  assign n6841 = n54036 & n6826;
  assign n6842 = n6288 & n54038;
  assign n6843 = n54035 & n6842;
  assign n6844 = n964 & n6843;
  assign n6845 = n4470 & n6844;
  assign n6846 = n53611 & n6845;
  assign n6847 = n343 & n6846;
  assign n6848 = n53998 & n6847;
  assign n6849 = n6806 & n6848;
  assign n6850 = n6535 & n6849;
  assign n6851 = n2367 & n6850;
  assign n6852 = n3776 & n6851;
  assign n6853 = ~n105 & n6852;
  assign n6854 = ~n1337 & n6853;
  assign n6855 = ~n513 & n6854;
  assign n6856 = ~n451 & n6855;
  assign n6857 = ~n646 & n6856;
  assign n6858 = n53998 & n54039;
  assign n6859 = n2053 & n6614;
  assign n6860 = ~n631 & ~n740;
  assign n6861 = n2092 & n6860;
  assign n6862 = n2092 & n6614;
  assign n6863 = n2053 & n6860;
  assign n6864 = n6862 & n6863;
  assign n6865 = n6859 & n6861;
  assign n6866 = ~n2201 & n4002;
  assign n6867 = ~n269 & ~n1088;
  assign n6868 = ~n1059 & ~n1088;
  assign n6869 = ~n269 & n6868;
  assign n6870 = ~n269 & ~n1059;
  assign n6871 = ~n1088 & n6870;
  assign n6872 = ~n1059 & n6867;
  assign n6873 = ~n274 & ~n848;
  assign n6874 = n2852 & n6873;
  assign n6875 = n54042 & n6874;
  assign n6876 = ~n822 & ~n2201;
  assign n6877 = ~n274 & n6876;
  assign n6878 = ~n409 & ~n848;
  assign n6879 = n4002 & n6878;
  assign n6880 = n6866 & n6874;
  assign n6881 = n6877 & n6879;
  assign n6882 = n54042 & n54043;
  assign n6883 = n6866 & n6875;
  assign n6884 = n2053 & n2852;
  assign n6885 = n6862 & n6884;
  assign n6886 = n6860 & n6873;
  assign n6887 = n54042 & n6886;
  assign n6888 = n6866 & n6887;
  assign n6889 = n6885 & n6888;
  assign n6890 = n54041 & n54044;
  assign n6891 = ~n319 & ~n360;
  assign n6892 = ~n360 & ~n493;
  assign n6893 = ~n319 & n6892;
  assign n6894 = ~n319 & ~n493;
  assign n6895 = ~n360 & n6894;
  assign n6896 = ~n493 & n6891;
  assign n6897 = ~n459 & ~n1486;
  assign n6898 = n421 & n2093;
  assign n6899 = n2093 & n6897;
  assign n6900 = n421 & n6899;
  assign n6901 = n6897 & n6898;
  assign n6902 = ~n493 & n54047;
  assign n6903 = ~n319 & n6902;
  assign n6904 = ~n360 & n6903;
  assign n6905 = n54046 & n54047;
  assign n6906 = n53572 & n54048;
  assign n6907 = n53572 & n53601;
  assign n6908 = n54048 & n6907;
  assign n6909 = n53601 & n6906;
  assign n6910 = n54045 & n54049;
  assign n6911 = n53591 & n6910;
  assign n6912 = n6863 & n54048;
  assign n6913 = n54040 & n6912;
  assign n6914 = n53601 & n6913;
  assign n6915 = n53572 & n6914;
  assign n6916 = n53591 & n6915;
  assign n6917 = n2092 & n6916;
  assign n6918 = n54042 & n6917;
  assign n6919 = n4002 & n6918;
  assign n6920 = n6614 & n6919;
  assign n6921 = ~n848 & n6920;
  assign n6922 = ~n822 & n6921;
  assign n6923 = ~n274 & n6922;
  assign n6924 = ~n409 & n6923;
  assign n6925 = ~n2201 & n6924;
  assign n6926 = n54040 & n6910;
  assign n6927 = n53591 & n6926;
  assign n6928 = n54040 & n6911;
  assign n6929 = ~n54034 & ~n54050;
  assign n6930 = n2454 & n2949;
  assign n6931 = n2949 & n2975;
  assign n6932 = n2454 & n6931;
  assign n6933 = n2975 & n6930;
  assign n6934 = n347 & ~n1658;
  assign n6935 = ~n310 & ~n788;
  assign n6936 = ~n310 & ~n902;
  assign n6937 = ~n788 & n6936;
  assign n6938 = ~n788 & ~n902;
  assign n6939 = ~n310 & n6938;
  assign n6940 = ~n902 & n6935;
  assign n6941 = n53809 & n54052;
  assign n6942 = n6934 & n6941;
  assign n6943 = n2454 & n6934;
  assign n6944 = n2949 & n6943;
  assign n6945 = n2975 & n6944;
  assign n6946 = n53809 & n6945;
  assign n6947 = ~n902 & n6946;
  assign n6948 = ~n310 & n6947;
  assign n6949 = ~n788 & n6948;
  assign n6950 = n54051 & n6942;
  assign n6951 = n3819 & n4261;
  assign n6952 = n814 & n5021;
  assign n6953 = n6951 & n6952;
  assign n6954 = ~n562 & ~n1491;
  assign n6955 = ~n1196 & ~n1466;
  assign n6956 = ~n1466 & ~n1491;
  assign n6957 = ~n562 & ~n1196;
  assign n6958 = n6956 & n6957;
  assign n6959 = n6954 & n6955;
  assign n6960 = n3389 & n3670;
  assign n6961 = n54054 & n6960;
  assign n6962 = ~n419 & ~n459;
  assign n6963 = ~n419 & ~n742;
  assign n6964 = ~n459 & n6963;
  assign n6965 = ~n459 & ~n742;
  assign n6966 = ~n419 & n6965;
  assign n6967 = ~n742 & n6962;
  assign n6968 = n54007 & n54055;
  assign n6969 = n6961 & n6968;
  assign n6970 = n3670 & n3819;
  assign n6971 = n4261 & n5021;
  assign n6972 = n6970 & n6971;
  assign n6973 = n814 & n3389;
  assign n6974 = n54054 & n6973;
  assign n6975 = n6968 & n6974;
  assign n6976 = n6972 & n6975;
  assign n6977 = n814 & n3670;
  assign n6978 = n3819 & n5021;
  assign n6979 = n6977 & n6978;
  assign n6980 = n6952 & n6970;
  assign n6981 = n3389 & n4261;
  assign n6982 = n54054 & n6981;
  assign n6983 = n6968 & n6982;
  assign n6984 = n54057 & n6983;
  assign n6985 = n6953 & n6969;
  assign n6986 = n3819 & n6968;
  assign n6987 = n54053 & n6986;
  assign n6988 = n814 & n6987;
  assign n6989 = n4261 & n6988;
  assign n6990 = n3670 & n6989;
  assign n6991 = n5021 & n6990;
  assign n6992 = n3389 & n6991;
  assign n6993 = ~n1466 & n6992;
  assign n6994 = ~n1491 & n6993;
  assign n6995 = ~n1196 & n6994;
  assign n6996 = ~n562 & n6995;
  assign n6997 = n54053 & n54056;
  assign n6998 = ~n256 & ~n564;
  assign n6999 = ~n911 & ~n1189;
  assign n7000 = ~n564 & ~n911;
  assign n7001 = ~n256 & ~n1189;
  assign n7002 = n7000 & n7001;
  assign n7003 = n6998 & n6999;
  assign n7004 = ~n498 & ~n628;
  assign n7005 = ~n1090 & ~n1478;
  assign n7006 = n4376 & n7005;
  assign n7007 = n7004 & n7005;
  assign n7008 = n4376 & n7007;
  assign n7009 = n7004 & n7006;
  assign n7010 = ~n256 & n54060;
  assign n7011 = ~n564 & n7010;
  assign n7012 = ~n1189 & n7011;
  assign n7013 = ~n911 & n7012;
  assign n7014 = n54059 & n54060;
  assign n7015 = ~n161 & ~n423;
  assign n7016 = ~n409 & ~n1062;
  assign n7017 = n7015 & n7016;
  assign n7018 = ~n275 & ~n554;
  assign n7019 = n1936 & n7018;
  assign n7020 = n1936 & n7016;
  assign n7021 = n7015 & n7018;
  assign n7022 = n7020 & n7021;
  assign n7023 = n7017 & n7019;
  assign n7024 = ~n852 & ~n1065;
  assign n7025 = ~n410 & n7024;
  assign n7026 = n2102 & n5157;
  assign n7027 = n7025 & n7026;
  assign n7028 = n2102 & n7018;
  assign n7029 = n7020 & n7028;
  assign n7030 = ~n161 & ~n776;
  assign n7031 = ~n423 & ~n611;
  assign n7032 = n7030 & n7031;
  assign n7033 = n7025 & n7032;
  assign n7034 = n7029 & n7033;
  assign n7035 = ~n161 & ~n611;
  assign n7036 = ~n776 & ~n1124;
  assign n7037 = n7035 & n7036;
  assign n7038 = ~n423 & ~n568;
  assign n7039 = n7016 & n7038;
  assign n7040 = n7037 & n7039;
  assign n7041 = n7025 & n7028;
  assign n7042 = n7040 & n7041;
  assign n7043 = n54062 & n7027;
  assign n7044 = ~n567 & ~n1034;
  assign n7045 = ~n450 & ~n1280;
  assign n7046 = ~n292 & ~n415;
  assign n7047 = n7045 & n7046;
  assign n7048 = ~n415 & n7045;
  assign n7049 = ~n567 & n7048;
  assign n7050 = ~n292 & n7049;
  assign n7051 = ~n1034 & n7050;
  assign n7052 = ~n415 & ~n1034;
  assign n7053 = ~n292 & ~n567;
  assign n7054 = n7052 & n7053;
  assign n7055 = n7045 & n7054;
  assign n7056 = n7044 & n7047;
  assign n7057 = ~n590 & ~n614;
  assign n7058 = ~n493 & ~n1127;
  assign n7059 = ~n1127 & ~n1703;
  assign n7060 = ~n493 & n7059;
  assign n7061 = ~n1703 & n7058;
  assign n7062 = ~n614 & n54065;
  assign n7063 = ~n590 & n7062;
  assign n7064 = ~n493 & ~n614;
  assign n7065 = ~n590 & ~n1703;
  assign n7066 = ~n1127 & n7065;
  assign n7067 = n7064 & n7066;
  assign n7068 = ~n614 & ~n1127;
  assign n7069 = ~n493 & n7068;
  assign n7070 = n7065 & n7069;
  assign n7071 = ~n614 & ~n1703;
  assign n7072 = ~n590 & n7058;
  assign n7073 = n7071 & n7072;
  assign n7074 = n7057 & n54065;
  assign n7075 = n54064 & n54066;
  assign n7076 = n54063 & n7075;
  assign n7077 = n7025 & n54066;
  assign n7078 = n54064 & n7077;
  assign n7079 = n54061 & n7078;
  assign n7080 = n7016 & n7079;
  assign n7081 = ~n1124 & n7080;
  assign n7082 = ~n1486 & n7081;
  assign n7083 = ~n161 & n7082;
  assign n7084 = ~n568 & n7083;
  assign n7085 = ~n554 & n7084;
  assign n7086 = ~n275 & n7085;
  assign n7087 = ~n611 & n7086;
  assign n7088 = ~n423 & n7087;
  assign n7089 = ~n360 & n7088;
  assign n7090 = ~n776 & n7089;
  assign n7091 = n54061 & n7076;
  assign n7092 = ~n560 & ~n1059;
  assign n7093 = ~n443 & ~n1081;
  assign n7094 = ~n956 & ~n1195;
  assign n7095 = n7093 & n7094;
  assign n7096 = n7092 & n7095;
  assign n7097 = n3561 & n3671;
  assign n7098 = n4530 & n6734;
  assign n7099 = n7097 & n7098;
  assign n7100 = n7096 & n7099;
  assign n7101 = ~n848 & ~n922;
  assign n7102 = ~n552 & ~n659;
  assign n7103 = ~n747 & ~n1079;
  assign n7104 = ~n659 & ~n1079;
  assign n7105 = ~n552 & ~n747;
  assign n7106 = n7104 & n7105;
  assign n7107 = n7102 & n7103;
  assign n7108 = ~n1079 & n7101;
  assign n7109 = ~n659 & n7108;
  assign n7110 = ~n552 & n7109;
  assign n7111 = ~n747 & n7110;
  assign n7112 = n7101 & n54068;
  assign n7113 = ~n212 & ~n495;
  assign n7114 = ~n495 & n53765;
  assign n7115 = n2338 & n7113;
  assign n7116 = n54069 & n54070;
  assign n7117 = n7100 & n7116;
  assign n7118 = ~n105 & ~n1088;
  assign n7119 = ~n461 & n7118;
  assign n7120 = ~n465 & n7119;
  assign n7121 = ~n105 & ~n465;
  assign n7122 = ~n461 & ~n1088;
  assign n7123 = n7121 & n7122;
  assign n7124 = n1760 & n7118;
  assign n7125 = n175 & ~n340;
  assign n7126 = n1274 & n3475;
  assign n7127 = n7125 & n7126;
  assign n7128 = n54071 & n7127;
  assign n7129 = n53869 & n7128;
  assign n7130 = ~n560 & ~n664;
  assign n7131 = ~n460 & ~n1059;
  assign n7132 = n7130 & n7131;
  assign n7133 = n7093 & n7132;
  assign n7134 = n3561 & n4530;
  assign n7135 = n6734 & n7094;
  assign n7136 = n7134 & n7135;
  assign n7137 = n7133 & n7136;
  assign n7138 = n7116 & n7137;
  assign n7139 = n3475 & n3671;
  assign n7140 = n7125 & n7139;
  assign n7141 = n54071 & n7140;
  assign n7142 = n53869 & n7141;
  assign n7143 = n7138 & n7142;
  assign n7144 = ~n460 & ~n1081;
  assign n7145 = n175 & n7094;
  assign n7146 = n7144 & n7145;
  assign n7147 = n3475 & n7130;
  assign n7148 = n3671 & n4530;
  assign n7149 = n7147 & n7148;
  assign n7150 = n7146 & n7149;
  assign n7151 = n7116 & n7150;
  assign n7152 = ~n443 & ~n1059;
  assign n7153 = ~n740 & n7152;
  assign n7154 = ~n340 & ~n405;
  assign n7155 = n3561 & n7154;
  assign n7156 = n7153 & n7155;
  assign n7157 = n54071 & n7156;
  assign n7158 = n53869 & n7157;
  assign n7159 = n7151 & n7158;
  assign n7160 = n3671 & n7144;
  assign n7161 = n7130 & n7160;
  assign n7162 = n175 & n3475;
  assign n7163 = n7134 & n7162;
  assign n7164 = n7161 & n7163;
  assign n7165 = n54069 & n7164;
  assign n7166 = ~n740 & ~n1195;
  assign n7167 = ~n956 & n7166;
  assign n7168 = ~n340 & ~n1059;
  assign n7169 = ~n405 & ~n443;
  assign n7170 = n7168 & n7169;
  assign n7171 = n7167 & n7170;
  assign n7172 = n54070 & n54071;
  assign n7173 = n7171 & n7172;
  assign n7174 = n53869 & n7173;
  assign n7175 = n7165 & n7174;
  assign n7176 = n7117 & n7129;
  assign n7177 = n54067 & n54072;
  assign n7178 = n54070 & n7130;
  assign n7179 = n54071 & n7178;
  assign n7180 = n54069 & n7179;
  assign n7181 = n54067 & n7180;
  assign n7182 = n3671 & n7181;
  assign n7183 = n54058 & n7182;
  assign n7184 = n7144 & n7183;
  assign n7185 = n4530 & n7184;
  assign n7186 = n53869 & n7185;
  assign n7187 = n175 & n7186;
  assign n7188 = n3475 & n7187;
  assign n7189 = n3561 & n7188;
  assign n7190 = ~n1195 & n7189;
  assign n7191 = ~n405 & n7190;
  assign n7192 = ~n1059 & n7191;
  assign n7193 = ~n956 & n7192;
  assign n7194 = ~n443 & n7193;
  assign n7195 = ~n340 & n7194;
  assign n7196 = ~n740 & n7195;
  assign n7197 = n54058 & n54072;
  assign n7198 = n54067 & n7197;
  assign n7199 = n54058 & n7177;
  assign n7200 = ~n54050 & ~n54073;
  assign n7201 = ~n568 & ~n631;
  assign n7202 = ~n466 & ~n591;
  assign n7203 = n5180 & n7202;
  assign n7204 = n7201 & n7203;
  assign n7205 = ~n1042 & ~n1455;
  assign n7206 = ~n894 & ~n1769;
  assign n7207 = n7205 & n7206;
  assign n7208 = n54042 & n7207;
  assign n7209 = ~n499 & ~n625;
  assign n7210 = ~n625 & n5203;
  assign n7211 = ~n788 & n7209;
  assign n7212 = ~n1065 & n5390;
  assign n7213 = n54074 & n7212;
  assign n7214 = n7208 & n7213;
  assign n7215 = n53883 & n54074;
  assign n7216 = n5390 & n7215;
  assign n7217 = n54042 & n7216;
  assign n7218 = n7201 & n7217;
  assign n7219 = ~n1065 & n7218;
  assign n7220 = ~n1455 & n7219;
  assign n7221 = ~n1042 & n7220;
  assign n7222 = ~n591 & n7221;
  assign n7223 = ~n466 & n7222;
  assign n7224 = ~n1769 & n7223;
  assign n7225 = n5180 & n5390;
  assign n7226 = n7201 & n7225;
  assign n7227 = n54042 & n54074;
  assign n7228 = ~n466 & ~n1769;
  assign n7229 = ~n591 & n7228;
  assign n7230 = ~n894 & ~n1455;
  assign n7231 = ~n1042 & ~n1065;
  assign n7232 = n7230 & n7231;
  assign n7233 = n7229 & n7232;
  assign n7234 = n7227 & n7233;
  assign n7235 = n7226 & n7234;
  assign n7236 = ~n591 & ~n1065;
  assign n7237 = n5390 & n7236;
  assign n7238 = n7201 & n7237;
  assign n7239 = n7205 & n7228;
  assign n7240 = n53883 & n7239;
  assign n7241 = n7227 & n7240;
  assign n7242 = n7238 & n7241;
  assign n7243 = n7204 & n7214;
  assign n7244 = ~n275 & ~n622;
  assign n7245 = ~n258 & ~n275;
  assign n7246 = ~n622 & n7245;
  assign n7247 = ~n258 & ~n622;
  assign n7248 = ~n275 & n7247;
  assign n7249 = ~n258 & n7244;
  assign n7250 = ~n141 & ~n651;
  assign n7251 = ~n141 & n1956;
  assign n7252 = ~n651 & n7251;
  assign n7253 = n1956 & n7250;
  assign n7254 = ~n268 & ~n627;
  assign n7255 = n1076 & n7254;
  assign n7256 = n54077 & n7255;
  assign n7257 = n54076 & n7256;
  assign n7258 = ~n291 & ~n553;
  assign n7259 = ~n491 & ~n852;
  assign n7260 = ~n1476 & n7259;
  assign n7261 = ~n291 & ~n1476;
  assign n7262 = ~n553 & n7261;
  assign n7263 = ~n852 & n7262;
  assign n7264 = ~n491 & n7263;
  assign n7265 = ~n291 & ~n491;
  assign n7266 = ~n553 & ~n852;
  assign n7267 = ~n1476 & n7266;
  assign n7268 = n7265 & n7267;
  assign n7269 = n7259 & n7262;
  assign n7270 = ~n291 & ~n852;
  assign n7271 = ~n553 & ~n1476;
  assign n7272 = ~n491 & n7271;
  assign n7273 = n7270 & n7272;
  assign n7274 = n7258 & n7260;
  assign n7275 = ~n408 & ~n2201;
  assign n7276 = ~n588 & ~n617;
  assign n7277 = ~n562 & ~n1472;
  assign n7278 = n7276 & n7277;
  assign n7279 = n7275 & n7276;
  assign n7280 = n7277 & n7279;
  assign n7281 = n7275 & n7278;
  assign n7282 = n54078 & n54079;
  assign n7283 = ~n627 & ~n1472;
  assign n7284 = ~n268 & ~n562;
  assign n7285 = n7254 & n7277;
  assign n7286 = n7283 & n7284;
  assign n7287 = n54077 & n54080;
  assign n7288 = n54076 & n7287;
  assign n7289 = n1076 & n7276;
  assign n7290 = n7275 & n7289;
  assign n7291 = n54078 & n7290;
  assign n7292 = n7288 & n7291;
  assign n7293 = n7257 & n7282;
  assign n7294 = n53718 & n54081;
  assign n7295 = n54076 & n54077;
  assign n7296 = n1076 & n7295;
  assign n7297 = n7275 & n7296;
  assign n7298 = n54078 & n7297;
  assign n7299 = n53718 & n7298;
  assign n7300 = n54075 & n7299;
  assign n7301 = n7276 & n7300;
  assign n7302 = ~n1472 & n7301;
  assign n7303 = ~n562 & n7302;
  assign n7304 = ~n268 & n7303;
  assign n7305 = ~n627 & n7304;
  assign n7306 = n54075 & n7294;
  assign n7307 = ~n630 & ~n832;
  assign n7308 = ~n207 & ~n1646;
  assign n7309 = n1819 & n7308;
  assign n7310 = n7307 & n7309;
  assign n7311 = ~n402 & ~n1681;
  assign n7312 = ~n1191 & n7311;
  assign n7313 = n976 & n6309;
  assign n7314 = n7312 & n7313;
  assign n7315 = n7307 & n7313;
  assign n7316 = ~n402 & ~n1191;
  assign n7317 = ~n565 & n7316;
  assign n7318 = ~n735 & ~n1681;
  assign n7319 = n7308 & n7318;
  assign n7320 = n7317 & n7319;
  assign n7321 = n7315 & n7320;
  assign n7322 = n7310 & n7314;
  assign n7323 = n6309 & n7307;
  assign n7324 = n54082 & n7323;
  assign n7325 = n976 & n7324;
  assign n7326 = ~n1681 & n7325;
  assign n7327 = ~n1191 & n7326;
  assign n7328 = ~n207 & n7327;
  assign n7329 = ~n565 & n7328;
  assign n7330 = ~n402 & n7329;
  assign n7331 = ~n1646 & n7330;
  assign n7332 = ~n735 & n7331;
  assign n7333 = n54082 & n54083;
  assign n7334 = ~n443 & ~n464;
  assign n7335 = ~n1196 & ~n1469;
  assign n7336 = n7334 & n7335;
  assign n7337 = ~n174 & ~n308;
  assign n7338 = n561 & n7337;
  assign n7339 = n7335 & n7337;
  assign n7340 = n561 & n7334;
  assign n7341 = n7339 & n7340;
  assign n7342 = n7336 & n7338;
  assign n7343 = ~n663 & ~n747;
  assign n7344 = ~n663 & n7005;
  assign n7345 = ~n747 & n7344;
  assign n7346 = n7005 & n7343;
  assign n7347 = n54027 & n54086;
  assign n7348 = n54085 & n7347;
  assign n7349 = n2916 & n4319;
  assign n7350 = ~n292 & ~n833;
  assign n7351 = n1532 & n7350;
  assign n7352 = n7349 & n7351;
  assign n7353 = n53542 & n7352;
  assign n7354 = n53510 & n7353;
  assign n7355 = n1532 & n2916;
  assign n7356 = n7350 & n7355;
  assign n7357 = n54086 & n7356;
  assign n7358 = n54027 & n7357;
  assign n7359 = n53510 & n7358;
  assign n7360 = n53542 & n7359;
  assign n7361 = n561 & n7360;
  assign n7362 = n4319 & n7361;
  assign n7363 = ~n464 & n7362;
  assign n7364 = ~n1469 & n7363;
  assign n7365 = ~n1196 & n7364;
  assign n7366 = ~n174 & n7365;
  assign n7367 = ~n308 & n7366;
  assign n7368 = ~n443 & n7367;
  assign n7369 = ~n443 & ~n1469;
  assign n7370 = ~n308 & ~n1196;
  assign n7371 = n7369 & n7370;
  assign n7372 = ~n174 & ~n464;
  assign n7373 = n4319 & n7372;
  assign n7374 = ~n308 & ~n464;
  assign n7375 = n7369 & n7374;
  assign n7376 = ~n174 & ~n1196;
  assign n7377 = n4319 & n7376;
  assign n7378 = n7375 & n7377;
  assign n7379 = n7371 & n7373;
  assign n7380 = n7347 & n54088;
  assign n7381 = n561 & n7350;
  assign n7382 = n561 & n2916;
  assign n7383 = n7351 & n7382;
  assign n7384 = n7355 & n7381;
  assign n7385 = n53542 & n54089;
  assign n7386 = n53510 & n7385;
  assign n7387 = n7380 & n7386;
  assign n7388 = n7348 & n7354;
  assign n7389 = ~n342 & ~n420;
  assign n7390 = ~n342 & ~n1658;
  assign n7391 = ~n420 & n7390;
  assign n7392 = ~n420 & ~n1658;
  assign n7393 = ~n342 & n7392;
  assign n7394 = ~n1658 & n7389;
  assign n7395 = ~n415 & ~n957;
  assign n7396 = ~n415 & ~n984;
  assign n7397 = ~n957 & n7396;
  assign n7398 = ~n984 & n7395;
  assign n7399 = n53997 & n54091;
  assign n7400 = n53997 & n54090;
  assign n7401 = ~n984 & n7400;
  assign n7402 = ~n415 & n7401;
  assign n7403 = ~n957 & n7402;
  assign n7404 = n54090 & n7399;
  assign n7405 = ~n742 & ~n748;
  assign n7406 = ~n742 & ~n774;
  assign n7407 = ~n748 & n7406;
  assign n7408 = ~n774 & n7405;
  assign n7409 = ~n256 & ~n618;
  assign n7410 = n2333 & n7409;
  assign n7411 = n54093 & n7410;
  assign n7412 = ~n948 & ~n1061;
  assign n7413 = n850 & ~n948;
  assign n7414 = ~n1061 & n7413;
  assign n7415 = n850 & n7412;
  assign n7416 = n4915 & n54094;
  assign n7417 = n7411 & n7416;
  assign n7418 = ~n144 & ~n296;
  assign n7419 = ~n410 & ~n585;
  assign n7420 = ~n504 & ~n1644;
  assign n7421 = ~n410 & ~n504;
  assign n7422 = ~n585 & ~n1644;
  assign n7423 = n7421 & n7422;
  assign n7424 = n7419 & n7420;
  assign n7425 = ~n504 & n7418;
  assign n7426 = ~n1644 & n7425;
  assign n7427 = ~n410 & n7426;
  assign n7428 = ~n585 & n7427;
  assign n7429 = n7418 & n54095;
  assign n7430 = n1128 & n2914;
  assign n7431 = n1078 & n7430;
  assign n7432 = n54096 & n7431;
  assign n7433 = n1128 & n7409;
  assign n7434 = n54093 & n7433;
  assign n7435 = n7416 & n7434;
  assign n7436 = n2333 & n2914;
  assign n7437 = n1078 & n7436;
  assign n7438 = n54096 & n7437;
  assign n7439 = n7435 & n7438;
  assign n7440 = n2914 & n7405;
  assign n7441 = n4915 & n7440;
  assign n7442 = ~n256 & ~n774;
  assign n7443 = ~n618 & n7442;
  assign n7444 = n54094 & n7443;
  assign n7445 = n7441 & n7444;
  assign n7446 = n1078 & n1128;
  assign n7447 = n2333 & n7446;
  assign n7448 = n54096 & n7447;
  assign n7449 = n7445 & n7448;
  assign n7450 = n7417 & n7432;
  assign n7451 = n54092 & n54097;
  assign n7452 = n54087 & n7451;
  assign n7453 = n2333 & n54094;
  assign n7454 = n4914 & n7453;
  assign n7455 = n54096 & n7454;
  assign n7456 = n54087 & n7455;
  assign n7457 = n1078 & n7456;
  assign n7458 = n54092 & n7457;
  assign n7459 = n54084 & n7458;
  assign n7460 = n1128 & n7459;
  assign n7461 = n2367 & n7460;
  assign n7462 = ~n1680 & n7461;
  assign n7463 = ~n256 & n7462;
  assign n7464 = ~n618 & n7463;
  assign n7465 = ~n742 & n7464;
  assign n7466 = ~n748 & n7465;
  assign n7467 = ~n774 & n7466;
  assign n7468 = ~n623 & n7467;
  assign n7469 = n54084 & n7452;
  assign n7470 = ~n54073 & ~n54098;
  assign n7471 = ~n650 & ~n789;
  assign n7472 = n7276 & n7471;
  assign n7473 = ~n174 & ~n221;
  assign n7474 = n1957 & n7473;
  assign n7475 = n7472 & n7474;
  assign n7476 = ~n184 & ~n466;
  assign n7477 = ~n1337 & n7476;
  assign n7478 = n2058 & n2925;
  assign n7479 = n7477 & n7478;
  assign n7480 = n1957 & n2058;
  assign n7481 = n7276 & n7473;
  assign n7482 = n1957 & n7481;
  assign n7483 = n2058 & n7482;
  assign n7484 = n2058 & n7276;
  assign n7485 = n7474 & n7484;
  assign n7486 = n7480 & n7481;
  assign n7487 = ~n184 & n54099;
  assign n7488 = ~n246 & n7487;
  assign n7489 = ~n1337 & n7488;
  assign n7490 = ~n466 & n7489;
  assign n7491 = ~n650 & n7490;
  assign n7492 = ~n789 & n7491;
  assign n7493 = ~n614 & n7492;
  assign n7494 = ~n246 & ~n466;
  assign n7495 = ~n184 & n7494;
  assign n7496 = ~n614 & ~n1337;
  assign n7497 = n7471 & n7496;
  assign n7498 = ~n789 & n2925;
  assign n7499 = ~n650 & ~n1337;
  assign n7500 = n7476 & n7499;
  assign n7501 = n7498 & n7500;
  assign n7502 = n7495 & n7497;
  assign n7503 = n54099 & n54101;
  assign n7504 = n7475 & n7479;
  assign n7505 = ~n662 & ~n894;
  assign n7506 = n2577 & n7505;
  assign n7507 = n1277 & n3217;
  assign n7508 = n3670 & n4026;
  assign n7509 = n7507 & n7508;
  assign n7510 = n7506 & n7509;
  assign n7511 = ~n317 & ~n1492;
  assign n7512 = n2675 & n7511;
  assign n7513 = ~n498 & ~n957;
  assign n7514 = n3000 & n7513;
  assign n7515 = n2675 & n3000;
  assign n7516 = ~n957 & n7515;
  assign n7517 = ~n1492 & n7516;
  assign n7518 = ~n317 & n7517;
  assign n7519 = ~n498 & n7518;
  assign n7520 = ~n317 & ~n957;
  assign n7521 = ~n498 & ~n1492;
  assign n7522 = n7520 & n7521;
  assign n7523 = n7515 & n7522;
  assign n7524 = n7512 & n7514;
  assign n7525 = ~n108 & ~n420;
  assign n7526 = ~n1127 & ~n1487;
  assign n7527 = n1671 & n7526;
  assign n7528 = n7525 & n7527;
  assign n7529 = n54102 & n7528;
  assign n7530 = ~n108 & ~n662;
  assign n7531 = ~n420 & ~n894;
  assign n7532 = n7530 & n7531;
  assign n7533 = n1277 & n2577;
  assign n7534 = n3217 & n3670;
  assign n7535 = n7533 & n7534;
  assign n7536 = n7532 & n7535;
  assign n7537 = n1671 & n4026;
  assign n7538 = n7526 & n7537;
  assign n7539 = n54102 & n7538;
  assign n7540 = n7536 & n7539;
  assign n7541 = n7525 & n7526;
  assign n7542 = n3217 & n4026;
  assign n7543 = n7506 & n7542;
  assign n7544 = n7541 & n7543;
  assign n7545 = n1277 & n1671;
  assign n7546 = n3670 & n7545;
  assign n7547 = n54102 & n7546;
  assign n7548 = n7544 & n7547;
  assign n7549 = ~n662 & ~n1127;
  assign n7550 = ~n420 & ~n1487;
  assign n7551 = n7549 & n7550;
  assign n7552 = ~n108 & ~n894;
  assign n7553 = n4026 & n7552;
  assign n7554 = n1671 & n2577;
  assign n7555 = n7553 & n7554;
  assign n7556 = n7551 & n7555;
  assign n7557 = n1277 & n3670;
  assign n7558 = n3217 & n7557;
  assign n7559 = n54102 & n7558;
  assign n7560 = n7556 & n7559;
  assign n7561 = n7510 & n7529;
  assign n7562 = n54100 & n54102;
  assign n7563 = n3217 & n7562;
  assign n7564 = n2577 & n7563;
  assign n7565 = n3670 & n7564;
  assign n7566 = n1671 & n7565;
  assign n7567 = n4026 & n7566;
  assign n7568 = n1277 & n7567;
  assign n7569 = ~n894 & n7568;
  assign n7570 = ~n1127 & n7569;
  assign n7571 = ~n1487 & n7570;
  assign n7572 = ~n108 & n7571;
  assign n7573 = ~n662 & n7572;
  assign n7574 = ~n420 & n7573;
  assign n7575 = n54100 & n54103;
  assign n7576 = ~n404 & ~n1280;
  assign n7577 = ~n404 & n54104;
  assign n7578 = ~n1280 & n7577;
  assign n7579 = n54104 & n7576;
  assign n7580 = ~n659 & ~n1034;
  assign n7581 = ~n659 & ~n1465;
  assign n7582 = ~n1034 & n7581;
  assign n7583 = ~n1034 & ~n1465;
  assign n7584 = ~n659 & n7583;
  assign n7585 = ~n1465 & n7580;
  assign n7586 = ~n268 & ~n311;
  assign n7587 = ~n513 & ~n1457;
  assign n7588 = ~n268 & ~n1457;
  assign n7589 = ~n311 & ~n513;
  assign n7590 = n7588 & n7589;
  assign n7591 = n7586 & n7587;
  assign n7592 = n1642 & n3932;
  assign n7593 = n54107 & n7592;
  assign n7594 = n54106 & n7593;
  assign n7595 = ~n101 & ~n172;
  assign n7596 = ~n212 & ~n622;
  assign n7597 = ~n182 & n7596;
  assign n7598 = ~n212 & n7595;
  assign n7599 = ~n182 & n7598;
  assign n7600 = ~n622 & n7599;
  assign n7601 = n7595 & n7597;
  assign n7602 = ~n459 & ~n1125;
  assign n7603 = n4753 & n7602;
  assign n7604 = ~n660 & ~n1196;
  assign n7605 = n2043 & n7604;
  assign n7606 = n7603 & n7605;
  assign n7607 = n54108 & n7606;
  assign n7608 = ~n268 & ~n1196;
  assign n7609 = ~n311 & ~n1457;
  assign n7610 = ~n311 & ~n1196;
  assign n7611 = n7588 & n7610;
  assign n7612 = n7608 & n7609;
  assign n7613 = n1391 & n4753;
  assign n7614 = n54109 & n7613;
  assign n7615 = n54106 & n7614;
  assign n7616 = ~n459 & ~n2042;
  assign n7617 = ~n751 & ~n1125;
  assign n7618 = n2043 & n7602;
  assign n7619 = n7616 & n7617;
  assign n7620 = n7592 & n54110;
  assign n7621 = n54108 & n7620;
  assign n7622 = n7615 & n7621;
  assign n7623 = n54109 & n54110;
  assign n7624 = n54106 & n7623;
  assign n7625 = n1642 & n4753;
  assign n7626 = n1391 & n3932;
  assign n7627 = n7625 & n7626;
  assign n7628 = n54108 & n7627;
  assign n7629 = n7624 & n7628;
  assign n7630 = n7594 & n7607;
  assign n7631 = n3932 & n54106;
  assign n7632 = n4753 & n7631;
  assign n7633 = n54108 & n7632;
  assign n7634 = n53917 & n7633;
  assign n7635 = n1391 & n7634;
  assign n7636 = n1642 & n7635;
  assign n7637 = ~n1125 & n7636;
  assign n7638 = ~n1196 & n7637;
  assign n7639 = ~n311 & n7638;
  assign n7640 = ~n1457 & n7639;
  assign n7641 = ~n459 & n7640;
  assign n7642 = ~n268 & n7641;
  assign n7643 = ~n751 & n7642;
  assign n7644 = ~n2042 & n7643;
  assign n7645 = n53917 & n54111;
  assign n7646 = ~n361 & ~n1476;
  assign n7647 = ~n206 & ~n495;
  assign n7648 = ~n168 & ~n216;
  assign n7649 = n7647 & n7648;
  assign n7650 = n7646 & n7647;
  assign n7651 = n7648 & n7650;
  assign n7652 = n7646 & n7649;
  assign n7653 = n512 & ~n849;
  assign n7654 = n5277 & n7418;
  assign n7655 = n7653 & n7654;
  assign n7656 = n2771 & n7655;
  assign n7657 = n512 & n2771;
  assign n7658 = n5277 & n7657;
  assign n7659 = n7646 & n7658;
  assign n7660 = ~n168 & n7659;
  assign n7661 = n7418 & n7660;
  assign n7662 = ~n206 & n7661;
  assign n7663 = ~n216 & n7662;
  assign n7664 = ~n495 & n7663;
  assign n7665 = ~n849 & n7664;
  assign n7666 = n512 & n7646;
  assign n7667 = n7647 & n7666;
  assign n7668 = ~n849 & n7648;
  assign n7669 = n7654 & n7668;
  assign n7670 = n2771 & n7669;
  assign n7671 = n7667 & n7670;
  assign n7672 = n512 & n7654;
  assign n7673 = ~n216 & n7647;
  assign n7674 = ~n168 & ~n849;
  assign n7675 = n7646 & n7674;
  assign n7676 = n7673 & n7675;
  assign n7677 = n2771 & n7676;
  assign n7678 = n7672 & n7677;
  assign n7679 = n54113 & n7656;
  assign n7680 = ~n215 & ~n562;
  assign n7681 = ~n747 & ~n1681;
  assign n7682 = ~n215 & ~n747;
  assign n7683 = ~n562 & ~n1681;
  assign n7684 = n7682 & n7683;
  assign n7685 = n7680 & n7681;
  assign n7686 = n755 & n2093;
  assign n7687 = n54115 & n7686;
  assign n7688 = n586 & n712;
  assign n7689 = ~n255 & ~n651;
  assign n7690 = ~n255 & ~n416;
  assign n7691 = ~n651 & n7690;
  assign n7692 = ~n416 & n7689;
  assign n7693 = n7688 & n54116;
  assign n7694 = n7687 & n7693;
  assign n7695 = ~n222 & ~n623;
  assign n7696 = ~n163 & ~n740;
  assign n7697 = ~n948 & ~n1491;
  assign n7698 = n7696 & n7697;
  assign n7699 = ~n163 & n7697;
  assign n7700 = ~n222 & n7699;
  assign n7701 = ~n740 & n7700;
  assign n7702 = ~n623 & n7701;
  assign n7703 = ~n163 & ~n948;
  assign n7704 = ~n623 & ~n740;
  assign n7705 = ~n222 & ~n1491;
  assign n7706 = n7704 & n7705;
  assign n7707 = n7703 & n7706;
  assign n7708 = ~n623 & ~n948;
  assign n7709 = ~n163 & ~n1491;
  assign n7710 = ~n222 & ~n740;
  assign n7711 = n7709 & n7710;
  assign n7712 = n7708 & n7711;
  assign n7713 = n7695 & n7698;
  assign n7714 = n1082 & n4710;
  assign n7715 = n5639 & n7714;
  assign n7716 = n53788 & n7715;
  assign n7717 = n54117 & n7716;
  assign n7718 = n54115 & n54116;
  assign n7719 = n2093 & n4710;
  assign n7720 = n755 & n5639;
  assign n7721 = n7719 & n7720;
  assign n7722 = n7718 & n7721;
  assign n7723 = n712 & n1082;
  assign n7724 = n586 & n7723;
  assign n7725 = n53788 & n7724;
  assign n7726 = n54117 & n7725;
  assign n7727 = n7722 & n7726;
  assign n7728 = n7719 & n7723;
  assign n7729 = n7718 & n7728;
  assign n7730 = n586 & n7720;
  assign n7731 = n54117 & n7730;
  assign n7732 = n53788 & n7731;
  assign n7733 = n7729 & n7732;
  assign n7734 = n7694 & n7717;
  assign n7735 = n54114 & n54118;
  assign n7736 = n54112 & n7735;
  assign n7737 = n54105 & n54116;
  assign n7738 = n1082 & n7737;
  assign n7739 = n53788 & n7738;
  assign n7740 = n54117 & n7739;
  assign n7741 = n54112 & n7740;
  assign n7742 = n54114 & n7741;
  assign n7743 = n755 & n7742;
  assign n7744 = n586 & n7743;
  assign n7745 = n712 & n7744;
  assign n7746 = n2093 & n7745;
  assign n7747 = n4710 & n7746;
  assign n7748 = n5639 & n7747;
  assign n7749 = ~n1681 & n7748;
  assign n7750 = ~n215 & n7749;
  assign n7751 = ~n562 & n7750;
  assign n7752 = ~n747 & n7751;
  assign n7753 = n54105 & n7736;
  assign n7754 = ~n54098 & ~n54119;
  assign n7755 = ~n295 & ~n1478;
  assign n7756 = ~n250 & n1708;
  assign n7757 = n1708 & n7755;
  assign n7758 = ~n250 & n7757;
  assign n7759 = n7755 & n7756;
  assign n7760 = ~n112 & ~n247;
  assign n7761 = ~n1079 & ~n1646;
  assign n7762 = ~n112 & ~n1079;
  assign n7763 = ~n247 & n7762;
  assign n7764 = ~n1646 & n7763;
  assign n7765 = ~n112 & ~n1646;
  assign n7766 = ~n247 & ~n1079;
  assign n7767 = n7765 & n7766;
  assign n7768 = n7760 & n7761;
  assign n7769 = ~n269 & ~n664;
  assign n7770 = ~n269 & ~n771;
  assign n7771 = ~n664 & n7770;
  assign n7772 = ~n664 & ~n771;
  assign n7773 = ~n269 & n7772;
  assign n7774 = ~n771 & n7769;
  assign n7775 = ~n664 & n54121;
  assign n7776 = ~n269 & n7775;
  assign n7777 = ~n771 & n7776;
  assign n7778 = n54121 & n54122;
  assign n7779 = n3671 & n4022;
  assign n7780 = n2092 & n4022;
  assign n7781 = n3671 & n7780;
  assign n7782 = n2092 & n7779;
  assign n7783 = n54123 & n54124;
  assign n7784 = n54120 & n54124;
  assign n7785 = n54123 & n7784;
  assign n7786 = n54120 & n7783;
  assign n7787 = ~n587 & n2094;
  assign n7788 = ~n830 & ~n1658;
  assign n7789 = ~n465 & ~n896;
  assign n7790 = n7788 & n7789;
  assign n7791 = n6577 & n7788;
  assign n7792 = n7789 & n7791;
  assign n7793 = n6577 & n7790;
  assign n7794 = n2094 & n6577;
  assign n7795 = n2094 & n7791;
  assign n7796 = n7788 & n7794;
  assign n7797 = ~n896 & n54127;
  assign n7798 = ~n587 & n7797;
  assign n7799 = ~n465 & n7798;
  assign n7800 = ~n587 & n7788;
  assign n7801 = n7789 & n7794;
  assign n7802 = n7800 & n7801;
  assign n7803 = ~n587 & n7789;
  assign n7804 = n54127 & n7803;
  assign n7805 = n7787 & n54126;
  assign n7806 = ~n317 & ~n565;
  assign n7807 = ~n317 & ~n1485;
  assign n7808 = ~n565 & n7807;
  assign n7809 = ~n1485 & n7806;
  assign n7810 = n54076 & n54129;
  assign n7811 = ~n441 & ~n1125;
  assign n7812 = ~n419 & ~n562;
  assign n7813 = ~n562 & ~n1125;
  assign n7814 = ~n441 & n7813;
  assign n7815 = ~n419 & n7814;
  assign n7816 = n7811 & n7812;
  assign n7817 = ~n735 & ~n753;
  assign n7818 = ~n735 & ~n1468;
  assign n7819 = ~n753 & n7818;
  assign n7820 = ~n753 & ~n1468;
  assign n7821 = ~n735 & n7820;
  assign n7822 = ~n1468 & n7817;
  assign n7823 = n54130 & n54131;
  assign n7824 = n7810 & n7823;
  assign n7825 = n53969 & n7824;
  assign n7826 = n54128 & n7825;
  assign n7827 = n54125 & n7826;
  assign n7828 = n53921 & n53995;
  assign n7829 = n54120 & n54131;
  assign n7830 = n54076 & n7829;
  assign n7831 = n53995 & n7830;
  assign n7832 = n53969 & n7831;
  assign n7833 = n53921 & n7832;
  assign n7834 = n3671 & n7833;
  assign n7835 = n2092 & n7834;
  assign n7836 = n54130 & n7835;
  assign n7837 = n54123 & n7836;
  assign n7838 = n54128 & n7837;
  assign n7839 = ~n1485 & n7838;
  assign n7840 = ~n211 & n7839;
  assign n7841 = ~n317 & n7840;
  assign n7842 = ~n565 & n7841;
  assign n7843 = ~n361 & n7842;
  assign n7844 = n7827 & n7828;
  assign n7845 = ~n54119 & ~n54132;
  assign n7846 = ~n307 & ~n499;
  assign n7847 = ~n307 & n53733;
  assign n7848 = ~n499 & n7847;
  assign n7849 = n53733 & n7846;
  assign n7850 = ~n161 & ~n1469;
  assign n7851 = ~n268 & n4094;
  assign n7852 = ~n1469 & n4094;
  assign n7853 = ~n161 & n7852;
  assign n7854 = ~n268 & n7853;
  assign n7855 = ~n268 & n7850;
  assign n7856 = n4094 & n7855;
  assign n7857 = n7850 & n7851;
  assign n7858 = ~n461 & ~n1491;
  assign n7859 = n106 & n7858;
  assign n7860 = n3933 & n5378;
  assign n7861 = n6535 & n6860;
  assign n7862 = n7860 & n7861;
  assign n7863 = ~n101 & ~n1491;
  assign n7864 = n3933 & n7863;
  assign n7865 = ~n105 & ~n461;
  assign n7866 = n6535 & n7865;
  assign n7867 = n5378 & n6860;
  assign n7868 = n7866 & n7867;
  assign n7869 = n7864 & n7868;
  assign n7870 = ~n101 & ~n461;
  assign n7871 = n3933 & n7870;
  assign n7872 = ~n105 & ~n1491;
  assign n7873 = n5378 & n7872;
  assign n7874 = n7861 & n7873;
  assign n7875 = n7871 & n7874;
  assign n7876 = n7859 & n7862;
  assign n7877 = n6860 & n54134;
  assign n7878 = n5378 & n7877;
  assign n7879 = n6535 & n7878;
  assign n7880 = ~n1491 & n7879;
  assign n7881 = ~n101 & n7880;
  assign n7882 = ~n105 & n7881;
  assign n7883 = ~n461 & n7882;
  assign n7884 = ~n360 & n7883;
  assign n7885 = ~n774 & n7884;
  assign n7886 = n54134 & n54135;
  assign n7887 = ~n247 & ~n552;
  assign n7888 = ~n247 & ~n1124;
  assign n7889 = ~n552 & n7888;
  assign n7890 = ~n552 & ~n1124;
  assign n7891 = ~n247 & n7890;
  assign n7892 = ~n1124 & n7887;
  assign n7893 = ~n321 & ~n340;
  assign n7894 = ~n321 & ~n440;
  assign n7895 = ~n340 & n7894;
  assign n7896 = ~n340 & ~n440;
  assign n7897 = ~n321 & n7896;
  assign n7898 = ~n440 & n7893;
  assign n7899 = n53720 & n54138;
  assign n7900 = n53720 & n54137;
  assign n7901 = n54138 & n7900;
  assign n7902 = n54137 & n7899;
  assign n7903 = ~n510 & ~n829;
  assign n7904 = ~n294 & ~n1644;
  assign n7905 = n5485 & n7904;
  assign n7906 = n7903 & n7905;
  assign n7907 = ~n269 & ~n448;
  assign n7908 = ~n450 & ~n2109;
  assign n7909 = ~n269 & ~n2109;
  assign n7910 = ~n448 & ~n450;
  assign n7911 = n7909 & n7910;
  assign n7912 = n7907 & n7908;
  assign n7913 = n276 & n5652;
  assign n7914 = n54140 & n7913;
  assign n7915 = n5652 & n7904;
  assign n7916 = n7903 & n7915;
  assign n7917 = n276 & n5485;
  assign n7918 = n54140 & n7917;
  assign n7919 = n7916 & n7918;
  assign n7920 = n5652 & n7917;
  assign n7921 = n5485 & n7913;
  assign n7922 = ~n829 & ~n1644;
  assign n7923 = n7909 & n7922;
  assign n7924 = ~n294 & ~n450;
  assign n7925 = ~n448 & ~n510;
  assign n7926 = n7924 & n7925;
  assign n7927 = ~n269 & ~n829;
  assign n7928 = n7904 & n7927;
  assign n7929 = ~n448 & ~n2109;
  assign n7930 = ~n450 & ~n510;
  assign n7931 = n7929 & n7930;
  assign n7932 = n7928 & n7931;
  assign n7933 = n7923 & n7926;
  assign n7934 = n54142 & n54143;
  assign n7935 = n7906 & n7914;
  assign n7936 = n54139 & n54141;
  assign n7937 = n5485 & n54138;
  assign n7938 = n54137 & n7937;
  assign n7939 = n54136 & n7938;
  assign n7940 = n53720 & n7939;
  assign n7941 = n5652 & n7940;
  assign n7942 = n276 & n7941;
  assign n7943 = ~n294 & n7942;
  assign n7944 = ~n829 & n7943;
  assign n7945 = ~n269 & n7944;
  assign n7946 = ~n1644 & n7945;
  assign n7947 = ~n510 & n7946;
  assign n7948 = ~n450 & n7947;
  assign n7949 = ~n448 & n7948;
  assign n7950 = ~n2109 & n7949;
  assign n7951 = n54136 & n7936;
  assign n7952 = ~n553 & ~n646;
  assign n7953 = n347 & n7952;
  assign n7954 = n5277 & n7953;
  assign n7955 = n1067 & n4585;
  assign n7956 = ~n255 & ~n750;
  assign n7957 = ~n902 & n7956;
  assign n7958 = n53734 & n7957;
  assign n7959 = n7955 & n7958;
  assign n7960 = n347 & n53734;
  assign n7961 = n4585 & n7960;
  assign n7962 = n1067 & n7961;
  assign n7963 = n5277 & n7962;
  assign n7964 = ~n902 & n7963;
  assign n7965 = ~n255 & n7964;
  assign n7966 = ~n553 & n7965;
  assign n7967 = ~n646 & n7966;
  assign n7968 = ~n750 & n7967;
  assign n7969 = ~n255 & ~n646;
  assign n7970 = n347 & n7969;
  assign n7971 = n5277 & n7970;
  assign n7972 = ~n553 & ~n750;
  assign n7973 = ~n902 & n7972;
  assign n7974 = n53734 & n7973;
  assign n7975 = n7955 & n7974;
  assign n7976 = n7971 & n7975;
  assign n7977 = ~n646 & ~n750;
  assign n7978 = n347 & n7977;
  assign n7979 = n5277 & n7978;
  assign n7980 = ~n255 & ~n553;
  assign n7981 = ~n255 & ~n902;
  assign n7982 = ~n553 & n7981;
  assign n7983 = ~n902 & n7980;
  assign n7984 = n53734 & n54146;
  assign n7985 = n7955 & n7984;
  assign n7986 = n7979 & n7985;
  assign n7987 = n347 & n7955;
  assign n7988 = n5277 & n7977;
  assign n7989 = n54146 & n7988;
  assign n7990 = n53734 & n7989;
  assign n7991 = n7987 & n7990;
  assign n7992 = n7954 & n7959;
  assign n7993 = ~n1127 & ~n1997;
  assign n7994 = ~n881 & ~n1997;
  assign n7995 = ~n1127 & n7994;
  assign n7996 = ~n881 & n7993;
  assign n7997 = ~n112 & ~n363;
  assign n7998 = ~n401 & ~n617;
  assign n7999 = ~n451 & ~n1455;
  assign n8000 = ~n451 & ~n617;
  assign n8001 = ~n401 & ~n1455;
  assign n8002 = n8000 & n8001;
  assign n8003 = n7998 & n7999;
  assign n8004 = n7997 & n54148;
  assign n8005 = ~n112 & n54147;
  assign n8006 = ~n401 & n8005;
  assign n8007 = ~n1455 & n8006;
  assign n8008 = ~n617 & n8007;
  assign n8009 = ~n363 & n8008;
  assign n8010 = ~n451 & n8009;
  assign n8011 = ~n112 & ~n1455;
  assign n8012 = ~n1127 & n8011;
  assign n8013 = ~n617 & ~n1997;
  assign n8014 = ~n401 & ~n881;
  assign n8015 = ~n363 & ~n451;
  assign n8016 = n8014 & n8015;
  assign n8017 = n8013 & n8016;
  assign n8018 = n8012 & n8017;
  assign n8019 = n54147 & n8004;
  assign n8020 = n1391 & n3086;
  assign n8021 = n3475 & n4472;
  assign n8022 = n8020 & n8021;
  assign n8023 = ~n1337 & ~n1457;
  assign n8024 = ~n1486 & ~n1881;
  assign n8025 = n8023 & n8024;
  assign n8026 = ~n554 & ~n753;
  assign n8027 = n217 & n8026;
  assign n8028 = n8025 & n8027;
  assign n8029 = ~n1457 & ~n1478;
  assign n8030 = ~n554 & ~n1486;
  assign n8031 = n8029 & n8030;
  assign n8032 = ~n753 & ~n848;
  assign n8033 = ~n1337 & ~n1881;
  assign n8034 = n8032 & n8033;
  assign n8035 = ~n1457 & ~n1486;
  assign n8036 = n4472 & n8035;
  assign n8037 = ~n753 & ~n1337;
  assign n8038 = ~n554 & ~n1881;
  assign n8039 = n8037 & n8038;
  assign n8040 = n8036 & n8039;
  assign n8041 = n8031 & n8034;
  assign n8042 = n217 & n3475;
  assign n8043 = n8020 & n8042;
  assign n8044 = n54150 & n8043;
  assign n8045 = n8022 & n8028;
  assign n8046 = n175 & ~n741;
  assign n8047 = n175 & n3742;
  assign n8048 = ~n741 & n8047;
  assign n8049 = ~n741 & n3742;
  assign n8050 = n175 & n8049;
  assign n8051 = n3742 & n8046;
  assign n8052 = ~n466 & ~n1061;
  assign n8053 = n4799 & n5362;
  assign n8054 = n8052 & n8053;
  assign n8055 = n54152 & n8054;
  assign n8056 = n1391 & n4799;
  assign n8057 = n3475 & n5362;
  assign n8058 = n8056 & n8057;
  assign n8059 = n54150 & n8058;
  assign n8060 = n217 & n8052;
  assign n8061 = n3086 & n8060;
  assign n8062 = n54152 & n8061;
  assign n8063 = n8059 & n8062;
  assign n8064 = n54151 & n8055;
  assign n8065 = n54149 & n54153;
  assign n8066 = n54145 & n8065;
  assign n8067 = n54144 & n8066;
  assign n8068 = n54133 & n54152;
  assign n8069 = n4799 & n8068;
  assign n8070 = n5362 & n8069;
  assign n8071 = n54145 & n8070;
  assign n8072 = n54144 & n8071;
  assign n8073 = n54149 & n8072;
  assign n8074 = n3086 & n8073;
  assign n8075 = n217 & n8074;
  assign n8076 = n8052 & n8075;
  assign n8077 = n1391 & n8076;
  assign n8078 = n3475 & n8077;
  assign n8079 = ~n1486 & n8078;
  assign n8080 = ~n1478 & n8079;
  assign n8081 = ~n554 & n8080;
  assign n8082 = ~n1457 & n8081;
  assign n8083 = ~n1337 & n8082;
  assign n8084 = ~n848 & n8083;
  assign n8085 = ~n753 & n8084;
  assign n8086 = ~n1881 & n8085;
  assign n8087 = n54133 & n8067;
  assign n8088 = ~n54132 & ~n54154;
  assign n8089 = ~n348 & ~n623;
  assign n8090 = n5198 & n8089;
  assign n8091 = ~n401 & ~n1485;
  assign n8092 = ~n776 & ~n975;
  assign n8093 = n8091 & n8092;
  assign n8094 = n5198 & n8091;
  assign n8095 = n8089 & n8092;
  assign n8096 = n8094 & n8095;
  assign n8097 = n8090 & n8093;
  assign n8098 = ~n591 & ~n883;
  assign n8099 = ~n883 & ~n1472;
  assign n8100 = ~n591 & n8099;
  assign n8101 = ~n591 & ~n1472;
  assign n8102 = ~n883 & n8101;
  assign n8103 = ~n1472 & n8098;
  assign n8104 = ~n174 & ~n822;
  assign n8105 = n4383 & n8104;
  assign n8106 = n54131 & n8105;
  assign n8107 = n54156 & n8106;
  assign n8108 = n54131 & n54156;
  assign n8109 = n5198 & n8108;
  assign n8110 = n4383 & n8109;
  assign n8111 = n8091 & n8110;
  assign n8112 = ~n174 & n8111;
  assign n8113 = ~n822 & n8112;
  assign n8114 = ~n975 & n8113;
  assign n8115 = ~n348 & n8114;
  assign n8116 = ~n776 & n8115;
  assign n8117 = ~n623 & n8116;
  assign n8118 = n4383 & n5198;
  assign n8119 = n8093 & n8118;
  assign n8120 = n8089 & n8104;
  assign n8121 = n54131 & n8120;
  assign n8122 = n54156 & n8121;
  assign n8123 = n8119 & n8122;
  assign n8124 = ~n174 & ~n623;
  assign n8125 = n8091 & n8124;
  assign n8126 = n8118 & n8125;
  assign n8127 = ~n348 & ~n822;
  assign n8128 = n8092 & n8127;
  assign n8129 = n54131 & n8128;
  assign n8130 = n54156 & n8129;
  assign n8131 = n8126 & n8130;
  assign n8132 = n54155 & n8107;
  assign n8133 = ~n246 & ~n848;
  assign n8134 = ~n1486 & n8133;
  assign n8135 = n5024 & n8134;
  assign n8136 = n53620 & n8135;
  assign n8137 = n1067 & n1820;
  assign n8138 = ~n564 & ~n1912;
  assign n8139 = n7595 & n8138;
  assign n8140 = n8137 & n8139;
  assign n8141 = n53738 & n8140;
  assign n8142 = ~n268 & n2326;
  assign n8143 = n2326 & n4224;
  assign n8144 = ~n268 & n8143;
  assign n8145 = ~n268 & n4224;
  assign n8146 = n2326 & n8145;
  assign n8147 = n4224 & n8142;
  assign n8148 = ~n319 & n629;
  assign n8149 = n343 & n831;
  assign n8150 = n629 & n831;
  assign n8151 = n343 & n8150;
  assign n8152 = ~n319 & n8151;
  assign n8153 = ~n319 & n343;
  assign n8154 = n8150 & n8153;
  assign n8155 = n8148 & n8149;
  assign n8156 = n54158 & n54159;
  assign n8157 = n8141 & n8156;
  assign n8158 = ~n246 & ~n983;
  assign n8159 = ~n357 & ~n848;
  assign n8160 = n8158 & n8159;
  assign n8161 = ~n163 & ~n1486;
  assign n8162 = n749 & n8161;
  assign n8163 = n8160 & n8162;
  assign n8164 = n53620 & n8163;
  assign n8165 = n1067 & n7595;
  assign n8166 = n8138 & n8165;
  assign n8167 = n53738 & n8166;
  assign n8168 = n8156 & n8167;
  assign n8169 = n8164 & n8168;
  assign n8170 = ~n163 & ~n246;
  assign n8171 = ~n983 & ~n1486;
  assign n8172 = n8170 & n8171;
  assign n8173 = ~n848 & ~n1912;
  assign n8174 = ~n357 & ~n564;
  assign n8175 = n8173 & n8174;
  assign n8176 = n8172 & n8175;
  assign n8177 = n53620 & n8176;
  assign n8178 = n749 & n1067;
  assign n8179 = n7595 & n8178;
  assign n8180 = n53738 & n8179;
  assign n8181 = n8156 & n8180;
  assign n8182 = n8177 & n8181;
  assign n8183 = n8136 & n8157;
  assign n8184 = n54157 & n54160;
  assign n8185 = ~n1085 & ~n1641;
  assign n8186 = ~n356 & ~n402;
  assign n8187 = ~n402 & ~n1085;
  assign n8188 = ~n1641 & n8187;
  assign n8189 = ~n356 & n8188;
  assign n8190 = n8185 & n8186;
  assign n8191 = ~n444 & ~n659;
  assign n8192 = ~n1535 & n8191;
  assign n8193 = n53836 & n8192;
  assign n8194 = n54161 & n8193;
  assign n8195 = n3214 & n6309;
  assign n8196 = ~n1034 & ~n2109;
  assign n8197 = n7201 & n8196;
  assign n8198 = n8195 & n8197;
  assign n8199 = n1361 & n3639;
  assign n8200 = n3535 & n4083;
  assign n8201 = n8199 & n8200;
  assign n8202 = n8198 & n8201;
  assign n8203 = n54078 & n8202;
  assign n8204 = n6309 & n8196;
  assign n8205 = n53836 & n8204;
  assign n8206 = n54161 & n8205;
  assign n8207 = n54078 & n8206;
  assign n8208 = n3639 & n8207;
  assign n8209 = n3535 & n8208;
  assign n8210 = n3214 & n8209;
  assign n8211 = n7201 & n8210;
  assign n8212 = n4083 & n8211;
  assign n8213 = ~n659 & n8212;
  assign n8214 = ~n1535 & n8213;
  assign n8215 = ~n611 & n8214;
  assign n8216 = ~n444 & n8215;
  assign n8217 = ~n789 & n8216;
  assign n8218 = ~n659 & ~n789;
  assign n8219 = ~n611 & n8218;
  assign n8220 = n53836 & n8219;
  assign n8221 = n54161 & n8220;
  assign n8222 = n4083 & n6309;
  assign n8223 = n8197 & n8222;
  assign n8224 = ~n444 & ~n1535;
  assign n8225 = n3214 & n8224;
  assign n8226 = n3535 & n3639;
  assign n8227 = n8225 & n8226;
  assign n8228 = n8223 & n8227;
  assign n8229 = n54078 & n8228;
  assign n8230 = n8221 & n8229;
  assign n8231 = ~n789 & ~n1535;
  assign n8232 = ~n444 & n8231;
  assign n8233 = n53836 & n8232;
  assign n8234 = n54161 & n8233;
  assign n8235 = n3535 & n7201;
  assign n8236 = n3639 & n8196;
  assign n8237 = n8235 & n8236;
  assign n8238 = ~n611 & ~n659;
  assign n8239 = n4083 & n8238;
  assign n8240 = n8195 & n8239;
  assign n8241 = n8237 & n8240;
  assign n8242 = n54078 & n8241;
  assign n8243 = n8234 & n8242;
  assign n8244 = n8194 & n8203;
  assign n8245 = n54058 & n54162;
  assign n8246 = n53620 & n54162;
  assign n8247 = n54159 & n8246;
  assign n8248 = n54058 & n8247;
  assign n8249 = n54158 & n8248;
  assign n8250 = n1067 & n8249;
  assign n8251 = n53738 & n8250;
  assign n8252 = n54157 & n8251;
  assign n8253 = n749 & n8252;
  assign n8254 = ~n1486 & n8253;
  assign n8255 = ~n983 & n8254;
  assign n8256 = ~n163 & n8255;
  assign n8257 = n7595 & n8256;
  assign n8258 = ~n246 & n8257;
  assign n8259 = ~n564 & n8258;
  assign n8260 = ~n848 & n8259;
  assign n8261 = ~n357 & n8260;
  assign n8262 = ~n1912 & n8261;
  assign n8263 = n8184 & n8245;
  assign n8264 = ~n54154 & ~n54163;
  assign n8265 = ~n268 & ~n646;
  assign n8266 = n6198 & n8265;
  assign n8267 = ~n212 & ~n587;
  assign n8268 = ~n168 & ~n1234;
  assign n8269 = n8267 & n8268;
  assign n8270 = n6198 & n8268;
  assign n8271 = n8265 & n8267;
  assign n8272 = n8270 & n8271;
  assign n8273 = n8266 & n8269;
  assign n8274 = ~n1085 & n5874;
  assign n8275 = ~n491 & ~n748;
  assign n8276 = ~n491 & ~n1492;
  assign n8277 = ~n748 & n8276;
  assign n8278 = ~n1492 & n8275;
  assign n8279 = n3715 & n3878;
  assign n8280 = n54165 & n8279;
  assign n8281 = n8274 & n8280;
  assign n8282 = n3878 & n8268;
  assign n8283 = n3715 & n8267;
  assign n8284 = n3715 & n8269;
  assign n8285 = n3878 & n8284;
  assign n8286 = n8282 & n8283;
  assign n8287 = n8274 & n54166;
  assign n8288 = ~n1127 & n8287;
  assign n8289 = ~n1492 & n8288;
  assign n8290 = ~n247 & n8289;
  assign n8291 = ~n748 & n8290;
  assign n8292 = ~n268 & n8291;
  assign n8293 = ~n491 & n8292;
  assign n8294 = ~n646 & n8293;
  assign n8295 = ~n1492 & n6198;
  assign n8296 = n8265 & n8275;
  assign n8297 = n8295 & n8296;
  assign n8298 = n8274 & n8297;
  assign n8299 = n54166 & n8298;
  assign n8300 = n54164 & n8281;
  assign n8301 = ~n405 & ~n408;
  assign n8302 = ~n789 & ~n1195;
  assign n8303 = n8301 & n8302;
  assign n8304 = n629 & n7245;
  assign n8305 = n185 & n2340;
  assign n8306 = n8304 & n8305;
  assign n8307 = n8303 & n8306;
  assign n8308 = ~n423 & ~n1646;
  assign n8309 = ~n216 & ~n883;
  assign n8310 = n963 & n8309;
  assign n8311 = ~n1646 & n8309;
  assign n8312 = ~n443 & n8311;
  assign n8313 = ~n423 & n8312;
  assign n8314 = ~n615 & n8313;
  assign n8315 = n8308 & n8309;
  assign n8316 = n963 & n8315;
  assign n8317 = n8308 & n8310;
  assign n8318 = n4261 & n4529;
  assign n8319 = ~n440 & ~n585;
  assign n8320 = ~n161 & ~n271;
  assign n8321 = n8319 & n8320;
  assign n8322 = n8318 & n8321;
  assign n8323 = n53984 & n8322;
  assign n8324 = n54168 & n8323;
  assign n8325 = ~n258 & ~n440;
  assign n8326 = ~n585 & ~n789;
  assign n8327 = n8325 & n8326;
  assign n8328 = n2340 & n4261;
  assign n8329 = ~n405 & ~n1195;
  assign n8330 = ~n275 & ~n408;
  assign n8331 = n8329 & n8330;
  assign n8332 = n8328 & n8331;
  assign n8333 = n8327 & n8332;
  assign n8334 = n629 & n4529;
  assign n8335 = n185 & n8320;
  assign n8336 = n8334 & n8335;
  assign n8337 = n54168 & n8336;
  assign n8338 = n53984 & n8337;
  assign n8339 = n8333 & n8338;
  assign n8340 = ~n585 & ~n1195;
  assign n8341 = ~n275 & ~n440;
  assign n8342 = n8340 & n8341;
  assign n8343 = ~n161 & ~n408;
  assign n8344 = ~n405 & ~n789;
  assign n8345 = n8343 & n8344;
  assign n8346 = ~n258 & ~n271;
  assign n8347 = n4261 & n8346;
  assign n8348 = n8345 & n8347;
  assign n8349 = n8342 & n8348;
  assign n8350 = n2340 & n4529;
  assign n8351 = n185 & n629;
  assign n8352 = n8350 & n8351;
  assign n8353 = n53984 & n8352;
  assign n8354 = n54168 & n8353;
  assign n8355 = n8349 & n8354;
  assign n8356 = n8307 & n8324;
  assign n8357 = n54167 & n54169;
  assign n8358 = ~n207 & ~n881;
  assign n8359 = ~n881 & n5873;
  assign n8360 = ~n207 & n8359;
  assign n8361 = n5873 & n8358;
  assign n8362 = ~n211 & n3737;
  assign n8363 = n54071 & n8362;
  assign n8364 = n54170 & n8363;
  assign n8365 = ~n416 & ~n911;
  assign n8366 = ~n1469 & ~n1477;
  assign n8367 = n8365 & n8366;
  assign n8368 = ~n460 & ~n1490;
  assign n8369 = ~n179 & ~n295;
  assign n8370 = n8368 & n8369;
  assign n8371 = ~n295 & ~n416;
  assign n8372 = ~n1469 & n8371;
  assign n8373 = ~n1490 & n8372;
  assign n8374 = ~n1477 & n8373;
  assign n8375 = ~n179 & n8374;
  assign n8376 = ~n911 & n8375;
  assign n8377 = ~n460 & n8376;
  assign n8378 = ~n295 & ~n1469;
  assign n8379 = n8365 & n8378;
  assign n8380 = ~n179 & ~n1477;
  assign n8381 = n8368 & n8380;
  assign n8382 = n8379 & n8381;
  assign n8383 = ~n911 & ~n1490;
  assign n8384 = ~n179 & ~n460;
  assign n8385 = n8383 & n8384;
  assign n8386 = n8366 & n8371;
  assign n8387 = n8385 & n8386;
  assign n8388 = n8367 & n8370;
  assign n8389 = ~n163 & ~n562;
  assign n8390 = n5943 & n7788;
  assign n8391 = n8389 & n8390;
  assign n8392 = n3535 & n3607;
  assign n8393 = n4258 & n5538;
  assign n8394 = n8392 & n8393;
  assign n8395 = n8391 & n8394;
  assign n8396 = n54171 & n8395;
  assign n8397 = n3607 & n54170;
  assign n8398 = n54071 & n8397;
  assign n8399 = n7788 & n8398;
  assign n8400 = n5538 & n8399;
  assign n8401 = n54171 & n8400;
  assign n8402 = n3535 & n8401;
  assign n8403 = n5943 & n8402;
  assign n8404 = n4258 & n8403;
  assign n8405 = ~n163 & n8404;
  assign n8406 = n3737 & n8405;
  assign n8407 = ~n211 & n8406;
  assign n8408 = ~n562 & n8407;
  assign n8409 = ~n211 & ~n562;
  assign n8410 = ~n211 & n8389;
  assign n8411 = ~n163 & n8409;
  assign n8412 = n54071 & n54173;
  assign n8413 = n54170 & n8412;
  assign n8414 = n3535 & n3737;
  assign n8415 = n3607 & n8414;
  assign n8416 = n8390 & n8393;
  assign n8417 = n5943 & n8393;
  assign n8418 = n3737 & n7788;
  assign n8419 = n8392 & n8418;
  assign n8420 = n8417 & n8419;
  assign n8421 = n8415 & n8416;
  assign n8422 = n54171 & n54174;
  assign n8423 = n8413 & n8422;
  assign n8424 = n8364 & n8396;
  assign n8425 = n175 & ~n901;
  assign n8426 = n905 & n6564;
  assign n8427 = n175 & n905;
  assign n8428 = ~n1191 & n8427;
  assign n8429 = ~n901 & n8428;
  assign n8430 = ~n776 & n8429;
  assign n8431 = ~n776 & ~n901;
  assign n8432 = ~n1191 & n8431;
  assign n8433 = n8427 & n8432;
  assign n8434 = n8425 & n8426;
  assign n8435 = n3369 & n5058;
  assign n8436 = n472 & n8435;
  assign n8437 = ~n259 & ~n317;
  assign n8438 = ~n852 & ~n2103;
  assign n8439 = ~n259 & ~n852;
  assign n8440 = ~n317 & ~n2103;
  assign n8441 = n8439 & n8440;
  assign n8442 = n8437 & n8438;
  assign n8443 = n1391 & n2981;
  assign n8444 = n54176 & n8443;
  assign n8445 = n472 & n5058;
  assign n8446 = n2981 & n8445;
  assign n8447 = n1391 & n3369;
  assign n8448 = n54176 & n8447;
  assign n8449 = n8446 & n8448;
  assign n8450 = n8436 & n8444;
  assign n8451 = n54175 & n54177;
  assign n8452 = ~n112 & ~n1192;
  assign n8453 = ~n1090 & ~n1681;
  assign n8454 = n5332 & n8453;
  assign n8455 = n8452 & n8454;
  assign n8456 = ~n441 & ~n504;
  assign n8457 = ~n1189 & n8456;
  assign n8458 = ~n614 & ~n663;
  assign n8459 = n4974 & n8458;
  assign n8460 = ~n1189 & n8458;
  assign n8461 = n4974 & n8456;
  assign n8462 = n8460 & n8461;
  assign n8463 = n8457 & n8459;
  assign n8464 = n2058 & n4974;
  assign n8465 = n4974 & n8453;
  assign n8466 = n2058 & n8465;
  assign n8467 = n8453 & n8464;
  assign n8468 = ~n1192 & n54179;
  assign n8469 = ~n112 & n8468;
  assign n8470 = ~n1189 & n8469;
  assign n8471 = ~n504 & n8470;
  assign n8472 = ~n441 & n8471;
  assign n8473 = ~n614 & n8472;
  assign n8474 = ~n1715 & n8473;
  assign n8475 = n2058 & n8452;
  assign n8476 = n8453 & n8475;
  assign n8477 = ~n504 & ~n614;
  assign n8478 = ~n1189 & n8477;
  assign n8479 = ~n441 & ~n1715;
  assign n8480 = n4974 & n8479;
  assign n8481 = n8478 & n8480;
  assign n8482 = n8476 & n8481;
  assign n8483 = ~n1189 & n8452;
  assign n8484 = ~n614 & ~n1715;
  assign n8485 = n8456 & n8484;
  assign n8486 = n8483 & n8485;
  assign n8487 = n54179 & n8486;
  assign n8488 = n8455 & n54178;
  assign n8489 = ~n141 & ~n340;
  assign n8490 = ~n141 & n293;
  assign n8491 = ~n340 & n8490;
  assign n8492 = n293 & n8489;
  assign n8493 = n2771 & n53896;
  assign n8494 = n54181 & n8493;
  assign n8495 = n54180 & n8494;
  assign n8496 = n2771 & n54181;
  assign n8497 = n5058 & n8496;
  assign n8498 = n2981 & n8497;
  assign n8499 = n3369 & n8498;
  assign n8500 = n472 & n8499;
  assign n8501 = n53896 & n8500;
  assign n8502 = n54175 & n8501;
  assign n8503 = n54180 & n8502;
  assign n8504 = n1391 & n8503;
  assign n8505 = ~n2103 & n8504;
  assign n8506 = ~n317 & n8505;
  assign n8507 = ~n259 & n8506;
  assign n8508 = ~n852 & n8507;
  assign n8509 = n8451 & n8495;
  assign n8510 = n54172 & n54182;
  assign n8511 = n185 & n8334;
  assign n8512 = n54168 & n8511;
  assign n8513 = n54172 & n8512;
  assign n8514 = n54167 & n8513;
  assign n8515 = n53984 & n8514;
  assign n8516 = n4261 & n8515;
  assign n8517 = n54182 & n8516;
  assign n8518 = n2340 & n8517;
  assign n8519 = ~n408 & n8518;
  assign n8520 = ~n1195 & n8519;
  assign n8521 = ~n258 & n8520;
  assign n8522 = ~n271 & n8521;
  assign n8523 = ~n161 & n8522;
  assign n8524 = ~n405 & n8523;
  assign n8525 = ~n275 & n8524;
  assign n8526 = ~n440 & n8525;
  assign n8527 = ~n789 & n8526;
  assign n8528 = ~n585 & n8527;
  assign n8529 = n8357 & n8510;
  assign n8530 = ~n54163 & ~n54183;
  assign n8531 = n304 & ~n881;
  assign n8532 = n293 & n2172;
  assign n8533 = ~n271 & ~n415;
  assign n8534 = ~n415 & ~n1634;
  assign n8535 = ~n271 & n8534;
  assign n8536 = ~n1634 & n8533;
  assign n8537 = n6615 & n54185;
  assign n8538 = n54184 & n8537;
  assign n8539 = ~n1033 & ~n1487;
  assign n8540 = n1075 & n1670;
  assign n8541 = n1670 & n8539;
  assign n8542 = n1075 & n8541;
  assign n8543 = n8539 & n8540;
  assign n8544 = n53989 & n54186;
  assign n8545 = n54123 & n8544;
  assign n8546 = n2172 & n53989;
  assign n8547 = n54123 & n8546;
  assign n8548 = n6614 & n8547;
  assign n8549 = n5873 & n8548;
  assign n8550 = n293 & n8549;
  assign n8551 = n1670 & n8550;
  assign n8552 = ~n1033 & n8551;
  assign n8553 = ~n415 & n8552;
  assign n8554 = ~n1487 & n8553;
  assign n8555 = ~n271 & n8554;
  assign n8556 = ~n660 & n8555;
  assign n8557 = ~n1634 & n8556;
  assign n8558 = ~n740 & n8557;
  assign n8559 = n8537 & n54186;
  assign n8560 = n53989 & n54184;
  assign n8561 = n54123 & n8560;
  assign n8562 = n8559 & n8561;
  assign n8563 = n1075 & ~n1487;
  assign n8564 = ~n271 & ~n1634;
  assign n8565 = ~n415 & ~n1033;
  assign n8566 = n8564 & n8565;
  assign n8567 = n1670 & n5873;
  assign n8568 = n8566 & n8567;
  assign n8569 = n8563 & n8568;
  assign n8570 = n293 & n6614;
  assign n8571 = n2172 & n8570;
  assign n8572 = n53989 & n8571;
  assign n8573 = n54123 & n8572;
  assign n8574 = n8569 & n8573;
  assign n8575 = n8538 & n8545;
  assign n8576 = ~n559 & n3389;
  assign n8577 = n3389 & n54130;
  assign n8578 = ~n559 & n8577;
  assign n8579 = n54130 & n8576;
  assign n8580 = n403 & n2693;
  assign n8581 = n403 & n1091;
  assign n8582 = n2693 & n8581;
  assign n8583 = n1091 & n8580;
  assign n8584 = ~n206 & n494;
  assign n8585 = n494 & n2340;
  assign n8586 = ~n206 & n8585;
  assign n8587 = ~n206 & n2340;
  assign n8588 = n494 & n8587;
  assign n8589 = n2340 & n8584;
  assign n8590 = n54189 & n54190;
  assign n8591 = n54188 & n54189;
  assign n8592 = n54190 & n8591;
  assign n8593 = n54188 & n54190;
  assign n8594 = n54189 & n8593;
  assign n8595 = n54188 & n8590;
  assign n8596 = n2094 & n4530;
  assign n8597 = n7201 & n8596;
  assign n8598 = ~n101 & ~n646;
  assign n8599 = ~n646 & ~n1280;
  assign n8600 = ~n101 & n8599;
  assign n8601 = ~n101 & ~n1280;
  assign n8602 = ~n646 & n8601;
  assign n8603 = ~n1280 & n8598;
  assign n8604 = ~n833 & ~n1997;
  assign n8605 = n4070 & n8604;
  assign n8606 = n54192 & n8605;
  assign n8607 = n2094 & n4070;
  assign n8608 = n7201 & n8607;
  assign n8609 = n4530 & n8604;
  assign n8610 = n54192 & n8609;
  assign n8611 = n8608 & n8610;
  assign n8612 = n8597 & n8606;
  assign n8613 = n53851 & n53863;
  assign n8614 = n54193 & n8613;
  assign n8615 = n54191 & n8614;
  assign n8616 = n54187 & n8615;
  assign n8617 = n54016 & n54189;
  assign n8618 = n54188 & n8617;
  assign n8619 = n54190 & n8618;
  assign n8620 = n53863 & n8619;
  assign n8621 = n53851 & n8620;
  assign n8622 = n54192 & n8621;
  assign n8623 = n7201 & n8622;
  assign n8624 = n4530 & n8623;
  assign n8625 = n54187 & n8624;
  assign n8626 = n2094 & n8625;
  assign n8627 = n4070 & n8626;
  assign n8628 = ~n1997 & n8627;
  assign n8629 = ~n833 & n8628;
  assign n8630 = n54016 & n8616;
  assign n8631 = ~n54183 & ~n54194;
  assign n8632 = ~n956 & ~n1487;
  assign n8633 = n3522 & n8632;
  assign n8634 = n4884 & n7308;
  assign n8635 = ~n255 & ~n1062;
  assign n8636 = n8267 & n8635;
  assign n8637 = n8634 & n8636;
  assign n8638 = ~n207 & ~n255;
  assign n8639 = n8632 & n8638;
  assign n8640 = ~n1062 & ~n1646;
  assign n8641 = n4884 & n8640;
  assign n8642 = n3522 & n8267;
  assign n8643 = n8641 & n8642;
  assign n8644 = n8639 & n8643;
  assign n8645 = n8633 & n8637;
  assign n8646 = n3522 & n4884;
  assign n8647 = n8267 & n8646;
  assign n8648 = n53954 & n8647;
  assign n8649 = ~n1062 & n8648;
  assign n8650 = ~n1487 & n8649;
  assign n8651 = ~n255 & n8650;
  assign n8652 = ~n207 & n8651;
  assign n8653 = ~n956 & n8652;
  assign n8654 = ~n1646 & n8653;
  assign n8655 = n53954 & n54195;
  assign n8656 = ~n311 & ~n1476;
  assign n8657 = n4020 & n4972;
  assign n8658 = n8656 & n8657;
  assign n8659 = ~n296 & n1577;
  assign n8660 = n54137 & n8659;
  assign n8661 = n1577 & n4020;
  assign n8662 = n54137 & n8661;
  assign n8663 = ~n296 & n8662;
  assign n8664 = ~n1476 & n8663;
  assign n8665 = ~n311 & n8664;
  assign n8666 = ~n319 & n8665;
  assign n8667 = ~n503 & n8666;
  assign n8668 = n8656 & n8661;
  assign n8669 = ~n296 & ~n503;
  assign n8670 = ~n319 & n8669;
  assign n8671 = n54137 & n8670;
  assign n8672 = n8668 & n8671;
  assign n8673 = n1577 & n8657;
  assign n8674 = ~n296 & n8656;
  assign n8675 = n54137 & n8674;
  assign n8676 = n8673 & n8675;
  assign n8677 = n8658 & n8660;
  assign n8678 = n53877 & n54094;
  assign n8679 = ~n166 & ~n618;
  assign n8680 = n164 & n8679;
  assign n8681 = ~n172 & ~n316;
  assign n8682 = ~n511 & ~n1337;
  assign n8683 = ~n1337 & n8681;
  assign n8684 = ~n511 & n8683;
  assign n8685 = ~n316 & ~n1337;
  assign n8686 = ~n172 & ~n511;
  assign n8687 = n8685 & n8686;
  assign n8688 = ~n172 & ~n1337;
  assign n8689 = ~n316 & ~n511;
  assign n8690 = n8688 & n8689;
  assign n8691 = n8681 & n8682;
  assign n8692 = n8680 & n54198;
  assign n8693 = n8678 & n8692;
  assign n8694 = ~n141 & ~n272;
  assign n8695 = n3014 & n8694;
  assign n8696 = ~n246 & ~n259;
  assign n8697 = n8091 & n8696;
  assign n8698 = n8695 & n8697;
  assign n8699 = ~n443 & ~n1997;
  assign n8700 = ~n1125 & ~n1491;
  assign n8701 = n8699 & n8700;
  assign n8702 = n53777 & n8701;
  assign n8703 = n3014 & n8091;
  assign n8704 = ~n272 & ~n443;
  assign n8705 = n8696 & n8704;
  assign n8706 = n8703 & n8705;
  assign n8707 = ~n141 & ~n1997;
  assign n8708 = n8700 & n8707;
  assign n8709 = n53777 & n8708;
  assign n8710 = n8706 & n8709;
  assign n8711 = ~n259 & ~n1125;
  assign n8712 = n8699 & n8711;
  assign n8713 = n8703 & n8712;
  assign n8714 = ~n246 & ~n1491;
  assign n8715 = n8694 & n8714;
  assign n8716 = n53777 & n8715;
  assign n8717 = n8713 & n8716;
  assign n8718 = n8698 & n8702;
  assign n8719 = n53877 & n54198;
  assign n8720 = n53777 & n54094;
  assign n8721 = n8719 & n8720;
  assign n8722 = n8680 & n8703;
  assign n8723 = ~n443 & ~n1125;
  assign n8724 = ~n141 & ~n246;
  assign n8725 = n8723 & n8724;
  assign n8726 = ~n259 & ~n272;
  assign n8727 = ~n1491 & ~n1997;
  assign n8728 = n8726 & n8727;
  assign n8729 = n8725 & n8728;
  assign n8730 = n8722 & n8729;
  assign n8731 = n8721 & n8730;
  assign n8732 = n8693 & n54199;
  assign n8733 = n54197 & n54200;
  assign n8734 = n54094 & n8679;
  assign n8735 = n54198 & n8734;
  assign n8736 = n54197 & n8735;
  assign n8737 = n53877 & n8736;
  assign n8738 = n54196 & n8737;
  assign n8739 = n8091 & n8738;
  assign n8740 = n53777 & n8739;
  assign n8741 = n3014 & n8740;
  assign n8742 = n164 & n8741;
  assign n8743 = ~n1125 & n8742;
  assign n8744 = ~n1997 & n8743;
  assign n8745 = ~n1491 & n8744;
  assign n8746 = ~n272 & n8745;
  assign n8747 = ~n259 & n8746;
  assign n8748 = ~n141 & n8747;
  assign n8749 = ~n246 & n8748;
  assign n8750 = ~n443 & n8749;
  assign n8751 = n54196 & n8733;
  assign n8752 = ~n310 & ~n514;
  assign n8753 = ~n506 & ~n1471;
  assign n8754 = ~n174 & ~n504;
  assign n8755 = n8753 & n8754;
  assign n8756 = n8752 & n8754;
  assign n8757 = n8753 & n8756;
  assign n8758 = n8752 & n8755;
  assign n8759 = ~n1079 & n4026;
  assign n8760 = n2162 & n6897;
  assign n8761 = n8759 & n8760;
  assign n8762 = n54184 & n8761;
  assign n8763 = n2172 & n8753;
  assign n8764 = n2172 & n8755;
  assign n8765 = n8754 & n8763;
  assign n8766 = n4026 & n54203;
  assign n8767 = n6897 & n8766;
  assign n8768 = n293 & n8767;
  assign n8769 = ~n1090 & n8768;
  assign n8770 = ~n1079 & n8769;
  assign n8771 = ~n307 & n8770;
  assign n8772 = ~n310 & n8771;
  assign n8773 = ~n514 & n8772;
  assign n8774 = n8752 & n8753;
  assign n8775 = n2162 & n8774;
  assign n8776 = n6897 & n8754;
  assign n8777 = n8759 & n8776;
  assign n8778 = n54184 & n8777;
  assign n8779 = n8775 & n8778;
  assign n8780 = n54202 & n8761;
  assign n8781 = n54184 & n8780;
  assign n8782 = ~n1079 & n8752;
  assign n8783 = n2162 & n4026;
  assign n8784 = n293 & n6897;
  assign n8785 = n8783 & n8784;
  assign n8786 = n8782 & n8785;
  assign n8787 = n54203 & n8786;
  assign n8788 = n54202 & n8762;
  assign n8789 = n4013 & n4259;
  assign n8790 = n4259 & n4584;
  assign n8791 = n4013 & n8790;
  assign n8792 = n4584 & n8789;
  assign n8793 = ~n852 & ~n1189;
  assign n8794 = ~n660 & ~n1681;
  assign n8795 = ~n1681 & n8793;
  assign n8796 = ~n660 & n8795;
  assign n8797 = n8793 & n8794;
  assign n8798 = ~n901 & ~n957;
  assign n8799 = ~n957 & ~n1703;
  assign n8800 = ~n901 & n8799;
  assign n8801 = ~n1703 & n8798;
  assign n8802 = n54206 & n54207;
  assign n8803 = n54205 & n8802;
  assign n8804 = ~n182 & n1708;
  assign n8805 = n1957 & n2202;
  assign n8806 = n1708 & n1957;
  assign n8807 = ~n215 & n8806;
  assign n8808 = ~n182 & n8807;
  assign n8809 = ~n2201 & n8808;
  assign n8810 = ~n182 & ~n2201;
  assign n8811 = ~n182 & n2202;
  assign n8812 = ~n215 & n8810;
  assign n8813 = n8806 & n54209;
  assign n8814 = n8804 & n8805;
  assign n8815 = n53982 & n54208;
  assign n8816 = n8803 & n8815;
  assign n8817 = ~n1455 & ~n2103;
  assign n8818 = ~n977 & ~n1455;
  assign n8819 = ~n2103 & n8818;
  assign n8820 = ~n977 & n8817;
  assign n8821 = ~n108 & ~n560;
  assign n8822 = n2635 & n8821;
  assign n8823 = ~n612 & ~n823;
  assign n8824 = ~n250 & ~n1535;
  assign n8825 = n8823 & n8824;
  assign n8826 = n8822 & n8825;
  assign n8827 = n2635 & n8825;
  assign n8828 = ~n977 & n8827;
  assign n8829 = ~n2103 & n8828;
  assign n8830 = ~n108 & n8829;
  assign n8831 = ~n560 & n8830;
  assign n8832 = ~n1455 & n8831;
  assign n8833 = ~n977 & ~n2103;
  assign n8834 = ~n108 & n8833;
  assign n8835 = ~n560 & ~n1455;
  assign n8836 = n2635 & n8835;
  assign n8837 = n8825 & n8836;
  assign n8838 = n8834 & n8837;
  assign n8839 = n54210 & n8826;
  assign n8840 = n53496 & n54211;
  assign n8841 = n8816 & n8840;
  assign n8842 = n54204 & n8841;
  assign n8843 = n53493 & n8842;
  assign n8844 = n53493 & n54206;
  assign n8845 = n4259 & n8844;
  assign n8846 = n4013 & n8845;
  assign n8847 = n54208 & n8846;
  assign n8848 = n53982 & n8847;
  assign n8849 = n54201 & n8848;
  assign n8850 = n54211 & n8849;
  assign n8851 = n53496 & n8850;
  assign n8852 = n54204 & n8851;
  assign n8853 = n4584 & n8852;
  assign n8854 = ~n957 & n8853;
  assign n8855 = ~n901 & n8854;
  assign n8856 = ~n1703 & n8855;
  assign n8857 = n54201 & n8843;
  assign n8858 = ~n54194 & ~n54212;
  assign n8859 = n4313 & n6117;
  assign n8860 = ~n415 & ~n591;
  assign n8861 = n7101 & n8860;
  assign n8862 = n8859 & n8861;
  assign n8863 = ~n559 & n1578;
  assign n8864 = ~n211 & ~n651;
  assign n8865 = ~n914 & ~n1485;
  assign n8866 = ~n211 & ~n914;
  assign n8867 = ~n651 & ~n1485;
  assign n8868 = n8866 & n8867;
  assign n8869 = n8864 & n8865;
  assign n8870 = n613 & n2916;
  assign n8871 = n54213 & n8870;
  assign n8872 = n8863 & n8871;
  assign n8873 = n2916 & n7101;
  assign n8874 = n8860 & n8873;
  assign n8875 = n613 & n8874;
  assign n8876 = n4313 & n8875;
  assign n8877 = ~n1485 & n8876;
  assign n8878 = n8863 & n8877;
  assign n8879 = ~n567 & n8878;
  assign n8880 = ~n211 & n8879;
  assign n8881 = ~n914 & n8880;
  assign n8882 = ~n510 & n8881;
  assign n8883 = ~n651 & n8882;
  assign n8884 = n4313 & n7101;
  assign n8885 = n8870 & n8884;
  assign n8886 = ~n567 & ~n1485;
  assign n8887 = ~n651 & ~n914;
  assign n8888 = n8886 & n8887;
  assign n8889 = ~n211 & ~n510;
  assign n8890 = n8860 & n8889;
  assign n8891 = n8888 & n8890;
  assign n8892 = n8863 & n8891;
  assign n8893 = n8885 & n8892;
  assign n8894 = n8862 & n8872;
  assign n8895 = ~n408 & ~n568;
  assign n8896 = ~n568 & ~n1634;
  assign n8897 = ~n408 & n8896;
  assign n8898 = ~n1634 & n8895;
  assign n8899 = ~n499 & ~n750;
  assign n8900 = ~n977 & ~n1644;
  assign n8901 = n8899 & n8900;
  assign n8902 = ~n250 & ~n623;
  assign n8903 = n3134 & n8902;
  assign n8904 = ~n250 & ~n750;
  assign n8905 = n8900 & n8904;
  assign n8906 = ~n499 & ~n623;
  assign n8907 = n3134 & n8906;
  assign n8908 = n8905 & n8907;
  assign n8909 = ~n499 & ~n977;
  assign n8910 = ~n623 & ~n1644;
  assign n8911 = n8909 & n8910;
  assign n8912 = n3134 & n8904;
  assign n8913 = n8911 & n8912;
  assign n8914 = ~n250 & ~n1644;
  assign n8915 = n8909 & n8914;
  assign n8916 = ~n623 & ~n750;
  assign n8917 = n3134 & n8916;
  assign n8918 = n8915 & n8917;
  assign n8919 = n8901 & n8903;
  assign n8920 = n3134 & n54215;
  assign n8921 = ~n977 & n8920;
  assign n8922 = ~n250 & n8921;
  assign n8923 = ~n1644 & n8922;
  assign n8924 = ~n499 & n8923;
  assign n8925 = ~n750 & n8924;
  assign n8926 = ~n623 & n8925;
  assign n8927 = n54215 & n54216;
  assign n8928 = n905 & n5578;
  assign n8929 = ~n789 & ~n1081;
  assign n8930 = n7276 & n8929;
  assign n8931 = n8928 & n8930;
  assign n8932 = ~n565 & ~n631;
  assign n8933 = n2675 & n8932;
  assign n8934 = n1035 & n5198;
  assign n8935 = n8933 & n8934;
  assign n8936 = ~n506 & ~n751;
  assign n8937 = ~n774 & ~n1769;
  assign n8938 = n8936 & n8937;
  assign n8939 = n53815 & n8938;
  assign n8940 = ~n506 & ~n631;
  assign n8941 = n2675 & n8940;
  assign n8942 = n8934 & n8941;
  assign n8943 = ~n565 & ~n774;
  assign n8944 = ~n751 & ~n1769;
  assign n8945 = n8943 & n8944;
  assign n8946 = n53815 & n8945;
  assign n8947 = n8942 & n8946;
  assign n8948 = ~n751 & ~n774;
  assign n8949 = n2675 & n8948;
  assign n8950 = n8934 & n8949;
  assign n8951 = ~n506 & ~n1769;
  assign n8952 = n8932 & n8951;
  assign n8953 = n53815 & n8952;
  assign n8954 = n8950 & n8953;
  assign n8955 = n8935 & n8939;
  assign n8956 = n8930 & n8934;
  assign n8957 = n2675 & n8936;
  assign n8958 = n8928 & n8957;
  assign n8959 = n8932 & n8937;
  assign n8960 = n53815 & n8959;
  assign n8961 = n8958 & n8960;
  assign n8962 = n8956 & n8961;
  assign n8963 = n8931 & n54218;
  assign n8964 = n54217 & n54219;
  assign n8965 = n54214 & n8964;
  assign n8966 = ~n748 & ~n1062;
  assign n8967 = ~n1062 & ~n1196;
  assign n8968 = ~n748 & n8967;
  assign n8969 = ~n1196 & n8966;
  assign n8970 = ~n443 & ~n1478;
  assign n8971 = ~n272 & ~n1535;
  assign n8972 = ~n310 & ~n554;
  assign n8973 = n8971 & n8972;
  assign n8974 = n8970 & n8973;
  assign n8975 = ~n1478 & n8967;
  assign n8976 = ~n310 & n8975;
  assign n8977 = ~n272 & n8976;
  assign n8978 = ~n554 & n8977;
  assign n8979 = ~n1535 & n8978;
  assign n8980 = ~n748 & n8979;
  assign n8981 = ~n443 & n8980;
  assign n8982 = ~n310 & ~n1478;
  assign n8983 = ~n554 & n8982;
  assign n8984 = ~n272 & ~n1062;
  assign n8985 = ~n443 & ~n1196;
  assign n8986 = ~n748 & ~n1535;
  assign n8987 = n8985 & n8986;
  assign n8988 = n8984 & n8987;
  assign n8989 = n8983 & n8988;
  assign n8990 = n54220 & n8974;
  assign n8991 = ~n363 & ~n495;
  assign n8992 = ~n495 & ~n1234;
  assign n8993 = ~n363 & n8992;
  assign n8994 = ~n363 & ~n1234;
  assign n8995 = ~n495 & n8994;
  assign n8996 = ~n1234 & n8991;
  assign n8997 = ~n295 & ~n614;
  assign n8998 = ~n295 & ~n852;
  assign n8999 = ~n614 & n8998;
  assign n9000 = ~n852 & n8997;
  assign n9001 = ~n258 & ~n316;
  assign n9002 = ~n348 & ~n879;
  assign n9003 = ~n316 & ~n348;
  assign n9004 = ~n258 & ~n879;
  assign n9005 = n9003 & n9004;
  assign n9006 = ~n258 & ~n348;
  assign n9007 = ~n316 & ~n879;
  assign n9008 = n9006 & n9007;
  assign n9009 = n9001 & n9002;
  assign n9010 = n54223 & n54224;
  assign n9011 = n54222 & n9010;
  assign n9012 = ~n364 & ~n2042;
  assign n9013 = ~n1124 & n9012;
  assign n9014 = ~n105 & ~n660;
  assign n9015 = n3678 & n9014;
  assign n9016 = ~n1124 & n3678;
  assign n9017 = ~n105 & n9016;
  assign n9018 = ~n660 & n9017;
  assign n9019 = ~n364 & n9018;
  assign n9020 = ~n2042 & n9019;
  assign n9021 = ~n105 & ~n2042;
  assign n9022 = ~n1124 & n9021;
  assign n9023 = ~n364 & ~n660;
  assign n9024 = n3678 & n9023;
  assign n9025 = n9022 & n9024;
  assign n9026 = ~n364 & ~n1124;
  assign n9027 = ~n660 & n9026;
  assign n9028 = n3678 & n9021;
  assign n9029 = n9027 & n9028;
  assign n9030 = n9013 & n9015;
  assign n9031 = n1032 & n2635;
  assign n9032 = n1705 & n5277;
  assign n9033 = n1032 & n5277;
  assign n9034 = n1705 & n2635;
  assign n9035 = n9033 & n9034;
  assign n9036 = n9031 & n9032;
  assign n9037 = n54225 & n54226;
  assign n9038 = n9011 & n9037;
  assign n9039 = n2635 & n54222;
  assign n9040 = n54223 & n9039;
  assign n9041 = n1705 & n9040;
  assign n9042 = n54225 & n9041;
  assign n9043 = n1032 & n9042;
  assign n9044 = n54221 & n9043;
  assign n9045 = n5277 & n9044;
  assign n9046 = ~n316 & n9045;
  assign n9047 = ~n879 & n9046;
  assign n9048 = ~n258 & n9047;
  assign n9049 = ~n348 & n9048;
  assign n9050 = n54221 & n9038;
  assign n9051 = n355 & ~n894;
  assign n9052 = ~n246 & ~n1492;
  assign n9053 = n208 & n9052;
  assign n9054 = n208 & n355;
  assign n9055 = ~n894 & n9054;
  assign n9056 = ~n1492 & n9055;
  assign n9057 = ~n246 & n9056;
  assign n9058 = ~n894 & ~n1492;
  assign n9059 = ~n246 & ~n894;
  assign n9060 = ~n1492 & n9059;
  assign n9061 = ~n246 & n9058;
  assign n9062 = n9054 & n54229;
  assign n9063 = n9051 & n9053;
  assign n9064 = ~n1044 & n2092;
  assign n9065 = n2092 & n53944;
  assign n9066 = ~n1044 & n9065;
  assign n9067 = n53944 & n9064;
  assign n9068 = ~n274 & ~n560;
  assign n9069 = ~n274 & ~n357;
  assign n9070 = ~n560 & n9069;
  assign n9071 = ~n357 & ~n560;
  assign n9072 = ~n274 & n9071;
  assign n9073 = ~n357 & n9068;
  assign n9074 = ~n560 & n2854;
  assign n9075 = ~n274 & n9074;
  assign n9076 = ~n357 & n9075;
  assign n9077 = n2854 & n54231;
  assign n9078 = n54230 & n54232;
  assign n9079 = n54228 & n54230;
  assign n9080 = n54232 & n9079;
  assign n9081 = n54228 & n54232;
  assign n9082 = n54230 & n9081;
  assign n9083 = n54228 & n9078;
  assign n9084 = ~n340 & ~n416;
  assign n9085 = ~n498 & n9084;
  assign n9086 = ~n562 & ~n664;
  assign n9087 = n3369 & n9086;
  assign n9088 = ~n416 & ~n562;
  assign n9089 = ~n416 & ~n664;
  assign n9090 = ~n562 & n9089;
  assign n9091 = ~n664 & n9088;
  assign n9092 = ~n340 & ~n498;
  assign n9093 = n3369 & n9092;
  assign n9094 = n54234 & n9093;
  assign n9095 = n9085 & n9087;
  assign n9096 = n53874 & n54192;
  assign n9097 = n54235 & n9096;
  assign n9098 = n3715 & n4026;
  assign n9099 = n5588 & n9098;
  assign n9100 = n54038 & n9099;
  assign n9101 = ~n498 & n9086;
  assign n9102 = n4026 & n9084;
  assign n9103 = n4026 & n9092;
  assign n9104 = n54234 & n9103;
  assign n9105 = n9101 & n9102;
  assign n9106 = n9096 & n54236;
  assign n9107 = n3369 & n5588;
  assign n9108 = n3369 & n3715;
  assign n9109 = n5588 & n9108;
  assign n9110 = n3715 & n9107;
  assign n9111 = n54038 & n54237;
  assign n9112 = n9106 & n9111;
  assign n9113 = n9097 & n9100;
  assign n9114 = n5588 & n54230;
  assign n9115 = n54038 & n9114;
  assign n9116 = n53874 & n9115;
  assign n9117 = n3369 & n9116;
  assign n9118 = n3715 & n9117;
  assign n9119 = n54228 & n9118;
  assign n9120 = n54232 & n9119;
  assign n9121 = n54192 & n9120;
  assign n9122 = n4026 & n9121;
  assign n9123 = ~n416 & n9122;
  assign n9124 = ~n664 & n9123;
  assign n9125 = ~n562 & n9124;
  assign n9126 = ~n498 & n9125;
  assign n9127 = ~n340 & n9126;
  assign n9128 = n54233 & n54238;
  assign n9129 = n54227 & n54239;
  assign n9130 = n2675 & n5198;
  assign n9131 = n53815 & n9130;
  assign n9132 = n8929 & n9131;
  assign n9133 = n54217 & n9132;
  assign n9134 = n54214 & n9133;
  assign n9135 = n54227 & n9134;
  assign n9136 = n54239 & n9135;
  assign n9137 = n7276 & n9136;
  assign n9138 = n1035 & n9137;
  assign n9139 = n905 & n9138;
  assign n9140 = ~n631 & n9139;
  assign n9141 = n5578 & n9140;
  assign n9142 = ~n565 & n9141;
  assign n9143 = ~n506 & n9142;
  assign n9144 = ~n774 & n9143;
  assign n9145 = ~n751 & n9144;
  assign n9146 = ~n1769 & n9145;
  assign n9147 = n8965 & n9129;
  assign n9148 = ~n54212 & ~n54240;
  assign n9149 = ~n268 & ~n591;
  assign n9150 = ~n404 & ~n824;
  assign n9151 = ~n268 & ~n404;
  assign n9152 = ~n591 & ~n824;
  assign n9153 = n9151 & n9152;
  assign n9154 = n9149 & n9150;
  assign n9155 = ~n250 & ~n740;
  assign n9156 = n2005 & n6300;
  assign n9157 = n9155 & n9156;
  assign n9158 = n6300 & n9155;
  assign n9159 = ~n404 & n9158;
  assign n9160 = ~n584 & n9159;
  assign n9161 = ~n824 & n9160;
  assign n9162 = ~n829 & n9161;
  assign n9163 = ~n268 & n9162;
  assign n9164 = ~n591 & n9163;
  assign n9165 = ~n268 & ~n829;
  assign n9166 = ~n584 & ~n591;
  assign n9167 = n9165 & n9166;
  assign n9168 = n6300 & n9150;
  assign n9169 = n9155 & n9168;
  assign n9170 = n9167 & n9169;
  assign n9171 = ~n404 & ~n584;
  assign n9172 = ~n268 & ~n824;
  assign n9173 = n9171 & n9172;
  assign n9174 = ~n591 & ~n829;
  assign n9175 = n6300 & n9174;
  assign n9176 = n9155 & n9175;
  assign n9177 = n9173 & n9176;
  assign n9178 = n54241 & n9157;
  assign n9179 = ~n440 & ~n983;
  assign n9180 = ~n983 & ~n1031;
  assign n9181 = ~n440 & n9180;
  assign n9182 = ~n1031 & n9179;
  assign n9183 = n53707 & n54243;
  assign n9184 = ~n496 & n3389;
  assign n9185 = n53944 & n9184;
  assign n9186 = n9183 & n9185;
  assign n9187 = ~n822 & ~n1485;
  assign n9188 = ~n292 & ~n357;
  assign n9189 = ~n361 & ~n510;
  assign n9190 = n9188 & n9189;
  assign n9191 = ~n292 & ~n510;
  assign n9192 = ~n292 & ~n1485;
  assign n9193 = ~n822 & n9192;
  assign n9194 = ~n510 & n9193;
  assign n9195 = n9187 & n9191;
  assign n9196 = ~n357 & n54244;
  assign n9197 = ~n361 & n9196;
  assign n9198 = ~n357 & ~n361;
  assign n9199 = n54244 & n9198;
  assign n9200 = ~n357 & ~n822;
  assign n9201 = n9192 & n9200;
  assign n9202 = n9189 & n9201;
  assign n9203 = ~n510 & ~n822;
  assign n9204 = ~n361 & ~n1485;
  assign n9205 = n9188 & n9204;
  assign n9206 = n9203 & n9205;
  assign n9207 = n9187 & n9190;
  assign n9208 = ~n414 & ~n590;
  assign n9209 = n2094 & n9208;
  assign n9210 = ~n777 & ~n1634;
  assign n9211 = ~n212 & ~n317;
  assign n9212 = n9210 & n9211;
  assign n9213 = n9209 & n9212;
  assign n9214 = n54245 & n9213;
  assign n9215 = ~n590 & ~n983;
  assign n9216 = ~n1031 & n9215;
  assign n9217 = n53707 & n9216;
  assign n9218 = n9185 & n9217;
  assign n9219 = ~n414 & ~n440;
  assign n9220 = n2094 & n9219;
  assign n9221 = n9212 & n9220;
  assign n9222 = n54245 & n9221;
  assign n9223 = n9218 & n9222;
  assign n9224 = ~n440 & ~n590;
  assign n9225 = ~n983 & n9224;
  assign n9226 = n53944 & n9225;
  assign n9227 = n53707 & n9184;
  assign n9228 = n9226 & n9227;
  assign n9229 = ~n414 & ~n1031;
  assign n9230 = n2094 & n9229;
  assign n9231 = n9212 & n9230;
  assign n9232 = n54245 & n9231;
  assign n9233 = n9228 & n9232;
  assign n9234 = n9186 & n9214;
  assign n9235 = n9211 & n9227;
  assign n9236 = n9210 & n9235;
  assign n9237 = n54245 & n9236;
  assign n9238 = n53944 & n9237;
  assign n9239 = n54242 & n9238;
  assign n9240 = n2094 & n9239;
  assign n9241 = ~n1031 & n9240;
  assign n9242 = ~n414 & n9241;
  assign n9243 = ~n983 & n9242;
  assign n9244 = ~n440 & n9243;
  assign n9245 = ~n590 & n9244;
  assign n9246 = n54242 & n54246;
  assign n9247 = n4002 & n54247;
  assign n9248 = ~n2201 & n9247;
  assign n9249 = n6866 & n54247;
  assign n9250 = ~n348 & ~n1468;
  assign n9251 = n850 & n9250;
  assign n9252 = n1267 & n5748;
  assign n9253 = n1803 & n7788;
  assign n9254 = n9252 & n9253;
  assign n9255 = n9251 & n9254;
  assign n9256 = ~n246 & ~n274;
  assign n9257 = ~n647 & ~n984;
  assign n9258 = n9256 & n9257;
  assign n9259 = ~n294 & ~n664;
  assign n9260 = ~n311 & ~n420;
  assign n9261 = n9259 & n9260;
  assign n9262 = n9258 & n9261;
  assign n9263 = n53800 & n9262;
  assign n9264 = n850 & n1803;
  assign n9265 = n1267 & n7788;
  assign n9266 = n9264 & n9265;
  assign n9267 = n1267 & n53800;
  assign n9268 = n7788 & n9267;
  assign n9269 = n1803 & n9268;
  assign n9270 = n850 & n9269;
  assign n9271 = n53800 & n9266;
  assign n9272 = ~n984 & n54249;
  assign n9273 = n5748 & n9272;
  assign n9274 = ~n1468 & n9273;
  assign n9275 = ~n294 & n9274;
  assign n9276 = ~n311 & n9275;
  assign n9277 = ~n246 & n9276;
  assign n9278 = ~n664 & n9277;
  assign n9279 = ~n274 & n9278;
  assign n9280 = ~n420 & n9279;
  assign n9281 = ~n647 & n9280;
  assign n9282 = ~n348 & n9281;
  assign n9283 = ~n984 & ~n1468;
  assign n9284 = n9256 & n9283;
  assign n9285 = ~n348 & ~n647;
  assign n9286 = n850 & n9285;
  assign n9287 = n9252 & n9286;
  assign n9288 = n9284 & n9287;
  assign n9289 = n9253 & n9261;
  assign n9290 = n53800 & n9289;
  assign n9291 = n9288 & n9290;
  assign n9292 = ~n246 & ~n664;
  assign n9293 = ~n274 & ~n984;
  assign n9294 = n9292 & n9293;
  assign n9295 = ~n294 & ~n647;
  assign n9296 = n9250 & n9295;
  assign n9297 = n7788 & n9260;
  assign n9298 = n9296 & n9297;
  assign n9299 = n9294 & n9298;
  assign n9300 = n850 & n1267;
  assign n9301 = n1803 & n5748;
  assign n9302 = n9300 & n9301;
  assign n9303 = n53800 & n9302;
  assign n9304 = n9299 & n9303;
  assign n9305 = ~n311 & ~n1468;
  assign n9306 = ~n246 & ~n420;
  assign n9307 = n9305 & n9306;
  assign n9308 = ~n274 & ~n348;
  assign n9309 = ~n664 & ~n984;
  assign n9310 = n9308 & n9309;
  assign n9311 = n5748 & n9295;
  assign n9312 = n9310 & n9311;
  assign n9313 = n9307 & n9312;
  assign n9314 = n54249 & n9313;
  assign n9315 = n9255 & n9263;
  assign n9316 = ~n144 & ~n615;
  assign n9317 = n500 & n9316;
  assign n9318 = n846 & n3273;
  assign n9319 = n9317 & n9318;
  assign n9320 = ~n447 & ~n506;
  assign n9321 = ~n754 & ~n1997;
  assign n9322 = n9320 & n9321;
  assign n9323 = n53791 & n9322;
  assign n9324 = n500 & n9320;
  assign n9325 = n9318 & n9324;
  assign n9326 = n9316 & n9321;
  assign n9327 = n53791 & n9326;
  assign n9328 = n9325 & n9327;
  assign n9329 = n9319 & n9323;
  assign n9330 = ~n465 & ~n1124;
  assign n9331 = ~n1644 & n9330;
  assign n9332 = ~n364 & ~n1042;
  assign n9333 = ~n1042 & n9331;
  assign n9334 = ~n364 & n9333;
  assign n9335 = n9331 & n9332;
  assign n9336 = n4710 & n7015;
  assign n9337 = ~n344 & ~n587;
  assign n9338 = n7276 & n9337;
  assign n9339 = n9336 & n9338;
  assign n9340 = n54252 & n9339;
  assign n9341 = ~n161 & ~n754;
  assign n9342 = ~n144 & ~n447;
  assign n9343 = n9341 & n9342;
  assign n9344 = n4710 & n9337;
  assign n9345 = n9343 & n9344;
  assign n9346 = ~n615 & ~n1997;
  assign n9347 = ~n423 & ~n506;
  assign n9348 = n9346 & n9347;
  assign n9349 = n53791 & n9348;
  assign n9350 = n9345 & n9349;
  assign n9351 = n846 & n7276;
  assign n9352 = n500 & n3273;
  assign n9353 = n9351 & n9352;
  assign n9354 = n54252 & n9353;
  assign n9355 = n9350 & n9354;
  assign n9356 = ~n423 & ~n615;
  assign n9357 = ~n447 & ~n1997;
  assign n9358 = n9356 & n9357;
  assign n9359 = n3273 & n9337;
  assign n9360 = n9358 & n9359;
  assign n9361 = ~n161 & ~n506;
  assign n9362 = ~n144 & ~n754;
  assign n9363 = n9361 & n9362;
  assign n9364 = n53791 & n9363;
  assign n9365 = n9360 & n9364;
  assign n9366 = n500 & n4710;
  assign n9367 = n9351 & n9366;
  assign n9368 = n54252 & n9367;
  assign n9369 = n9365 & n9368;
  assign n9370 = n54251 & n9340;
  assign n9371 = n54180 & n54253;
  assign n9372 = n54250 & n9371;
  assign n9373 = n54162 & n9372;
  assign n9374 = n54248 & n54252;
  assign n9375 = n53791 & n9374;
  assign n9376 = n3273 & n9375;
  assign n9377 = n54162 & n9376;
  assign n9378 = n846 & n9377;
  assign n9379 = n500 & n9378;
  assign n9380 = n9337 & n9379;
  assign n9381 = n7276 & n9380;
  assign n9382 = n4710 & n9381;
  assign n9383 = n54180 & n9382;
  assign n9384 = n54250 & n9383;
  assign n9385 = ~n1997 & n9384;
  assign n9386 = ~n144 & n9385;
  assign n9387 = ~n161 & n9386;
  assign n9388 = ~n506 & n9387;
  assign n9389 = ~n423 & n9388;
  assign n9390 = ~n615 & n9389;
  assign n9391 = ~n447 & n9390;
  assign n9392 = ~n754 & n9391;
  assign n9393 = n54248 & n9373;
  assign n9394 = ~n54240 & ~n54254;
  assign n9395 = n1704 & n4259;
  assign n9396 = ~n346 & ~n450;
  assign n9397 = n8052 & n9396;
  assign n9398 = n9395 & n9397;
  assign n9399 = ~n112 & ~n307;
  assign n9400 = ~n881 & ~n1065;
  assign n9401 = ~n307 & ~n1065;
  assign n9402 = ~n112 & ~n881;
  assign n9403 = n9401 & n9402;
  assign n9404 = n9399 & n9400;
  assign n9405 = n2477 & n3001;
  assign n9406 = n54255 & n9405;
  assign n9407 = ~n552 & ~n663;
  assign n9408 = ~n101 & ~n498;
  assign n9409 = ~n101 & ~n663;
  assign n9410 = ~n552 & n9409;
  assign n9411 = ~n498 & n9410;
  assign n9412 = ~n101 & ~n552;
  assign n9413 = ~n498 & ~n663;
  assign n9414 = n9412 & n9413;
  assign n9415 = n9407 & n9408;
  assign n9416 = n5278 & n54256;
  assign n9417 = n9406 & n9416;
  assign n9418 = n2477 & n4259;
  assign n9419 = n3001 & n9418;
  assign n9420 = n54256 & n9419;
  assign n9421 = n8052 & n9420;
  assign n9422 = n1704 & n9421;
  assign n9423 = n5277 & n9422;
  assign n9424 = n1458 & n9423;
  assign n9425 = ~n881 & n9424;
  assign n9426 = ~n1065 & n9425;
  assign n9427 = ~n112 & n9426;
  assign n9428 = ~n307 & n9427;
  assign n9429 = ~n450 & n9428;
  assign n9430 = ~n346 & n9429;
  assign n9431 = n9397 & n9418;
  assign n9432 = n1704 & n3001;
  assign n9433 = n54255 & n9432;
  assign n9434 = n9416 & n9433;
  assign n9435 = n9431 & n9434;
  assign n9436 = n1458 & n1704;
  assign n9437 = n2477 & n8052;
  assign n9438 = n9436 & n9437;
  assign n9439 = ~n307 & ~n450;
  assign n9440 = n5277 & n9439;
  assign n9441 = n3001 & n4259;
  assign n9442 = n9440 & n9441;
  assign n9443 = ~n112 & ~n346;
  assign n9444 = n9400 & n9443;
  assign n9445 = n54256 & n9444;
  assign n9446 = n9442 & n9445;
  assign n9447 = n9438 & n9446;
  assign n9448 = n9398 & n9417;
  assign n9449 = ~n211 & ~n402;
  assign n9450 = ~n211 & ~n833;
  assign n9451 = ~n402 & n9450;
  assign n9452 = ~n833 & n9449;
  assign n9453 = ~n206 & ~n364;
  assign n9454 = n411 & n9453;
  assign n9455 = ~n206 & ~n211;
  assign n9456 = ~n402 & n9455;
  assign n9457 = ~n833 & n9456;
  assign n9458 = ~n364 & n9457;
  assign n9459 = ~n409 & n9458;
  assign n9460 = ~n410 & n9459;
  assign n9461 = ~n402 & ~n833;
  assign n9462 = ~n364 & n9461;
  assign n9463 = n411 & n9455;
  assign n9464 = n9462 & n9463;
  assign n9465 = n54258 & n9454;
  assign n9466 = ~n1769 & ~n1997;
  assign n9467 = ~n1192 & n2093;
  assign n9468 = ~n1997 & n9467;
  assign n9469 = ~n1769 & n9468;
  assign n9470 = ~n1192 & n9466;
  assign n9471 = n2093 & n9470;
  assign n9472 = n9466 & n9467;
  assign n9473 = n53674 & n54260;
  assign n9474 = n53674 & n54259;
  assign n9475 = n54260 & n9474;
  assign n9476 = n54259 & n9473;
  assign n9477 = ~n914 & ~n1234;
  assign n9478 = n8656 & n9477;
  assign n9479 = ~n221 & ~n354;
  assign n9480 = n1955 & n9479;
  assign n9481 = n9478 & n9480;
  assign n9482 = ~n215 & ~n618;
  assign n9483 = ~n753 & n9482;
  assign n9484 = n749 & n1645;
  assign n9485 = ~n753 & ~n1644;
  assign n9486 = ~n1034 & n9485;
  assign n9487 = n749 & n9482;
  assign n9488 = n9486 & n9487;
  assign n9489 = n9483 & n9484;
  assign n9490 = n749 & n8656;
  assign n9491 = n9477 & n9479;
  assign n9492 = n9490 & n9491;
  assign n9493 = ~n618 & ~n1644;
  assign n9494 = ~n215 & n9493;
  assign n9495 = ~n753 & ~n1034;
  assign n9496 = n1955 & n9495;
  assign n9497 = n9494 & n9496;
  assign n9498 = n9492 & n9497;
  assign n9499 = n1955 & n9477;
  assign n9500 = n9484 & n9499;
  assign n9501 = ~n618 & n9479;
  assign n9502 = ~n215 & ~n753;
  assign n9503 = n8656 & n9502;
  assign n9504 = n9501 & n9503;
  assign n9505 = n9500 & n9504;
  assign n9506 = n9481 & n54262;
  assign n9507 = n53805 & n54263;
  assign n9508 = n54261 & n9507;
  assign n9509 = n54257 & n9508;
  assign n9510 = ~n356 & ~n849;
  assign n9511 = ~n222 & ~n344;
  assign n9512 = n8696 & n9511;
  assign n9513 = n9510 & n9512;
  assign n9514 = n613 & n1642;
  assign n9515 = n903 & n3947;
  assign n9516 = n9514 & n9515;
  assign n9517 = ~n585 & ~n646;
  assign n9518 = ~n269 & ~n735;
  assign n9519 = n9517 & n9518;
  assign n9520 = n53647 & n9519;
  assign n9521 = n9516 & n9520;
  assign n9522 = n3947 & n9510;
  assign n9523 = n3947 & n9511;
  assign n9524 = n9510 & n9523;
  assign n9525 = n9511 & n9522;
  assign n9526 = ~n269 & ~n585;
  assign n9527 = ~n246 & ~n735;
  assign n9528 = ~n246 & ~n585;
  assign n9529 = n9518 & n9528;
  assign n9530 = n9526 & n9527;
  assign n9531 = n53647 & n54265;
  assign n9532 = n613 & n903;
  assign n9533 = ~n259 & ~n646;
  assign n9534 = n1642 & n9533;
  assign n9535 = n9532 & n9534;
  assign n9536 = ~n269 & ~n646;
  assign n9537 = n613 & n9536;
  assign n9538 = n903 & n1642;
  assign n9539 = n9537 & n9538;
  assign n9540 = ~n585 & ~n735;
  assign n9541 = n8696 & n9540;
  assign n9542 = n53647 & n9541;
  assign n9543 = n9539 & n9542;
  assign n9544 = n9531 & n9535;
  assign n9545 = n54264 & n54266;
  assign n9546 = n9511 & n9532;
  assign n9547 = n9510 & n9533;
  assign n9548 = n1642 & n3947;
  assign n9549 = n9547 & n9548;
  assign n9550 = n9531 & n9549;
  assign n9551 = n9546 & n9550;
  assign n9552 = n9513 & n9521;
  assign n9553 = n53647 & n3947;
  assign n9554 = n53891 & n9553;
  assign n9555 = n9510 & n9554;
  assign n9556 = n613 & n9555;
  assign n9557 = n9511 & n9556;
  assign n9558 = n1642 & n9557;
  assign n9559 = n903 & n9558;
  assign n9560 = ~n259 & n9559;
  assign n9561 = ~n246 & n9560;
  assign n9562 = ~n269 & n9561;
  assign n9563 = ~n646 & n9562;
  assign n9564 = ~n735 & n9563;
  assign n9565 = ~n585 & n9564;
  assign n9566 = n53891 & n54267;
  assign n9567 = n54247 & n54268;
  assign n9568 = n53805 & n54260;
  assign n9569 = n53674 & n9568;
  assign n9570 = n1955 & n9569;
  assign n9571 = n54247 & n9570;
  assign n9572 = n54259 & n9571;
  assign n9573 = n54257 & n9572;
  assign n9574 = n9477 & n9573;
  assign n9575 = n749 & n9574;
  assign n9576 = n54268 & n9575;
  assign n9577 = ~n1476 & n9576;
  assign n9578 = ~n215 & n9577;
  assign n9579 = ~n311 & n9578;
  assign n9580 = ~n221 & n9579;
  assign n9581 = ~n1034 & n9580;
  assign n9582 = ~n618 & n9581;
  assign n9583 = ~n1644 & n9582;
  assign n9584 = ~n354 & n9583;
  assign n9585 = ~n753 & n9584;
  assign n9586 = n9509 & n9567;
  assign n9587 = ~n54254 & ~n54269;
  assign n9588 = ~n650 & ~n1769;
  assign n9589 = n897 & n2163;
  assign n9590 = n9588 & n9589;
  assign n9591 = ~n414 & ~n506;
  assign n9592 = ~n414 & ~n1337;
  assign n9593 = ~n506 & n9592;
  assign n9594 = ~n1337 & n9591;
  assign n9595 = ~n513 & ~n659;
  assign n9596 = n494 & n9595;
  assign n9597 = n9184 & n9596;
  assign n9598 = n54270 & n9597;
  assign n9599 = n9184 & n54270;
  assign n9600 = n897 & n9599;
  assign n9601 = n494 & n9600;
  assign n9602 = ~n901 & n9601;
  assign n9603 = ~n659 & n9602;
  assign n9604 = ~n562 & n9603;
  assign n9605 = ~n513 & n9604;
  assign n9606 = ~n650 & n9605;
  assign n9607 = ~n1769 & n9606;
  assign n9608 = n494 & n9588;
  assign n9609 = n2163 & n9608;
  assign n9610 = n897 & n9595;
  assign n9611 = n9184 & n9610;
  assign n9612 = n54270 & n9611;
  assign n9613 = n9609 & n9612;
  assign n9614 = n897 & n9596;
  assign n9615 = ~n650 & ~n901;
  assign n9616 = ~n562 & ~n1769;
  assign n9617 = n9615 & n9616;
  assign n9618 = n9184 & n9617;
  assign n9619 = n54270 & n9618;
  assign n9620 = n9614 & n9619;
  assign n9621 = n9590 & n9598;
  assign n9622 = ~n141 & ~n461;
  assign n9623 = ~n141 & ~n567;
  assign n9624 = ~n568 & n9623;
  assign n9625 = ~n461 & n9624;
  assign n9626 = n569 & n9622;
  assign n9627 = ~n363 & ~n440;
  assign n9628 = ~n363 & ~n733;
  assign n9629 = ~n440 & n9628;
  assign n9630 = ~n733 & n9627;
  assign n9631 = ~n612 & ~n741;
  assign n9632 = n1682 & n9631;
  assign n9633 = ~n363 & ~n612;
  assign n9634 = ~n440 & n9633;
  assign n9635 = ~n733 & ~n741;
  assign n9636 = n1682 & n9635;
  assign n9637 = n9634 & n9636;
  assign n9638 = n54273 & n9632;
  assign n9639 = n1682 & n54272;
  assign n9640 = ~n612 & n9639;
  assign n9641 = ~n440 & n9640;
  assign n9642 = ~n733 & n9641;
  assign n9643 = ~n363 & n9642;
  assign n9644 = ~n741 & n9643;
  assign n9645 = n54272 & n54274;
  assign n9646 = ~n296 & ~n1455;
  assign n9647 = n1869 & n7788;
  assign n9648 = n9646 & n9647;
  assign n9649 = ~n166 & ~n883;
  assign n9650 = n164 & n9649;
  assign n9651 = n1702 & n2691;
  assign n9652 = n5485 & n6614;
  assign n9653 = n9651 & n9652;
  assign n9654 = n9650 & n9653;
  assign n9655 = n1869 & n6614;
  assign n9656 = n9646 & n9655;
  assign n9657 = n7788 & n9649;
  assign n9658 = n164 & n2691;
  assign n9659 = n1702 & n5485;
  assign n9660 = n9658 & n9659;
  assign n9661 = n9657 & n9660;
  assign n9662 = n9656 & n9661;
  assign n9663 = n164 & n7788;
  assign n9664 = n2691 & n9663;
  assign n9665 = ~n166 & ~n789;
  assign n9666 = ~n179 & ~n296;
  assign n9667 = n9665 & n9666;
  assign n9668 = ~n883 & ~n1455;
  assign n9669 = n1702 & n9668;
  assign n9670 = n9652 & n9669;
  assign n9671 = n9667 & n9670;
  assign n9672 = n9664 & n9671;
  assign n9673 = n9648 & n9654;
  assign n9674 = n54275 & n54276;
  assign n9675 = n54271 & n9674;
  assign n9676 = n53531 & n53880;
  assign n9677 = n5485 & n9651;
  assign n9678 = n7788 & n9677;
  assign n9679 = n53880 & n9678;
  assign n9680 = n53531 & n9679;
  assign n9681 = n54271 & n9680;
  assign n9682 = n54275 & n9681;
  assign n9683 = n6614 & n9682;
  assign n9684 = n164 & n9683;
  assign n9685 = ~n883 & n9684;
  assign n9686 = ~n296 & n9685;
  assign n9687 = ~n179 & n9686;
  assign n9688 = ~n166 & n9687;
  assign n9689 = ~n1455 & n9688;
  assign n9690 = ~n789 & n9689;
  assign n9691 = n9675 & n9676;
  assign n9692 = ~n54269 & ~n54277;
  assign n9693 = ~n741 & n2975;
  assign n9694 = n2975 & n3950;
  assign n9695 = ~n741 & n9694;
  assign n9696 = n3950 & n9693;
  assign n9697 = n449 & n2675;
  assign n9698 = n5652 & n8860;
  assign n9699 = n2675 & n5652;
  assign n9700 = n449 & n8860;
  assign n9701 = n9699 & n9700;
  assign n9702 = n449 & n5652;
  assign n9703 = n2675 & n8860;
  assign n9704 = n9702 & n9703;
  assign n9705 = n9697 & n9698;
  assign n9706 = ~n829 & ~n1646;
  assign n9707 = ~n510 & n9706;
  assign n9708 = ~n510 & ~n1646;
  assign n9709 = ~n829 & n9708;
  assign n9710 = ~n1646 & n7903;
  assign n9711 = ~n101 & ~n271;
  assign n9712 = ~n733 & ~n1477;
  assign n9713 = ~n271 & ~n733;
  assign n9714 = ~n101 & ~n1477;
  assign n9715 = n9713 & n9714;
  assign n9716 = n9711 & n9712;
  assign n9717 = n54280 & n54281;
  assign n9718 = n54279 & n9717;
  assign n9719 = n54278 & n54280;
  assign n9720 = n8860 & n9719;
  assign n9721 = n2675 & n9720;
  assign n9722 = n5652 & n9721;
  assign n9723 = ~n1477 & n9722;
  assign n9724 = ~n101 & n9723;
  assign n9725 = ~n271 & n9724;
  assign n9726 = ~n733 & n9725;
  assign n9727 = ~n447 & n9726;
  assign n9728 = ~n448 & n9727;
  assign n9729 = n54278 & n9718;
  assign n9730 = ~n212 & ~n627;
  assign n9731 = ~n348 & ~n1059;
  assign n9732 = ~n212 & ~n1059;
  assign n9733 = ~n348 & ~n627;
  assign n9734 = n9732 & n9733;
  assign n9735 = ~n212 & ~n348;
  assign n9736 = ~n627 & ~n1059;
  assign n9737 = n9735 & n9736;
  assign n9738 = n9730 & n9731;
  assign n9739 = ~n611 & ~n896;
  assign n9740 = ~n559 & ~n894;
  assign n9741 = n3878 & n9740;
  assign n9742 = n3878 & n9739;
  assign n9743 = ~n894 & n9742;
  assign n9744 = ~n559 & n9743;
  assign n9745 = n9739 & n9741;
  assign n9746 = ~n212 & n54284;
  assign n9747 = ~n1059 & n9746;
  assign n9748 = ~n627 & n9747;
  assign n9749 = ~n348 & n9748;
  assign n9750 = n9732 & n9740;
  assign n9751 = n3878 & n9733;
  assign n9752 = n9739 & n9751;
  assign n9753 = n9750 & n9752;
  assign n9754 = n54283 & n54284;
  assign n9755 = ~n274 & ~n646;
  assign n9756 = ~n274 & ~n291;
  assign n9757 = ~n646 & n9756;
  assign n9758 = ~n291 & ~n646;
  assign n9759 = ~n274 & n9758;
  assign n9760 = ~n291 & n9755;
  assign n9761 = ~n848 & ~n851;
  assign n9762 = ~n1085 & ~n1472;
  assign n9763 = n9761 & n9762;
  assign n9764 = n54106 & n9763;
  assign n9765 = n54286 & n9764;
  assign n9766 = ~n161 & ~n742;
  assign n9767 = ~n172 & ~n294;
  assign n9768 = n7016 & n9767;
  assign n9769 = n7016 & n9766;
  assign n9770 = n9767 & n9769;
  assign n9771 = n9766 & n9768;
  assign n9772 = n424 & n624;
  assign n9773 = n3273 & n4884;
  assign n9774 = n9772 & n9773;
  assign n9775 = n424 & n9766;
  assign n9776 = n9767 & n9775;
  assign n9777 = n624 & n3273;
  assign n9778 = n4884 & n7016;
  assign n9779 = n9777 & n9778;
  assign n9780 = n9776 & n9779;
  assign n9781 = n54287 & n9774;
  assign n9782 = n9762 & n9767;
  assign n9783 = n54286 & n9782;
  assign n9784 = n54106 & n9783;
  assign n9785 = n9766 & n9773;
  assign n9786 = n624 & n9761;
  assign n9787 = n424 & n7016;
  assign n9788 = n9786 & n9787;
  assign n9789 = n9785 & n9788;
  assign n9790 = n9784 & n9789;
  assign n9791 = n9765 & n54288;
  assign n9792 = n54285 & n54289;
  assign n9793 = n54106 & n9766;
  assign n9794 = n54286 & n9793;
  assign n9795 = n4884 & n9794;
  assign n9796 = n3273 & n9795;
  assign n9797 = n54282 & n9796;
  assign n9798 = n54285 & n9797;
  assign n9799 = n7016 & n9798;
  assign n9800 = n424 & n9799;
  assign n9801 = n624 & n9800;
  assign n9802 = ~n1085 & n9801;
  assign n9803 = ~n1472 & n9802;
  assign n9804 = ~n172 & n9803;
  assign n9805 = ~n294 & n9804;
  assign n9806 = ~n848 & n9805;
  assign n9807 = ~n851 & n9806;
  assign n9808 = n54282 & n9792;
  assign n9809 = n1265 & n5060;
  assign n9810 = n5390 & n7350;
  assign n9811 = n9809 & n9810;
  assign n9812 = ~n585 & ~n649;
  assign n9813 = ~n649 & ~n883;
  assign n9814 = ~n585 & n9813;
  assign n9815 = ~n883 & n9812;
  assign n9816 = n6934 & n54291;
  assign n9817 = n9811 & n9816;
  assign n9818 = ~n402 & ~n750;
  assign n9819 = ~n402 & n53518;
  assign n9820 = ~n750 & n9819;
  assign n9821 = n53518 & n9818;
  assign n9822 = n7473 & n8138;
  assign n9823 = n9477 & n9822;
  assign n9824 = n54292 & n9823;
  assign n9825 = n1265 & n9813;
  assign n9826 = n5060 & n5390;
  assign n9827 = n9825 & n9826;
  assign n9828 = ~n585 & ~n1912;
  assign n9829 = ~n564 & n9828;
  assign n9830 = n6934 & n9829;
  assign n9831 = n9827 & n9830;
  assign n9832 = n7350 & n7473;
  assign n9833 = n9477 & n9832;
  assign n9834 = n54292 & n9833;
  assign n9835 = n9831 & n9834;
  assign n9836 = n9817 & n9824;
  assign n9837 = n6934 & n7473;
  assign n9838 = n54292 & n9837;
  assign n9839 = n7350 & n9838;
  assign n9840 = n54032 & n9839;
  assign n9841 = n5060 & n9840;
  assign n9842 = n1265 & n9841;
  assign n9843 = n5390 & n9842;
  assign n9844 = n9477 & n9843;
  assign n9845 = ~n883 & n9844;
  assign n9846 = ~n564 & n9845;
  assign n9847 = ~n649 & n9846;
  assign n9848 = ~n1912 & n9847;
  assign n9849 = ~n585 & n9848;
  assign n9850 = n54032 & n54293;
  assign n9851 = ~n440 & ~n1468;
  assign n9852 = ~n1468 & n4916;
  assign n9853 = ~n440 & n9852;
  assign n9854 = n4916 & n9851;
  assign n9855 = ~n823 & ~n1486;
  assign n9856 = ~n823 & ~n1033;
  assign n9857 = ~n1486 & n9856;
  assign n9858 = ~n1033 & ~n1486;
  assign n9859 = ~n823 & n9858;
  assign n9860 = ~n1033 & n9855;
  assign n9861 = ~n414 & ~n660;
  assign n9862 = ~n465 & n8929;
  assign n9863 = ~n414 & ~n465;
  assign n9864 = ~n660 & n9863;
  assign n9865 = n8929 & n9864;
  assign n9866 = n9861 & n9862;
  assign n9867 = n54296 & n54297;
  assign n9868 = n54295 & n54296;
  assign n9869 = n8929 & n9868;
  assign n9870 = ~n414 & n9869;
  assign n9871 = ~n660 & n9870;
  assign n9872 = ~n465 & n9871;
  assign n9873 = n54295 & n9867;
  assign n9874 = ~n902 & n5059;
  assign n9875 = n5115 & n6867;
  assign n9876 = n8092 & n9875;
  assign n9877 = ~n902 & ~n1088;
  assign n9878 = ~n1466 & n9877;
  assign n9879 = ~n1487 & n9878;
  assign n9880 = ~n560 & n9879;
  assign n9881 = ~n975 & n9880;
  assign n9882 = ~n269 & n9881;
  assign n9883 = ~n356 & n9882;
  assign n9884 = ~n776 & n9883;
  assign n9885 = ~n902 & ~n1487;
  assign n9886 = ~n1466 & n9885;
  assign n9887 = n5059 & n6867;
  assign n9888 = n8092 & n9887;
  assign n9889 = n9886 & n9888;
  assign n9890 = ~n1487 & n6867;
  assign n9891 = ~n560 & ~n1466;
  assign n9892 = ~n356 & ~n975;
  assign n9893 = ~n776 & ~n902;
  assign n9894 = n9892 & n9893;
  assign n9895 = n9891 & n9894;
  assign n9896 = n9890 & n9895;
  assign n9897 = n9874 & n9876;
  assign n9898 = ~n353 & ~n408;
  assign n9899 = ~n353 & ~n360;
  assign n9900 = ~n408 & ~n493;
  assign n9901 = n9899 & n9900;
  assign n9902 = n6892 & n9898;
  assign n9903 = n749 & n775;
  assign n9904 = n54300 & n9903;
  assign n9905 = ~n316 & ~n499;
  assign n9906 = ~n316 & ~n1490;
  assign n9907 = ~n514 & n9906;
  assign n9908 = ~n499 & n9907;
  assign n9909 = n1868 & n9905;
  assign n9910 = ~n1703 & ~n2042;
  assign n9911 = ~n948 & n9910;
  assign n9912 = n54301 & n9911;
  assign n9913 = ~n948 & ~n2042;
  assign n9914 = ~n360 & ~n1703;
  assign n9915 = n9913 & n9914;
  assign n9916 = n9903 & n9915;
  assign n9917 = ~n493 & n9898;
  assign n9918 = n54301 & n9917;
  assign n9919 = n9916 & n9918;
  assign n9920 = n9904 & n9912;
  assign n9921 = ~n216 & n2093;
  assign n9922 = n2093 & n3780;
  assign n9923 = ~n216 & n9922;
  assign n9924 = ~n216 & n3780;
  assign n9925 = n2093 & n9924;
  assign n9926 = n3780 & n9921;
  assign n9927 = n882 & n2476;
  assign n9928 = n9588 & n9927;
  assign n9929 = n54303 & n9928;
  assign n9930 = ~n408 & ~n881;
  assign n9931 = ~n353 & ~n650;
  assign n9932 = n9930 & n9931;
  assign n9933 = n2326 & n9913;
  assign n9934 = n9932 & n9933;
  assign n9935 = ~n493 & ~n1769;
  assign n9936 = ~n360 & n9935;
  assign n9937 = n54301 & n9936;
  assign n9938 = n9934 & n9937;
  assign n9939 = n749 & n2476;
  assign n9940 = n775 & n9939;
  assign n9941 = n54303 & n9940;
  assign n9942 = n9938 & n9941;
  assign n9943 = n54302 & n9929;
  assign n9944 = n54299 & n54304;
  assign n9945 = n54298 & n9944;
  assign n9946 = n54294 & n9945;
  assign n9947 = n54301 & n54303;
  assign n9948 = n54294 & n9947;
  assign n9949 = n54298 & n9948;
  assign n9950 = n54290 & n9949;
  assign n9951 = n54299 & n9950;
  assign n9952 = n775 & n9951;
  assign n9953 = n2476 & n9952;
  assign n9954 = n2326 & n9953;
  assign n9955 = n749 & n9954;
  assign n9956 = ~n881 & n9955;
  assign n9957 = ~n948 & n9956;
  assign n9958 = ~n408 & n9957;
  assign n9959 = ~n493 & n9958;
  assign n9960 = ~n360 & n9959;
  assign n9961 = ~n353 & n9960;
  assign n9962 = ~n650 & n9961;
  assign n9963 = ~n2042 & n9962;
  assign n9964 = ~n1769 & n9963;
  assign n9965 = n54290 & n9946;
  assign n9966 = ~n54277 & ~n54305;
  assign n9967 = n54277 & n54305;
  assign n9968 = ~n9966 & ~n9967;
  assign n9969 = ~n491 & ~n776;
  assign n9970 = n1391 & n9969;
  assign n9971 = n3371 & n9970;
  assign n9972 = n6482 & n8091;
  assign n9973 = ~n1280 & ~n1646;
  assign n9974 = ~n1280 & n3742;
  assign n9975 = ~n1646 & n9974;
  assign n9976 = n3742 & n9973;
  assign n9977 = n9972 & n54306;
  assign n9978 = n9971 & n9977;
  assign n9979 = ~n628 & ~n650;
  assign n9980 = ~n1044 & n9979;
  assign n9981 = ~n222 & ~n410;
  assign n9982 = ~n218 & ~n584;
  assign n9983 = n9981 & n9982;
  assign n9984 = ~n628 & ~n1044;
  assign n9985 = ~n218 & n9984;
  assign n9986 = ~n222 & n9985;
  assign n9987 = ~n584 & n9986;
  assign n9988 = ~n410 & n9987;
  assign n9989 = ~n650 & n9988;
  assign n9990 = ~n410 & ~n1044;
  assign n9991 = ~n628 & n9990;
  assign n9992 = ~n222 & ~n650;
  assign n9993 = n9982 & n9992;
  assign n9994 = n9991 & n9993;
  assign n9995 = ~n222 & ~n1044;
  assign n9996 = ~n1044 & n9981;
  assign n9997 = ~n410 & n9995;
  assign n9998 = n9979 & n9982;
  assign n9999 = n54308 & n9998;
  assign n10000 = n9980 & n9983;
  assign n10001 = ~n554 & ~n823;
  assign n10002 = n1705 & n1716;
  assign n10003 = n10001 & n10002;
  assign n10004 = n54307 & n10003;
  assign n10005 = n9969 & n10001;
  assign n10006 = n9972 & n10005;
  assign n10007 = n3371 & n54306;
  assign n10008 = n3371 & n10005;
  assign n10009 = n9977 & n10008;
  assign n10010 = n10006 & n10007;
  assign n10011 = n1391 & n1705;
  assign n10012 = n1391 & n1716;
  assign n10013 = n1705 & n10012;
  assign n10014 = n1716 & n10011;
  assign n10015 = n54307 & n54310;
  assign n10016 = n54309 & n10015;
  assign n10017 = n9978 & n10004;
  assign n10018 = n1705 & n54306;
  assign n10019 = n3371 & n10018;
  assign n10020 = n53594 & n10019;
  assign n10021 = n54307 & n10020;
  assign n10022 = n8091 & n10021;
  assign n10023 = n1391 & n10022;
  assign n10024 = n6482 & n10023;
  assign n10025 = n1716 & n10024;
  assign n10026 = ~n554 & n10025;
  assign n10027 = ~n823 & n10026;
  assign n10028 = ~n491 & n10027;
  assign n10029 = ~n776 & n10028;
  assign n10030 = n53594 & n54311;
  assign n10031 = ~n902 & ~n1681;
  assign n10032 = ~n294 & n6326;
  assign n10033 = ~n294 & n10031;
  assign n10034 = n6326 & n10033;
  assign n10035 = n10031 & n10032;
  assign n10036 = n6150 & n6479;
  assign n10037 = ~n321 & ~n1059;
  assign n10038 = n897 & n10037;
  assign n10039 = n10036 & n10038;
  assign n10040 = n54252 & n10039;
  assign n10041 = n54313 & n10040;
  assign n10042 = n180 & n1197;
  assign n10043 = n5873 & n7997;
  assign n10044 = n10042 & n10043;
  assign n10045 = ~n623 & ~n957;
  assign n10046 = ~n957 & n5113;
  assign n10047 = ~n623 & n10046;
  assign n10048 = n5113 & n10045;
  assign n10049 = ~n212 & ~n565;
  assign n10050 = ~n1034 & ~n1680;
  assign n10051 = ~n212 & ~n1034;
  assign n10052 = ~n565 & ~n1680;
  assign n10053 = n10051 & n10052;
  assign n10054 = n10049 & n10050;
  assign n10055 = n54314 & n54315;
  assign n10056 = n1197 & n54314;
  assign n10057 = n180 & n10056;
  assign n10058 = n5873 & n10057;
  assign n10059 = ~n1680 & n10058;
  assign n10060 = ~n112 & n10059;
  assign n10061 = ~n212 & n10060;
  assign n10062 = ~n565 & n10061;
  assign n10063 = ~n1034 & n10062;
  assign n10064 = ~n363 & n10063;
  assign n10065 = ~n212 & ~n1680;
  assign n10066 = n5873 & n10065;
  assign n10067 = n10042 & n10066;
  assign n10068 = ~n363 & ~n1034;
  assign n10069 = ~n112 & ~n565;
  assign n10070 = n10068 & n10069;
  assign n10071 = n54314 & n10070;
  assign n10072 = n10067 & n10071;
  assign n10073 = n10044 & n10055;
  assign n10074 = ~n833 & ~n1466;
  assign n10075 = n417 & n10074;
  assign n10076 = n445 & n4587;
  assign n10077 = n10075 & n10076;
  assign n10078 = ~n256 & n2577;
  assign n10079 = n3780 & n4753;
  assign n10080 = n10078 & n10079;
  assign n10081 = n417 & n3780;
  assign n10082 = n4587 & n4753;
  assign n10083 = n10081 & n10082;
  assign n10084 = n445 & n10074;
  assign n10085 = n10078 & n10084;
  assign n10086 = n10083 & n10085;
  assign n10087 = n10077 & n10080;
  assign n10088 = n54316 & n54317;
  assign n10089 = n445 & n10078;
  assign n10090 = n54252 & n10089;
  assign n10091 = n897 & n10090;
  assign n10092 = n4753 & n10091;
  assign n10093 = n54313 & n10092;
  assign n10094 = n54316 & n10093;
  assign n10095 = n417 & n10094;
  assign n10096 = n6150 & n10095;
  assign n10097 = n3780 & n10096;
  assign n10098 = n4587 & n10097;
  assign n10099 = ~n1466 & n10098;
  assign n10100 = ~n1081 & n10099;
  assign n10101 = ~n321 & n10100;
  assign n10102 = ~n1059 & n10101;
  assign n10103 = ~n833 & n10102;
  assign n10104 = ~n466 & n10103;
  assign n10105 = n4753 & n6479;
  assign n10106 = n897 & n6150;
  assign n10107 = n10105 & n10106;
  assign n10108 = n54313 & n10107;
  assign n10109 = n54252 & n10108;
  assign n10110 = n417 & n10037;
  assign n10111 = n10076 & n10110;
  assign n10112 = n3780 & n10074;
  assign n10113 = n10078 & n10112;
  assign n10114 = n10111 & n10113;
  assign n10115 = n54316 & n10114;
  assign n10116 = n10109 & n10115;
  assign n10117 = n897 & n3780;
  assign n10118 = n417 & n445;
  assign n10119 = n10117 & n10118;
  assign n10120 = n54252 & n10119;
  assign n10121 = n54313 & n10120;
  assign n10122 = ~n1059 & ~n1466;
  assign n10123 = n4753 & n10122;
  assign n10124 = n4587 & n6150;
  assign n10125 = n10123 & n10124;
  assign n10126 = ~n321 & ~n833;
  assign n10127 = n6479 & n10126;
  assign n10128 = n10078 & n10127;
  assign n10129 = n10125 & n10128;
  assign n10130 = n54316 & n10129;
  assign n10131 = n10121 & n10130;
  assign n10132 = n10041 & n10088;
  assign n10133 = n6535 & n7016;
  assign n10134 = n2257 & n8319;
  assign n10135 = n10133 & n10134;
  assign n10136 = ~n646 & ~n771;
  assign n10137 = ~n881 & n10136;
  assign n10138 = n4833 & n5588;
  assign n10139 = n10137 & n10138;
  assign n10140 = n4833 & n7016;
  assign n10141 = n5588 & n6535;
  assign n10142 = n5588 & n7016;
  assign n10143 = n6535 & n10142;
  assign n10144 = n4833 & n10143;
  assign n10145 = n10140 & n10141;
  assign n10146 = ~n881 & n54319;
  assign n10147 = ~n422 & n10146;
  assign n10148 = ~n250 & n10147;
  assign n10149 = ~n440 & n10148;
  assign n10150 = ~n646 & n10149;
  assign n10151 = ~n771 & n10150;
  assign n10152 = ~n585 & n10151;
  assign n10153 = n2257 & n7016;
  assign n10154 = n10138 & n10153;
  assign n10155 = ~n440 & ~n881;
  assign n10156 = ~n585 & n10155;
  assign n10157 = n6535 & n10136;
  assign n10158 = n10156 & n10157;
  assign n10159 = n10154 & n10158;
  assign n10160 = ~n585 & ~n771;
  assign n10161 = ~n440 & n10160;
  assign n10162 = ~n646 & ~n881;
  assign n10163 = n2257 & n10162;
  assign n10164 = n10161 & n10163;
  assign n10165 = n54319 & n10164;
  assign n10166 = n10135 & n10139;
  assign n10167 = n318 & n712;
  assign n10168 = n2454 & n3086;
  assign n10169 = n10167 & n10168;
  assign n10170 = ~n360 & ~n748;
  assign n10171 = n293 & ~n748;
  assign n10172 = ~n360 & n10171;
  assign n10173 = n293 & n10170;
  assign n10174 = ~n207 & ~n459;
  assign n10175 = ~n495 & ~n983;
  assign n10176 = ~n207 & ~n983;
  assign n10177 = ~n459 & ~n495;
  assign n10178 = n10176 & n10177;
  assign n10179 = n10174 & n10175;
  assign n10180 = n54321 & n54322;
  assign n10181 = n10169 & n10180;
  assign n10182 = ~n268 & ~n753;
  assign n10183 = ~n617 & ~n774;
  assign n10184 = ~n751 & ~n1033;
  assign n10185 = n10183 & n10184;
  assign n10186 = n10182 & n10183;
  assign n10187 = n10184 & n10186;
  assign n10188 = n10182 & n10185;
  assign n10189 = n5199 & n7307;
  assign n10190 = n7473 & n8793;
  assign n10191 = n10189 & n10190;
  assign n10192 = n54323 & n10191;
  assign n10193 = n318 & n5199;
  assign n10194 = n712 & n2454;
  assign n10195 = n10193 & n10194;
  assign n10196 = n10180 & n10195;
  assign n10197 = n7307 & n7473;
  assign n10198 = n3086 & n8793;
  assign n10199 = n10197 & n10198;
  assign n10200 = n54323 & n10199;
  assign n10201 = n10196 & n10200;
  assign n10202 = n10181 & n10192;
  assign n10203 = n54320 & n54324;
  assign n10204 = n54318 & n10203;
  assign n10205 = n7473 & n54321;
  assign n10206 = n10182 & n10205;
  assign n10207 = n10184 & n10206;
  assign n10208 = n10183 & n10207;
  assign n10209 = n7307 & n10208;
  assign n10210 = n54320 & n10209;
  assign n10211 = n54312 & n10210;
  assign n10212 = n54318 & n10211;
  assign n10213 = n5199 & n10212;
  assign n10214 = n2454 & n10213;
  assign n10215 = n3086 & n10214;
  assign n10216 = n712 & n10215;
  assign n10217 = n318 & n10216;
  assign n10218 = n8793 & n10217;
  assign n10219 = ~n983 & n10218;
  assign n10220 = ~n207 & n10219;
  assign n10221 = ~n495 & n10220;
  assign n10222 = ~n459 & n10221;
  assign n10223 = n54312 & n10203;
  assign n10224 = n54318 & n10223;
  assign n10225 = n54312 & n10204;
  assign n10226 = n54305 & n54325;
  assign n10227 = n185 & n1267;
  assign n10228 = n1128 & n4071;
  assign n10229 = n1128 & n1267;
  assign n10230 = n185 & n4071;
  assign n10231 = n10229 & n10230;
  assign n10232 = n10227 & n10228;
  assign n10233 = ~n259 & ~n291;
  assign n10234 = ~n259 & ~n773;
  assign n10235 = ~n291 & n10234;
  assign n10236 = ~n773 & n10233;
  assign n10237 = n54018 & n54327;
  assign n10238 = ~n562 & ~n2109;
  assign n10239 = ~n1477 & n10238;
  assign n10240 = n424 & n2326;
  assign n10241 = n10239 & n10240;
  assign n10242 = n10237 & n10241;
  assign n10243 = n1128 & n2326;
  assign n10244 = n10227 & n10243;
  assign n10245 = ~n291 & n4071;
  assign n10246 = n424 & n10234;
  assign n10247 = n10245 & n10246;
  assign n10248 = n54018 & n10239;
  assign n10249 = n10247 & n10248;
  assign n10250 = n10244 & n10249;
  assign n10251 = n54326 & n10242;
  assign n10252 = ~n466 & ~n510;
  assign n10253 = ~n466 & ~n498;
  assign n10254 = ~n510 & n10253;
  assign n10255 = ~n498 & ~n510;
  assign n10256 = ~n466 & n10255;
  assign n10257 = ~n498 & n10252;
  assign n10258 = n772 & n54329;
  assign n10259 = n772 & n53935;
  assign n10260 = ~n498 & n10259;
  assign n10261 = ~n510 & n10260;
  assign n10262 = ~n466 & n10261;
  assign n10263 = n53935 & n10258;
  assign n10264 = n54221 & n54330;
  assign n10265 = n1267 & n10239;
  assign n10266 = n185 & n10265;
  assign n10267 = n54018 & n10266;
  assign n10268 = n54330 & n10267;
  assign n10269 = n54221 & n10268;
  assign n10270 = n1128 & n10269;
  assign n10271 = n2326 & n10270;
  assign n10272 = n424 & n10271;
  assign n10273 = ~n291 & n10272;
  assign n10274 = ~n259 & n10273;
  assign n10275 = ~n340 & n10274;
  assign n10276 = ~n773 & n10275;
  assign n10277 = ~n741 & n10276;
  assign n10278 = n54328 & n10264;
  assign n10279 = n1035 & n2537;
  assign n10280 = n1067 & n4020;
  assign n10281 = n10279 & n10280;
  assign n10282 = n53448 & n10281;
  assign n10283 = ~n319 & ~n588;
  assign n10284 = ~n513 & ~n588;
  assign n10285 = ~n319 & n10284;
  assign n10286 = ~n319 & ~n513;
  assign n10287 = ~n588 & n10286;
  assign n10288 = ~n513 & n10283;
  assign n10289 = ~n319 & n7646;
  assign n10290 = ~n513 & n10289;
  assign n10291 = ~n588 & n10290;
  assign n10292 = n7646 & n54332;
  assign n10293 = n54230 & n54333;
  assign n10294 = n54230 & n10281;
  assign n10295 = n53448 & n54333;
  assign n10296 = n10294 & n10295;
  assign n10297 = n10282 & n10293;
  assign n10298 = ~n662 & ~n751;
  assign n10299 = n1955 & n10298;
  assign n10300 = ~n354 & ~n559;
  assign n10301 = ~n623 & ~n852;
  assign n10302 = n10300 & n10301;
  assign n10303 = n1955 & n10300;
  assign n10304 = n10298 & n10301;
  assign n10305 = n10303 & n10304;
  assign n10306 = n10299 & n10302;
  assign n10307 = ~n256 & ~n628;
  assign n10308 = ~n503 & ~n1881;
  assign n10309 = ~n256 & ~n1881;
  assign n10310 = ~n503 & ~n628;
  assign n10311 = n10309 & n10310;
  assign n10312 = n10307 & n10308;
  assign n10313 = n7101 & n9259;
  assign n10314 = n54336 & n10313;
  assign n10315 = n1955 & n7101;
  assign n10316 = n7101 & n10300;
  assign n10317 = n10301 & n10316;
  assign n10318 = n1955 & n10317;
  assign n10319 = n10302 & n10315;
  assign n10320 = ~n628 & n54337;
  assign n10321 = ~n662 & n10320;
  assign n10322 = ~n294 & n10321;
  assign n10323 = ~n256 & n10322;
  assign n10324 = ~n664 & n10323;
  assign n10325 = ~n503 & n10324;
  assign n10326 = ~n751 & n10325;
  assign n10327 = ~n1881 & n10326;
  assign n10328 = n7101 & n10298;
  assign n10329 = n10302 & n10328;
  assign n10330 = ~n294 & ~n503;
  assign n10331 = ~n628 & ~n664;
  assign n10332 = n10330 & n10331;
  assign n10333 = n1955 & n10309;
  assign n10334 = n10332 & n10333;
  assign n10335 = n10329 & n10334;
  assign n10336 = ~n628 & ~n662;
  assign n10337 = ~n256 & ~n664;
  assign n10338 = n10336 & n10337;
  assign n10339 = ~n751 & ~n1881;
  assign n10340 = n10330 & n10339;
  assign n10341 = n10338 & n10340;
  assign n10342 = n54337 & n10341;
  assign n10343 = n54335 & n10314;
  assign n10344 = ~n451 & ~n742;
  assign n10345 = ~n742 & ~n957;
  assign n10346 = ~n829 & n10345;
  assign n10347 = ~n451 & n10346;
  assign n10348 = ~n742 & ~n829;
  assign n10349 = ~n451 & ~n957;
  assign n10350 = n10348 & n10349;
  assign n10351 = n3951 & n10344;
  assign n10352 = ~n618 & ~n788;
  assign n10353 = ~n618 & ~n901;
  assign n10354 = ~n788 & n10353;
  assign n10355 = ~n788 & ~n901;
  assign n10356 = ~n618 & n10355;
  assign n10357 = ~n901 & n10352;
  assign n10358 = ~n404 & ~n659;
  assign n10359 = ~n420 & ~n450;
  assign n10360 = ~n450 & ~n659;
  assign n10361 = ~n404 & ~n420;
  assign n10362 = n10360 & n10361;
  assign n10363 = n10358 & n10359;
  assign n10364 = n54340 & n54341;
  assign n10365 = n54339 & n54341;
  assign n10366 = n54340 & n10365;
  assign n10367 = n54339 & n10364;
  assign n10368 = n54338 & n54342;
  assign n10369 = n1067 & n10361;
  assign n10370 = n1035 & n4020;
  assign n10371 = n10369 & n10370;
  assign n10372 = n53448 & n10371;
  assign n10373 = n10293 & n10372;
  assign n10374 = n2537 & n10360;
  assign n10375 = n54340 & n10374;
  assign n10376 = n54339 & n10375;
  assign n10377 = n54338 & n10376;
  assign n10378 = n10373 & n10377;
  assign n10379 = n2537 & n4020;
  assign n10380 = n10369 & n10379;
  assign n10381 = n54230 & n10380;
  assign n10382 = n10295 & n10381;
  assign n10383 = n1035 & n10360;
  assign n10384 = n54339 & n10383;
  assign n10385 = n54340 & n10384;
  assign n10386 = n54338 & n10385;
  assign n10387 = n10382 & n10386;
  assign n10388 = n54334 & n10368;
  assign n10389 = n54294 & n54343;
  assign n10390 = n54230 & n54340;
  assign n10391 = n4020 & n10390;
  assign n10392 = n54333 & n10391;
  assign n10393 = n54294 & n10392;
  assign n10394 = n54338 & n10393;
  assign n10395 = n53448 & n10394;
  assign n10396 = n2537 & n10395;
  assign n10397 = n1067 & n10396;
  assign n10398 = n54331 & n10397;
  assign n10399 = n54339 & n10398;
  assign n10400 = n1035 & n10399;
  assign n10401 = ~n659 & n10400;
  assign n10402 = ~n404 & n10401;
  assign n10403 = ~n420 & n10402;
  assign n10404 = ~n450 & n10403;
  assign n10405 = n54331 & n10389;
  assign n10406 = ~n54305 & ~n54344;
  assign n10407 = ~n54325 & ~n54344;
  assign n10408 = n54305 & ~n54344;
  assign n10409 = ~n54325 & n10408;
  assign n10410 = n54305 & n10407;
  assign n10411 = ~n10406 & ~n54345;
  assign n10412 = ~n10226 & ~n54344;
  assign n10413 = n9968 & ~n54346;
  assign n10414 = ~n9966 & ~n10413;
  assign n10415 = n54269 & n54277;
  assign n10416 = ~n9692 & ~n10415;
  assign n10417 = ~n10414 & n10416;
  assign n10418 = ~n9692 & ~n10417;
  assign n10419 = n54254 & n54269;
  assign n10420 = ~n9587 & ~n10419;
  assign n10421 = ~n10418 & n10420;
  assign n10422 = ~n9587 & ~n10421;
  assign n10423 = n54240 & n54254;
  assign n10424 = ~n9394 & ~n10423;
  assign n10425 = ~n10422 & n10424;
  assign n10426 = ~n9394 & ~n10425;
  assign n10427 = n54212 & n54240;
  assign n10428 = ~n9148 & ~n10427;
  assign n10429 = ~n10426 & n10428;
  assign n10430 = ~n9148 & ~n10429;
  assign n10431 = n54194 & n54212;
  assign n10432 = ~n8858 & ~n10431;
  assign n10433 = ~n10430 & n10432;
  assign n10434 = ~n8858 & ~n10433;
  assign n10435 = n54183 & n54194;
  assign n10436 = ~n8631 & ~n10435;
  assign n10437 = ~n10434 & n10436;
  assign n10438 = ~n8631 & ~n10437;
  assign n10439 = n54163 & n54183;
  assign n10440 = ~n8530 & ~n10439;
  assign n10441 = ~n10438 & n10440;
  assign n10442 = ~n8530 & ~n10441;
  assign n10443 = n54154 & n54163;
  assign n10444 = ~n8264 & ~n10443;
  assign n10445 = ~n10442 & n10444;
  assign n10446 = ~n8264 & ~n10445;
  assign n10447 = n54132 & n54154;
  assign n10448 = ~n8088 & ~n10447;
  assign n10449 = ~n10446 & n10448;
  assign n10450 = ~n8088 & ~n10449;
  assign n10451 = n54119 & n54132;
  assign n10452 = ~n7845 & ~n10451;
  assign n10453 = ~n10450 & n10452;
  assign n10454 = ~n7845 & ~n10453;
  assign n10455 = n54098 & n54119;
  assign n10456 = ~n7754 & ~n10455;
  assign n10457 = ~n10454 & n10456;
  assign n10458 = ~n7754 & ~n10457;
  assign n10459 = n54073 & n54098;
  assign n10460 = ~n7470 & ~n10459;
  assign n10461 = ~n10458 & n10460;
  assign n10462 = ~n7470 & ~n10461;
  assign n10463 = n54050 & n54073;
  assign n10464 = ~n7200 & ~n10463;
  assign n10465 = ~n10462 & n10464;
  assign n10466 = ~n7200 & ~n10465;
  assign n10467 = n54034 & n54050;
  assign n10468 = ~n6929 & ~n10467;
  assign n10469 = ~n10466 & n10468;
  assign n10470 = ~n6929 & ~n10469;
  assign n10471 = n54005 & n54034;
  assign n10472 = ~n6794 & ~n10471;
  assign n10473 = ~n10470 & n10472;
  assign n10474 = ~n6794 & ~n10473;
  assign n10475 = n53970 & n54005;
  assign n10476 = ~n6529 & ~n10475;
  assign n10477 = ~n10474 & n10476;
  assign n10478 = ~n6529 & ~n10477;
  assign n10479 = n53962 & n53970;
  assign n10480 = ~n6149 & ~n10479;
  assign n10481 = ~n10478 & n10480;
  assign n10482 = ~n6149 & ~n10481;
  assign n10483 = n53930 & n53962;
  assign n10484 = ~n6052 & ~n10483;
  assign n10485 = ~n10482 & n10484;
  assign n10486 = ~n6052 & ~n10485;
  assign n10487 = n53907 & n53930;
  assign n10488 = ~n5732 & ~n10487;
  assign n10489 = ~n10486 & n10488;
  assign n10490 = ~n5732 & ~n10489;
  assign n10491 = n53888 & n53907;
  assign n10492 = ~n5440 & ~n10491;
  assign n10493 = ~n10490 & n10492;
  assign n10494 = ~n5440 & ~n10493;
  assign n10495 = n53860 & n53888;
  assign n10496 = ~n5255 & ~n10495;
  assign n10497 = ~n10494 & n10496;
  assign n10498 = ~n5255 & ~n10497;
  assign n10499 = n53845 & n53860;
  assign n10500 = ~n4951 & ~n10499;
  assign n10501 = ~n10498 & n10500;
  assign n10502 = ~n4951 & ~n10501;
  assign n10503 = n53819 & n53845;
  assign n10504 = ~n4785 & ~n10503;
  assign n10505 = ~n10502 & n10504;
  assign n10506 = ~n4785 & ~n10505;
  assign n10507 = n53799 & n53819;
  assign n10508 = ~n4456 & ~n10507;
  assign n10509 = ~n10506 & n10508;
  assign n10510 = ~n4456 & ~n10509;
  assign n10511 = n53774 & n53799;
  assign n10512 = ~n4196 & ~n10511;
  assign n10513 = ~n10510 & n10512;
  assign n10514 = ~n4196 & ~n10513;
  assign n10515 = n53741 & n53774;
  assign n10516 = ~n3876 & ~n10515;
  assign n10517 = ~n10514 & n10516;
  assign n10518 = ~n3876 & ~n10517;
  assign n10519 = n53712 & n53741;
  assign n10520 = ~n3521 & ~n10519;
  assign n10521 = ~n10518 & n10520;
  assign n10522 = ~n3521 & ~n10521;
  assign n10523 = n53685 & n53712;
  assign n10524 = ~n3213 & ~n10523;
  assign n10525 = ~n10522 & n10524;
  assign n10526 = ~n3213 & ~n10525;
  assign n10527 = n53657 & n53685;
  assign n10528 = ~n2891 & ~n10527;
  assign n10529 = ~n10526 & n10528;
  assign n10530 = ~n2891 & ~n10529;
  assign n10531 = n53650 & n53657;
  assign n10532 = ~n2626 & ~n10531;
  assign n10533 = ~n10530 & n10532;
  assign n10534 = ~n2626 & ~n10533;
  assign n10535 = n53634 & n53650;
  assign n10536 = ~n2536 & ~n10535;
  assign n10537 = ~n10534 & n10536;
  assign n10538 = ~n2536 & ~n10537;
  assign n10539 = ~n53565 & n53634;
  assign n10540 = n2325 & ~n53634;
  assign n10541 = ~n2325 & ~n53634;
  assign n10542 = n53565 & n53634;
  assign n10543 = n2325 & n53634;
  assign n10544 = ~n10541 & ~n54347;
  assign n10545 = ~n10539 & ~n10540;
  assign n10546 = ~n10538 & n54348;
  assign n10547 = n53634 & ~n10546;
  assign n10548 = ~n2325 & n10547;
  assign n10549 = n2325 & n10546;
  assign n10550 = ~n10538 & n10540;
  assign n10551 = ~n2325 & ~n10547;
  assign n10552 = ~n10541 & ~n10546;
  assign n10553 = n2325 & n10552;
  assign n10554 = n2325 & ~n10546;
  assign n10555 = ~n10551 & ~n54350;
  assign n10556 = ~n10548 & ~n54349;
  assign n10557 = n1576 & n54351;
  assign n10558 = pi30  & pi31 ;
  assign n10559 = ~pi30  & ~pi31 ;
  assign n10560 = pi30  & ~pi31 ;
  assign n10561 = ~pi30  & pi31 ;
  assign n10562 = ~n10560 & ~n10561;
  assign n10563 = ~n10558 & ~n10559;
  assign n10564 = n94 & ~n54352;
  assign n10565 = ~n2325 & n10564;
  assign n10566 = ~n10557 & ~n10565;
  assign n10567 = ~n1575 & ~n10566;
  assign n10568 = ~n1574 & n10566;
  assign n10569 = ~n1575 & ~n10568;
  assign n10570 = ~n1574 & ~n1575;
  assign n10571 = ~n10566 & n10570;
  assign n10572 = ~n1574 & ~n10571;
  assign n10573 = ~n1574 & ~n10567;
  assign n10574 = n877 & n54353;
  assign n10575 = ~n877 & ~n54353;
  assign n10576 = ~n10574 & ~n10575;
  assign n10577 = ~n465 & ~n1125;
  assign n10578 = ~n1485 & n10577;
  assign n10579 = n4319 & n5116;
  assign n10580 = n10578 & n10579;
  assign n10581 = ~n348 & ~n1031;
  assign n10582 = ~n623 & n10581;
  assign n10583 = ~n1031 & n8089;
  assign n10584 = ~n163 & ~n447;
  assign n10585 = ~n163 & ~n1644;
  assign n10586 = ~n447 & n10585;
  assign n10587 = ~n447 & ~n1644;
  assign n10588 = ~n163 & n10587;
  assign n10589 = ~n1644 & n10584;
  assign n10590 = n54354 & n54355;
  assign n10591 = n10580 & n10590;
  assign n10592 = n1458 & n4710;
  assign n10593 = ~n295 & ~n1476;
  assign n10594 = n915 & n10593;
  assign n10595 = n10592 & n10594;
  assign n10596 = n54168 & n10595;
  assign n10597 = n54228 & n10596;
  assign n10598 = ~n465 & ~n1476;
  assign n10599 = ~n1485 & n10598;
  assign n10600 = ~n295 & ~n1125;
  assign n10601 = n4319 & n10600;
  assign n10602 = n4319 & n10593;
  assign n10603 = n10578 & n10602;
  assign n10604 = n10599 & n10601;
  assign n10605 = n10590 & n54356;
  assign n10606 = n4710 & n5116;
  assign n10607 = n915 & n1458;
  assign n10608 = n915 & n5116;
  assign n10609 = n10592 & n10608;
  assign n10610 = n10606 & n10607;
  assign n10611 = n54168 & n54357;
  assign n10612 = n54228 & n10611;
  assign n10613 = n10605 & n10612;
  assign n10614 = n10591 & n10597;
  assign n10615 = n915 & n10590;
  assign n10616 = n54168 & n10615;
  assign n10617 = n54228 & n10616;
  assign n10618 = n54204 & n10617;
  assign n10619 = n5116 & n10618;
  assign n10620 = n4710 & n10619;
  assign n10621 = n4319 & n10620;
  assign n10622 = n1458 & n10621;
  assign n10623 = ~n1125 & n10622;
  assign n10624 = ~n295 & n10623;
  assign n10625 = ~n1485 & n10624;
  assign n10626 = ~n1476 & n10625;
  assign n10627 = ~n465 & n10626;
  assign n10628 = n54204 & n54358;
  assign n10629 = ~n553 & ~n776;
  assign n10630 = ~n553 & ~n1658;
  assign n10631 = ~n776 & n10630;
  assign n10632 = ~n776 & ~n1658;
  assign n10633 = ~n553 & n10632;
  assign n10634 = ~n1658 & n10629;
  assign n10635 = ~n349 & ~n832;
  assign n10636 = ~n1062 & ~n1337;
  assign n10637 = n10635 & n10636;
  assign n10638 = n53946 & n10637;
  assign n10639 = n54360 & n10638;
  assign n10640 = ~n218 & ~n296;
  assign n10641 = n5639 & n9631;
  assign n10642 = n10640 & n10641;
  assign n10643 = n358 & n561;
  assign n10644 = n1094 & n4002;
  assign n10645 = n10643 & n10644;
  assign n10646 = n10642 & n10645;
  assign n10647 = n53946 & n54360;
  assign n10648 = n1094 & n10647;
  assign n10649 = n4002 & n10648;
  assign n10650 = n358 & n10649;
  assign n10651 = n561 & n10650;
  assign n10652 = n5639 & n10651;
  assign n10653 = ~n296 & n10652;
  assign n10654 = ~n1062 & n10653;
  assign n10655 = ~n218 & n10654;
  assign n10656 = ~n1337 & n10655;
  assign n10657 = ~n832 & n10656;
  assign n10658 = ~n612 & n10657;
  assign n10659 = ~n349 & n10658;
  assign n10660 = ~n741 & n10659;
  assign n10661 = ~n296 & ~n1062;
  assign n10662 = n5790 & n10661;
  assign n10663 = n53946 & n10662;
  assign n10664 = n54360 & n10663;
  assign n10665 = n5639 & n10643;
  assign n10666 = ~n832 & ~n1337;
  assign n10667 = n9631 & n10666;
  assign n10668 = n10644 & n10667;
  assign n10669 = n10665 & n10668;
  assign n10670 = n10664 & n10669;
  assign n10671 = ~n296 & ~n612;
  assign n10672 = n10635 & n10671;
  assign n10673 = n53946 & n10672;
  assign n10674 = n54360 & n10673;
  assign n10675 = n1094 & n5639;
  assign n10676 = n561 & n10675;
  assign n10677 = ~n218 & ~n1062;
  assign n10678 = ~n741 & ~n1337;
  assign n10679 = n10677 & n10678;
  assign n10680 = n358 & n4002;
  assign n10681 = n10679 & n10680;
  assign n10682 = n10676 & n10681;
  assign n10683 = n10674 & n10682;
  assign n10684 = n10639 & n10646;
  assign n10685 = ~n748 & ~n824;
  assign n10686 = ~n630 & n10685;
  assign n10687 = ~n344 & ~n622;
  assign n10688 = ~n344 & ~n496;
  assign n10689 = ~n622 & n10688;
  assign n10690 = ~n496 & ~n622;
  assign n10691 = ~n344 & n10690;
  assign n10692 = ~n496 & n10687;
  assign n10693 = n2740 & n54362;
  assign n10694 = n10686 & n54362;
  assign n10695 = n2740 & n10694;
  assign n10696 = n10686 & n10693;
  assign n10697 = ~n319 & ~n565;
  assign n10698 = ~n460 & ~n742;
  assign n10699 = n10697 & n10698;
  assign n10700 = n755 & n4753;
  assign n10701 = n10699 & n10700;
  assign n10702 = ~n1059 & ~n1280;
  assign n10703 = ~n1061 & n10702;
  assign n10704 = n2339 & n10703;
  assign n10705 = n755 & n10697;
  assign n10706 = n4753 & n7131;
  assign n10707 = n10705 & n10706;
  assign n10708 = ~n742 & ~n1280;
  assign n10709 = ~n1061 & n10708;
  assign n10710 = n2339 & n10709;
  assign n10711 = n10707 & n10710;
  assign n10712 = n2338 & n4753;
  assign n10713 = n755 & n1682;
  assign n10714 = n2339 & n10700;
  assign n10715 = n10712 & n10713;
  assign n10716 = ~n460 & ~n1061;
  assign n10717 = ~n565 & n10716;
  assign n10718 = ~n319 & ~n1280;
  assign n10719 = ~n742 & ~n1059;
  assign n10720 = n10718 & n10719;
  assign n10721 = ~n319 & n10698;
  assign n10722 = ~n565 & ~n1280;
  assign n10723 = ~n1059 & ~n1061;
  assign n10724 = n10722 & n10723;
  assign n10725 = n10721 & n10724;
  assign n10726 = n10717 & n10720;
  assign n10727 = n54365 & n54366;
  assign n10728 = n10701 & n10704;
  assign n10729 = n54363 & n54364;
  assign n10730 = n1671 & n5154;
  assign n10731 = n5815 & n9260;
  assign n10732 = n10730 & n10731;
  assign n10733 = ~n255 & ~n568;
  assign n10734 = ~n255 & ~n1081;
  assign n10735 = ~n568 & n10734;
  assign n10736 = ~n1081 & n10733;
  assign n10737 = n1704 & n3801;
  assign n10738 = n54367 & n10737;
  assign n10739 = n1671 & n10737;
  assign n10740 = ~n1997 & n10739;
  assign n10741 = ~n1195 & n10740;
  assign n10742 = ~n1081 & n10741;
  assign n10743 = ~n311 & n10742;
  assign n10744 = ~n255 & n10743;
  assign n10745 = ~n568 & n10744;
  assign n10746 = ~n617 & n10745;
  assign n10747 = ~n420 & n10746;
  assign n10748 = ~n585 & n10747;
  assign n10749 = n1671 & n3801;
  assign n10750 = n10731 & n10749;
  assign n10751 = n1704 & n5154;
  assign n10752 = n54367 & n10751;
  assign n10753 = n10750 & n10752;
  assign n10754 = ~n568 & ~n617;
  assign n10755 = n1704 & n10754;
  assign n10756 = n10749 & n10755;
  assign n10757 = ~n420 & ~n1195;
  assign n10758 = ~n1081 & n10757;
  assign n10759 = ~n255 & ~n1997;
  assign n10760 = ~n311 & ~n585;
  assign n10761 = n10759 & n10760;
  assign n10762 = n10758 & n10761;
  assign n10763 = n10756 & n10762;
  assign n10764 = n10732 & n10738;
  assign n10765 = n53794 & n54368;
  assign n10766 = n10729 & n10765;
  assign n10767 = n54361 & n10766;
  assign n10768 = n1682 & n10693;
  assign n10769 = n4753 & n10768;
  assign n10770 = n53794 & n10769;
  assign n10771 = n54368 & n10770;
  assign n10772 = n54361 & n10771;
  assign n10773 = n10686 & n10772;
  assign n10774 = n54359 & n10773;
  assign n10775 = n2338 & n10774;
  assign n10776 = n755 & n10775;
  assign n10777 = ~n1061 & n10776;
  assign n10778 = ~n565 & n10777;
  assign n10779 = ~n1059 & n10778;
  assign n10780 = ~n1280 & n10779;
  assign n10781 = ~n742 & n10780;
  assign n10782 = ~n319 & n10781;
  assign n10783 = ~n460 & n10782;
  assign n10784 = n54359 & n10767;
  assign n10785 = n53537 & ~n54369;
  assign n10786 = ~n53537 & n54369;
  assign n10787 = ~n10785 & ~n10786;
  assign n10788 = ~n247 & ~n612;
  assign n10789 = ~n735 & n10788;
  assign n10790 = ~n788 & ~n1472;
  assign n10791 = ~n414 & ~n562;
  assign n10792 = n10790 & n10791;
  assign n10793 = n6223 & n7277;
  assign n10794 = ~n247 & ~n788;
  assign n10795 = ~n735 & n10794;
  assign n10796 = ~n414 & ~n612;
  assign n10797 = n7277 & n10796;
  assign n10798 = n10795 & n10797;
  assign n10799 = n10789 & n54370;
  assign n10800 = ~n163 & ~n1081;
  assign n10801 = ~n977 & ~n1081;
  assign n10802 = ~n163 & n10801;
  assign n10803 = ~n163 & ~n977;
  assign n10804 = ~n1081 & n10803;
  assign n10805 = ~n977 & n10800;
  assign n10806 = ~n771 & ~n914;
  assign n10807 = ~n914 & ~n1085;
  assign n10808 = ~n771 & n10807;
  assign n10809 = ~n771 & ~n1085;
  assign n10810 = ~n914 & n10809;
  assign n10811 = ~n1085 & n10806;
  assign n10812 = n54372 & n54373;
  assign n10813 = ~n414 & n10812;
  assign n10814 = ~n1472 & n10813;
  assign n10815 = ~n247 & n10814;
  assign n10816 = ~n562 & n10815;
  assign n10817 = ~n612 & n10816;
  assign n10818 = ~n788 & n10817;
  assign n10819 = ~n735 & n10818;
  assign n10820 = n54371 & n10812;
  assign n10821 = ~n1476 & ~n1490;
  assign n10822 = ~n1195 & ~n1490;
  assign n10823 = ~n1476 & n10822;
  assign n10824 = ~n1195 & n10821;
  assign n10825 = ~n348 & ~n504;
  assign n10826 = ~n1703 & n10825;
  assign n10827 = n4214 & n4319;
  assign n10828 = n10826 & n10827;
  assign n10829 = n54375 & n10828;
  assign n10830 = ~n560 & ~n1125;
  assign n10831 = ~n310 & ~n1468;
  assign n10832 = n10830 & n10831;
  assign n10833 = ~n1125 & n54362;
  assign n10834 = ~n1468 & n10833;
  assign n10835 = ~n310 & n10834;
  assign n10836 = ~n560 & n10835;
  assign n10837 = n54362 & n10832;
  assign n10838 = n6482 & n7648;
  assign n10839 = n7846 & n10031;
  assign n10840 = n10838 & n10839;
  assign n10841 = n54376 & n10840;
  assign n10842 = ~n504 & ~n1703;
  assign n10843 = ~n216 & n10842;
  assign n10844 = ~n168 & ~n348;
  assign n10845 = n4214 & n10844;
  assign n10846 = n10843 & n10845;
  assign n10847 = n54375 & n10846;
  assign n10848 = n6482 & n10031;
  assign n10849 = n4319 & n7846;
  assign n10850 = n10848 & n10849;
  assign n10851 = n54376 & n10850;
  assign n10852 = n10847 & n10851;
  assign n10853 = ~n499 & ~n1703;
  assign n10854 = ~n216 & n10853;
  assign n10855 = ~n307 & ~n348;
  assign n10856 = ~n168 & ~n504;
  assign n10857 = n10855 & n10856;
  assign n10858 = n10854 & n10857;
  assign n10859 = n54375 & n10858;
  assign n10860 = n4214 & n6482;
  assign n10861 = n4319 & n10031;
  assign n10862 = n10860 & n10861;
  assign n10863 = n54376 & n10862;
  assign n10864 = n10859 & n10863;
  assign n10865 = n10829 & n10841;
  assign n10866 = n54375 & n54376;
  assign n10867 = n54374 & n10866;
  assign n10868 = n6482 & n10867;
  assign n10869 = n4319 & n10868;
  assign n10870 = n4214 & n10869;
  assign n10871 = n10031 & n10870;
  assign n10872 = ~n1703 & n10871;
  assign n10873 = ~n168 & n10872;
  assign n10874 = ~n307 & n10873;
  assign n10875 = ~n216 & n10874;
  assign n10876 = ~n504 & n10875;
  assign n10877 = ~n499 & n10876;
  assign n10878 = ~n348 & n10877;
  assign n10879 = n54374 & n54377;
  assign n10880 = ~n174 & ~n317;
  assign n10881 = ~n364 & ~n503;
  assign n10882 = ~n174 & ~n503;
  assign n10883 = ~n317 & ~n364;
  assign n10884 = n10882 & n10883;
  assign n10885 = n10880 & n10881;
  assign n10886 = n3335 & n8539;
  assign n10887 = ~n291 & ~n1033;
  assign n10888 = ~n1487 & n10887;
  assign n10889 = ~n174 & n10888;
  assign n10890 = ~n317 & n10889;
  assign n10891 = ~n503 & n10890;
  assign n10892 = ~n364 & n10891;
  assign n10893 = ~n409 & n10892;
  assign n10894 = ~n291 & ~n317;
  assign n10895 = n8539 & n10894;
  assign n10896 = ~n174 & ~n409;
  assign n10897 = n10881 & n10896;
  assign n10898 = n10895 & n10897;
  assign n10899 = n54379 & n10886;
  assign n10900 = n4261 & n7788;
  assign n10901 = ~n255 & ~n1465;
  assign n10902 = n1955 & n10901;
  assign n10903 = n10900 & n10902;
  assign n10904 = n566 & n775;
  assign n10905 = n2454 & n3134;
  assign n10906 = n10904 & n10905;
  assign n10907 = n10903 & n10906;
  assign n10908 = n54380 & n10907;
  assign n10909 = n3650 & n7045;
  assign n10910 = ~n256 & ~n1535;
  assign n10911 = n10001 & n10910;
  assign n10912 = n10909 & n10911;
  assign n10913 = ~n311 & ~n618;
  assign n10914 = ~n833 & n10913;
  assign n10915 = n4502 & n10914;
  assign n10916 = n4501 & n7045;
  assign n10917 = ~n316 & n10916;
  assign n10918 = ~n184 & n10917;
  assign n10919 = ~n311 & n10918;
  assign n10920 = ~n256 & n10919;
  assign n10921 = ~n554 & n10920;
  assign n10922 = ~n1535 & n10921;
  assign n10923 = ~n618 & n10922;
  assign n10924 = ~n1042 & n10923;
  assign n10925 = ~n823 & n10924;
  assign n10926 = ~n833 & n10925;
  assign n10927 = n7045 & n10001;
  assign n10928 = n10910 & n10927;
  assign n10929 = ~n316 & ~n618;
  assign n10930 = ~n311 & ~n833;
  assign n10931 = n10929 & n10930;
  assign n10932 = n3650 & n4501;
  assign n10933 = n10931 & n10932;
  assign n10934 = n10928 & n10933;
  assign n10935 = n4501 & n10910;
  assign n10936 = n10001 & n10935;
  assign n10937 = n10909 & n10931;
  assign n10938 = n10936 & n10937;
  assign n10939 = ~n1042 & ~n1535;
  assign n10940 = n7045 & n10939;
  assign n10941 = n4501 & n10940;
  assign n10942 = ~n184 & ~n618;
  assign n10943 = n10001 & n10942;
  assign n10944 = ~n311 & ~n316;
  assign n10945 = ~n256 & ~n833;
  assign n10946 = n10944 & n10945;
  assign n10947 = n10943 & n10946;
  assign n10948 = n10941 & n10947;
  assign n10949 = n10912 & n10915;
  assign n10950 = n2340 & n3014;
  assign n10951 = ~n491 & ~n1192;
  assign n10952 = ~n419 & n10951;
  assign n10953 = ~n320 & ~n360;
  assign n10954 = ~n320 & ~n1881;
  assign n10955 = ~n360 & n10954;
  assign n10956 = ~n1881 & n10953;
  assign n10957 = n10952 & n54382;
  assign n10958 = n10950 & n10957;
  assign n10959 = n54381 & n10958;
  assign n10960 = n3134 & n4261;
  assign n10961 = n1955 & n2340;
  assign n10962 = n10960 & n10961;
  assign n10963 = n2454 & n3014;
  assign n10964 = n7788 & n10901;
  assign n10965 = n10963 & n10964;
  assign n10966 = n10962 & n10965;
  assign n10967 = n54380 & n10966;
  assign n10968 = n10904 & n54382;
  assign n10969 = n10952 & n10968;
  assign n10970 = n54381 & n10969;
  assign n10971 = n10967 & n10970;
  assign n10972 = n1955 & n3134;
  assign n10973 = n775 & n10901;
  assign n10974 = n10972 & n10973;
  assign n10975 = n2454 & n7788;
  assign n10976 = n8328 & n10975;
  assign n10977 = n10974 & n10976;
  assign n10978 = n54380 & n10977;
  assign n10979 = ~n565 & n10953;
  assign n10980 = ~n564 & ~n1881;
  assign n10981 = n3014 & n10980;
  assign n10982 = n10979 & n10981;
  assign n10983 = n10952 & n10982;
  assign n10984 = n54381 & n10983;
  assign n10985 = n10978 & n10984;
  assign n10986 = n10908 & n10959;
  assign n10987 = n54378 & n54383;
  assign n10988 = n3134 & n10952;
  assign n10989 = n7788 & n10988;
  assign n10990 = n54381 & n10989;
  assign n10991 = n54378 & n10990;
  assign n10992 = n54040 & n10991;
  assign n10993 = n1955 & n10992;
  assign n10994 = n2454 & n10993;
  assign n10995 = n775 & n10994;
  assign n10996 = n54380 & n10995;
  assign n10997 = n4261 & n10996;
  assign n10998 = n10901 & n10997;
  assign n10999 = n2340 & n10998;
  assign n11000 = n3014 & n10999;
  assign n11001 = ~n320 & n11000;
  assign n11002 = ~n565 & n11001;
  assign n11003 = ~n564 & n11002;
  assign n11004 = ~n360 & n11003;
  assign n11005 = ~n1881 & n11004;
  assign n11006 = n54040 & n10987;
  assign n11007 = ~n215 & ~n222;
  assign n11008 = ~n292 & ~n1090;
  assign n11009 = ~n222 & ~n292;
  assign n11010 = ~n215 & ~n1090;
  assign n11011 = n11009 & n11010;
  assign n11012 = n11007 & n11008;
  assign n11013 = n5539 & n6535;
  assign n11014 = n7130 & n11013;
  assign n11015 = n6535 & n7130;
  assign n11016 = ~n1090 & n11015;
  assign n11017 = ~n215 & n11016;
  assign n11018 = ~n292 & n11017;
  assign n11019 = ~n222 & n11018;
  assign n11020 = ~n440 & n11019;
  assign n11021 = ~n450 & n11020;
  assign n11022 = ~n215 & ~n292;
  assign n11023 = ~n222 & ~n440;
  assign n11024 = ~n292 & ~n440;
  assign n11025 = n11007 & n11024;
  assign n11026 = n11022 & n11023;
  assign n11027 = ~n450 & ~n1090;
  assign n11028 = n6535 & n11027;
  assign n11029 = n7130 & n11028;
  assign n11030 = n54387 & n11029;
  assign n11031 = n54385 & n11014;
  assign n11032 = ~n207 & ~n771;
  assign n11033 = ~n207 & ~n1997;
  assign n11034 = ~n771 & n11033;
  assign n11035 = ~n771 & ~n1997;
  assign n11036 = ~n207 & n11035;
  assign n11037 = ~n1997 & n11032;
  assign n11038 = n3476 & n4378;
  assign n11039 = n1489 & n11038;
  assign n11040 = n54388 & n11039;
  assign n11041 = n906 & n1536;
  assign n11042 = ~n562 & ~n663;
  assign n11043 = ~n354 & ~n553;
  assign n11044 = n11042 & n11043;
  assign n11045 = n11041 & n11044;
  assign n11046 = ~n754 & n1366;
  assign n11047 = n4026 & n4893;
  assign n11048 = n11046 & n11047;
  assign n11049 = n11045 & n11048;
  assign n11050 = ~n754 & ~n1485;
  assign n11051 = n1366 & n11050;
  assign n11052 = n1488 & n3476;
  assign n11053 = n11051 & n11052;
  assign n11054 = n54388 & n11053;
  assign n11055 = n906 & n4026;
  assign n11056 = n4378 & n11055;
  assign n11057 = n4893 & n11042;
  assign n11058 = n1536 & n11043;
  assign n11059 = n11057 & n11058;
  assign n11060 = n11042 & n11058;
  assign n11061 = n4026 & n4378;
  assign n11062 = n906 & n4893;
  assign n11063 = n11061 & n11062;
  assign n11064 = n11060 & n11063;
  assign n11065 = n11056 & n11059;
  assign n11066 = n11054 & n54389;
  assign n11067 = ~n754 & ~n922;
  assign n11068 = n11042 & n11067;
  assign n11069 = ~n1485 & ~n1535;
  assign n11070 = ~n911 & ~n1031;
  assign n11071 = n11069 & n11070;
  assign n11072 = n11068 & n11071;
  assign n11073 = n54388 & n11072;
  assign n11074 = n906 & n3476;
  assign n11075 = n11043 & n11074;
  assign n11076 = n1488 & n4893;
  assign n11077 = n11061 & n11076;
  assign n11078 = n11075 & n11077;
  assign n11079 = n11073 & n11078;
  assign n11080 = n11040 & n11049;
  assign n11081 = n4893 & n54388;
  assign n11082 = n11043 & n11081;
  assign n11083 = n54386 & n11082;
  assign n11084 = n1488 & n11083;
  assign n11085 = n3476 & n11084;
  assign n11086 = n4378 & n11085;
  assign n11087 = n4026 & n11086;
  assign n11088 = n906 & n11087;
  assign n11089 = ~n1031 & n11088;
  assign n11090 = ~n922 & n11089;
  assign n11091 = ~n1485 & n11090;
  assign n11092 = ~n562 & n11091;
  assign n11093 = ~n663 & n11092;
  assign n11094 = ~n1535 & n11093;
  assign n11095 = ~n911 & n11094;
  assign n11096 = ~n754 & n11095;
  assign n11097 = n54386 & n54390;
  assign n11098 = ~n513 & n1578;
  assign n11099 = ~n246 & ~n1658;
  assign n11100 = ~n246 & n1578;
  assign n11101 = ~n1658 & n11100;
  assign n11102 = ~n513 & n11101;
  assign n11103 = ~n513 & ~n1658;
  assign n11104 = ~n246 & n11103;
  assign n11105 = n1578 & n11104;
  assign n11106 = n11098 & n11099;
  assign n11107 = ~n172 & ~n504;
  assign n11108 = ~n774 & n11107;
  assign n11109 = n3217 & n11108;
  assign n11110 = ~n310 & ~n588;
  assign n11111 = ~n612 & ~n822;
  assign n11112 = ~n310 & ~n822;
  assign n11113 = ~n612 & n11112;
  assign n11114 = ~n588 & n11113;
  assign n11115 = n11110 & n11111;
  assign n11116 = n4503 & n54393;
  assign n11117 = ~n590 & ~n774;
  assign n11118 = n11107 & n11117;
  assign n11119 = n3217 & n3742;
  assign n11120 = n11118 & n11119;
  assign n11121 = n54393 & n11120;
  assign n11122 = n11109 & n11116;
  assign n11123 = n54392 & n54393;
  assign n11124 = n3217 & n11123;
  assign n11125 = n3742 & n11124;
  assign n11126 = ~n172 & n11125;
  assign n11127 = ~n504 & n11126;
  assign n11128 = ~n774 & n11127;
  assign n11129 = ~n590 & n11128;
  assign n11130 = n54392 & n54394;
  assign n11131 = n3389 & n3878;
  assign n11132 = n3214 & n4381;
  assign n11133 = n11131 & n11132;
  assign n11134 = ~n564 & ~n753;
  assign n11135 = ~n498 & ~n1065;
  assign n11136 = ~n1065 & n11134;
  assign n11137 = ~n498 & n11136;
  assign n11138 = n11134 & n11135;
  assign n11139 = ~n567 & ~n830;
  assign n11140 = ~n824 & ~n1192;
  assign n11141 = ~n567 & ~n824;
  assign n11142 = ~n830 & ~n1192;
  assign n11143 = n11141 & n11142;
  assign n11144 = n11139 & n11140;
  assign n11145 = n54396 & n54397;
  assign n11146 = n11133 & n11145;
  assign n11147 = ~n356 & ~n625;
  assign n11148 = ~n625 & ~n770;
  assign n11149 = ~n356 & n11148;
  assign n11150 = ~n770 & n11147;
  assign n11151 = ~n356 & n2367;
  assign n11152 = ~n770 & n11151;
  assign n11153 = ~n625 & n11152;
  assign n11154 = n2367 & n54398;
  assign n11155 = ~n511 & ~n617;
  assign n11156 = n6860 & n9337;
  assign n11157 = n11155 & n11156;
  assign n11158 = n54399 & n11157;
  assign n11159 = n3214 & n6860;
  assign n11160 = n3878 & n4381;
  assign n11161 = n11159 & n11160;
  assign n11162 = n3389 & n11142;
  assign n11163 = n54396 & n11162;
  assign n11164 = n11161 & n11163;
  assign n11165 = n9337 & n11155;
  assign n11166 = n11141 & n11165;
  assign n11167 = n54399 & n11166;
  assign n11168 = n11164 & n11167;
  assign n11169 = n11141 & n11155;
  assign n11170 = n11156 & n11169;
  assign n11171 = n3214 & n11142;
  assign n11172 = n54396 & n11171;
  assign n11173 = n11170 & n11172;
  assign n11174 = n3389 & n4381;
  assign n11175 = n3878 & n11174;
  assign n11176 = n54399 & n11175;
  assign n11177 = n11173 & n11176;
  assign n11178 = n3878 & n9337;
  assign n11179 = n11174 & n11178;
  assign n11180 = n11145 & n11179;
  assign n11181 = n11155 & n11159;
  assign n11182 = n54399 & n11181;
  assign n11183 = n11180 & n11182;
  assign n11184 = n11146 & n11158;
  assign n11185 = n54395 & n54400;
  assign n11186 = n54318 & n11185;
  assign n11187 = n54396 & n11155;
  assign n11188 = n6860 & n11187;
  assign n11189 = n54399 & n11188;
  assign n11190 = n54318 & n11189;
  assign n11191 = n54391 & n11190;
  assign n11192 = n54395 & n11191;
  assign n11193 = n3878 & n11192;
  assign n11194 = n3214 & n11193;
  assign n11195 = n9337 & n11194;
  assign n11196 = n3389 & n11195;
  assign n11197 = n4381 & n11196;
  assign n11198 = ~n1192 & n11197;
  assign n11199 = ~n567 & n11198;
  assign n11200 = ~n824 & n11199;
  assign n11201 = ~n830 & n11200;
  assign n11202 = n54391 & n11186;
  assign n11203 = ~n54384 & ~n54401;
  assign n11204 = n54384 & n54401;
  assign n11205 = ~pi26  & ~n11203;
  assign n11206 = ~n11203 & ~n11204;
  assign n11207 = ~pi26  & n11206;
  assign n11208 = ~n11204 & n11205;
  assign n11209 = ~n11203 & ~n54402;
  assign n11210 = n54369 & ~n11209;
  assign n11211 = ~n54369 & n11209;
  assign n11212 = n10530 & ~n10532;
  assign n11213 = ~n10533 & ~n11212;
  assign n11214 = n1576 & n11213;
  assign n11215 = ~pi31  & ~n94;
  assign n11216 = ~n53650 & n11215;
  assign n11217 = n94 & n10558;
  assign n11218 = pi31  & n53443;
  assign n11219 = ~n53685 & n54403;
  assign n11220 = ~n53657 & n10564;
  assign n11221 = ~n11219 & ~n11220;
  assign n11222 = ~n11216 & n11221;
  assign n11223 = ~n11214 & n11222;
  assign n11224 = ~n11211 & ~n11223;
  assign n11225 = ~n11210 & n11223;
  assign n11226 = ~n11211 & ~n11225;
  assign n11227 = ~n11210 & ~n11211;
  assign n11228 = ~n11223 & n11227;
  assign n11229 = ~n11210 & ~n11228;
  assign n11230 = ~n11210 & ~n11224;
  assign n11231 = ~n10785 & n54404;
  assign n11232 = ~n10786 & n11231;
  assign n11233 = n10787 & n54404;
  assign n11234 = ~n10785 & ~n54405;
  assign n11235 = ~pi29  & ~n53560;
  assign n11236 = ~n1568 & n1573;
  assign n11237 = ~n11235 & ~n11236;
  assign n11238 = ~n11234 & ~n11237;
  assign n11239 = n11234 & n11237;
  assign n11240 = ~n11238 & ~n11239;
  assign n11241 = n10538 & ~n54348;
  assign n11242 = ~n10546 & ~n11241;
  assign n11243 = n1576 & n11242;
  assign n11244 = ~n53650 & n54403;
  assign n11245 = ~n53634 & n10564;
  assign n11246 = ~n11244 & ~n11245;
  assign n11247 = ~n11243 & n11246;
  assign n11248 = n11240 & ~n11247;
  assign n11249 = ~n11238 & ~n11248;
  assign n11250 = n10566 & ~n10570;
  assign n11251 = ~n10566 & ~n10571;
  assign n11252 = n10570 & ~n10571;
  assign n11253 = ~n11251 & ~n11252;
  assign n11254 = ~n10571 & ~n11250;
  assign n11255 = ~n11249 & ~n54406;
  assign n11256 = n11249 & n54406;
  assign n11257 = ~n11255 & ~n11256;
  assign n11258 = ~n11240 & n11247;
  assign n11259 = ~n11248 & ~n11258;
  assign n11260 = ~n209 & ~n289;
  assign n11261 = pi26  & ~pi27 ;
  assign n11262 = ~pi26  & pi27 ;
  assign n11263 = ~pi26  & ~pi27 ;
  assign n11264 = pi26  & pi27 ;
  assign n11265 = ~n11263 & ~n11264;
  assign n11266 = ~n11261 & ~n11262;
  assign n11267 = n11260 & ~n54407;
  assign n11268 = ~n54407 & ~n11267;
  assign n11269 = ~n11260 & ~n54407;
  assign n11270 = pi28  & ~pi29 ;
  assign n11271 = ~pi28  & pi29 ;
  assign n11272 = ~pi28  & ~pi29 ;
  assign n11273 = pi28  & pi29 ;
  assign n11274 = ~n11272 & ~n11273;
  assign n11275 = ~n11270 & ~n11271;
  assign n11276 = ~n54407 & n54409;
  assign n11277 = ~n11260 & n11276;
  assign n11278 = n54408 & n54409;
  assign n11279 = n54407 & n54409;
  assign n11280 = ~n10547 & n11279;
  assign n11281 = ~n54410 & ~n11280;
  assign n11282 = ~n2325 & ~n11281;
  assign n11283 = ~n2325 & n54410;
  assign n11284 = ~pi29  & ~n54411;
  assign n11285 = n10534 & ~n10536;
  assign n11286 = ~n10537 & ~n11285;
  assign n11287 = n1576 & n11286;
  assign n11288 = ~n53650 & n10564;
  assign n11289 = ~n53657 & n54403;
  assign n11290 = ~n53634 & n11215;
  assign n11291 = ~n11289 & ~n11290;
  assign n11292 = ~n11288 & ~n11289;
  assign n11293 = ~n11290 & n11292;
  assign n11294 = ~n11288 & n11291;
  assign n11295 = ~n11287 & n54412;
  assign n11296 = n11284 & n11295;
  assign n11297 = ~n11284 & ~n11295;
  assign n11298 = ~n10787 & ~n54404;
  assign n11299 = n54404 & ~n54405;
  assign n11300 = ~n10786 & n11234;
  assign n11301 = ~n11299 & ~n11300;
  assign n11302 = ~n54405 & ~n11298;
  assign n11303 = ~n11297 & n54413;
  assign n11304 = ~n11284 & ~n11297;
  assign n11305 = ~n11295 & ~n11297;
  assign n11306 = ~n11304 & ~n11305;
  assign n11307 = ~n11296 & ~n11297;
  assign n11308 = ~n54413 & ~n54414;
  assign n11309 = ~n11297 & ~n11308;
  assign n11310 = ~n11296 & ~n11303;
  assign n11311 = n11259 & ~n54415;
  assign n11312 = n1273 & n7276;
  assign n11313 = n1653 & n11043;
  assign n11314 = n1273 & n1653;
  assign n11315 = n7276 & n11043;
  assign n11316 = n11314 & n11315;
  assign n11317 = n11312 & n11313;
  assign n11318 = ~n179 & ~n271;
  assign n11319 = ~n179 & ~n363;
  assign n11320 = ~n271 & n11319;
  assign n11321 = ~n271 & ~n363;
  assign n11322 = ~n179 & n11321;
  assign n11323 = ~n363 & n11318;
  assign n11324 = ~n651 & ~n1658;
  assign n11325 = ~n975 & ~n983;
  assign n11326 = ~n975 & ~n1658;
  assign n11327 = ~n651 & ~n983;
  assign n11328 = n11326 & n11327;
  assign n11329 = ~n651 & ~n975;
  assign n11330 = ~n983 & ~n1658;
  assign n11331 = n11329 & n11330;
  assign n11332 = n11324 & n11325;
  assign n11333 = n5984 & n54418;
  assign n11334 = n54417 & n11333;
  assign n11335 = n1653 & n7276;
  assign n11336 = n5984 & n11335;
  assign n11337 = n1273 & n11043;
  assign n11338 = n54418 & n11337;
  assign n11339 = n54417 & n11338;
  assign n11340 = n11336 & n11339;
  assign n11341 = n54416 & n11334;
  assign n11342 = n53579 & n54419;
  assign n11343 = n1653 & n54417;
  assign n11344 = n11043 & n11343;
  assign n11345 = n53617 & n11344;
  assign n11346 = n53579 & n11345;
  assign n11347 = n1273 & n11346;
  assign n11348 = n2476 & n11347;
  assign n11349 = n7276 & n11348;
  assign n11350 = n3672 & n11349;
  assign n11351 = ~n983 & n11350;
  assign n11352 = ~n975 & n11351;
  assign n11353 = ~n1658 & n11352;
  assign n11354 = ~n651 & n11353;
  assign n11355 = n53617 & n11342;
  assign n11356 = n54384 & ~n54420;
  assign n11357 = ~n54384 & n54420;
  assign n11358 = ~n11356 & ~n11357;
  assign n11359 = n10522 & ~n10524;
  assign n11360 = ~n10525 & ~n11359;
  assign n11361 = n1576 & n11360;
  assign n11362 = ~n53685 & n11215;
  assign n11363 = ~n53741 & n54403;
  assign n11364 = ~n53712 & n10564;
  assign n11365 = ~n11363 & ~n11364;
  assign n11366 = ~n11362 & ~n11363;
  assign n11367 = ~n11364 & n11366;
  assign n11368 = ~n11362 & n11365;
  assign n11369 = ~n11361 & n54421;
  assign n11370 = ~n11356 & ~n11369;
  assign n11371 = ~n11357 & n11370;
  assign n11372 = n11358 & ~n11369;
  assign n11373 = ~n11356 & ~n54422;
  assign n11374 = ~pi26  & ~n54402;
  assign n11375 = ~n11204 & n11209;
  assign n11376 = ~n11374 & ~n11375;
  assign n11377 = ~n11373 & ~n11376;
  assign n11378 = n11373 & n11376;
  assign n11379 = n10526 & ~n10528;
  assign n11380 = ~n10529 & ~n11379;
  assign n11381 = n1576 & n11380;
  assign n11382 = ~n53685 & n10564;
  assign n11383 = ~n53657 & n11215;
  assign n11384 = ~n53712 & n54403;
  assign n11385 = ~n11383 & ~n11384;
  assign n11386 = ~n11382 & ~n11384;
  assign n11387 = ~n11383 & n11386;
  assign n11388 = ~n11382 & n11385;
  assign n11389 = ~n11381 & n54423;
  assign n11390 = ~n11378 & ~n11389;
  assign n11391 = ~n11377 & ~n11378;
  assign n11392 = ~n11389 & n11391;
  assign n11393 = ~n11377 & ~n11392;
  assign n11394 = ~n11377 & ~n11390;
  assign n11395 = n11223 & ~n11227;
  assign n11396 = ~n11223 & ~n11228;
  assign n11397 = n11227 & ~n11228;
  assign n11398 = ~n11396 & ~n11397;
  assign n11399 = ~n11228 & ~n11395;
  assign n11400 = ~n54424 & ~n54425;
  assign n11401 = n54424 & n54425;
  assign n11402 = n54351 & n11279;
  assign n11403 = ~n53634 & n54410;
  assign n11404 = ~n2325 & n11267;
  assign n11405 = ~n11403 & ~n11404;
  assign n11406 = ~n11402 & n11405;
  assign n11407 = pi29  & ~n11406;
  assign n11408 = pi29  & ~n11407;
  assign n11409 = pi29  & n11406;
  assign n11410 = ~n11406 & ~n11407;
  assign n11411 = ~pi29  & ~n11406;
  assign n11412 = ~n54426 & ~n54427;
  assign n11413 = ~n11401 & ~n11412;
  assign n11414 = ~n11400 & ~n11401;
  assign n11415 = ~n11412 & n11414;
  assign n11416 = ~n11400 & ~n11415;
  assign n11417 = ~n11400 & ~n11413;
  assign n11418 = n54413 & ~n54414;
  assign n11419 = ~n54413 & n54414;
  assign n11420 = ~n11418 & ~n11419;
  assign n11421 = ~n54428 & ~n11420;
  assign n11422 = ~n11358 & n11369;
  assign n11423 = ~n11369 & ~n54422;
  assign n11424 = ~n11357 & n11373;
  assign n11425 = ~n11423 & ~n11424;
  assign n11426 = ~n54422 & ~n11422;
  assign n11427 = ~n321 & ~n1192;
  assign n11428 = ~n221 & ~n514;
  assign n11429 = n7604 & n11428;
  assign n11430 = n11427 & n11429;
  assign n11431 = ~n275 & ~n552;
  assign n11432 = ~n1715 & n11431;
  assign n11433 = n3218 & n3932;
  assign n11434 = n11432 & n11433;
  assign n11435 = n53760 & n54021;
  assign n11436 = n11434 & n11435;
  assign n11437 = n3932 & n54021;
  assign n11438 = n53760 & n11437;
  assign n11439 = n11428 & n11438;
  assign n11440 = ~n896 & n11439;
  assign n11441 = ~n1192 & n11440;
  assign n11442 = ~n1196 & n11441;
  assign n11443 = ~n321 & n11442;
  assign n11444 = ~n660 & n11443;
  assign n11445 = ~n552 & n11444;
  assign n11446 = ~n275 & n11445;
  assign n11447 = ~n741 & n11446;
  assign n11448 = ~n1715 & n11447;
  assign n11449 = n3932 & n11427;
  assign n11450 = n11428 & n11449;
  assign n11451 = ~n275 & ~n1196;
  assign n11452 = ~n552 & n11451;
  assign n11453 = ~n660 & ~n1715;
  assign n11454 = n3218 & n11453;
  assign n11455 = n11452 & n11454;
  assign n11456 = n11435 & n11455;
  assign n11457 = n11450 & n11456;
  assign n11458 = ~n552 & ~n1715;
  assign n11459 = n3932 & n11458;
  assign n11460 = n11428 & n11459;
  assign n11461 = ~n321 & ~n660;
  assign n11462 = ~n275 & n11461;
  assign n11463 = ~n1192 & ~n1196;
  assign n11464 = n3218 & n11463;
  assign n11465 = n11462 & n11464;
  assign n11466 = n11435 & n11465;
  assign n11467 = n11460 & n11466;
  assign n11468 = n11430 & n11436;
  assign n11469 = ~n585 & ~n615;
  assign n11470 = n4313 & n11469;
  assign n11471 = n7602 & n11470;
  assign n11472 = ~n659 & n755;
  assign n11473 = ~n832 & ~n1042;
  assign n11474 = ~n1641 & n11473;
  assign n11475 = n11472 & n11474;
  assign n11476 = n4313 & n11473;
  assign n11477 = n7602 & n11476;
  assign n11478 = ~n1641 & n11469;
  assign n11479 = n11472 & n11478;
  assign n11480 = n11477 & n11479;
  assign n11481 = ~n615 & ~n1641;
  assign n11482 = n7602 & n11481;
  assign n11483 = n4313 & n11482;
  assign n11484 = ~n585 & n11473;
  assign n11485 = n11472 & n11484;
  assign n11486 = n11483 & n11485;
  assign n11487 = n11471 & n11475;
  assign n11488 = n54299 & n54431;
  assign n11489 = ~n177 & ~n219;
  assign n11490 = ~n184 & ~n1646;
  assign n11491 = n11489 & n11490;
  assign n11492 = ~n255 & ~n1468;
  assign n11493 = n3676 & n6395;
  assign n11494 = n11492 & n11493;
  assign n11495 = ~n422 & n3676;
  assign n11496 = ~n1468 & n11495;
  assign n11497 = ~n184 & n11496;
  assign n11498 = ~n177 & n11497;
  assign n11499 = ~n219 & n11498;
  assign n11500 = ~n255 & n11499;
  assign n11501 = ~n1646 & n11500;
  assign n11502 = ~n448 & n11501;
  assign n11503 = ~n177 & ~n184;
  assign n11504 = n11492 & n11503;
  assign n11505 = ~n219 & ~n1646;
  assign n11506 = n6395 & n11505;
  assign n11507 = n3676 & n11506;
  assign n11508 = n11504 & n11507;
  assign n11509 = n11491 & n11494;
  assign n11510 = ~n559 & ~n833;
  assign n11511 = ~n833 & ~n879;
  assign n11512 = ~n559 & n11511;
  assign n11513 = ~n879 & n11510;
  assign n11514 = ~n789 & ~n2103;
  assign n11515 = n421 & n11155;
  assign n11516 = n11514 & n11515;
  assign n11517 = ~n2103 & n11515;
  assign n11518 = ~n879 & n11517;
  assign n11519 = ~n559 & n11518;
  assign n11520 = ~n833 & n11519;
  assign n11521 = ~n789 & n11520;
  assign n11522 = ~n789 & ~n833;
  assign n11523 = ~n2103 & n11522;
  assign n11524 = ~n559 & ~n879;
  assign n11525 = n421 & n11524;
  assign n11526 = n11155 & n11525;
  assign n11527 = n11523 & n11526;
  assign n11528 = n54433 & n11516;
  assign n11529 = n54432 & n54434;
  assign n11530 = n11488 & n11529;
  assign n11531 = n54430 & n54434;
  assign n11532 = n54299 & n11531;
  assign n11533 = n54432 & n11532;
  assign n11534 = n4313 & n11533;
  assign n11535 = ~n1125 & n11534;
  assign n11536 = n11472 & n11535;
  assign n11537 = ~n1042 & n11536;
  assign n11538 = ~n459 & n11537;
  assign n11539 = ~n832 & n11538;
  assign n11540 = ~n1641 & n11539;
  assign n11541 = ~n615 & n11540;
  assign n11542 = ~n585 & n11541;
  assign n11543 = n54430 & n11530;
  assign n11544 = ~n161 & ~n363;
  assign n11545 = ~n881 & n11544;
  assign n11546 = ~n416 & ~n554;
  assign n11547 = ~n310 & ~n510;
  assign n11548 = n11546 & n11547;
  assign n11549 = ~n416 & ~n881;
  assign n11550 = ~n310 & n11549;
  assign n11551 = ~n161 & n11550;
  assign n11552 = ~n554 & n11551;
  assign n11553 = ~n510 & n11552;
  assign n11554 = ~n363 & n11553;
  assign n11555 = ~n310 & ~n363;
  assign n11556 = ~n554 & n11555;
  assign n11557 = ~n416 & ~n510;
  assign n11558 = ~n161 & ~n881;
  assign n11559 = n11557 & n11558;
  assign n11560 = n11556 & n11559;
  assign n11561 = n11545 & n11548;
  assign n11562 = ~n513 & ~n647;
  assign n11563 = ~n742 & ~n2109;
  assign n11564 = ~n742 & ~n1491;
  assign n11565 = ~n2109 & n11564;
  assign n11566 = ~n1491 & n11563;
  assign n11567 = ~n513 & n11564;
  assign n11568 = ~n647 & n11567;
  assign n11569 = ~n2109 & n11568;
  assign n11570 = n11562 & n54437;
  assign n11571 = n906 & n964;
  assign n11572 = n8052 & n11571;
  assign n11573 = n54438 & n11572;
  assign n11574 = n54436 & n11573;
  assign n11575 = ~n402 & ~n1658;
  assign n11576 = ~n894 & ~n1195;
  assign n11577 = n11575 & n11576;
  assign n11578 = ~n291 & ~n294;
  assign n11579 = n1541 & n11578;
  assign n11580 = n11577 & n11579;
  assign n11581 = ~n450 & ~n499;
  assign n11582 = ~n499 & n1803;
  assign n11583 = ~n450 & n11582;
  assign n11584 = n1803 & n11581;
  assign n11585 = n9184 & n54439;
  assign n11586 = n11580 & n11585;
  assign n11587 = n53991 & n11586;
  assign n11588 = n906 & n1541;
  assign n11589 = n8052 & n11588;
  assign n11590 = n54436 & n11589;
  assign n11591 = n54438 & n11589;
  assign n11592 = n54436 & n11591;
  assign n11593 = n54438 & n11590;
  assign n11594 = ~n291 & ~n1195;
  assign n11595 = n11575 & n11594;
  assign n11596 = ~n294 & ~n894;
  assign n11597 = n964 & n11596;
  assign n11598 = ~n294 & ~n1658;
  assign n11599 = ~n291 & ~n402;
  assign n11600 = n11598 & n11599;
  assign n11601 = n964 & n11576;
  assign n11602 = n11600 & n11601;
  assign n11603 = n11595 & n11597;
  assign n11604 = n11585 & n54441;
  assign n11605 = n53991 & n11604;
  assign n11606 = n54440 & n11605;
  assign n11607 = n11574 & n11587;
  assign n11608 = n964 & n11585;
  assign n11609 = n54438 & n11608;
  assign n11610 = n53991 & n11609;
  assign n11611 = n54436 & n11610;
  assign n11612 = n54435 & n11611;
  assign n11613 = n8052 & n11612;
  assign n11614 = n1541 & n11613;
  assign n11615 = n906 & n11614;
  assign n11616 = ~n291 & n11615;
  assign n11617 = ~n894 & n11616;
  assign n11618 = ~n1195 & n11617;
  assign n11619 = ~n294 & n11618;
  assign n11620 = ~n402 & n11619;
  assign n11621 = ~n1658 & n11620;
  assign n11622 = n54435 & n54442;
  assign n11623 = ~n498 & ~n1641;
  assign n11624 = ~n498 & ~n1455;
  assign n11625 = ~n1641 & n11624;
  assign n11626 = ~n1455 & n11623;
  assign n11627 = n54375 & n54444;
  assign n11628 = ~n409 & ~n2109;
  assign n11629 = ~n451 & ~n466;
  assign n11630 = ~n409 & ~n466;
  assign n11631 = ~n451 & n11630;
  assign n11632 = ~n2109 & n11631;
  assign n11633 = ~n451 & ~n2109;
  assign n11634 = n11630 & n11633;
  assign n11635 = ~n409 & ~n451;
  assign n11636 = ~n466 & ~n2109;
  assign n11637 = n11635 & n11636;
  assign n11638 = n11628 & n11629;
  assign n11639 = ~n559 & ~n590;
  assign n11640 = ~n319 & ~n590;
  assign n11641 = ~n559 & n11640;
  assign n11642 = ~n319 & ~n559;
  assign n11643 = ~n590 & n11642;
  assign n11644 = ~n319 & n11639;
  assign n11645 = n54445 & n54446;
  assign n11646 = n11627 & n11645;
  assign n11647 = n2975 & n4501;
  assign n11648 = n1082 & n11647;
  assign n11649 = n293 & n417;
  assign n11650 = n1277 & n1336;
  assign n11651 = n11649 & n11650;
  assign n11652 = n1277 & n2975;
  assign n11653 = n1082 & n11652;
  assign n11654 = n417 & n4501;
  assign n11655 = n293 & n1336;
  assign n11656 = n11654 & n11655;
  assign n11657 = n11653 & n11656;
  assign n11658 = n11648 & n11651;
  assign n11659 = n53738 & n54447;
  assign n11660 = n54375 & n54446;
  assign n11661 = n1082 & n11660;
  assign n11662 = n4501 & n11661;
  assign n11663 = n54445 & n11662;
  assign n11664 = n417 & n11663;
  assign n11665 = n2975 & n11664;
  assign n11666 = n53738 & n11665;
  assign n11667 = n1277 & n11666;
  assign n11668 = n293 & n11667;
  assign n11669 = ~n1455 & n11668;
  assign n11670 = ~n1641 & n11669;
  assign n11671 = ~n503 & n11670;
  assign n11672 = ~n498 & n11671;
  assign n11673 = ~n773 & n11672;
  assign n11674 = ~n503 & ~n1455;
  assign n11675 = ~n498 & n11674;
  assign n11676 = n54446 & n11675;
  assign n11677 = n54375 & n54445;
  assign n11678 = n11676 & n11677;
  assign n11679 = n293 & n1277;
  assign n11680 = n417 & n11679;
  assign n11681 = ~n773 & ~n1641;
  assign n11682 = n2975 & n11681;
  assign n11683 = n1082 & n4501;
  assign n11684 = n11682 & n11683;
  assign n11685 = n11680 & n11684;
  assign n11686 = n53738 & n11685;
  assign n11687 = n11678 & n11686;
  assign n11688 = n11646 & n11659;
  assign n11689 = n1458 & n6150;
  assign n11690 = n7130 & n8091;
  assign n11691 = n11689 & n11690;
  assign n11692 = n53785 & n11691;
  assign n11693 = ~n163 & ~n1033;
  assign n11694 = n251 & n11693;
  assign n11695 = n712 & n5956;
  assign n11696 = ~n1033 & n11695;
  assign n11697 = ~n163 & n11696;
  assign n11698 = ~n250 & n11697;
  assign n11699 = ~n249 & n11698;
  assign n11700 = n712 & n11693;
  assign n11701 = n251 & n5956;
  assign n11702 = n11700 & n11701;
  assign n11703 = n11694 & n11695;
  assign n11704 = n54392 & n54449;
  assign n11705 = n11692 & n11704;
  assign n11706 = ~n957 & ~n1471;
  assign n11707 = ~n894 & ~n957;
  assign n11708 = ~n1471 & n11707;
  assign n11709 = ~n894 & n11706;
  assign n11710 = ~n344 & ~n848;
  assign n11711 = n4213 & n11710;
  assign n11712 = n1078 & n5060;
  assign n11713 = n11711 & n11712;
  assign n11714 = n54450 & n11713;
  assign n11715 = n53587 & n11714;
  assign n11716 = n7130 & n54392;
  assign n11717 = n54449 & n11716;
  assign n11718 = n53587 & n11717;
  assign n11719 = n53785 & n11718;
  assign n11720 = n5060 & n11719;
  assign n11721 = n1078 & n11720;
  assign n11722 = n6150 & n11721;
  assign n11723 = n8091 & n11722;
  assign n11724 = n1458 & n11723;
  assign n11725 = ~n1471 & n11724;
  assign n11726 = ~n894 & n11725;
  assign n11727 = ~n957 & n11726;
  assign n11728 = ~n568 & n11727;
  assign n11729 = ~n848 & n11728;
  assign n11730 = ~n344 & n11729;
  assign n11731 = ~n448 & n11730;
  assign n11732 = n1078 & n8091;
  assign n11733 = n4213 & n5060;
  assign n11734 = n11732 & n11733;
  assign n11735 = n54392 & n11734;
  assign n11736 = n53785 & n54449;
  assign n11737 = n11735 & n11736;
  assign n11738 = ~n344 & ~n957;
  assign n11739 = ~n848 & n11738;
  assign n11740 = ~n894 & ~n1471;
  assign n11741 = n6150 & n11740;
  assign n11742 = n1458 & n7130;
  assign n11743 = n11741 & n11742;
  assign n11744 = n11739 & n11743;
  assign n11745 = n53587 & n11744;
  assign n11746 = n11737 & n11745;
  assign n11747 = n1458 & n5060;
  assign n11748 = n6150 & n7130;
  assign n11749 = n11747 & n11748;
  assign n11750 = n53785 & n11749;
  assign n11751 = n11704 & n11750;
  assign n11752 = ~n344 & ~n1471;
  assign n11753 = ~n957 & n11752;
  assign n11754 = ~n848 & ~n894;
  assign n11755 = n4213 & n11754;
  assign n11756 = n11732 & n11755;
  assign n11757 = n11753 & n11756;
  assign n11758 = n53587 & n11757;
  assign n11759 = n11751 & n11758;
  assign n11760 = n11705 & n11715;
  assign n11761 = n54448 & n54451;
  assign n11762 = n2646 & n4002;
  assign n11763 = n4002 & n8793;
  assign n11764 = ~n984 & n11763;
  assign n11765 = ~n1769 & n11764;
  assign n11766 = n8793 & n11762;
  assign n11767 = ~n255 & ~n662;
  assign n11768 = ~n662 & ~n822;
  assign n11769 = ~n255 & n11768;
  assign n11770 = ~n822 & n11767;
  assign n11771 = ~n662 & n4070;
  assign n11772 = ~n255 & n11771;
  assign n11773 = ~n822 & n11772;
  assign n11774 = n4070 & n54453;
  assign n11775 = ~n307 & ~n511;
  assign n11776 = ~n307 & ~n1196;
  assign n11777 = ~n511 & n11776;
  assign n11778 = ~n1196 & n11775;
  assign n11779 = n624 & n9739;
  assign n11780 = n54455 & n11779;
  assign n11781 = n54454 & n11780;
  assign n11782 = n9739 & n54454;
  assign n11783 = n54452 & n11782;
  assign n11784 = n624 & n11783;
  assign n11785 = ~n1196 & n11784;
  assign n11786 = ~n307 & n11785;
  assign n11787 = ~n511 & n11786;
  assign n11788 = n54452 & n11780;
  assign n11789 = n54454 & n11788;
  assign n11790 = n54452 & n11781;
  assign n11791 = ~n1065 & ~n1191;
  assign n11792 = n6204 & n11791;
  assign n11793 = ~n357 & ~n740;
  assign n11794 = n916 & n6897;
  assign n11795 = n11793 & n11794;
  assign n11796 = ~n1065 & n11794;
  assign n11797 = ~n1191 & n11796;
  assign n11798 = ~n1469 & n11797;
  assign n11799 = ~n496 & n11798;
  assign n11800 = ~n357 & n11799;
  assign n11801 = ~n740 & n11800;
  assign n11802 = n6897 & n11791;
  assign n11803 = n916 & n6204;
  assign n11804 = n11793 & n11803;
  assign n11805 = n11802 & n11804;
  assign n11806 = ~n496 & ~n1191;
  assign n11807 = n11793 & n11806;
  assign n11808 = ~n1065 & ~n1469;
  assign n11809 = n6897 & n11808;
  assign n11810 = n916 & n11809;
  assign n11811 = n11807 & n11810;
  assign n11812 = n11792 & n11795;
  assign n11813 = ~n108 & ~n777;
  assign n11814 = ~n2201 & n11813;
  assign n11815 = ~n177 & ~n660;
  assign n11816 = n1816 & n11815;
  assign n11817 = n11814 & n11816;
  assign n11818 = ~n353 & ~n1634;
  assign n11819 = ~n1124 & ~n1715;
  assign n11820 = ~n1124 & ~n1634;
  assign n11821 = ~n353 & n11820;
  assign n11822 = ~n1715 & n11821;
  assign n11823 = ~n1634 & ~n1715;
  assign n11824 = ~n353 & ~n1124;
  assign n11825 = n11823 & n11824;
  assign n11826 = n11818 & n11819;
  assign n11827 = n53514 & n54458;
  assign n11828 = n11817 & n11827;
  assign n11829 = ~n1042 & ~n1472;
  assign n11830 = ~n922 & ~n1192;
  assign n11831 = n7471 & n11830;
  assign n11832 = n11829 & n11831;
  assign n11833 = n53940 & n11832;
  assign n11834 = ~n650 & ~n777;
  assign n11835 = ~n789 & n11834;
  assign n11836 = ~n777 & n11815;
  assign n11837 = n1816 & n7471;
  assign n11838 = n11836 & n11837;
  assign n11839 = n11816 & n11835;
  assign n11840 = n11827 & n54459;
  assign n11841 = ~n108 & ~n2201;
  assign n11842 = n11829 & n11830;
  assign n11843 = n11829 & n11841;
  assign n11844 = n11830 & n11843;
  assign n11845 = n11841 & n11842;
  assign n11846 = n53940 & n54460;
  assign n11847 = n11840 & n11846;
  assign n11848 = ~n922 & n11815;
  assign n11849 = ~n789 & ~n1192;
  assign n11850 = n11813 & n11849;
  assign n11851 = n11848 & n11850;
  assign n11852 = n11827 & n11851;
  assign n11853 = ~n650 & ~n2201;
  assign n11854 = n1816 & n11853;
  assign n11855 = n11829 & n11854;
  assign n11856 = n53940 & n11855;
  assign n11857 = n11852 & n11856;
  assign n11858 = n11828 & n11833;
  assign n11859 = n54457 & n54461;
  assign n11860 = n54456 & n11859;
  assign n11861 = n53514 & n1816;
  assign n11862 = n53940 & n11861;
  assign n11863 = n54458 & n11862;
  assign n11864 = n54451 & n11863;
  assign n11865 = n54457 & n11864;
  assign n11866 = n54448 & n11865;
  assign n11867 = n54456 & n11866;
  assign n11868 = n11829 & n11867;
  assign n11869 = ~n922 & n11868;
  assign n11870 = ~n1192 & n11869;
  assign n11871 = ~n108 & n11870;
  assign n11872 = ~n177 & n11871;
  assign n11873 = ~n660 & n11872;
  assign n11874 = ~n650 & n11873;
  assign n11875 = ~n777 & n11874;
  assign n11876 = ~n789 & n11875;
  assign n11877 = ~n2201 & n11876;
  assign n11878 = n11761 & n11860;
  assign n11879 = ~n54443 & ~n54462;
  assign n11880 = n54443 & n54462;
  assign n11881 = ~pi23  & ~n11879;
  assign n11882 = ~n11879 & ~n11880;
  assign n11883 = ~pi23  & n11882;
  assign n11884 = ~n11880 & n11881;
  assign n11885 = ~n11879 & ~n54463;
  assign n11886 = ~n54384 & n11885;
  assign n11887 = n54384 & ~n11885;
  assign n11888 = n10518 & ~n10520;
  assign n11889 = ~n10521 & ~n11888;
  assign n11890 = n1576 & n11889;
  assign n11891 = ~n53712 & n11215;
  assign n11892 = ~n53774 & n54403;
  assign n11893 = ~n53741 & n10564;
  assign n11894 = ~n11892 & ~n11893;
  assign n11895 = ~n11891 & ~n11892;
  assign n11896 = ~n11893 & n11895;
  assign n11897 = ~n11891 & n11894;
  assign n11898 = ~n11890 & n54464;
  assign n11899 = ~n11887 & n11898;
  assign n11900 = ~n11886 & ~n11898;
  assign n11901 = ~n11887 & ~n11900;
  assign n11902 = ~n11886 & ~n11887;
  assign n11903 = ~n11898 & n11902;
  assign n11904 = ~n11887 & ~n11903;
  assign n11905 = ~n11886 & ~n11899;
  assign n11906 = ~n54429 & ~n54465;
  assign n11907 = n54429 & n54465;
  assign n11908 = ~n11906 & ~n11907;
  assign n11909 = ~pi23  & ~n54463;
  assign n11910 = ~n11880 & n11885;
  assign n11911 = ~n11909 & ~n11910;
  assign n11912 = n10514 & ~n10516;
  assign n11913 = ~n10517 & ~n11912;
  assign n11914 = n1576 & n11913;
  assign n11915 = ~n53741 & n11215;
  assign n11916 = ~n53774 & n10564;
  assign n11917 = ~n53799 & n54403;
  assign n11918 = ~n11916 & ~n11917;
  assign n11919 = ~n11915 & ~n11916;
  assign n11920 = ~n11917 & n11919;
  assign n11921 = ~n11915 & n11918;
  assign n11922 = ~n11914 & ~n11917;
  assign n11923 = ~n11916 & n11922;
  assign n11924 = ~n11915 & n11923;
  assign n11925 = ~n11914 & n54466;
  assign n11926 = ~n11911 & ~n54467;
  assign n11927 = ~n292 & ~n296;
  assign n11928 = ~n296 & ~n1491;
  assign n11929 = ~n292 & n11928;
  assign n11930 = ~n292 & ~n1491;
  assign n11931 = ~n296 & n11930;
  assign n11932 = ~n1491 & n11927;
  assign n11933 = ~n450 & ~n883;
  assign n11934 = ~n450 & ~n1471;
  assign n11935 = ~n663 & ~n883;
  assign n11936 = n11934 & n11935;
  assign n11937 = n5850 & n11933;
  assign n11938 = n6289 & n11935;
  assign n11939 = n11934 & n11938;
  assign n11940 = n6289 & n54469;
  assign n11941 = ~n1471 & n54468;
  assign n11942 = ~n883 & n11941;
  assign n11943 = ~n663 & n11942;
  assign n11944 = ~n420 & n11943;
  assign n11945 = ~n409 & n11944;
  assign n11946 = ~n450 & n11945;
  assign n11947 = n54468 & n54470;
  assign n11948 = n4262 & n4798;
  assign n11949 = n5113 & n6577;
  assign n11950 = n11948 & n11949;
  assign n11951 = ~n163 & ~n829;
  assign n11952 = ~n1485 & n11951;
  assign n11953 = n10079 & n11952;
  assign n11954 = n4262 & n4753;
  assign n11955 = n11949 & n11954;
  assign n11956 = ~n1485 & n4798;
  assign n11957 = n3780 & n11951;
  assign n11958 = n11956 & n11957;
  assign n11959 = n11955 & n11958;
  assign n11960 = n4262 & n6577;
  assign n11961 = n10079 & n11960;
  assign n11962 = ~n1088 & ~n1485;
  assign n11963 = ~n829 & n11962;
  assign n11964 = ~n163 & ~n879;
  assign n11965 = n5113 & n11964;
  assign n11966 = n11963 & n11965;
  assign n11967 = n11961 & n11966;
  assign n11968 = n4753 & n5113;
  assign n11969 = n3780 & n6577;
  assign n11970 = n11968 & n11969;
  assign n11971 = ~n1088 & n11964;
  assign n11972 = ~n829 & ~n1485;
  assign n11973 = n4262 & n11972;
  assign n11974 = n11971 & n11973;
  assign n11975 = n11970 & n11974;
  assign n11976 = n11950 & n11953;
  assign n11977 = ~n415 & ~n1680;
  assign n11978 = n1265 & ~n1912;
  assign n11979 = ~n415 & n1265;
  assign n11980 = ~n1680 & n11979;
  assign n11981 = ~n1912 & n11980;
  assign n11982 = ~n1912 & n11977;
  assign n11983 = n1265 & n11982;
  assign n11984 = n11977 & n11978;
  assign n11985 = n4667 & n54473;
  assign n11986 = n54472 & n11985;
  assign n11987 = n54471 & n11986;
  assign n11988 = n53898 & n11987;
  assign n11989 = ~n776 & n8308;
  assign n11990 = ~n310 & ~n660;
  assign n11991 = n898 & n11990;
  assign n11992 = ~n310 & ~n776;
  assign n11993 = ~n660 & n11992;
  assign n11994 = n898 & n8308;
  assign n11995 = n11993 & n11994;
  assign n11996 = n11989 & n11991;
  assign n11997 = ~n310 & n54313;
  assign n11998 = ~n272 & n11997;
  assign n11999 = ~n660 & n11998;
  assign n12000 = ~n459 & n11999;
  assign n12001 = ~n1646 & n12000;
  assign n12002 = ~n423 & n12001;
  assign n12003 = ~n776 & n12002;
  assign n12004 = n54313 & n54474;
  assign n12005 = ~n618 & ~n956;
  assign n12006 = n4378 & n12005;
  assign n12007 = ~n216 & ~n1090;
  assign n12008 = ~n177 & ~n2042;
  assign n12009 = n12007 & n12008;
  assign n12010 = n4378 & n12007;
  assign n12011 = n12005 & n12008;
  assign n12012 = n12010 & n12011;
  assign n12013 = n12006 & n12009;
  assign n12014 = ~n295 & ~n319;
  assign n12015 = ~n422 & n12014;
  assign n12016 = n1266 & n2693;
  assign n12017 = n12015 & n12016;
  assign n12018 = ~n256 & ~n975;
  assign n12019 = ~n256 & ~n1997;
  assign n12020 = ~n975 & n12019;
  assign n12021 = ~n975 & ~n1997;
  assign n12022 = ~n256 & n12021;
  assign n12023 = ~n1997 & n12018;
  assign n12024 = n7688 & n54477;
  assign n12025 = n12017 & n12024;
  assign n12026 = n7688 & n12009;
  assign n12027 = ~n295 & ~n422;
  assign n12028 = ~n422 & ~n618;
  assign n12029 = ~n295 & n12028;
  assign n12030 = ~n618 & n12027;
  assign n12031 = n54477 & n54478;
  assign n12032 = n1266 & n2814;
  assign n12033 = n2693 & n4378;
  assign n12034 = n12032 & n12033;
  assign n12035 = n12031 & n12034;
  assign n12036 = n12026 & n12035;
  assign n12037 = n12009 & n12032;
  assign n12038 = n712 & n4378;
  assign n12039 = n586 & n2693;
  assign n12040 = n12038 & n12039;
  assign n12041 = n12031 & n12040;
  assign n12042 = n12037 & n12041;
  assign n12043 = n54476 & n12025;
  assign n12044 = n12007 & n54477;
  assign n12045 = n12008 & n12044;
  assign n12046 = n1266 & n12045;
  assign n12047 = n2814 & n12046;
  assign n12048 = n586 & n12047;
  assign n12049 = n4378 & n12048;
  assign n12050 = n54475 & n12049;
  assign n12051 = n712 & n12050;
  assign n12052 = n2693 & n12051;
  assign n12053 = ~n422 & n12052;
  assign n12054 = ~n295 & n12053;
  assign n12055 = ~n618 & n12054;
  assign n12056 = n54475 & n54479;
  assign n12057 = n54239 & n54480;
  assign n12058 = n4262 & n4667;
  assign n12059 = n6577 & n12058;
  assign n12060 = n54473 & n12059;
  assign n12061 = n4753 & n12060;
  assign n12062 = n53898 & n12061;
  assign n12063 = n54239 & n12062;
  assign n12064 = n3780 & n12063;
  assign n12065 = n54471 & n12064;
  assign n12066 = n54480 & n12065;
  assign n12067 = n5113 & n12066;
  assign n12068 = ~n1088 & n12067;
  assign n12069 = ~n879 & n12068;
  assign n12070 = ~n1485 & n12069;
  assign n12071 = ~n163 & n12070;
  assign n12072 = ~n829 & n12071;
  assign n12073 = n11988 & n12057;
  assign n12074 = n54443 & ~n54481;
  assign n12075 = ~n54443 & n54481;
  assign n12076 = ~n12074 & ~n12075;
  assign n12077 = n1670 & n4470;
  assign n12078 = n2038 & n4585;
  assign n12079 = n9972 & n12078;
  assign n12080 = n9972 & n12077;
  assign n12081 = n12078 & n12080;
  assign n12082 = n12077 & n12079;
  assign n12083 = n2980 & n3715;
  assign n12084 = n4892 & n12083;
  assign n12085 = ~n161 & ~n511;
  assign n12086 = ~n740 & ~n922;
  assign n12087 = n12085 & n12086;
  assign n12088 = n2404 & n12087;
  assign n12089 = n12084 & n12088;
  assign n12090 = n9972 & n12087;
  assign n12091 = n2404 & n12090;
  assign n12092 = n4585 & n4892;
  assign n12093 = n2038 & n12092;
  assign n12094 = n2980 & n4470;
  assign n12095 = n1670 & n3715;
  assign n12096 = n12094 & n12095;
  assign n12097 = n12093 & n12096;
  assign n12098 = n12091 & n12097;
  assign n12099 = n2980 & n8091;
  assign n12100 = n12087 & n12099;
  assign n12101 = n2404 & n12100;
  assign n12102 = n2038 & n4892;
  assign n12103 = n3715 & n12102;
  assign n12104 = n4585 & n6482;
  assign n12105 = n12077 & n12104;
  assign n12106 = n12103 & n12105;
  assign n12107 = n12101 & n12106;
  assign n12108 = n54482 & n12089;
  assign n12109 = n53938 & n54483;
  assign n12110 = n53584 & n12109;
  assign n12111 = n1957 & n4751;
  assign n12112 = ~n460 & ~n1337;
  assign n12113 = n10830 & n12112;
  assign n12114 = n12111 & n12113;
  assign n12115 = ~n294 & ~n562;
  assign n12116 = ~n308 & ~n754;
  assign n12117 = ~n294 & ~n308;
  assign n12118 = ~n562 & ~n754;
  assign n12119 = n12117 & n12118;
  assign n12120 = n12115 & n12116;
  assign n12121 = n775 & n2537;
  assign n12122 = n54484 & n12121;
  assign n12123 = n54468 & n12122;
  assign n12124 = n2537 & n10830;
  assign n12125 = n12111 & n12124;
  assign n12126 = ~n308 & ~n460;
  assign n12127 = n12115 & n12126;
  assign n12128 = ~n754 & ~n1337;
  assign n12129 = n775 & n12128;
  assign n12130 = n12127 & n12129;
  assign n12131 = n54468 & n12130;
  assign n12132 = n12125 & n12131;
  assign n12133 = n12111 & n12121;
  assign n12134 = ~n460 & ~n562;
  assign n12135 = n12116 & n12134;
  assign n12136 = ~n294 & ~n560;
  assign n12137 = ~n1125 & ~n1337;
  assign n12138 = n12136 & n12137;
  assign n12139 = n12135 & n12138;
  assign n12140 = n54468 & n12139;
  assign n12141 = n12133 & n12140;
  assign n12142 = n12114 & n12123;
  assign n12143 = ~n246 & ~n612;
  assign n12144 = n3675 & n12143;
  assign n12145 = n964 & n11977;
  assign n12146 = n12144 & n12145;
  assign n12147 = ~n750 & ~n1634;
  assign n12148 = ~n1081 & n12147;
  assign n12149 = n54355 & n12148;
  assign n12150 = n964 & n54355;
  assign n12151 = n3675 & n12150;
  assign n12152 = ~n415 & n12151;
  assign n12153 = ~n1680 & n12152;
  assign n12154 = ~n1081 & n12153;
  assign n12155 = ~n246 & n12154;
  assign n12156 = ~n612 & n12155;
  assign n12157 = ~n1634 & n12156;
  assign n12158 = ~n750 & n12157;
  assign n12159 = ~n750 & ~n1081;
  assign n12160 = n964 & n12159;
  assign n12161 = n3675 & n11977;
  assign n12162 = n12160 & n12161;
  assign n12163 = ~n1634 & n12143;
  assign n12164 = n54355 & n12163;
  assign n12165 = n12162 & n12164;
  assign n12166 = ~n750 & ~n1680;
  assign n12167 = n8534 & n12166;
  assign n12168 = n964 & n3675;
  assign n12169 = n12167 & n12168;
  assign n12170 = ~n1081 & n12143;
  assign n12171 = n54355 & n12170;
  assign n12172 = n12169 & n12171;
  assign n12173 = n12146 & n12149;
  assign n12174 = n54128 & n54486;
  assign n12175 = n4751 & n54468;
  assign n12176 = n54486 & n12175;
  assign n12177 = n2537 & n12176;
  assign n12178 = n775 & n12177;
  assign n12179 = n1957 & n12178;
  assign n12180 = n54128 & n12179;
  assign n12181 = ~n1125 & n12180;
  assign n12182 = ~n308 & n12181;
  assign n12183 = ~n294 & n12182;
  assign n12184 = ~n560 & n12183;
  assign n12185 = ~n562 & n12184;
  assign n12186 = ~n1337 & n12185;
  assign n12187 = ~n460 & n12186;
  assign n12188 = ~n754 & n12187;
  assign n12189 = n54485 & n12174;
  assign n12190 = n2740 & n53987;
  assign n12191 = n53987 & n54339;
  assign n12192 = n2740 & n12191;
  assign n12193 = n54339 & n12190;
  assign n12194 = n906 & n3086;
  assign n12195 = n586 & n906;
  assign n12196 = n3086 & n12195;
  assign n12197 = n586 & n12194;
  assign n12198 = ~n414 & ~n771;
  assign n12199 = ~n414 & ~n975;
  assign n12200 = ~n771 & n12199;
  assign n12201 = ~n975 & n12198;
  assign n12202 = n175 & n2981;
  assign n12203 = n54490 & n12202;
  assign n12204 = n586 & n12202;
  assign n12205 = n12194 & n54490;
  assign n12206 = n12204 & n12205;
  assign n12207 = n54489 & n12203;
  assign n12208 = ~n310 & n8863;
  assign n12209 = ~n510 & ~n631;
  assign n12210 = ~n510 & ~n514;
  assign n12211 = ~n631 & n12210;
  assign n12212 = ~n514 & n12209;
  assign n12213 = n2334 & n8753;
  assign n12214 = ~n631 & n8753;
  assign n12215 = ~n1997 & n12214;
  assign n12216 = ~n977 & n12215;
  assign n12217 = ~n514 & n12216;
  assign n12218 = ~n510 & n12217;
  assign n12219 = ~n514 & ~n977;
  assign n12220 = ~n631 & n12219;
  assign n12221 = ~n510 & ~n1997;
  assign n12222 = n8753 & n12221;
  assign n12223 = n12220 & n12222;
  assign n12224 = n54492 & n12213;
  assign n12225 = n12208 & n54493;
  assign n12226 = n54491 & n12225;
  assign n12227 = n12190 & n12208;
  assign n12228 = n2981 & n12227;
  assign n12229 = n54493 & n12228;
  assign n12230 = n3086 & n12229;
  assign n12231 = n54339 & n12230;
  assign n12232 = n586 & n12231;
  assign n12233 = n906 & n12232;
  assign n12234 = n175 & n12233;
  assign n12235 = ~n414 & n12234;
  assign n12236 = ~n975 & n12235;
  assign n12237 = ~n771 & n12236;
  assign n12238 = n54488 & n12226;
  assign n12239 = n54487 & n54494;
  assign n12240 = n2038 & n2404;
  assign n12241 = n4470 & n12240;
  assign n12242 = n4892 & n12241;
  assign n12243 = n3715 & n12242;
  assign n12244 = n53938 & n12243;
  assign n12245 = n53584 & n12244;
  assign n12246 = n54494 & n12245;
  assign n12247 = n4585 & n12246;
  assign n12248 = n54487 & n12247;
  assign n12249 = n8091 & n12248;
  assign n12250 = n6482 & n12249;
  assign n12251 = n1670 & n12250;
  assign n12252 = ~n922 & n12251;
  assign n12253 = ~n161 & n12252;
  assign n12254 = ~n249 & n12253;
  assign n12255 = ~n1280 & n12254;
  assign n12256 = ~n511 & n12255;
  assign n12257 = ~n740 & n12256;
  assign n12258 = n12110 & n12239;
  assign n12259 = ~n901 & ~n1125;
  assign n12260 = n846 & n12259;
  assign n12261 = n1265 & n3062;
  assign n12262 = n12260 & n12261;
  assign n12263 = ~n450 & ~n465;
  assign n12264 = n403 & ~n465;
  assign n12265 = ~n450 & n12264;
  assign n12266 = n403 & n12263;
  assign n12267 = ~n651 & ~n2109;
  assign n12268 = ~n651 & n11829;
  assign n12269 = ~n2109 & n12268;
  assign n12270 = n11829 & n12267;
  assign n12271 = n54496 & n54497;
  assign n12272 = n12262 & n12271;
  assign n12273 = ~n206 & ~n218;
  assign n12274 = ~n1124 & n12273;
  assign n12275 = ~n182 & ~n441;
  assign n12276 = n10184 & n12275;
  assign n12277 = n5361 & n10184;
  assign n12278 = ~n218 & n12277;
  assign n12279 = ~n206 & n12278;
  assign n12280 = ~n441 & n12279;
  assign n12281 = ~n206 & ~n441;
  assign n12282 = ~n218 & n12281;
  assign n12283 = ~n441 & n12273;
  assign n12284 = n12277 & n54499;
  assign n12285 = n12274 & n12276;
  assign n12286 = ~n774 & ~n1487;
  assign n12287 = n2039 & n8860;
  assign n12288 = n12286 & n12287;
  assign n12289 = n1670 & n5113;
  assign n12290 = n1672 & n5943;
  assign n12291 = n12289 & n12290;
  assign n12292 = n12288 & n12291;
  assign n12293 = n54498 & n12292;
  assign n12294 = n8860 & n54497;
  assign n12295 = n54496 & n12294;
  assign n12296 = n12286 & n12295;
  assign n12297 = n846 & n12296;
  assign n12298 = n1265 & n12297;
  assign n12299 = n5943 & n12298;
  assign n12300 = n1672 & n12299;
  assign n12301 = n5113 & n12300;
  assign n12302 = n54498 & n12301;
  assign n12303 = n3062 & n12302;
  assign n12304 = n1670 & n12303;
  assign n12305 = ~n1125 & n12304;
  assign n12306 = ~n901 & n12305;
  assign n12307 = ~n177 & n12306;
  assign n12308 = ~n311 & n12307;
  assign n12309 = n5113 & n12259;
  assign n12310 = n12261 & n12309;
  assign n12311 = n12271 & n12310;
  assign n12312 = n846 & n1670;
  assign n12313 = n12290 & n12312;
  assign n12314 = n12288 & n12313;
  assign n12315 = n54498 & n12314;
  assign n12316 = n12311 & n12315;
  assign n12317 = n2039 & n12259;
  assign n12318 = n1265 & n8860;
  assign n12319 = n12317 & n12318;
  assign n12320 = n12271 & n12319;
  assign n12321 = n12286 & n12290;
  assign n12322 = n3062 & n5113;
  assign n12323 = n12312 & n12322;
  assign n12324 = n12321 & n12323;
  assign n12325 = n54498 & n12324;
  assign n12326 = n12320 & n12325;
  assign n12327 = n12272 & n12293;
  assign n12328 = ~n587 & n4021;
  assign n12329 = ~n101 & ~n1634;
  assign n12330 = n12328 & n12329;
  assign n12331 = n905 & n4026;
  assign n12332 = ~n464 & ~n1681;
  assign n12333 = ~n1471 & ~n1681;
  assign n12334 = ~n464 & n12333;
  assign n12335 = ~n464 & ~n1471;
  assign n12336 = ~n1681 & n12335;
  assign n12337 = ~n1471 & n12332;
  assign n12338 = n12331 & n54501;
  assign n12339 = ~n628 & n4587;
  assign n12340 = ~n567 & n5021;
  assign n12341 = n12339 & n12340;
  assign n12342 = n12338 & n12341;
  assign n12343 = ~n101 & ~n567;
  assign n12344 = ~n1634 & n12343;
  assign n12345 = n5021 & n12344;
  assign n12346 = n12331 & n12339;
  assign n12347 = n12328 & n54501;
  assign n12348 = n12346 & n12347;
  assign n12349 = n12345 & n12348;
  assign n12350 = n4021 & n5021;
  assign n12351 = n4021 & n4026;
  assign n12352 = n905 & n5021;
  assign n12353 = n12351 & n12352;
  assign n12354 = n12331 & n12350;
  assign n12355 = ~n567 & ~n587;
  assign n12356 = n12329 & n12355;
  assign n12357 = n12339 & n12356;
  assign n12358 = n54501 & n12356;
  assign n12359 = n12339 & n12358;
  assign n12360 = n54501 & n12357;
  assign n12361 = n54503 & n54504;
  assign n12362 = n12330 & n12342;
  assign n12363 = n1642 & n2690;
  assign n12364 = n4377 & n4584;
  assign n12365 = n12363 & n12364;
  assign n12366 = ~n511 & ~n733;
  assign n12367 = ~n1065 & n12366;
  assign n12368 = ~n275 & ~n649;
  assign n12369 = ~n163 & ~n354;
  assign n12370 = n12368 & n12369;
  assign n12371 = ~n163 & ~n733;
  assign n12372 = ~n1065 & n12371;
  assign n12373 = ~n354 & ~n511;
  assign n12374 = n12368 & n12373;
  assign n12375 = n12372 & n12374;
  assign n12376 = n12367 & n12370;
  assign n12377 = n2690 & n4584;
  assign n12378 = n1642 & n12377;
  assign n12379 = ~n1065 & n12378;
  assign n12380 = ~n163 & n12379;
  assign n12381 = ~n275 & n12380;
  assign n12382 = ~n511 & n12381;
  assign n12383 = ~n461 & n12382;
  assign n12384 = ~n649 & n12383;
  assign n12385 = ~n733 & n12384;
  assign n12386 = ~n354 & n12385;
  assign n12387 = ~n1881 & n12386;
  assign n12388 = ~n461 & ~n649;
  assign n12389 = n2690 & n12388;
  assign n12390 = n1642 & n4584;
  assign n12391 = n12389 & n12390;
  assign n12392 = ~n275 & ~n511;
  assign n12393 = ~n354 & n12392;
  assign n12394 = ~n733 & ~n1881;
  assign n12395 = ~n163 & ~n1065;
  assign n12396 = n12394 & n12395;
  assign n12397 = n12393 & n12396;
  assign n12398 = n12391 & n12397;
  assign n12399 = ~n733 & ~n1065;
  assign n12400 = n1642 & n12399;
  assign n12401 = n12377 & n12400;
  assign n12402 = ~n275 & n1401;
  assign n12403 = ~n649 & ~n1881;
  assign n12404 = ~n163 & ~n511;
  assign n12405 = n12403 & n12404;
  assign n12406 = n12402 & n12405;
  assign n12407 = n12401 & n12406;
  assign n12408 = n12365 & n54505;
  assign n12409 = n54048 & n54506;
  assign n12410 = n54501 & n12339;
  assign n12411 = n4021 & n12410;
  assign n12412 = n54048 & n12411;
  assign n12413 = n54506 & n12412;
  assign n12414 = n4026 & n12413;
  assign n12415 = n5021 & n12414;
  assign n12416 = n905 & n12415;
  assign n12417 = ~n101 & n12416;
  assign n12418 = ~n567 & n12417;
  assign n12419 = ~n1634 & n12418;
  assign n12420 = ~n587 & n12419;
  assign n12421 = n54502 & n12409;
  assign n12422 = n3475 & n3676;
  assign n12423 = n1704 & n4261;
  assign n12424 = n12422 & n12423;
  assign n12425 = ~n588 & ~n735;
  assign n12426 = ~n750 & ~n1997;
  assign n12427 = ~n735 & ~n750;
  assign n12428 = ~n588 & ~n1997;
  assign n12429 = n12427 & n12428;
  assign n12430 = n12425 & n12426;
  assign n12431 = n54223 & n54508;
  assign n12432 = n12424 & n12431;
  assign n12433 = n53711 & n12432;
  assign n12434 = ~n564 & ~n615;
  assign n12435 = n2328 & n12434;
  assign n12436 = ~n174 & ~n296;
  assign n12437 = n5476 & n12436;
  assign n12438 = n12435 & n12437;
  assign n12439 = ~n1644 & ~n2042;
  assign n12440 = ~n1031 & n12439;
  assign n12441 = ~n141 & ~n316;
  assign n12442 = ~n361 & ~n1234;
  assign n12443 = n12441 & n12442;
  assign n12444 = n12440 & n12443;
  assign n12445 = ~n902 & n2328;
  assign n12446 = ~n1031 & n12445;
  assign n12447 = ~n316 & n12446;
  assign n12448 = ~n296 & n12447;
  assign n12449 = ~n174 & n12448;
  assign n12450 = ~n141 & n12449;
  assign n12451 = ~n564 & n12450;
  assign n12452 = ~n584 & n12451;
  assign n12453 = ~n1234 & n12452;
  assign n12454 = ~n1644 & n12453;
  assign n12455 = ~n615 & n12454;
  assign n12456 = ~n361 & n12455;
  assign n12457 = ~n2042 & n12456;
  assign n12458 = ~n361 & ~n615;
  assign n12459 = n2328 & n12458;
  assign n12460 = n12437 & n12459;
  assign n12461 = ~n564 & ~n1234;
  assign n12462 = n12441 & n12461;
  assign n12463 = n12440 & n12462;
  assign n12464 = n12460 & n12463;
  assign n12465 = ~n1234 & ~n2042;
  assign n12466 = ~n316 & ~n361;
  assign n12467 = n12465 & n12466;
  assign n12468 = n2328 & n5476;
  assign n12469 = n12467 & n12468;
  assign n12470 = ~n296 & ~n615;
  assign n12471 = ~n141 & n12470;
  assign n12472 = ~n174 & ~n564;
  assign n12473 = ~n1031 & ~n1644;
  assign n12474 = n12472 & n12473;
  assign n12475 = n12471 & n12474;
  assign n12476 = n12469 & n12475;
  assign n12477 = ~n584 & ~n1234;
  assign n12478 = n12439 & n12477;
  assign n12479 = ~n174 & ~n615;
  assign n12480 = n2328 & n12479;
  assign n12481 = n12478 & n12480;
  assign n12482 = ~n316 & ~n564;
  assign n12483 = ~n296 & n12482;
  assign n12484 = ~n361 & ~n1031;
  assign n12485 = ~n141 & ~n902;
  assign n12486 = n12484 & n12485;
  assign n12487 = n12483 & n12486;
  assign n12488 = n12481 & n12487;
  assign n12489 = n12438 & n12444;
  assign n12490 = ~n747 & ~n832;
  assign n12491 = n772 & n9511;
  assign n12492 = n12490 & n12491;
  assign n12493 = ~n179 & ~n631;
  assign n12494 = ~n466 & ~n631;
  assign n12495 = ~n179 & n12494;
  assign n12496 = ~n179 & ~n466;
  assign n12497 = ~n631 & n12496;
  assign n12498 = ~n466 & n12493;
  assign n12499 = ~n342 & ~n622;
  assign n12500 = ~n342 & ~n1337;
  assign n12501 = ~n622 & n12500;
  assign n12502 = ~n1337 & n12499;
  assign n12503 = n54510 & n54511;
  assign n12504 = n772 & n54510;
  assign n12505 = n9511 & n12504;
  assign n12506 = ~n1337 & n12505;
  assign n12507 = ~n832 & n12506;
  assign n12508 = ~n342 & n12507;
  assign n12509 = ~n747 & n12508;
  assign n12510 = ~n622 & n12509;
  assign n12511 = ~n622 & ~n1337;
  assign n12512 = n772 & n12511;
  assign n12513 = n9511 & n12512;
  assign n12514 = ~n342 & n12490;
  assign n12515 = n54510 & n12514;
  assign n12516 = n12513 & n12515;
  assign n12517 = n12492 & n12503;
  assign n12518 = n54509 & n54512;
  assign n12519 = n12432 & n54512;
  assign n12520 = n53711 & n54509;
  assign n12521 = n12519 & n12520;
  assign n12522 = n12433 & n12518;
  assign n12523 = n54507 & n54513;
  assign n12524 = n3676 & n54223;
  assign n12525 = n53711 & n12524;
  assign n12526 = n54509 & n12525;
  assign n12527 = n54507 & n12526;
  assign n12528 = n54500 & n12527;
  assign n12529 = n54512 & n12528;
  assign n12530 = n4261 & n12529;
  assign n12531 = n1704 & n12530;
  assign n12532 = n3475 & n12531;
  assign n12533 = ~n1997 & n12532;
  assign n12534 = ~n750 & n12533;
  assign n12535 = ~n735 & n12534;
  assign n12536 = ~n588 & n12535;
  assign n12537 = n54500 & n54513;
  assign n12538 = n54507 & n12537;
  assign n12539 = n54500 & n12523;
  assign n12540 = ~n54495 & ~n54514;
  assign n12541 = n54495 & n54514;
  assign n12542 = ~pi20  & ~n12540;
  assign n12543 = ~n12540 & ~n12541;
  assign n12544 = ~pi20  & n12543;
  assign n12545 = ~n12541 & n12542;
  assign n12546 = ~n12540 & ~n54515;
  assign n12547 = ~n54481 & n12546;
  assign n12548 = n54481 & ~n12546;
  assign n12549 = n10506 & ~n10508;
  assign n12550 = ~n10509 & ~n12549;
  assign n12551 = n1576 & n12550;
  assign n12552 = ~n53819 & n10564;
  assign n12553 = ~n53845 & n54403;
  assign n12554 = ~n53799 & n11215;
  assign n12555 = ~n12553 & ~n12554;
  assign n12556 = ~n12552 & ~n12553;
  assign n12557 = ~n12554 & n12556;
  assign n12558 = ~n12552 & n12555;
  assign n12559 = ~n12551 & n54516;
  assign n12560 = ~n12548 & n12559;
  assign n12561 = ~n12547 & ~n12559;
  assign n12562 = ~n12548 & ~n12561;
  assign n12563 = ~n12547 & ~n12548;
  assign n12564 = ~n12559 & n12563;
  assign n12565 = ~n12548 & ~n12564;
  assign n12566 = ~n12547 & ~n12560;
  assign n12567 = ~n12074 & ~n54517;
  assign n12568 = ~n12075 & n12567;
  assign n12569 = n12076 & ~n54517;
  assign n12570 = ~n12074 & ~n54518;
  assign n12571 = n11911 & n54467;
  assign n12572 = ~n11926 & ~n12571;
  assign n12573 = ~n12570 & n12572;
  assign n12574 = ~n11926 & ~n12573;
  assign n12575 = n11898 & ~n11902;
  assign n12576 = ~n11898 & ~n11903;
  assign n12577 = n11902 & ~n11903;
  assign n12578 = ~n12576 & ~n12577;
  assign n12579 = ~n11903 & ~n12575;
  assign n12580 = ~n12574 & ~n54519;
  assign n12581 = n12574 & n54519;
  assign n12582 = ~n12580 & ~n12581;
  assign n12583 = n11213 & n11279;
  assign n12584 = n54407 & ~n54409;
  assign n12585 = ~n53650 & n12584;
  assign n12586 = ~n53685 & n54410;
  assign n12587 = ~n53657 & n11267;
  assign n12588 = ~n12586 & ~n12587;
  assign n12589 = ~n12585 & n12588;
  assign n12590 = ~n11279 & n12589;
  assign n12591 = ~n11213 & n12589;
  assign n12592 = ~n12590 & ~n12591;
  assign n12593 = ~n12583 & n12589;
  assign n12594 = pi29  & ~n54520;
  assign n12595 = ~pi29  & n54520;
  assign n12596 = ~n12594 & ~n12595;
  assign n12597 = n12582 & ~n12596;
  assign n12598 = ~n12580 & ~n12597;
  assign n12599 = n11908 & ~n12598;
  assign n12600 = ~n11906 & ~n12599;
  assign n12601 = n11389 & ~n11391;
  assign n12602 = ~n11389 & ~n11392;
  assign n12603 = n11391 & ~n11392;
  assign n12604 = ~n12602 & ~n12603;
  assign n12605 = ~n11392 & ~n12601;
  assign n12606 = ~n12600 & ~n54521;
  assign n12607 = n11242 & n11279;
  assign n12608 = ~n53650 & n54410;
  assign n12609 = ~n2325 & n12584;
  assign n12610 = ~n53634 & n11267;
  assign n12611 = ~n12609 & ~n12610;
  assign n12612 = ~n12608 & ~n12610;
  assign n12613 = ~n12609 & n12612;
  assign n12614 = ~n12608 & n12611;
  assign n12615 = ~n12607 & n54522;
  assign n12616 = pi29  & ~n12615;
  assign n12617 = pi29  & ~n12616;
  assign n12618 = pi29  & n12615;
  assign n12619 = ~n12615 & ~n12616;
  assign n12620 = ~pi29  & ~n12615;
  assign n12621 = ~n54523 & ~n54524;
  assign n12622 = n12600 & n54521;
  assign n12623 = ~n12600 & ~n12606;
  assign n12624 = ~n54521 & ~n12606;
  assign n12625 = ~n12623 & ~n12624;
  assign n12626 = ~n12606 & ~n12622;
  assign n12627 = ~n12621 & ~n54525;
  assign n12628 = ~n12606 & ~n12627;
  assign n12629 = n11412 & ~n11414;
  assign n12630 = n11414 & ~n11415;
  assign n12631 = n11412 & n11414;
  assign n12632 = ~n11412 & ~n11415;
  assign n12633 = ~n11412 & ~n11414;
  assign n12634 = ~n54526 & ~n54527;
  assign n12635 = ~n11415 & ~n12629;
  assign n12636 = ~n12628 & ~n54528;
  assign n12637 = n12628 & n54528;
  assign n12638 = ~n12636 & ~n12637;
  assign n12639 = n123 & ~n10547;
  assign n12640 = ~n53444 & ~n12639;
  assign n12641 = n123 & n10551;
  assign n12642 = n53444 & ~n2325;
  assign n12643 = ~n12641 & ~n12642;
  assign n12644 = ~n2325 & ~n12640;
  assign n12645 = pi26  & ~n54529;
  assign n12646 = ~n54529 & ~n12645;
  assign n12647 = ~pi26  & ~n54529;
  assign n12648 = pi26  & ~n12645;
  assign n12649 = pi26  & n54529;
  assign n12650 = ~n54530 & ~n54531;
  assign n12651 = n11279 & n11286;
  assign n12652 = ~n53650 & n11267;
  assign n12653 = ~n53657 & n54410;
  assign n12654 = ~n53634 & n12584;
  assign n12655 = ~n12653 & ~n12654;
  assign n12656 = ~n12652 & ~n12653;
  assign n12657 = ~n12654 & n12656;
  assign n12658 = ~n12652 & n12655;
  assign n12659 = ~n12651 & n54532;
  assign n12660 = pi29  & ~n12659;
  assign n12661 = pi29  & ~n12660;
  assign n12662 = pi29  & n12659;
  assign n12663 = ~n12659 & ~n12660;
  assign n12664 = ~pi29  & ~n12659;
  assign n12665 = ~n54533 & ~n54534;
  assign n12666 = ~n12650 & ~n12665;
  assign n12667 = ~n11908 & n12598;
  assign n12668 = ~n12599 & ~n12667;
  assign n12669 = n12650 & n12665;
  assign n12670 = ~n12650 & ~n12666;
  assign n12671 = ~n12665 & ~n12666;
  assign n12672 = ~n12670 & ~n12671;
  assign n12673 = ~n12666 & ~n12669;
  assign n12674 = n12668 & ~n54535;
  assign n12675 = ~n12666 & ~n12674;
  assign n12676 = n12621 & n54525;
  assign n12677 = ~n54525 & ~n12627;
  assign n12678 = ~n12621 & ~n12627;
  assign n12679 = ~n12677 & ~n12678;
  assign n12680 = ~n12627 & ~n12676;
  assign n12681 = ~n12675 & ~n54536;
  assign n12682 = ~n12582 & n12596;
  assign n12683 = ~n12597 & ~n12682;
  assign n12684 = ~n12076 & n54517;
  assign n12685 = ~n54517 & ~n54518;
  assign n12686 = ~n12075 & n12570;
  assign n12687 = ~n12685 & ~n12686;
  assign n12688 = ~n54518 & ~n12684;
  assign n12689 = n10510 & ~n10512;
  assign n12690 = ~n10513 & ~n12689;
  assign n12691 = n1576 & n12690;
  assign n12692 = ~n53819 & n54403;
  assign n12693 = ~n53799 & n10564;
  assign n12694 = ~n53774 & n11215;
  assign n12695 = ~n12693 & ~n12694;
  assign n12696 = ~n12692 & n12695;
  assign n12697 = ~n12691 & ~n12692;
  assign n12698 = ~n12693 & n12697;
  assign n12699 = ~n12694 & n12698;
  assign n12700 = ~n12691 & n12696;
  assign n12701 = ~n54537 & ~n54538;
  assign n12702 = ~n461 & ~n901;
  assign n12703 = ~n901 & n6621;
  assign n12704 = ~n461 & n12703;
  assign n12705 = n6621 & n12702;
  assign n12706 = n1673 & n4197;
  assign n12707 = n1091 & n5538;
  assign n12708 = n12706 & n12707;
  assign n12709 = n54539 & n12708;
  assign n12710 = ~n733 & n5873;
  assign n12711 = n5873 & n5943;
  assign n12712 = ~n733 & n12711;
  assign n12713 = ~n733 & n5943;
  assign n12714 = n5873 & n12713;
  assign n12715 = n5943 & n12710;
  assign n12716 = ~n754 & ~n1061;
  assign n12717 = ~n1062 & n12716;
  assign n12718 = ~n754 & n1063;
  assign n12719 = n802 & ~n1062;
  assign n12720 = ~n1061 & n12719;
  assign n12721 = ~n754 & n12720;
  assign n12722 = n802 & n54541;
  assign n12723 = n54540 & n54542;
  assign n12724 = n12708 & n54540;
  assign n12725 = n54539 & n54542;
  assign n12726 = n12724 & n12725;
  assign n12727 = n12709 & n12723;
  assign n12728 = ~n977 & ~n1535;
  assign n12729 = ~n896 & n12728;
  assign n12730 = ~n320 & ~n1644;
  assign n12731 = ~n177 & ~n292;
  assign n12732 = n10300 & n12731;
  assign n12733 = n12730 & n12732;
  assign n12734 = ~n896 & n10300;
  assign n12735 = ~n320 & n12734;
  assign n12736 = ~n977 & n12735;
  assign n12737 = ~n177 & n12736;
  assign n12738 = ~n292 & n12737;
  assign n12739 = ~n1535 & n12738;
  assign n12740 = ~n1644 & n12739;
  assign n12741 = ~n896 & ~n977;
  assign n12742 = ~n292 & n12741;
  assign n12743 = ~n177 & ~n1535;
  assign n12744 = n10300 & n12743;
  assign n12745 = n12730 & n12744;
  assign n12746 = n12742 & n12745;
  assign n12747 = ~n320 & ~n977;
  assign n12748 = ~n177 & n12747;
  assign n12749 = ~n896 & ~n1644;
  assign n12750 = ~n292 & ~n1535;
  assign n12751 = n12749 & n12750;
  assign n12752 = n10300 & n12751;
  assign n12753 = n12748 & n12752;
  assign n12754 = n12729 & n12733;
  assign n12755 = ~n618 & ~n2042;
  assign n12756 = ~n1491 & ~n1715;
  assign n12757 = ~n618 & ~n1715;
  assign n12758 = ~n1491 & ~n2042;
  assign n12759 = n12757 & n12758;
  assign n12760 = ~n1715 & ~n2042;
  assign n12761 = ~n618 & ~n1491;
  assign n12762 = n12760 & n12761;
  assign n12763 = n12755 & n12756;
  assign n12764 = n53699 & n54545;
  assign n12765 = n53775 & n12764;
  assign n12766 = n54544 & n12765;
  assign n12767 = n53699 & n54540;
  assign n12768 = n54542 & n12767;
  assign n12769 = n53775 & n12768;
  assign n12770 = n5538 & n12769;
  assign n12771 = n54539 & n12770;
  assign n12772 = n54544 & n12771;
  assign n12773 = n1091 & n12772;
  assign n12774 = n1673 & n12773;
  assign n12775 = ~n879 & n12774;
  assign n12776 = ~n1491 & n12775;
  assign n12777 = ~n172 & n12776;
  assign n12778 = ~n618 & n12777;
  assign n12779 = ~n1715 & n12778;
  assign n12780 = ~n2042 & n12779;
  assign n12781 = n1673 & n12760;
  assign n12782 = n12707 & n12781;
  assign n12783 = n54539 & n12782;
  assign n12784 = n12723 & n12783;
  assign n12785 = n4197 & n12761;
  assign n12786 = n53775 & n12785;
  assign n12787 = n53699 & n12786;
  assign n12788 = n54544 & n12787;
  assign n12789 = n12784 & n12788;
  assign n12790 = n54543 & n12766;
  assign n12791 = ~n1881 & ~n2103;
  assign n12792 = ~n1487 & n12791;
  assign n12793 = ~n179 & ~n216;
  assign n12794 = ~n415 & ~n646;
  assign n12795 = n5156 & n12794;
  assign n12796 = n12793 & n12795;
  assign n12797 = ~n415 & ~n1487;
  assign n12798 = ~n415 & ~n2103;
  assign n12799 = ~n1487 & n12798;
  assign n12800 = ~n2103 & n12797;
  assign n12801 = ~n179 & n54547;
  assign n12802 = ~n321 & n12801;
  assign n12803 = ~n216 & n12802;
  assign n12804 = ~n404 & n12803;
  assign n12805 = ~n646 & n12804;
  assign n12806 = ~n1881 & n12805;
  assign n12807 = ~n646 & ~n1881;
  assign n12808 = n5156 & n12807;
  assign n12809 = n12793 & n12808;
  assign n12810 = n54547 & n12809;
  assign n12811 = ~n1487 & n12793;
  assign n12812 = ~n404 & ~n1881;
  assign n12813 = ~n321 & ~n2103;
  assign n12814 = n12812 & n12813;
  assign n12815 = n12794 & n12814;
  assign n12816 = n12811 & n12815;
  assign n12817 = n12792 & n12796;
  assign n12818 = ~n344 & ~n491;
  assign n12819 = ~n1769 & n12818;
  assign n12820 = n53766 & n12819;
  assign n12821 = n4530 & n5021;
  assign n12822 = n54360 & n12821;
  assign n12823 = n54360 & n12819;
  assign n12824 = n53766 & n12821;
  assign n12825 = n12823 & n12824;
  assign n12826 = n12820 & n12822;
  assign n12827 = ~n466 & ~n496;
  assign n12828 = ~n1478 & ~n1634;
  assign n12829 = n12827 & n12828;
  assign n12830 = ~n565 & ~n612;
  assign n12831 = n749 & n12830;
  assign n12832 = n749 & ~n1478;
  assign n12833 = ~n565 & n12832;
  assign n12834 = ~n612 & n12833;
  assign n12835 = ~n1634 & n12834;
  assign n12836 = ~n496 & n12835;
  assign n12837 = ~n466 & n12836;
  assign n12838 = n12828 & n12830;
  assign n12839 = n749 & n12827;
  assign n12840 = n12838 & n12839;
  assign n12841 = ~n466 & ~n612;
  assign n12842 = n12828 & n12841;
  assign n12843 = ~n496 & ~n565;
  assign n12844 = n749 & n12843;
  assign n12845 = n12842 & n12844;
  assign n12846 = ~n466 & ~n1478;
  assign n12847 = n12843 & n12846;
  assign n12848 = ~n612 & ~n1634;
  assign n12849 = n749 & n12848;
  assign n12850 = n12847 & n12849;
  assign n12851 = n12829 & n12831;
  assign n12852 = n772 & n1273;
  assign n12853 = n4587 & n6806;
  assign n12854 = n12852 & n12853;
  assign n12855 = n54550 & n12854;
  assign n12856 = n772 & n6806;
  assign n12857 = n12819 & n12856;
  assign n12858 = n53766 & n54360;
  assign n12859 = n12857 & n12858;
  assign n12860 = n4530 & n4587;
  assign n12861 = n1273 & n5021;
  assign n12862 = n12860 & n12861;
  assign n12863 = n54550 & n12862;
  assign n12864 = n12859 & n12863;
  assign n12865 = n54549 & n12855;
  assign n12866 = n54550 & n12858;
  assign n12867 = n6806 & n12866;
  assign n12868 = n54548 & n12867;
  assign n12869 = n1273 & n12868;
  assign n12870 = n772 & n12869;
  assign n12871 = n4530 & n12870;
  assign n12872 = n5021 & n12871;
  assign n12873 = n4587 & n12872;
  assign n12874 = ~n491 & n12873;
  assign n12875 = ~n344 & n12874;
  assign n12876 = ~n1769 & n12875;
  assign n12877 = n54548 & n54551;
  assign n12878 = ~n271 & ~n1034;
  assign n12879 = ~n271 & ~n883;
  assign n12880 = ~n1034 & n12879;
  assign n12881 = ~n883 & ~n1034;
  assign n12882 = ~n271 & n12881;
  assign n12883 = ~n883 & n12878;
  assign n12884 = ~n144 & ~n211;
  assign n12885 = ~n144 & ~n735;
  assign n12886 = ~n211 & n12885;
  assign n12887 = ~n735 & n12884;
  assign n12888 = n53673 & n54554;
  assign n12889 = n54553 & n12888;
  assign n12890 = n3672 & n5113;
  assign n12891 = n5956 & n11428;
  assign n12892 = n12890 & n12891;
  assign n12893 = n54134 & n12892;
  assign n12894 = n12889 & n12893;
  assign n12895 = n53835 & n54197;
  assign n12896 = n12894 & n12895;
  assign n12897 = n54552 & n12896;
  assign n12898 = n5956 & n54553;
  assign n12899 = n54134 & n12898;
  assign n12900 = n53835 & n12899;
  assign n12901 = n54197 & n12900;
  assign n12902 = n54552 & n12901;
  assign n12903 = n54546 & n12902;
  assign n12904 = n53673 & n12903;
  assign n12905 = n11428 & n12904;
  assign n12906 = n5113 & n12905;
  assign n12907 = n3672 & n12906;
  assign n12908 = ~n144 & n12907;
  assign n12909 = ~n211 & n12908;
  assign n12910 = ~n735 & n12909;
  assign n12911 = n54546 & n12896;
  assign n12912 = n54552 & n12911;
  assign n12913 = n54546 & n12897;
  assign n12914 = n54495 & ~n54555;
  assign n12915 = ~n54495 & n54555;
  assign n12916 = ~n12914 & ~n12915;
  assign n12917 = n10498 & ~n10500;
  assign n12918 = ~n10501 & ~n12917;
  assign n12919 = n1576 & n12918;
  assign n12920 = ~n53860 & n10564;
  assign n12921 = ~n53888 & n54403;
  assign n12922 = ~n53845 & n11215;
  assign n12923 = ~n12921 & ~n12922;
  assign n12924 = ~n12920 & ~n12921;
  assign n12925 = ~n12922 & n12924;
  assign n12926 = ~n12920 & n12923;
  assign n12927 = ~n12919 & n54556;
  assign n12928 = ~n12914 & ~n12927;
  assign n12929 = ~n12915 & n12928;
  assign n12930 = n12916 & ~n12927;
  assign n12931 = ~n12914 & ~n54557;
  assign n12932 = ~pi20  & ~n54515;
  assign n12933 = ~n12541 & n12546;
  assign n12934 = ~n12932 & ~n12933;
  assign n12935 = ~n12931 & ~n12934;
  assign n12936 = n12931 & n12934;
  assign n12937 = n10502 & ~n10504;
  assign n12938 = ~n10505 & ~n12937;
  assign n12939 = n1576 & n12938;
  assign n12940 = ~n53819 & n11215;
  assign n12941 = ~n53860 & n54403;
  assign n12942 = ~n53845 & n10564;
  assign n12943 = ~n12941 & ~n12942;
  assign n12944 = ~n12940 & ~n12941;
  assign n12945 = ~n12942 & n12944;
  assign n12946 = ~n12940 & n12943;
  assign n12947 = ~n12939 & n54558;
  assign n12948 = ~n12936 & ~n12947;
  assign n12949 = ~n12935 & ~n12936;
  assign n12950 = ~n12947 & n12949;
  assign n12951 = ~n12935 & ~n12950;
  assign n12952 = ~n12935 & ~n12948;
  assign n12953 = n12559 & ~n12563;
  assign n12954 = ~n12559 & ~n12564;
  assign n12955 = n12563 & ~n12564;
  assign n12956 = ~n12954 & ~n12955;
  assign n12957 = ~n12564 & ~n12953;
  assign n12958 = ~n54559 & ~n54560;
  assign n12959 = n54559 & n54560;
  assign n12960 = ~n12958 & ~n12959;
  assign n12961 = n11279 & n11889;
  assign n12962 = ~n53712 & n12584;
  assign n12963 = ~n53774 & n54410;
  assign n12964 = ~n53741 & n11267;
  assign n12965 = ~n12963 & ~n12964;
  assign n12966 = ~n12962 & ~n12963;
  assign n12967 = ~n12964 & n12966;
  assign n12968 = ~n12962 & n12965;
  assign n12969 = ~n11279 & n54561;
  assign n12970 = ~n11889 & n54561;
  assign n12971 = ~n12969 & ~n12970;
  assign n12972 = ~n12961 & n54561;
  assign n12973 = pi29  & ~n54562;
  assign n12974 = ~pi29  & n54562;
  assign n12975 = ~n12973 & ~n12974;
  assign n12976 = n12960 & ~n12975;
  assign n12977 = ~n12958 & ~n12976;
  assign n12978 = n54537 & n54538;
  assign n12979 = ~n54537 & ~n12701;
  assign n12980 = ~n54537 & n54538;
  assign n12981 = ~n54538 & ~n12701;
  assign n12982 = n54537 & ~n54538;
  assign n12983 = ~n54563 & ~n54564;
  assign n12984 = ~n12701 & ~n12978;
  assign n12985 = ~n12977 & ~n54565;
  assign n12986 = ~n12701 & ~n12985;
  assign n12987 = n12570 & ~n12572;
  assign n12988 = ~n12573 & ~n12987;
  assign n12989 = n12986 & ~n12988;
  assign n12990 = ~n12986 & n12988;
  assign n12991 = n11279 & n11380;
  assign n12992 = ~n53685 & n11267;
  assign n12993 = ~n53657 & n12584;
  assign n12994 = ~n53712 & n54410;
  assign n12995 = ~n12993 & ~n12994;
  assign n12996 = ~n12992 & ~n12994;
  assign n12997 = ~n12993 & n12996;
  assign n12998 = ~n12992 & n12995;
  assign n12999 = ~n12991 & n54566;
  assign n13000 = pi29  & ~n12999;
  assign n13001 = pi29  & ~n13000;
  assign n13002 = pi29  & n12999;
  assign n13003 = ~n12999 & ~n13000;
  assign n13004 = ~pi29  & ~n12999;
  assign n13005 = ~n54567 & ~n54568;
  assign n13006 = ~n12990 & n13005;
  assign n13007 = ~n12989 & ~n12990;
  assign n13008 = ~n13005 & n13007;
  assign n13009 = ~n12990 & ~n13008;
  assign n13010 = ~n12989 & ~n13006;
  assign n13011 = n12683 & ~n54569;
  assign n13012 = n123 & n54351;
  assign n13013 = n53444 & ~n53634;
  assign n13014 = n127 & ~n2325;
  assign n13015 = ~n13013 & ~n13014;
  assign n13016 = ~n13012 & n13015;
  assign n13017 = pi26  & ~n13016;
  assign n13018 = ~n13016 & ~n13017;
  assign n13019 = ~pi26  & ~n13016;
  assign n13020 = pi26  & ~n13017;
  assign n13021 = pi26  & n13016;
  assign n13022 = ~n54570 & ~n54571;
  assign n13023 = ~n12683 & n54569;
  assign n13024 = ~n54569 & ~n13011;
  assign n13025 = n12683 & ~n13011;
  assign n13026 = ~n13024 & ~n13025;
  assign n13027 = ~n13011 & ~n13023;
  assign n13028 = ~n13022 & ~n54572;
  assign n13029 = ~n13011 & ~n13028;
  assign n13030 = ~n12668 & n54535;
  assign n13031 = ~n12674 & ~n13030;
  assign n13032 = ~n13029 & n13031;
  assign n13033 = n123 & n11242;
  assign n13034 = n53444 & ~n53650;
  assign n13035 = n128 & ~n2325;
  assign n13036 = n127 & ~n53634;
  assign n13037 = ~n13035 & ~n13036;
  assign n13038 = ~n13034 & ~n13036;
  assign n13039 = ~n13035 & n13038;
  assign n13040 = ~n13034 & n13037;
  assign n13041 = ~n123 & n54573;
  assign n13042 = ~n11242 & n54573;
  assign n13043 = ~n13041 & ~n13042;
  assign n13044 = ~n13033 & n54573;
  assign n13045 = pi26  & ~n54574;
  assign n13046 = ~pi26  & n54574;
  assign n13047 = ~n13045 & ~n13046;
  assign n13048 = n11279 & n11360;
  assign n13049 = ~n53685 & n12584;
  assign n13050 = ~n53741 & n54410;
  assign n13051 = ~n53712 & n11267;
  assign n13052 = ~n13050 & ~n13051;
  assign n13053 = ~n13049 & ~n13050;
  assign n13054 = ~n13051 & n13053;
  assign n13055 = ~n13049 & n13052;
  assign n13056 = ~n11279 & n54575;
  assign n13057 = ~n11360 & n54575;
  assign n13058 = ~n13056 & ~n13057;
  assign n13059 = ~n13048 & n54575;
  assign n13060 = pi29  & ~n54576;
  assign n13061 = ~pi29  & n54576;
  assign n13062 = ~n13060 & ~n13061;
  assign n13063 = n12977 & n54565;
  assign n13064 = ~n12977 & ~n12985;
  assign n13065 = ~n54565 & ~n12985;
  assign n13066 = ~n13064 & ~n13065;
  assign n13067 = ~n12985 & ~n13063;
  assign n13068 = n13062 & n54577;
  assign n13069 = ~n13062 & ~n54577;
  assign n13070 = n123 & n11286;
  assign n13071 = n127 & ~n53650;
  assign n13072 = n53444 & ~n53657;
  assign n13073 = n128 & ~n53634;
  assign n13074 = ~n13072 & ~n13073;
  assign n13075 = ~n13071 & ~n13072;
  assign n13076 = ~n13073 & n13075;
  assign n13077 = ~n13071 & n13074;
  assign n13078 = ~n13070 & n54578;
  assign n13079 = pi26  & ~n13078;
  assign n13080 = pi26  & ~n13079;
  assign n13081 = pi26  & n13078;
  assign n13082 = ~n13078 & ~n13079;
  assign n13083 = ~pi26  & ~n13078;
  assign n13084 = ~n54579 & ~n54580;
  assign n13085 = ~n13069 & n13084;
  assign n13086 = ~n13068 & ~n13069;
  assign n13087 = ~n13084 & n13086;
  assign n13088 = ~n13069 & ~n13087;
  assign n13089 = ~n13068 & ~n13085;
  assign n13090 = ~n13047 & ~n54581;
  assign n13091 = n13047 & n54581;
  assign n13092 = ~n54581 & ~n13090;
  assign n13093 = n13047 & ~n54581;
  assign n13094 = ~n13047 & ~n13090;
  assign n13095 = ~n13047 & n54581;
  assign n13096 = ~n54582 & ~n54583;
  assign n13097 = ~n13090 & ~n13091;
  assign n13098 = n13007 & ~n13008;
  assign n13099 = n13005 & n13007;
  assign n13100 = ~n13005 & ~n13008;
  assign n13101 = ~n13005 & ~n13007;
  assign n13102 = ~n54585 & ~n54586;
  assign n13103 = ~n54584 & ~n13102;
  assign n13104 = ~n13090 & ~n13103;
  assign n13105 = n13022 & ~n13025;
  assign n13106 = ~n13024 & n13105;
  assign n13107 = n13022 & n54572;
  assign n13108 = ~n13028 & ~n54587;
  assign n13109 = ~n13104 & n13108;
  assign n13110 = ~n54583 & n13102;
  assign n13111 = ~n54582 & n13110;
  assign n13112 = ~n54582 & n13102;
  assign n13113 = ~n54583 & n13112;
  assign n13114 = n54584 & n13102;
  assign n13115 = ~n13103 & ~n54588;
  assign n13116 = n11279 & n11913;
  assign n13117 = ~n53774 & n11267;
  assign n13118 = ~n53799 & n54410;
  assign n13119 = ~n53741 & n12584;
  assign n13120 = ~n13118 & ~n13119;
  assign n13121 = ~n13117 & ~n13118;
  assign n13122 = ~n13119 & n13121;
  assign n13123 = ~n13117 & n13120;
  assign n13124 = ~n13116 & n54589;
  assign n13125 = pi29  & ~n13124;
  assign n13126 = ~n13124 & ~n13125;
  assign n13127 = ~pi29  & ~n13124;
  assign n13128 = pi29  & ~n13125;
  assign n13129 = pi29  & n13124;
  assign n13130 = ~n54590 & ~n54591;
  assign n13131 = n12947 & ~n12949;
  assign n13132 = ~n12947 & ~n12950;
  assign n13133 = n12949 & ~n12950;
  assign n13134 = ~n13132 & ~n13133;
  assign n13135 = ~n12950 & ~n13131;
  assign n13136 = ~n13130 & ~n54592;
  assign n13137 = ~n12916 & n12927;
  assign n13138 = ~n12927 & ~n54557;
  assign n13139 = ~n12915 & n12931;
  assign n13140 = ~n13138 & ~n13139;
  assign n13141 = ~n54557 & ~n13137;
  assign n13142 = n2333 & n3716;
  assign n13143 = n4314 & n4587;
  assign n13144 = n13142 & n13143;
  assign n13145 = ~n308 & ~n628;
  assign n13146 = ~n628 & ~n1062;
  assign n13147 = ~n308 & n13146;
  assign n13148 = ~n255 & n13147;
  assign n13149 = ~n255 & ~n308;
  assign n13150 = n13146 & n13149;
  assign n13151 = n8635 & n13145;
  assign n13152 = ~n272 & ~n567;
  assign n13153 = ~n340 & ~n956;
  assign n13154 = ~n340 & ~n567;
  assign n13155 = ~n272 & ~n956;
  assign n13156 = n13154 & n13155;
  assign n13157 = ~n272 & ~n340;
  assign n13158 = ~n567 & ~n956;
  assign n13159 = n13157 & n13158;
  assign n13160 = n13152 & n13153;
  assign n13161 = n54594 & n54595;
  assign n13162 = n13144 & n13161;
  assign n13163 = n1067 & n5362;
  assign n13164 = ~n211 & ~n553;
  assign n13165 = n8754 & n13164;
  assign n13166 = n13163 & n13165;
  assign n13167 = n53778 & n13166;
  assign n13168 = n4587 & n8754;
  assign n13169 = n13142 & n13168;
  assign n13170 = n13161 & n13169;
  assign n13171 = n4314 & n5362;
  assign n13172 = n1067 & n13164;
  assign n13173 = n13171 & n13172;
  assign n13174 = n53778 & n13173;
  assign n13175 = n13170 & n13174;
  assign n13176 = n1067 & n4314;
  assign n13177 = n3716 & n4587;
  assign n13178 = n13176 & n13177;
  assign n13179 = n13161 & n13178;
  assign n13180 = n2333 & n5362;
  assign n13181 = n13165 & n13180;
  assign n13182 = n53778 & n13181;
  assign n13183 = n13179 & n13182;
  assign n13184 = n13162 & n13167;
  assign n13185 = n54211 & n54596;
  assign n13186 = n53538 & n54257;
  assign n13187 = n13185 & n13186;
  assign n13188 = n2333 & n4314;
  assign n13189 = n3716 & n13188;
  assign n13190 = n8754 & n13189;
  assign n13191 = n54594 & n13190;
  assign n13192 = n53778 & n13191;
  assign n13193 = n5362 & n13192;
  assign n13194 = n54211 & n13193;
  assign n13195 = n53693 & n13194;
  assign n13196 = n53538 & n13195;
  assign n13197 = n54257 & n13196;
  assign n13198 = n1067 & n13197;
  assign n13199 = n4587 & n13198;
  assign n13200 = n13164 & n13199;
  assign n13201 = ~n567 & n13200;
  assign n13202 = ~n272 & n13201;
  assign n13203 = ~n956 & n13202;
  assign n13204 = ~n340 & n13203;
  assign n13205 = n53693 & n13187;
  assign n13206 = ~n211 & ~n984;
  assign n13207 = n2693 & n13206;
  assign n13208 = n2896 & n3082;
  assign n13209 = n13207 & n13208;
  assign n13210 = ~n218 & ~n554;
  assign n13211 = ~n218 & n2949;
  assign n13212 = ~n554 & n13211;
  assign n13213 = n2949 & n13210;
  assign n13214 = n3011 & n54598;
  assign n13215 = n13209 & n13214;
  assign n13216 = n5058 & n7275;
  assign n13217 = ~n174 & ~n340;
  assign n13218 = n12793 & n13217;
  assign n13219 = n13216 & n13218;
  assign n13220 = n53984 & n13219;
  assign n13221 = ~n493 & ~n496;
  assign n13222 = ~n507 & ~n830;
  assign n13223 = ~n496 & ~n507;
  assign n13224 = ~n493 & ~n830;
  assign n13225 = n13223 & n13224;
  assign n13226 = ~n493 & ~n507;
  assign n13227 = ~n496 & ~n830;
  assign n13228 = n13226 & n13227;
  assign n13229 = n13221 & n13222;
  assign n13230 = ~n553 & ~n788;
  assign n13231 = n5952 & n13230;
  assign n13232 = ~n553 & n5952;
  assign n13233 = ~n493 & n13232;
  assign n13234 = ~n830 & n13233;
  assign n13235 = ~n496 & n13234;
  assign n13236 = ~n507 & n13235;
  assign n13237 = ~n788 & n13236;
  assign n13238 = n54599 & n13231;
  assign n13239 = ~n414 & ~n1912;
  assign n13240 = n1672 & n13239;
  assign n13241 = n586 & n1672;
  assign n13242 = ~n414 & n13241;
  assign n13243 = ~n1912 & n13242;
  assign n13244 = n586 & n13240;
  assign n13245 = n54600 & n54601;
  assign n13246 = n13220 & n13245;
  assign n13247 = n5058 & n13214;
  assign n13248 = n7275 & n13247;
  assign n13249 = n54601 & n13248;
  assign n13250 = n54600 & n13249;
  assign n13251 = n3082 & n13250;
  assign n13252 = n53984 & n13251;
  assign n13253 = n2693 & n13252;
  assign n13254 = ~n984 & n13253;
  assign n13255 = ~n179 & n13254;
  assign n13256 = ~n174 & n13255;
  assign n13257 = ~n211 & n13256;
  assign n13258 = ~n216 & n13257;
  assign n13259 = ~n849 & n13258;
  assign n13260 = ~n420 & n13259;
  assign n13261 = ~n340 & n13260;
  assign n13262 = n2896 & n12793;
  assign n13263 = n13206 & n13217;
  assign n13264 = n13262 & n13263;
  assign n13265 = n13214 & n13264;
  assign n13266 = n3082 & n5058;
  assign n13267 = n2693 & n7275;
  assign n13268 = n13266 & n13267;
  assign n13269 = n53984 & n13268;
  assign n13270 = n13245 & n13269;
  assign n13271 = n13265 & n13270;
  assign n13272 = n13215 & n13246;
  assign n13273 = ~n405 & ~n419;
  assign n13274 = ~n883 & ~n1062;
  assign n13275 = n13273 & n13274;
  assign n13276 = n53809 & n13275;
  assign n13277 = ~n503 & ~n591;
  assign n13278 = ~n591 & n4381;
  assign n13279 = ~n503 & n13278;
  assign n13280 = n4381 & n13277;
  assign n13281 = n53602 & n54603;
  assign n13282 = n13276 & n13281;
  assign n13283 = n2152 & n7044;
  assign n13284 = n8929 & n13283;
  assign n13285 = n1091 & n1659;
  assign n13286 = n5639 & n6620;
  assign n13287 = n13285 & n13286;
  assign n13288 = n6620 & n7044;
  assign n13289 = n8929 & n13288;
  assign n13290 = n2152 & n5639;
  assign n13291 = n13285 & n13290;
  assign n13292 = n13289 & n13291;
  assign n13293 = n13284 & n13287;
  assign n13294 = n53459 & n54604;
  assign n13295 = ~n883 & ~n1485;
  assign n13296 = n13273 & n13295;
  assign n13297 = n53809 & n13296;
  assign n13298 = n13281 & n13297;
  assign n13299 = n8929 & n13290;
  assign n13300 = ~n249 & ~n1062;
  assign n13301 = n7044 & n13300;
  assign n13302 = n13285 & n13301;
  assign n13303 = n13299 & n13302;
  assign n13304 = n53459 & n13303;
  assign n13305 = n13298 & n13304;
  assign n13306 = n13282 & n13294;
  assign n13307 = n54602 & n54605;
  assign n13308 = n8929 & n13281;
  assign n13309 = n53754 & n13308;
  assign n13310 = n54602 & n13309;
  assign n13311 = n53459 & n13310;
  assign n13312 = n1091 & n13311;
  assign n13313 = n53809 & n13312;
  assign n13314 = n1659 & n13313;
  assign n13315 = n5639 & n13314;
  assign n13316 = ~n883 & n13315;
  assign n13317 = ~n1062 & n13316;
  assign n13318 = ~n1485 & n13317;
  assign n13319 = ~n567 & n13318;
  assign n13320 = ~n249 & n13319;
  assign n13321 = n2152 & n13320;
  assign n13322 = ~n405 & n13321;
  assign n13323 = ~n1034 & n13322;
  assign n13324 = ~n419 & n13323;
  assign n13325 = n53754 & n13307;
  assign n13326 = ~n54597 & ~n54606;
  assign n13327 = n54597 & n54606;
  assign n13328 = ~pi17  & ~n13326;
  assign n13329 = ~n13326 & ~n13327;
  assign n13330 = ~pi17  & n13329;
  assign n13331 = ~n13327 & n13328;
  assign n13332 = ~n13326 & ~n54607;
  assign n13333 = n54495 & ~n13332;
  assign n13334 = ~n54495 & n13332;
  assign n13335 = n10494 & ~n10496;
  assign n13336 = ~n10497 & ~n13335;
  assign n13337 = n1576 & n13336;
  assign n13338 = ~n53888 & n10564;
  assign n13339 = ~n53907 & n54403;
  assign n13340 = ~n53860 & n11215;
  assign n13341 = ~n13339 & ~n13340;
  assign n13342 = ~n13338 & ~n13339;
  assign n13343 = ~n13340 & n13342;
  assign n13344 = ~n13338 & n13341;
  assign n13345 = ~n13337 & n54608;
  assign n13346 = ~n13334 & ~n13345;
  assign n13347 = ~n13333 & n13345;
  assign n13348 = ~n13334 & ~n13347;
  assign n13349 = ~n13333 & ~n13334;
  assign n13350 = ~n13345 & n13349;
  assign n13351 = ~n13333 & ~n13350;
  assign n13352 = ~n13333 & ~n13346;
  assign n13353 = ~n54593 & n54609;
  assign n13354 = n54593 & ~n54609;
  assign n13355 = ~n13353 & ~n13354;
  assign n13356 = ~pi17  & ~n54607;
  assign n13357 = ~n13327 & n13332;
  assign n13358 = ~n13356 & ~n13357;
  assign n13359 = n10490 & ~n10492;
  assign n13360 = ~n10493 & ~n13359;
  assign n13361 = n1576 & n13360;
  assign n13362 = ~n53930 & n54403;
  assign n13363 = ~n53907 & n10564;
  assign n13364 = ~n53888 & n11215;
  assign n13365 = ~n13363 & ~n13364;
  assign n13366 = ~n13362 & ~n13363;
  assign n13367 = ~n13364 & n13366;
  assign n13368 = ~n13362 & n13365;
  assign n13369 = ~n13361 & ~n13362;
  assign n13370 = ~n13363 & n13369;
  assign n13371 = ~n13364 & n13370;
  assign n13372 = ~n13361 & n54610;
  assign n13373 = ~n13358 & ~n54611;
  assign n13374 = n586 & n8679;
  assign n13375 = ~n405 & ~n751;
  assign n13376 = n1955 & n13375;
  assign n13377 = n13374 & n13376;
  assign n13378 = n53833 & n13377;
  assign n13379 = n54225 & n13378;
  assign n13380 = ~n346 & ~n560;
  assign n13381 = ~n754 & ~n1088;
  assign n13382 = n13380 & n13381;
  assign n13383 = n5323 & n6322;
  assign n13384 = n13382 & n13383;
  assign n13385 = n53518 & n13384;
  assign n13386 = n54330 & n13385;
  assign n13387 = n586 & n5323;
  assign n13388 = n8679 & n13375;
  assign n13389 = n13387 & n13388;
  assign n13390 = n53833 & n13389;
  assign n13391 = n54225 & n13390;
  assign n13392 = ~n560 & ~n823;
  assign n13393 = ~n346 & ~n1088;
  assign n13394 = n13392 & n13393;
  assign n13395 = ~n451 & ~n754;
  assign n13396 = n1955 & n13395;
  assign n13397 = n13394 & n13396;
  assign n13398 = n53518 & n13397;
  assign n13399 = n54330 & n13398;
  assign n13400 = n13391 & n13399;
  assign n13401 = ~n161 & ~n560;
  assign n13402 = n586 & n13401;
  assign n13403 = n1955 & n8679;
  assign n13404 = n13402 & n13403;
  assign n13405 = n53833 & n13404;
  assign n13406 = n54225 & n13405;
  assign n13407 = ~n405 & ~n1088;
  assign n13408 = ~n754 & ~n823;
  assign n13409 = n13407 & n13408;
  assign n13410 = ~n553 & ~n751;
  assign n13411 = n3296 & n13410;
  assign n13412 = n13409 & n13411;
  assign n13413 = n53518 & n13412;
  assign n13414 = n54330 & n13413;
  assign n13415 = n13406 & n13414;
  assign n13416 = n13379 & n13386;
  assign n13417 = ~n773 & ~n1189;
  assign n13418 = ~n1189 & n9510;
  assign n13419 = ~n773 & n13418;
  assign n13420 = n9510 & n13417;
  assign n13421 = ~n144 & ~n513;
  assign n13422 = n1197 & n13421;
  assign n13423 = n1076 & n3389;
  assign n13424 = n13422 & n13423;
  assign n13425 = n54613 & n13424;
  assign n13426 = n1043 & n1653;
  assign n13427 = ~n404 & ~n879;
  assign n13428 = ~n984 & ~n1477;
  assign n13429 = n13427 & n13428;
  assign n13430 = n13426 & n13429;
  assign n13431 = n54159 & n13430;
  assign n13432 = n1653 & n54613;
  assign n13433 = n1076 & n13432;
  assign n13434 = n54159 & n13433;
  assign n13435 = n1197 & n13434;
  assign n13436 = n3389 & n13435;
  assign n13437 = ~n984 & n13436;
  assign n13438 = ~n879 & n13437;
  assign n13439 = ~n1477 & n13438;
  assign n13440 = ~n144 & n13439;
  assign n13441 = ~n404 & n13440;
  assign n13442 = ~n1042 & n13441;
  assign n13443 = ~n587 & n13442;
  assign n13444 = ~n513 & n13443;
  assign n13445 = n1653 & n13421;
  assign n13446 = n1197 & n3389;
  assign n13447 = n13445 & n13446;
  assign n13448 = n54613 & n13447;
  assign n13449 = n1043 & n1076;
  assign n13450 = n13429 & n13449;
  assign n13451 = n54159 & n13450;
  assign n13452 = n13448 & n13451;
  assign n13453 = ~n513 & ~n1042;
  assign n13454 = ~n144 & ~n587;
  assign n13455 = n13453 & n13454;
  assign n13456 = n1197 & n13427;
  assign n13457 = n13455 & n13456;
  assign n13458 = n54613 & n13457;
  assign n13459 = n1653 & n13428;
  assign n13460 = n13423 & n13459;
  assign n13461 = n54159 & n13460;
  assign n13462 = n13458 & n13461;
  assign n13463 = ~n587 & ~n879;
  assign n13464 = ~n144 & ~n1042;
  assign n13465 = n13463 & n13464;
  assign n13466 = ~n513 & ~n1477;
  assign n13467 = ~n404 & ~n984;
  assign n13468 = n13466 & n13467;
  assign n13469 = n13465 & n13468;
  assign n13470 = n54613 & n13469;
  assign n13471 = n1197 & n1653;
  assign n13472 = n13423 & n13471;
  assign n13473 = n54159 & n13472;
  assign n13474 = n13470 & n13473;
  assign n13475 = n13425 & n13431;
  assign n13476 = ~n590 & n5652;
  assign n13477 = n613 & n3878;
  assign n13478 = n4975 & n13477;
  assign n13479 = ~n590 & n3878;
  assign n13480 = n613 & n4975;
  assign n13481 = n5652 & n13480;
  assign n13482 = n13479 & n13481;
  assign n13483 = ~n590 & n4975;
  assign n13484 = n3878 & n5652;
  assign n13485 = n613 & n13484;
  assign n13486 = n13483 & n13485;
  assign n13487 = n13476 & n13478;
  assign n13488 = n613 & n54260;
  assign n13489 = n5652 & n13488;
  assign n13490 = n3878 & n13489;
  assign n13491 = ~n741 & n13490;
  assign n13492 = ~n622 & n13491;
  assign n13493 = ~n590 & n13492;
  assign n13494 = n54260 & n54615;
  assign n13495 = n54614 & n54616;
  assign n13496 = n54612 & n13495;
  assign n13497 = n53833 & n8679;
  assign n13498 = n54225 & n13497;
  assign n13499 = n1955 & n13498;
  assign n13500 = n54614 & n13499;
  assign n13501 = n54359 & n13500;
  assign n13502 = n54616 & n13501;
  assign n13503 = n53518 & n13502;
  assign n13504 = n54330 & n13503;
  assign n13505 = n586 & n13504;
  assign n13506 = ~n1088 & n13505;
  assign n13507 = ~n161 & n13506;
  assign n13508 = ~n560 & n13507;
  assign n13509 = ~n405 & n13508;
  assign n13510 = ~n553 & n13509;
  assign n13511 = ~n823 & n13510;
  assign n13512 = ~n451 & n13511;
  assign n13513 = ~n754 & n13512;
  assign n13514 = ~n751 & n13513;
  assign n13515 = ~n346 & n13514;
  assign n13516 = n54359 & n13496;
  assign n13517 = n54597 & ~n54617;
  assign n13518 = ~n54597 & n54617;
  assign n13519 = ~n13517 & ~n13518;
  assign n13520 = ~n207 & ~n564;
  assign n13521 = ~n207 & ~n222;
  assign n13522 = ~n564 & n13521;
  assign n13523 = ~n222 & n13520;
  assign n13524 = n3086 & n4092;
  assign n13525 = n54618 & n13524;
  assign n13526 = n54138 & n10239;
  assign n13527 = n13525 & n13526;
  assign n13528 = ~n625 & ~n914;
  assign n13529 = n4314 & n13528;
  assign n13530 = ~n258 & ~n1492;
  assign n13531 = n10640 & n13530;
  assign n13532 = n4314 & n13530;
  assign n13533 = ~n296 & n13532;
  assign n13534 = ~n218 & n13533;
  assign n13535 = ~n914 & n13534;
  assign n13536 = ~n625 & n13535;
  assign n13537 = ~n218 & ~n625;
  assign n13538 = ~n296 & ~n914;
  assign n13539 = n10640 & n13528;
  assign n13540 = n13537 & n13538;
  assign n13541 = n13532 & n54620;
  assign n13542 = n13529 & n13531;
  assign n13543 = ~n249 & ~n848;
  assign n13544 = n4832 & n13543;
  assign n13545 = ~n317 & ~n1471;
  assign n13546 = ~n249 & n13545;
  assign n13547 = ~n848 & n13546;
  assign n13548 = ~n460 & n13547;
  assign n13549 = ~n773 & n13548;
  assign n13550 = n5661 & n13544;
  assign n13551 = ~n496 & ~n1079;
  assign n13552 = n1091 & n6482;
  assign n13553 = n13551 & n13552;
  assign n13554 = n54621 & n13553;
  assign n13555 = n54619 & n13554;
  assign n13556 = n3086 & n6482;
  assign n13557 = n54618 & n13556;
  assign n13558 = n13526 & n13557;
  assign n13559 = n1091 & n4092;
  assign n13560 = n13551 & n13559;
  assign n13561 = n54621 & n13560;
  assign n13562 = n54619 & n13561;
  assign n13563 = n13558 & n13562;
  assign n13564 = ~n222 & ~n1079;
  assign n13565 = ~n496 & n13564;
  assign n13566 = ~n207 & ~n650;
  assign n13567 = ~n420 & ~n564;
  assign n13568 = n13566 & n13567;
  assign n13569 = n13565 & n13568;
  assign n13570 = n13526 & n13569;
  assign n13571 = n3086 & n13552;
  assign n13572 = n54619 & n13571;
  assign n13573 = n54621 & n13572;
  assign n13574 = n13570 & n13573;
  assign n13575 = n13527 & n13555;
  assign n13576 = n13526 & n54621;
  assign n13577 = n54616 & n13576;
  assign n13578 = n54619 & n13577;
  assign n13579 = n3086 & n13578;
  assign n13580 = n1091 & n13579;
  assign n13581 = n6482 & n13580;
  assign n13582 = ~n1079 & n13581;
  assign n13583 = ~n222 & n13582;
  assign n13584 = ~n207 & n13583;
  assign n13585 = ~n564 & n13584;
  assign n13586 = ~n496 & n13585;
  assign n13587 = ~n420 & n13586;
  assign n13588 = ~n650 & n13587;
  assign n13589 = n54616 & n54622;
  assign n13590 = ~n464 & ~n587;
  assign n13591 = ~n506 & n13590;
  assign n13592 = ~n357 & n13591;
  assign n13593 = ~n464 & ~n506;
  assign n13594 = ~n357 & ~n587;
  assign n13595 = n13593 & n13594;
  assign n13596 = n6302 & n13590;
  assign n13597 = ~n105 & ~n552;
  assign n13598 = ~n615 & n13597;
  assign n13599 = n54354 & n13598;
  assign n13600 = n54624 & n13599;
  assign n13601 = ~n216 & ~n219;
  assign n13602 = ~n353 & ~n461;
  assign n13603 = n13601 & n13602;
  assign n13604 = n417 & n13603;
  assign n13605 = ~n742 & ~n984;
  assign n13606 = ~n742 & ~n1486;
  assign n13607 = ~n984 & n13606;
  assign n13608 = ~n1486 & n13605;
  assign n13609 = n5690 & n54625;
  assign n13610 = n13604 & n13609;
  assign n13611 = n53769 & n54292;
  assign n13612 = n13610 & n13611;
  assign n13613 = n5690 & n54292;
  assign n13614 = n54354 & n13613;
  assign n13615 = n54624 & n13614;
  assign n13616 = n53769 & n13615;
  assign n13617 = n417 & n13616;
  assign n13618 = n13598 & n13617;
  assign n13619 = ~n984 & n13618;
  assign n13620 = ~n1486 & n13619;
  assign n13621 = ~n219 & n13620;
  assign n13622 = ~n216 & n13621;
  assign n13623 = ~n742 & n13622;
  assign n13624 = ~n461 & n13623;
  assign n13625 = ~n353 & n13624;
  assign n13626 = n5690 & n13598;
  assign n13627 = n54624 & n13626;
  assign n13628 = ~n219 & ~n461;
  assign n13629 = ~n216 & ~n1486;
  assign n13630 = n13628 & n13629;
  assign n13631 = n417 & n13630;
  assign n13632 = ~n353 & ~n742;
  assign n13633 = ~n984 & n13632;
  assign n13634 = n54354 & n13633;
  assign n13635 = n13631 & n13634;
  assign n13636 = n13611 & n13635;
  assign n13637 = n13627 & n13636;
  assign n13638 = n5690 & n54354;
  assign n13639 = n54624 & n13638;
  assign n13640 = ~n219 & ~n353;
  assign n13641 = n13605 & n13640;
  assign n13642 = n417 & n13641;
  assign n13643 = ~n216 & ~n461;
  assign n13644 = ~n1486 & n13643;
  assign n13645 = n13598 & n13644;
  assign n13646 = n13642 & n13645;
  assign n13647 = n13611 & n13646;
  assign n13648 = n13639 & n13647;
  assign n13649 = n13600 & n13612;
  assign n13650 = ~n405 & ~n441;
  assign n13651 = n7016 & n12730;
  assign n13652 = n13650 & n13651;
  assign n13653 = ~n1658 & ~n1680;
  assign n13654 = ~n269 & n13653;
  assign n13655 = ~n269 & ~n1680;
  assign n13656 = ~n1658 & n13655;
  assign n13657 = ~n1680 & n2579;
  assign n13658 = ~n211 & ~n259;
  assign n13659 = ~n307 & ~n1042;
  assign n13660 = n13658 & n13659;
  assign n13661 = ~n659 & ~n664;
  assign n13662 = n3523 & n13661;
  assign n13663 = n13660 & n13662;
  assign n13664 = n54627 & n13663;
  assign n13665 = n3523 & n54627;
  assign n13666 = n7016 & n13665;
  assign n13667 = ~n320 & n13666;
  assign n13668 = ~n659 & n13667;
  assign n13669 = ~n307 & n13668;
  assign n13670 = ~n211 & n13669;
  assign n13671 = ~n259 & n13670;
  assign n13672 = ~n664 & n13671;
  assign n13673 = ~n405 & n13672;
  assign n13674 = ~n1042 & n13673;
  assign n13675 = ~n441 & n13674;
  assign n13676 = ~n1644 & n13675;
  assign n13677 = n3523 & n7016;
  assign n13678 = n12730 & n13677;
  assign n13679 = ~n211 & ~n307;
  assign n13680 = n13661 & n13679;
  assign n13681 = ~n259 & ~n405;
  assign n13682 = ~n441 & ~n1042;
  assign n13683 = n13681 & n13682;
  assign n13684 = ~n405 & ~n1042;
  assign n13685 = n13658 & n13684;
  assign n13686 = ~n441 & ~n664;
  assign n13687 = ~n307 & ~n659;
  assign n13688 = n13686 & n13687;
  assign n13689 = n13685 & n13688;
  assign n13690 = n13680 & n13683;
  assign n13691 = n54627 & n54629;
  assign n13692 = n13678 & n13691;
  assign n13693 = ~n259 & ~n307;
  assign n13694 = n7016 & n13693;
  assign n13695 = n3523 & n13694;
  assign n13696 = ~n664 & ~n1042;
  assign n13697 = ~n320 & ~n405;
  assign n13698 = n13696 & n13697;
  assign n13699 = ~n211 & ~n659;
  assign n13700 = ~n441 & ~n1644;
  assign n13701 = n13699 & n13700;
  assign n13702 = n13698 & n13701;
  assign n13703 = n54627 & n13702;
  assign n13704 = n13695 & n13703;
  assign n13705 = n13652 & n13664;
  assign n13706 = ~n459 & ~n1715;
  assign n13707 = ~n459 & ~n1469;
  assign n13708 = ~n1715 & n13707;
  assign n13709 = ~n1469 & ~n1715;
  assign n13710 = ~n459 & n13709;
  assign n13711 = ~n1469 & n13706;
  assign n13712 = ~n177 & ~n364;
  assign n13713 = ~n177 & ~n1468;
  assign n13714 = ~n364 & n13713;
  assign n13715 = ~n364 & ~n1468;
  assign n13716 = ~n177 & n13715;
  assign n13717 = ~n1468 & n13712;
  assign n13718 = n293 & n8929;
  assign n13719 = n54631 & n13718;
  assign n13720 = n8929 & n54630;
  assign n13721 = n293 & n13720;
  assign n13722 = ~n1468 & n13721;
  assign n13723 = ~n177 & n13722;
  assign n13724 = ~n364 & n13723;
  assign n13725 = n54630 & n13719;
  assign n13726 = ~n294 & ~n410;
  assign n13727 = ~n788 & ~n2042;
  assign n13728 = n13726 & n13727;
  assign n13729 = n1197 & n3082;
  assign n13730 = n13728 & n13729;
  assign n13731 = ~n422 & ~n627;
  assign n13732 = ~n422 & ~n1535;
  assign n13733 = ~n627 & n13732;
  assign n13734 = ~n1535 & n13731;
  assign n13735 = n54192 & n54633;
  assign n13736 = n13730 & n13735;
  assign n13737 = ~n144 & ~n565;
  assign n13738 = ~n360 & ~n849;
  assign n13739 = n1128 & n13738;
  assign n13740 = n1128 & n13737;
  assign n13741 = n13738 & n13740;
  assign n13742 = n13737 & n13739;
  assign n13743 = n12208 & n54634;
  assign n13744 = n1128 & n1197;
  assign n13745 = n13728 & n13744;
  assign n13746 = n13735 & n13745;
  assign n13747 = n3082 & n13738;
  assign n13748 = n13737 & n13747;
  assign n13749 = n12208 & n13748;
  assign n13750 = n13746 & n13749;
  assign n13751 = ~n788 & ~n849;
  assign n13752 = ~n360 & ~n410;
  assign n13753 = n13751 & n13752;
  assign n13754 = ~n294 & ~n2042;
  assign n13755 = n3082 & n13754;
  assign n13756 = n13753 & n13755;
  assign n13757 = n13735 & n13756;
  assign n13758 = n13737 & n13744;
  assign n13759 = n12208 & n13758;
  assign n13760 = n13757 & n13759;
  assign n13761 = n13736 & n13743;
  assign n13762 = n54632 & n54635;
  assign n13763 = n54628 & n13762;
  assign n13764 = n54626 & n13763;
  assign n13765 = n12208 & n13737;
  assign n13766 = n54633 & n13765;
  assign n13767 = n54632 & n13766;
  assign n13768 = n1197 & n13767;
  assign n13769 = n54192 & n13768;
  assign n13770 = n54628 & n13769;
  assign n13771 = n54626 & n13770;
  assign n13772 = n54623 & n13771;
  assign n13773 = n3082 & n13772;
  assign n13774 = n1128 & n13773;
  assign n13775 = ~n294 & n13774;
  assign n13776 = ~n849 & n13775;
  assign n13777 = ~n360 & n13776;
  assign n13778 = ~n410 & n13777;
  assign n13779 = ~n788 & n13778;
  assign n13780 = ~n2042 & n13779;
  assign n13781 = n54623 & n13764;
  assign n13782 = n8824 & n10183;
  assign n13783 = n11134 & n13782;
  assign n13784 = ~n271 & ~n291;
  assign n13785 = ~n291 & ~n1090;
  assign n13786 = ~n271 & n13785;
  assign n13787 = ~n271 & ~n1090;
  assign n13788 = ~n291 & n13787;
  assign n13789 = ~n1090 & n13784;
  assign n13790 = n629 & n5361;
  assign n13791 = n54637 & n13790;
  assign n13792 = n54603 & n13791;
  assign n13793 = n5361 & n8824;
  assign n13794 = n54603 & n13793;
  assign n13795 = n629 & n13794;
  assign n13796 = n10183 & n13795;
  assign n13797 = n11134 & n13796;
  assign n13798 = ~n291 & n13797;
  assign n13799 = ~n1090 & n13798;
  assign n13800 = ~n271 & n13799;
  assign n13801 = n10183 & n13793;
  assign n13802 = n629 & n11134;
  assign n13803 = n54637 & n13802;
  assign n13804 = n54603 & n13803;
  assign n13805 = n13801 & n13804;
  assign n13806 = n13783 & n13792;
  assign n13807 = ~n316 & ~n493;
  assign n13808 = n6205 & n6897;
  assign n13809 = n13807 & n13808;
  assign n13810 = ~n419 & ~n740;
  assign n13811 = ~n1088 & ~n1457;
  assign n13812 = n13810 & n13811;
  assign n13813 = ~n207 & ~n588;
  assign n13814 = n4470 & n13813;
  assign n13815 = ~n588 & ~n740;
  assign n13816 = n13811 & n13815;
  assign n13817 = ~n207 & ~n419;
  assign n13818 = n4470 & n13817;
  assign n13819 = n13816 & n13818;
  assign n13820 = n13812 & n13814;
  assign n13821 = n54613 & n54639;
  assign n13822 = n4470 & n6205;
  assign n13823 = n6897 & n13822;
  assign n13824 = n13807 & n13813;
  assign n13825 = n13812 & n13824;
  assign n13826 = n54613 & n13825;
  assign n13827 = n13823 & n13826;
  assign n13828 = n13809 & n13821;
  assign n13829 = n53708 & n54640;
  assign n13830 = n6205 & n54613;
  assign n13831 = n4470 & n13830;
  assign n13832 = n54638 & n13831;
  assign n13833 = n53708 & n13832;
  assign n13834 = n6897 & n13833;
  assign n13835 = ~n1088 & n13834;
  assign n13836 = ~n316 & n13835;
  assign n13837 = ~n207 & n13836;
  assign n13838 = ~n1457 & n13837;
  assign n13839 = ~n493 & n13838;
  assign n13840 = ~n419 & n13839;
  assign n13841 = ~n740 & n13840;
  assign n13842 = ~n588 & n13841;
  assign n13843 = n54638 & n13829;
  assign n13844 = ~n292 & ~n852;
  assign n13845 = ~n1468 & ~n1681;
  assign n13846 = n13844 & n13845;
  assign n13847 = ~n166 & ~n211;
  assign n13848 = n406 & n13847;
  assign n13849 = n2367 & n3675;
  assign n13850 = n13848 & n13849;
  assign n13851 = n13846 & n13850;
  assign n13852 = ~n295 & ~n615;
  assign n13853 = n5198 & n7513;
  assign n13854 = n13852 & n13853;
  assign n13855 = n54232 & n13854;
  assign n13856 = ~n751 & n9051;
  assign n13857 = n355 & n3214;
  assign n13858 = n54550 & n54642;
  assign n13859 = n13855 & n13858;
  assign n13860 = n5198 & n54550;
  assign n13861 = n54232 & n13860;
  assign n13862 = n3675 & n13861;
  assign n13863 = n3214 & n13862;
  assign n13864 = n355 & n13863;
  assign n13865 = n406 & n13864;
  assign n13866 = n2367 & n13865;
  assign n13867 = ~n295 & n13866;
  assign n13868 = ~n957 & n13867;
  assign n13869 = ~n1681 & n13868;
  assign n13870 = ~n1468 & n13869;
  assign n13871 = ~n211 & n13870;
  assign n13872 = ~n292 & n13871;
  assign n13873 = ~n166 & n13872;
  assign n13874 = ~n852 & n13873;
  assign n13875 = ~n498 & n13874;
  assign n13876 = ~n615 & n13875;
  assign n13877 = ~n852 & ~n1468;
  assign n13878 = n2367 & n13877;
  assign n13879 = n406 & n3675;
  assign n13880 = n13878 & n13879;
  assign n13881 = ~n211 & ~n1681;
  assign n13882 = ~n166 & ~n292;
  assign n13883 = n13881 & n13882;
  assign n13884 = n54642 & n13883;
  assign n13885 = ~n211 & ~n292;
  assign n13886 = n406 & n13885;
  assign n13887 = n13849 & n13886;
  assign n13888 = ~n166 & ~n852;
  assign n13889 = n13845 & n13888;
  assign n13890 = n54642 & n13889;
  assign n13891 = n13887 & n13890;
  assign n13892 = n13880 & n13884;
  assign n13893 = n54550 & n13855;
  assign n13894 = n54644 & n13893;
  assign n13895 = n2367 & n13852;
  assign n13896 = n3675 & n5198;
  assign n13897 = n13895 & n13896;
  assign n13898 = ~n498 & ~n1468;
  assign n13899 = ~n166 & ~n1681;
  assign n13900 = n13898 & n13899;
  assign n13901 = ~n211 & ~n852;
  assign n13902 = ~n292 & ~n957;
  assign n13903 = n13901 & n13902;
  assign n13904 = n13900 & n13903;
  assign n13905 = n13897 & n13904;
  assign n13906 = n355 & n406;
  assign n13907 = n3214 & n13906;
  assign n13908 = n54232 & n13907;
  assign n13909 = n54550 & n13908;
  assign n13910 = n13905 & n13909;
  assign n13911 = n13851 & n13859;
  assign n13912 = ~n851 & ~n922;
  assign n13913 = n5639 & n8452;
  assign n13914 = n13912 & n13913;
  assign n13915 = ~n215 & ~n268;
  assign n13916 = ~n163 & ~n901;
  assign n13917 = ~n163 & ~n215;
  assign n13918 = ~n268 & ~n901;
  assign n13919 = n13917 & n13918;
  assign n13920 = n13915 & n13916;
  assign n13921 = n53942 & n54645;
  assign n13922 = n54222 & n13921;
  assign n13923 = n53942 & n54222;
  assign n13924 = n13912 & n13923;
  assign n13925 = n5639 & n13924;
  assign n13926 = ~n1192 & n13925;
  assign n13927 = ~n901 & n13926;
  assign n13928 = ~n163 & n13927;
  assign n13929 = ~n112 & n13928;
  assign n13930 = ~n215 & n13929;
  assign n13931 = ~n268 & n13930;
  assign n13932 = n5639 & n13915;
  assign n13933 = n13912 & n13932;
  assign n13934 = ~n112 & ~n901;
  assign n13935 = ~n163 & ~n1192;
  assign n13936 = n13934 & n13935;
  assign n13937 = n53942 & n13936;
  assign n13938 = n54222 & n13937;
  assign n13939 = n13933 & n13938;
  assign n13940 = n13914 & n13922;
  assign n13941 = ~n415 & ~n1191;
  assign n13942 = ~n622 & n4791;
  assign n13943 = ~n415 & ~n622;
  assign n13944 = ~n1191 & n13943;
  assign n13945 = n4791 & n13944;
  assign n13946 = ~n1191 & n4791;
  assign n13947 = n13943 & n13946;
  assign n13948 = n13941 & n13942;
  assign n13949 = ~n415 & n54074;
  assign n13950 = ~n1191 & n13949;
  assign n13951 = ~n161 & n13950;
  assign n13952 = ~n622 & n13951;
  assign n13953 = ~n1912 & n13952;
  assign n13954 = n54074 & n54647;
  assign n13955 = n1078 & n6481;
  assign n13956 = n3015 & n53913;
  assign n13957 = n13955 & n13956;
  assign n13958 = ~n510 & ~n1465;
  assign n13959 = n3256 & n4378;
  assign n13960 = n13958 & n13959;
  assign n13961 = ~n511 & ~n618;
  assign n13962 = ~n883 & n13961;
  assign n13963 = n831 & n2537;
  assign n13964 = n13962 & n13963;
  assign n13965 = n2537 & n3256;
  assign n13966 = n4378 & n13965;
  assign n13967 = n512 & n831;
  assign n13968 = ~n618 & ~n883;
  assign n13969 = ~n1465 & n13968;
  assign n13970 = n13967 & n13969;
  assign n13971 = n13966 & n13970;
  assign n13972 = n512 & n2537;
  assign n13973 = n831 & n13972;
  assign n13974 = n2537 & n13967;
  assign n13975 = ~n883 & ~n1465;
  assign n13976 = ~n1031 & n13975;
  assign n13977 = ~n618 & ~n776;
  assign n13978 = n4378 & n13977;
  assign n13979 = n13976 & n13978;
  assign n13980 = n54650 & n13979;
  assign n13981 = n13960 & n13964;
  assign n13982 = ~n618 & n3256;
  assign n13983 = n53913 & n13982;
  assign n13984 = n3015 & n13983;
  assign n13985 = n4378 & n13975;
  assign n13986 = n13955 & n13985;
  assign n13987 = n54650 & n13986;
  assign n13988 = n13984 & n13987;
  assign n13989 = n13957 & n54649;
  assign n13990 = n54648 & n54651;
  assign n13991 = n54646 & n13990;
  assign n13992 = n54643 & n13991;
  assign n13993 = n831 & n3015;
  assign n13994 = n6481 & n13993;
  assign n13995 = n53913 & n13994;
  assign n13996 = n512 & n13995;
  assign n13997 = n54643 & n13996;
  assign n13998 = n54641 & n13997;
  assign n13999 = n54646 & n13998;
  assign n14000 = n54648 & n13999;
  assign n14001 = n1078 & n14000;
  assign n14002 = n2537 & n14001;
  assign n14003 = n4378 & n14002;
  assign n14004 = ~n1031 & n14003;
  assign n14005 = ~n883 & n14004;
  assign n14006 = ~n1465 & n14005;
  assign n14007 = ~n618 & n14006;
  assign n14008 = ~n776 & n14007;
  assign n14009 = n54641 & n13992;
  assign n14010 = ~n54636 & ~n54652;
  assign n14011 = n54636 & n54652;
  assign n14012 = ~pi14  & ~n14010;
  assign n14013 = ~n14010 & ~n14011;
  assign n14014 = ~pi14  & n14013;
  assign n14015 = ~n14011 & n14012;
  assign n14016 = ~n14010 & ~n54653;
  assign n14017 = n54617 & ~n14016;
  assign n14018 = ~n54617 & n14016;
  assign n14019 = n10482 & ~n10484;
  assign n14020 = ~n10485 & ~n14019;
  assign n14021 = n1576 & n14020;
  assign n14022 = ~n53962 & n10564;
  assign n14023 = ~n53970 & n54403;
  assign n14024 = ~n53930 & n11215;
  assign n14025 = ~n14023 & ~n14024;
  assign n14026 = ~n14022 & ~n14023;
  assign n14027 = ~n14024 & n14026;
  assign n14028 = ~n14022 & n14025;
  assign n14029 = ~n14021 & n54654;
  assign n14030 = ~n14018 & ~n14029;
  assign n14031 = ~n14017 & n14029;
  assign n14032 = ~n14018 & ~n14031;
  assign n14033 = ~n14017 & ~n14018;
  assign n14034 = ~n14029 & n14033;
  assign n14035 = ~n14017 & ~n14034;
  assign n14036 = ~n14017 & ~n14030;
  assign n14037 = ~n13517 & n54655;
  assign n14038 = ~n13518 & n14037;
  assign n14039 = n13519 & n54655;
  assign n14040 = ~n13517 & ~n54656;
  assign n14041 = n13358 & n54611;
  assign n14042 = ~n13373 & ~n14041;
  assign n14043 = ~n14040 & n14042;
  assign n14044 = ~n13373 & ~n14043;
  assign n14045 = n13345 & ~n13349;
  assign n14046 = ~n13345 & ~n13350;
  assign n14047 = n13349 & ~n13350;
  assign n14048 = ~n14046 & ~n14047;
  assign n14049 = ~n13350 & ~n14045;
  assign n14050 = ~n14044 & ~n54657;
  assign n14051 = n14044 & n54657;
  assign n14052 = ~n14050 & ~n14051;
  assign n14053 = n11279 & n12550;
  assign n14054 = ~n53819 & n11267;
  assign n14055 = ~n53845 & n54410;
  assign n14056 = ~n53799 & n12584;
  assign n14057 = ~n14055 & ~n14056;
  assign n14058 = ~n14054 & ~n14055;
  assign n14059 = ~n14056 & n14058;
  assign n14060 = ~n14054 & n14057;
  assign n14061 = ~n11279 & n54658;
  assign n14062 = ~n12550 & n54658;
  assign n14063 = ~n14061 & ~n14062;
  assign n14064 = ~n14053 & n54658;
  assign n14065 = pi29  & ~n54659;
  assign n14066 = ~pi29  & n54659;
  assign n14067 = ~n14065 & ~n14066;
  assign n14068 = n14052 & ~n14067;
  assign n14069 = ~n14050 & ~n14068;
  assign n14070 = n13355 & ~n14069;
  assign n14071 = ~n13353 & ~n14070;
  assign n14072 = n13130 & n54592;
  assign n14073 = ~n13130 & ~n13136;
  assign n14074 = ~n13130 & n54592;
  assign n14075 = ~n54592 & ~n13136;
  assign n14076 = n13130 & ~n54592;
  assign n14077 = ~n54660 & ~n54661;
  assign n14078 = ~n13136 & ~n14072;
  assign n14079 = ~n14071 & ~n54662;
  assign n14080 = ~n13136 & ~n14079;
  assign n14081 = ~n12960 & n12975;
  assign n14082 = ~n12976 & ~n14081;
  assign n14083 = ~n14080 & n14082;
  assign n14084 = n123 & n11213;
  assign n14085 = n128 & ~n53650;
  assign n14086 = n53444 & ~n53685;
  assign n14087 = n127 & ~n53657;
  assign n14088 = ~n14086 & ~n14087;
  assign n14089 = ~n14085 & n14088;
  assign n14090 = ~n14084 & n14089;
  assign n14091 = pi26  & ~n14090;
  assign n14092 = ~n14090 & ~n14091;
  assign n14093 = ~pi26  & ~n14090;
  assign n14094 = pi26  & ~n14091;
  assign n14095 = pi26  & n14090;
  assign n14096 = ~n54663 & ~n54664;
  assign n14097 = n14080 & ~n14082;
  assign n14098 = ~n14080 & ~n14083;
  assign n14099 = n14082 & ~n14083;
  assign n14100 = ~n14098 & ~n14099;
  assign n14101 = ~n14083 & ~n14097;
  assign n14102 = ~n14096 & ~n54665;
  assign n14103 = ~n14083 & ~n14102;
  assign n14104 = pi21  & ~pi22 ;
  assign n14105 = ~pi21  & pi22 ;
  assign n14106 = ~pi21  & ~pi22 ;
  assign n14107 = pi21  & pi22 ;
  assign n14108 = ~n14106 & ~n14107;
  assign n14109 = ~n14104 & ~n14105;
  assign n14110 = ~n53441 & ~n54666;
  assign n14111 = ~n53441 & n53442;
  assign n14112 = ~n54666 & n14111;
  assign n14113 = n53442 & n14110;
  assign n14114 = n90 & ~n10547;
  assign n14115 = ~n54667 & ~n14114;
  assign n14116 = ~n2325 & n54667;
  assign n14117 = ~n10551 & ~n14116;
  assign n14118 = ~n90 & ~n14116;
  assign n14119 = ~n14117 & ~n14118;
  assign n14120 = ~n2325 & ~n14115;
  assign n14121 = pi23  & ~n54668;
  assign n14122 = ~pi23  & n54668;
  assign n14123 = ~n14121 & ~n14122;
  assign n14124 = n14103 & n14123;
  assign n14125 = ~n14103 & ~n14123;
  assign n14126 = n13086 & ~n13087;
  assign n14127 = n13084 & n13086;
  assign n14128 = ~n13084 & ~n13087;
  assign n14129 = ~n13084 & ~n13086;
  assign n14130 = ~n54669 & ~n54670;
  assign n14131 = ~n14125 & n14130;
  assign n14132 = ~n14124 & ~n14125;
  assign n14133 = ~n14130 & n14132;
  assign n14134 = ~n14125 & ~n14133;
  assign n14135 = ~n14124 & ~n14131;
  assign n14136 = n13115 & ~n54671;
  assign n14137 = n14071 & n54662;
  assign n14138 = ~n14079 & ~n14137;
  assign n14139 = n123 & n11380;
  assign n14140 = n127 & ~n53685;
  assign n14141 = n128 & ~n53657;
  assign n14142 = n53444 & ~n53712;
  assign n14143 = ~n14141 & ~n14142;
  assign n14144 = ~n14140 & ~n14142;
  assign n14145 = ~n14141 & n14144;
  assign n14146 = ~n14140 & n14143;
  assign n14147 = ~n123 & n54672;
  assign n14148 = ~n11380 & n54672;
  assign n14149 = ~n14147 & ~n14148;
  assign n14150 = ~n14139 & n54672;
  assign n14151 = pi26  & ~n54673;
  assign n14152 = ~pi26  & n54673;
  assign n14153 = ~n14151 & ~n14152;
  assign n14154 = n14138 & ~n14153;
  assign n14155 = ~n13355 & n14069;
  assign n14156 = ~n14070 & ~n14155;
  assign n14157 = n11279 & n12690;
  assign n14158 = ~n53774 & n12584;
  assign n14159 = ~n53819 & n54410;
  assign n14160 = ~n53799 & n11267;
  assign n14161 = ~n14159 & ~n14160;
  assign n14162 = ~n14158 & ~n14159;
  assign n14163 = ~n14160 & n14162;
  assign n14164 = ~n14158 & n14161;
  assign n14165 = ~n11279 & n54674;
  assign n14166 = ~n12690 & n54674;
  assign n14167 = ~n14165 & ~n14166;
  assign n14168 = ~n14157 & n54674;
  assign n14169 = pi29  & ~n54675;
  assign n14170 = ~pi29  & n54675;
  assign n14171 = ~n14169 & ~n14170;
  assign n14172 = n14156 & ~n14171;
  assign n14173 = n123 & n11360;
  assign n14174 = n128 & ~n53685;
  assign n14175 = n53444 & ~n53741;
  assign n14176 = n127 & ~n53712;
  assign n14177 = ~n14175 & ~n14176;
  assign n14178 = ~n14174 & ~n14175;
  assign n14179 = ~n14176 & n14178;
  assign n14180 = ~n14174 & n14177;
  assign n14181 = ~n14173 & n54676;
  assign n14182 = pi26  & ~n14181;
  assign n14183 = pi26  & ~n14182;
  assign n14184 = pi26  & n14181;
  assign n14185 = ~n14181 & ~n14182;
  assign n14186 = ~pi26  & ~n14181;
  assign n14187 = ~n54677 & ~n54678;
  assign n14188 = ~n14156 & n14171;
  assign n14189 = ~n14187 & ~n14188;
  assign n14190 = ~n14172 & ~n14188;
  assign n14191 = ~n14187 & n14190;
  assign n14192 = ~n14172 & ~n14191;
  assign n14193 = ~n14172 & ~n14189;
  assign n14194 = ~n14138 & n14153;
  assign n14195 = n14138 & ~n14154;
  assign n14196 = n14138 & n14153;
  assign n14197 = ~n14153 & ~n14154;
  assign n14198 = ~n14138 & ~n14153;
  assign n14199 = ~n54680 & ~n54681;
  assign n14200 = ~n14154 & ~n14194;
  assign n14201 = ~n54679 & ~n54682;
  assign n14202 = ~n14154 & ~n14201;
  assign n14203 = n14096 & ~n14099;
  assign n14204 = ~n14098 & n14203;
  assign n14205 = n14096 & n54665;
  assign n14206 = ~n14102 & ~n54683;
  assign n14207 = ~n14202 & n14206;
  assign n14208 = n90 & n54351;
  assign n14209 = ~n53634 & n54667;
  assign n14210 = ~n53441 & n54666;
  assign n14211 = ~n2325 & n14210;
  assign n14212 = ~n14209 & ~n14211;
  assign n14213 = ~n14208 & n14212;
  assign n14214 = pi23  & ~n14213;
  assign n14215 = ~n14213 & ~n14214;
  assign n14216 = ~pi23  & ~n14213;
  assign n14217 = pi23  & ~n14214;
  assign n14218 = pi23  & n14213;
  assign n14219 = ~n54684 & ~n54685;
  assign n14220 = n14202 & ~n14206;
  assign n14221 = ~n14207 & ~n14220;
  assign n14222 = ~n14219 & n14221;
  assign n14223 = ~n14207 & ~n14222;
  assign n14224 = n14130 & ~n14132;
  assign n14225 = ~n14130 & ~n14133;
  assign n14226 = n14132 & ~n14133;
  assign n14227 = ~n14225 & ~n14226;
  assign n14228 = ~n14133 & ~n14224;
  assign n14229 = ~n14223 & ~n54686;
  assign n14230 = n14223 & n54686;
  assign n14231 = ~n14229 & ~n14230;
  assign n14232 = n14219 & ~n14221;
  assign n14233 = ~n14222 & ~n14232;
  assign n14234 = n90 & n11242;
  assign n14235 = ~n53650 & n54667;
  assign n14236 = n53441 & ~n53442;
  assign n14237 = ~n2325 & n14236;
  assign n14238 = ~n53634 & n14210;
  assign n14239 = ~n14237 & ~n14238;
  assign n14240 = ~n14235 & ~n14238;
  assign n14241 = ~n14237 & n14240;
  assign n14242 = ~n14235 & n14239;
  assign n14243 = ~n90 & n54687;
  assign n14244 = ~n11242 & n54687;
  assign n14245 = ~n14243 & ~n14244;
  assign n14246 = ~n14234 & n54687;
  assign n14247 = pi23  & ~n54688;
  assign n14248 = ~pi23  & n54688;
  assign n14249 = ~n14247 & ~n14248;
  assign n14250 = n14187 & ~n14190;
  assign n14251 = n14190 & ~n14191;
  assign n14252 = ~n14187 & ~n14191;
  assign n14253 = ~n14251 & ~n14252;
  assign n14254 = ~n14191 & ~n14250;
  assign n14255 = ~n14052 & n14067;
  assign n14256 = ~n14068 & ~n14255;
  assign n14257 = ~n13519 & ~n54655;
  assign n14258 = n54655 & ~n54656;
  assign n14259 = ~n13518 & n14040;
  assign n14260 = ~n14258 & ~n14259;
  assign n14261 = ~n54656 & ~n14257;
  assign n14262 = n10486 & ~n10488;
  assign n14263 = ~n10489 & ~n14262;
  assign n14264 = n1576 & n14263;
  assign n14265 = ~n53962 & n54403;
  assign n14266 = ~n53930 & n10564;
  assign n14267 = ~n53907 & n11215;
  assign n14268 = ~n14266 & ~n14267;
  assign n14269 = ~n14265 & ~n14266;
  assign n14270 = ~n14267 & n14269;
  assign n14271 = ~n14265 & n14268;
  assign n14272 = ~n14264 & ~n14265;
  assign n14273 = ~n14266 & n14272;
  assign n14274 = ~n14267 & n14273;
  assign n14275 = ~n14264 & n54691;
  assign n14276 = ~n54690 & ~n54692;
  assign n14277 = n11279 & n12918;
  assign n14278 = ~n53860 & n11267;
  assign n14279 = ~n53888 & n54410;
  assign n14280 = ~n53845 & n12584;
  assign n14281 = ~n14279 & ~n14280;
  assign n14282 = ~n14278 & ~n14279;
  assign n14283 = ~n14280 & n14282;
  assign n14284 = ~n14278 & n14281;
  assign n14285 = ~n14277 & n54693;
  assign n14286 = pi29  & ~n14285;
  assign n14287 = ~n14285 & ~n14286;
  assign n14288 = ~pi29  & ~n14285;
  assign n14289 = pi29  & ~n14286;
  assign n14290 = pi29  & n14285;
  assign n14291 = ~n54694 & ~n54695;
  assign n14292 = n54690 & n54692;
  assign n14293 = ~n54690 & ~n14276;
  assign n14294 = ~n54690 & n54692;
  assign n14295 = ~n54692 & ~n14276;
  assign n14296 = n54690 & ~n54692;
  assign n14297 = ~n54696 & ~n54697;
  assign n14298 = ~n14276 & ~n14292;
  assign n14299 = ~n14291 & ~n54698;
  assign n14300 = ~n14276 & ~n14299;
  assign n14301 = n14040 & ~n14042;
  assign n14302 = ~n14043 & ~n14301;
  assign n14303 = ~n14300 & n14302;
  assign n14304 = n14300 & ~n14302;
  assign n14305 = n11279 & n12938;
  assign n14306 = ~n53819 & n12584;
  assign n14307 = ~n53860 & n54410;
  assign n14308 = ~n53845 & n11267;
  assign n14309 = ~n14307 & ~n14308;
  assign n14310 = ~n14306 & ~n14307;
  assign n14311 = ~n14308 & n14310;
  assign n14312 = ~n14306 & n14309;
  assign n14313 = ~n14305 & n54699;
  assign n14314 = pi29  & ~n14313;
  assign n14315 = pi29  & ~n14314;
  assign n14316 = pi29  & n14313;
  assign n14317 = ~n14313 & ~n14314;
  assign n14318 = ~pi29  & ~n14313;
  assign n14319 = ~n54700 & ~n54701;
  assign n14320 = ~n14304 & ~n14319;
  assign n14321 = ~n14303 & ~n14304;
  assign n14322 = ~n14319 & n14321;
  assign n14323 = ~n14303 & ~n14322;
  assign n14324 = ~n14303 & ~n14320;
  assign n14325 = n14256 & ~n54702;
  assign n14326 = ~n14256 & n54702;
  assign n14327 = n123 & n11889;
  assign n14328 = n128 & ~n53712;
  assign n14329 = n53444 & ~n53774;
  assign n14330 = n127 & ~n53741;
  assign n14331 = ~n14329 & ~n14330;
  assign n14332 = ~n14328 & ~n14329;
  assign n14333 = ~n14330 & n14332;
  assign n14334 = ~n14328 & n14331;
  assign n14335 = ~n14327 & n54703;
  assign n14336 = pi26  & ~n14335;
  assign n14337 = pi26  & ~n14336;
  assign n14338 = pi26  & n14335;
  assign n14339 = ~n14335 & ~n14336;
  assign n14340 = ~pi26  & ~n14335;
  assign n14341 = ~n54704 & ~n54705;
  assign n14342 = ~n14326 & ~n14341;
  assign n14343 = ~n14325 & ~n14326;
  assign n14344 = ~n14341 & n14343;
  assign n14345 = ~n14325 & ~n14344;
  assign n14346 = ~n14325 & ~n14342;
  assign n14347 = ~n54689 & ~n54706;
  assign n14348 = n54689 & n54706;
  assign n14349 = n90 & n11286;
  assign n14350 = ~n53650 & n14210;
  assign n14351 = ~n53657 & n54667;
  assign n14352 = ~n53634 & n14236;
  assign n14353 = ~n14351 & ~n14352;
  assign n14354 = ~n14350 & ~n14351;
  assign n14355 = ~n14352 & n14354;
  assign n14356 = ~n14350 & n14353;
  assign n14357 = ~n14349 & n54707;
  assign n14358 = pi23  & ~n14357;
  assign n14359 = pi23  & ~n14358;
  assign n14360 = pi23  & n14357;
  assign n14361 = ~n14357 & ~n14358;
  assign n14362 = ~pi23  & ~n14357;
  assign n14363 = ~n54708 & ~n54709;
  assign n14364 = ~n14348 & ~n14363;
  assign n14365 = ~n14347 & ~n14348;
  assign n14366 = ~n14363 & n14365;
  assign n14367 = ~n14347 & ~n14366;
  assign n14368 = ~n14347 & ~n14364;
  assign n14369 = ~n14249 & ~n54710;
  assign n14370 = n14249 & n54710;
  assign n14371 = n54679 & n54682;
  assign n14372 = ~n54679 & ~n14201;
  assign n14373 = ~n54679 & n54682;
  assign n14374 = ~n54682 & ~n14201;
  assign n14375 = n54679 & ~n54682;
  assign n14376 = ~n54711 & ~n54712;
  assign n14377 = ~n14201 & ~n14371;
  assign n14378 = ~n14370 & ~n54713;
  assign n14379 = ~n14369 & ~n14370;
  assign n14380 = ~n54713 & n14379;
  assign n14381 = ~n14369 & ~n14380;
  assign n14382 = ~n14369 & ~n14378;
  assign n14383 = n14233 & ~n54714;
  assign n14384 = n54713 & ~n14379;
  assign n14385 = n14379 & ~n14380;
  assign n14386 = ~n54713 & ~n14380;
  assign n14387 = ~n14385 & ~n14386;
  assign n14388 = ~n14380 & ~n14384;
  assign n14389 = pi19  & ~pi20 ;
  assign n14390 = ~pi19  & pi20 ;
  assign n14391 = ~pi19  & ~pi20 ;
  assign n14392 = pi19  & pi20 ;
  assign n14393 = ~n14391 & ~n14392;
  assign n14394 = ~n14389 & ~n14390;
  assign n14395 = pi17  & ~pi18 ;
  assign n14396 = ~pi17  & pi18 ;
  assign n14397 = ~pi17  & ~pi18 ;
  assign n14398 = pi17  & pi18 ;
  assign n14399 = ~n14397 & ~n14398;
  assign n14400 = ~n14395 & ~n14396;
  assign n14401 = pi18  & ~pi19 ;
  assign n14402 = ~pi18  & pi19 ;
  assign n14403 = ~pi18  & ~pi19 ;
  assign n14404 = pi18  & pi19 ;
  assign n14405 = ~n14403 & ~n14404;
  assign n14406 = ~n14401 & ~n14402;
  assign n14407 = ~n54717 & ~n54718;
  assign n14408 = n54716 & ~n54717;
  assign n14409 = ~n54718 & n14408;
  assign n14410 = n54716 & ~n54718;
  assign n14411 = ~n54717 & n14410;
  assign n14412 = n54716 & n14407;
  assign n14413 = n54716 & n54717;
  assign n14414 = ~n10547 & n14413;
  assign n14415 = ~n54719 & ~n14414;
  assign n14416 = ~n2325 & n54719;
  assign n14417 = ~n10551 & ~n14416;
  assign n14418 = ~n14413 & ~n14416;
  assign n14419 = ~n14417 & ~n14418;
  assign n14420 = ~n2325 & ~n14415;
  assign n14421 = pi20  & ~n54720;
  assign n14422 = ~pi20  & n54720;
  assign n14423 = ~n14421 & ~n14422;
  assign n14424 = n123 & n11913;
  assign n14425 = n127 & ~n53774;
  assign n14426 = n53444 & ~n53799;
  assign n14427 = n128 & ~n53741;
  assign n14428 = ~n14426 & ~n14427;
  assign n14429 = ~n14425 & ~n14426;
  assign n14430 = ~n14427 & n14429;
  assign n14431 = ~n14425 & n14428;
  assign n14432 = ~n123 & n54721;
  assign n14433 = ~n11913 & n54721;
  assign n14434 = ~n14432 & ~n14433;
  assign n14435 = ~n14424 & n54721;
  assign n14436 = pi26  & ~n54722;
  assign n14437 = ~pi26  & n54722;
  assign n14438 = ~n14436 & ~n14437;
  assign n14439 = n14319 & ~n14321;
  assign n14440 = n14321 & ~n14322;
  assign n14441 = ~n14319 & ~n14322;
  assign n14442 = ~n14440 & ~n14441;
  assign n14443 = ~n14322 & ~n14439;
  assign n14444 = ~n14438 & ~n54723;
  assign n14445 = n14438 & n54723;
  assign n14446 = ~n14444 & ~n14445;
  assign n14447 = ~n274 & ~n420;
  assign n14448 = ~n410 & ~n748;
  assign n14449 = ~n1486 & n14448;
  assign n14450 = ~n748 & ~n1486;
  assign n14451 = ~n274 & n14450;
  assign n14452 = ~n420 & n14451;
  assign n14453 = ~n410 & n14452;
  assign n14454 = ~n420 & ~n1486;
  assign n14455 = ~n274 & ~n748;
  assign n14456 = ~n410 & n14455;
  assign n14457 = n14454 & n14456;
  assign n14458 = ~n410 & n14454;
  assign n14459 = n14455 & n14458;
  assign n14460 = n14447 & n14449;
  assign n14461 = n561 & n3672;
  assign n14462 = n3672 & n9739;
  assign n14463 = n561 & n14462;
  assign n14464 = n9739 & n14461;
  assign n14465 = ~n246 & ~n628;
  assign n14466 = ~n491 & ~n911;
  assign n14467 = ~n491 & ~n628;
  assign n14468 = ~n246 & ~n911;
  assign n14469 = n14467 & n14468;
  assign n14470 = ~n628 & ~n911;
  assign n14471 = ~n246 & ~n491;
  assign n14472 = n14470 & n14471;
  assign n14473 = n14465 & n14466;
  assign n14474 = n54340 & n54726;
  assign n14475 = n54725 & n14474;
  assign n14476 = n9739 & n54340;
  assign n14477 = n54724 & n14476;
  assign n14478 = n561 & n14477;
  assign n14479 = n3672 & n14478;
  assign n14480 = ~n628 & n14479;
  assign n14481 = ~n246 & n14480;
  assign n14482 = ~n911 & n14481;
  assign n14483 = ~n491 & n14482;
  assign n14484 = n54724 & n14475;
  assign n14485 = ~n269 & ~n833;
  assign n14486 = ~n740 & ~n833;
  assign n14487 = ~n269 & n14486;
  assign n14488 = ~n740 & n14485;
  assign n14489 = ~n630 & ~n649;
  assign n14490 = n3670 & n14489;
  assign n14491 = n54728 & n14490;
  assign n14492 = n53720 & n14491;
  assign n14493 = ~n754 & ~n1081;
  assign n14494 = ~n902 & ~n1491;
  assign n14495 = n14493 & n14494;
  assign n14496 = ~n320 & ~n503;
  assign n14497 = n12007 & n14496;
  assign n14498 = ~n902 & n12007;
  assign n14499 = ~n320 & n14498;
  assign n14500 = ~n1491 & n14499;
  assign n14501 = ~n1081 & n14500;
  assign n14502 = ~n503 & n14501;
  assign n14503 = ~n754 & n14502;
  assign n14504 = ~n902 & ~n1081;
  assign n14505 = n14496 & n14504;
  assign n14506 = n5070 & n12007;
  assign n14507 = n14505 & n14506;
  assign n14508 = ~n503 & ~n1491;
  assign n14509 = n14504 & n14508;
  assign n14510 = ~n320 & ~n754;
  assign n14511 = n12007 & n14510;
  assign n14512 = n14509 & n14511;
  assign n14513 = ~n320 & ~n902;
  assign n14514 = n14493 & n14513;
  assign n14515 = n12007 & n14508;
  assign n14516 = n14514 & n14515;
  assign n14517 = n14495 & n14497;
  assign n14518 = n4530 & n9511;
  assign n14519 = ~n295 & ~n568;
  assign n14520 = ~n247 & ~n1189;
  assign n14521 = n14519 & n14520;
  assign n14522 = n14518 & n14521;
  assign n14523 = n54152 & n14522;
  assign n14524 = n54729 & n14523;
  assign n14525 = n14489 & n14519;
  assign n14526 = n54728 & n14525;
  assign n14527 = n53720 & n14526;
  assign n14528 = n3670 & n4530;
  assign n14529 = n9511 & n14520;
  assign n14530 = n14528 & n14529;
  assign n14531 = n54152 & n14530;
  assign n14532 = n54729 & n14531;
  assign n14533 = n14527 & n14532;
  assign n14534 = n14492 & n14524;
  assign n14535 = n54727 & n54730;
  assign n14536 = n799 & n3134;
  assign n14537 = n2949 & n5378;
  assign n14538 = n14536 & n14537;
  assign n14539 = ~n353 & ~n751;
  assign n14540 = ~n353 & n3525;
  assign n14541 = ~n751 & n14540;
  assign n14542 = n3525 & n14539;
  assign n14543 = ~n363 & ~n591;
  assign n14544 = n424 & n14543;
  assign n14545 = n54731 & n14544;
  assign n14546 = n14538 & n14545;
  assign n14547 = n164 & ~n590;
  assign n14548 = n164 & n4223;
  assign n14549 = ~n590 & n14548;
  assign n14550 = ~n590 & n4223;
  assign n14551 = n164 & n14550;
  assign n14552 = n4223 & n14547;
  assign n14553 = n1957 & n11428;
  assign n14554 = ~n291 & ~n956;
  assign n14555 = n13164 & n14554;
  assign n14556 = n14553 & n14555;
  assign n14557 = n53801 & n14556;
  assign n14558 = n54732 & n14557;
  assign n14559 = n3134 & n54732;
  assign n14560 = n54731 & n14559;
  assign n14561 = n53801 & n14560;
  assign n14562 = n2949 & n14561;
  assign n14563 = n5378 & n14562;
  assign n14564 = n799 & n14563;
  assign n14565 = n11428 & n14564;
  assign n14566 = n1957 & n14565;
  assign n14567 = n424 & n14566;
  assign n14568 = n13164 & n14567;
  assign n14569 = ~n291 & n14568;
  assign n14570 = ~n956 & n14569;
  assign n14571 = ~n591 & n14570;
  assign n14572 = ~n363 & n14571;
  assign n14573 = n799 & n2949;
  assign n14574 = n1957 & n5378;
  assign n14575 = n14573 & n14574;
  assign n14576 = n3134 & n14543;
  assign n14577 = n54731 & n14576;
  assign n14578 = n14575 & n14577;
  assign n14579 = n424 & n11428;
  assign n14580 = n14555 & n14579;
  assign n14581 = n53801 & n14580;
  assign n14582 = n54732 & n14581;
  assign n14583 = n14578 & n14582;
  assign n14584 = n424 & n1957;
  assign n14585 = n799 & n5378;
  assign n14586 = n14584 & n14585;
  assign n14587 = ~n291 & ~n591;
  assign n14588 = ~n363 & ~n956;
  assign n14589 = n14587 & n14588;
  assign n14590 = n54731 & n14589;
  assign n14591 = n14586 & n14590;
  assign n14592 = n2949 & n3134;
  assign n14593 = n11428 & n13164;
  assign n14594 = n14592 & n14593;
  assign n14595 = n53801 & n14594;
  assign n14596 = n54732 & n14595;
  assign n14597 = n14591 & n14596;
  assign n14598 = n14546 & n14558;
  assign n14599 = ~n565 & n850;
  assign n14600 = n850 & n11134;
  assign n14601 = ~n565 & n14600;
  assign n14602 = ~n565 & n11134;
  assign n14603 = n850 & n14602;
  assign n14604 = n11134 & n14599;
  assign n14605 = ~n975 & ~n2103;
  assign n14606 = ~n554 & ~n1644;
  assign n14607 = n10901 & n14606;
  assign n14608 = n10901 & n14605;
  assign n14609 = n14606 & n14608;
  assign n14610 = n14605 & n14607;
  assign n14611 = ~n948 & ~n1492;
  assign n14612 = n2752 & n14611;
  assign n14613 = n4383 & n5390;
  assign n14614 = n14612 & n14613;
  assign n14615 = n54735 & n14614;
  assign n14616 = n54734 & n14615;
  assign n14617 = n53777 & n54393;
  assign n14618 = n12077 & n14617;
  assign n14619 = n53614 & n14618;
  assign n14620 = n54393 & n54734;
  assign n14621 = n4383 & n14620;
  assign n14622 = n4470 & n14621;
  assign n14623 = n53614 & n14622;
  assign n14624 = n10901 & n14623;
  assign n14625 = n5390 & n14624;
  assign n14626 = n53777 & n14625;
  assign n14627 = n1670 & n14626;
  assign n14628 = ~n948 & n14627;
  assign n14629 = ~n1471 & n14628;
  assign n14630 = ~n2103 & n14629;
  assign n14631 = ~n1490 & n14630;
  assign n14632 = ~n1492 & n14631;
  assign n14633 = ~n554 & n14632;
  assign n14634 = ~n975 & n14633;
  assign n14635 = ~n1644 & n14634;
  assign n14636 = n14605 & n14613;
  assign n14637 = n4470 & n10901;
  assign n14638 = n1670 & n2752;
  assign n14639 = n14637 & n14638;
  assign n14640 = n14636 & n14639;
  assign n14641 = n54734 & n14640;
  assign n14642 = ~n554 & ~n948;
  assign n14643 = ~n1492 & ~n1644;
  assign n14644 = n14642 & n14643;
  assign n14645 = n54393 & n14644;
  assign n14646 = n53777 & n14645;
  assign n14647 = n53614 & n14646;
  assign n14648 = n14641 & n14647;
  assign n14649 = n4470 & n5390;
  assign n14650 = n10901 & n14649;
  assign n14651 = ~n948 & ~n1471;
  assign n14652 = ~n1490 & ~n1644;
  assign n14653 = n14651 & n14652;
  assign n14654 = n1670 & n4383;
  assign n14655 = n14653 & n14654;
  assign n14656 = n14650 & n14655;
  assign n14657 = n54734 & n14656;
  assign n14658 = ~n975 & ~n1492;
  assign n14659 = ~n554 & ~n2103;
  assign n14660 = n14658 & n14659;
  assign n14661 = n53777 & n14660;
  assign n14662 = n54393 & n14661;
  assign n14663 = n53614 & n14662;
  assign n14664 = n14657 & n14663;
  assign n14665 = n14616 & n14619;
  assign n14666 = n54733 & n54736;
  assign n14667 = n54152 & n14520;
  assign n14668 = n54727 & n14667;
  assign n14669 = n54736 & n14668;
  assign n14670 = n53720 & n14669;
  assign n14671 = n54733 & n14670;
  assign n14672 = n54729 & n14671;
  assign n14673 = n3670 & n14672;
  assign n14674 = n4530 & n14673;
  assign n14675 = n9511 & n14674;
  assign n14676 = ~n295 & n14675;
  assign n14677 = ~n568 & n14676;
  assign n14678 = ~n833 & n14677;
  assign n14679 = ~n630 & n14678;
  assign n14680 = ~n269 & n14679;
  assign n14681 = ~n649 & n14680;
  assign n14682 = ~n740 & n14681;
  assign n14683 = n14535 & n14666;
  assign n14684 = n54636 & ~n54737;
  assign n14685 = ~n54636 & n54737;
  assign n14686 = ~n14684 & ~n14685;
  assign n14687 = n10474 & ~n10476;
  assign n14688 = ~n10477 & ~n14687;
  assign n14689 = n1576 & n14688;
  assign n14690 = ~n54005 & n10564;
  assign n14691 = ~n54034 & n54403;
  assign n14692 = ~n53970 & n11215;
  assign n14693 = ~n14691 & ~n14692;
  assign n14694 = ~n14690 & ~n14691;
  assign n14695 = ~n14692 & n14694;
  assign n14696 = ~n14690 & n14693;
  assign n14697 = ~n14689 & n54738;
  assign n14698 = ~n14684 & ~n14697;
  assign n14699 = ~n14685 & n14698;
  assign n14700 = n14686 & ~n14697;
  assign n14701 = ~n14684 & ~n54739;
  assign n14702 = ~pi14  & ~n54653;
  assign n14703 = ~n14011 & n14016;
  assign n14704 = ~n14702 & ~n14703;
  assign n14705 = ~n14701 & ~n14704;
  assign n14706 = n14701 & n14704;
  assign n14707 = n10478 & ~n10480;
  assign n14708 = ~n10481 & ~n14707;
  assign n14709 = n1576 & n14708;
  assign n14710 = ~n54005 & n54403;
  assign n14711 = ~n53970 & n10564;
  assign n14712 = ~n53962 & n11215;
  assign n14713 = ~n14711 & ~n14712;
  assign n14714 = ~n14710 & ~n14711;
  assign n14715 = ~n14712 & n14714;
  assign n14716 = ~n14710 & n14713;
  assign n14717 = ~n14709 & n54740;
  assign n14718 = ~n14706 & ~n14717;
  assign n14719 = ~n14705 & ~n14706;
  assign n14720 = ~n14717 & n14719;
  assign n14721 = ~n14705 & ~n14720;
  assign n14722 = ~n14705 & ~n14718;
  assign n14723 = n14029 & ~n14033;
  assign n14724 = ~n14029 & ~n14034;
  assign n14725 = n14033 & ~n14034;
  assign n14726 = ~n14724 & ~n14725;
  assign n14727 = ~n14034 & ~n14723;
  assign n14728 = ~n54741 & ~n54742;
  assign n14729 = n54741 & n54742;
  assign n14730 = ~n14728 & ~n14729;
  assign n14731 = n11279 & n13336;
  assign n14732 = ~n53888 & n11267;
  assign n14733 = ~n53907 & n54410;
  assign n14734 = ~n53860 & n12584;
  assign n14735 = ~n14733 & ~n14734;
  assign n14736 = ~n14732 & ~n14733;
  assign n14737 = ~n14734 & n14736;
  assign n14738 = ~n14732 & n14735;
  assign n14739 = ~n11279 & n54743;
  assign n14740 = ~n13336 & n54743;
  assign n14741 = ~n14739 & ~n14740;
  assign n14742 = ~n14731 & n54743;
  assign n14743 = pi29  & ~n54744;
  assign n14744 = ~pi29  & n54744;
  assign n14745 = ~n14743 & ~n14744;
  assign n14746 = n14730 & ~n14745;
  assign n14747 = ~n14728 & ~n14746;
  assign n14748 = n14291 & n54698;
  assign n14749 = ~n14291 & ~n14299;
  assign n14750 = ~n54698 & ~n14299;
  assign n14751 = ~n14749 & ~n14750;
  assign n14752 = ~n14299 & ~n14748;
  assign n14753 = ~n14747 & ~n54745;
  assign n14754 = n14747 & n54745;
  assign n14755 = n123 & n12690;
  assign n14756 = n128 & ~n53774;
  assign n14757 = n53444 & ~n53819;
  assign n14758 = n127 & ~n53799;
  assign n14759 = ~n14757 & ~n14758;
  assign n14760 = ~n14756 & ~n14757;
  assign n14761 = ~n14758 & n14760;
  assign n14762 = ~n14756 & n14759;
  assign n14763 = ~n14755 & n54746;
  assign n14764 = pi26  & ~n14763;
  assign n14765 = pi26  & ~n14764;
  assign n14766 = pi26  & n14763;
  assign n14767 = ~n14763 & ~n14764;
  assign n14768 = ~pi26  & ~n14763;
  assign n14769 = ~n54747 & ~n54748;
  assign n14770 = ~n14754 & ~n14769;
  assign n14771 = ~n14753 & ~n14754;
  assign n14772 = ~n14769 & n14771;
  assign n14773 = ~n14753 & ~n14772;
  assign n14774 = ~n14753 & ~n14770;
  assign n14775 = n14446 & ~n54749;
  assign n14776 = ~n14444 & ~n14775;
  assign n14777 = n14341 & ~n14343;
  assign n14778 = n14343 & ~n14344;
  assign n14779 = ~n14341 & ~n14344;
  assign n14780 = ~n14778 & ~n14779;
  assign n14781 = ~n14344 & ~n14777;
  assign n14782 = ~n14776 & ~n54750;
  assign n14783 = n14776 & n54750;
  assign n14784 = n90 & n11213;
  assign n14785 = ~n53650 & n14236;
  assign n14786 = ~n53685 & n54667;
  assign n14787 = ~n53657 & n14210;
  assign n14788 = ~n14786 & ~n14787;
  assign n14789 = ~n14785 & n14788;
  assign n14790 = ~n14784 & n14789;
  assign n14791 = pi23  & ~n14790;
  assign n14792 = pi23  & ~n14791;
  assign n14793 = pi23  & n14790;
  assign n14794 = ~n14790 & ~n14791;
  assign n14795 = ~pi23  & ~n14790;
  assign n14796 = ~n54751 & ~n54752;
  assign n14797 = ~n14783 & ~n14796;
  assign n14798 = ~n14782 & ~n14783;
  assign n14799 = ~n14796 & n14798;
  assign n14800 = ~n14782 & ~n14799;
  assign n14801 = ~n14782 & ~n14797;
  assign n14802 = ~n14423 & ~n54753;
  assign n14803 = n14423 & n54753;
  assign n14804 = n14363 & ~n14365;
  assign n14805 = n14365 & ~n14366;
  assign n14806 = ~n14363 & ~n14366;
  assign n14807 = ~n14805 & ~n14806;
  assign n14808 = ~n14366 & ~n14804;
  assign n14809 = ~n14803 & ~n54754;
  assign n14810 = ~n14802 & ~n14803;
  assign n14811 = ~n54754 & n14810;
  assign n14812 = ~n14802 & ~n14811;
  assign n14813 = ~n14802 & ~n14809;
  assign n14814 = ~n54715 & ~n54755;
  assign n14815 = n54715 & n54755;
  assign n14816 = ~n14814 & ~n14815;
  assign n14817 = n54754 & ~n14810;
  assign n14818 = ~n54754 & ~n14811;
  assign n14819 = n14810 & ~n14811;
  assign n14820 = ~n14818 & ~n14819;
  assign n14821 = ~n14811 & ~n14817;
  assign n14822 = n90 & n11380;
  assign n14823 = ~n53685 & n14210;
  assign n14824 = ~n53657 & n14236;
  assign n14825 = ~n53712 & n54667;
  assign n14826 = ~n14824 & ~n14825;
  assign n14827 = ~n14823 & ~n14825;
  assign n14828 = ~n14824 & n14827;
  assign n14829 = ~n14823 & n14826;
  assign n14830 = ~n14822 & n54757;
  assign n14831 = pi23  & ~n14830;
  assign n14832 = ~n14830 & ~n14831;
  assign n14833 = ~pi23  & ~n14830;
  assign n14834 = pi23  & ~n14831;
  assign n14835 = pi23  & n14830;
  assign n14836 = ~n54758 & ~n54759;
  assign n14837 = ~n14446 & n54749;
  assign n14838 = ~n14775 & ~n14837;
  assign n14839 = ~n14836 & n14838;
  assign n14840 = n14836 & ~n14838;
  assign n14841 = ~n14836 & ~n14839;
  assign n14842 = ~n14836 & ~n14838;
  assign n14843 = n14838 & ~n14839;
  assign n14844 = n14836 & n14838;
  assign n14845 = ~n54760 & ~n54761;
  assign n14846 = ~n14839 & ~n14840;
  assign n14847 = n14769 & ~n14771;
  assign n14848 = n14771 & ~n14772;
  assign n14849 = ~n14769 & ~n14772;
  assign n14850 = ~n14848 & ~n14849;
  assign n14851 = ~n14772 & ~n14847;
  assign n14852 = n11279 & n13360;
  assign n14853 = ~n53907 & n11267;
  assign n14854 = ~n53930 & n54410;
  assign n14855 = ~n53888 & n12584;
  assign n14856 = ~n14854 & ~n14855;
  assign n14857 = ~n14853 & ~n14854;
  assign n14858 = ~n14855 & n14857;
  assign n14859 = ~n14853 & n14856;
  assign n14860 = ~n14852 & n54764;
  assign n14861 = pi29  & ~n14860;
  assign n14862 = ~n14860 & ~n14861;
  assign n14863 = ~pi29  & ~n14860;
  assign n14864 = pi29  & ~n14861;
  assign n14865 = pi29  & n14860;
  assign n14866 = ~n54765 & ~n54766;
  assign n14867 = n14717 & ~n14719;
  assign n14868 = ~n14717 & ~n14720;
  assign n14869 = n14719 & ~n14720;
  assign n14870 = ~n14868 & ~n14869;
  assign n14871 = ~n14720 & ~n14867;
  assign n14872 = ~n14866 & ~n54767;
  assign n14873 = ~n14686 & n14697;
  assign n14874 = ~n14697 & ~n54739;
  assign n14875 = ~n14685 & n14701;
  assign n14876 = ~n14874 & ~n14875;
  assign n14877 = ~n54739 & ~n14873;
  assign n14878 = ~n881 & n2326;
  assign n14879 = n2326 & n9337;
  assign n14880 = ~n881 & n14879;
  assign n14881 = ~n881 & n9337;
  assign n14882 = n2326 & n14881;
  assign n14883 = n9337 & n14878;
  assign n14884 = ~n419 & ~n1912;
  assign n14885 = n5058 & n14884;
  assign n14886 = n915 & n12436;
  assign n14887 = ~n174 & ~n1912;
  assign n14888 = ~n296 & ~n419;
  assign n14889 = n12436 & n14884;
  assign n14890 = n14887 & n14888;
  assign n14891 = n915 & n5058;
  assign n14892 = n54770 & n14891;
  assign n14893 = n14885 & n14886;
  assign n14894 = ~n182 & ~n451;
  assign n14895 = ~n451 & ~n747;
  assign n14896 = ~n182 & n14895;
  assign n14897 = ~n182 & ~n747;
  assign n14898 = ~n451 & n14897;
  assign n14899 = ~n747 & n14894;
  assign n14900 = ~n105 & ~n269;
  assign n14901 = ~n105 & ~n896;
  assign n14902 = ~n269 & n14901;
  assign n14903 = ~n896 & n14900;
  assign n14904 = n54772 & n54773;
  assign n14905 = n54771 & n14904;
  assign n14906 = n54769 & n14905;
  assign n14907 = n54061 & n54632;
  assign n14908 = n14906 & n14907;
  assign n14909 = ~n246 & ~n320;
  assign n14910 = ~n1485 & ~n1769;
  assign n14911 = ~n246 & ~n1769;
  assign n14912 = ~n320 & ~n1485;
  assign n14913 = n14911 & n14912;
  assign n14914 = n14909 & n14910;
  assign n14915 = n6288 & n54774;
  assign n14916 = ~n342 & ~n584;
  assign n14917 = ~n460 & ~n584;
  assign n14918 = ~n342 & n14917;
  assign n14919 = ~n460 & n14916;
  assign n14920 = n54116 & n54775;
  assign n14921 = n14915 & n14920;
  assign n14922 = ~n307 & ~n440;
  assign n14923 = n7307 & n14922;
  assign n14924 = ~n735 & ~n774;
  assign n14925 = n8185 & n14924;
  assign n14926 = ~n1085 & n7307;
  assign n14927 = ~n307 & n14926;
  assign n14928 = ~n1641 & n14927;
  assign n14929 = ~n440 & n14928;
  assign n14930 = ~n774 & n14929;
  assign n14931 = ~n735 & n14930;
  assign n14932 = n14922 & n14924;
  assign n14933 = n7307 & n8185;
  assign n14934 = n14932 & n14933;
  assign n14935 = n14923 & n14925;
  assign n14936 = n3255 & n5060;
  assign n14937 = ~n218 & ~n552;
  assign n14938 = n11829 & n14937;
  assign n14939 = n14936 & n14938;
  assign n14940 = n54776 & n14939;
  assign n14941 = n6288 & n54116;
  assign n14942 = n54775 & n14941;
  assign n14943 = n5060 & n14942;
  assign n14944 = n54776 & n14943;
  assign n14945 = n11829 & n14944;
  assign n14946 = ~n320 & n14945;
  assign n14947 = ~n1680 & n14946;
  assign n14948 = ~n1485 & n14947;
  assign n14949 = ~n218 & n14948;
  assign n14950 = ~n246 & n14949;
  assign n14951 = ~n552 & n14950;
  assign n14952 = ~n849 & n14951;
  assign n14953 = ~n1769 & n14952;
  assign n14954 = ~n320 & ~n849;
  assign n14955 = n14911 & n14954;
  assign n14956 = n6288 & n14955;
  assign n14957 = n14920 & n14956;
  assign n14958 = ~n1485 & ~n1680;
  assign n14959 = n14937 & n14958;
  assign n14960 = n5060 & n11829;
  assign n14961 = n14959 & n14960;
  assign n14962 = n54776 & n14961;
  assign n14963 = n14957 & n14962;
  assign n14964 = n14921 & n14940;
  assign n14965 = ~n184 & ~n503;
  assign n14966 = n3083 & n6482;
  assign n14967 = n14965 & n14966;
  assign n14968 = ~n222 & ~n401;
  assign n14969 = ~n401 & ~n773;
  assign n14970 = ~n222 & n14969;
  assign n14971 = ~n773 & n14968;
  assign n14972 = n318 & n1583;
  assign n14973 = n54778 & n14972;
  assign n14974 = n1278 & n13912;
  assign n14975 = n54270 & n14974;
  assign n14976 = n14973 & n14975;
  assign n14977 = n54270 & n14965;
  assign n14978 = n13912 & n14977;
  assign n14979 = n3083 & n14978;
  assign n14980 = n1278 & n14979;
  assign n14981 = n318 & n14980;
  assign n14982 = n6482 & n14981;
  assign n14983 = ~n222 & n14982;
  assign n14984 = ~n401 & n14983;
  assign n14985 = ~n591 & n14984;
  assign n14986 = ~n611 & n14985;
  assign n14987 = ~n773 & n14986;
  assign n14988 = n14965 & n14972;
  assign n14989 = n14966 & n54778;
  assign n14990 = n14975 & n14989;
  assign n14991 = n14988 & n14990;
  assign n14992 = n14965 & n14974;
  assign n14993 = ~n611 & ~n773;
  assign n14994 = n6482 & n14993;
  assign n14995 = n318 & n3083;
  assign n14996 = n14994 & n14995;
  assign n14997 = ~n401 & ~n591;
  assign n14998 = ~n222 & n14997;
  assign n14999 = n54270 & n14998;
  assign n15000 = n14996 & n14999;
  assign n15001 = n14992 & n15000;
  assign n15002 = n14967 & n14976;
  assign n15003 = n54777 & n54779;
  assign n15004 = n14908 & n15003;
  assign n15005 = n5058 & n54769;
  assign n15006 = n54773 & n15005;
  assign n15007 = n54772 & n15006;
  assign n15008 = n915 & n15007;
  assign n15009 = n54632 & n15008;
  assign n15010 = n54061 & n15009;
  assign n15011 = n53787 & n15010;
  assign n15012 = n54777 & n15011;
  assign n15013 = n54779 & n15012;
  assign n15014 = ~n296 & n15013;
  assign n15015 = ~n174 & n15014;
  assign n15016 = ~n419 & n15015;
  assign n15017 = ~n1912 & n15016;
  assign n15018 = n53787 & n15004;
  assign n15019 = n1704 & n5277;
  assign n15020 = n9766 & n12007;
  assign n15021 = n5277 & n9766;
  assign n15022 = n1704 & n12007;
  assign n15023 = n15021 & n15022;
  assign n15024 = n15019 & n15020;
  assign n15025 = ~n269 & ~n1912;
  assign n15026 = ~n1044 & ~n1468;
  assign n15027 = ~n269 & n15026;
  assign n15028 = ~n1912 & n15027;
  assign n15029 = ~n1468 & ~n1912;
  assign n15030 = ~n269 & ~n1044;
  assign n15031 = n15029 & n15030;
  assign n15032 = n15025 & n15026;
  assign n15033 = ~n249 & ~n554;
  assign n15034 = ~n504 & ~n554;
  assign n15035 = ~n249 & n15034;
  assign n15036 = ~n249 & ~n504;
  assign n15037 = ~n554 & n15036;
  assign n15038 = ~n504 & n15033;
  assign n15039 = n54782 & n54783;
  assign n15040 = n15020 & n54782;
  assign n15041 = n1704 & n15040;
  assign n15042 = n5277 & n15041;
  assign n15043 = ~n249 & n15042;
  assign n15044 = ~n554 & n15043;
  assign n15045 = ~n504 & n15044;
  assign n15046 = n54781 & n15039;
  assign n15047 = n1542 & n7201;
  assign n15048 = n7276 & n7526;
  assign n15049 = n15047 & n15048;
  assign n15050 = ~n218 & ~n1478;
  assign n15051 = ~n894 & ~n1478;
  assign n15052 = ~n218 & n15051;
  assign n15053 = ~n218 & ~n894;
  assign n15054 = ~n1478 & n15053;
  assign n15055 = ~n894 & n15050;
  assign n15056 = n2340 & n5639;
  assign n15057 = n54785 & n15056;
  assign n15058 = n15049 & n15057;
  assign n15059 = n1456 & n13958;
  assign n15060 = ~n507 & ~n735;
  assign n15061 = ~n291 & ~n902;
  assign n15062 = n15060 & n15061;
  assign n15063 = n15059 & n15062;
  assign n15064 = n53848 & n15063;
  assign n15065 = n1542 & n5639;
  assign n15066 = n7201 & n7276;
  assign n15067 = n15065 & n15066;
  assign n15068 = n2340 & n13958;
  assign n15069 = n54785 & n15068;
  assign n15070 = n15067 & n15069;
  assign n15071 = n1456 & n7526;
  assign n15072 = n15062 & n15071;
  assign n15073 = n53848 & n15072;
  assign n15074 = n15070 & n15073;
  assign n15075 = n2340 & n15060;
  assign n15076 = n15065 & n15075;
  assign n15077 = n7526 & n13958;
  assign n15078 = n54785 & n15077;
  assign n15079 = n15076 & n15078;
  assign n15080 = n1456 & n15061;
  assign n15081 = n15066 & n15080;
  assign n15082 = n53848 & n15081;
  assign n15083 = n15079 & n15082;
  assign n15084 = ~n291 & ~n510;
  assign n15085 = ~n507 & ~n1465;
  assign n15086 = n15084 & n15085;
  assign n15087 = n1542 & n2340;
  assign n15088 = n15086 & n15087;
  assign n15089 = ~n902 & ~n1127;
  assign n15090 = ~n735 & ~n1487;
  assign n15091 = n15089 & n15090;
  assign n15092 = n54785 & n15091;
  assign n15093 = n15088 & n15092;
  assign n15094 = n5639 & n7276;
  assign n15095 = n1456 & n7201;
  assign n15096 = n15094 & n15095;
  assign n15097 = n53848 & n15096;
  assign n15098 = n15093 & n15097;
  assign n15099 = n15058 & n15064;
  assign n15100 = n1456 & n54785;
  assign n15101 = n1542 & n15100;
  assign n15102 = n54784 & n15101;
  assign n15103 = n53848 & n15102;
  assign n15104 = n7201 & n15103;
  assign n15105 = n7276 & n15104;
  assign n15106 = n2340 & n15105;
  assign n15107 = n5639 & n15106;
  assign n15108 = ~n902 & n15107;
  assign n15109 = ~n291 & n15108;
  assign n15110 = ~n1127 & n15109;
  assign n15111 = ~n1465 & n15110;
  assign n15112 = ~n1487 & n15111;
  assign n15113 = ~n510 & n15112;
  assign n15114 = ~n507 & n15113;
  assign n15115 = ~n735 & n15114;
  assign n15116 = n54784 & n54786;
  assign n15117 = ~n168 & ~n848;
  assign n15118 = ~n956 & n15117;
  assign n15119 = ~n614 & ~n627;
  assign n15120 = n494 & n15119;
  assign n15121 = n15118 & n15120;
  assign n15122 = n53519 & n53932;
  assign n15123 = n15121 & n15122;
  assign n15124 = n5060 & n5199;
  assign n15125 = n5538 & n13551;
  assign n15126 = n15124 & n15125;
  assign n15127 = n2636 & n3014;
  assign n15128 = n3742 & n4070;
  assign n15129 = n15127 & n15128;
  assign n15130 = n15126 & n15129;
  assign n15131 = ~n848 & n15119;
  assign n15132 = ~n168 & ~n956;
  assign n15133 = n3014 & n15132;
  assign n15134 = n15131 & n15133;
  assign n15135 = n15122 & n15134;
  assign n15136 = n5199 & n5538;
  assign n15137 = n494 & n13551;
  assign n15138 = n15136 & n15137;
  assign n15139 = n4070 & n5060;
  assign n15140 = n2636 & n3742;
  assign n15141 = n15139 & n15140;
  assign n15142 = n15138 & n15141;
  assign n15143 = n15135 & n15142;
  assign n15144 = ~n956 & ~n1079;
  assign n15145 = ~n496 & n15144;
  assign n15146 = ~n627 & ~n2201;
  assign n15147 = ~n168 & ~n211;
  assign n15148 = n15146 & n15147;
  assign n15149 = n15145 & n15148;
  assign n15150 = n15122 & n15149;
  assign n15151 = n494 & n5538;
  assign n15152 = n15139 & n15151;
  assign n15153 = ~n614 & ~n848;
  assign n15154 = n5199 & n15153;
  assign n15155 = n3014 & n3742;
  assign n15156 = n15154 & n15155;
  assign n15157 = n15152 & n15156;
  assign n15158 = n15150 & n15157;
  assign n15159 = n15123 & n15130;
  assign n15160 = n54486 & n54788;
  assign n15161 = n54430 & n54779;
  assign n15162 = n15160 & n15161;
  assign n15163 = n5538 & n53932;
  assign n15164 = n54430 & n15163;
  assign n15165 = n5199 & n15164;
  assign n15166 = n5060 & n15165;
  assign n15167 = n54486 & n15166;
  assign n15168 = n53519 & n15167;
  assign n15169 = n494 & n15168;
  assign n15170 = n54787 & n15169;
  assign n15171 = n54779 & n15170;
  assign n15172 = n4070 & n15171;
  assign n15173 = n3014 & n15172;
  assign n15174 = n3742 & n15173;
  assign n15175 = ~n1079 & n15174;
  assign n15176 = ~n168 & n15175;
  assign n15177 = ~n211 & n15176;
  assign n15178 = ~n956 & n15177;
  assign n15179 = ~n848 & n15178;
  assign n15180 = ~n496 & n15179;
  assign n15181 = ~n627 & n15180;
  assign n15182 = ~n614 & n15181;
  assign n15183 = ~n2201 & n15182;
  assign n15184 = n54787 & n15162;
  assign n15185 = ~n54780 & ~n54789;
  assign n15186 = n54780 & n54789;
  assign n15187 = ~pi11  & ~n15185;
  assign n15188 = ~n15185 & ~n15186;
  assign n15189 = ~pi11  & n15188;
  assign n15190 = ~n15186 & n15187;
  assign n15191 = ~n15185 & ~n54790;
  assign n15192 = n54636 & ~n15191;
  assign n15193 = ~n54636 & n15191;
  assign n15194 = n10470 & ~n10472;
  assign n15195 = ~n10473 & ~n15194;
  assign n15196 = n1576 & n15195;
  assign n15197 = ~n54050 & n54403;
  assign n15198 = ~n54005 & n11215;
  assign n15199 = ~n54034 & n10564;
  assign n15200 = ~n15198 & ~n15199;
  assign n15201 = ~n15197 & ~n15199;
  assign n15202 = ~n15198 & n15201;
  assign n15203 = ~n15197 & n15200;
  assign n15204 = ~n15196 & n54791;
  assign n15205 = ~n15193 & ~n15204;
  assign n15206 = ~n15192 & n15204;
  assign n15207 = ~n15193 & ~n15206;
  assign n15208 = ~n15192 & ~n15193;
  assign n15209 = ~n15204 & n15208;
  assign n15210 = ~n15192 & ~n15209;
  assign n15211 = ~n15192 & ~n15205;
  assign n15212 = ~n54768 & n54792;
  assign n15213 = n54768 & ~n54792;
  assign n15214 = ~n15212 & ~n15213;
  assign n15215 = ~pi11  & ~n54790;
  assign n15216 = ~n15186 & n15191;
  assign n15217 = ~n15215 & ~n15216;
  assign n15218 = n10466 & ~n10468;
  assign n15219 = ~n10469 & ~n15218;
  assign n15220 = n1576 & n15219;
  assign n15221 = ~n54050 & n10564;
  assign n15222 = ~n54034 & n11215;
  assign n15223 = ~n54073 & n54403;
  assign n15224 = ~n15222 & ~n15223;
  assign n15225 = ~n15221 & n15224;
  assign n15226 = ~n15220 & ~n15223;
  assign n15227 = ~n15221 & n15226;
  assign n15228 = ~n15222 & n15227;
  assign n15229 = ~n15220 & n15225;
  assign n15230 = ~n15217 & ~n54793;
  assign n15231 = ~n774 & ~n851;
  assign n15232 = ~n881 & n15231;
  assign n15233 = n53895 & n15232;
  assign n15234 = ~n625 & ~n1881;
  assign n15235 = ~n625 & n6806;
  assign n15236 = ~n1881 & n15235;
  assign n15237 = n6806 & n15234;
  assign n15238 = ~n363 & ~n1472;
  assign n15239 = ~n1472 & n3214;
  assign n15240 = ~n363 & n15239;
  assign n15241 = n3214 & n15238;
  assign n15242 = n54794 & n54795;
  assign n15243 = n15233 & n15242;
  assign n15244 = ~n166 & ~n353;
  assign n15245 = ~n822 & ~n1477;
  assign n15246 = n1067 & n15245;
  assign n15247 = n1067 & ~n1477;
  assign n15248 = ~n166 & n15247;
  assign n15249 = ~n822 & n15248;
  assign n15250 = ~n353 & n15249;
  assign n15251 = n15244 & n15245;
  assign n15252 = n1067 & n15251;
  assign n15253 = n15244 & n15246;
  assign n15254 = ~n101 & ~n584;
  assign n15255 = n8052 & n15254;
  assign n15256 = n9256 & n9477;
  assign n15257 = n8052 & n9477;
  assign n15258 = n9256 & n15254;
  assign n15259 = n15257 & n15258;
  assign n15260 = n15255 & n15256;
  assign n15261 = n54796 & n54797;
  assign n15262 = ~n274 & ~n881;
  assign n15263 = ~n584 & n15262;
  assign n15264 = n53895 & n15263;
  assign n15265 = n15242 & n15264;
  assign n15266 = ~n101 & ~n246;
  assign n15267 = n15231 & n15266;
  assign n15268 = n15257 & n15267;
  assign n15269 = n54796 & n15268;
  assign n15270 = n15265 & n15269;
  assign n15271 = ~n246 & ~n881;
  assign n15272 = ~n774 & n15271;
  assign n15273 = n53895 & n15272;
  assign n15274 = n15242 & n15273;
  assign n15275 = ~n101 & ~n851;
  assign n15276 = ~n274 & ~n584;
  assign n15277 = n15275 & n15276;
  assign n15278 = n15257 & n15277;
  assign n15279 = n54796 & n15278;
  assign n15280 = n15274 & n15279;
  assign n15281 = n15243 & n15261;
  assign n15282 = n54434 & n54798;
  assign n15283 = n54053 & n15282;
  assign n15284 = n54067 & n15283;
  assign n15285 = n53895 & n15242;
  assign n15286 = n54796 & n15285;
  assign n15287 = n54067 & n15286;
  assign n15288 = n54434 & n15287;
  assign n15289 = n54053 & n15288;
  assign n15290 = n8052 & n15289;
  assign n15291 = n9477 & n15290;
  assign n15292 = n53872 & n15291;
  assign n15293 = ~n881 & n15292;
  assign n15294 = ~n101 & n15293;
  assign n15295 = ~n246 & n15294;
  assign n15296 = ~n584 & n15295;
  assign n15297 = ~n851 & n15296;
  assign n15298 = ~n274 & n15297;
  assign n15299 = ~n774 & n15298;
  assign n15300 = n53872 & n15284;
  assign n15301 = n54780 & ~n54799;
  assign n15302 = ~n54780 & n54799;
  assign n15303 = ~n15301 & ~n15302;
  assign n15304 = ~n291 & ~n631;
  assign n15305 = ~n956 & n15304;
  assign n15306 = ~n631 & n14554;
  assign n15307 = ~n567 & ~n628;
  assign n15308 = n9210 & n15307;
  assign n15309 = n9210 & n54800;
  assign n15310 = ~n628 & n15309;
  assign n15311 = ~n567 & n15310;
  assign n15312 = n54800 & n15308;
  assign n15313 = ~n824 & ~n1490;
  assign n15314 = ~n174 & ~n1997;
  assign n15315 = n6323 & n15314;
  assign n15316 = n15313 & n15315;
  assign n15317 = n54117 & n15316;
  assign n15318 = n54801 & n15317;
  assign n15319 = ~n216 & ~n735;
  assign n15320 = ~n901 & n15319;
  assign n15321 = n185 & n882;
  assign n15322 = n11427 & n15321;
  assign n15323 = ~n1192 & n15321;
  assign n15324 = ~n901 & n15323;
  assign n15325 = ~n321 & n15324;
  assign n15326 = ~n216 & n15325;
  assign n15327 = ~n735 & n15326;
  assign n15328 = ~n216 & n11427;
  assign n15329 = ~n735 & ~n901;
  assign n15330 = n882 & n15329;
  assign n15331 = n185 & n15330;
  assign n15332 = n15328 & n15331;
  assign n15333 = n15320 & n15322;
  assign n15334 = ~n754 & n4457;
  assign n15335 = n53573 & n15334;
  assign n15336 = n54785 & n15335;
  assign n15337 = n53470 & n15336;
  assign n15338 = n54802 & n15337;
  assign n15339 = ~n105 & ~n754;
  assign n15340 = n15314 & n15339;
  assign n15341 = n15313 & n15340;
  assign n15342 = n54117 & n15341;
  assign n15343 = n54801 & n15342;
  assign n15344 = ~n419 & ~n614;
  assign n15345 = ~n2201 & n15344;
  assign n15346 = n53573 & n15345;
  assign n15347 = n54785 & n15346;
  assign n15348 = n53470 & n15347;
  assign n15349 = n54802 & n15348;
  assign n15350 = n15343 & n15349;
  assign n15351 = ~n824 & ~n2201;
  assign n15352 = n6323 & n15351;
  assign n15353 = n15314 & n15352;
  assign n15354 = n54117 & n15353;
  assign n15355 = n54801 & n15354;
  assign n15356 = ~n419 & ~n1490;
  assign n15357 = ~n754 & n15356;
  assign n15358 = n53573 & n15357;
  assign n15359 = n54785 & n15358;
  assign n15360 = n53470 & n15359;
  assign n15361 = n54802 & n15360;
  assign n15362 = n15355 & n15361;
  assign n15363 = n15318 & n15338;
  assign n15364 = ~n562 & ~n1081;
  assign n15365 = ~n1081 & n5873;
  assign n15366 = ~n562 & n15365;
  assign n15367 = n5873 & n15364;
  assign n15368 = n54206 & n12078;
  assign n15369 = n54804 & n15368;
  assign n15370 = n9257 & n9479;
  assign n15371 = n11829 & n15370;
  assign n15372 = ~n259 & ~n404;
  assign n15373 = ~n493 & ~n770;
  assign n15374 = n15372 & n15373;
  assign n15375 = n2340 & n7525;
  assign n15376 = n15374 & n15375;
  assign n15377 = n9479 & n10361;
  assign n15378 = n11829 & n15377;
  assign n15379 = ~n108 & ~n493;
  assign n15380 = ~n259 & ~n647;
  assign n15381 = ~n493 & ~n647;
  assign n15382 = ~n108 & ~n259;
  assign n15383 = n15381 & n15382;
  assign n15384 = n15379 & n15380;
  assign n15385 = n2340 & n4833;
  assign n15386 = n54805 & n15385;
  assign n15387 = n15378 & n15386;
  assign n15388 = n15371 & n15376;
  assign n15389 = n54206 & n54805;
  assign n15390 = n54804 & n15389;
  assign n15391 = n2038 & n4833;
  assign n15392 = n2340 & n4585;
  assign n15393 = n15391 & n15392;
  assign n15394 = n15378 & n15393;
  assign n15395 = n15390 & n15394;
  assign n15396 = n9479 & n15379;
  assign n15397 = n54206 & n15396;
  assign n15398 = n54804 & n15397;
  assign n15399 = n11829 & n15391;
  assign n15400 = n10361 & n15380;
  assign n15401 = n15392 & n15400;
  assign n15402 = n15399 & n15401;
  assign n15403 = n15398 & n15402;
  assign n15404 = n15369 & n54806;
  assign n15405 = n54206 & n54804;
  assign n15406 = n2038 & n15405;
  assign n15407 = n54648 & n15406;
  assign n15408 = n4585 & n15407;
  assign n15409 = n4833 & n15408;
  assign n15410 = n2340 & n15409;
  assign n15411 = n11829 & n15410;
  assign n15412 = ~n108 & n15411;
  assign n15413 = ~n259 & n15412;
  assign n15414 = ~n221 & n15413;
  assign n15415 = ~n404 & n15414;
  assign n15416 = ~n493 & n15415;
  assign n15417 = ~n420 & n15416;
  assign n15418 = ~n647 & n15417;
  assign n15419 = ~n354 & n15418;
  assign n15420 = n54648 & n54807;
  assign n15421 = ~n789 & ~n1234;
  assign n15422 = ~n1065 & n15421;
  assign n15423 = ~n311 & ~n340;
  assign n15424 = ~n423 & ~n514;
  assign n15425 = ~n340 & ~n514;
  assign n15426 = ~n311 & ~n423;
  assign n15427 = n15425 & n15426;
  assign n15428 = n15423 & n15424;
  assign n15429 = ~n789 & n15424;
  assign n15430 = ~n340 & ~n1234;
  assign n15431 = ~n311 & ~n1065;
  assign n15432 = n15430 & n15431;
  assign n15433 = n15429 & n15432;
  assign n15434 = n15422 & n54809;
  assign n15435 = n53944 & n54627;
  assign n15436 = n54810 & n15435;
  assign n15437 = n208 & n2853;
  assign n15438 = n2256 & n15437;
  assign n15439 = n53919 & n15438;
  assign n15440 = ~n514 & ~n651;
  assign n15441 = ~n311 & n15440;
  assign n15442 = ~n1065 & ~n1234;
  assign n15443 = ~n789 & ~n1703;
  assign n15444 = n15442 & n15443;
  assign n15445 = n15441 & n15444;
  assign n15446 = n15435 & n15445;
  assign n15447 = ~n340 & ~n423;
  assign n15448 = n2256 & n15447;
  assign n15449 = n208 & n15448;
  assign n15450 = n53919 & n15449;
  assign n15451 = n15446 & n15450;
  assign n15452 = n15436 & n15439;
  assign n15453 = ~n1031 & ~n1034;
  assign n15454 = ~n1044 & ~n1492;
  assign n15455 = n15453 & n15454;
  assign n15456 = ~n268 & ~n585;
  assign n15457 = ~n416 & ~n833;
  assign n15458 = ~n585 & ~n833;
  assign n15459 = ~n268 & ~n416;
  assign n15460 = n15458 & n15459;
  assign n15461 = n15456 & n15457;
  assign n15462 = ~n268 & ~n1492;
  assign n15463 = ~n585 & ~n1044;
  assign n15464 = n15462 & n15463;
  assign n15465 = ~n833 & ~n1034;
  assign n15466 = ~n416 & ~n1031;
  assign n15467 = n15465 & n15466;
  assign n15468 = n15464 & n15467;
  assign n15469 = n15454 & n15458;
  assign n15470 = ~n416 & ~n1034;
  assign n15471 = ~n268 & ~n1031;
  assign n15472 = n15470 & n15471;
  assign n15473 = n15469 & n15472;
  assign n15474 = n15455 & n54812;
  assign n15475 = ~n1031 & n54446;
  assign n15476 = ~n1044 & n15475;
  assign n15477 = ~n416 & n15476;
  assign n15478 = ~n1492 & n15477;
  assign n15479 = ~n1034 & n15478;
  assign n15480 = ~n833 & n15479;
  assign n15481 = ~n268 & n15480;
  assign n15482 = ~n585 & n15481;
  assign n15483 = n54446 & n54813;
  assign n15484 = ~n356 & ~n612;
  assign n15485 = ~n498 & ~n851;
  assign n15486 = ~n356 & ~n498;
  assign n15487 = ~n612 & ~n851;
  assign n15488 = n15486 & n15487;
  assign n15489 = ~n498 & ~n612;
  assign n15490 = ~n356 & ~n851;
  assign n15491 = n15489 & n15490;
  assign n15492 = n15484 & n15485;
  assign n15493 = ~n751 & ~n851;
  assign n15494 = ~n405 & ~n612;
  assign n15495 = n15486 & n15494;
  assign n15496 = n15493 & n15495;
  assign n15497 = n13375 & n54815;
  assign n15498 = ~n405 & n54198;
  assign n15499 = ~n851 & n15498;
  assign n15500 = ~n612 & n15499;
  assign n15501 = ~n498 & n15500;
  assign n15502 = ~n356 & n15501;
  assign n15503 = ~n751 & n15502;
  assign n15504 = n54198 & n54816;
  assign n15505 = n54814 & n54817;
  assign n15506 = n208 & n54627;
  assign n15507 = n2256 & n15506;
  assign n15508 = n53919 & n15507;
  assign n15509 = n53944 & n15508;
  assign n15510 = n54814 & n15509;
  assign n15511 = n54817 & n15510;
  assign n15512 = ~n1065 & n15511;
  assign n15513 = ~n1703 & n15512;
  assign n15514 = ~n311 & n15513;
  assign n15515 = ~n1234 & n15514;
  assign n15516 = ~n514 & n15515;
  assign n15517 = ~n423 & n15516;
  assign n15518 = ~n340 & n15517;
  assign n15519 = ~n651 & n15518;
  assign n15520 = ~n789 & n15519;
  assign n15521 = n54811 & n15505;
  assign n15522 = n54808 & n54818;
  assign n15523 = n53573 & n54785;
  assign n15524 = n54117 & n15523;
  assign n15525 = n54802 & n15524;
  assign n15526 = n53470 & n15525;
  assign n15527 = n54818 & n15526;
  assign n15528 = n54801 & n15527;
  assign n15529 = n54808 & n15528;
  assign n15530 = ~n1490 & n15529;
  assign n15531 = n15314 & n15530;
  assign n15532 = ~n105 & n15531;
  assign n15533 = ~n824 & n15532;
  assign n15534 = ~n419 & n15533;
  assign n15535 = ~n754 & n15534;
  assign n15536 = ~n614 & n15535;
  assign n15537 = ~n2201 & n15536;
  assign n15538 = n54803 & n15522;
  assign n15539 = n1704 & n5651;
  assign n15540 = n7144 & n15539;
  assign n15541 = ~n342 & ~n983;
  assign n15542 = ~n922 & n15541;
  assign n15543 = n2256 & n2975;
  assign n15544 = n15542 & n15543;
  assign n15545 = n1704 & n2256;
  assign n15546 = n7144 & n15545;
  assign n15547 = ~n983 & ~n1042;
  assign n15548 = ~n922 & n15547;
  assign n15549 = ~n342 & ~n506;
  assign n15550 = n2975 & n15549;
  assign n15551 = n15548 & n15550;
  assign n15552 = n15546 & n15551;
  assign n15553 = n15540 & n15544;
  assign n15554 = ~n829 & ~n2042;
  assign n15555 = n1035 & n15554;
  assign n15556 = n1716 & n11110;
  assign n15557 = n1035 & n1716;
  assign n15558 = ~n310 & n15557;
  assign n15559 = ~n829 & n15558;
  assign n15560 = ~n2042 & n15559;
  assign n15561 = ~n588 & n15560;
  assign n15562 = n11110 & n15554;
  assign n15563 = n15557 & n15562;
  assign n15564 = n15555 & n15556;
  assign n15565 = n54540 & n54821;
  assign n15566 = n54820 & n15565;
  assign n15567 = n2814 & n3535;
  assign n15568 = n2814 & n9211;
  assign n15569 = n3535 & n15568;
  assign n15570 = n3535 & n9211;
  assign n15571 = n2814 & n15570;
  assign n15572 = n9211 & n15567;
  assign n15573 = ~n957 & ~n1681;
  assign n15574 = ~n1085 & ~n1477;
  assign n15575 = n15573 & n15574;
  assign n15576 = ~n247 & ~n590;
  assign n15577 = ~n340 & ~n975;
  assign n15578 = ~n590 & ~n975;
  assign n15579 = ~n247 & ~n340;
  assign n15580 = n15578 & n15579;
  assign n15581 = n15576 & n15577;
  assign n15582 = ~n957 & ~n1477;
  assign n15583 = ~n247 & ~n1085;
  assign n15584 = n15582 & n15583;
  assign n15585 = ~n340 & ~n1681;
  assign n15586 = n15578 & n15585;
  assign n15587 = n15584 & n15586;
  assign n15588 = ~n247 & ~n1681;
  assign n15589 = n15578 & n15588;
  assign n15590 = ~n340 & ~n1085;
  assign n15591 = n15582 & n15590;
  assign n15592 = n15589 & n15591;
  assign n15593 = n15575 & n54823;
  assign n15594 = ~n1085 & n54822;
  assign n15595 = ~n957 & n15594;
  assign n15596 = ~n1681 & n15595;
  assign n15597 = ~n1477 & n15596;
  assign n15598 = ~n247 & n15597;
  assign n15599 = ~n975 & n15598;
  assign n15600 = ~n340 & n15599;
  assign n15601 = ~n590 & n15600;
  assign n15602 = n54822 & n54824;
  assign n15603 = ~n182 & ~n625;
  assign n15604 = ~n182 & n421;
  assign n15605 = ~n625 & n15604;
  assign n15606 = n421 & n15603;
  assign n15607 = n53673 & n11098;
  assign n15608 = n54826 & n15607;
  assign n15609 = n54825 & n15608;
  assign n15610 = n54540 & n54826;
  assign n15611 = n2256 & n15610;
  assign n15612 = n54821 & n15611;
  assign n15613 = n54825 & n15612;
  assign n15614 = n2975 & n15613;
  assign n15615 = n53673 & n15614;
  assign n15616 = n1578 & n15615;
  assign n15617 = n7144 & n15616;
  assign n15618 = n1704 & n15617;
  assign n15619 = ~n922 & n15618;
  assign n15620 = ~n983 & n15619;
  assign n15621 = ~n1042 & n15620;
  assign n15622 = ~n513 & n15621;
  assign n15623 = ~n506 & n15622;
  assign n15624 = ~n342 & n15623;
  assign n15625 = n527 & n7144;
  assign n15626 = n15543 & n15625;
  assign n15627 = n54540 & n15626;
  assign n15628 = n54821 & n15627;
  assign n15629 = n53673 & n54826;
  assign n15630 = ~n342 & ~n922;
  assign n15631 = ~n342 & ~n1042;
  assign n15632 = ~n922 & ~n983;
  assign n15633 = n15631 & n15632;
  assign n15634 = n15547 & n15630;
  assign n15635 = n1578 & n1704;
  assign n15636 = n54828 & n15635;
  assign n15637 = n15629 & n15636;
  assign n15638 = n54825 & n15637;
  assign n15639 = n15628 & n15638;
  assign n15640 = n1578 & n7144;
  assign n15641 = n15545 & n15640;
  assign n15642 = n54540 & n15641;
  assign n15643 = n54821 & n15642;
  assign n15644 = n527 & n2975;
  assign n15645 = n54828 & n15644;
  assign n15646 = n15629 & n15645;
  assign n15647 = n54825 & n15646;
  assign n15648 = n15643 & n15647;
  assign n15649 = n15566 & n15609;
  assign n15650 = ~n1457 & ~n1535;
  assign n15651 = ~n1465 & ~n2201;
  assign n15652 = ~n1465 & ~n1535;
  assign n15653 = ~n1457 & ~n2201;
  assign n15654 = n15652 & n15653;
  assign n15655 = n15650 & n15651;
  assign n15656 = n2338 & n2454;
  assign n15657 = n54829 & n15656;
  assign n15658 = n54296 & n15657;
  assign n15659 = n3085 & n3675;
  assign n15660 = n4214 & n9982;
  assign n15661 = n15659 & n15660;
  assign n15662 = n54542 & n15661;
  assign n15663 = n2454 & n4214;
  assign n15664 = n54829 & n15663;
  assign n15665 = n54296 & n15664;
  assign n15666 = n2338 & n3085;
  assign n15667 = n3675 & n9982;
  assign n15668 = n15666 & n15667;
  assign n15669 = n54542 & n15668;
  assign n15670 = n15665 & n15669;
  assign n15671 = n2338 & n9982;
  assign n15672 = n54829 & n15671;
  assign n15673 = n54296 & n15672;
  assign n15674 = n3085 & n4214;
  assign n15675 = n2454 & n3675;
  assign n15676 = n15674 & n15675;
  assign n15677 = n54542 & n15676;
  assign n15678 = n15673 & n15677;
  assign n15679 = n15658 & n15662;
  assign n15680 = ~n353 & ~n465;
  assign n15681 = ~n750 & ~n1079;
  assign n15682 = n15680 & n15681;
  assign n15683 = ~n320 & ~n591;
  assign n15684 = n175 & n15683;
  assign n15685 = n13852 & n15684;
  assign n15686 = n175 & ~n320;
  assign n15687 = ~n295 & n15686;
  assign n15688 = ~n1079 & n15687;
  assign n15689 = ~n591 & n15688;
  assign n15690 = ~n465 & n15689;
  assign n15691 = ~n615 & n15690;
  assign n15692 = ~n353 & n15691;
  assign n15693 = ~n750 & n15692;
  assign n15694 = n15681 & n15683;
  assign n15695 = n175 & n15680;
  assign n15696 = n13852 & n15695;
  assign n15697 = n15694 & n15696;
  assign n15698 = ~n465 & ~n1079;
  assign n15699 = ~n353 & ~n591;
  assign n15700 = n15698 & n15699;
  assign n15701 = ~n320 & ~n750;
  assign n15702 = n175 & n15701;
  assign n15703 = n13852 & n15702;
  assign n15704 = n15700 & n15703;
  assign n15705 = ~n320 & ~n1079;
  assign n15706 = n15680 & n15705;
  assign n15707 = ~n591 & ~n750;
  assign n15708 = n13852 & n15707;
  assign n15709 = n175 & n15708;
  assign n15710 = n15706 & n15709;
  assign n15711 = n15682 & n15685;
  assign n15712 = n2783 & n5733;
  assign n15713 = n7004 & n11042;
  assign n15714 = n15712 & n15713;
  assign n15715 = ~n360 & ~n507;
  assign n15716 = ~n984 & n15715;
  assign n15717 = ~n166 & ~n222;
  assign n15718 = n846 & n15717;
  assign n15719 = ~n222 & ~n984;
  assign n15720 = ~n984 & n15717;
  assign n15721 = ~n166 & n15719;
  assign n15722 = n846 & n15715;
  assign n15723 = n54832 & n15722;
  assign n15724 = n15716 & n15718;
  assign n15725 = n846 & n5733;
  assign n15726 = n2783 & n7004;
  assign n15727 = n5733 & n15726;
  assign n15728 = n846 & n15727;
  assign n15729 = n846 & n2783;
  assign n15730 = n5733 & n7004;
  assign n15731 = n15729 & n15730;
  assign n15732 = n15725 & n15726;
  assign n15733 = ~n984 & n54834;
  assign n15734 = ~n166 & n15733;
  assign n15735 = ~n222 & n15734;
  assign n15736 = ~n562 & n15735;
  assign n15737 = ~n663 & n15736;
  assign n15738 = ~n507 & n15737;
  assign n15739 = ~n360 & n15738;
  assign n15740 = ~n166 & ~n360;
  assign n15741 = ~n222 & n15740;
  assign n15742 = ~n507 & ~n984;
  assign n15743 = n11042 & n15742;
  assign n15744 = n11042 & n15715;
  assign n15745 = n54832 & n15744;
  assign n15746 = n15741 & n15743;
  assign n15747 = n54834 & n54836;
  assign n15748 = n15714 & n54833;
  assign n15749 = n54831 & n54835;
  assign n15750 = n54830 & n15749;
  assign n15751 = n54552 & n15750;
  assign n15752 = n54296 & n54542;
  assign n15753 = n54552 & n15752;
  assign n15754 = n54831 & n15753;
  assign n15755 = n2454 & n15754;
  assign n15756 = n3085 & n15755;
  assign n15757 = n54835 & n15756;
  assign n15758 = n2338 & n15757;
  assign n15759 = n3675 & n15758;
  assign n15760 = n54827 & n15759;
  assign n15761 = n4214 & n15760;
  assign n15762 = ~n1465 & n15761;
  assign n15763 = ~n218 & n15762;
  assign n15764 = ~n584 & n15763;
  assign n15765 = ~n1457 & n15764;
  assign n15766 = ~n1535 & n15765;
  assign n15767 = ~n2201 & n15766;
  assign n15768 = n54827 & n15751;
  assign n15769 = ~n54819 & ~n54837;
  assign n15770 = n54819 & n54837;
  assign n15771 = ~pi8  & ~n15769;
  assign n15772 = ~n15769 & ~n15770;
  assign n15773 = ~pi8  & n15772;
  assign n15774 = ~n15770 & n15771;
  assign n15775 = ~n15769 & ~n54838;
  assign n15776 = n54780 & ~n15775;
  assign n15777 = ~n54780 & n15775;
  assign n15778 = n10458 & ~n10460;
  assign n15779 = ~n10461 & ~n15778;
  assign n15780 = n1576 & n15779;
  assign n15781 = ~n54098 & n10564;
  assign n15782 = ~n54119 & n54403;
  assign n15783 = ~n54073 & n11215;
  assign n15784 = ~n15782 & ~n15783;
  assign n15785 = ~n15781 & ~n15782;
  assign n15786 = ~n15783 & n15785;
  assign n15787 = ~n15781 & ~n15783;
  assign n15788 = ~n15782 & n15787;
  assign n15789 = ~n15781 & n15784;
  assign n15790 = ~n15780 & n54839;
  assign n15791 = ~n15777 & ~n15790;
  assign n15792 = ~n15776 & n15790;
  assign n15793 = ~n15777 & ~n15792;
  assign n15794 = ~n15776 & ~n15777;
  assign n15795 = ~n15790 & n15794;
  assign n15796 = ~n15776 & ~n15795;
  assign n15797 = ~n15776 & ~n15791;
  assign n15798 = ~n15301 & n54840;
  assign n15799 = ~n15302 & n15798;
  assign n15800 = n15303 & n54840;
  assign n15801 = ~n15301 & ~n54841;
  assign n15802 = n15217 & n54793;
  assign n15803 = ~n15230 & ~n15802;
  assign n15804 = ~n15801 & n15803;
  assign n15805 = ~n15230 & ~n15804;
  assign n15806 = n15204 & ~n15208;
  assign n15807 = ~n15204 & ~n15209;
  assign n15808 = n15208 & ~n15209;
  assign n15809 = ~n15807 & ~n15808;
  assign n15810 = ~n15209 & ~n15806;
  assign n15811 = ~n15805 & ~n54842;
  assign n15812 = n15805 & n54842;
  assign n15813 = ~n15811 & ~n15812;
  assign n15814 = n11279 & n14020;
  assign n15815 = ~n53962 & n11267;
  assign n15816 = ~n53970 & n54410;
  assign n15817 = ~n53930 & n12584;
  assign n15818 = ~n15816 & ~n15817;
  assign n15819 = ~n15815 & ~n15816;
  assign n15820 = ~n15817 & n15819;
  assign n15821 = ~n15815 & n15818;
  assign n15822 = ~n11279 & n54843;
  assign n15823 = ~n14020 & n54843;
  assign n15824 = ~n15822 & ~n15823;
  assign n15825 = ~n15814 & n54843;
  assign n15826 = pi29  & ~n54844;
  assign n15827 = ~pi29  & n54844;
  assign n15828 = ~n15826 & ~n15827;
  assign n15829 = n15813 & ~n15828;
  assign n15830 = ~n15811 & ~n15829;
  assign n15831 = n15214 & ~n15830;
  assign n15832 = ~n15212 & ~n15831;
  assign n15833 = n14866 & n54767;
  assign n15834 = ~n14866 & ~n14872;
  assign n15835 = ~n14866 & n54767;
  assign n15836 = ~n54767 & ~n14872;
  assign n15837 = n14866 & ~n54767;
  assign n15838 = ~n54845 & ~n54846;
  assign n15839 = ~n14872 & ~n15833;
  assign n15840 = ~n15832 & ~n54847;
  assign n15841 = ~n14872 & ~n15840;
  assign n15842 = ~n14730 & n14745;
  assign n15843 = ~n14746 & ~n15842;
  assign n15844 = ~n15841 & n15843;
  assign n15845 = n15841 & ~n15843;
  assign n15846 = n123 & n12550;
  assign n15847 = n127 & ~n53819;
  assign n15848 = n53444 & ~n53845;
  assign n15849 = n128 & ~n53799;
  assign n15850 = ~n15848 & ~n15849;
  assign n15851 = ~n15847 & ~n15848;
  assign n15852 = ~n15849 & n15851;
  assign n15853 = ~n15847 & n15850;
  assign n15854 = ~n15846 & n54848;
  assign n15855 = pi26  & ~n15854;
  assign n15856 = pi26  & ~n15855;
  assign n15857 = pi26  & n15854;
  assign n15858 = ~n15854 & ~n15855;
  assign n15859 = ~pi26  & ~n15854;
  assign n15860 = ~n54849 & ~n54850;
  assign n15861 = ~n15845 & ~n15860;
  assign n15862 = ~n15844 & ~n15845;
  assign n15863 = ~n15860 & n15862;
  assign n15864 = ~n15844 & ~n15863;
  assign n15865 = ~n15844 & ~n15861;
  assign n15866 = ~n54763 & ~n54851;
  assign n15867 = n54763 & n54851;
  assign n15868 = n90 & n11360;
  assign n15869 = ~n53685 & n14236;
  assign n15870 = ~n53741 & n54667;
  assign n15871 = ~n53712 & n14210;
  assign n15872 = ~n15870 & ~n15871;
  assign n15873 = ~n15869 & ~n15870;
  assign n15874 = ~n15871 & n15873;
  assign n15875 = ~n15869 & n15872;
  assign n15876 = ~n15868 & n54852;
  assign n15877 = pi23  & ~n15876;
  assign n15878 = pi23  & ~n15877;
  assign n15879 = pi23  & n15876;
  assign n15880 = ~n15876 & ~n15877;
  assign n15881 = ~pi23  & ~n15876;
  assign n15882 = ~n54853 & ~n54854;
  assign n15883 = ~n15867 & ~n15882;
  assign n15884 = ~n15866 & ~n15867;
  assign n15885 = ~n15882 & n15884;
  assign n15886 = ~n15866 & ~n15885;
  assign n15887 = ~n15866 & ~n15883;
  assign n15888 = ~n54762 & ~n54855;
  assign n15889 = ~n14839 & ~n15888;
  assign n15890 = n14798 & ~n14799;
  assign n15891 = n14796 & n14798;
  assign n15892 = ~n14796 & ~n14799;
  assign n15893 = ~n14796 & ~n14798;
  assign n15894 = n14796 & ~n14798;
  assign n15895 = ~n14799 & ~n15894;
  assign n15896 = ~n54856 & ~n54857;
  assign n15897 = ~n15889 & n54858;
  assign n15898 = n15889 & ~n54858;
  assign n15899 = n54351 & n14413;
  assign n15900 = ~n53634 & n54719;
  assign n15901 = ~n54717 & n54718;
  assign n15902 = ~n2325 & n15901;
  assign n15903 = ~n15900 & ~n15902;
  assign n15904 = ~n15899 & n15903;
  assign n15905 = pi20  & ~n15904;
  assign n15906 = pi20  & ~n15905;
  assign n15907 = pi20  & n15904;
  assign n15908 = ~n15904 & ~n15905;
  assign n15909 = ~pi20  & ~n15904;
  assign n15910 = ~n54859 & ~n54860;
  assign n15911 = ~n15898 & ~n15910;
  assign n15912 = ~n15897 & ~n15898;
  assign n15913 = ~n15910 & n15912;
  assign n15914 = ~n15897 & ~n15913;
  assign n15915 = ~n15897 & ~n15911;
  assign n15916 = ~n54756 & ~n54861;
  assign n15917 = n54756 & n54861;
  assign n15918 = ~n15916 & ~n15917;
  assign n15919 = n11242 & n14413;
  assign n15920 = ~n53650 & n54719;
  assign n15921 = ~n54716 & n54717;
  assign n15922 = ~n2325 & n15921;
  assign n15923 = ~n53634 & n15901;
  assign n15924 = ~n15922 & ~n15923;
  assign n15925 = ~n15920 & ~n15923;
  assign n15926 = ~n15922 & n15925;
  assign n15927 = ~n15920 & n15924;
  assign n15928 = ~n14413 & n54862;
  assign n15929 = ~n11242 & n54862;
  assign n15930 = ~n15928 & ~n15929;
  assign n15931 = ~n15919 & n54862;
  assign n15932 = pi20  & ~n54863;
  assign n15933 = ~pi20  & n54863;
  assign n15934 = ~n15932 & ~n15933;
  assign n15935 = n15882 & ~n15884;
  assign n15936 = n15884 & ~n15885;
  assign n15937 = ~n15882 & ~n15885;
  assign n15938 = ~n15936 & ~n15937;
  assign n15939 = ~n15885 & ~n15935;
  assign n15940 = n15832 & n54847;
  assign n15941 = ~n15840 & ~n15940;
  assign n15942 = n123 & n12938;
  assign n15943 = n128 & ~n53819;
  assign n15944 = n53444 & ~n53860;
  assign n15945 = n127 & ~n53845;
  assign n15946 = ~n15944 & ~n15945;
  assign n15947 = ~n15943 & ~n15944;
  assign n15948 = ~n15945 & n15947;
  assign n15949 = ~n15943 & n15946;
  assign n15950 = ~n123 & n54865;
  assign n15951 = ~n12938 & n54865;
  assign n15952 = ~n15950 & ~n15951;
  assign n15953 = ~n15942 & n54865;
  assign n15954 = pi26  & ~n54866;
  assign n15955 = ~pi26  & n54866;
  assign n15956 = ~n15954 & ~n15955;
  assign n15957 = n15941 & ~n15956;
  assign n15958 = ~n15941 & n15956;
  assign n15959 = ~n15957 & ~n15958;
  assign n15960 = ~n15214 & n15830;
  assign n15961 = ~n15831 & ~n15960;
  assign n15962 = n11279 & n14263;
  assign n15963 = ~n53930 & n11267;
  assign n15964 = ~n53962 & n54410;
  assign n15965 = ~n53907 & n12584;
  assign n15966 = ~n15964 & ~n15965;
  assign n15967 = ~n15963 & ~n15964;
  assign n15968 = ~n15965 & n15967;
  assign n15969 = ~n15963 & n15966;
  assign n15970 = ~n11279 & n54867;
  assign n15971 = ~n14263 & n54867;
  assign n15972 = ~n15970 & ~n15971;
  assign n15973 = ~n15962 & n54867;
  assign n15974 = pi29  & ~n54868;
  assign n15975 = ~pi29  & n54868;
  assign n15976 = ~n15974 & ~n15975;
  assign n15977 = n15961 & ~n15976;
  assign n15978 = n123 & n12918;
  assign n15979 = n127 & ~n53860;
  assign n15980 = n53444 & ~n53888;
  assign n15981 = n128 & ~n53845;
  assign n15982 = ~n15980 & ~n15981;
  assign n15983 = ~n15979 & ~n15980;
  assign n15984 = ~n15981 & n15983;
  assign n15985 = ~n15979 & n15982;
  assign n15986 = ~n15978 & n54869;
  assign n15987 = pi26  & ~n15986;
  assign n15988 = pi26  & ~n15987;
  assign n15989 = pi26  & n15986;
  assign n15990 = ~n15986 & ~n15987;
  assign n15991 = ~pi26  & ~n15986;
  assign n15992 = ~n54870 & ~n54871;
  assign n15993 = ~n15961 & n15976;
  assign n15994 = ~n15992 & ~n15993;
  assign n15995 = ~n15977 & ~n15993;
  assign n15996 = ~n15992 & n15995;
  assign n15997 = ~n15977 & ~n15996;
  assign n15998 = ~n15977 & ~n15994;
  assign n15999 = n15959 & ~n54872;
  assign n16000 = ~n15957 & ~n15999;
  assign n16001 = n15860 & ~n15862;
  assign n16002 = n15862 & ~n15863;
  assign n16003 = ~n15860 & ~n15863;
  assign n16004 = ~n16002 & ~n16003;
  assign n16005 = ~n15863 & ~n16001;
  assign n16006 = ~n16000 & ~n54873;
  assign n16007 = n16000 & n54873;
  assign n16008 = n90 & n11889;
  assign n16009 = ~n53712 & n14236;
  assign n16010 = ~n53774 & n54667;
  assign n16011 = ~n53741 & n14210;
  assign n16012 = ~n16010 & ~n16011;
  assign n16013 = ~n16009 & ~n16010;
  assign n16014 = ~n16011 & n16013;
  assign n16015 = ~n16009 & n16012;
  assign n16016 = ~n16008 & n54874;
  assign n16017 = pi23  & ~n16016;
  assign n16018 = pi23  & ~n16017;
  assign n16019 = pi23  & n16016;
  assign n16020 = ~n16016 & ~n16017;
  assign n16021 = ~pi23  & ~n16016;
  assign n16022 = ~n54875 & ~n54876;
  assign n16023 = ~n16007 & ~n16022;
  assign n16024 = ~n16006 & ~n16007;
  assign n16025 = ~n16022 & n16024;
  assign n16026 = ~n16006 & ~n16025;
  assign n16027 = ~n16006 & ~n16023;
  assign n16028 = ~n54864 & ~n54877;
  assign n16029 = n54864 & n54877;
  assign n16030 = n11286 & n14413;
  assign n16031 = ~n53650 & n15901;
  assign n16032 = ~n53657 & n54719;
  assign n16033 = ~n53634 & n15921;
  assign n16034 = ~n16032 & ~n16033;
  assign n16035 = ~n16031 & ~n16032;
  assign n16036 = ~n16033 & n16035;
  assign n16037 = ~n16031 & n16034;
  assign n16038 = ~n16030 & n54878;
  assign n16039 = pi20  & ~n16038;
  assign n16040 = pi20  & ~n16039;
  assign n16041 = pi20  & n16038;
  assign n16042 = ~n16038 & ~n16039;
  assign n16043 = ~pi20  & ~n16038;
  assign n16044 = ~n54879 & ~n54880;
  assign n16045 = ~n16029 & ~n16044;
  assign n16046 = ~n16028 & ~n16029;
  assign n16047 = ~n16044 & n16046;
  assign n16048 = ~n16028 & ~n16047;
  assign n16049 = ~n16028 & ~n16045;
  assign n16050 = ~n15934 & ~n54881;
  assign n16051 = n54762 & n54855;
  assign n16052 = ~n15888 & ~n16051;
  assign n16053 = n15934 & n54881;
  assign n16054 = ~n16050 & ~n16053;
  assign n16055 = n16052 & n16054;
  assign n16056 = ~n16050 & ~n16055;
  assign n16057 = n15910 & ~n15912;
  assign n16058 = n15912 & ~n15913;
  assign n16059 = ~n15910 & ~n15913;
  assign n16060 = ~n16058 & ~n16059;
  assign n16061 = ~n15913 & ~n16057;
  assign n16062 = ~n16056 & ~n54882;
  assign n16063 = n16056 & n54882;
  assign n16064 = ~n16062 & ~n16063;
  assign n16065 = ~n16052 & ~n16054;
  assign n16066 = ~n16055 & ~n16065;
  assign n16067 = pi14  & ~pi15 ;
  assign n16068 = ~pi14  & pi15 ;
  assign n16069 = ~pi14  & ~pi15 ;
  assign n16070 = pi14  & pi15 ;
  assign n16071 = ~n16069 & ~n16070;
  assign n16072 = ~n16067 & ~n16068;
  assign n16073 = pi16  & ~pi17 ;
  assign n16074 = ~pi16  & pi17 ;
  assign n16075 = ~pi16  & ~pi17 ;
  assign n16076 = pi16  & pi17 ;
  assign n16077 = ~n16075 & ~n16076;
  assign n16078 = ~n16073 & ~n16074;
  assign n16079 = n54883 & n54884;
  assign n16080 = ~n10547 & n16079;
  assign n16081 = pi15  & ~pi16 ;
  assign n16082 = ~pi15  & pi16 ;
  assign n16083 = ~pi15  & ~pi16 ;
  assign n16084 = pi15  & pi16 ;
  assign n16085 = ~n16083 & ~n16084;
  assign n16086 = ~n16081 & ~n16082;
  assign n16087 = ~n54883 & ~n54885;
  assign n16088 = ~n54883 & n54884;
  assign n16089 = ~n54885 & n16088;
  assign n16090 = n54884 & n16087;
  assign n16091 = ~n16080 & ~n54886;
  assign n16092 = ~n2325 & n54886;
  assign n16093 = ~n10551 & ~n16092;
  assign n16094 = ~n16079 & ~n16092;
  assign n16095 = ~n16093 & ~n16094;
  assign n16096 = ~n2325 & ~n16091;
  assign n16097 = pi17  & ~n54887;
  assign n16098 = ~pi17  & n54887;
  assign n16099 = ~n16097 & ~n16098;
  assign n16100 = n90 & n11913;
  assign n16101 = ~n53774 & n14210;
  assign n16102 = ~n53799 & n54667;
  assign n16103 = ~n53741 & n14236;
  assign n16104 = ~n16102 & ~n16103;
  assign n16105 = ~n16101 & ~n16102;
  assign n16106 = ~n16103 & n16105;
  assign n16107 = ~n16101 & n16104;
  assign n16108 = ~n16100 & n54888;
  assign n16109 = pi23  & ~n16108;
  assign n16110 = ~n16108 & ~n16109;
  assign n16111 = ~pi23  & ~n16108;
  assign n16112 = pi23  & ~n16109;
  assign n16113 = pi23  & n16108;
  assign n16114 = ~n54889 & ~n54890;
  assign n16115 = ~n15959 & n54872;
  assign n16116 = ~n15999 & ~n16115;
  assign n16117 = ~n16114 & n16116;
  assign n16118 = n16114 & ~n16116;
  assign n16119 = ~n16114 & ~n16117;
  assign n16120 = ~n16114 & ~n16116;
  assign n16121 = n16116 & ~n16117;
  assign n16122 = n16114 & n16116;
  assign n16123 = ~n54891 & ~n54892;
  assign n16124 = ~n16117 & ~n16118;
  assign n16125 = n15992 & ~n15995;
  assign n16126 = n15995 & ~n15996;
  assign n16127 = ~n15992 & ~n15996;
  assign n16128 = ~n16126 & ~n16127;
  assign n16129 = ~n15996 & ~n16125;
  assign n16130 = ~n15813 & n15828;
  assign n16131 = ~n15829 & ~n16130;
  assign n16132 = ~n15303 & ~n54840;
  assign n16133 = n54840 & ~n54841;
  assign n16134 = ~n15302 & n15801;
  assign n16135 = ~n16133 & ~n16134;
  assign n16136 = ~n54841 & ~n16132;
  assign n16137 = n10462 & ~n10464;
  assign n16138 = ~n10465 & ~n16137;
  assign n16139 = n1576 & n16138;
  assign n16140 = ~n54098 & n54403;
  assign n16141 = ~n54050 & n11215;
  assign n16142 = ~n54073 & n10564;
  assign n16143 = ~n16141 & ~n16142;
  assign n16144 = ~n16140 & n16143;
  assign n16145 = ~n16139 & ~n16140;
  assign n16146 = ~n16142 & n16145;
  assign n16147 = ~n16141 & n16146;
  assign n16148 = ~n16139 & n16144;
  assign n16149 = ~n54895 & ~n54896;
  assign n16150 = n11279 & n14688;
  assign n16151 = ~n54005 & n11267;
  assign n16152 = ~n54034 & n54410;
  assign n16153 = ~n53970 & n12584;
  assign n16154 = ~n16152 & ~n16153;
  assign n16155 = ~n16151 & ~n16152;
  assign n16156 = ~n16153 & n16155;
  assign n16157 = ~n16151 & n16154;
  assign n16158 = ~n16150 & n54897;
  assign n16159 = pi29  & ~n16158;
  assign n16160 = ~n16158 & ~n16159;
  assign n16161 = ~pi29  & ~n16158;
  assign n16162 = pi29  & ~n16159;
  assign n16163 = pi29  & n16158;
  assign n16164 = ~n54898 & ~n54899;
  assign n16165 = n54895 & n54896;
  assign n16166 = ~n54895 & ~n16149;
  assign n16167 = ~n54895 & n54896;
  assign n16168 = ~n54896 & ~n16149;
  assign n16169 = n54895 & ~n54896;
  assign n16170 = ~n54900 & ~n54901;
  assign n16171 = ~n16149 & ~n16165;
  assign n16172 = ~n16164 & ~n54902;
  assign n16173 = ~n16149 & ~n16172;
  assign n16174 = n15801 & ~n15803;
  assign n16175 = ~n15804 & ~n16174;
  assign n16176 = ~n16173 & n16175;
  assign n16177 = n16173 & ~n16175;
  assign n16178 = n11279 & n14708;
  assign n16179 = ~n54005 & n54410;
  assign n16180 = ~n53970 & n11267;
  assign n16181 = ~n53962 & n12584;
  assign n16182 = ~n16180 & ~n16181;
  assign n16183 = ~n16179 & ~n16180;
  assign n16184 = ~n16181 & n16183;
  assign n16185 = ~n16179 & n16182;
  assign n16186 = ~n16178 & n54903;
  assign n16187 = pi29  & ~n16186;
  assign n16188 = pi29  & ~n16187;
  assign n16189 = pi29  & n16186;
  assign n16190 = ~n16186 & ~n16187;
  assign n16191 = ~pi29  & ~n16186;
  assign n16192 = ~n54904 & ~n54905;
  assign n16193 = ~n16177 & ~n16192;
  assign n16194 = ~n16176 & ~n16177;
  assign n16195 = ~n16192 & n16194;
  assign n16196 = ~n16176 & ~n16195;
  assign n16197 = ~n16176 & ~n16193;
  assign n16198 = n16131 & ~n54906;
  assign n16199 = ~n16131 & n54906;
  assign n16200 = n123 & n13336;
  assign n16201 = n127 & ~n53888;
  assign n16202 = n53444 & ~n53907;
  assign n16203 = n128 & ~n53860;
  assign n16204 = ~n16202 & ~n16203;
  assign n16205 = ~n16201 & ~n16202;
  assign n16206 = ~n16203 & n16205;
  assign n16207 = ~n16201 & n16204;
  assign n16208 = ~n16200 & n54907;
  assign n16209 = pi26  & ~n16208;
  assign n16210 = pi26  & ~n16209;
  assign n16211 = pi26  & n16208;
  assign n16212 = ~n16208 & ~n16209;
  assign n16213 = ~pi26  & ~n16208;
  assign n16214 = ~n54908 & ~n54909;
  assign n16215 = ~n16199 & ~n16214;
  assign n16216 = ~n16198 & ~n16199;
  assign n16217 = ~n16214 & n16216;
  assign n16218 = ~n16198 & ~n16217;
  assign n16219 = ~n16198 & ~n16215;
  assign n16220 = ~n54894 & ~n54910;
  assign n16221 = n54894 & n54910;
  assign n16222 = n90 & n12690;
  assign n16223 = ~n53774 & n14236;
  assign n16224 = ~n53819 & n54667;
  assign n16225 = ~n53799 & n14210;
  assign n16226 = ~n16224 & ~n16225;
  assign n16227 = ~n16223 & ~n16224;
  assign n16228 = ~n16225 & n16227;
  assign n16229 = ~n16223 & n16226;
  assign n16230 = ~n16222 & n54911;
  assign n16231 = pi23  & ~n16230;
  assign n16232 = pi23  & ~n16231;
  assign n16233 = pi23  & n16230;
  assign n16234 = ~n16230 & ~n16231;
  assign n16235 = ~pi23  & ~n16230;
  assign n16236 = ~n54912 & ~n54913;
  assign n16237 = ~n16221 & ~n16236;
  assign n16238 = ~n16220 & ~n16221;
  assign n16239 = ~n16236 & n16238;
  assign n16240 = ~n16220 & ~n16239;
  assign n16241 = ~n16220 & ~n16237;
  assign n16242 = ~n54893 & ~n54914;
  assign n16243 = ~n16117 & ~n16242;
  assign n16244 = n16024 & ~n16025;
  assign n16245 = n16022 & n16024;
  assign n16246 = ~n16022 & ~n16025;
  assign n16247 = ~n16022 & ~n16024;
  assign n16248 = n16022 & ~n16024;
  assign n16249 = ~n16025 & ~n16248;
  assign n16250 = ~n54915 & ~n54916;
  assign n16251 = ~n16243 & n54917;
  assign n16252 = n16243 & ~n54917;
  assign n16253 = n11213 & n14413;
  assign n16254 = ~n53650 & n15921;
  assign n16255 = ~n53685 & n54719;
  assign n16256 = ~n53657 & n15901;
  assign n16257 = ~n16255 & ~n16256;
  assign n16258 = ~n16254 & n16257;
  assign n16259 = ~n16253 & n16258;
  assign n16260 = pi20  & ~n16259;
  assign n16261 = pi20  & ~n16260;
  assign n16262 = pi20  & n16259;
  assign n16263 = ~n16259 & ~n16260;
  assign n16264 = ~pi20  & ~n16259;
  assign n16265 = ~n54918 & ~n54919;
  assign n16266 = ~n16252 & ~n16265;
  assign n16267 = ~n16251 & ~n16252;
  assign n16268 = ~n16265 & n16267;
  assign n16269 = ~n16251 & ~n16268;
  assign n16270 = ~n16251 & ~n16266;
  assign n16271 = ~n16099 & ~n54920;
  assign n16272 = n16099 & n54920;
  assign n16273 = n16044 & ~n16046;
  assign n16274 = n16046 & ~n16047;
  assign n16275 = ~n16044 & ~n16047;
  assign n16276 = ~n16274 & ~n16275;
  assign n16277 = ~n16047 & ~n16273;
  assign n16278 = ~n16272 & ~n54921;
  assign n16279 = ~n16271 & ~n16272;
  assign n16280 = ~n54921 & n16279;
  assign n16281 = ~n16271 & ~n16280;
  assign n16282 = ~n16271 & ~n16278;
  assign n16283 = n16066 & ~n54922;
  assign n16284 = n54921 & ~n16279;
  assign n16285 = ~n54921 & ~n16280;
  assign n16286 = n16279 & ~n16280;
  assign n16287 = ~n16285 & ~n16286;
  assign n16288 = ~n16280 & ~n16284;
  assign n16289 = n54893 & n54914;
  assign n16290 = ~n16242 & ~n16289;
  assign n16291 = n11380 & n14413;
  assign n16292 = ~n53685 & n15901;
  assign n16293 = ~n53657 & n15921;
  assign n16294 = ~n53712 & n54719;
  assign n16295 = ~n16293 & ~n16294;
  assign n16296 = ~n16292 & ~n16294;
  assign n16297 = ~n16293 & n16296;
  assign n16298 = ~n16292 & n16295;
  assign n16299 = ~n14413 & n54924;
  assign n16300 = ~n11380 & n54924;
  assign n16301 = ~n16299 & ~n16300;
  assign n16302 = ~n16291 & n54924;
  assign n16303 = pi20  & ~n54925;
  assign n16304 = ~pi20  & n54925;
  assign n16305 = ~n16303 & ~n16304;
  assign n16306 = n16290 & ~n16305;
  assign n16307 = ~n16290 & n16305;
  assign n16308 = ~n16306 & ~n16307;
  assign n16309 = n16236 & ~n16238;
  assign n16310 = n16238 & ~n16239;
  assign n16311 = ~n16236 & ~n16239;
  assign n16312 = ~n16310 & ~n16311;
  assign n16313 = ~n16239 & ~n16309;
  assign n16314 = n123 & n13360;
  assign n16315 = n127 & ~n53907;
  assign n16316 = n53444 & ~n53930;
  assign n16317 = n128 & ~n53888;
  assign n16318 = ~n16316 & ~n16317;
  assign n16319 = ~n16315 & ~n16316;
  assign n16320 = ~n16317 & n16319;
  assign n16321 = ~n16315 & n16318;
  assign n16322 = ~n123 & n54927;
  assign n16323 = ~n13360 & n54927;
  assign n16324 = ~n16322 & ~n16323;
  assign n16325 = ~n16314 & n54927;
  assign n16326 = pi26  & ~n54928;
  assign n16327 = ~pi26  & n54928;
  assign n16328 = ~n16326 & ~n16327;
  assign n16329 = n16192 & ~n16194;
  assign n16330 = n16194 & ~n16195;
  assign n16331 = ~n16192 & ~n16195;
  assign n16332 = ~n16330 & ~n16331;
  assign n16333 = ~n16195 & ~n16329;
  assign n16334 = ~n16328 & ~n54929;
  assign n16335 = n16328 & n54929;
  assign n16336 = ~n16334 & ~n16335;
  assign n16337 = ~n562 & ~n1191;
  assign n16338 = ~n1085 & ~n1191;
  assign n16339 = ~n562 & n16338;
  assign n16340 = ~n562 & ~n1085;
  assign n16341 = ~n1191 & n16340;
  assign n16342 = ~n1085 & n16337;
  assign n16343 = ~n618 & ~n660;
  assign n16344 = ~n269 & ~n308;
  assign n16345 = n16343 & n16344;
  assign n16346 = n3672 & n4258;
  assign n16347 = n16345 & n16346;
  assign n16348 = n54930 & n16347;
  assign n16349 = n4799 & n5273;
  assign n16350 = ~n514 & ~n852;
  assign n16351 = n13428 & n16350;
  assign n16352 = n16349 & n16351;
  assign n16353 = n54821 & n16352;
  assign n16354 = ~n1062 & ~n1477;
  assign n16355 = n16350 & n16354;
  assign n16356 = n16345 & n16355;
  assign n16357 = n54930 & n16356;
  assign n16358 = n1265 & n4258;
  assign n16359 = n3672 & n4799;
  assign n16360 = n16358 & n16359;
  assign n16361 = n54821 & n16360;
  assign n16362 = n16357 & n16361;
  assign n16363 = n16348 & n16353;
  assign n16364 = n54802 & n54931;
  assign n16365 = ~n247 & ~n510;
  assign n16366 = ~n948 & n16365;
  assign n16367 = n53719 & n16366;
  assign n16368 = n54439 & n13476;
  assign n16369 = n16367 & n16368;
  assign n16370 = n712 & ~n1457;
  assign n16371 = n712 & n2058;
  assign n16372 = ~n1457 & n16371;
  assign n16373 = ~n1457 & n2058;
  assign n16374 = n712 & n16373;
  assign n16375 = n2058 & n16370;
  assign n16376 = ~n274 & ~n585;
  assign n16377 = n6530 & n16376;
  assign n16378 = n7144 & n12286;
  assign n16379 = n16377 & n16378;
  assign n16380 = n54932 & n16379;
  assign n16381 = n54439 & n54932;
  assign n16382 = n53719 & n16381;
  assign n16383 = n6530 & n16382;
  assign n16384 = n12286 & n16383;
  assign n16385 = n5652 & n16384;
  assign n16386 = n7144 & n16385;
  assign n16387 = ~n948 & n16386;
  assign n16388 = ~n247 & n16387;
  assign n16389 = ~n274 & n16388;
  assign n16390 = ~n510 & n16389;
  assign n16391 = ~n590 & n16390;
  assign n16392 = ~n585 & n16391;
  assign n16393 = ~n247 & ~n585;
  assign n16394 = ~n948 & n16393;
  assign n16395 = n53719 & n16394;
  assign n16396 = n16368 & n16395;
  assign n16397 = ~n274 & ~n510;
  assign n16398 = n6530 & n16397;
  assign n16399 = n16378 & n16398;
  assign n16400 = n54932 & n16399;
  assign n16401 = n16396 & n16400;
  assign n16402 = n15576 & n16376;
  assign n16403 = ~n510 & ~n948;
  assign n16404 = n5652 & n16403;
  assign n16405 = n16365 & n16376;
  assign n16406 = ~n590 & ~n948;
  assign n16407 = n5652 & n16406;
  assign n16408 = n16405 & n16407;
  assign n16409 = n16402 & n16404;
  assign n16410 = n53719 & n54439;
  assign n16411 = n54934 & n16410;
  assign n16412 = n6530 & n7144;
  assign n16413 = n12286 & n16412;
  assign n16414 = n54932 & n16413;
  assign n16415 = n16411 & n16414;
  assign n16416 = n16369 & n16380;
  assign n16417 = n53876 & n54933;
  assign n16418 = n16364 & n16417;
  assign n16419 = n4799 & n54930;
  assign n16420 = n54821 & n16419;
  assign n16421 = n53876 & n16420;
  assign n16422 = n54802 & n16421;
  assign n16423 = n54507 & n16422;
  assign n16424 = n54933 & n16423;
  assign n16425 = n1265 & n16424;
  assign n16426 = n4258 & n16425;
  assign n16427 = n3672 & n16426;
  assign n16428 = ~n1062 & n16427;
  assign n16429 = ~n1477 & n16428;
  assign n16430 = ~n308 & n16429;
  assign n16431 = ~n660 & n16430;
  assign n16432 = ~n618 & n16431;
  assign n16433 = ~n514 & n16432;
  assign n16434 = ~n852 & n16433;
  assign n16435 = ~n269 & n16434;
  assign n16436 = n54507 & n16418;
  assign n16437 = n54819 & ~n54935;
  assign n16438 = ~n54819 & n54935;
  assign n16439 = ~n16437 & ~n16438;
  assign n16440 = ~n423 & ~n448;
  assign n16441 = ~n448 & ~n911;
  assign n16442 = ~n423 & n16441;
  assign n16443 = ~n911 & n16440;
  assign n16444 = n2577 & n3638;
  assign n16445 = n54936 & n16444;
  assign n16446 = n53606 & n4916;
  assign n16447 = n16445 & n16446;
  assign n16448 = n3780 & n7647;
  assign n16449 = n9466 & n16448;
  assign n16450 = n53789 & n16449;
  assign n16451 = n2577 & n3780;
  assign n16452 = n54936 & n16451;
  assign n16453 = n16446 & n16452;
  assign n16454 = n3638 & n7647;
  assign n16455 = n9466 & n16454;
  assign n16456 = n53789 & n16455;
  assign n16457 = n16453 & n16456;
  assign n16458 = ~n495 & ~n911;
  assign n16459 = ~n1769 & n16458;
  assign n16460 = ~n448 & ~n1997;
  assign n16461 = ~n206 & ~n1196;
  assign n16462 = n16460 & n16461;
  assign n16463 = n16459 & n16462;
  assign n16464 = n16446 & n16463;
  assign n16465 = ~n423 & ~n894;
  assign n16466 = n2577 & n16465;
  assign n16467 = n3780 & n16466;
  assign n16468 = n53789 & n16467;
  assign n16469 = n16464 & n16468;
  assign n16470 = n16447 & n16450;
  assign n16471 = ~n742 & ~n822;
  assign n16472 = ~n742 & ~n754;
  assign n16473 = ~n822 & n16472;
  assign n16474 = ~n754 & n16471;
  assign n16475 = ~n274 & ~n1031;
  assign n16476 = n1866 & n3821;
  assign n16477 = n16475 & n16476;
  assign n16478 = ~n1031 & n16476;
  assign n16479 = ~n742 & n16478;
  assign n16480 = ~n822 & n16479;
  assign n16481 = ~n274 & n16480;
  assign n16482 = ~n754 & n16481;
  assign n16483 = ~n742 & ~n1031;
  assign n16484 = ~n754 & n16483;
  assign n16485 = ~n274 & ~n822;
  assign n16486 = n1866 & n16485;
  assign n16487 = n3821 & n16486;
  assign n16488 = n16484 & n16487;
  assign n16489 = n54938 & n16477;
  assign n16490 = n53776 & n54939;
  assign n16491 = n54937 & n16490;
  assign n16492 = n54378 & n16491;
  assign n16493 = n53606 & n53789;
  assign n16494 = n54378 & n16493;
  assign n16495 = n54641 & n16494;
  assign n16496 = n4916 & n16495;
  assign n16497 = n54939 & n16496;
  assign n16498 = n3780 & n16497;
  assign n16499 = n53776 & n16498;
  assign n16500 = n2577 & n16499;
  assign n16501 = ~n894 & n16500;
  assign n16502 = ~n1997 & n16501;
  assign n16503 = ~n1196 & n16502;
  assign n16504 = ~n206 & n16503;
  assign n16505 = ~n495 & n16504;
  assign n16506 = ~n911 & n16505;
  assign n16507 = ~n423 & n16506;
  assign n16508 = ~n448 & n16507;
  assign n16509 = ~n1769 & n16508;
  assign n16510 = n54641 & n16492;
  assign n16511 = ~pi2  & ~n54940;
  assign n16512 = pi2  & n54940;
  assign n16513 = pi2  & ~n54940;
  assign n16514 = ~pi2  & n54940;
  assign n16515 = ~n16513 & ~n16514;
  assign n16516 = ~n16511 & ~n16512;
  assign n16517 = ~pi5  & ~n54941;
  assign n16518 = ~n16511 & ~n16517;
  assign n16519 = n54819 & ~n16518;
  assign n16520 = ~n54819 & n16518;
  assign n16521 = n10446 & ~n10448;
  assign n16522 = ~n10449 & ~n16521;
  assign n16523 = n1576 & n16522;
  assign n16524 = ~n54154 & n10564;
  assign n16525 = ~n54132 & n11215;
  assign n16526 = ~n54163 & n54403;
  assign n16527 = ~n16525 & ~n16526;
  assign n16528 = ~n16524 & ~n16526;
  assign n16529 = ~n16525 & n16528;
  assign n16530 = ~n16524 & n16527;
  assign n16531 = ~n16523 & n54942;
  assign n16532 = ~n16520 & ~n16531;
  assign n16533 = ~n16519 & ~n16520;
  assign n16534 = ~n16531 & n16533;
  assign n16535 = ~n16519 & ~n16534;
  assign n16536 = ~n16519 & ~n16532;
  assign n16537 = ~n16437 & ~n54943;
  assign n16538 = ~n16438 & n16537;
  assign n16539 = n16439 & ~n54943;
  assign n16540 = ~n16437 & ~n54944;
  assign n16541 = ~pi8  & ~n54838;
  assign n16542 = ~n15770 & n15775;
  assign n16543 = ~n16541 & ~n16542;
  assign n16544 = ~n16540 & ~n16543;
  assign n16545 = n16540 & n16543;
  assign n16546 = n10454 & ~n10456;
  assign n16547 = ~n10457 & ~n16546;
  assign n16548 = n1576 & n16547;
  assign n16549 = ~n54119 & n10564;
  assign n16550 = ~n54098 & n11215;
  assign n16551 = ~n54132 & n54403;
  assign n16552 = ~n16550 & ~n16551;
  assign n16553 = ~n16549 & ~n16551;
  assign n16554 = ~n16550 & n16553;
  assign n16555 = ~n16549 & n16552;
  assign n16556 = ~n16548 & n54945;
  assign n16557 = ~n16545 & ~n16556;
  assign n16558 = ~n16544 & ~n16545;
  assign n16559 = ~n16556 & n16558;
  assign n16560 = ~n16544 & ~n16559;
  assign n16561 = ~n16544 & ~n16557;
  assign n16562 = n15790 & ~n15794;
  assign n16563 = ~n15790 & ~n15795;
  assign n16564 = n15794 & ~n15795;
  assign n16565 = ~n16563 & ~n16564;
  assign n16566 = ~n15795 & ~n16562;
  assign n16567 = ~n54946 & ~n54947;
  assign n16568 = n54946 & n54947;
  assign n16569 = ~n16567 & ~n16568;
  assign n16570 = n11279 & n15195;
  assign n16571 = ~n54050 & n54410;
  assign n16572 = ~n54005 & n12584;
  assign n16573 = ~n54034 & n11267;
  assign n16574 = ~n16572 & ~n16573;
  assign n16575 = ~n16571 & ~n16573;
  assign n16576 = ~n16572 & n16575;
  assign n16577 = ~n16571 & n16574;
  assign n16578 = ~n11279 & n54948;
  assign n16579 = ~n15195 & n54948;
  assign n16580 = ~n16578 & ~n16579;
  assign n16581 = ~n16570 & n54948;
  assign n16582 = pi29  & ~n54949;
  assign n16583 = ~pi29  & n54949;
  assign n16584 = ~n16582 & ~n16583;
  assign n16585 = n16569 & ~n16584;
  assign n16586 = ~n16567 & ~n16585;
  assign n16587 = n16164 & n54902;
  assign n16588 = ~n16164 & ~n16172;
  assign n16589 = ~n54902 & ~n16172;
  assign n16590 = ~n16588 & ~n16589;
  assign n16591 = ~n16172 & ~n16587;
  assign n16592 = ~n16586 & ~n54950;
  assign n16593 = n16586 & n54950;
  assign n16594 = n123 & n14263;
  assign n16595 = n127 & ~n53930;
  assign n16596 = n53444 & ~n53962;
  assign n16597 = n128 & ~n53907;
  assign n16598 = ~n16596 & ~n16597;
  assign n16599 = ~n16595 & ~n16596;
  assign n16600 = ~n16597 & n16599;
  assign n16601 = ~n16595 & n16598;
  assign n16602 = ~n16594 & n54951;
  assign n16603 = pi26  & ~n16602;
  assign n16604 = pi26  & ~n16603;
  assign n16605 = pi26  & n16602;
  assign n16606 = ~n16602 & ~n16603;
  assign n16607 = ~pi26  & ~n16602;
  assign n16608 = ~n54952 & ~n54953;
  assign n16609 = ~n16593 & ~n16608;
  assign n16610 = ~n16592 & ~n16593;
  assign n16611 = ~n16608 & n16610;
  assign n16612 = ~n16592 & ~n16611;
  assign n16613 = ~n16592 & ~n16609;
  assign n16614 = n16336 & ~n54954;
  assign n16615 = ~n16334 & ~n16614;
  assign n16616 = n16214 & ~n16216;
  assign n16617 = n16216 & ~n16217;
  assign n16618 = ~n16214 & ~n16217;
  assign n16619 = ~n16617 & ~n16618;
  assign n16620 = ~n16217 & ~n16616;
  assign n16621 = ~n16615 & ~n54955;
  assign n16622 = n16615 & n54955;
  assign n16623 = n90 & n12550;
  assign n16624 = ~n53819 & n14210;
  assign n16625 = ~n53845 & n54667;
  assign n16626 = ~n53799 & n14236;
  assign n16627 = ~n16625 & ~n16626;
  assign n16628 = ~n16624 & ~n16625;
  assign n16629 = ~n16626 & n16628;
  assign n16630 = ~n16624 & n16627;
  assign n16631 = ~n16623 & n54956;
  assign n16632 = pi23  & ~n16631;
  assign n16633 = pi23  & ~n16632;
  assign n16634 = pi23  & n16631;
  assign n16635 = ~n16631 & ~n16632;
  assign n16636 = ~pi23  & ~n16631;
  assign n16637 = ~n54957 & ~n54958;
  assign n16638 = ~n16622 & ~n16637;
  assign n16639 = ~n16621 & ~n16622;
  assign n16640 = ~n16637 & n16639;
  assign n16641 = ~n16621 & ~n16640;
  assign n16642 = ~n16621 & ~n16638;
  assign n16643 = ~n54926 & ~n54959;
  assign n16644 = n54926 & n54959;
  assign n16645 = n11360 & n14413;
  assign n16646 = ~n53685 & n15921;
  assign n16647 = ~n53741 & n54719;
  assign n16648 = ~n53712 & n15901;
  assign n16649 = ~n16647 & ~n16648;
  assign n16650 = ~n16646 & ~n16647;
  assign n16651 = ~n16648 & n16650;
  assign n16652 = ~n16646 & n16649;
  assign n16653 = ~n16645 & n54960;
  assign n16654 = pi20  & ~n16653;
  assign n16655 = pi20  & ~n16654;
  assign n16656 = pi20  & n16653;
  assign n16657 = ~n16653 & ~n16654;
  assign n16658 = ~pi20  & ~n16653;
  assign n16659 = ~n54961 & ~n54962;
  assign n16660 = ~n16644 & ~n16659;
  assign n16661 = ~n16643 & ~n16644;
  assign n16662 = ~n16659 & n16661;
  assign n16663 = ~n16643 & ~n16662;
  assign n16664 = ~n16643 & ~n16660;
  assign n16665 = n16308 & ~n54963;
  assign n16666 = ~n16306 & ~n16665;
  assign n16667 = n16265 & ~n16267;
  assign n16668 = n16267 & ~n16268;
  assign n16669 = ~n16265 & ~n16268;
  assign n16670 = ~n16668 & ~n16669;
  assign n16671 = ~n16268 & ~n16667;
  assign n16672 = ~n16666 & ~n54964;
  assign n16673 = n16666 & n54964;
  assign n16674 = n54351 & n16079;
  assign n16675 = ~n53634 & n54886;
  assign n16676 = ~n54883 & n54885;
  assign n16677 = ~n2325 & n16676;
  assign n16678 = ~n16675 & ~n16677;
  assign n16679 = ~n16674 & n16678;
  assign n16680 = pi17  & ~n16679;
  assign n16681 = pi17  & ~n16680;
  assign n16682 = pi17  & n16679;
  assign n16683 = ~n16679 & ~n16680;
  assign n16684 = ~pi17  & ~n16679;
  assign n16685 = ~n54965 & ~n54966;
  assign n16686 = ~n16673 & ~n16685;
  assign n16687 = ~n16672 & ~n16673;
  assign n16688 = ~n16685 & n16687;
  assign n16689 = ~n16672 & ~n16688;
  assign n16690 = ~n16672 & ~n16686;
  assign n16691 = ~n54923 & ~n54967;
  assign n16692 = n54923 & n54967;
  assign n16693 = ~n16691 & ~n16692;
  assign n16694 = n11242 & n16079;
  assign n16695 = ~n53650 & n54886;
  assign n16696 = n54883 & ~n54884;
  assign n16697 = ~n2325 & n16696;
  assign n16698 = ~n53634 & n16676;
  assign n16699 = ~n16697 & ~n16698;
  assign n16700 = ~n16695 & ~n16698;
  assign n16701 = ~n16697 & n16700;
  assign n16702 = ~n16695 & n16699;
  assign n16703 = ~n16079 & n54968;
  assign n16704 = ~n11242 & n54968;
  assign n16705 = ~n16703 & ~n16704;
  assign n16706 = ~n16694 & n54968;
  assign n16707 = pi17  & ~n54969;
  assign n16708 = ~pi17  & n54969;
  assign n16709 = ~n16707 & ~n16708;
  assign n16710 = n16659 & ~n16661;
  assign n16711 = n16661 & ~n16662;
  assign n16712 = ~n16659 & ~n16662;
  assign n16713 = ~n16711 & ~n16712;
  assign n16714 = ~n16662 & ~n16710;
  assign n16715 = n90 & n12938;
  assign n16716 = ~n53819 & n14236;
  assign n16717 = ~n53860 & n54667;
  assign n16718 = ~n53845 & n14210;
  assign n16719 = ~n16717 & ~n16718;
  assign n16720 = ~n16716 & ~n16717;
  assign n16721 = ~n16718 & n16720;
  assign n16722 = ~n16716 & n16719;
  assign n16723 = ~n16715 & n54971;
  assign n16724 = pi23  & ~n16723;
  assign n16725 = ~n16723 & ~n16724;
  assign n16726 = ~pi23  & ~n16723;
  assign n16727 = pi23  & ~n16724;
  assign n16728 = pi23  & n16723;
  assign n16729 = ~n54972 & ~n54973;
  assign n16730 = ~n16336 & n54954;
  assign n16731 = ~n16614 & ~n16730;
  assign n16732 = ~n16729 & n16731;
  assign n16733 = n16729 & ~n16731;
  assign n16734 = ~n16729 & ~n16732;
  assign n16735 = ~n16729 & ~n16731;
  assign n16736 = n16731 & ~n16732;
  assign n16737 = n16729 & n16731;
  assign n16738 = ~n54974 & ~n54975;
  assign n16739 = ~n16732 & ~n16733;
  assign n16740 = n16608 & ~n16610;
  assign n16741 = n16610 & ~n16611;
  assign n16742 = ~n16608 & ~n16611;
  assign n16743 = ~n16741 & ~n16742;
  assign n16744 = ~n16611 & ~n16740;
  assign n16745 = n11279 & n15219;
  assign n16746 = ~n54050 & n11267;
  assign n16747 = ~n54034 & n12584;
  assign n16748 = ~n54073 & n54410;
  assign n16749 = ~n16747 & ~n16748;
  assign n16750 = ~n16746 & ~n16748;
  assign n16751 = ~n16747 & n16750;
  assign n16752 = ~n16746 & n16749;
  assign n16753 = ~n16745 & n54978;
  assign n16754 = pi29  & ~n16753;
  assign n16755 = ~n16753 & ~n16754;
  assign n16756 = ~pi29  & ~n16753;
  assign n16757 = pi29  & ~n16754;
  assign n16758 = pi29  & n16753;
  assign n16759 = ~n54979 & ~n54980;
  assign n16760 = n16556 & ~n16558;
  assign n16761 = ~n16556 & ~n16559;
  assign n16762 = n16558 & ~n16559;
  assign n16763 = ~n16761 & ~n16762;
  assign n16764 = ~n16559 & ~n16760;
  assign n16765 = ~n16759 & ~n54981;
  assign n16766 = ~n16439 & n54943;
  assign n16767 = ~n54943 & ~n54944;
  assign n16768 = ~n16438 & n16540;
  assign n16769 = ~n16767 & ~n16768;
  assign n16770 = ~n54944 & ~n16766;
  assign n16771 = n10450 & ~n10452;
  assign n16772 = ~n10453 & ~n16771;
  assign n16773 = n1576 & n16772;
  assign n16774 = ~n54154 & n54403;
  assign n16775 = ~n54119 & n11215;
  assign n16776 = ~n54132 & n10564;
  assign n16777 = ~n16775 & ~n16776;
  assign n16778 = ~n16774 & ~n16776;
  assign n16779 = ~n16775 & n16778;
  assign n16780 = ~n16774 & n16777;
  assign n16781 = ~n16773 & ~n16774;
  assign n16782 = ~n16776 & n16781;
  assign n16783 = ~n16775 & n16782;
  assign n16784 = ~n16773 & n54983;
  assign n16785 = ~n54982 & ~n54984;
  assign n16786 = n16531 & ~n16533;
  assign n16787 = ~n16531 & ~n16534;
  assign n16788 = n16533 & ~n16534;
  assign n16789 = ~n16787 & ~n16788;
  assign n16790 = ~n16534 & ~n16786;
  assign n16791 = ~n503 & ~n1191;
  assign n16792 = ~n503 & ~n1703;
  assign n16793 = ~n1191 & n16792;
  assign n16794 = ~n1703 & n16791;
  assign n16795 = n3073 & n8453;
  assign n16796 = ~n1191 & n8453;
  assign n16797 = ~n1703 & n16796;
  assign n16798 = ~n172 & n16797;
  assign n16799 = ~n503 & n16798;
  assign n16800 = ~n498 & n16799;
  assign n16801 = ~n498 & ~n1703;
  assign n16802 = ~n1191 & n16801;
  assign n16803 = ~n172 & ~n503;
  assign n16804 = n8453 & n16803;
  assign n16805 = n16802 & n16804;
  assign n16806 = n54986 & n16795;
  assign n16807 = n2161 & n10901;
  assign n16808 = n13737 & n16807;
  assign n16809 = n53955 & n16808;
  assign n16810 = n54987 & n16809;
  assign n16811 = ~n464 & ~n832;
  assign n16812 = ~n832 & ~n1881;
  assign n16813 = ~n464 & n16812;
  assign n16814 = ~n464 & ~n1881;
  assign n16815 = ~n832 & n16814;
  assign n16816 = ~n1881 & n16811;
  assign n16817 = n1346 & n2691;
  assign n16818 = n3261 & n10300;
  assign n16819 = n1346 & n3261;
  assign n16820 = n2691 & n10300;
  assign n16821 = n16819 & n16820;
  assign n16822 = n16817 & n16818;
  assign n16823 = n1346 & n10300;
  assign n16824 = n2691 & n16823;
  assign n16825 = ~n464 & n16824;
  assign n16826 = ~n832 & n16825;
  assign n16827 = n3261 & n16826;
  assign n16828 = ~n1881 & n16827;
  assign n16829 = n54988 & n54989;
  assign n16830 = ~n448 & ~n771;
  assign n16831 = n1708 & n16830;
  assign n16832 = n1675 & n16831;
  assign n16833 = n54782 & n54795;
  assign n16834 = n16832 & n16833;
  assign n16835 = n54990 & n16834;
  assign n16836 = n1708 & n2161;
  assign n16837 = n13737 & n16836;
  assign n16838 = n53955 & n16837;
  assign n16839 = n54987 & n16838;
  assign n16840 = n10901 & n16830;
  assign n16841 = n1675 & n16840;
  assign n16842 = n16833 & n16841;
  assign n16843 = n54990 & n16842;
  assign n16844 = n16839 & n16843;
  assign n16845 = n1708 & n13737;
  assign n16846 = n10901 & n16845;
  assign n16847 = n53955 & n16846;
  assign n16848 = n54987 & n16847;
  assign n16849 = n2161 & n16830;
  assign n16850 = n1675 & n16849;
  assign n16851 = n16833 & n16850;
  assign n16852 = n54990 & n16851;
  assign n16853 = n16848 & n16852;
  assign n16854 = n16810 & n16835;
  assign n16855 = n53485 & n54991;
  assign n16856 = n54172 & n54247;
  assign n16857 = n13737 & n54795;
  assign n16858 = n54782 & n16857;
  assign n16859 = n53955 & n16858;
  assign n16860 = n54172 & n16859;
  assign n16861 = n53485 & n16860;
  assign n16862 = n54990 & n16861;
  assign n16863 = n54247 & n16862;
  assign n16864 = n54987 & n16863;
  assign n16865 = n1675 & n16864;
  assign n16866 = n10901 & n16865;
  assign n16867 = n1708 & n16866;
  assign n16868 = ~n833 & n16867;
  assign n16869 = ~n342 & n16868;
  assign n16870 = ~n771 & n16869;
  assign n16871 = ~n448 & n16870;
  assign n16872 = n16855 & n16856;
  assign n16873 = pi2  & ~n54992;
  assign n16874 = ~n751 & ~n1644;
  assign n16875 = n6614 & n14520;
  assign n16876 = n16874 & n16875;
  assign n16877 = n53785 & n16876;
  assign n16878 = n1708 & n4892;
  assign n16879 = n4892 & n11428;
  assign n16880 = n1708 & n16879;
  assign n16881 = n11428 & n16878;
  assign n16882 = n54619 & n54993;
  assign n16883 = n16877 & n16882;
  assign n16884 = ~n219 & ~n590;
  assign n16885 = ~n361 & ~n911;
  assign n16886 = ~n219 & ~n361;
  assign n16887 = ~n590 & ~n911;
  assign n16888 = n16886 & n16887;
  assign n16889 = ~n361 & ~n590;
  assign n16890 = ~n219 & ~n911;
  assign n16891 = n16889 & n16890;
  assign n16892 = n16884 & n16885;
  assign n16893 = n500 & n1659;
  assign n16894 = n54994 & n16893;
  assign n16895 = n3371 & n12821;
  assign n16896 = n16894 & n16895;
  assign n16897 = n54381 & n16896;
  assign n16898 = n5021 & n6614;
  assign n16899 = n14520 & n16898;
  assign n16900 = n53785 & n16899;
  assign n16901 = n16882 & n16900;
  assign n16902 = n4530 & n16874;
  assign n16903 = n16893 & n16902;
  assign n16904 = n3371 & n54994;
  assign n16905 = n16903 & n16904;
  assign n16906 = n54381 & n16905;
  assign n16907 = n16901 & n16906;
  assign n16908 = n16883 & n16897;
  assign n16909 = n53818 & n54995;
  assign n16910 = n14520 & n54993;
  assign n16911 = n3371 & n16910;
  assign n16912 = n53818 & n16911;
  assign n16913 = n54381 & n16912;
  assign n16914 = n54290 & n16913;
  assign n16915 = n53785 & n16914;
  assign n16916 = n54619 & n16915;
  assign n16917 = n500 & n16916;
  assign n16918 = n1659 & n16917;
  assign n16919 = n4530 & n16918;
  assign n16920 = n5021 & n16919;
  assign n16921 = n6614 & n16920;
  assign n16922 = ~n219 & n16921;
  assign n16923 = ~n911 & n16922;
  assign n16924 = ~n1644 & n16923;
  assign n16925 = ~n361 & n16924;
  assign n16926 = ~n751 & n16925;
  assign n16927 = ~n590 & n16926;
  assign n16928 = n54290 & n16909;
  assign n16929 = pi2  & ~n54996;
  assign n16930 = n1675 & n54280;
  assign n16931 = n54794 & n16930;
  assign n16932 = n2326 & n3671;
  assign n16933 = n6577 & n11043;
  assign n16934 = n16932 & n16933;
  assign n16935 = ~n310 & ~n344;
  assign n16936 = ~n1061 & n16935;
  assign n16937 = ~n221 & ~n296;
  assign n16938 = n1659 & n16937;
  assign n16939 = ~n221 & ~n310;
  assign n16940 = ~n1061 & n16939;
  assign n16941 = ~n296 & ~n344;
  assign n16942 = n1659 & n16941;
  assign n16943 = n16940 & n16942;
  assign n16944 = n16936 & n16938;
  assign n16945 = n1659 & n3671;
  assign n16946 = n2326 & n6577;
  assign n16947 = n16945 & n16946;
  assign n16948 = ~n221 & ~n1061;
  assign n16949 = ~n296 & n16948;
  assign n16950 = n11043 & n16935;
  assign n16951 = n16949 & n16950;
  assign n16952 = n16947 & n16951;
  assign n16953 = n1659 & n6577;
  assign n16954 = n3671 & n11043;
  assign n16955 = n16953 & n16954;
  assign n16956 = ~n296 & n16939;
  assign n16957 = ~n344 & ~n1061;
  assign n16958 = n2326 & n16957;
  assign n16959 = n16956 & n16958;
  assign n16960 = n16955 & n16959;
  assign n16961 = n16934 & n54997;
  assign n16962 = n54801 & n54998;
  assign n16963 = n54280 & n54794;
  assign n16964 = n6577 & n16963;
  assign n16965 = n11043 & n16964;
  assign n16966 = n54801 & n16965;
  assign n16967 = n3671 & n16966;
  assign n16968 = n1675 & n16967;
  assign n16969 = n1659 & n16968;
  assign n16970 = n2326 & n16969;
  assign n16971 = ~n296 & n16970;
  assign n16972 = ~n1061 & n16971;
  assign n16973 = ~n310 & n16972;
  assign n16974 = ~n221 & n16973;
  assign n16975 = ~n344 & n16974;
  assign n16976 = n16931 & n16962;
  assign n16977 = ~n419 & ~n776;
  assign n16978 = n4223 & n16977;
  assign n16979 = n8679 & n10183;
  assign n16980 = n16978 & n16979;
  assign n16981 = n54396 & n16980;
  assign n16982 = ~n402 & ~n823;
  assign n16983 = ~n881 & n16982;
  assign n16984 = ~n651 & ~n849;
  assign n16985 = n2367 & n16984;
  assign n16986 = ~n881 & n2367;
  assign n16987 = ~n402 & n16986;
  assign n16988 = ~n823 & n16987;
  assign n16989 = ~n849 & n16988;
  assign n16990 = ~n651 & n16989;
  assign n16991 = ~n402 & ~n651;
  assign n16992 = ~n849 & n16991;
  assign n16993 = ~n823 & ~n881;
  assign n16994 = n2367 & n16993;
  assign n16995 = n16992 & n16994;
  assign n16996 = ~n823 & n16991;
  assign n16997 = ~n849 & ~n881;
  assign n16998 = n2367 & n16997;
  assign n16999 = n16996 & n16998;
  assign n17000 = n16983 & n16985;
  assign n17001 = n10901 & n13530;
  assign n17002 = n14539 & n17001;
  assign n17003 = n55000 & n17002;
  assign n17004 = n4223 & n8679;
  assign n17005 = n10901 & n16977;
  assign n17006 = n17004 & n17005;
  assign n17007 = n54396 & n17006;
  assign n17008 = n10183 & n13530;
  assign n17009 = n14539 & n17008;
  assign n17010 = n55000 & n17009;
  assign n17011 = n17007 & n17010;
  assign n17012 = n14539 & n16977;
  assign n17013 = n17004 & n17012;
  assign n17014 = n54396 & n17013;
  assign n17015 = n10901 & n17008;
  assign n17016 = n55000 & n17015;
  assign n17017 = n17014 & n17016;
  assign n17018 = n16981 & n17003;
  assign n17019 = n54316 & n54386;
  assign n17020 = n55001 & n17019;
  assign n17021 = n54999 & n17020;
  assign n17022 = n54396 & n13530;
  assign n17023 = n8679 & n17022;
  assign n17024 = n10183 & n17023;
  assign n17025 = n55000 & n17024;
  assign n17026 = n54316 & n17025;
  assign n17027 = n54999 & n17026;
  assign n17028 = n54386 & n17027;
  assign n17029 = n4223 & n17028;
  assign n17030 = n53986 & n17029;
  assign n17031 = n10901 & n17030;
  assign n17032 = ~n419 & n17031;
  assign n17033 = ~n353 & n17032;
  assign n17034 = ~n776 & n17033;
  assign n17035 = ~n751 & n17034;
  assign n17036 = n53986 & n17021;
  assign n17037 = pi2  & ~n55002;
  assign n17038 = ~pi2  & n55002;
  assign n17039 = ~n17037 & ~n17038;
  assign n17040 = n10430 & ~n10432;
  assign n17041 = ~n10433 & ~n17040;
  assign n17042 = n1576 & n17041;
  assign n17043 = ~n54212 & n10564;
  assign n17044 = ~n54194 & n11215;
  assign n17045 = ~n54240 & n54403;
  assign n17046 = ~n17044 & ~n17045;
  assign n17047 = ~n17043 & ~n17045;
  assign n17048 = ~n17044 & n17047;
  assign n17049 = ~n17043 & n17046;
  assign n17050 = ~n17042 & n55003;
  assign n17051 = ~n17037 & ~n17050;
  assign n17052 = ~n17038 & n17051;
  assign n17053 = n17039 & ~n17050;
  assign n17054 = ~n17037 & ~n55004;
  assign n17055 = ~pi2  & n54996;
  assign n17056 = ~n16929 & ~n17055;
  assign n17057 = ~n16929 & ~n17054;
  assign n17058 = ~n17055 & n17057;
  assign n17059 = ~n17054 & n17056;
  assign n17060 = ~n16929 & ~n55005;
  assign n17061 = ~pi2  & n54992;
  assign n17062 = ~n16873 & ~n17061;
  assign n17063 = ~n16873 & ~n17060;
  assign n17064 = ~n17061 & n17063;
  assign n17065 = ~n17060 & n17062;
  assign n17066 = ~n16873 & ~n55006;
  assign n17067 = pi5  & n54941;
  assign n17068 = ~n16517 & ~n17067;
  assign n17069 = ~n17066 & n17068;
  assign n17070 = n17066 & ~n17068;
  assign n17071 = n10442 & ~n10444;
  assign n17072 = ~n10445 & ~n17071;
  assign n17073 = n1576 & n17072;
  assign n17074 = ~n54154 & n11215;
  assign n17075 = ~n54183 & n54403;
  assign n17076 = ~n54163 & n10564;
  assign n17077 = ~n17075 & ~n17076;
  assign n17078 = ~n17074 & n17077;
  assign n17079 = ~n17073 & n17078;
  assign n17080 = ~n17070 & ~n17079;
  assign n17081 = ~n17069 & ~n17070;
  assign n17082 = ~n17079 & n17081;
  assign n17083 = ~n17069 & ~n17082;
  assign n17084 = ~n17069 & ~n17080;
  assign n17085 = ~n54985 & ~n55007;
  assign n17086 = n54985 & n55007;
  assign n17087 = ~n17085 & ~n17086;
  assign n17088 = n11279 & n15779;
  assign n17089 = ~n54098 & n11267;
  assign n17090 = ~n54119 & n54410;
  assign n17091 = ~n54073 & n12584;
  assign n17092 = ~n17090 & ~n17091;
  assign n17093 = ~n17089 & ~n17090;
  assign n17094 = ~n17091 & n17093;
  assign n17095 = ~n17089 & ~n17091;
  assign n17096 = ~n17090 & n17095;
  assign n17097 = ~n17089 & n17092;
  assign n17098 = ~n11279 & n55008;
  assign n17099 = ~n15779 & n55008;
  assign n17100 = ~n17098 & ~n17099;
  assign n17101 = ~n17088 & n55008;
  assign n17102 = pi29  & ~n55009;
  assign n17103 = ~pi29  & n55009;
  assign n17104 = ~n17102 & ~n17103;
  assign n17105 = n17087 & ~n17104;
  assign n17106 = ~n17085 & ~n17105;
  assign n17107 = n54982 & n54984;
  assign n17108 = ~n54982 & ~n16785;
  assign n17109 = ~n54982 & n54984;
  assign n17110 = ~n54984 & ~n16785;
  assign n17111 = n54982 & ~n54984;
  assign n17112 = ~n55010 & ~n55011;
  assign n17113 = ~n16785 & ~n17107;
  assign n17114 = ~n17106 & ~n55012;
  assign n17115 = ~n16785 & ~n17114;
  assign n17116 = n16759 & n54981;
  assign n17117 = ~n16759 & ~n16765;
  assign n17118 = ~n16759 & n54981;
  assign n17119 = ~n54981 & ~n16765;
  assign n17120 = n16759 & ~n54981;
  assign n17121 = ~n55013 & ~n55014;
  assign n17122 = ~n16765 & ~n17116;
  assign n17123 = ~n17115 & ~n55015;
  assign n17124 = ~n16765 & ~n17123;
  assign n17125 = ~n16569 & n16584;
  assign n17126 = ~n16585 & ~n17125;
  assign n17127 = ~n17124 & n17126;
  assign n17128 = n17124 & ~n17126;
  assign n17129 = n123 & n14020;
  assign n17130 = n127 & ~n53962;
  assign n17131 = n53444 & ~n53970;
  assign n17132 = n128 & ~n53930;
  assign n17133 = ~n17131 & ~n17132;
  assign n17134 = ~n17130 & ~n17131;
  assign n17135 = ~n17132 & n17134;
  assign n17136 = ~n17130 & n17133;
  assign n17137 = ~n17129 & n55016;
  assign n17138 = pi26  & ~n17137;
  assign n17139 = pi26  & ~n17138;
  assign n17140 = pi26  & n17137;
  assign n17141 = ~n17137 & ~n17138;
  assign n17142 = ~pi26  & ~n17137;
  assign n17143 = ~n55017 & ~n55018;
  assign n17144 = ~n17128 & ~n17143;
  assign n17145 = ~n17127 & ~n17128;
  assign n17146 = ~n17143 & n17145;
  assign n17147 = ~n17127 & ~n17146;
  assign n17148 = ~n17127 & ~n17144;
  assign n17149 = ~n54977 & ~n55019;
  assign n17150 = n54977 & n55019;
  assign n17151 = n90 & n12918;
  assign n17152 = ~n53860 & n14210;
  assign n17153 = ~n53888 & n54667;
  assign n17154 = ~n53845 & n14236;
  assign n17155 = ~n17153 & ~n17154;
  assign n17156 = ~n17152 & ~n17153;
  assign n17157 = ~n17154 & n17156;
  assign n17158 = ~n17152 & n17155;
  assign n17159 = ~n17151 & n55020;
  assign n17160 = pi23  & ~n17159;
  assign n17161 = pi23  & ~n17160;
  assign n17162 = pi23  & n17159;
  assign n17163 = ~n17159 & ~n17160;
  assign n17164 = ~pi23  & ~n17159;
  assign n17165 = ~n55021 & ~n55022;
  assign n17166 = ~n17150 & ~n17165;
  assign n17167 = ~n17149 & ~n17150;
  assign n17168 = ~n17165 & n17167;
  assign n17169 = ~n17149 & ~n17168;
  assign n17170 = ~n17149 & ~n17166;
  assign n17171 = ~n54976 & ~n55023;
  assign n17172 = ~n16732 & ~n17171;
  assign n17173 = n16639 & ~n16640;
  assign n17174 = n16637 & n16639;
  assign n17175 = ~n16637 & ~n16640;
  assign n17176 = ~n16637 & ~n16639;
  assign n17177 = n16637 & ~n16639;
  assign n17178 = ~n16640 & ~n17177;
  assign n17179 = ~n55024 & ~n55025;
  assign n17180 = ~n17172 & n55026;
  assign n17181 = n17172 & ~n55026;
  assign n17182 = n11889 & n14413;
  assign n17183 = ~n53712 & n15921;
  assign n17184 = ~n53774 & n54719;
  assign n17185 = ~n53741 & n15901;
  assign n17186 = ~n17184 & ~n17185;
  assign n17187 = ~n17183 & ~n17184;
  assign n17188 = ~n17185 & n17187;
  assign n17189 = ~n17183 & n17186;
  assign n17190 = ~n17182 & n55027;
  assign n17191 = pi20  & ~n17190;
  assign n17192 = pi20  & ~n17191;
  assign n17193 = pi20  & n17190;
  assign n17194 = ~n17190 & ~n17191;
  assign n17195 = ~pi20  & ~n17190;
  assign n17196 = ~n55028 & ~n55029;
  assign n17197 = ~n17181 & ~n17196;
  assign n17198 = ~n17180 & ~n17181;
  assign n17199 = ~n17196 & n17198;
  assign n17200 = ~n17180 & ~n17199;
  assign n17201 = ~n17180 & ~n17197;
  assign n17202 = ~n54970 & ~n55030;
  assign n17203 = n54970 & n55030;
  assign n17204 = n11286 & n16079;
  assign n17205 = ~n53650 & n16676;
  assign n17206 = ~n53657 & n54886;
  assign n17207 = ~n53634 & n16696;
  assign n17208 = ~n17206 & ~n17207;
  assign n17209 = ~n17205 & ~n17206;
  assign n17210 = ~n17207 & n17209;
  assign n17211 = ~n17205 & n17208;
  assign n17212 = ~n17204 & n55031;
  assign n17213 = pi17  & ~n17212;
  assign n17214 = pi17  & ~n17213;
  assign n17215 = pi17  & n17212;
  assign n17216 = ~n17212 & ~n17213;
  assign n17217 = ~pi17  & ~n17212;
  assign n17218 = ~n55032 & ~n55033;
  assign n17219 = ~n17203 & ~n17218;
  assign n17220 = ~n17202 & ~n17203;
  assign n17221 = ~n17218 & n17220;
  assign n17222 = ~n17202 & ~n17221;
  assign n17223 = ~n17202 & ~n17219;
  assign n17224 = ~n16709 & ~n55034;
  assign n17225 = n16709 & n55034;
  assign n17226 = ~n17224 & ~n17225;
  assign n17227 = ~n16308 & n54963;
  assign n17228 = ~n16665 & ~n17227;
  assign n17229 = n17226 & n17228;
  assign n17230 = ~n17224 & ~n17229;
  assign n17231 = n16687 & ~n16688;
  assign n17232 = n16685 & n16687;
  assign n17233 = ~n16685 & ~n16688;
  assign n17234 = ~n16685 & ~n16687;
  assign n17235 = n16685 & ~n16687;
  assign n17236 = ~n16688 & ~n17235;
  assign n17237 = ~n55035 & ~n55036;
  assign n17238 = ~n17230 & n55037;
  assign n17239 = n17230 & ~n55037;
  assign n17240 = ~n17238 & ~n17239;
  assign n17241 = ~n17226 & ~n17228;
  assign n17242 = ~n17229 & ~n17241;
  assign n17243 = pi12  & ~pi13 ;
  assign n17244 = ~pi12  & pi13 ;
  assign n17245 = ~pi12  & ~pi13 ;
  assign n17246 = pi12  & pi13 ;
  assign n17247 = ~n17245 & ~n17246;
  assign n17248 = ~n17243 & ~n17244;
  assign n17249 = pi11  & ~pi12 ;
  assign n17250 = ~pi11  & pi12 ;
  assign n17251 = ~pi11  & ~pi12 ;
  assign n17252 = pi11  & pi12 ;
  assign n17253 = ~n17251 & ~n17252;
  assign n17254 = ~n17249 & ~n17250;
  assign n17255 = ~n55038 & ~n55039;
  assign n17256 = pi13  & ~pi14 ;
  assign n17257 = ~pi13  & pi14 ;
  assign n17258 = ~pi13  & ~pi14 ;
  assign n17259 = pi13  & pi14 ;
  assign n17260 = ~n17258 & ~n17259;
  assign n17261 = ~n17256 & ~n17257;
  assign n17262 = ~n55039 & n55040;
  assign n17263 = ~n55038 & n17262;
  assign n17264 = n17255 & n55040;
  assign n17265 = n55039 & n55040;
  assign n17266 = ~n10547 & n17265;
  assign n17267 = ~n55041 & ~n17266;
  assign n17268 = ~n2325 & n55041;
  assign n17269 = ~n17265 & ~n17268;
  assign n17270 = ~n10551 & ~n17268;
  assign n17271 = ~n17269 & ~n17270;
  assign n17272 = ~n2325 & ~n17267;
  assign n17273 = pi14  & ~n55042;
  assign n17274 = ~pi14  & n55042;
  assign n17275 = ~n17273 & ~n17274;
  assign n17276 = n54976 & n55023;
  assign n17277 = ~n17171 & ~n17276;
  assign n17278 = n11913 & n14413;
  assign n17279 = ~n53774 & n15901;
  assign n17280 = ~n53799 & n54719;
  assign n17281 = ~n53741 & n15921;
  assign n17282 = ~n17280 & ~n17281;
  assign n17283 = ~n17279 & ~n17280;
  assign n17284 = ~n17281 & n17283;
  assign n17285 = ~n17279 & n17282;
  assign n17286 = ~n14413 & n55043;
  assign n17287 = ~n11913 & n55043;
  assign n17288 = ~n17286 & ~n17287;
  assign n17289 = ~n17278 & n55043;
  assign n17290 = pi20  & ~n55044;
  assign n17291 = ~pi20  & n55044;
  assign n17292 = ~n17290 & ~n17291;
  assign n17293 = n17277 & ~n17292;
  assign n17294 = ~n17277 & n17292;
  assign n17295 = ~n17293 & ~n17294;
  assign n17296 = n17165 & ~n17167;
  assign n17297 = n17167 & ~n17168;
  assign n17298 = ~n17165 & ~n17168;
  assign n17299 = ~n17297 & ~n17298;
  assign n17300 = ~n17168 & ~n17296;
  assign n17301 = n17115 & n55015;
  assign n17302 = ~n17123 & ~n17301;
  assign n17303 = n123 & n14708;
  assign n17304 = n53444 & ~n54005;
  assign n17305 = n127 & ~n53970;
  assign n17306 = n128 & ~n53962;
  assign n17307 = ~n17305 & ~n17306;
  assign n17308 = ~n17304 & ~n17305;
  assign n17309 = ~n17306 & n17308;
  assign n17310 = ~n17304 & n17307;
  assign n17311 = ~n123 & n55046;
  assign n17312 = ~n14708 & n55046;
  assign n17313 = ~n17311 & ~n17312;
  assign n17314 = ~n17303 & n55046;
  assign n17315 = pi26  & ~n55047;
  assign n17316 = ~pi26  & n55047;
  assign n17317 = ~n17315 & ~n17316;
  assign n17318 = n17302 & ~n17317;
  assign n17319 = ~n17302 & n17317;
  assign n17320 = ~n17318 & ~n17319;
  assign n17321 = n11279 & n16138;
  assign n17322 = ~n54098 & n54410;
  assign n17323 = ~n54050 & n12584;
  assign n17324 = ~n54073 & n11267;
  assign n17325 = ~n17323 & ~n17324;
  assign n17326 = ~n17322 & ~n17324;
  assign n17327 = ~n17323 & n17326;
  assign n17328 = ~n17322 & n17325;
  assign n17329 = ~n11279 & n55048;
  assign n17330 = ~n16138 & n55048;
  assign n17331 = ~n17329 & ~n17330;
  assign n17332 = ~n17321 & n55048;
  assign n17333 = pi29  & ~n55049;
  assign n17334 = ~pi29  & n55049;
  assign n17335 = ~n17333 & ~n17334;
  assign n17336 = n17106 & n55012;
  assign n17337 = ~n17106 & ~n17114;
  assign n17338 = ~n55012 & ~n17114;
  assign n17339 = ~n17337 & ~n17338;
  assign n17340 = ~n17114 & ~n17336;
  assign n17341 = ~n17335 & ~n55050;
  assign n17342 = n17335 & n55050;
  assign n17343 = n123 & n14688;
  assign n17344 = n127 & ~n54005;
  assign n17345 = n53444 & ~n54034;
  assign n17346 = n128 & ~n53970;
  assign n17347 = ~n17345 & ~n17346;
  assign n17348 = ~n17344 & ~n17345;
  assign n17349 = ~n17346 & n17348;
  assign n17350 = ~n17344 & n17347;
  assign n17351 = ~n17343 & n55051;
  assign n17352 = pi26  & ~n17351;
  assign n17353 = pi26  & ~n17352;
  assign n17354 = pi26  & n17351;
  assign n17355 = ~n17351 & ~n17352;
  assign n17356 = ~pi26  & ~n17351;
  assign n17357 = ~n55052 & ~n55053;
  assign n17358 = ~n17342 & ~n17357;
  assign n17359 = ~n17341 & ~n17342;
  assign n17360 = ~n17357 & n17359;
  assign n17361 = ~n17341 & ~n17360;
  assign n17362 = ~n17341 & ~n17358;
  assign n17363 = n17320 & ~n55054;
  assign n17364 = ~n17318 & ~n17363;
  assign n17365 = n17143 & ~n17145;
  assign n17366 = n17145 & ~n17146;
  assign n17367 = ~n17143 & ~n17146;
  assign n17368 = ~n17366 & ~n17367;
  assign n17369 = ~n17146 & ~n17365;
  assign n17370 = ~n17364 & ~n55055;
  assign n17371 = n17364 & n55055;
  assign n17372 = n90 & n13336;
  assign n17373 = ~n53888 & n14210;
  assign n17374 = ~n53907 & n54667;
  assign n17375 = ~n53860 & n14236;
  assign n17376 = ~n17374 & ~n17375;
  assign n17377 = ~n17373 & ~n17374;
  assign n17378 = ~n17375 & n17377;
  assign n17379 = ~n17373 & n17376;
  assign n17380 = ~n17372 & n55056;
  assign n17381 = pi23  & ~n17380;
  assign n17382 = pi23  & ~n17381;
  assign n17383 = pi23  & n17380;
  assign n17384 = ~n17380 & ~n17381;
  assign n17385 = ~pi23  & ~n17380;
  assign n17386 = ~n55057 & ~n55058;
  assign n17387 = ~n17371 & ~n17386;
  assign n17388 = ~n17370 & ~n17371;
  assign n17389 = ~n17386 & n17388;
  assign n17390 = ~n17370 & ~n17389;
  assign n17391 = ~n17370 & ~n17387;
  assign n17392 = ~n55045 & ~n55059;
  assign n17393 = n55045 & n55059;
  assign n17394 = n12690 & n14413;
  assign n17395 = ~n53774 & n15921;
  assign n17396 = ~n53819 & n54719;
  assign n17397 = ~n53799 & n15901;
  assign n17398 = ~n17396 & ~n17397;
  assign n17399 = ~n17395 & ~n17396;
  assign n17400 = ~n17397 & n17399;
  assign n17401 = ~n17395 & n17398;
  assign n17402 = ~n17394 & n55060;
  assign n17403 = pi20  & ~n17402;
  assign n17404 = pi20  & ~n17403;
  assign n17405 = pi20  & n17402;
  assign n17406 = ~n17402 & ~n17403;
  assign n17407 = ~pi20  & ~n17402;
  assign n17408 = ~n55061 & ~n55062;
  assign n17409 = ~n17393 & ~n17408;
  assign n17410 = ~n17392 & ~n17393;
  assign n17411 = ~n17408 & n17410;
  assign n17412 = ~n17392 & ~n17411;
  assign n17413 = ~n17392 & ~n17409;
  assign n17414 = n17295 & ~n55063;
  assign n17415 = ~n17293 & ~n17414;
  assign n17416 = n17196 & ~n17198;
  assign n17417 = n17198 & ~n17199;
  assign n17418 = ~n17196 & ~n17199;
  assign n17419 = ~n17417 & ~n17418;
  assign n17420 = ~n17199 & ~n17416;
  assign n17421 = ~n17415 & ~n55064;
  assign n17422 = n17415 & n55064;
  assign n17423 = n11213 & n16079;
  assign n17424 = ~n53650 & n16696;
  assign n17425 = ~n53685 & n54886;
  assign n17426 = ~n53657 & n16676;
  assign n17427 = ~n17425 & ~n17426;
  assign n17428 = ~n17424 & n17427;
  assign n17429 = ~n17423 & n17428;
  assign n17430 = pi17  & ~n17429;
  assign n17431 = pi17  & ~n17430;
  assign n17432 = pi17  & n17429;
  assign n17433 = ~n17429 & ~n17430;
  assign n17434 = ~pi17  & ~n17429;
  assign n17435 = ~n55065 & ~n55066;
  assign n17436 = ~n17422 & ~n17435;
  assign n17437 = ~n17421 & ~n17422;
  assign n17438 = ~n17435 & n17437;
  assign n17439 = ~n17421 & ~n17438;
  assign n17440 = ~n17421 & ~n17436;
  assign n17441 = ~n17275 & ~n55067;
  assign n17442 = n17275 & n55067;
  assign n17443 = n17218 & ~n17220;
  assign n17444 = n17220 & ~n17221;
  assign n17445 = ~n17218 & ~n17221;
  assign n17446 = ~n17444 & ~n17445;
  assign n17447 = ~n17221 & ~n17443;
  assign n17448 = ~n17442 & ~n55068;
  assign n17449 = ~n17441 & ~n17442;
  assign n17450 = ~n55068 & n17449;
  assign n17451 = ~n17441 & ~n17450;
  assign n17452 = ~n17441 & ~n17448;
  assign n17453 = n17242 & ~n55069;
  assign n17454 = ~n17242 & n55069;
  assign n17455 = ~n17453 & ~n17454;
  assign n17456 = n11380 & n16079;
  assign n17457 = ~n53685 & n16676;
  assign n17458 = ~n53657 & n16696;
  assign n17459 = ~n53712 & n54886;
  assign n17460 = ~n17458 & ~n17459;
  assign n17461 = ~n17457 & ~n17459;
  assign n17462 = ~n17458 & n17461;
  assign n17463 = ~n17457 & n17460;
  assign n17464 = ~n17456 & n55070;
  assign n17465 = pi17  & ~n17464;
  assign n17466 = ~n17464 & ~n17465;
  assign n17467 = ~pi17  & ~n17464;
  assign n17468 = pi17  & ~n17465;
  assign n17469 = pi17  & n17464;
  assign n17470 = ~n55071 & ~n55072;
  assign n17471 = ~n17295 & n55063;
  assign n17472 = ~n17414 & ~n17471;
  assign n17473 = ~n17470 & n17472;
  assign n17474 = n17470 & ~n17472;
  assign n17475 = ~n17470 & ~n17473;
  assign n17476 = ~n17470 & ~n17472;
  assign n17477 = n17472 & ~n17473;
  assign n17478 = n17470 & n17472;
  assign n17479 = ~n55073 & ~n55074;
  assign n17480 = ~n17473 & ~n17474;
  assign n17481 = n17408 & ~n17410;
  assign n17482 = n17410 & ~n17411;
  assign n17483 = ~n17408 & ~n17411;
  assign n17484 = ~n17482 & ~n17483;
  assign n17485 = ~n17411 & ~n17481;
  assign n17486 = n90 & n13360;
  assign n17487 = ~n53907 & n14210;
  assign n17488 = ~n53930 & n54667;
  assign n17489 = ~n53888 & n14236;
  assign n17490 = ~n17488 & ~n17489;
  assign n17491 = ~n17487 & ~n17488;
  assign n17492 = ~n17489 & n17491;
  assign n17493 = ~n17487 & n17490;
  assign n17494 = ~n17486 & n55077;
  assign n17495 = pi23  & ~n17494;
  assign n17496 = ~n17494 & ~n17495;
  assign n17497 = ~pi23  & ~n17494;
  assign n17498 = pi23  & ~n17495;
  assign n17499 = pi23  & n17494;
  assign n17500 = ~n55078 & ~n55079;
  assign n17501 = ~n17320 & n55054;
  assign n17502 = ~n17363 & ~n17501;
  assign n17503 = ~n17500 & n17502;
  assign n17504 = n17500 & ~n17502;
  assign n17505 = ~n17500 & ~n17503;
  assign n17506 = ~n17500 & ~n17502;
  assign n17507 = n17502 & ~n17503;
  assign n17508 = n17500 & n17502;
  assign n17509 = ~n55080 & ~n55081;
  assign n17510 = ~n17503 & ~n17504;
  assign n17511 = n17357 & ~n17359;
  assign n17512 = n17359 & ~n17360;
  assign n17513 = ~n17357 & ~n17360;
  assign n17514 = ~n17512 & ~n17513;
  assign n17515 = ~n17360 & ~n17511;
  assign n17516 = ~n17087 & n17104;
  assign n17517 = ~n17105 & ~n17516;
  assign n17518 = n17060 & ~n17062;
  assign n17519 = ~n17060 & ~n55006;
  assign n17520 = ~n17061 & n17066;
  assign n17521 = ~n17519 & ~n17520;
  assign n17522 = ~n55006 & ~n17518;
  assign n17523 = n10438 & ~n10440;
  assign n17524 = ~n10441 & ~n17523;
  assign n17525 = n1576 & n17524;
  assign n17526 = ~n54194 & n54403;
  assign n17527 = ~n54183 & n10564;
  assign n17528 = ~n54163 & n11215;
  assign n17529 = ~n17527 & ~n17528;
  assign n17530 = ~n17526 & ~n17527;
  assign n17531 = ~n17528 & n17530;
  assign n17532 = ~n17526 & n17529;
  assign n17533 = ~n17525 & ~n17526;
  assign n17534 = ~n17527 & n17533;
  assign n17535 = ~n17528 & n17534;
  assign n17536 = ~n17525 & n55085;
  assign n17537 = ~n55084 & ~n55086;
  assign n17538 = n17054 & ~n17056;
  assign n17539 = ~n17054 & ~n55005;
  assign n17540 = ~n17055 & n17060;
  assign n17541 = ~n17539 & ~n17540;
  assign n17542 = ~n55005 & ~n17538;
  assign n17543 = n10434 & ~n10436;
  assign n17544 = ~n10437 & ~n17543;
  assign n17545 = n1576 & n17544;
  assign n17546 = ~n54212 & n54403;
  assign n17547 = ~n54183 & n11215;
  assign n17548 = ~n54194 & n10564;
  assign n17549 = ~n17547 & ~n17548;
  assign n17550 = ~n17546 & n17549;
  assign n17551 = ~n17545 & ~n17546;
  assign n17552 = ~n17548 & n17551;
  assign n17553 = ~n17547 & n17552;
  assign n17554 = ~n17545 & n17550;
  assign n17555 = ~n55087 & ~n55088;
  assign n17556 = ~n506 & ~n1881;
  assign n17557 = ~n506 & n2405;
  assign n17558 = ~n1881 & n17557;
  assign n17559 = n2405 & n17556;
  assign n17560 = n5387 & n54373;
  assign n17561 = n55089 & n17560;
  assign n17562 = ~n559 & ~n585;
  assign n17563 = ~n402 & n17562;
  assign n17564 = ~n559 & n3882;
  assign n17565 = ~n559 & n15314;
  assign n17566 = ~n402 & n17565;
  assign n17567 = ~n585 & n17566;
  assign n17568 = n15314 & n55090;
  assign n17569 = n5021 & n7307;
  assign n17570 = n7811 & n9622;
  assign n17571 = n17569 & n17570;
  assign n17572 = n3821 & n4893;
  assign n17573 = n53474 & n17572;
  assign n17574 = n17571 & n17573;
  assign n17575 = n55091 & n17574;
  assign n17576 = n53474 & n55089;
  assign n17577 = n53474 & n54373;
  assign n17578 = n55089 & n17577;
  assign n17579 = n54373 & n17576;
  assign n17580 = n4893 & n5021;
  assign n17581 = n3821 & n7307;
  assign n17582 = n17580 & n17581;
  assign n17583 = ~n444 & n9622;
  assign n17584 = n1659 & n7811;
  assign n17585 = n17583 & n17584;
  assign n17586 = ~n444 & n4893;
  assign n17587 = n1659 & n3821;
  assign n17588 = n5387 & n17572;
  assign n17589 = n17586 & n17587;
  assign n17590 = n17571 & n55093;
  assign n17591 = n17582 & n17585;
  assign n17592 = n55091 & n55094;
  assign n17593 = n55092 & n17592;
  assign n17594 = n17561 & n17575;
  assign n17595 = n54638 & n55095;
  assign n17596 = n1488 & n3014;
  assign n17597 = n1672 & n5378;
  assign n17598 = n3014 & n5378;
  assign n17599 = n1488 & n1672;
  assign n17600 = n17598 & n17599;
  assign n17601 = n17596 & n17597;
  assign n17602 = ~n1466 & ~n1644;
  assign n17603 = ~n902 & ~n1644;
  assign n17604 = ~n1466 & n17603;
  assign n17605 = ~n902 & n17602;
  assign n17606 = ~n112 & ~n275;
  assign n17607 = n309 & n17606;
  assign n17608 = n55097 & n17607;
  assign n17609 = n309 & n1488;
  assign n17610 = n17597 & n17609;
  assign n17611 = ~n275 & n17602;
  assign n17612 = ~n112 & ~n902;
  assign n17613 = n3014 & n17612;
  assign n17614 = n17611 & n17613;
  assign n17615 = n17610 & n17614;
  assign n17616 = n55096 & n17608;
  assign n17617 = n9766 & n13912;
  assign n17618 = n14520 & n17617;
  assign n17619 = n54621 & n17618;
  assign n17620 = ~n275 & n17612;
  assign n17621 = n9766 & n17602;
  assign n17622 = n17620 & n17621;
  assign n17623 = n55096 & n17622;
  assign n17624 = n309 & n13912;
  assign n17625 = n14520 & n17624;
  assign n17626 = n54621 & n17625;
  assign n17627 = n17623 & n17626;
  assign n17628 = n55098 & n17619;
  assign n17629 = n54114 & n17619;
  assign n17630 = n1488 & n17629;
  assign n17631 = n5378 & n17630;
  assign n17632 = n1672 & n17631;
  assign n17633 = n309 & n17632;
  assign n17634 = n3014 & n17633;
  assign n17635 = ~n902 & n17634;
  assign n17636 = ~n1466 & n17635;
  assign n17637 = ~n112 & n17636;
  assign n17638 = ~n275 & n17637;
  assign n17639 = ~n1644 & n17638;
  assign n17640 = n54114 & n55099;
  assign n17641 = n54643 & n55100;
  assign n17642 = n3821 & n54373;
  assign n17643 = n4893 & n17642;
  assign n17644 = n55089 & n17643;
  assign n17645 = n55091 & n17644;
  assign n17646 = n7307 & n17645;
  assign n17647 = n54643 & n17646;
  assign n17648 = n54638 & n17647;
  assign n17649 = n55100 & n17648;
  assign n17650 = n1659 & n17649;
  assign n17651 = n5021 & n17650;
  assign n17652 = n53474 & n17651;
  assign n17653 = ~n1125 & n17652;
  assign n17654 = ~n141 & n17653;
  assign n17655 = ~n441 & n17654;
  assign n17656 = ~n461 & n17655;
  assign n17657 = ~n444 & n17656;
  assign n17658 = n17595 & n17641;
  assign n17659 = n10426 & ~n10428;
  assign n17660 = ~n10429 & ~n17659;
  assign n17661 = n1576 & n17660;
  assign n17662 = ~n54254 & n54403;
  assign n17663 = ~n54212 & n11215;
  assign n17664 = ~n54240 & n10564;
  assign n17665 = ~n17663 & ~n17664;
  assign n17666 = ~n17662 & ~n17664;
  assign n17667 = ~n17663 & n17666;
  assign n17668 = ~n17662 & n17665;
  assign n17669 = ~n17661 & ~n17662;
  assign n17670 = ~n17664 & n17669;
  assign n17671 = ~n17663 & n17670;
  assign n17672 = ~n17661 & n55102;
  assign n17673 = ~n55101 & ~n55103;
  assign n17674 = ~n247 & ~n646;
  assign n17675 = n4530 & n17674;
  assign n17676 = ~n184 & n4530;
  assign n17677 = ~n247 & n17676;
  assign n17678 = ~n441 & n17677;
  assign n17679 = ~n646 & n17678;
  assign n17680 = ~n441 & ~n646;
  assign n17681 = ~n184 & ~n247;
  assign n17682 = n17680 & n17681;
  assign n17683 = n4530 & n17682;
  assign n17684 = n5942 & n17675;
  assign n17685 = n7307 & n8752;
  assign n17686 = n11134 & n17685;
  assign n17687 = n4538 & n5362;
  assign n17688 = n1532 & n7275;
  assign n17689 = n17687 & n17688;
  assign n17690 = n17686 & n17689;
  assign n17691 = n55104 & n17690;
  assign n17692 = ~n420 & ~n499;
  assign n17693 = ~n1033 & ~n1195;
  assign n17694 = ~n420 & ~n1033;
  assign n17695 = ~n499 & ~n1195;
  assign n17696 = n17694 & n17695;
  assign n17697 = n17692 & n17693;
  assign n17698 = n850 & n3522;
  assign n17699 = n55105 & n17698;
  assign n17700 = ~n206 & ~n983;
  assign n17701 = ~n983 & n5873;
  assign n17702 = ~n206 & n17701;
  assign n17703 = n5873 & n17700;
  assign n17704 = n3015 & n55106;
  assign n17705 = n17699 & n17704;
  assign n17706 = n54784 & n17705;
  assign n17707 = n1532 & n7307;
  assign n17708 = n7275 & n17707;
  assign n17709 = n17687 & n17698;
  assign n17710 = n17708 & n17709;
  assign n17711 = n55104 & n17710;
  assign n17712 = n8752 & n11134;
  assign n17713 = n55105 & n17712;
  assign n17714 = n17704 & n17713;
  assign n17715 = n54784 & n17714;
  assign n17716 = n17711 & n17715;
  assign n17717 = n11134 & n17698;
  assign n17718 = n5362 & n7275;
  assign n17719 = n17707 & n17718;
  assign n17720 = n17717 & n17719;
  assign n17721 = n55104 & n17720;
  assign n17722 = n4538 & n8752;
  assign n17723 = n55105 & n17722;
  assign n17724 = n17704 & n17723;
  assign n17725 = n54784 & n17724;
  assign n17726 = n17721 & n17725;
  assign n17727 = n17691 & n17706;
  assign n17728 = n512 & ~n664;
  assign n17729 = n3819 & n4214;
  assign n17730 = n17728 & n17729;
  assign n17731 = ~n259 & ~n447;
  assign n17732 = ~n259 & ~n1079;
  assign n17733 = ~n447 & n17732;
  assign n17734 = ~n1079 & n17731;
  assign n17735 = n54775 & n55108;
  assign n17736 = n17730 & n17735;
  assign n17737 = n5069 & n6395;
  assign n17738 = n10593 & n15244;
  assign n17739 = n17737 & n17738;
  assign n17740 = n54600 & n17739;
  assign n17741 = n512 & n17735;
  assign n17742 = n3819 & n17741;
  assign n17743 = n54600 & n17742;
  assign n17744 = n424 & n17743;
  assign n17745 = n4214 & n17744;
  assign n17746 = ~n295 & n17745;
  assign n17747 = ~n1491 & n17746;
  assign n17748 = ~n1476 & n17747;
  assign n17749 = ~n166 & n17748;
  assign n17750 = ~n664 & n17749;
  assign n17751 = ~n353 & n17750;
  assign n17752 = ~n448 & n17751;
  assign n17753 = n512 & n3819;
  assign n17754 = ~n423 & ~n664;
  assign n17755 = ~n1491 & n17754;
  assign n17756 = n17753 & n17755;
  assign n17757 = n17735 & n17756;
  assign n17758 = n4214 & n6395;
  assign n17759 = n17738 & n17758;
  assign n17760 = n54600 & n17759;
  assign n17761 = n17757 & n17760;
  assign n17762 = ~n664 & n6395;
  assign n17763 = n4214 & n10593;
  assign n17764 = n17762 & n17763;
  assign n17765 = n17735 & n17764;
  assign n17766 = n3819 & n5069;
  assign n17767 = n512 & n15244;
  assign n17768 = n17766 & n17767;
  assign n17769 = n54600 & n17768;
  assign n17770 = n17765 & n17769;
  assign n17771 = ~n664 & n15244;
  assign n17772 = ~n295 & ~n1491;
  assign n17773 = ~n448 & ~n1476;
  assign n17774 = n17772 & n17773;
  assign n17775 = n17771 & n17774;
  assign n17776 = n17735 & n17775;
  assign n17777 = n424 & n4214;
  assign n17778 = n17753 & n17777;
  assign n17779 = n54600 & n17778;
  assign n17780 = n17776 & n17779;
  assign n17781 = n17736 & n17740;
  assign n17782 = n53814 & n55109;
  assign n17783 = n1532 & n3015;
  assign n17784 = n3522 & n17783;
  assign n17785 = n55106 & n17784;
  assign n17786 = n7275 & n17785;
  assign n17787 = n55104 & n17786;
  assign n17788 = n5362 & n17787;
  assign n17789 = n7307 & n17788;
  assign n17790 = n53814 & n17789;
  assign n17791 = n11134 & n17790;
  assign n17792 = n55109 & n17791;
  assign n17793 = n54784 & n17792;
  assign n17794 = n4538 & n17793;
  assign n17795 = n850 & n17794;
  assign n17796 = ~n1033 & n17795;
  assign n17797 = ~n1195 & n17796;
  assign n17798 = ~n310 & n17797;
  assign n17799 = ~n514 & n17798;
  assign n17800 = ~n499 & n17799;
  assign n17801 = ~n420 & n17800;
  assign n17802 = n55107 & n17782;
  assign n17803 = n10422 & ~n10424;
  assign n17804 = ~n10425 & ~n17803;
  assign n17805 = n1576 & n17804;
  assign n17806 = ~n54254 & n10564;
  assign n17807 = ~n54240 & n11215;
  assign n17808 = ~n54269 & n54403;
  assign n17809 = ~n17807 & ~n17808;
  assign n17810 = ~n17806 & n17809;
  assign n17811 = ~n17805 & ~n17808;
  assign n17812 = ~n17806 & n17811;
  assign n17813 = ~n17807 & n17812;
  assign n17814 = ~n17805 & n17810;
  assign n17815 = ~n55110 & ~n55111;
  assign n17816 = ~n105 & ~n567;
  assign n17817 = ~n1486 & n17816;
  assign n17818 = ~n1486 & n54192;
  assign n17819 = ~n105 & n17818;
  assign n17820 = ~n567 & n17819;
  assign n17821 = n54192 & n17817;
  assign n17822 = ~n255 & ~n584;
  assign n17823 = ~n733 & ~n879;
  assign n17824 = n17822 & n17823;
  assign n17825 = n3334 & n6396;
  assign n17826 = n1866 & n17825;
  assign n17827 = ~n879 & ~n975;
  assign n17828 = ~n255 & ~n444;
  assign n17829 = n17827 & n17828;
  assign n17830 = ~n584 & ~n733;
  assign n17831 = n3334 & n17830;
  assign n17832 = n1866 & n17831;
  assign n17833 = n17829 & n17832;
  assign n17834 = n17824 & n17826;
  assign n17835 = n55112 & n55113;
  assign n17836 = n4214 & n4381;
  assign n17837 = ~n911 & ~n1191;
  assign n17838 = n8753 & n17837;
  assign n17839 = n17836 & n17838;
  assign n17840 = ~n410 & ~n832;
  assign n17841 = ~n832 & ~n1487;
  assign n17842 = ~n410 & n17841;
  assign n17843 = ~n1487 & n17840;
  assign n17844 = n53896 & n55114;
  assign n17845 = n53896 & n8753;
  assign n17846 = n4381 & n17845;
  assign n17847 = n4214 & n17846;
  assign n17848 = ~n1191 & n17847;
  assign n17849 = ~n1487 & n17848;
  assign n17850 = ~n911 & n17849;
  assign n17851 = ~n832 & n17850;
  assign n17852 = ~n410 & n17851;
  assign n17853 = ~n832 & ~n911;
  assign n17854 = n4214 & n17853;
  assign n17855 = n4381 & n8753;
  assign n17856 = n17854 & n17855;
  assign n17857 = ~n410 & ~n1191;
  assign n17858 = ~n1487 & n17857;
  assign n17859 = n53896 & n17858;
  assign n17860 = n17856 & n17859;
  assign n17861 = n17839 & n17844;
  assign n17862 = n53669 & n54217;
  assign n17863 = n55115 & n17862;
  assign n17864 = n17835 & n17863;
  assign n17865 = ~n647 & ~n664;
  assign n17866 = ~n647 & ~n1062;
  assign n17867 = ~n664 & n17866;
  assign n17868 = ~n1062 & n17865;
  assign n17869 = n749 & n1716;
  assign n17870 = n55116 & n17869;
  assign n17871 = n54055 & n17870;
  assign n17872 = n6530 & n7018;
  assign n17873 = ~n496 & ~n1681;
  assign n17874 = n7789 & n17873;
  assign n17875 = n17872 & n17874;
  assign n17876 = n54796 & n17875;
  assign n17877 = ~n776 & n1277;
  assign n17878 = ~n296 & n1277;
  assign n17879 = ~n1455 & n17878;
  assign n17880 = ~n776 & n17879;
  assign n17881 = ~n776 & ~n1455;
  assign n17882 = ~n296 & n17881;
  assign n17883 = n1277 & n17882;
  assign n17884 = n9646 & n17877;
  assign n17885 = n53619 & n55117;
  assign n17886 = n17876 & n17885;
  assign n17887 = n6530 & n54055;
  assign n17888 = n55117 & n17887;
  assign n17889 = n53619 & n17888;
  assign n17890 = n54796 & n17889;
  assign n17891 = n749 & n17890;
  assign n17892 = n1716 & n17891;
  assign n17893 = ~n896 & n17892;
  assign n17894 = ~n1681 & n17893;
  assign n17895 = ~n1062 & n17894;
  assign n17896 = ~n664 & n17895;
  assign n17897 = ~n554 & n17896;
  assign n17898 = ~n275 & n17897;
  assign n17899 = ~n496 & n17898;
  assign n17900 = ~n647 & n17899;
  assign n17901 = ~n465 & n17900;
  assign n17902 = n749 & n17873;
  assign n17903 = n55116 & n17902;
  assign n17904 = n54055 & n17903;
  assign n17905 = n1716 & n6530;
  assign n17906 = n7018 & n7789;
  assign n17907 = n17905 & n17906;
  assign n17908 = n54796 & n17907;
  assign n17909 = n17885 & n17908;
  assign n17910 = n17904 & n17909;
  assign n17911 = ~n496 & n7018;
  assign n17912 = ~n664 & ~n1681;
  assign n17913 = n7789 & n17912;
  assign n17914 = n17911 & n17913;
  assign n17915 = n54055 & n17914;
  assign n17916 = n1716 & n17866;
  assign n17917 = n749 & n6530;
  assign n17918 = n17916 & n17917;
  assign n17919 = n54796 & n17918;
  assign n17920 = n17885 & n17919;
  assign n17921 = n17915 & n17920;
  assign n17922 = n17871 & n17886;
  assign n17923 = n54818 & n55118;
  assign n17924 = n1866 & n3334;
  assign n17925 = n55112 & n17924;
  assign n17926 = n54217 & n17925;
  assign n17927 = n53669 & n17926;
  assign n17928 = n54818 & n17927;
  assign n17929 = n55118 & n17928;
  assign n17930 = n55115 & n17929;
  assign n17931 = ~n879 & n17930;
  assign n17932 = ~n255 & n17931;
  assign n17933 = ~n584 & n17932;
  assign n17934 = ~n975 & n17933;
  assign n17935 = ~n733 & n17934;
  assign n17936 = ~n444 & n17935;
  assign n17937 = n17864 & n17923;
  assign n17938 = n10418 & ~n10420;
  assign n17939 = ~n10421 & ~n17938;
  assign n17940 = n1576 & n17939;
  assign n17941 = ~n54254 & n11215;
  assign n17942 = ~n54277 & n54403;
  assign n17943 = ~n54269 & n10564;
  assign n17944 = ~n17942 & ~n17943;
  assign n17945 = ~n17941 & n17944;
  assign n17946 = ~n17940 & ~n17942;
  assign n17947 = ~n17943 & n17946;
  assign n17948 = ~n17941 & n17947;
  assign n17949 = ~n17940 & n17945;
  assign n17950 = ~n55119 & ~n55120;
  assign n17951 = n343 & n1467;
  assign n17952 = n3474 & n6806;
  assign n17953 = n343 & n6806;
  assign n17954 = n1467 & n3474;
  assign n17955 = n17953 & n17954;
  assign n17956 = n17951 & n17952;
  assign n17957 = ~n1088 & ~n1127;
  assign n17958 = ~n984 & n17957;
  assign n17959 = ~n218 & ~n627;
  assign n17960 = ~n914 & ~n1081;
  assign n17961 = n17959 & n17960;
  assign n17962 = ~n984 & n17959;
  assign n17963 = n17957 & n17960;
  assign n17964 = n17962 & n17963;
  assign n17965 = ~n1081 & ~n1088;
  assign n17966 = ~n914 & n17965;
  assign n17967 = ~n984 & ~n1127;
  assign n17968 = n17959 & n17967;
  assign n17969 = n17966 & n17968;
  assign n17970 = n17958 & n17961;
  assign n17971 = n54553 & n55122;
  assign n17972 = n3474 & n54553;
  assign n17973 = n1467 & n17972;
  assign n17974 = n343 & n17973;
  assign n17975 = n6806 & n17974;
  assign n17976 = ~n984 & n17975;
  assign n17977 = ~n1088 & n17976;
  assign n17978 = ~n1127 & n17977;
  assign n17979 = ~n1081 & n17978;
  assign n17980 = ~n218 & n17979;
  assign n17981 = ~n914 & n17980;
  assign n17982 = ~n627 & n17981;
  assign n17983 = n55121 & n17971;
  assign n17984 = ~n423 & ~n663;
  assign n17985 = ~n748 & ~n879;
  assign n17986 = ~n663 & ~n879;
  assign n17987 = ~n423 & ~n748;
  assign n17988 = n17986 & n17987;
  assign n17989 = n17984 & n17985;
  assign n17990 = n6934 & n55124;
  assign n17991 = ~n349 & ~n1478;
  assign n17992 = n500 & ~n1478;
  assign n17993 = ~n349 & n17992;
  assign n17994 = n500 & n17991;
  assign n17995 = n54445 & n55125;
  assign n17996 = n17990 & n17995;
  assign n17997 = ~n513 & ~n735;
  assign n17998 = n355 & n17997;
  assign n17999 = n355 & n53621;
  assign n18000 = ~n513 & n17999;
  assign n18001 = ~n735 & n18000;
  assign n18002 = n53621 & n17998;
  assign n18003 = n976 & n5116;
  assign n18004 = n10037 & n13530;
  assign n18005 = n18003 & n18004;
  assign n18006 = n406 & n755;
  assign n18007 = n775 & n2693;
  assign n18008 = n755 & n2693;
  assign n18009 = n406 & n775;
  assign n18010 = n18008 & n18009;
  assign n18011 = n18006 & n18007;
  assign n18012 = n406 & n2693;
  assign n18013 = n976 & n13530;
  assign n18014 = n18012 & n18013;
  assign n18015 = n755 & n775;
  assign n18016 = n5116 & n10037;
  assign n18017 = n18015 & n18016;
  assign n18018 = n18014 & n18017;
  assign n18019 = n18005 & n55127;
  assign n18020 = n55126 & n55128;
  assign n18021 = ~n321 & ~n663;
  assign n18022 = n17985 & n18021;
  assign n18023 = n6934 & n18022;
  assign n18024 = n17995 & n18023;
  assign n18025 = n775 & n13530;
  assign n18026 = n18008 & n18025;
  assign n18027 = ~n423 & ~n1059;
  assign n18028 = n976 & n18027;
  assign n18029 = n406 & n5116;
  assign n18030 = n18028 & n18029;
  assign n18031 = n18026 & n18030;
  assign n18032 = n55126 & n18031;
  assign n18033 = n18024 & n18032;
  assign n18034 = n17996 & n18020;
  assign n18035 = n55123 & n55129;
  assign n18036 = n6934 & n55125;
  assign n18037 = n13530 & n18036;
  assign n18038 = n54445 & n18037;
  assign n18039 = n55126 & n18038;
  assign n18040 = n54201 & n18039;
  assign n18041 = n55123 & n18040;
  assign n18042 = n5116 & n18041;
  assign n18043 = n775 & n18042;
  assign n18044 = n755 & n18043;
  assign n18045 = n2693 & n18044;
  assign n18046 = n406 & n18045;
  assign n18047 = n976 & n18046;
  assign n18048 = ~n879 & n18047;
  assign n18049 = ~n321 & n18048;
  assign n18050 = ~n663 & n18049;
  assign n18051 = ~n1059 & n18050;
  assign n18052 = ~n748 & n18051;
  assign n18053 = ~n423 & n18052;
  assign n18054 = n54201 & n18035;
  assign n18055 = n10414 & ~n10416;
  assign n18056 = ~n10417 & ~n18055;
  assign n18057 = n1576 & n18056;
  assign n18058 = ~n54305 & n54403;
  assign n18059 = ~n54277 & n10564;
  assign n18060 = ~n54269 & n11215;
  assign n18061 = ~n18059 & ~n18060;
  assign n18062 = ~n18058 & n18061;
  assign n18063 = ~n18057 & ~n18058;
  assign n18064 = ~n18059 & n18063;
  assign n18065 = ~n18060 & n18064;
  assign n18066 = ~n18057 & n18062;
  assign n18067 = ~n55130 & ~n55131;
  assign n18068 = ~n495 & ~n552;
  assign n18069 = ~n922 & ~n1065;
  assign n18070 = n18068 & n18069;
  assign n18071 = ~n618 & ~n650;
  assign n18072 = n3001 & n18071;
  assign n18073 = n10301 & n18072;
  assign n18074 = n3001 & n10301;
  assign n18075 = ~n1065 & n18074;
  assign n18076 = ~n922 & n18075;
  assign n18077 = ~n552 & n18076;
  assign n18078 = ~n618 & n18077;
  assign n18079 = ~n495 & n18078;
  assign n18080 = ~n650 & n18079;
  assign n18081 = ~n552 & ~n650;
  assign n18082 = n18069 & n18081;
  assign n18083 = ~n495 & ~n618;
  assign n18084 = n3001 & n18083;
  assign n18085 = n10301 & n18084;
  assign n18086 = n18082 & n18085;
  assign n18087 = ~n495 & ~n650;
  assign n18088 = ~n618 & ~n922;
  assign n18089 = n18087 & n18088;
  assign n18090 = ~n552 & ~n1065;
  assign n18091 = n3001 & n18090;
  assign n18092 = n10301 & n18091;
  assign n18093 = n18089 & n18092;
  assign n18094 = n18070 & n18073;
  assign n18095 = ~n163 & ~n664;
  assign n18096 = ~n1031 & ~n1466;
  assign n18097 = ~n163 & ~n1466;
  assign n18098 = ~n664 & ~n1031;
  assign n18099 = n18097 & n18098;
  assign n18100 = n18095 & n18096;
  assign n18101 = n3819 & n4584;
  assign n18102 = n55133 & n18101;
  assign n18103 = n3062 & n4974;
  assign n18104 = n4003 & n18103;
  assign n18105 = n18102 & n18104;
  assign n18106 = ~n348 & ~n1715;
  assign n18107 = ~n348 & n11472;
  assign n18108 = ~n1715 & n18107;
  assign n18109 = n11472 & n18106;
  assign n18110 = n5377 & n7201;
  assign n18111 = n11492 & n17837;
  assign n18112 = n18110 & n18111;
  assign n18113 = n55134 & n18112;
  assign n18114 = n4002 & n4584;
  assign n18115 = n18103 & n18114;
  assign n18116 = ~n163 & ~n1191;
  assign n18117 = n11492 & n18116;
  assign n18118 = ~n664 & ~n911;
  assign n18119 = n18096 & n18118;
  assign n18120 = n18117 & n18119;
  assign n18121 = n18115 & n18120;
  assign n18122 = n3819 & n5377;
  assign n18123 = n903 & n7201;
  assign n18124 = n18122 & n18123;
  assign n18125 = n55134 & n18124;
  assign n18126 = n18121 & n18125;
  assign n18127 = n18105 & n18113;
  assign n18128 = n55132 & n55135;
  assign n18129 = n54167 & n18128;
  assign n18130 = n54448 & n54602;
  assign n18131 = n3819 & n4974;
  assign n18132 = n55134 & n18131;
  assign n18133 = n54602 & n18132;
  assign n18134 = n54167 & n18133;
  assign n18135 = n54448 & n18134;
  assign n18136 = n55132 & n18135;
  assign n18137 = n4584 & n18136;
  assign n18138 = n7201 & n18137;
  assign n18139 = n4002 & n18138;
  assign n18140 = n5377 & n18139;
  assign n18141 = n903 & n18140;
  assign n18142 = n3062 & n18141;
  assign n18143 = ~n1031 & n18142;
  assign n18144 = ~n1191 & n18143;
  assign n18145 = ~n1466 & n18144;
  assign n18146 = ~n1468 & n18145;
  assign n18147 = ~n163 & n18146;
  assign n18148 = ~n255 & n18147;
  assign n18149 = ~n664 & n18148;
  assign n18150 = ~n911 & n18149;
  assign n18151 = n18129 & n18130;
  assign n18152 = n54325 & ~n54344;
  assign n18153 = n54305 & ~n18152;
  assign n18154 = n54325 & n10406;
  assign n18155 = ~n54305 & n18152;
  assign n18156 = ~n18153 & ~n55137;
  assign n18157 = n1576 & n18156;
  assign n18158 = ~n54305 & n11215;
  assign n18159 = ~n54344 & n10564;
  assign n18160 = ~n54325 & n54403;
  assign n18161 = ~n18159 & ~n18160;
  assign n18162 = ~n18158 & n18161;
  assign n18163 = ~n18157 & ~n18160;
  assign n18164 = ~n18159 & n18163;
  assign n18165 = ~n18158 & n18164;
  assign n18166 = ~n18157 & n18162;
  assign n18167 = ~n55136 & ~n55138;
  assign n18168 = ~n340 & ~n344;
  assign n18169 = ~n495 & ~n1912;
  assign n18170 = n18168 & n18169;
  assign n18171 = ~n585 & ~n647;
  assign n18172 = n3535 & n18171;
  assign n18173 = ~n495 & ~n647;
  assign n18174 = n9828 & n18173;
  assign n18175 = n3535 & n18168;
  assign n18176 = n18174 & n18175;
  assign n18177 = ~n495 & ~n585;
  assign n18178 = ~n344 & ~n647;
  assign n18179 = n18177 & n18178;
  assign n18180 = ~n340 & ~n1912;
  assign n18181 = n3535 & n18180;
  assign n18182 = n18179 & n18181;
  assign n18183 = ~n344 & ~n1912;
  assign n18184 = n18177 & n18183;
  assign n18185 = ~n340 & ~n647;
  assign n18186 = n3535 & n18185;
  assign n18187 = n18184 & n18186;
  assign n18188 = n18170 & n18172;
  assign n18189 = n53964 & n10686;
  assign n18190 = n55139 & n18189;
  assign n18191 = ~n321 & ~n1124;
  assign n18192 = ~n1485 & n18191;
  assign n18193 = n8389 & n13650;
  assign n18194 = ~n1124 & ~n1485;
  assign n18195 = ~n1124 & n3001;
  assign n18196 = ~n1485 & n18195;
  assign n18197 = n3001 & n18194;
  assign n18198 = ~n163 & n55140;
  assign n18199 = ~n405 & n18198;
  assign n18200 = ~n562 & n18199;
  assign n18201 = ~n405 & ~n1124;
  assign n18202 = ~n1485 & n18201;
  assign n18203 = n3001 & n8389;
  assign n18204 = n18202 & n18203;
  assign n18205 = ~n562 & ~n1124;
  assign n18206 = ~n1485 & n18205;
  assign n18207 = ~n163 & ~n405;
  assign n18208 = n3001 & n18207;
  assign n18209 = n18206 & n18208;
  assign n18210 = ~n405 & ~n562;
  assign n18211 = ~n163 & n18210;
  assign n18212 = n55140 & n18211;
  assign n18213 = n18192 & n18193;
  assign n18214 = ~n144 & ~n504;
  assign n18215 = ~n144 & n1459;
  assign n18216 = ~n144 & n1458;
  assign n18217 = ~n504 & n18216;
  assign n18218 = n1458 & n18214;
  assign n18219 = n54064 & n55142;
  assign n18220 = n54064 & n55141;
  assign n18221 = n55142 & n18220;
  assign n18222 = n55141 & n18219;
  assign n18223 = n18189 & n55142;
  assign n18224 = n54064 & n55139;
  assign n18225 = n55141 & n18224;
  assign n18226 = n18223 & n18225;
  assign n18227 = n18190 & n55143;
  assign n18228 = n54298 & n55144;
  assign n18229 = n1265 & n1278;
  assign n18230 = n1265 & n2974;
  assign n18231 = n1278 & n18230;
  assign n18232 = n2974 & n18229;
  assign n18233 = ~n268 & ~n565;
  assign n18234 = ~n356 & ~n1715;
  assign n18235 = ~n565 & ~n1715;
  assign n18236 = ~n268 & ~n356;
  assign n18237 = n18235 & n18236;
  assign n18238 = ~n268 & ~n1715;
  assign n18239 = ~n356 & ~n565;
  assign n18240 = n18238 & n18239;
  assign n18241 = n18233 & n18234;
  assign n18242 = n7025 & n55146;
  assign n18243 = n2974 & n7025;
  assign n18244 = n1265 & n18243;
  assign n18245 = n1278 & n18244;
  assign n18246 = ~n565 & n18245;
  assign n18247 = ~n268 & n18246;
  assign n18248 = ~n356 & n18247;
  assign n18249 = ~n1715 & n18248;
  assign n18250 = n55145 & n18242;
  assign n18251 = ~n174 & ~n651;
  assign n18252 = n755 & n18251;
  assign n18253 = n846 & n4319;
  assign n18254 = n18252 & n18253;
  assign n18255 = ~n419 & ~n617;
  assign n18256 = ~n617 & n3283;
  assign n18257 = ~n419 & n18256;
  assign n18258 = n3283 & n18255;
  assign n18259 = ~n408 & ~n447;
  assign n18260 = ~n496 & ~n1535;
  assign n18261 = n18259 & n18260;
  assign n18262 = n55148 & n18261;
  assign n18263 = ~n447 & ~n496;
  assign n18264 = n755 & n18263;
  assign n18265 = n18253 & n18264;
  assign n18266 = ~n408 & ~n1535;
  assign n18267 = n18251 & n18266;
  assign n18268 = n55148 & n18267;
  assign n18269 = n18265 & n18268;
  assign n18270 = n18254 & n18262;
  assign n18271 = ~n2103 & n8274;
  assign n18272 = n1671 & n2038;
  assign n18273 = n2092 & n9210;
  assign n18274 = n18272 & n18273;
  assign n18275 = n18271 & n18274;
  assign n18276 = n755 & n18260;
  assign n18277 = n1671 & n4319;
  assign n18278 = n18276 & n18277;
  assign n18279 = ~n174 & ~n447;
  assign n18280 = ~n408 & ~n651;
  assign n18281 = n18279 & n18280;
  assign n18282 = n55148 & n18281;
  assign n18283 = n18278 & n18282;
  assign n18284 = n846 & n2038;
  assign n18285 = n18273 & n18284;
  assign n18286 = n18271 & n18285;
  assign n18287 = n18283 & n18286;
  assign n18288 = n4319 & n18279;
  assign n18289 = n846 & n1671;
  assign n18290 = n18288 & n18289;
  assign n18291 = ~n496 & ~n651;
  assign n18292 = n18266 & n18291;
  assign n18293 = n55148 & n18292;
  assign n18294 = n18290 & n18293;
  assign n18295 = n2038 & n2092;
  assign n18296 = n755 & n9210;
  assign n18297 = n18295 & n18296;
  assign n18298 = n18271 & n18297;
  assign n18299 = n18294 & n18298;
  assign n18300 = n55149 & n18275;
  assign n18301 = n9210 & n18271;
  assign n18302 = n55148 & n18301;
  assign n18303 = n2038 & n18302;
  assign n18304 = n2092 & n18303;
  assign n18305 = n846 & n18304;
  assign n18306 = n55147 & n18305;
  assign n18307 = n755 & n18306;
  assign n18308 = n1671 & n18307;
  assign n18309 = n4319 & n18308;
  assign n18310 = ~n408 & n18309;
  assign n18311 = ~n174 & n18310;
  assign n18312 = ~n1535 & n18311;
  assign n18313 = ~n496 & n18312;
  assign n18314 = ~n651 & n18313;
  assign n18315 = ~n447 & n18314;
  assign n18316 = n55147 & n55150;
  assign n18317 = n54015 & n55151;
  assign n18318 = n53964 & n55142;
  assign n18319 = n54064 & n18318;
  assign n18320 = n54298 & n18319;
  assign n18321 = n54015 & n18320;
  assign n18322 = n55151 & n18321;
  assign n18323 = n10686 & n18322;
  assign n18324 = n3535 & n18323;
  assign n18325 = n55141 & n18324;
  assign n18326 = ~n495 & n18325;
  assign n18327 = ~n647 & n18326;
  assign n18328 = ~n344 & n18327;
  assign n18329 = ~n340 & n18328;
  assign n18330 = ~n1912 & n18329;
  assign n18331 = ~n585 & n18330;
  assign n18332 = n18228 & n18317;
  assign n18333 = n18167 & ~n55152;
  assign n18334 = ~n18167 & n55152;
  assign n18335 = ~n9968 & n54346;
  assign n18336 = ~n10413 & ~n18335;
  assign n18337 = n1576 & n18336;
  assign n18338 = ~n54305 & n10564;
  assign n18339 = ~n54277 & n11215;
  assign n18340 = ~n54344 & n54403;
  assign n18341 = ~n18339 & ~n18340;
  assign n18342 = ~n18338 & ~n18340;
  assign n18343 = ~n18339 & n18342;
  assign n18344 = ~n18338 & n18341;
  assign n18345 = ~n18337 & n55153;
  assign n18346 = ~n18334 & ~n18345;
  assign n18347 = ~n18333 & ~n18334;
  assign n18348 = ~n18345 & n18347;
  assign n18349 = ~n18333 & ~n18348;
  assign n18350 = ~n18333 & ~n18346;
  assign n18351 = n55130 & n55131;
  assign n18352 = ~n55130 & ~n18067;
  assign n18353 = ~n55130 & n55131;
  assign n18354 = ~n55131 & ~n18067;
  assign n18355 = n55130 & ~n55131;
  assign n18356 = ~n55155 & ~n55156;
  assign n18357 = ~n18067 & ~n18351;
  assign n18358 = ~n55154 & ~n55157;
  assign n18359 = ~n18067 & ~n18358;
  assign n18360 = n55119 & n55120;
  assign n18361 = ~n55119 & ~n17950;
  assign n18362 = ~n55119 & n55120;
  assign n18363 = ~n55120 & ~n17950;
  assign n18364 = n55119 & ~n55120;
  assign n18365 = ~n55158 & ~n55159;
  assign n18366 = ~n17950 & ~n18360;
  assign n18367 = ~n18359 & ~n55160;
  assign n18368 = ~n17950 & ~n18367;
  assign n18369 = n55110 & n55111;
  assign n18370 = ~n55110 & ~n17815;
  assign n18371 = ~n55110 & n55111;
  assign n18372 = ~n55111 & ~n17815;
  assign n18373 = n55110 & ~n55111;
  assign n18374 = ~n55161 & ~n55162;
  assign n18375 = ~n17815 & ~n18369;
  assign n18376 = ~n18368 & ~n55163;
  assign n18377 = ~n17815 & ~n18376;
  assign n18378 = n55101 & n55103;
  assign n18379 = ~n55101 & ~n17673;
  assign n18380 = ~n55101 & n55103;
  assign n18381 = ~n55103 & ~n17673;
  assign n18382 = n55101 & ~n55103;
  assign n18383 = ~n55164 & ~n55165;
  assign n18384 = ~n17673 & ~n18378;
  assign n18385 = ~n18377 & ~n55166;
  assign n18386 = ~n17673 & ~n18385;
  assign n18387 = ~n17039 & n17050;
  assign n18388 = ~n17050 & ~n55004;
  assign n18389 = ~n17038 & n17054;
  assign n18390 = ~n18388 & ~n18389;
  assign n18391 = ~n55004 & ~n18387;
  assign n18392 = ~n18386 & ~n55167;
  assign n18393 = n18386 & n55167;
  assign n18394 = ~n18392 & ~n18393;
  assign n18395 = n11279 & n17072;
  assign n18396 = ~n54154 & n12584;
  assign n18397 = ~n54183 & n54410;
  assign n18398 = ~n54163 & n11267;
  assign n18399 = ~n18397 & ~n18398;
  assign n18400 = ~n18396 & n18399;
  assign n18401 = ~n11279 & n18400;
  assign n18402 = ~n17072 & n18400;
  assign n18403 = ~n18401 & ~n18402;
  assign n18404 = ~n18395 & n18400;
  assign n18405 = pi29  & ~n55168;
  assign n18406 = ~pi29  & n55168;
  assign n18407 = ~n18405 & ~n18406;
  assign n18408 = n18394 & ~n18407;
  assign n18409 = ~n18392 & ~n18408;
  assign n18410 = n55087 & n55088;
  assign n18411 = ~n55087 & ~n17555;
  assign n18412 = ~n55087 & n55088;
  assign n18413 = ~n55088 & ~n17555;
  assign n18414 = n55087 & ~n55088;
  assign n18415 = ~n55169 & ~n55170;
  assign n18416 = ~n17555 & ~n18410;
  assign n18417 = ~n18409 & ~n55171;
  assign n18418 = ~n17555 & ~n18417;
  assign n18419 = n55084 & n55086;
  assign n18420 = ~n55084 & ~n17537;
  assign n18421 = ~n55084 & n55086;
  assign n18422 = ~n55086 & ~n17537;
  assign n18423 = n55084 & ~n55086;
  assign n18424 = ~n55172 & ~n55173;
  assign n18425 = ~n17537 & ~n18419;
  assign n18426 = ~n18418 & ~n55174;
  assign n18427 = ~n17537 & ~n18426;
  assign n18428 = n17079 & ~n17081;
  assign n18429 = n17081 & ~n17082;
  assign n18430 = ~n17079 & ~n17082;
  assign n18431 = ~n18429 & ~n18430;
  assign n18432 = ~n17082 & ~n18428;
  assign n18433 = ~n18427 & ~n55175;
  assign n18434 = n18427 & n55175;
  assign n18435 = n11279 & n16547;
  assign n18436 = ~n54119 & n11267;
  assign n18437 = ~n54098 & n12584;
  assign n18438 = ~n54132 & n54410;
  assign n18439 = ~n18437 & ~n18438;
  assign n18440 = ~n18436 & ~n18438;
  assign n18441 = ~n18437 & n18440;
  assign n18442 = ~n18436 & n18439;
  assign n18443 = ~n18435 & n55176;
  assign n18444 = pi29  & ~n18443;
  assign n18445 = pi29  & ~n18444;
  assign n18446 = pi29  & n18443;
  assign n18447 = ~n18443 & ~n18444;
  assign n18448 = ~pi29  & ~n18443;
  assign n18449 = ~n55177 & ~n55178;
  assign n18450 = ~n18434 & ~n18449;
  assign n18451 = ~n18433 & ~n18434;
  assign n18452 = ~n18449 & n18451;
  assign n18453 = ~n18433 & ~n18452;
  assign n18454 = ~n18433 & ~n18450;
  assign n18455 = n17517 & ~n55179;
  assign n18456 = ~n17517 & n55179;
  assign n18457 = n123 & n15195;
  assign n18458 = n53444 & ~n54050;
  assign n18459 = n128 & ~n54005;
  assign n18460 = n127 & ~n54034;
  assign n18461 = ~n18459 & ~n18460;
  assign n18462 = ~n18458 & ~n18460;
  assign n18463 = ~n18459 & n18462;
  assign n18464 = ~n18458 & n18461;
  assign n18465 = ~n18457 & n55180;
  assign n18466 = pi26  & ~n18465;
  assign n18467 = pi26  & ~n18466;
  assign n18468 = pi26  & n18465;
  assign n18469 = ~n18465 & ~n18466;
  assign n18470 = ~pi26  & ~n18465;
  assign n18471 = ~n55181 & ~n55182;
  assign n18472 = ~n18456 & ~n18471;
  assign n18473 = ~n18455 & ~n18456;
  assign n18474 = ~n18471 & n18473;
  assign n18475 = ~n18455 & ~n18474;
  assign n18476 = ~n18455 & ~n18472;
  assign n18477 = ~n55083 & ~n55183;
  assign n18478 = n55083 & n55183;
  assign n18479 = n90 & n14263;
  assign n18480 = ~n53930 & n14210;
  assign n18481 = ~n53962 & n54667;
  assign n18482 = ~n53907 & n14236;
  assign n18483 = ~n18481 & ~n18482;
  assign n18484 = ~n18480 & ~n18481;
  assign n18485 = ~n18482 & n18484;
  assign n18486 = ~n18480 & n18483;
  assign n18487 = ~n18479 & n55184;
  assign n18488 = pi23  & ~n18487;
  assign n18489 = pi23  & ~n18488;
  assign n18490 = pi23  & n18487;
  assign n18491 = ~n18487 & ~n18488;
  assign n18492 = ~pi23  & ~n18487;
  assign n18493 = ~n55185 & ~n55186;
  assign n18494 = ~n18478 & ~n18493;
  assign n18495 = ~n18477 & ~n18478;
  assign n18496 = ~n18493 & n18495;
  assign n18497 = ~n18477 & ~n18496;
  assign n18498 = ~n18477 & ~n18494;
  assign n18499 = ~n55082 & ~n55187;
  assign n18500 = ~n17503 & ~n18499;
  assign n18501 = n17388 & ~n17389;
  assign n18502 = n17386 & n17388;
  assign n18503 = ~n17386 & ~n17389;
  assign n18504 = ~n17386 & ~n17388;
  assign n18505 = n17386 & ~n17388;
  assign n18506 = ~n17389 & ~n18505;
  assign n18507 = ~n55188 & ~n55189;
  assign n18508 = ~n18500 & n55190;
  assign n18509 = n18500 & ~n55190;
  assign n18510 = n12550 & n14413;
  assign n18511 = ~n53819 & n15901;
  assign n18512 = ~n53845 & n54719;
  assign n18513 = ~n53799 & n15921;
  assign n18514 = ~n18512 & ~n18513;
  assign n18515 = ~n18511 & ~n18512;
  assign n18516 = ~n18513 & n18515;
  assign n18517 = ~n18511 & n18514;
  assign n18518 = ~n18510 & n55191;
  assign n18519 = pi20  & ~n18518;
  assign n18520 = pi20  & ~n18519;
  assign n18521 = pi20  & n18518;
  assign n18522 = ~n18518 & ~n18519;
  assign n18523 = ~pi20  & ~n18518;
  assign n18524 = ~n55192 & ~n55193;
  assign n18525 = ~n18509 & ~n18524;
  assign n18526 = ~n18508 & ~n18509;
  assign n18527 = ~n18524 & n18526;
  assign n18528 = ~n18508 & ~n18527;
  assign n18529 = ~n18508 & ~n18525;
  assign n18530 = ~n55076 & ~n55194;
  assign n18531 = n55076 & n55194;
  assign n18532 = n11360 & n16079;
  assign n18533 = ~n53685 & n16696;
  assign n18534 = ~n53741 & n54886;
  assign n18535 = ~n53712 & n16676;
  assign n18536 = ~n18534 & ~n18535;
  assign n18537 = ~n18533 & ~n18534;
  assign n18538 = ~n18535 & n18537;
  assign n18539 = ~n18533 & n18536;
  assign n18540 = ~n18532 & n55195;
  assign n18541 = pi17  & ~n18540;
  assign n18542 = pi17  & ~n18541;
  assign n18543 = pi17  & n18540;
  assign n18544 = ~n18540 & ~n18541;
  assign n18545 = ~pi17  & ~n18540;
  assign n18546 = ~n55196 & ~n55197;
  assign n18547 = ~n18531 & ~n18546;
  assign n18548 = ~n18530 & ~n18531;
  assign n18549 = ~n18546 & n18548;
  assign n18550 = ~n18530 & ~n18549;
  assign n18551 = ~n18530 & ~n18547;
  assign n18552 = ~n55075 & ~n55198;
  assign n18553 = ~n17473 & ~n18552;
  assign n18554 = n54351 & n17265;
  assign n18555 = ~n53634 & n55041;
  assign n18556 = n55038 & ~n55039;
  assign n18557 = ~n2325 & n18556;
  assign n18558 = ~n18555 & ~n18557;
  assign n18559 = ~n17265 & n18558;
  assign n18560 = ~n54351 & n18558;
  assign n18561 = ~n18559 & ~n18560;
  assign n18562 = ~n18554 & n18558;
  assign n18563 = pi14  & ~n55199;
  assign n18564 = ~pi14  & n55199;
  assign n18565 = ~n18563 & ~n18564;
  assign n18566 = ~n18553 & ~n18565;
  assign n18567 = n18553 & n18565;
  assign n18568 = ~n18566 & ~n18567;
  assign n18569 = n17437 & ~n17438;
  assign n18570 = n17435 & n17437;
  assign n18571 = ~n17435 & ~n17438;
  assign n18572 = ~n17435 & ~n17437;
  assign n18573 = n17435 & ~n17437;
  assign n18574 = ~n17438 & ~n18573;
  assign n18575 = ~n55200 & ~n55201;
  assign n18576 = n18568 & n55202;
  assign n18577 = ~n18566 & ~n18576;
  assign n18578 = n55068 & ~n17449;
  assign n18579 = ~n55068 & ~n17450;
  assign n18580 = n17449 & ~n17450;
  assign n18581 = ~n18579 & ~n18580;
  assign n18582 = ~n17450 & ~n18578;
  assign n18583 = ~n18577 & ~n55203;
  assign n18584 = n18577 & n55203;
  assign n18585 = ~n18583 & ~n18584;
  assign n18586 = n11242 & n17265;
  assign n18587 = ~n53650 & n55041;
  assign n18588 = n55039 & ~n55040;
  assign n18589 = ~n2325 & n18588;
  assign n18590 = ~n53634 & n18556;
  assign n18591 = ~n18589 & ~n18590;
  assign n18592 = ~n18587 & ~n18590;
  assign n18593 = ~n18589 & n18592;
  assign n18594 = ~n18587 & n18591;
  assign n18595 = ~n17265 & n55204;
  assign n18596 = ~n11242 & n55204;
  assign n18597 = ~n18595 & ~n18596;
  assign n18598 = ~n18586 & n55204;
  assign n18599 = pi14  & ~n55205;
  assign n18600 = ~pi14  & n55205;
  assign n18601 = ~n18599 & ~n18600;
  assign n18602 = n18546 & ~n18548;
  assign n18603 = n18548 & ~n18549;
  assign n18604 = ~n18546 & ~n18549;
  assign n18605 = ~n18603 & ~n18604;
  assign n18606 = ~n18549 & ~n18602;
  assign n18607 = n55082 & n55187;
  assign n18608 = ~n18499 & ~n18607;
  assign n18609 = n12938 & n14413;
  assign n18610 = ~n53819 & n15921;
  assign n18611 = ~n53860 & n54719;
  assign n18612 = ~n53845 & n15901;
  assign n18613 = ~n18611 & ~n18612;
  assign n18614 = ~n18610 & ~n18611;
  assign n18615 = ~n18612 & n18614;
  assign n18616 = ~n18610 & n18613;
  assign n18617 = ~n14413 & n55207;
  assign n18618 = ~n12938 & n55207;
  assign n18619 = ~n18617 & ~n18618;
  assign n18620 = ~n18609 & n55207;
  assign n18621 = pi20  & ~n55208;
  assign n18622 = ~pi20  & n55208;
  assign n18623 = ~n18621 & ~n18622;
  assign n18624 = n18608 & ~n18623;
  assign n18625 = ~n18608 & n18623;
  assign n18626 = ~n18624 & ~n18625;
  assign n18627 = n18493 & ~n18495;
  assign n18628 = n18495 & ~n18496;
  assign n18629 = ~n18493 & ~n18496;
  assign n18630 = ~n18628 & ~n18629;
  assign n18631 = ~n18496 & ~n18627;
  assign n18632 = n123 & n15219;
  assign n18633 = n127 & ~n54050;
  assign n18634 = n128 & ~n54034;
  assign n18635 = n53444 & ~n54073;
  assign n18636 = ~n18634 & ~n18635;
  assign n18637 = ~n18633 & ~n18635;
  assign n18638 = ~n18634 & n18637;
  assign n18639 = ~n18633 & n18636;
  assign n18640 = ~n123 & n55210;
  assign n18641 = ~n15219 & n55210;
  assign n18642 = ~n18640 & ~n18641;
  assign n18643 = ~n18632 & n55210;
  assign n18644 = pi26  & ~n55211;
  assign n18645 = ~pi26  & n55211;
  assign n18646 = ~n18644 & ~n18645;
  assign n18647 = n18451 & ~n18452;
  assign n18648 = n18449 & n18451;
  assign n18649 = ~n18449 & ~n18452;
  assign n18650 = ~n18449 & ~n18451;
  assign n18651 = n18449 & ~n18451;
  assign n18652 = ~n18452 & ~n18651;
  assign n18653 = ~n55212 & ~n55213;
  assign n18654 = ~n18646 & n55214;
  assign n18655 = n18646 & ~n55214;
  assign n18656 = ~n18654 & ~n18655;
  assign n18657 = n11279 & n16772;
  assign n18658 = ~n54154 & n54410;
  assign n18659 = ~n54119 & n12584;
  assign n18660 = ~n54132 & n11267;
  assign n18661 = ~n18659 & ~n18660;
  assign n18662 = ~n18658 & ~n18660;
  assign n18663 = ~n18659 & n18662;
  assign n18664 = ~n18658 & n18661;
  assign n18665 = ~n11279 & n55215;
  assign n18666 = ~n16772 & n55215;
  assign n18667 = ~n18665 & ~n18666;
  assign n18668 = ~n18657 & n55215;
  assign n18669 = pi29  & ~n55216;
  assign n18670 = ~pi29  & n55216;
  assign n18671 = ~n18669 & ~n18670;
  assign n18672 = n18418 & n55174;
  assign n18673 = ~n18418 & ~n18426;
  assign n18674 = ~n55174 & ~n18426;
  assign n18675 = ~n18673 & ~n18674;
  assign n18676 = ~n18426 & ~n18672;
  assign n18677 = ~n18671 & ~n55217;
  assign n18678 = n18671 & n55217;
  assign n18679 = n123 & n16138;
  assign n18680 = n53444 & ~n54098;
  assign n18681 = n128 & ~n54050;
  assign n18682 = n127 & ~n54073;
  assign n18683 = ~n18681 & ~n18682;
  assign n18684 = ~n18680 & ~n18682;
  assign n18685 = ~n18681 & n18684;
  assign n18686 = ~n18680 & n18683;
  assign n18687 = ~n18679 & n55218;
  assign n18688 = pi26  & ~n18687;
  assign n18689 = pi26  & ~n18688;
  assign n18690 = pi26  & n18687;
  assign n18691 = ~n18687 & ~n18688;
  assign n18692 = ~pi26  & ~n18687;
  assign n18693 = ~n55219 & ~n55220;
  assign n18694 = ~n18678 & ~n18693;
  assign n18695 = ~n18677 & ~n18678;
  assign n18696 = ~n18693 & n18695;
  assign n18697 = ~n18677 & ~n18696;
  assign n18698 = ~n18677 & ~n18694;
  assign n18699 = n18656 & ~n55221;
  assign n18700 = ~n18654 & ~n18699;
  assign n18701 = n18471 & ~n18473;
  assign n18702 = n18473 & ~n18474;
  assign n18703 = ~n18471 & ~n18474;
  assign n18704 = ~n18702 & ~n18703;
  assign n18705 = ~n18474 & ~n18701;
  assign n18706 = ~n18700 & ~n55222;
  assign n18707 = n18700 & n55222;
  assign n18708 = n90 & n14020;
  assign n18709 = ~n53962 & n14210;
  assign n18710 = ~n53970 & n54667;
  assign n18711 = ~n53930 & n14236;
  assign n18712 = ~n18710 & ~n18711;
  assign n18713 = ~n18709 & ~n18710;
  assign n18714 = ~n18711 & n18713;
  assign n18715 = ~n18709 & n18712;
  assign n18716 = ~n18708 & n55223;
  assign n18717 = pi23  & ~n18716;
  assign n18718 = pi23  & ~n18717;
  assign n18719 = pi23  & n18716;
  assign n18720 = ~n18716 & ~n18717;
  assign n18721 = ~pi23  & ~n18716;
  assign n18722 = ~n55224 & ~n55225;
  assign n18723 = ~n18707 & ~n18722;
  assign n18724 = ~n18706 & ~n18707;
  assign n18725 = ~n18722 & n18724;
  assign n18726 = ~n18706 & ~n18725;
  assign n18727 = ~n18706 & ~n18723;
  assign n18728 = ~n55209 & ~n55226;
  assign n18729 = n55209 & n55226;
  assign n18730 = n12918 & n14413;
  assign n18731 = ~n53860 & n15901;
  assign n18732 = ~n53888 & n54719;
  assign n18733 = ~n53845 & n15921;
  assign n18734 = ~n18732 & ~n18733;
  assign n18735 = ~n18731 & ~n18732;
  assign n18736 = ~n18733 & n18735;
  assign n18737 = ~n18731 & n18734;
  assign n18738 = ~n18730 & n55227;
  assign n18739 = pi20  & ~n18738;
  assign n18740 = pi20  & ~n18739;
  assign n18741 = pi20  & n18738;
  assign n18742 = ~n18738 & ~n18739;
  assign n18743 = ~pi20  & ~n18738;
  assign n18744 = ~n55228 & ~n55229;
  assign n18745 = ~n18729 & ~n18744;
  assign n18746 = ~n18728 & ~n18729;
  assign n18747 = ~n18744 & n18746;
  assign n18748 = ~n18728 & ~n18747;
  assign n18749 = ~n18728 & ~n18745;
  assign n18750 = n18626 & ~n55230;
  assign n18751 = ~n18624 & ~n18750;
  assign n18752 = n18524 & ~n18526;
  assign n18753 = n18526 & ~n18527;
  assign n18754 = ~n18524 & ~n18527;
  assign n18755 = ~n18753 & ~n18754;
  assign n18756 = ~n18527 & ~n18752;
  assign n18757 = ~n18751 & ~n55231;
  assign n18758 = n18751 & n55231;
  assign n18759 = n11889 & n16079;
  assign n18760 = ~n53712 & n16696;
  assign n18761 = ~n53774 & n54886;
  assign n18762 = ~n53741 & n16676;
  assign n18763 = ~n18761 & ~n18762;
  assign n18764 = ~n18760 & ~n18761;
  assign n18765 = ~n18762 & n18764;
  assign n18766 = ~n18760 & n18763;
  assign n18767 = ~n18759 & n55232;
  assign n18768 = pi17  & ~n18767;
  assign n18769 = pi17  & ~n18768;
  assign n18770 = pi17  & n18767;
  assign n18771 = ~n18767 & ~n18768;
  assign n18772 = ~pi17  & ~n18767;
  assign n18773 = ~n55233 & ~n55234;
  assign n18774 = ~n18758 & ~n18773;
  assign n18775 = ~n18757 & ~n18758;
  assign n18776 = ~n18773 & n18775;
  assign n18777 = ~n18757 & ~n18776;
  assign n18778 = ~n18757 & ~n18774;
  assign n18779 = ~n55206 & ~n55235;
  assign n18780 = n55206 & n55235;
  assign n18781 = n11286 & n17265;
  assign n18782 = ~n53650 & n18556;
  assign n18783 = ~n53657 & n55041;
  assign n18784 = ~n53634 & n18588;
  assign n18785 = ~n18783 & ~n18784;
  assign n18786 = ~n18782 & ~n18783;
  assign n18787 = ~n18784 & n18786;
  assign n18788 = ~n18782 & n18785;
  assign n18789 = ~n18781 & n55236;
  assign n18790 = pi14  & ~n18789;
  assign n18791 = pi14  & ~n18790;
  assign n18792 = pi14  & n18789;
  assign n18793 = ~n18789 & ~n18790;
  assign n18794 = ~pi14  & ~n18789;
  assign n18795 = ~n55237 & ~n55238;
  assign n18796 = ~n18780 & ~n18795;
  assign n18797 = ~n18779 & ~n18780;
  assign n18798 = ~n18795 & n18797;
  assign n18799 = ~n18779 & ~n18798;
  assign n18800 = ~n18779 & ~n18796;
  assign n18801 = ~n18601 & ~n55239;
  assign n18802 = n55075 & n55198;
  assign n18803 = ~n18552 & ~n18802;
  assign n18804 = n18601 & n55239;
  assign n18805 = ~n55239 & ~n18801;
  assign n18806 = n18601 & ~n55239;
  assign n18807 = ~n18601 & ~n18801;
  assign n18808 = ~n18601 & n55239;
  assign n18809 = ~n55240 & ~n55241;
  assign n18810 = ~n18801 & ~n18804;
  assign n18811 = n18803 & ~n55242;
  assign n18812 = ~n18801 & ~n18811;
  assign n18813 = ~n18568 & ~n55202;
  assign n18814 = ~n18576 & ~n18813;
  assign n18815 = ~n18812 & n18814;
  assign n18816 = ~n18803 & ~n55241;
  assign n18817 = ~n55240 & n18816;
  assign n18818 = ~n18803 & ~n55240;
  assign n18819 = ~n55241 & n18818;
  assign n18820 = ~n18803 & n55242;
  assign n18821 = ~n18811 & ~n55243;
  assign n18822 = pi8  & ~pi9 ;
  assign n18823 = ~pi8  & pi9 ;
  assign n18824 = ~pi8  & ~pi9 ;
  assign n18825 = pi8  & pi9 ;
  assign n18826 = ~n18824 & ~n18825;
  assign n18827 = ~n18822 & ~n18823;
  assign n18828 = pi9  & ~pi10 ;
  assign n18829 = ~pi9  & pi10 ;
  assign n18830 = ~pi9  & ~pi10 ;
  assign n18831 = pi9  & pi10 ;
  assign n18832 = ~n18830 & ~n18831;
  assign n18833 = ~n18828 & ~n18829;
  assign n18834 = ~n55244 & ~n55245;
  assign n18835 = pi10  & ~pi11 ;
  assign n18836 = ~pi10  & pi11 ;
  assign n18837 = ~pi10  & ~pi11 ;
  assign n18838 = pi10  & pi11 ;
  assign n18839 = ~n18837 & ~n18838;
  assign n18840 = ~n18835 & ~n18836;
  assign n18841 = ~n55244 & n55246;
  assign n18842 = ~n55245 & n18841;
  assign n18843 = ~n55245 & n55246;
  assign n18844 = ~n55244 & n18843;
  assign n18845 = n18834 & n55246;
  assign n18846 = n55244 & n55246;
  assign n18847 = ~n10547 & n18846;
  assign n18848 = ~n55247 & ~n18847;
  assign n18849 = ~n2325 & n55247;
  assign n18850 = ~n10551 & ~n18849;
  assign n18851 = ~n18846 & ~n18849;
  assign n18852 = ~n18850 & ~n18851;
  assign n18853 = ~n2325 & ~n18848;
  assign n18854 = pi11  & ~n55248;
  assign n18855 = ~pi11  & n55248;
  assign n18856 = ~n18854 & ~n18855;
  assign n18857 = n11913 & n16079;
  assign n18858 = ~n53774 & n16676;
  assign n18859 = ~n53799 & n54886;
  assign n18860 = ~n53741 & n16696;
  assign n18861 = ~n18859 & ~n18860;
  assign n18862 = ~n18858 & ~n18859;
  assign n18863 = ~n18860 & n18862;
  assign n18864 = ~n18858 & n18861;
  assign n18865 = ~n18857 & n55249;
  assign n18866 = pi17  & ~n18865;
  assign n18867 = ~n18865 & ~n18866;
  assign n18868 = ~pi17  & ~n18865;
  assign n18869 = pi17  & ~n18866;
  assign n18870 = pi17  & n18865;
  assign n18871 = ~n55250 & ~n55251;
  assign n18872 = ~n18626 & n55230;
  assign n18873 = ~n18750 & ~n18872;
  assign n18874 = ~n18871 & n18873;
  assign n18875 = n18871 & ~n18873;
  assign n18876 = ~n18871 & ~n18874;
  assign n18877 = ~n18871 & ~n18873;
  assign n18878 = n18873 & ~n18874;
  assign n18879 = n18871 & n18873;
  assign n18880 = ~n55252 & ~n55253;
  assign n18881 = ~n18874 & ~n18875;
  assign n18882 = n18744 & ~n18746;
  assign n18883 = n18746 & ~n18747;
  assign n18884 = ~n18744 & ~n18747;
  assign n18885 = ~n18883 & ~n18884;
  assign n18886 = ~n18747 & ~n18882;
  assign n18887 = n90 & n14708;
  assign n18888 = ~n54005 & n54667;
  assign n18889 = ~n53970 & n14210;
  assign n18890 = ~n53962 & n14236;
  assign n18891 = ~n18889 & ~n18890;
  assign n18892 = ~n18888 & ~n18889;
  assign n18893 = ~n18890 & n18892;
  assign n18894 = ~n18888 & n18891;
  assign n18895 = ~n18887 & n55256;
  assign n18896 = pi23  & ~n18895;
  assign n18897 = ~n18895 & ~n18896;
  assign n18898 = ~pi23  & ~n18895;
  assign n18899 = pi23  & ~n18896;
  assign n18900 = pi23  & n18895;
  assign n18901 = ~n55257 & ~n55258;
  assign n18902 = ~n18656 & n55221;
  assign n18903 = ~n18699 & ~n18902;
  assign n18904 = ~n18901 & n18903;
  assign n18905 = n18901 & ~n18903;
  assign n18906 = ~n18901 & ~n18904;
  assign n18907 = ~n18901 & ~n18903;
  assign n18908 = n18903 & ~n18904;
  assign n18909 = n18901 & n18903;
  assign n18910 = ~n55259 & ~n55260;
  assign n18911 = ~n18904 & ~n18905;
  assign n18912 = n18693 & ~n18695;
  assign n18913 = n18695 & ~n18696;
  assign n18914 = ~n18693 & ~n18696;
  assign n18915 = ~n18913 & ~n18914;
  assign n18916 = ~n18696 & ~n18912;
  assign n18917 = n11279 & n16522;
  assign n18918 = ~n54154 & n11267;
  assign n18919 = ~n54132 & n12584;
  assign n18920 = ~n54163 & n54410;
  assign n18921 = ~n18919 & ~n18920;
  assign n18922 = ~n18918 & ~n18920;
  assign n18923 = ~n18919 & n18922;
  assign n18924 = ~n18918 & n18921;
  assign n18925 = ~n11279 & n55263;
  assign n18926 = ~n16522 & n55263;
  assign n18927 = ~n18925 & ~n18926;
  assign n18928 = ~n18917 & n55263;
  assign n18929 = pi29  & ~n55264;
  assign n18930 = ~pi29  & n55264;
  assign n18931 = ~n18929 & ~n18930;
  assign n18932 = n18409 & n55171;
  assign n18933 = ~n18409 & ~n18417;
  assign n18934 = ~n55171 & ~n18417;
  assign n18935 = ~n18933 & ~n18934;
  assign n18936 = ~n18417 & ~n18932;
  assign n18937 = ~n18931 & ~n55265;
  assign n18938 = n18931 & n55265;
  assign n18939 = n123 & n15779;
  assign n18940 = n127 & ~n54098;
  assign n18941 = n53444 & ~n54119;
  assign n18942 = n128 & ~n54073;
  assign n18943 = ~n18941 & ~n18942;
  assign n18944 = ~n18940 & ~n18941;
  assign n18945 = ~n18942 & n18944;
  assign n18946 = ~n18940 & ~n18942;
  assign n18947 = ~n18941 & n18946;
  assign n18948 = ~n18940 & n18943;
  assign n18949 = ~n18939 & n55266;
  assign n18950 = pi26  & ~n18949;
  assign n18951 = pi26  & ~n18950;
  assign n18952 = pi26  & n18949;
  assign n18953 = ~n18949 & ~n18950;
  assign n18954 = ~pi26  & ~n18949;
  assign n18955 = ~n55267 & ~n55268;
  assign n18956 = ~n18938 & ~n18955;
  assign n18957 = ~n18937 & ~n18938;
  assign n18958 = ~n18955 & n18957;
  assign n18959 = ~n18937 & ~n18958;
  assign n18960 = ~n18937 & ~n18956;
  assign n18961 = ~n55262 & ~n55269;
  assign n18962 = n55262 & n55269;
  assign n18963 = n90 & n14688;
  assign n18964 = ~n54005 & n14210;
  assign n18965 = ~n54034 & n54667;
  assign n18966 = ~n53970 & n14236;
  assign n18967 = ~n18965 & ~n18966;
  assign n18968 = ~n18964 & ~n18965;
  assign n18969 = ~n18966 & n18968;
  assign n18970 = ~n18964 & n18967;
  assign n18971 = ~n18963 & n55270;
  assign n18972 = pi23  & ~n18971;
  assign n18973 = pi23  & ~n18972;
  assign n18974 = pi23  & n18971;
  assign n18975 = ~n18971 & ~n18972;
  assign n18976 = ~pi23  & ~n18971;
  assign n18977 = ~n55271 & ~n55272;
  assign n18978 = ~n18962 & ~n18977;
  assign n18979 = ~n18961 & ~n18962;
  assign n18980 = ~n18977 & n18979;
  assign n18981 = ~n18961 & ~n18980;
  assign n18982 = ~n18961 & ~n18978;
  assign n18983 = ~n55261 & ~n55273;
  assign n18984 = ~n18904 & ~n18983;
  assign n18985 = n18724 & ~n18725;
  assign n18986 = n18722 & n18724;
  assign n18987 = ~n18722 & ~n18725;
  assign n18988 = ~n18722 & ~n18724;
  assign n18989 = n18722 & ~n18724;
  assign n18990 = ~n18725 & ~n18989;
  assign n18991 = ~n55274 & ~n55275;
  assign n18992 = ~n18984 & n55276;
  assign n18993 = n18984 & ~n55276;
  assign n18994 = n13336 & n14413;
  assign n18995 = ~n53888 & n15901;
  assign n18996 = ~n53907 & n54719;
  assign n18997 = ~n53860 & n15921;
  assign n18998 = ~n18996 & ~n18997;
  assign n18999 = ~n18995 & ~n18996;
  assign n19000 = ~n18997 & n18999;
  assign n19001 = ~n18995 & n18998;
  assign n19002 = ~n18994 & n55277;
  assign n19003 = pi20  & ~n19002;
  assign n19004 = pi20  & ~n19003;
  assign n19005 = pi20  & n19002;
  assign n19006 = ~n19002 & ~n19003;
  assign n19007 = ~pi20  & ~n19002;
  assign n19008 = ~n55278 & ~n55279;
  assign n19009 = ~n18993 & ~n19008;
  assign n19010 = ~n18992 & ~n18993;
  assign n19011 = ~n19008 & n19010;
  assign n19012 = ~n18992 & ~n19011;
  assign n19013 = ~n18992 & ~n19009;
  assign n19014 = ~n55255 & ~n55280;
  assign n19015 = n55255 & n55280;
  assign n19016 = n12690 & n16079;
  assign n19017 = ~n53774 & n16696;
  assign n19018 = ~n53819 & n54886;
  assign n19019 = ~n53799 & n16676;
  assign n19020 = ~n19018 & ~n19019;
  assign n19021 = ~n19017 & ~n19018;
  assign n19022 = ~n19019 & n19021;
  assign n19023 = ~n19017 & n19020;
  assign n19024 = ~n19016 & n55281;
  assign n19025 = pi17  & ~n19024;
  assign n19026 = pi17  & ~n19025;
  assign n19027 = pi17  & n19024;
  assign n19028 = ~n19024 & ~n19025;
  assign n19029 = ~pi17  & ~n19024;
  assign n19030 = ~n55282 & ~n55283;
  assign n19031 = ~n19015 & ~n19030;
  assign n19032 = ~n19014 & ~n19015;
  assign n19033 = ~n19030 & n19032;
  assign n19034 = ~n19014 & ~n19033;
  assign n19035 = ~n19014 & ~n19031;
  assign n19036 = ~n55254 & ~n55284;
  assign n19037 = ~n18874 & ~n19036;
  assign n19038 = n18775 & ~n18776;
  assign n19039 = n18773 & n18775;
  assign n19040 = ~n18773 & ~n18776;
  assign n19041 = ~n18773 & ~n18775;
  assign n19042 = n18773 & ~n18775;
  assign n19043 = ~n18776 & ~n19042;
  assign n19044 = ~n55285 & ~n55286;
  assign n19045 = ~n19037 & n55287;
  assign n19046 = n19037 & ~n55287;
  assign n19047 = n11213 & n17265;
  assign n19048 = ~n53650 & n18588;
  assign n19049 = ~n53685 & n55041;
  assign n19050 = ~n53657 & n18556;
  assign n19051 = ~n19049 & ~n19050;
  assign n19052 = ~n19048 & n19051;
  assign n19053 = ~n19047 & n19052;
  assign n19054 = pi14  & ~n19053;
  assign n19055 = pi14  & ~n19054;
  assign n19056 = pi14  & n19053;
  assign n19057 = ~n19053 & ~n19054;
  assign n19058 = ~pi14  & ~n19053;
  assign n19059 = ~n55288 & ~n55289;
  assign n19060 = ~n19046 & ~n19059;
  assign n19061 = ~n19045 & ~n19046;
  assign n19062 = ~n19059 & n19061;
  assign n19063 = ~n19045 & ~n19062;
  assign n19064 = ~n19045 & ~n19060;
  assign n19065 = ~n18856 & ~n55290;
  assign n19066 = n18856 & n55290;
  assign n19067 = n18795 & ~n18797;
  assign n19068 = n18797 & ~n18798;
  assign n19069 = ~n18795 & ~n18798;
  assign n19070 = ~n19068 & ~n19069;
  assign n19071 = ~n18798 & ~n19067;
  assign n19072 = ~n19066 & ~n55291;
  assign n19073 = ~n19065 & ~n19066;
  assign n19074 = ~n55291 & n19073;
  assign n19075 = ~n19065 & ~n19074;
  assign n19076 = ~n19065 & ~n19072;
  assign n19077 = n18821 & ~n55292;
  assign n19078 = n55254 & n55284;
  assign n19079 = ~n19036 & ~n19078;
  assign n19080 = n11380 & n17265;
  assign n19081 = ~n53685 & n18556;
  assign n19082 = ~n53657 & n18588;
  assign n19083 = ~n53712 & n55041;
  assign n19084 = ~n19082 & ~n19083;
  assign n19085 = ~n19081 & ~n19083;
  assign n19086 = ~n19082 & n19085;
  assign n19087 = ~n19081 & n19084;
  assign n19088 = ~n17265 & n55293;
  assign n19089 = ~n11380 & n55293;
  assign n19090 = ~n19088 & ~n19089;
  assign n19091 = ~n19080 & n55293;
  assign n19092 = pi14  & ~n55294;
  assign n19093 = ~pi14  & n55294;
  assign n19094 = ~n19092 & ~n19093;
  assign n19095 = n19079 & ~n19094;
  assign n19096 = ~n19079 & n19094;
  assign n19097 = n19079 & ~n19095;
  assign n19098 = n19079 & n19094;
  assign n19099 = ~n19094 & ~n19095;
  assign n19100 = ~n19079 & ~n19094;
  assign n19101 = ~n55295 & ~n55296;
  assign n19102 = ~n19095 & ~n19096;
  assign n19103 = n19030 & ~n19032;
  assign n19104 = n19032 & ~n19033;
  assign n19105 = ~n19030 & ~n19033;
  assign n19106 = ~n19104 & ~n19105;
  assign n19107 = ~n19033 & ~n19103;
  assign n19108 = n55261 & n55273;
  assign n19109 = ~n18983 & ~n19108;
  assign n19110 = n13360 & n14413;
  assign n19111 = ~n53907 & n15901;
  assign n19112 = ~n53930 & n54719;
  assign n19113 = ~n53888 & n15921;
  assign n19114 = ~n19112 & ~n19113;
  assign n19115 = ~n19111 & ~n19112;
  assign n19116 = ~n19113 & n19115;
  assign n19117 = ~n19111 & n19114;
  assign n19118 = ~n14413 & n55299;
  assign n19119 = ~n13360 & n55299;
  assign n19120 = ~n19118 & ~n19119;
  assign n19121 = ~n19110 & n55299;
  assign n19122 = pi20  & ~n55300;
  assign n19123 = ~pi20  & n55300;
  assign n19124 = ~n19122 & ~n19123;
  assign n19125 = n19109 & ~n19124;
  assign n19126 = ~n19109 & n19124;
  assign n19127 = ~n19125 & ~n19126;
  assign n19128 = n18977 & ~n18979;
  assign n19129 = n18979 & ~n18980;
  assign n19130 = ~n18977 & ~n18980;
  assign n19131 = ~n19129 & ~n19130;
  assign n19132 = ~n18980 & ~n19128;
  assign n19133 = n11279 & n17524;
  assign n19134 = ~n54183 & n11267;
  assign n19135 = ~n54194 & n54410;
  assign n19136 = ~n54163 & n12584;
  assign n19137 = ~n19135 & ~n19136;
  assign n19138 = ~n19134 & ~n19135;
  assign n19139 = ~n19136 & n19138;
  assign n19140 = ~n19134 & n19137;
  assign n19141 = ~n11279 & n55302;
  assign n19142 = ~n17524 & n55302;
  assign n19143 = ~n19141 & ~n19142;
  assign n19144 = ~n19133 & n55302;
  assign n19145 = pi29  & ~n55303;
  assign n19146 = ~pi29  & n55303;
  assign n19147 = ~n19145 & ~n19146;
  assign n19148 = n18377 & n55166;
  assign n19149 = ~n18377 & ~n18385;
  assign n19150 = ~n55166 & ~n18385;
  assign n19151 = ~n19149 & ~n19150;
  assign n19152 = ~n18385 & ~n19148;
  assign n19153 = ~n19147 & ~n55304;
  assign n19154 = n11279 & n17544;
  assign n19155 = ~n54212 & n54410;
  assign n19156 = ~n54183 & n12584;
  assign n19157 = ~n54194 & n11267;
  assign n19158 = ~n19156 & ~n19157;
  assign n19159 = ~n19155 & ~n19157;
  assign n19160 = ~n19156 & n19159;
  assign n19161 = ~n19155 & n19158;
  assign n19162 = ~n11279 & n55305;
  assign n19163 = ~n17544 & n55305;
  assign n19164 = ~n19162 & ~n19163;
  assign n19165 = ~n19154 & n55305;
  assign n19166 = pi29  & ~n55306;
  assign n19167 = ~pi29  & n55306;
  assign n19168 = ~n19166 & ~n19167;
  assign n19169 = n18368 & n55163;
  assign n19170 = ~n18368 & ~n18376;
  assign n19171 = ~n55163 & ~n18376;
  assign n19172 = ~n19170 & ~n19171;
  assign n19173 = ~n18376 & ~n19169;
  assign n19174 = ~n19168 & ~n55307;
  assign n19175 = n11279 & n17041;
  assign n19176 = ~n54212 & n11267;
  assign n19177 = ~n54194 & n12584;
  assign n19178 = ~n54240 & n54410;
  assign n19179 = ~n19177 & ~n19178;
  assign n19180 = ~n19176 & ~n19178;
  assign n19181 = ~n19177 & n19180;
  assign n19182 = ~n19176 & n19179;
  assign n19183 = ~n19175 & n55308;
  assign n19184 = pi29  & ~n19183;
  assign n19185 = ~n19183 & ~n19184;
  assign n19186 = ~pi29  & ~n19183;
  assign n19187 = pi29  & ~n19184;
  assign n19188 = pi29  & n19183;
  assign n19189 = ~n55309 & ~n55310;
  assign n19190 = n18359 & n55160;
  assign n19191 = ~n18359 & ~n18367;
  assign n19192 = ~n55160 & ~n18367;
  assign n19193 = ~n19191 & ~n19192;
  assign n19194 = ~n18367 & ~n19190;
  assign n19195 = ~n19189 & ~n55311;
  assign n19196 = n11279 & n17660;
  assign n19197 = ~n54254 & n54410;
  assign n19198 = ~n54212 & n12584;
  assign n19199 = ~n54240 & n11267;
  assign n19200 = ~n19198 & ~n19199;
  assign n19201 = ~n19197 & ~n19199;
  assign n19202 = ~n19198 & n19201;
  assign n19203 = ~n19197 & n19200;
  assign n19204 = ~n19196 & n55312;
  assign n19205 = pi29  & ~n19204;
  assign n19206 = ~n19204 & ~n19205;
  assign n19207 = ~pi29  & ~n19204;
  assign n19208 = pi29  & ~n19205;
  assign n19209 = pi29  & n19204;
  assign n19210 = ~n55313 & ~n55314;
  assign n19211 = n55154 & n55157;
  assign n19212 = ~n55154 & ~n18358;
  assign n19213 = ~n55157 & ~n18358;
  assign n19214 = ~n19212 & ~n19213;
  assign n19215 = ~n18358 & ~n19211;
  assign n19216 = ~n19210 & ~n55315;
  assign n19217 = n11279 & n17804;
  assign n19218 = ~n54254 & n11267;
  assign n19219 = ~n54240 & n12584;
  assign n19220 = ~n54269 & n54410;
  assign n19221 = ~n19219 & ~n19220;
  assign n19222 = ~n19218 & ~n19220;
  assign n19223 = ~n19219 & n19222;
  assign n19224 = ~n19218 & n19221;
  assign n19225 = ~n19217 & n55316;
  assign n19226 = pi29  & ~n19225;
  assign n19227 = ~n19225 & ~n19226;
  assign n19228 = ~pi29  & ~n19225;
  assign n19229 = pi29  & ~n19226;
  assign n19230 = pi29  & n19225;
  assign n19231 = ~n55317 & ~n55318;
  assign n19232 = n18345 & ~n18347;
  assign n19233 = ~n18345 & ~n18348;
  assign n19234 = n18347 & ~n18348;
  assign n19235 = ~n19233 & ~n19234;
  assign n19236 = ~n18348 & ~n19232;
  assign n19237 = ~n19231 & ~n55319;
  assign n19238 = n11279 & n17939;
  assign n19239 = ~n54254 & n12584;
  assign n19240 = ~n54277 & n54410;
  assign n19241 = ~n54269 & n11267;
  assign n19242 = ~n19240 & ~n19241;
  assign n19243 = ~n19239 & n19242;
  assign n19244 = ~n19238 & n19243;
  assign n19245 = pi29  & ~n19244;
  assign n19246 = ~n19244 & ~n19245;
  assign n19247 = ~pi29  & ~n19244;
  assign n19248 = pi29  & ~n19245;
  assign n19249 = pi29  & n19244;
  assign n19250 = ~n55320 & ~n55321;
  assign n19251 = n55136 & n55138;
  assign n19252 = ~n55136 & ~n18167;
  assign n19253 = ~n55136 & n55138;
  assign n19254 = ~n55138 & ~n18167;
  assign n19255 = n55136 & ~n55138;
  assign n19256 = ~n55322 & ~n55323;
  assign n19257 = ~n18167 & ~n19251;
  assign n19258 = ~n19250 & ~n55324;
  assign n19259 = n11279 & n18056;
  assign n19260 = ~n54305 & n54410;
  assign n19261 = ~n54277 & n11267;
  assign n19262 = ~n54269 & n12584;
  assign n19263 = ~n19261 & ~n19262;
  assign n19264 = ~n19260 & ~n19261;
  assign n19265 = ~n19262 & n19264;
  assign n19266 = ~n19260 & n19263;
  assign n19267 = ~n19259 & n55325;
  assign n19268 = pi29  & ~n19267;
  assign n19269 = ~n19267 & ~n19268;
  assign n19270 = ~pi29  & ~n19267;
  assign n19271 = pi29  & ~n19268;
  assign n19272 = pi29  & n19267;
  assign n19273 = ~n55326 & ~n55327;
  assign n19274 = ~n54325 & n54344;
  assign n19275 = ~n18152 & ~n19274;
  assign n19276 = n1576 & ~n19275;
  assign n19277 = ~n54325 & n10564;
  assign n19278 = ~n54344 & n11215;
  assign n19279 = ~n19277 & ~n19278;
  assign n19280 = ~n19276 & n19279;
  assign n19281 = ~n19273 & ~n19280;
  assign n19282 = ~n94 & ~n54325;
  assign n19283 = n11279 & ~n19275;
  assign n19284 = ~n54325 & n11267;
  assign n19285 = ~n54344 & n12584;
  assign n19286 = ~n19284 & ~n19285;
  assign n19287 = ~n19283 & n19286;
  assign n19288 = ~n54325 & n54407;
  assign n19289 = pi29  & ~n19288;
  assign n19290 = pi29  & ~n19287;
  assign n19291 = pi29  & ~n19290;
  assign n19292 = ~n19287 & ~n19290;
  assign n19293 = ~n19291 & ~n19292;
  assign n19294 = n19289 & ~n19293;
  assign n19295 = n19287 & n19289;
  assign n19296 = n11279 & n18156;
  assign n19297 = ~n54305 & n12584;
  assign n19298 = ~n54325 & n54410;
  assign n19299 = ~n54344 & n11267;
  assign n19300 = ~n19298 & ~n19299;
  assign n19301 = ~n19297 & n19300;
  assign n19302 = ~n11279 & n19301;
  assign n19303 = ~n18156 & n19301;
  assign n19304 = ~n19302 & ~n19303;
  assign n19305 = ~n19296 & n19301;
  assign n19306 = pi29  & ~n55329;
  assign n19307 = ~pi29  & n55329;
  assign n19308 = ~n19306 & ~n19307;
  assign n19309 = n55328 & ~n19308;
  assign n19310 = n55328 & ~n55329;
  assign n19311 = n19282 & n55330;
  assign n19312 = n11279 & n18336;
  assign n19313 = ~n54305 & n11267;
  assign n19314 = ~n54277 & n12584;
  assign n19315 = ~n54344 & n54410;
  assign n19316 = ~n19314 & ~n19315;
  assign n19317 = ~n19313 & ~n19315;
  assign n19318 = ~n19314 & n19317;
  assign n19319 = ~n19313 & n19316;
  assign n19320 = ~n19312 & n55331;
  assign n19321 = pi29  & ~n19320;
  assign n19322 = ~n19320 & ~n19321;
  assign n19323 = ~pi29  & ~n19320;
  assign n19324 = pi29  & ~n19321;
  assign n19325 = pi29  & n19320;
  assign n19326 = ~n55332 & ~n55333;
  assign n19327 = ~n19282 & ~n55330;
  assign n19328 = ~n19282 & n55330;
  assign n19329 = n19282 & ~n55330;
  assign n19330 = ~n19328 & ~n19329;
  assign n19331 = ~n19311 & ~n19327;
  assign n19332 = ~n19326 & ~n55334;
  assign n19333 = ~n19311 & ~n19332;
  assign n19334 = n19273 & n19280;
  assign n19335 = ~n19273 & ~n19281;
  assign n19336 = ~n19273 & n19280;
  assign n19337 = ~n19280 & ~n19281;
  assign n19338 = n19273 & ~n19280;
  assign n19339 = ~n55335 & ~n55336;
  assign n19340 = ~n19281 & ~n19334;
  assign n19341 = ~n19333 & ~n55337;
  assign n19342 = ~n19281 & ~n19341;
  assign n19343 = n19250 & n55324;
  assign n19344 = ~n19250 & ~n19258;
  assign n19345 = ~n55324 & ~n19258;
  assign n19346 = ~n19344 & ~n19345;
  assign n19347 = ~n19258 & ~n19343;
  assign n19348 = ~n19342 & ~n55338;
  assign n19349 = ~n19258 & ~n19348;
  assign n19350 = n19231 & n55319;
  assign n19351 = ~n19231 & ~n19237;
  assign n19352 = ~n55319 & ~n19237;
  assign n19353 = ~n19351 & ~n19352;
  assign n19354 = ~n19237 & ~n19350;
  assign n19355 = ~n19349 & ~n55339;
  assign n19356 = ~n19237 & ~n19355;
  assign n19357 = n19210 & n55315;
  assign n19358 = ~n19210 & ~n19216;
  assign n19359 = ~n19210 & n55315;
  assign n19360 = ~n55315 & ~n19216;
  assign n19361 = n19210 & ~n55315;
  assign n19362 = ~n55340 & ~n55341;
  assign n19363 = ~n19216 & ~n19357;
  assign n19364 = ~n19356 & ~n55342;
  assign n19365 = ~n19216 & ~n19364;
  assign n19366 = n19189 & n55311;
  assign n19367 = ~n19189 & ~n19195;
  assign n19368 = ~n19189 & n55311;
  assign n19369 = ~n55311 & ~n19195;
  assign n19370 = n19189 & ~n55311;
  assign n19371 = ~n55343 & ~n55344;
  assign n19372 = ~n19195 & ~n19366;
  assign n19373 = ~n19365 & ~n55345;
  assign n19374 = ~n19195 & ~n19373;
  assign n19375 = n19168 & n55307;
  assign n19376 = ~n19174 & ~n19375;
  assign n19377 = ~n19374 & n19376;
  assign n19378 = ~n19174 & ~n19377;
  assign n19379 = n19147 & n55304;
  assign n19380 = ~n19153 & ~n19379;
  assign n19381 = ~n19378 & n19380;
  assign n19382 = ~n19153 & ~n19381;
  assign n19383 = ~n18394 & n18407;
  assign n19384 = ~n18408 & ~n19383;
  assign n19385 = ~n19382 & n19384;
  assign n19386 = n123 & n16547;
  assign n19387 = n127 & ~n54119;
  assign n19388 = n128 & ~n54098;
  assign n19389 = n53444 & ~n54132;
  assign n19390 = ~n19388 & ~n19389;
  assign n19391 = ~n19387 & ~n19389;
  assign n19392 = ~n19388 & n19391;
  assign n19393 = ~n19387 & n19390;
  assign n19394 = ~n19386 & n55346;
  assign n19395 = pi26  & ~n19394;
  assign n19396 = ~n19394 & ~n19395;
  assign n19397 = ~pi26  & ~n19394;
  assign n19398 = pi26  & ~n19395;
  assign n19399 = pi26  & n19394;
  assign n19400 = ~n55347 & ~n55348;
  assign n19401 = n19382 & ~n19384;
  assign n19402 = ~n19385 & ~n19401;
  assign n19403 = ~n19400 & n19402;
  assign n19404 = ~n19385 & ~n19403;
  assign n19405 = n18955 & ~n18957;
  assign n19406 = n18957 & ~n18958;
  assign n19407 = ~n18955 & ~n18958;
  assign n19408 = ~n19406 & ~n19407;
  assign n19409 = ~n18958 & ~n19405;
  assign n19410 = ~n19404 & ~n55349;
  assign n19411 = n19404 & n55349;
  assign n19412 = n90 & n15195;
  assign n19413 = ~n54050 & n54667;
  assign n19414 = ~n54005 & n14236;
  assign n19415 = ~n54034 & n14210;
  assign n19416 = ~n19414 & ~n19415;
  assign n19417 = ~n19413 & ~n19415;
  assign n19418 = ~n19414 & n19417;
  assign n19419 = ~n19413 & n19416;
  assign n19420 = ~n19412 & n55350;
  assign n19421 = pi23  & ~n19420;
  assign n19422 = pi23  & ~n19421;
  assign n19423 = pi23  & n19420;
  assign n19424 = ~n19420 & ~n19421;
  assign n19425 = ~pi23  & ~n19420;
  assign n19426 = ~n55351 & ~n55352;
  assign n19427 = ~n19411 & ~n19426;
  assign n19428 = ~n19410 & ~n19411;
  assign n19429 = ~n19426 & n19428;
  assign n19430 = ~n19410 & ~n19429;
  assign n19431 = ~n19410 & ~n19427;
  assign n19432 = ~n55301 & ~n55353;
  assign n19433 = n55301 & n55353;
  assign n19434 = n14263 & n14413;
  assign n19435 = ~n53930 & n15901;
  assign n19436 = ~n53962 & n54719;
  assign n19437 = ~n53907 & n15921;
  assign n19438 = ~n19436 & ~n19437;
  assign n19439 = ~n19435 & ~n19436;
  assign n19440 = ~n19437 & n19439;
  assign n19441 = ~n19435 & n19438;
  assign n19442 = ~n19434 & n55354;
  assign n19443 = pi20  & ~n19442;
  assign n19444 = pi20  & ~n19443;
  assign n19445 = pi20  & n19442;
  assign n19446 = ~n19442 & ~n19443;
  assign n19447 = ~pi20  & ~n19442;
  assign n19448 = ~n55355 & ~n55356;
  assign n19449 = ~n19433 & ~n19448;
  assign n19450 = ~n19432 & ~n19433;
  assign n19451 = ~n19448 & n19450;
  assign n19452 = ~n19432 & ~n19451;
  assign n19453 = ~n19432 & ~n19449;
  assign n19454 = n19127 & ~n55357;
  assign n19455 = ~n19125 & ~n19454;
  assign n19456 = n19008 & ~n19010;
  assign n19457 = n19010 & ~n19011;
  assign n19458 = ~n19008 & ~n19011;
  assign n19459 = ~n19457 & ~n19458;
  assign n19460 = ~n19011 & ~n19456;
  assign n19461 = ~n19455 & ~n55358;
  assign n19462 = n19455 & n55358;
  assign n19463 = n12550 & n16079;
  assign n19464 = ~n53819 & n16676;
  assign n19465 = ~n53845 & n54886;
  assign n19466 = ~n53799 & n16696;
  assign n19467 = ~n19465 & ~n19466;
  assign n19468 = ~n19464 & ~n19465;
  assign n19469 = ~n19466 & n19468;
  assign n19470 = ~n19464 & n19467;
  assign n19471 = ~n19463 & n55359;
  assign n19472 = pi17  & ~n19471;
  assign n19473 = pi17  & ~n19472;
  assign n19474 = pi17  & n19471;
  assign n19475 = ~n19471 & ~n19472;
  assign n19476 = ~pi17  & ~n19471;
  assign n19477 = ~n55360 & ~n55361;
  assign n19478 = ~n19462 & ~n19477;
  assign n19479 = ~n19461 & ~n19462;
  assign n19480 = ~n19477 & n19479;
  assign n19481 = ~n19461 & ~n19480;
  assign n19482 = ~n19461 & ~n19478;
  assign n19483 = ~n55298 & ~n55362;
  assign n19484 = n55298 & n55362;
  assign n19485 = n11360 & n17265;
  assign n19486 = ~n53685 & n18588;
  assign n19487 = ~n53741 & n55041;
  assign n19488 = ~n53712 & n18556;
  assign n19489 = ~n19487 & ~n19488;
  assign n19490 = ~n19486 & ~n19487;
  assign n19491 = ~n19488 & n19490;
  assign n19492 = ~n19486 & n19489;
  assign n19493 = ~n19485 & n55363;
  assign n19494 = pi14  & ~n19493;
  assign n19495 = pi14  & ~n19494;
  assign n19496 = pi14  & n19493;
  assign n19497 = ~n19493 & ~n19494;
  assign n19498 = ~pi14  & ~n19493;
  assign n19499 = ~n55364 & ~n55365;
  assign n19500 = ~n19484 & ~n19499;
  assign n19501 = ~n19483 & ~n19484;
  assign n19502 = ~n19499 & n19501;
  assign n19503 = ~n19483 & ~n19502;
  assign n19504 = ~n19483 & ~n19500;
  assign n19505 = ~n55297 & ~n55366;
  assign n19506 = ~n19095 & ~n19505;
  assign n19507 = n54351 & n18846;
  assign n19508 = ~n53634 & n55247;
  assign n19509 = ~n55244 & n55245;
  assign n19510 = ~n2325 & n19509;
  assign n19511 = ~n19508 & ~n19510;
  assign n19512 = ~n18846 & n19511;
  assign n19513 = ~n54351 & n19511;
  assign n19514 = ~n19512 & ~n19513;
  assign n19515 = ~n19507 & n19511;
  assign n19516 = pi11  & ~n55367;
  assign n19517 = ~pi11  & n55367;
  assign n19518 = ~n19516 & ~n19517;
  assign n19519 = ~n19506 & ~n19518;
  assign n19520 = n19506 & n19518;
  assign n19521 = ~n19519 & ~n19520;
  assign n19522 = n19059 & ~n19061;
  assign n19523 = n19061 & ~n19062;
  assign n19524 = ~n19059 & ~n19062;
  assign n19525 = ~n19523 & ~n19524;
  assign n19526 = ~n19062 & ~n19522;
  assign n19527 = n19521 & ~n55368;
  assign n19528 = ~n19519 & ~n19527;
  assign n19529 = n55291 & ~n19073;
  assign n19530 = ~n55291 & ~n19074;
  assign n19531 = n19073 & ~n19074;
  assign n19532 = ~n19530 & ~n19531;
  assign n19533 = ~n19074 & ~n19529;
  assign n19534 = ~n19528 & ~n55369;
  assign n19535 = n19528 & n55369;
  assign n19536 = ~n19534 & ~n19535;
  assign n19537 = ~n19521 & n55368;
  assign n19538 = ~n19527 & ~n19537;
  assign n19539 = n11242 & n18846;
  assign n19540 = ~n53650 & n55247;
  assign n19541 = n55244 & ~n55246;
  assign n19542 = ~n2325 & n19541;
  assign n19543 = ~n53634 & n19509;
  assign n19544 = ~n19542 & ~n19543;
  assign n19545 = ~n19540 & ~n19543;
  assign n19546 = ~n19542 & n19545;
  assign n19547 = ~n19540 & n19544;
  assign n19548 = ~n18846 & n55370;
  assign n19549 = ~n11242 & n55370;
  assign n19550 = ~n19548 & ~n19549;
  assign n19551 = ~n19539 & n55370;
  assign n19552 = pi11  & ~n55371;
  assign n19553 = ~pi11  & n55371;
  assign n19554 = ~n19552 & ~n19553;
  assign n19555 = n19499 & ~n19501;
  assign n19556 = n19501 & ~n19502;
  assign n19557 = ~n19499 & ~n19502;
  assign n19558 = ~n19556 & ~n19557;
  assign n19559 = ~n19502 & ~n19555;
  assign n19560 = n12938 & n16079;
  assign n19561 = ~n53819 & n16696;
  assign n19562 = ~n53860 & n54886;
  assign n19563 = ~n53845 & n16676;
  assign n19564 = ~n19562 & ~n19563;
  assign n19565 = ~n19561 & ~n19562;
  assign n19566 = ~n19563 & n19565;
  assign n19567 = ~n19561 & n19564;
  assign n19568 = ~n19560 & n55373;
  assign n19569 = pi17  & ~n19568;
  assign n19570 = ~n19568 & ~n19569;
  assign n19571 = ~pi17  & ~n19568;
  assign n19572 = pi17  & ~n19569;
  assign n19573 = pi17  & n19568;
  assign n19574 = ~n55374 & ~n55375;
  assign n19575 = ~n19127 & n55357;
  assign n19576 = ~n19454 & ~n19575;
  assign n19577 = ~n19574 & n19576;
  assign n19578 = n19574 & ~n19576;
  assign n19579 = ~n19574 & ~n19577;
  assign n19580 = ~n19574 & ~n19576;
  assign n19581 = n19576 & ~n19577;
  assign n19582 = n19574 & n19576;
  assign n19583 = ~n55376 & ~n55377;
  assign n19584 = ~n19577 & ~n19578;
  assign n19585 = n19448 & ~n19450;
  assign n19586 = n19450 & ~n19451;
  assign n19587 = ~n19448 & ~n19451;
  assign n19588 = ~n19586 & ~n19587;
  assign n19589 = ~n19451 & ~n19585;
  assign n19590 = n19378 & ~n19380;
  assign n19591 = ~n19381 & ~n19590;
  assign n19592 = n123 & n16772;
  assign n19593 = n53444 & ~n54154;
  assign n19594 = n128 & ~n54119;
  assign n19595 = n127 & ~n54132;
  assign n19596 = ~n19594 & ~n19595;
  assign n19597 = ~n19593 & ~n19595;
  assign n19598 = ~n19594 & n19597;
  assign n19599 = ~n19593 & n19596;
  assign n19600 = ~n123 & n55380;
  assign n19601 = ~n16772 & n55380;
  assign n19602 = ~n19600 & ~n19601;
  assign n19603 = ~n19592 & n55380;
  assign n19604 = pi26  & ~n55381;
  assign n19605 = ~pi26  & n55381;
  assign n19606 = ~n19604 & ~n19605;
  assign n19607 = n19591 & ~n19606;
  assign n19608 = n19374 & ~n19376;
  assign n19609 = ~n19377 & ~n19608;
  assign n19610 = n123 & n16522;
  assign n19611 = n127 & ~n54154;
  assign n19612 = n128 & ~n54132;
  assign n19613 = n53444 & ~n54163;
  assign n19614 = ~n19612 & ~n19613;
  assign n19615 = ~n19611 & ~n19613;
  assign n19616 = ~n19612 & n19615;
  assign n19617 = ~n19611 & n19614;
  assign n19618 = ~n123 & n55382;
  assign n19619 = ~n16522 & n55382;
  assign n19620 = ~n19618 & ~n19619;
  assign n19621 = ~n19610 & n55382;
  assign n19622 = pi26  & ~n55383;
  assign n19623 = ~pi26  & n55383;
  assign n19624 = ~n19622 & ~n19623;
  assign n19625 = n19609 & ~n19624;
  assign n19626 = n19365 & n55345;
  assign n19627 = ~n19373 & ~n19626;
  assign n19628 = n123 & n17072;
  assign n19629 = n128 & ~n54154;
  assign n19630 = n53444 & ~n54183;
  assign n19631 = n127 & ~n54163;
  assign n19632 = ~n19630 & ~n19631;
  assign n19633 = ~n19629 & n19632;
  assign n19634 = ~n123 & n19633;
  assign n19635 = ~n17072 & n19633;
  assign n19636 = ~n19634 & ~n19635;
  assign n19637 = ~n19628 & n19633;
  assign n19638 = pi26  & ~n55384;
  assign n19639 = ~pi26  & n55384;
  assign n19640 = ~n19638 & ~n19639;
  assign n19641 = n19627 & ~n19640;
  assign n19642 = n19356 & n55342;
  assign n19643 = ~n19364 & ~n19642;
  assign n19644 = n123 & n17524;
  assign n19645 = n127 & ~n54183;
  assign n19646 = n53444 & ~n54194;
  assign n19647 = n128 & ~n54163;
  assign n19648 = ~n19646 & ~n19647;
  assign n19649 = ~n19645 & ~n19646;
  assign n19650 = ~n19647 & n19649;
  assign n19651 = ~n19645 & n19648;
  assign n19652 = ~n123 & n55385;
  assign n19653 = ~n17524 & n55385;
  assign n19654 = ~n19652 & ~n19653;
  assign n19655 = ~n19644 & n55385;
  assign n19656 = pi26  & ~n55386;
  assign n19657 = ~pi26  & n55386;
  assign n19658 = ~n19656 & ~n19657;
  assign n19659 = n19643 & ~n19658;
  assign n19660 = n19349 & n55339;
  assign n19661 = ~n19355 & ~n19660;
  assign n19662 = n123 & n17544;
  assign n19663 = n53444 & ~n54212;
  assign n19664 = n128 & ~n54183;
  assign n19665 = n127 & ~n54194;
  assign n19666 = ~n19664 & ~n19665;
  assign n19667 = ~n19663 & ~n19665;
  assign n19668 = ~n19664 & n19667;
  assign n19669 = ~n19663 & n19666;
  assign n19670 = ~n123 & n55387;
  assign n19671 = ~n17544 & n55387;
  assign n19672 = ~n19670 & ~n19671;
  assign n19673 = ~n19662 & n55387;
  assign n19674 = pi26  & ~n55388;
  assign n19675 = ~pi26  & n55388;
  assign n19676 = ~n19674 & ~n19675;
  assign n19677 = n19661 & ~n19676;
  assign n19678 = n19342 & n55338;
  assign n19679 = ~n19348 & ~n19678;
  assign n19680 = n123 & n17041;
  assign n19681 = n127 & ~n54212;
  assign n19682 = n128 & ~n54194;
  assign n19683 = n53444 & ~n54240;
  assign n19684 = ~n19682 & ~n19683;
  assign n19685 = ~n19681 & ~n19683;
  assign n19686 = ~n19682 & n19685;
  assign n19687 = ~n19681 & n19684;
  assign n19688 = ~n123 & n55389;
  assign n19689 = ~n17041 & n55389;
  assign n19690 = ~n19688 & ~n19689;
  assign n19691 = ~n19680 & n55389;
  assign n19692 = pi26  & ~n55390;
  assign n19693 = ~pi26  & n55390;
  assign n19694 = ~n19692 & ~n19693;
  assign n19695 = n19679 & ~n19694;
  assign n19696 = n123 & n17660;
  assign n19697 = n53444 & ~n54254;
  assign n19698 = n128 & ~n54212;
  assign n19699 = n127 & ~n54240;
  assign n19700 = ~n19698 & ~n19699;
  assign n19701 = ~n19697 & ~n19699;
  assign n19702 = ~n19698 & n19701;
  assign n19703 = ~n19697 & n19700;
  assign n19704 = ~n123 & n55391;
  assign n19705 = ~n17660 & n55391;
  assign n19706 = ~n19704 & ~n19705;
  assign n19707 = ~n19696 & n55391;
  assign n19708 = pi26  & ~n55392;
  assign n19709 = ~pi26  & n55392;
  assign n19710 = ~n19708 & ~n19709;
  assign n19711 = n19333 & n55337;
  assign n19712 = ~n55337 & ~n19341;
  assign n19713 = ~n19333 & ~n19341;
  assign n19714 = ~n19712 & ~n19713;
  assign n19715 = ~n19341 & ~n19711;
  assign n19716 = ~n19710 & ~n55393;
  assign n19717 = n123 & n17804;
  assign n19718 = n127 & ~n54254;
  assign n19719 = n128 & ~n54240;
  assign n19720 = n53444 & ~n54269;
  assign n19721 = ~n19719 & ~n19720;
  assign n19722 = ~n19718 & ~n19720;
  assign n19723 = ~n19719 & n19722;
  assign n19724 = ~n19718 & n19721;
  assign n19725 = ~n19717 & n55394;
  assign n19726 = pi26  & ~n19725;
  assign n19727 = ~n19725 & ~n19726;
  assign n19728 = ~pi26  & ~n19725;
  assign n19729 = pi26  & ~n19726;
  assign n19730 = pi26  & n19725;
  assign n19731 = ~n55395 & ~n55396;
  assign n19732 = n19326 & n55334;
  assign n19733 = ~n19332 & ~n19732;
  assign n19734 = ~n19731 & n19733;
  assign n19735 = n123 & n17939;
  assign n19736 = n128 & ~n54254;
  assign n19737 = n53444 & ~n54277;
  assign n19738 = n127 & ~n54269;
  assign n19739 = ~n19737 & ~n19738;
  assign n19740 = ~n19736 & n19739;
  assign n19741 = ~n19735 & n19740;
  assign n19742 = pi26  & ~n19741;
  assign n19743 = ~n19741 & ~n19742;
  assign n19744 = ~pi26  & ~n19741;
  assign n19745 = pi26  & ~n19742;
  assign n19746 = pi26  & n19741;
  assign n19747 = ~n55397 & ~n55398;
  assign n19748 = pi29  & ~n55328;
  assign n19749 = ~n55329 & ~n19748;
  assign n19750 = n55329 & n19748;
  assign n19751 = ~n55328 & n19308;
  assign n19752 = ~n55330 & ~n19751;
  assign n19753 = ~n19749 & ~n19750;
  assign n19754 = ~n19747 & n55399;
  assign n19755 = n123 & n18056;
  assign n19756 = n53444 & ~n54305;
  assign n19757 = n127 & ~n54277;
  assign n19758 = n128 & ~n54269;
  assign n19759 = ~n19757 & ~n19758;
  assign n19760 = ~n19756 & ~n19757;
  assign n19761 = ~n19758 & n19760;
  assign n19762 = ~n19756 & n19759;
  assign n19763 = ~n123 & n55400;
  assign n19764 = ~n18056 & n55400;
  assign n19765 = ~n19763 & ~n19764;
  assign n19766 = ~n19755 & n55400;
  assign n19767 = pi26  & ~n55401;
  assign n19768 = ~pi26  & n55401;
  assign n19769 = ~n19767 & ~n19768;
  assign n19770 = pi29  & n19288;
  assign n19771 = ~n19287 & n19770;
  assign n19772 = n19287 & ~n19770;
  assign n19773 = ~n19289 & n19293;
  assign n19774 = ~n55328 & ~n19773;
  assign n19775 = ~n19771 & ~n19772;
  assign n19776 = ~n19769 & n55402;
  assign n19777 = n123 & ~n19275;
  assign n19778 = n127 & ~n54325;
  assign n19779 = n128 & ~n54344;
  assign n19780 = ~n19778 & ~n19779;
  assign n19781 = ~n19777 & n19780;
  assign n19782 = ~n120 & ~n54325;
  assign n19783 = pi26  & ~n19782;
  assign n19784 = pi26  & ~n19781;
  assign n19785 = pi26  & ~n19784;
  assign n19786 = ~n19781 & ~n19784;
  assign n19787 = ~n19785 & ~n19786;
  assign n19788 = n19783 & ~n19787;
  assign n19789 = n19781 & n19783;
  assign n19790 = n123 & n18156;
  assign n19791 = n128 & ~n54305;
  assign n19792 = n53444 & ~n54325;
  assign n19793 = n127 & ~n54344;
  assign n19794 = ~n19792 & ~n19793;
  assign n19795 = ~n19791 & n19794;
  assign n19796 = ~n123 & n19795;
  assign n19797 = ~n18156 & n19795;
  assign n19798 = ~n19796 & ~n19797;
  assign n19799 = ~n19790 & n19795;
  assign n19800 = pi26  & ~n55404;
  assign n19801 = ~pi26  & n55404;
  assign n19802 = ~n19800 & ~n19801;
  assign n19803 = n55403 & ~n19802;
  assign n19804 = n55403 & ~n55404;
  assign n19805 = n19288 & n55405;
  assign n19806 = n123 & n18336;
  assign n19807 = n127 & ~n54305;
  assign n19808 = n128 & ~n54277;
  assign n19809 = n53444 & ~n54344;
  assign n19810 = ~n19808 & ~n19809;
  assign n19811 = ~n19807 & ~n19809;
  assign n19812 = ~n19808 & n19811;
  assign n19813 = ~n19807 & n19810;
  assign n19814 = ~n19806 & n55406;
  assign n19815 = pi26  & ~n19814;
  assign n19816 = pi26  & ~n19815;
  assign n19817 = pi26  & n19814;
  assign n19818 = ~n19814 & ~n19815;
  assign n19819 = ~pi26  & ~n19814;
  assign n19820 = ~n55407 & ~n55408;
  assign n19821 = ~n19288 & ~n55405;
  assign n19822 = n55405 & ~n19805;
  assign n19823 = ~n19288 & n55405;
  assign n19824 = n19288 & ~n19805;
  assign n19825 = n19288 & ~n55405;
  assign n19826 = ~n55409 & ~n55410;
  assign n19827 = ~n19805 & ~n19821;
  assign n19828 = ~n19820 & ~n55411;
  assign n19829 = ~n19805 & ~n19828;
  assign n19830 = n19769 & ~n55402;
  assign n19831 = ~n19776 & ~n19830;
  assign n19832 = ~n19829 & n19831;
  assign n19833 = ~n19776 & ~n19832;
  assign n19834 = n19747 & ~n55399;
  assign n19835 = ~n19747 & ~n19754;
  assign n19836 = ~n19747 & ~n55399;
  assign n19837 = n55399 & ~n19754;
  assign n19838 = n19747 & n55399;
  assign n19839 = ~n55412 & ~n55413;
  assign n19840 = ~n19754 & ~n19834;
  assign n19841 = ~n19833 & ~n55414;
  assign n19842 = ~n19754 & ~n19841;
  assign n19843 = n19731 & ~n19733;
  assign n19844 = ~n19731 & ~n19734;
  assign n19845 = ~n19731 & ~n19733;
  assign n19846 = n19733 & ~n19734;
  assign n19847 = n19731 & n19733;
  assign n19848 = ~n55415 & ~n55416;
  assign n19849 = ~n19734 & ~n19843;
  assign n19850 = ~n19842 & ~n55417;
  assign n19851 = ~n19734 & ~n19850;
  assign n19852 = n19710 & n55393;
  assign n19853 = ~n55393 & ~n19716;
  assign n19854 = n19710 & ~n55393;
  assign n19855 = ~n19710 & ~n19716;
  assign n19856 = ~n19710 & n55393;
  assign n19857 = ~n55418 & ~n55419;
  assign n19858 = ~n19716 & ~n19852;
  assign n19859 = ~n19851 & ~n55420;
  assign n19860 = ~n19716 & ~n19859;
  assign n19861 = ~n19679 & n19694;
  assign n19862 = n19679 & ~n19695;
  assign n19863 = n19679 & n19694;
  assign n19864 = ~n19694 & ~n19695;
  assign n19865 = ~n19679 & ~n19694;
  assign n19866 = ~n55421 & ~n55422;
  assign n19867 = ~n19695 & ~n19861;
  assign n19868 = ~n19860 & ~n55423;
  assign n19869 = ~n19695 & ~n19868;
  assign n19870 = ~n19661 & n19676;
  assign n19871 = n19661 & ~n19677;
  assign n19872 = n19661 & n19676;
  assign n19873 = ~n19676 & ~n19677;
  assign n19874 = ~n19661 & ~n19676;
  assign n19875 = ~n55424 & ~n55425;
  assign n19876 = ~n19677 & ~n19870;
  assign n19877 = ~n19869 & ~n55426;
  assign n19878 = ~n19677 & ~n19877;
  assign n19879 = ~n19643 & n19658;
  assign n19880 = n19643 & ~n19659;
  assign n19881 = n19643 & n19658;
  assign n19882 = ~n19658 & ~n19659;
  assign n19883 = ~n19643 & ~n19658;
  assign n19884 = ~n55427 & ~n55428;
  assign n19885 = ~n19659 & ~n19879;
  assign n19886 = ~n19878 & ~n55429;
  assign n19887 = ~n19659 & ~n19886;
  assign n19888 = ~n19627 & n19640;
  assign n19889 = n19627 & ~n19641;
  assign n19890 = n19627 & n19640;
  assign n19891 = ~n19640 & ~n19641;
  assign n19892 = ~n19627 & ~n19640;
  assign n19893 = ~n55430 & ~n55431;
  assign n19894 = ~n19641 & ~n19888;
  assign n19895 = ~n19887 & ~n55432;
  assign n19896 = ~n19641 & ~n19895;
  assign n19897 = ~n19609 & n19624;
  assign n19898 = n19609 & ~n19625;
  assign n19899 = n19609 & n19624;
  assign n19900 = ~n19624 & ~n19625;
  assign n19901 = ~n19609 & ~n19624;
  assign n19902 = ~n55433 & ~n55434;
  assign n19903 = ~n19625 & ~n19897;
  assign n19904 = ~n19896 & ~n55435;
  assign n19905 = ~n19625 & ~n19904;
  assign n19906 = ~n19591 & n19606;
  assign n19907 = n19591 & ~n19607;
  assign n19908 = n19591 & n19606;
  assign n19909 = ~n19606 & ~n19607;
  assign n19910 = ~n19591 & ~n19606;
  assign n19911 = ~n55436 & ~n55437;
  assign n19912 = ~n19607 & ~n19906;
  assign n19913 = ~n19905 & ~n55438;
  assign n19914 = ~n19607 & ~n19913;
  assign n19915 = n19400 & ~n19402;
  assign n19916 = ~n19403 & ~n19915;
  assign n19917 = ~n19914 & n19916;
  assign n19918 = n90 & n15219;
  assign n19919 = ~n54050 & n14210;
  assign n19920 = ~n54034 & n14236;
  assign n19921 = ~n54073 & n54667;
  assign n19922 = ~n19920 & ~n19921;
  assign n19923 = ~n19919 & ~n19921;
  assign n19924 = ~n19920 & n19923;
  assign n19925 = ~n19919 & n19922;
  assign n19926 = ~n19918 & n55439;
  assign n19927 = pi23  & ~n19926;
  assign n19928 = ~n19926 & ~n19927;
  assign n19929 = ~pi23  & ~n19926;
  assign n19930 = pi23  & ~n19927;
  assign n19931 = pi23  & n19926;
  assign n19932 = ~n55440 & ~n55441;
  assign n19933 = n19914 & ~n19916;
  assign n19934 = ~n19917 & ~n19933;
  assign n19935 = ~n19932 & n19934;
  assign n19936 = ~n19917 & ~n19935;
  assign n19937 = n19428 & ~n19429;
  assign n19938 = n19426 & n19428;
  assign n19939 = ~n19426 & ~n19429;
  assign n19940 = ~n19426 & ~n19428;
  assign n19941 = n19426 & ~n19428;
  assign n19942 = ~n19429 & ~n19941;
  assign n19943 = ~n55442 & ~n55443;
  assign n19944 = ~n19936 & n55444;
  assign n19945 = n19936 & ~n55444;
  assign n19946 = n14020 & n14413;
  assign n19947 = ~n53962 & n15901;
  assign n19948 = ~n53970 & n54719;
  assign n19949 = ~n53930 & n15921;
  assign n19950 = ~n19948 & ~n19949;
  assign n19951 = ~n19947 & ~n19948;
  assign n19952 = ~n19949 & n19951;
  assign n19953 = ~n19947 & n19950;
  assign n19954 = ~n19946 & n55445;
  assign n19955 = pi20  & ~n19954;
  assign n19956 = pi20  & ~n19955;
  assign n19957 = pi20  & n19954;
  assign n19958 = ~n19954 & ~n19955;
  assign n19959 = ~pi20  & ~n19954;
  assign n19960 = ~n55446 & ~n55447;
  assign n19961 = ~n19945 & ~n19960;
  assign n19962 = ~n19944 & ~n19945;
  assign n19963 = ~n19960 & n19962;
  assign n19964 = ~n19944 & ~n19963;
  assign n19965 = ~n19944 & ~n19961;
  assign n19966 = ~n55379 & ~n55448;
  assign n19967 = n55379 & n55448;
  assign n19968 = n12918 & n16079;
  assign n19969 = ~n53860 & n16676;
  assign n19970 = ~n53888 & n54886;
  assign n19971 = ~n53845 & n16696;
  assign n19972 = ~n19970 & ~n19971;
  assign n19973 = ~n19969 & ~n19970;
  assign n19974 = ~n19971 & n19973;
  assign n19975 = ~n19969 & n19972;
  assign n19976 = ~n19968 & n55449;
  assign n19977 = pi17  & ~n19976;
  assign n19978 = pi17  & ~n19977;
  assign n19979 = pi17  & n19976;
  assign n19980 = ~n19976 & ~n19977;
  assign n19981 = ~pi17  & ~n19976;
  assign n19982 = ~n55450 & ~n55451;
  assign n19983 = ~n19967 & ~n19982;
  assign n19984 = ~n19966 & ~n19967;
  assign n19985 = ~n19982 & n19984;
  assign n19986 = ~n19966 & ~n19985;
  assign n19987 = ~n19966 & ~n19983;
  assign n19988 = ~n55378 & ~n55452;
  assign n19989 = ~n19577 & ~n19988;
  assign n19990 = n19479 & ~n19480;
  assign n19991 = n19477 & n19479;
  assign n19992 = ~n19477 & ~n19480;
  assign n19993 = ~n19477 & ~n19479;
  assign n19994 = n19477 & ~n19479;
  assign n19995 = ~n19480 & ~n19994;
  assign n19996 = ~n55453 & ~n55454;
  assign n19997 = ~n19989 & n55455;
  assign n19998 = n19989 & ~n55455;
  assign n19999 = n11889 & n17265;
  assign n20000 = ~n53712 & n18588;
  assign n20001 = ~n53774 & n55041;
  assign n20002 = ~n53741 & n18556;
  assign n20003 = ~n20001 & ~n20002;
  assign n20004 = ~n20000 & ~n20001;
  assign n20005 = ~n20002 & n20004;
  assign n20006 = ~n20000 & n20003;
  assign n20007 = ~n19999 & n55456;
  assign n20008 = pi14  & ~n20007;
  assign n20009 = pi14  & ~n20008;
  assign n20010 = pi14  & n20007;
  assign n20011 = ~n20007 & ~n20008;
  assign n20012 = ~pi14  & ~n20007;
  assign n20013 = ~n55457 & ~n55458;
  assign n20014 = ~n19998 & ~n20013;
  assign n20015 = ~n19997 & ~n19998;
  assign n20016 = ~n20013 & n20015;
  assign n20017 = ~n19997 & ~n20016;
  assign n20018 = ~n19997 & ~n20014;
  assign n20019 = ~n55372 & ~n55459;
  assign n20020 = n55372 & n55459;
  assign n20021 = n11286 & n18846;
  assign n20022 = ~n53650 & n19509;
  assign n20023 = ~n53657 & n55247;
  assign n20024 = ~n53634 & n19541;
  assign n20025 = ~n20023 & ~n20024;
  assign n20026 = ~n20022 & ~n20023;
  assign n20027 = ~n20024 & n20026;
  assign n20028 = ~n20022 & n20025;
  assign n20029 = ~n20021 & n55460;
  assign n20030 = pi11  & ~n20029;
  assign n20031 = pi11  & ~n20030;
  assign n20032 = pi11  & n20029;
  assign n20033 = ~n20029 & ~n20030;
  assign n20034 = ~pi11  & ~n20029;
  assign n20035 = ~n55461 & ~n55462;
  assign n20036 = ~n20020 & ~n20035;
  assign n20037 = ~n20019 & ~n20020;
  assign n20038 = ~n20035 & n20037;
  assign n20039 = ~n20019 & ~n20038;
  assign n20040 = ~n20019 & ~n20036;
  assign n20041 = ~n19554 & ~n55463;
  assign n20042 = n19554 & n55463;
  assign n20043 = n55297 & n55366;
  assign n20044 = ~n55366 & ~n19505;
  assign n20045 = n55297 & ~n55366;
  assign n20046 = ~n55297 & ~n19505;
  assign n20047 = ~n55297 & n55366;
  assign n20048 = ~n55464 & ~n55465;
  assign n20049 = ~n19505 & ~n20043;
  assign n20050 = ~n20042 & ~n55466;
  assign n20051 = ~n20041 & ~n20042;
  assign n20052 = ~n55466 & n20051;
  assign n20053 = ~n20041 & ~n20052;
  assign n20054 = ~n20041 & ~n20050;
  assign n20055 = n19538 & ~n55467;
  assign n20056 = n55466 & ~n20051;
  assign n20057 = n20051 & ~n20052;
  assign n20058 = ~n55466 & ~n20052;
  assign n20059 = ~n20057 & ~n20058;
  assign n20060 = ~n20052 & ~n20056;
  assign n20061 = pi5  & ~pi6 ;
  assign n20062 = ~pi5  & pi6 ;
  assign n20063 = ~pi5  & ~pi6 ;
  assign n20064 = pi5  & pi6 ;
  assign n20065 = ~n20063 & ~n20064;
  assign n20066 = ~n20061 & ~n20062;
  assign n20067 = pi6  & ~pi7 ;
  assign n20068 = ~pi6  & pi7 ;
  assign n20069 = ~pi6  & ~pi7 ;
  assign n20070 = pi6  & pi7 ;
  assign n20071 = ~n20069 & ~n20070;
  assign n20072 = ~n20067 & ~n20068;
  assign n20073 = ~n55469 & ~n55470;
  assign n20074 = pi7  & ~pi8 ;
  assign n20075 = ~pi7  & pi8 ;
  assign n20076 = ~pi7  & ~pi8 ;
  assign n20077 = pi7  & pi8 ;
  assign n20078 = ~n20076 & ~n20077;
  assign n20079 = ~n20074 & ~n20075;
  assign n20080 = ~n55469 & n55471;
  assign n20081 = ~n55470 & n20080;
  assign n20082 = ~n55470 & n55471;
  assign n20083 = ~n55469 & n20082;
  assign n20084 = n20073 & n55471;
  assign n20085 = n55469 & n55471;
  assign n20086 = ~n10547 & n20085;
  assign n20087 = ~n55472 & ~n20086;
  assign n20088 = ~n2325 & n55472;
  assign n20089 = ~n10551 & ~n20088;
  assign n20090 = ~n20085 & ~n20088;
  assign n20091 = ~n20089 & ~n20090;
  assign n20092 = ~n2325 & ~n20087;
  assign n20093 = pi8  & ~n55473;
  assign n20094 = ~pi8  & n55473;
  assign n20095 = ~n20093 & ~n20094;
  assign n20096 = n55378 & n55452;
  assign n20097 = ~n19988 & ~n20096;
  assign n20098 = n11913 & n17265;
  assign n20099 = ~n53774 & n18556;
  assign n20100 = ~n53799 & n55041;
  assign n20101 = ~n53741 & n18588;
  assign n20102 = ~n20100 & ~n20101;
  assign n20103 = ~n20099 & ~n20100;
  assign n20104 = ~n20101 & n20103;
  assign n20105 = ~n20099 & n20102;
  assign n20106 = ~n17265 & n55474;
  assign n20107 = ~n11913 & n55474;
  assign n20108 = ~n20106 & ~n20107;
  assign n20109 = ~n20098 & n55474;
  assign n20110 = pi14  & ~n55475;
  assign n20111 = ~pi14  & n55475;
  assign n20112 = ~n20110 & ~n20111;
  assign n20113 = n20097 & ~n20112;
  assign n20114 = ~n20097 & n20112;
  assign n20115 = ~n20113 & ~n20114;
  assign n20116 = n19982 & ~n19984;
  assign n20117 = n19984 & ~n19985;
  assign n20118 = ~n19982 & ~n19985;
  assign n20119 = ~n20117 & ~n20118;
  assign n20120 = ~n19985 & ~n20116;
  assign n20121 = n90 & n16138;
  assign n20122 = ~n54098 & n54667;
  assign n20123 = ~n54050 & n14236;
  assign n20124 = ~n54073 & n14210;
  assign n20125 = ~n20123 & ~n20124;
  assign n20126 = ~n20122 & ~n20124;
  assign n20127 = ~n20123 & n20126;
  assign n20128 = ~n20122 & n20125;
  assign n20129 = ~n20121 & n55477;
  assign n20130 = pi23  & ~n20129;
  assign n20131 = ~n20129 & ~n20130;
  assign n20132 = ~pi23  & ~n20129;
  assign n20133 = pi23  & ~n20130;
  assign n20134 = pi23  & n20129;
  assign n20135 = ~n55478 & ~n55479;
  assign n20136 = n19905 & n55438;
  assign n20137 = ~n19905 & ~n19913;
  assign n20138 = ~n55438 & ~n19913;
  assign n20139 = ~n20137 & ~n20138;
  assign n20140 = ~n19913 & ~n20136;
  assign n20141 = ~n20135 & ~n55480;
  assign n20142 = n90 & n15779;
  assign n20143 = ~n54098 & n14210;
  assign n20144 = ~n54119 & n54667;
  assign n20145 = ~n54073 & n14236;
  assign n20146 = ~n20144 & ~n20145;
  assign n20147 = ~n20143 & ~n20144;
  assign n20148 = ~n20145 & n20147;
  assign n20149 = ~n20143 & ~n20145;
  assign n20150 = ~n20144 & n20149;
  assign n20151 = ~n20143 & n20146;
  assign n20152 = ~n20142 & n55481;
  assign n20153 = pi23  & ~n20152;
  assign n20154 = ~n20152 & ~n20153;
  assign n20155 = ~pi23  & ~n20152;
  assign n20156 = pi23  & ~n20153;
  assign n20157 = pi23  & n20152;
  assign n20158 = ~n55482 & ~n55483;
  assign n20159 = n19896 & n55435;
  assign n20160 = ~n19896 & ~n19904;
  assign n20161 = ~n55435 & ~n19904;
  assign n20162 = ~n20160 & ~n20161;
  assign n20163 = ~n19904 & ~n20159;
  assign n20164 = ~n20158 & ~n55484;
  assign n20165 = n90 & n16547;
  assign n20166 = ~n54119 & n14210;
  assign n20167 = ~n54098 & n14236;
  assign n20168 = ~n54132 & n54667;
  assign n20169 = ~n20167 & ~n20168;
  assign n20170 = ~n20166 & ~n20168;
  assign n20171 = ~n20167 & n20170;
  assign n20172 = ~n20166 & n20169;
  assign n20173 = ~n20165 & n55485;
  assign n20174 = pi23  & ~n20173;
  assign n20175 = ~n20173 & ~n20174;
  assign n20176 = ~pi23  & ~n20173;
  assign n20177 = pi23  & ~n20174;
  assign n20178 = pi23  & n20173;
  assign n20179 = ~n55486 & ~n55487;
  assign n20180 = n19887 & n55432;
  assign n20181 = ~n19887 & ~n19895;
  assign n20182 = ~n19887 & n55432;
  assign n20183 = ~n55432 & ~n19895;
  assign n20184 = n19887 & ~n55432;
  assign n20185 = ~n55488 & ~n55489;
  assign n20186 = ~n19895 & ~n20180;
  assign n20187 = ~n20179 & ~n55490;
  assign n20188 = n90 & n16772;
  assign n20189 = ~n54154 & n54667;
  assign n20190 = ~n54119 & n14236;
  assign n20191 = ~n54132 & n14210;
  assign n20192 = ~n20190 & ~n20191;
  assign n20193 = ~n20189 & ~n20191;
  assign n20194 = ~n20190 & n20193;
  assign n20195 = ~n20189 & n20192;
  assign n20196 = ~n20188 & n55491;
  assign n20197 = pi23  & ~n20196;
  assign n20198 = ~n20196 & ~n20197;
  assign n20199 = ~pi23  & ~n20196;
  assign n20200 = pi23  & ~n20197;
  assign n20201 = pi23  & n20196;
  assign n20202 = ~n55492 & ~n55493;
  assign n20203 = n19878 & n55429;
  assign n20204 = ~n19878 & ~n19886;
  assign n20205 = ~n19878 & n55429;
  assign n20206 = ~n55429 & ~n19886;
  assign n20207 = n19878 & ~n55429;
  assign n20208 = ~n55494 & ~n55495;
  assign n20209 = ~n19886 & ~n20203;
  assign n20210 = ~n20202 & ~n55496;
  assign n20211 = n90 & n16522;
  assign n20212 = ~n54154 & n14210;
  assign n20213 = ~n54132 & n14236;
  assign n20214 = ~n54163 & n54667;
  assign n20215 = ~n20213 & ~n20214;
  assign n20216 = ~n20212 & ~n20214;
  assign n20217 = ~n20213 & n20216;
  assign n20218 = ~n20212 & n20215;
  assign n20219 = ~n20211 & n55497;
  assign n20220 = pi23  & ~n20219;
  assign n20221 = ~n20219 & ~n20220;
  assign n20222 = ~pi23  & ~n20219;
  assign n20223 = pi23  & ~n20220;
  assign n20224 = pi23  & n20219;
  assign n20225 = ~n55498 & ~n55499;
  assign n20226 = n19869 & n55426;
  assign n20227 = ~n19869 & ~n19877;
  assign n20228 = ~n55426 & ~n19877;
  assign n20229 = ~n20227 & ~n20228;
  assign n20230 = ~n19877 & ~n20226;
  assign n20231 = ~n20225 & ~n55500;
  assign n20232 = n90 & n17072;
  assign n20233 = ~n54154 & n14236;
  assign n20234 = ~n54183 & n54667;
  assign n20235 = ~n54163 & n14210;
  assign n20236 = ~n20234 & ~n20235;
  assign n20237 = ~n20233 & n20236;
  assign n20238 = ~n20232 & n20237;
  assign n20239 = pi23  & ~n20238;
  assign n20240 = ~n20238 & ~n20239;
  assign n20241 = ~pi23  & ~n20238;
  assign n20242 = pi23  & ~n20239;
  assign n20243 = pi23  & n20238;
  assign n20244 = ~n55501 & ~n55502;
  assign n20245 = n19860 & n55423;
  assign n20246 = ~n19860 & ~n19868;
  assign n20247 = ~n55423 & ~n19868;
  assign n20248 = ~n20246 & ~n20247;
  assign n20249 = ~n19868 & ~n20245;
  assign n20250 = ~n20244 & ~n55503;
  assign n20251 = n90 & n17524;
  assign n20252 = ~n54183 & n14210;
  assign n20253 = ~n54194 & n54667;
  assign n20254 = ~n54163 & n14236;
  assign n20255 = ~n20253 & ~n20254;
  assign n20256 = ~n20252 & ~n20253;
  assign n20257 = ~n20254 & n20256;
  assign n20258 = ~n20252 & n20255;
  assign n20259 = ~n20251 & n55504;
  assign n20260 = pi23  & ~n20259;
  assign n20261 = ~n20259 & ~n20260;
  assign n20262 = ~pi23  & ~n20259;
  assign n20263 = pi23  & ~n20260;
  assign n20264 = pi23  & n20259;
  assign n20265 = ~n55505 & ~n55506;
  assign n20266 = n19851 & n55420;
  assign n20267 = ~n19851 & ~n19859;
  assign n20268 = ~n19851 & n55420;
  assign n20269 = ~n55420 & ~n19859;
  assign n20270 = n19851 & ~n55420;
  assign n20271 = ~n55507 & ~n55508;
  assign n20272 = ~n19859 & ~n20266;
  assign n20273 = ~n20265 & ~n55509;
  assign n20274 = n19842 & n55417;
  assign n20275 = ~n19850 & ~n20274;
  assign n20276 = n90 & n17544;
  assign n20277 = ~n54212 & n54667;
  assign n20278 = ~n54183 & n14236;
  assign n20279 = ~n54194 & n14210;
  assign n20280 = ~n20278 & ~n20279;
  assign n20281 = ~n20277 & ~n20279;
  assign n20282 = ~n20278 & n20281;
  assign n20283 = ~n20277 & n20280;
  assign n20284 = ~n90 & n55510;
  assign n20285 = ~n17544 & n55510;
  assign n20286 = ~n20284 & ~n20285;
  assign n20287 = ~n20276 & n55510;
  assign n20288 = pi23  & ~n55511;
  assign n20289 = ~pi23  & n55511;
  assign n20290 = ~n20288 & ~n20289;
  assign n20291 = n20275 & ~n20290;
  assign n20292 = n19833 & n55414;
  assign n20293 = ~n19841 & ~n20292;
  assign n20294 = n90 & n17041;
  assign n20295 = ~n54212 & n14210;
  assign n20296 = ~n54194 & n14236;
  assign n20297 = ~n54240 & n54667;
  assign n20298 = ~n20296 & ~n20297;
  assign n20299 = ~n20295 & ~n20297;
  assign n20300 = ~n20296 & n20299;
  assign n20301 = ~n20295 & n20298;
  assign n20302 = ~n90 & n55512;
  assign n20303 = ~n17041 & n55512;
  assign n20304 = ~n20302 & ~n20303;
  assign n20305 = ~n20294 & n55512;
  assign n20306 = pi23  & ~n55513;
  assign n20307 = ~pi23  & n55513;
  assign n20308 = ~n20306 & ~n20307;
  assign n20309 = n20293 & ~n20308;
  assign n20310 = n90 & n17660;
  assign n20311 = ~n54254 & n54667;
  assign n20312 = ~n54212 & n14236;
  assign n20313 = ~n54240 & n14210;
  assign n20314 = ~n20312 & ~n20313;
  assign n20315 = ~n20311 & ~n20313;
  assign n20316 = ~n20312 & n20315;
  assign n20317 = ~n20311 & n20314;
  assign n20318 = ~n20310 & n55514;
  assign n20319 = pi23  & ~n20318;
  assign n20320 = ~n20318 & ~n20319;
  assign n20321 = ~pi23  & ~n20318;
  assign n20322 = pi23  & ~n20319;
  assign n20323 = pi23  & n20318;
  assign n20324 = ~n55515 & ~n55516;
  assign n20325 = n19829 & ~n19831;
  assign n20326 = ~n19832 & ~n20325;
  assign n20327 = ~n20324 & n20326;
  assign n20328 = n90 & n17804;
  assign n20329 = ~n54254 & n14210;
  assign n20330 = ~n54240 & n14236;
  assign n20331 = ~n54269 & n54667;
  assign n20332 = ~n20330 & ~n20331;
  assign n20333 = ~n20329 & ~n20331;
  assign n20334 = ~n20330 & n20333;
  assign n20335 = ~n20329 & n20332;
  assign n20336 = ~n90 & n55517;
  assign n20337 = ~n17804 & n55517;
  assign n20338 = ~n20336 & ~n20337;
  assign n20339 = ~n20328 & n55517;
  assign n20340 = pi23  & ~n55518;
  assign n20341 = ~pi23  & n55518;
  assign n20342 = ~n20340 & ~n20341;
  assign n20343 = n19820 & n55411;
  assign n20344 = ~n55411 & ~n19828;
  assign n20345 = ~n19820 & ~n19828;
  assign n20346 = ~n20344 & ~n20345;
  assign n20347 = ~n19828 & ~n20343;
  assign n20348 = ~n20342 & ~n55519;
  assign n20349 = n90 & n17939;
  assign n20350 = ~n54254 & n14236;
  assign n20351 = ~n54277 & n54667;
  assign n20352 = ~n54269 & n14210;
  assign n20353 = ~n20351 & ~n20352;
  assign n20354 = ~n20350 & n20353;
  assign n20355 = ~n20349 & n20354;
  assign n20356 = pi23  & ~n20355;
  assign n20357 = ~n20355 & ~n20356;
  assign n20358 = ~pi23  & ~n20355;
  assign n20359 = pi23  & ~n20356;
  assign n20360 = pi23  & n20355;
  assign n20361 = ~n55520 & ~n55521;
  assign n20362 = pi26  & ~n55403;
  assign n20363 = ~n55404 & ~n20362;
  assign n20364 = n55404 & n20362;
  assign n20365 = ~n55403 & n19802;
  assign n20366 = ~n55405 & ~n20365;
  assign n20367 = ~n20363 & ~n20364;
  assign n20368 = ~n20361 & n55522;
  assign n20369 = n90 & n18056;
  assign n20370 = ~n54305 & n54667;
  assign n20371 = ~n54277 & n14210;
  assign n20372 = ~n54269 & n14236;
  assign n20373 = ~n20371 & ~n20372;
  assign n20374 = ~n20370 & ~n20371;
  assign n20375 = ~n20372 & n20374;
  assign n20376 = ~n20370 & n20373;
  assign n20377 = ~n90 & n55523;
  assign n20378 = ~n18056 & n55523;
  assign n20379 = ~n20377 & ~n20378;
  assign n20380 = ~n20369 & n55523;
  assign n20381 = pi23  & ~n55524;
  assign n20382 = ~pi23  & n55524;
  assign n20383 = ~n20381 & ~n20382;
  assign n20384 = pi26  & n19782;
  assign n20385 = ~n19781 & n20384;
  assign n20386 = n19781 & ~n20384;
  assign n20387 = ~n19783 & n19787;
  assign n20388 = ~n55403 & ~n20387;
  assign n20389 = ~n20385 & ~n20386;
  assign n20390 = ~n20383 & n55525;
  assign n20391 = n90 & ~n19275;
  assign n20392 = ~n54325 & n14210;
  assign n20393 = ~n54344 & n14236;
  assign n20394 = ~n20392 & ~n20393;
  assign n20395 = ~n20391 & n20394;
  assign n20396 = n53441 & ~n54325;
  assign n20397 = pi23  & ~n20396;
  assign n20398 = pi23  & ~n20395;
  assign n20399 = pi23  & ~n20398;
  assign n20400 = ~n20395 & ~n20398;
  assign n20401 = ~n20399 & ~n20400;
  assign n20402 = n20397 & ~n20401;
  assign n20403 = n20395 & n20397;
  assign n20404 = n90 & n18156;
  assign n20405 = ~n54305 & n14236;
  assign n20406 = ~n54325 & n54667;
  assign n20407 = ~n54344 & n14210;
  assign n20408 = ~n20406 & ~n20407;
  assign n20409 = ~n20405 & n20408;
  assign n20410 = ~n90 & n20409;
  assign n20411 = ~n18156 & n20409;
  assign n20412 = ~n20410 & ~n20411;
  assign n20413 = ~n20404 & n20409;
  assign n20414 = pi23  & ~n55527;
  assign n20415 = ~pi23  & n55527;
  assign n20416 = ~n20414 & ~n20415;
  assign n20417 = n55526 & ~n20416;
  assign n20418 = n55526 & ~n55527;
  assign n20419 = n19782 & n55528;
  assign n20420 = n90 & n18336;
  assign n20421 = ~n54305 & n14210;
  assign n20422 = ~n54277 & n14236;
  assign n20423 = ~n54344 & n54667;
  assign n20424 = ~n20422 & ~n20423;
  assign n20425 = ~n20421 & ~n20423;
  assign n20426 = ~n20422 & n20425;
  assign n20427 = ~n20421 & n20424;
  assign n20428 = ~n20420 & n55529;
  assign n20429 = pi23  & ~n20428;
  assign n20430 = pi23  & ~n20429;
  assign n20431 = pi23  & n20428;
  assign n20432 = ~n20428 & ~n20429;
  assign n20433 = ~pi23  & ~n20428;
  assign n20434 = ~n55530 & ~n55531;
  assign n20435 = ~n19782 & ~n55528;
  assign n20436 = n55528 & ~n20419;
  assign n20437 = ~n19782 & n55528;
  assign n20438 = n19782 & ~n20419;
  assign n20439 = n19782 & ~n55528;
  assign n20440 = ~n55532 & ~n55533;
  assign n20441 = ~n20419 & ~n20435;
  assign n20442 = ~n20434 & ~n55534;
  assign n20443 = ~n20419 & ~n20442;
  assign n20444 = n20383 & ~n55525;
  assign n20445 = ~n20390 & ~n20444;
  assign n20446 = ~n20443 & n20445;
  assign n20447 = ~n20390 & ~n20446;
  assign n20448 = n20361 & ~n55522;
  assign n20449 = ~n20361 & ~n20368;
  assign n20450 = ~n20361 & ~n55522;
  assign n20451 = n55522 & ~n20368;
  assign n20452 = n20361 & n55522;
  assign n20453 = ~n55535 & ~n55536;
  assign n20454 = ~n20368 & ~n20448;
  assign n20455 = ~n20447 & ~n55537;
  assign n20456 = ~n20368 & ~n20455;
  assign n20457 = n20342 & n55519;
  assign n20458 = ~n20348 & ~n20457;
  assign n20459 = ~n20456 & n20458;
  assign n20460 = ~n20348 & ~n20459;
  assign n20461 = n20324 & ~n20326;
  assign n20462 = ~n20324 & ~n20327;
  assign n20463 = ~n20324 & ~n20326;
  assign n20464 = n20326 & ~n20327;
  assign n20465 = n20324 & n20326;
  assign n20466 = ~n55538 & ~n55539;
  assign n20467 = ~n20327 & ~n20461;
  assign n20468 = ~n20460 & ~n55540;
  assign n20469 = ~n20327 & ~n20468;
  assign n20470 = ~n20293 & n20308;
  assign n20471 = n20293 & ~n20309;
  assign n20472 = n20293 & n20308;
  assign n20473 = ~n20308 & ~n20309;
  assign n20474 = ~n20293 & ~n20308;
  assign n20475 = ~n55541 & ~n55542;
  assign n20476 = ~n20309 & ~n20470;
  assign n20477 = ~n20469 & ~n55543;
  assign n20478 = ~n20309 & ~n20477;
  assign n20479 = ~n20275 & n20290;
  assign n20480 = ~n20291 & ~n20479;
  assign n20481 = ~n20478 & n20480;
  assign n20482 = ~n20291 & ~n20481;
  assign n20483 = n20265 & n55509;
  assign n20484 = ~n20265 & ~n20273;
  assign n20485 = ~n55509 & ~n20273;
  assign n20486 = ~n20484 & ~n20485;
  assign n20487 = ~n20273 & ~n20483;
  assign n20488 = ~n20482 & ~n55544;
  assign n20489 = ~n20273 & ~n20488;
  assign n20490 = n20244 & n55503;
  assign n20491 = ~n20244 & ~n20250;
  assign n20492 = ~n20244 & n55503;
  assign n20493 = ~n55503 & ~n20250;
  assign n20494 = n20244 & ~n55503;
  assign n20495 = ~n55545 & ~n55546;
  assign n20496 = ~n20250 & ~n20490;
  assign n20497 = ~n20489 & ~n55547;
  assign n20498 = ~n20250 & ~n20497;
  assign n20499 = n20225 & n55500;
  assign n20500 = ~n20225 & ~n20231;
  assign n20501 = ~n20225 & n55500;
  assign n20502 = ~n55500 & ~n20231;
  assign n20503 = n20225 & ~n55500;
  assign n20504 = ~n55548 & ~n55549;
  assign n20505 = ~n20231 & ~n20499;
  assign n20506 = ~n20498 & ~n55550;
  assign n20507 = ~n20231 & ~n20506;
  assign n20508 = n20202 & n55496;
  assign n20509 = ~n20202 & ~n20210;
  assign n20510 = ~n55496 & ~n20210;
  assign n20511 = ~n20509 & ~n20510;
  assign n20512 = ~n20210 & ~n20508;
  assign n20513 = ~n20507 & ~n55551;
  assign n20514 = ~n20210 & ~n20513;
  assign n20515 = n20179 & n55490;
  assign n20516 = ~n20179 & ~n20187;
  assign n20517 = ~n55490 & ~n20187;
  assign n20518 = ~n20516 & ~n20517;
  assign n20519 = ~n20187 & ~n20515;
  assign n20520 = ~n20514 & ~n55552;
  assign n20521 = ~n20187 & ~n20520;
  assign n20522 = n20158 & n55484;
  assign n20523 = ~n20158 & ~n20164;
  assign n20524 = ~n20158 & n55484;
  assign n20525 = ~n55484 & ~n20164;
  assign n20526 = n20158 & ~n55484;
  assign n20527 = ~n55553 & ~n55554;
  assign n20528 = ~n20164 & ~n20522;
  assign n20529 = ~n20521 & ~n55555;
  assign n20530 = ~n20164 & ~n20529;
  assign n20531 = n20135 & n55480;
  assign n20532 = ~n20135 & ~n20141;
  assign n20533 = ~n20135 & n55480;
  assign n20534 = ~n55480 & ~n20141;
  assign n20535 = n20135 & ~n55480;
  assign n20536 = ~n55556 & ~n55557;
  assign n20537 = ~n20141 & ~n20531;
  assign n20538 = ~n20530 & ~n55558;
  assign n20539 = ~n20141 & ~n20538;
  assign n20540 = n19932 & ~n19934;
  assign n20541 = ~n19935 & ~n20540;
  assign n20542 = ~n20539 & n20541;
  assign n20543 = n14413 & n14708;
  assign n20544 = ~n54005 & n54719;
  assign n20545 = ~n53970 & n15901;
  assign n20546 = ~n53962 & n15921;
  assign n20547 = ~n20545 & ~n20546;
  assign n20548 = ~n20544 & ~n20545;
  assign n20549 = ~n20546 & n20548;
  assign n20550 = ~n20544 & n20547;
  assign n20551 = ~n20543 & n55559;
  assign n20552 = pi20  & ~n20551;
  assign n20553 = ~n20551 & ~n20552;
  assign n20554 = ~pi20  & ~n20551;
  assign n20555 = pi20  & ~n20552;
  assign n20556 = pi20  & n20551;
  assign n20557 = ~n55560 & ~n55561;
  assign n20558 = n20539 & ~n20541;
  assign n20559 = ~n20542 & ~n20558;
  assign n20560 = ~n20557 & n20559;
  assign n20561 = ~n20542 & ~n20560;
  assign n20562 = n19960 & ~n19962;
  assign n20563 = n19962 & ~n19963;
  assign n20564 = ~n19960 & ~n19963;
  assign n20565 = ~n20563 & ~n20564;
  assign n20566 = ~n19963 & ~n20562;
  assign n20567 = ~n20561 & ~n55562;
  assign n20568 = n20561 & n55562;
  assign n20569 = n13336 & n16079;
  assign n20570 = ~n53888 & n16676;
  assign n20571 = ~n53907 & n54886;
  assign n20572 = ~n53860 & n16696;
  assign n20573 = ~n20571 & ~n20572;
  assign n20574 = ~n20570 & ~n20571;
  assign n20575 = ~n20572 & n20574;
  assign n20576 = ~n20570 & n20573;
  assign n20577 = ~n20569 & n55563;
  assign n20578 = pi17  & ~n20577;
  assign n20579 = pi17  & ~n20578;
  assign n20580 = pi17  & n20577;
  assign n20581 = ~n20577 & ~n20578;
  assign n20582 = ~pi17  & ~n20577;
  assign n20583 = ~n55564 & ~n55565;
  assign n20584 = ~n20568 & ~n20583;
  assign n20585 = ~n20567 & ~n20568;
  assign n20586 = ~n20583 & n20585;
  assign n20587 = ~n20567 & ~n20586;
  assign n20588 = ~n20567 & ~n20584;
  assign n20589 = ~n55476 & ~n55566;
  assign n20590 = n55476 & n55566;
  assign n20591 = n12690 & n17265;
  assign n20592 = ~n53774 & n18588;
  assign n20593 = ~n53819 & n55041;
  assign n20594 = ~n53799 & n18556;
  assign n20595 = ~n20593 & ~n20594;
  assign n20596 = ~n20592 & ~n20593;
  assign n20597 = ~n20594 & n20596;
  assign n20598 = ~n20592 & n20595;
  assign n20599 = ~n20591 & n55567;
  assign n20600 = pi14  & ~n20599;
  assign n20601 = pi14  & ~n20600;
  assign n20602 = pi14  & n20599;
  assign n20603 = ~n20599 & ~n20600;
  assign n20604 = ~pi14  & ~n20599;
  assign n20605 = ~n55568 & ~n55569;
  assign n20606 = ~n20590 & ~n20605;
  assign n20607 = ~n20589 & ~n20590;
  assign n20608 = ~n20605 & n20607;
  assign n20609 = ~n20589 & ~n20608;
  assign n20610 = ~n20589 & ~n20606;
  assign n20611 = n20115 & ~n55570;
  assign n20612 = ~n20113 & ~n20611;
  assign n20613 = n20013 & ~n20015;
  assign n20614 = n20015 & ~n20016;
  assign n20615 = ~n20013 & ~n20016;
  assign n20616 = ~n20614 & ~n20615;
  assign n20617 = ~n20016 & ~n20613;
  assign n20618 = ~n20612 & ~n55571;
  assign n20619 = n20612 & n55571;
  assign n20620 = n11213 & n18846;
  assign n20621 = ~n53650 & n19541;
  assign n20622 = ~n53685 & n55247;
  assign n20623 = ~n53657 & n19509;
  assign n20624 = ~n20622 & ~n20623;
  assign n20625 = ~n20621 & n20624;
  assign n20626 = ~n20620 & n20625;
  assign n20627 = pi11  & ~n20626;
  assign n20628 = pi11  & ~n20627;
  assign n20629 = pi11  & n20626;
  assign n20630 = ~n20626 & ~n20627;
  assign n20631 = ~pi11  & ~n20626;
  assign n20632 = ~n55572 & ~n55573;
  assign n20633 = ~n20619 & ~n20632;
  assign n20634 = ~n20618 & ~n20619;
  assign n20635 = ~n20632 & n20634;
  assign n20636 = ~n20618 & ~n20635;
  assign n20637 = ~n20618 & ~n20633;
  assign n20638 = ~n20095 & ~n55574;
  assign n20639 = n20095 & n55574;
  assign n20640 = n20035 & ~n20037;
  assign n20641 = n20037 & ~n20038;
  assign n20642 = ~n20035 & ~n20038;
  assign n20643 = ~n20641 & ~n20642;
  assign n20644 = ~n20038 & ~n20640;
  assign n20645 = ~n20639 & ~n55575;
  assign n20646 = ~n20638 & ~n20639;
  assign n20647 = ~n55575 & n20646;
  assign n20648 = ~n20638 & ~n20647;
  assign n20649 = ~n20638 & ~n20645;
  assign n20650 = ~n55468 & ~n55576;
  assign n20651 = n55468 & n55576;
  assign n20652 = ~n20650 & ~n20651;
  assign n20653 = n11380 & n18846;
  assign n20654 = ~n53685 & n19509;
  assign n20655 = ~n53657 & n19541;
  assign n20656 = ~n53712 & n55247;
  assign n20657 = ~n20655 & ~n20656;
  assign n20658 = ~n20654 & ~n20656;
  assign n20659 = ~n20655 & n20658;
  assign n20660 = ~n20654 & n20657;
  assign n20661 = ~n18846 & n55577;
  assign n20662 = ~n11380 & n55577;
  assign n20663 = ~n20661 & ~n20662;
  assign n20664 = ~n20653 & n55577;
  assign n20665 = pi11  & ~n55578;
  assign n20666 = ~pi11  & n55578;
  assign n20667 = ~n20665 & ~n20666;
  assign n20668 = n20605 & ~n20607;
  assign n20669 = n20607 & ~n20608;
  assign n20670 = ~n20605 & ~n20608;
  assign n20671 = ~n20669 & ~n20670;
  assign n20672 = ~n20608 & ~n20668;
  assign n20673 = n20530 & n55558;
  assign n20674 = ~n20538 & ~n20673;
  assign n20675 = n14413 & n14688;
  assign n20676 = ~n54005 & n15901;
  assign n20677 = ~n54034 & n54719;
  assign n20678 = ~n53970 & n15921;
  assign n20679 = ~n20677 & ~n20678;
  assign n20680 = ~n20676 & ~n20677;
  assign n20681 = ~n20678 & n20680;
  assign n20682 = ~n20676 & n20679;
  assign n20683 = ~n14413 & n55580;
  assign n20684 = ~n14688 & n55580;
  assign n20685 = ~n20683 & ~n20684;
  assign n20686 = ~n20675 & n55580;
  assign n20687 = pi20  & ~n55581;
  assign n20688 = ~pi20  & n55581;
  assign n20689 = ~n20687 & ~n20688;
  assign n20690 = n20674 & ~n20689;
  assign n20691 = n20521 & n55555;
  assign n20692 = ~n20529 & ~n20691;
  assign n20693 = n14413 & n15195;
  assign n20694 = ~n54050 & n54719;
  assign n20695 = ~n54005 & n15921;
  assign n20696 = ~n54034 & n15901;
  assign n20697 = ~n20695 & ~n20696;
  assign n20698 = ~n20694 & ~n20696;
  assign n20699 = ~n20695 & n20698;
  assign n20700 = ~n20694 & n20697;
  assign n20701 = ~n14413 & n55582;
  assign n20702 = ~n15195 & n55582;
  assign n20703 = ~n20701 & ~n20702;
  assign n20704 = ~n20693 & n55582;
  assign n20705 = pi20  & ~n55583;
  assign n20706 = ~pi20  & n55583;
  assign n20707 = ~n20705 & ~n20706;
  assign n20708 = n20692 & ~n20707;
  assign n20709 = n20514 & n55552;
  assign n20710 = ~n20520 & ~n20709;
  assign n20711 = n14413 & n15219;
  assign n20712 = ~n54050 & n15901;
  assign n20713 = ~n54034 & n15921;
  assign n20714 = ~n54073 & n54719;
  assign n20715 = ~n20713 & ~n20714;
  assign n20716 = ~n20712 & ~n20714;
  assign n20717 = ~n20713 & n20716;
  assign n20718 = ~n20712 & n20715;
  assign n20719 = ~n14413 & n55584;
  assign n20720 = ~n15219 & n55584;
  assign n20721 = ~n20719 & ~n20720;
  assign n20722 = ~n20711 & n55584;
  assign n20723 = pi20  & ~n55585;
  assign n20724 = ~pi20  & n55585;
  assign n20725 = ~n20723 & ~n20724;
  assign n20726 = n20710 & ~n20725;
  assign n20727 = n20507 & n55551;
  assign n20728 = ~n20513 & ~n20727;
  assign n20729 = n14413 & n16138;
  assign n20730 = ~n54098 & n54719;
  assign n20731 = ~n54050 & n15921;
  assign n20732 = ~n54073 & n15901;
  assign n20733 = ~n20731 & ~n20732;
  assign n20734 = ~n20730 & ~n20732;
  assign n20735 = ~n20731 & n20734;
  assign n20736 = ~n20730 & n20733;
  assign n20737 = ~n14413 & n55586;
  assign n20738 = ~n16138 & n55586;
  assign n20739 = ~n20737 & ~n20738;
  assign n20740 = ~n20729 & n55586;
  assign n20741 = pi20  & ~n55587;
  assign n20742 = ~pi20  & n55587;
  assign n20743 = ~n20741 & ~n20742;
  assign n20744 = n20728 & ~n20743;
  assign n20745 = n20498 & n55550;
  assign n20746 = ~n20506 & ~n20745;
  assign n20747 = n14413 & n15779;
  assign n20748 = ~n54098 & n15901;
  assign n20749 = ~n54119 & n54719;
  assign n20750 = ~n54073 & n15921;
  assign n20751 = ~n20749 & ~n20750;
  assign n20752 = ~n20748 & ~n20749;
  assign n20753 = ~n20750 & n20752;
  assign n20754 = ~n20748 & ~n20750;
  assign n20755 = ~n20749 & n20754;
  assign n20756 = ~n20748 & n20751;
  assign n20757 = ~n14413 & n55588;
  assign n20758 = ~n15779 & n55588;
  assign n20759 = ~n20757 & ~n20758;
  assign n20760 = ~n20747 & n55588;
  assign n20761 = pi20  & ~n55589;
  assign n20762 = ~pi20  & n55589;
  assign n20763 = ~n20761 & ~n20762;
  assign n20764 = n20746 & ~n20763;
  assign n20765 = n20489 & n55547;
  assign n20766 = ~n20497 & ~n20765;
  assign n20767 = n14413 & n16547;
  assign n20768 = ~n54119 & n15901;
  assign n20769 = ~n54098 & n15921;
  assign n20770 = ~n54132 & n54719;
  assign n20771 = ~n20769 & ~n20770;
  assign n20772 = ~n20768 & ~n20770;
  assign n20773 = ~n20769 & n20772;
  assign n20774 = ~n20768 & n20771;
  assign n20775 = ~n14413 & n55590;
  assign n20776 = ~n16547 & n55590;
  assign n20777 = ~n20775 & ~n20776;
  assign n20778 = ~n20767 & n55590;
  assign n20779 = pi20  & ~n55591;
  assign n20780 = ~pi20  & n55591;
  assign n20781 = ~n20779 & ~n20780;
  assign n20782 = n20766 & ~n20781;
  assign n20783 = n20482 & n55544;
  assign n20784 = ~n20488 & ~n20783;
  assign n20785 = n14413 & n16772;
  assign n20786 = ~n54154 & n54719;
  assign n20787 = ~n54119 & n15921;
  assign n20788 = ~n54132 & n15901;
  assign n20789 = ~n20787 & ~n20788;
  assign n20790 = ~n20786 & ~n20788;
  assign n20791 = ~n20787 & n20790;
  assign n20792 = ~n20786 & n20789;
  assign n20793 = ~n14413 & n55592;
  assign n20794 = ~n16772 & n55592;
  assign n20795 = ~n20793 & ~n20794;
  assign n20796 = ~n20785 & n55592;
  assign n20797 = pi20  & ~n55593;
  assign n20798 = ~pi20  & n55593;
  assign n20799 = ~n20797 & ~n20798;
  assign n20800 = n20784 & ~n20799;
  assign n20801 = n14413 & n16522;
  assign n20802 = ~n54154 & n15901;
  assign n20803 = ~n54132 & n15921;
  assign n20804 = ~n54163 & n54719;
  assign n20805 = ~n20803 & ~n20804;
  assign n20806 = ~n20802 & ~n20804;
  assign n20807 = ~n20803 & n20806;
  assign n20808 = ~n20802 & n20805;
  assign n20809 = ~n20801 & n55594;
  assign n20810 = pi20  & ~n20809;
  assign n20811 = ~n20809 & ~n20810;
  assign n20812 = ~pi20  & ~n20809;
  assign n20813 = pi20  & ~n20810;
  assign n20814 = pi20  & n20809;
  assign n20815 = ~n55595 & ~n55596;
  assign n20816 = n20478 & ~n20480;
  assign n20817 = ~n20481 & ~n20816;
  assign n20818 = ~n20815 & n20817;
  assign n20819 = n14413 & n17072;
  assign n20820 = ~n54154 & n15921;
  assign n20821 = ~n54183 & n54719;
  assign n20822 = ~n54163 & n15901;
  assign n20823 = ~n20821 & ~n20822;
  assign n20824 = ~n20820 & n20823;
  assign n20825 = ~n20819 & n20824;
  assign n20826 = pi20  & ~n20825;
  assign n20827 = ~n20825 & ~n20826;
  assign n20828 = ~pi20  & ~n20825;
  assign n20829 = pi20  & ~n20826;
  assign n20830 = pi20  & n20825;
  assign n20831 = ~n55597 & ~n55598;
  assign n20832 = n20469 & n55543;
  assign n20833 = ~n20469 & ~n20477;
  assign n20834 = ~n20469 & n55543;
  assign n20835 = ~n55543 & ~n20477;
  assign n20836 = n20469 & ~n55543;
  assign n20837 = ~n55599 & ~n55600;
  assign n20838 = ~n20477 & ~n20832;
  assign n20839 = ~n20831 & ~n55601;
  assign n20840 = n20460 & n55540;
  assign n20841 = ~n20468 & ~n20840;
  assign n20842 = n14413 & n17524;
  assign n20843 = ~n54183 & n15901;
  assign n20844 = ~n54194 & n54719;
  assign n20845 = ~n54163 & n15921;
  assign n20846 = ~n20844 & ~n20845;
  assign n20847 = ~n20843 & ~n20844;
  assign n20848 = ~n20845 & n20847;
  assign n20849 = ~n20843 & n20846;
  assign n20850 = ~n14413 & n55602;
  assign n20851 = ~n17524 & n55602;
  assign n20852 = ~n20850 & ~n20851;
  assign n20853 = ~n20842 & n55602;
  assign n20854 = pi20  & ~n55603;
  assign n20855 = ~pi20  & n55603;
  assign n20856 = ~n20854 & ~n20855;
  assign n20857 = n20841 & ~n20856;
  assign n20858 = n20456 & ~n20458;
  assign n20859 = ~n20459 & ~n20858;
  assign n20860 = n14413 & n17544;
  assign n20861 = ~n54212 & n54719;
  assign n20862 = ~n54183 & n15921;
  assign n20863 = ~n54194 & n15901;
  assign n20864 = ~n20862 & ~n20863;
  assign n20865 = ~n20861 & ~n20863;
  assign n20866 = ~n20862 & n20865;
  assign n20867 = ~n20861 & n20864;
  assign n20868 = ~n14413 & n55604;
  assign n20869 = ~n17544 & n55604;
  assign n20870 = ~n20868 & ~n20869;
  assign n20871 = ~n20860 & n55604;
  assign n20872 = pi20  & ~n55605;
  assign n20873 = ~pi20  & n55605;
  assign n20874 = ~n20872 & ~n20873;
  assign n20875 = n20859 & ~n20874;
  assign n20876 = n20447 & n55537;
  assign n20877 = ~n20455 & ~n20876;
  assign n20878 = n14413 & n17041;
  assign n20879 = ~n54212 & n15901;
  assign n20880 = ~n54194 & n15921;
  assign n20881 = ~n54240 & n54719;
  assign n20882 = ~n20880 & ~n20881;
  assign n20883 = ~n20879 & ~n20881;
  assign n20884 = ~n20880 & n20883;
  assign n20885 = ~n20879 & n20882;
  assign n20886 = ~n14413 & n55606;
  assign n20887 = ~n17041 & n55606;
  assign n20888 = ~n20886 & ~n20887;
  assign n20889 = ~n20878 & n55606;
  assign n20890 = pi20  & ~n55607;
  assign n20891 = ~pi20  & n55607;
  assign n20892 = ~n20890 & ~n20891;
  assign n20893 = n20877 & ~n20892;
  assign n20894 = n14413 & n17660;
  assign n20895 = ~n54254 & n54719;
  assign n20896 = ~n54212 & n15921;
  assign n20897 = ~n54240 & n15901;
  assign n20898 = ~n20896 & ~n20897;
  assign n20899 = ~n20895 & ~n20897;
  assign n20900 = ~n20896 & n20899;
  assign n20901 = ~n20895 & n20898;
  assign n20902 = ~n20894 & n55608;
  assign n20903 = pi20  & ~n20902;
  assign n20904 = ~n20902 & ~n20903;
  assign n20905 = ~pi20  & ~n20902;
  assign n20906 = pi20  & ~n20903;
  assign n20907 = pi20  & n20902;
  assign n20908 = ~n55609 & ~n55610;
  assign n20909 = n20443 & ~n20445;
  assign n20910 = ~n20446 & ~n20909;
  assign n20911 = ~n20908 & n20910;
  assign n20912 = n14413 & n17804;
  assign n20913 = ~n54254 & n15901;
  assign n20914 = ~n54240 & n15921;
  assign n20915 = ~n54269 & n54719;
  assign n20916 = ~n20914 & ~n20915;
  assign n20917 = ~n20913 & ~n20915;
  assign n20918 = ~n20914 & n20917;
  assign n20919 = ~n20913 & n20916;
  assign n20920 = ~n14413 & n55611;
  assign n20921 = ~n17804 & n55611;
  assign n20922 = ~n20920 & ~n20921;
  assign n20923 = ~n20912 & n55611;
  assign n20924 = pi20  & ~n55612;
  assign n20925 = ~pi20  & n55612;
  assign n20926 = ~n20924 & ~n20925;
  assign n20927 = n20434 & n55534;
  assign n20928 = ~n55534 & ~n20442;
  assign n20929 = ~n20434 & ~n20442;
  assign n20930 = ~n20928 & ~n20929;
  assign n20931 = ~n20442 & ~n20927;
  assign n20932 = ~n20926 & ~n55613;
  assign n20933 = n14413 & n17939;
  assign n20934 = ~n54254 & n15921;
  assign n20935 = ~n54277 & n54719;
  assign n20936 = ~n54269 & n15901;
  assign n20937 = ~n20935 & ~n20936;
  assign n20938 = ~n20934 & n20937;
  assign n20939 = ~n20933 & n20938;
  assign n20940 = pi20  & ~n20939;
  assign n20941 = ~n20939 & ~n20940;
  assign n20942 = ~pi20  & ~n20939;
  assign n20943 = pi20  & ~n20940;
  assign n20944 = pi20  & n20939;
  assign n20945 = ~n55614 & ~n55615;
  assign n20946 = pi23  & ~n55526;
  assign n20947 = ~n55527 & ~n20946;
  assign n20948 = n55527 & n20946;
  assign n20949 = ~n55526 & n20416;
  assign n20950 = ~n55528 & ~n20949;
  assign n20951 = ~n20947 & ~n20948;
  assign n20952 = ~n20945 & n55616;
  assign n20953 = n14413 & n18056;
  assign n20954 = ~n54305 & n54719;
  assign n20955 = ~n54277 & n15901;
  assign n20956 = ~n54269 & n15921;
  assign n20957 = ~n20955 & ~n20956;
  assign n20958 = ~n20954 & ~n20955;
  assign n20959 = ~n20956 & n20958;
  assign n20960 = ~n20954 & n20957;
  assign n20961 = ~n14413 & n55617;
  assign n20962 = ~n18056 & n55617;
  assign n20963 = ~n20961 & ~n20962;
  assign n20964 = ~n20953 & n55617;
  assign n20965 = pi20  & ~n55618;
  assign n20966 = ~pi20  & n55618;
  assign n20967 = ~n20965 & ~n20966;
  assign n20968 = pi23  & n20396;
  assign n20969 = ~n20395 & n20968;
  assign n20970 = n20395 & ~n20968;
  assign n20971 = ~n20397 & n20401;
  assign n20972 = ~n55526 & ~n20971;
  assign n20973 = ~n20969 & ~n20970;
  assign n20974 = ~n20967 & n55619;
  assign n20975 = n14413 & ~n19275;
  assign n20976 = ~n54325 & n15901;
  assign n20977 = ~n54344 & n15921;
  assign n20978 = ~n20976 & ~n20977;
  assign n20979 = ~n20975 & n20978;
  assign n20980 = ~n54325 & n54717;
  assign n20981 = pi20  & ~n20980;
  assign n20982 = pi20  & ~n20979;
  assign n20983 = pi20  & ~n20982;
  assign n20984 = ~n20979 & ~n20982;
  assign n20985 = ~n20983 & ~n20984;
  assign n20986 = n20981 & ~n20985;
  assign n20987 = n20979 & n20981;
  assign n20988 = n14413 & n18156;
  assign n20989 = ~n54305 & n15921;
  assign n20990 = ~n54325 & n54719;
  assign n20991 = ~n54344 & n15901;
  assign n20992 = ~n20990 & ~n20991;
  assign n20993 = ~n20989 & n20992;
  assign n20994 = ~n14413 & n20993;
  assign n20995 = ~n18156 & n20993;
  assign n20996 = ~n20994 & ~n20995;
  assign n20997 = ~n20988 & n20993;
  assign n20998 = pi20  & ~n55621;
  assign n20999 = ~pi20  & n55621;
  assign n21000 = ~n20998 & ~n20999;
  assign n21001 = n55620 & ~n21000;
  assign n21002 = n55620 & ~n55621;
  assign n21003 = n20396 & n55622;
  assign n21004 = n14413 & n18336;
  assign n21005 = ~n54305 & n15901;
  assign n21006 = ~n54277 & n15921;
  assign n21007 = ~n54344 & n54719;
  assign n21008 = ~n21006 & ~n21007;
  assign n21009 = ~n21005 & ~n21007;
  assign n21010 = ~n21006 & n21009;
  assign n21011 = ~n21005 & n21008;
  assign n21012 = ~n21004 & n55623;
  assign n21013 = pi20  & ~n21012;
  assign n21014 = pi20  & ~n21013;
  assign n21015 = pi20  & n21012;
  assign n21016 = ~n21012 & ~n21013;
  assign n21017 = ~pi20  & ~n21012;
  assign n21018 = ~n55624 & ~n55625;
  assign n21019 = ~n20396 & ~n55622;
  assign n21020 = n55622 & ~n21003;
  assign n21021 = ~n20396 & n55622;
  assign n21022 = n20396 & ~n21003;
  assign n21023 = n20396 & ~n55622;
  assign n21024 = ~n55626 & ~n55627;
  assign n21025 = ~n21003 & ~n21019;
  assign n21026 = ~n21018 & ~n55628;
  assign n21027 = ~n21003 & ~n21026;
  assign n21028 = n20967 & ~n55619;
  assign n21029 = ~n20974 & ~n21028;
  assign n21030 = ~n21027 & n21029;
  assign n21031 = ~n20974 & ~n21030;
  assign n21032 = n20945 & ~n55616;
  assign n21033 = ~n20945 & ~n20952;
  assign n21034 = ~n20945 & ~n55616;
  assign n21035 = n55616 & ~n20952;
  assign n21036 = n20945 & n55616;
  assign n21037 = ~n55629 & ~n55630;
  assign n21038 = ~n20952 & ~n21032;
  assign n21039 = ~n21031 & ~n55631;
  assign n21040 = ~n20952 & ~n21039;
  assign n21041 = n20926 & n55613;
  assign n21042 = ~n20932 & ~n21041;
  assign n21043 = ~n21040 & n21042;
  assign n21044 = ~n20932 & ~n21043;
  assign n21045 = n20908 & ~n20910;
  assign n21046 = ~n20908 & ~n20911;
  assign n21047 = ~n20908 & ~n20910;
  assign n21048 = n20910 & ~n20911;
  assign n21049 = n20908 & n20910;
  assign n21050 = ~n55632 & ~n55633;
  assign n21051 = ~n20911 & ~n21045;
  assign n21052 = ~n21044 & ~n55634;
  assign n21053 = ~n20911 & ~n21052;
  assign n21054 = ~n20877 & n20892;
  assign n21055 = n20877 & ~n20893;
  assign n21056 = n20877 & n20892;
  assign n21057 = ~n20892 & ~n20893;
  assign n21058 = ~n20877 & ~n20892;
  assign n21059 = ~n55635 & ~n55636;
  assign n21060 = ~n20893 & ~n21054;
  assign n21061 = ~n21053 & ~n55637;
  assign n21062 = ~n20893 & ~n21061;
  assign n21063 = ~n20859 & n20874;
  assign n21064 = n20859 & ~n20875;
  assign n21065 = n20859 & n20874;
  assign n21066 = ~n20874 & ~n20875;
  assign n21067 = ~n20859 & ~n20874;
  assign n21068 = ~n55638 & ~n55639;
  assign n21069 = ~n20875 & ~n21063;
  assign n21070 = ~n21062 & ~n55640;
  assign n21071 = ~n20875 & ~n21070;
  assign n21072 = ~n20841 & n20856;
  assign n21073 = ~n20857 & ~n21072;
  assign n21074 = ~n21071 & n21073;
  assign n21075 = ~n20857 & ~n21074;
  assign n21076 = n20831 & n55601;
  assign n21077 = ~n20831 & ~n20839;
  assign n21078 = ~n55601 & ~n20839;
  assign n21079 = ~n21077 & ~n21078;
  assign n21080 = ~n20839 & ~n21076;
  assign n21081 = ~n21075 & ~n55641;
  assign n21082 = ~n20839 & ~n21081;
  assign n21083 = n20815 & ~n20817;
  assign n21084 = ~n20815 & ~n20818;
  assign n21085 = ~n20815 & ~n20817;
  assign n21086 = n20817 & ~n20818;
  assign n21087 = n20815 & n20817;
  assign n21088 = ~n55642 & ~n55643;
  assign n21089 = ~n20818 & ~n21083;
  assign n21090 = ~n21082 & ~n55644;
  assign n21091 = ~n20818 & ~n21090;
  assign n21092 = ~n20784 & n20799;
  assign n21093 = n20784 & ~n20800;
  assign n21094 = n20784 & n20799;
  assign n21095 = ~n20799 & ~n20800;
  assign n21096 = ~n20784 & ~n20799;
  assign n21097 = ~n55645 & ~n55646;
  assign n21098 = ~n20800 & ~n21092;
  assign n21099 = ~n21091 & ~n55647;
  assign n21100 = ~n20800 & ~n21099;
  assign n21101 = ~n20766 & n20781;
  assign n21102 = n20766 & ~n20782;
  assign n21103 = n20766 & n20781;
  assign n21104 = ~n20781 & ~n20782;
  assign n21105 = ~n20766 & ~n20781;
  assign n21106 = ~n55648 & ~n55649;
  assign n21107 = ~n20782 & ~n21101;
  assign n21108 = ~n21100 & ~n55650;
  assign n21109 = ~n20782 & ~n21108;
  assign n21110 = ~n20746 & n20763;
  assign n21111 = n20746 & ~n20764;
  assign n21112 = n20746 & n20763;
  assign n21113 = ~n20763 & ~n20764;
  assign n21114 = ~n20746 & ~n20763;
  assign n21115 = ~n55651 & ~n55652;
  assign n21116 = ~n20764 & ~n21110;
  assign n21117 = ~n21109 & ~n55653;
  assign n21118 = ~n20764 & ~n21117;
  assign n21119 = ~n20728 & n20743;
  assign n21120 = n20728 & ~n20744;
  assign n21121 = n20728 & n20743;
  assign n21122 = ~n20743 & ~n20744;
  assign n21123 = ~n20728 & ~n20743;
  assign n21124 = ~n55654 & ~n55655;
  assign n21125 = ~n20744 & ~n21119;
  assign n21126 = ~n21118 & ~n55656;
  assign n21127 = ~n20744 & ~n21126;
  assign n21128 = ~n20710 & n20725;
  assign n21129 = n20710 & ~n20726;
  assign n21130 = n20710 & n20725;
  assign n21131 = ~n20725 & ~n20726;
  assign n21132 = ~n20710 & ~n20725;
  assign n21133 = ~n55657 & ~n55658;
  assign n21134 = ~n20726 & ~n21128;
  assign n21135 = ~n21127 & ~n55659;
  assign n21136 = ~n20726 & ~n21135;
  assign n21137 = ~n20692 & n20707;
  assign n21138 = n20692 & ~n20708;
  assign n21139 = n20692 & n20707;
  assign n21140 = ~n20707 & ~n20708;
  assign n21141 = ~n20692 & ~n20707;
  assign n21142 = ~n55660 & ~n55661;
  assign n21143 = ~n20708 & ~n21137;
  assign n21144 = ~n21136 & ~n55662;
  assign n21145 = ~n20708 & ~n21144;
  assign n21146 = ~n20674 & n20689;
  assign n21147 = n20674 & ~n20690;
  assign n21148 = n20674 & n20689;
  assign n21149 = ~n20689 & ~n20690;
  assign n21150 = ~n20674 & ~n20689;
  assign n21151 = ~n55663 & ~n55664;
  assign n21152 = ~n20690 & ~n21146;
  assign n21153 = ~n21145 & ~n55665;
  assign n21154 = ~n20690 & ~n21153;
  assign n21155 = n20557 & ~n20559;
  assign n21156 = ~n20560 & ~n21155;
  assign n21157 = ~n21154 & n21156;
  assign n21158 = n13360 & n16079;
  assign n21159 = ~n53907 & n16676;
  assign n21160 = ~n53930 & n54886;
  assign n21161 = ~n53888 & n16696;
  assign n21162 = ~n21160 & ~n21161;
  assign n21163 = ~n21159 & ~n21160;
  assign n21164 = ~n21161 & n21163;
  assign n21165 = ~n21159 & n21162;
  assign n21166 = ~n21158 & n55666;
  assign n21167 = pi17  & ~n21166;
  assign n21168 = ~n21166 & ~n21167;
  assign n21169 = ~pi17  & ~n21166;
  assign n21170 = pi17  & ~n21167;
  assign n21171 = pi17  & n21166;
  assign n21172 = ~n55667 & ~n55668;
  assign n21173 = n21154 & ~n21156;
  assign n21174 = ~n21157 & ~n21173;
  assign n21175 = ~n21172 & n21174;
  assign n21176 = ~n21157 & ~n21175;
  assign n21177 = n20585 & ~n20586;
  assign n21178 = n20583 & n20585;
  assign n21179 = ~n20583 & ~n20586;
  assign n21180 = ~n20583 & ~n20585;
  assign n21181 = n20583 & ~n20585;
  assign n21182 = ~n20586 & ~n21181;
  assign n21183 = ~n55669 & ~n55670;
  assign n21184 = ~n21176 & n55671;
  assign n21185 = n21176 & ~n55671;
  assign n21186 = n12550 & n17265;
  assign n21187 = ~n53819 & n18556;
  assign n21188 = ~n53845 & n55041;
  assign n21189 = ~n53799 & n18588;
  assign n21190 = ~n21188 & ~n21189;
  assign n21191 = ~n21187 & ~n21188;
  assign n21192 = ~n21189 & n21191;
  assign n21193 = ~n21187 & n21190;
  assign n21194 = ~n21186 & n55672;
  assign n21195 = pi14  & ~n21194;
  assign n21196 = pi14  & ~n21195;
  assign n21197 = pi14  & n21194;
  assign n21198 = ~n21194 & ~n21195;
  assign n21199 = ~pi14  & ~n21194;
  assign n21200 = ~n55673 & ~n55674;
  assign n21201 = ~n21185 & ~n21200;
  assign n21202 = ~n21184 & ~n21185;
  assign n21203 = ~n21200 & n21202;
  assign n21204 = ~n21184 & ~n21203;
  assign n21205 = ~n21184 & ~n21201;
  assign n21206 = ~n55579 & ~n55675;
  assign n21207 = n55579 & n55675;
  assign n21208 = n11360 & n18846;
  assign n21209 = ~n53685 & n19541;
  assign n21210 = ~n53741 & n55247;
  assign n21211 = ~n53712 & n19509;
  assign n21212 = ~n21210 & ~n21211;
  assign n21213 = ~n21209 & ~n21210;
  assign n21214 = ~n21211 & n21213;
  assign n21215 = ~n21209 & n21212;
  assign n21216 = ~n21208 & n55676;
  assign n21217 = pi11  & ~n21216;
  assign n21218 = pi11  & ~n21217;
  assign n21219 = pi11  & n21216;
  assign n21220 = ~n21216 & ~n21217;
  assign n21221 = ~pi11  & ~n21216;
  assign n21222 = ~n55677 & ~n55678;
  assign n21223 = ~n21207 & ~n21222;
  assign n21224 = ~n21206 & ~n21207;
  assign n21225 = ~n21222 & n21224;
  assign n21226 = ~n21206 & ~n21225;
  assign n21227 = ~n21206 & ~n21223;
  assign n21228 = ~n20667 & ~n55679;
  assign n21229 = n20667 & n55679;
  assign n21230 = ~n21228 & ~n21229;
  assign n21231 = ~n20115 & n55570;
  assign n21232 = ~n20611 & ~n21231;
  assign n21233 = n21230 & n21232;
  assign n21234 = ~n21228 & ~n21233;
  assign n21235 = n54351 & n20085;
  assign n21236 = ~n53634 & n55472;
  assign n21237 = ~n55469 & n55470;
  assign n21238 = ~n2325 & n21237;
  assign n21239 = ~n21236 & ~n21238;
  assign n21240 = ~n20085 & n21239;
  assign n21241 = ~n54351 & n21239;
  assign n21242 = ~n21240 & ~n21241;
  assign n21243 = ~n21235 & n21239;
  assign n21244 = pi8  & ~n55680;
  assign n21245 = ~pi8  & n55680;
  assign n21246 = ~n21244 & ~n21245;
  assign n21247 = ~n21234 & ~n21246;
  assign n21248 = n21234 & n21246;
  assign n21249 = ~n21247 & ~n21248;
  assign n21250 = n20634 & ~n20635;
  assign n21251 = n20632 & n20634;
  assign n21252 = ~n20632 & ~n20635;
  assign n21253 = ~n20632 & ~n20634;
  assign n21254 = n20632 & ~n20634;
  assign n21255 = ~n20635 & ~n21254;
  assign n21256 = ~n55681 & ~n55682;
  assign n21257 = n21249 & n55683;
  assign n21258 = ~n21247 & ~n21257;
  assign n21259 = n55575 & ~n20646;
  assign n21260 = ~n55575 & ~n20647;
  assign n21261 = n20646 & ~n20647;
  assign n21262 = ~n21260 & ~n21261;
  assign n21263 = ~n20647 & ~n21259;
  assign n21264 = ~n21258 & ~n55684;
  assign n21265 = n21258 & n55684;
  assign n21266 = ~n21264 & ~n21265;
  assign n21267 = n11242 & n20085;
  assign n21268 = ~n53650 & n55472;
  assign n21269 = n55469 & ~n55471;
  assign n21270 = ~n2325 & n21269;
  assign n21271 = ~n53634 & n21237;
  assign n21272 = ~n21270 & ~n21271;
  assign n21273 = ~n21268 & ~n21271;
  assign n21274 = ~n21270 & n21273;
  assign n21275 = ~n21268 & n21272;
  assign n21276 = ~n20085 & n55685;
  assign n21277 = ~n11242 & n55685;
  assign n21278 = ~n21276 & ~n21277;
  assign n21279 = ~n21267 & n55685;
  assign n21280 = pi8  & ~n55686;
  assign n21281 = ~pi8  & n55686;
  assign n21282 = ~n21280 & ~n21281;
  assign n21283 = n21222 & ~n21224;
  assign n21284 = n21224 & ~n21225;
  assign n21285 = ~n21222 & ~n21225;
  assign n21286 = ~n21284 & ~n21285;
  assign n21287 = ~n21225 & ~n21283;
  assign n21288 = n14263 & n16079;
  assign n21289 = ~n53930 & n16676;
  assign n21290 = ~n53962 & n54886;
  assign n21291 = ~n53907 & n16696;
  assign n21292 = ~n21290 & ~n21291;
  assign n21293 = ~n21289 & ~n21290;
  assign n21294 = ~n21291 & n21293;
  assign n21295 = ~n21289 & n21292;
  assign n21296 = ~n21288 & n55688;
  assign n21297 = pi17  & ~n21296;
  assign n21298 = ~n21296 & ~n21297;
  assign n21299 = ~pi17  & ~n21296;
  assign n21300 = pi17  & ~n21297;
  assign n21301 = pi17  & n21296;
  assign n21302 = ~n55689 & ~n55690;
  assign n21303 = n21145 & n55665;
  assign n21304 = ~n21145 & ~n21153;
  assign n21305 = ~n21145 & n55665;
  assign n21306 = ~n55665 & ~n21153;
  assign n21307 = n21145 & ~n55665;
  assign n21308 = ~n55691 & ~n55692;
  assign n21309 = ~n21153 & ~n21303;
  assign n21310 = ~n21302 & ~n55693;
  assign n21311 = n14020 & n16079;
  assign n21312 = ~n53962 & n16676;
  assign n21313 = ~n53970 & n54886;
  assign n21314 = ~n53930 & n16696;
  assign n21315 = ~n21313 & ~n21314;
  assign n21316 = ~n21312 & ~n21313;
  assign n21317 = ~n21314 & n21316;
  assign n21318 = ~n21312 & n21315;
  assign n21319 = ~n21311 & n55694;
  assign n21320 = pi17  & ~n21319;
  assign n21321 = ~n21319 & ~n21320;
  assign n21322 = ~pi17  & ~n21319;
  assign n21323 = pi17  & ~n21320;
  assign n21324 = pi17  & n21319;
  assign n21325 = ~n55695 & ~n55696;
  assign n21326 = n21136 & n55662;
  assign n21327 = ~n21136 & ~n21144;
  assign n21328 = ~n21136 & n55662;
  assign n21329 = ~n55662 & ~n21144;
  assign n21330 = n21136 & ~n55662;
  assign n21331 = ~n55697 & ~n55698;
  assign n21332 = ~n21144 & ~n21326;
  assign n21333 = ~n21325 & ~n55699;
  assign n21334 = n14708 & n16079;
  assign n21335 = ~n54005 & n54886;
  assign n21336 = ~n53970 & n16676;
  assign n21337 = ~n53962 & n16696;
  assign n21338 = ~n21336 & ~n21337;
  assign n21339 = ~n21335 & ~n21336;
  assign n21340 = ~n21337 & n21339;
  assign n21341 = ~n21335 & n21338;
  assign n21342 = ~n21334 & n55700;
  assign n21343 = pi17  & ~n21342;
  assign n21344 = ~n21342 & ~n21343;
  assign n21345 = ~pi17  & ~n21342;
  assign n21346 = pi17  & ~n21343;
  assign n21347 = pi17  & n21342;
  assign n21348 = ~n55701 & ~n55702;
  assign n21349 = n21127 & n55659;
  assign n21350 = ~n21127 & ~n21135;
  assign n21351 = ~n55659 & ~n21135;
  assign n21352 = ~n21350 & ~n21351;
  assign n21353 = ~n21135 & ~n21349;
  assign n21354 = ~n21348 & ~n55703;
  assign n21355 = n14688 & n16079;
  assign n21356 = ~n54005 & n16676;
  assign n21357 = ~n54034 & n54886;
  assign n21358 = ~n53970 & n16696;
  assign n21359 = ~n21357 & ~n21358;
  assign n21360 = ~n21356 & ~n21357;
  assign n21361 = ~n21358 & n21360;
  assign n21362 = ~n21356 & n21359;
  assign n21363 = ~n21355 & n55704;
  assign n21364 = pi17  & ~n21363;
  assign n21365 = ~n21363 & ~n21364;
  assign n21366 = ~pi17  & ~n21363;
  assign n21367 = pi17  & ~n21364;
  assign n21368 = pi17  & n21363;
  assign n21369 = ~n55705 & ~n55706;
  assign n21370 = n21118 & n55656;
  assign n21371 = ~n21118 & ~n21126;
  assign n21372 = ~n55656 & ~n21126;
  assign n21373 = ~n21371 & ~n21372;
  assign n21374 = ~n21126 & ~n21370;
  assign n21375 = ~n21369 & ~n55707;
  assign n21376 = n15195 & n16079;
  assign n21377 = ~n54050 & n54886;
  assign n21378 = ~n54005 & n16696;
  assign n21379 = ~n54034 & n16676;
  assign n21380 = ~n21378 & ~n21379;
  assign n21381 = ~n21377 & ~n21379;
  assign n21382 = ~n21378 & n21381;
  assign n21383 = ~n21377 & n21380;
  assign n21384 = ~n21376 & n55708;
  assign n21385 = pi17  & ~n21384;
  assign n21386 = ~n21384 & ~n21385;
  assign n21387 = ~pi17  & ~n21384;
  assign n21388 = pi17  & ~n21385;
  assign n21389 = pi17  & n21384;
  assign n21390 = ~n55709 & ~n55710;
  assign n21391 = n21109 & n55653;
  assign n21392 = ~n21109 & ~n21117;
  assign n21393 = ~n21109 & n55653;
  assign n21394 = ~n55653 & ~n21117;
  assign n21395 = n21109 & ~n55653;
  assign n21396 = ~n55711 & ~n55712;
  assign n21397 = ~n21117 & ~n21391;
  assign n21398 = ~n21390 & ~n55713;
  assign n21399 = n15219 & n16079;
  assign n21400 = ~n54050 & n16676;
  assign n21401 = ~n54034 & n16696;
  assign n21402 = ~n54073 & n54886;
  assign n21403 = ~n21401 & ~n21402;
  assign n21404 = ~n21400 & ~n21402;
  assign n21405 = ~n21401 & n21404;
  assign n21406 = ~n21400 & n21403;
  assign n21407 = ~n21399 & n55714;
  assign n21408 = pi17  & ~n21407;
  assign n21409 = ~n21407 & ~n21408;
  assign n21410 = ~pi17  & ~n21407;
  assign n21411 = pi17  & ~n21408;
  assign n21412 = pi17  & n21407;
  assign n21413 = ~n55715 & ~n55716;
  assign n21414 = n21100 & n55650;
  assign n21415 = ~n21100 & ~n21108;
  assign n21416 = ~n21100 & n55650;
  assign n21417 = ~n55650 & ~n21108;
  assign n21418 = n21100 & ~n55650;
  assign n21419 = ~n55717 & ~n55718;
  assign n21420 = ~n21108 & ~n21414;
  assign n21421 = ~n21413 & ~n55719;
  assign n21422 = n16079 & n16138;
  assign n21423 = ~n54098 & n54886;
  assign n21424 = ~n54050 & n16696;
  assign n21425 = ~n54073 & n16676;
  assign n21426 = ~n21424 & ~n21425;
  assign n21427 = ~n21423 & ~n21425;
  assign n21428 = ~n21424 & n21427;
  assign n21429 = ~n21423 & n21426;
  assign n21430 = ~n21422 & n55720;
  assign n21431 = pi17  & ~n21430;
  assign n21432 = ~n21430 & ~n21431;
  assign n21433 = ~pi17  & ~n21430;
  assign n21434 = pi17  & ~n21431;
  assign n21435 = pi17  & n21430;
  assign n21436 = ~n55721 & ~n55722;
  assign n21437 = n21091 & n55647;
  assign n21438 = ~n21091 & ~n21099;
  assign n21439 = ~n55647 & ~n21099;
  assign n21440 = ~n21438 & ~n21439;
  assign n21441 = ~n21099 & ~n21437;
  assign n21442 = ~n21436 & ~n55723;
  assign n21443 = n21082 & n55644;
  assign n21444 = ~n21090 & ~n21443;
  assign n21445 = n15779 & n16079;
  assign n21446 = ~n54098 & n16676;
  assign n21447 = ~n54119 & n54886;
  assign n21448 = ~n54073 & n16696;
  assign n21449 = ~n21447 & ~n21448;
  assign n21450 = ~n21446 & ~n21447;
  assign n21451 = ~n21448 & n21450;
  assign n21452 = ~n21446 & ~n21448;
  assign n21453 = ~n21447 & n21452;
  assign n21454 = ~n21446 & n21449;
  assign n21455 = ~n16079 & n55724;
  assign n21456 = ~n15779 & n55724;
  assign n21457 = ~n21455 & ~n21456;
  assign n21458 = ~n21445 & n55724;
  assign n21459 = pi17  & ~n55725;
  assign n21460 = ~pi17  & n55725;
  assign n21461 = ~n21459 & ~n21460;
  assign n21462 = n21444 & ~n21461;
  assign n21463 = n21075 & n55641;
  assign n21464 = ~n21081 & ~n21463;
  assign n21465 = n16079 & n16547;
  assign n21466 = ~n54119 & n16676;
  assign n21467 = ~n54098 & n16696;
  assign n21468 = ~n54132 & n54886;
  assign n21469 = ~n21467 & ~n21468;
  assign n21470 = ~n21466 & ~n21468;
  assign n21471 = ~n21467 & n21470;
  assign n21472 = ~n21466 & n21469;
  assign n21473 = ~n16079 & n55726;
  assign n21474 = ~n16547 & n55726;
  assign n21475 = ~n21473 & ~n21474;
  assign n21476 = ~n21465 & n55726;
  assign n21477 = pi17  & ~n55727;
  assign n21478 = ~pi17  & n55727;
  assign n21479 = ~n21477 & ~n21478;
  assign n21480 = n21464 & ~n21479;
  assign n21481 = n16079 & n16772;
  assign n21482 = ~n54154 & n54886;
  assign n21483 = ~n54119 & n16696;
  assign n21484 = ~n54132 & n16676;
  assign n21485 = ~n21483 & ~n21484;
  assign n21486 = ~n21482 & ~n21484;
  assign n21487 = ~n21483 & n21486;
  assign n21488 = ~n21482 & n21485;
  assign n21489 = ~n21481 & n55728;
  assign n21490 = pi17  & ~n21489;
  assign n21491 = ~n21489 & ~n21490;
  assign n21492 = ~pi17  & ~n21489;
  assign n21493 = pi17  & ~n21490;
  assign n21494 = pi17  & n21489;
  assign n21495 = ~n55729 & ~n55730;
  assign n21496 = n21071 & ~n21073;
  assign n21497 = ~n21074 & ~n21496;
  assign n21498 = ~n21495 & n21497;
  assign n21499 = n16079 & n16522;
  assign n21500 = ~n54154 & n16676;
  assign n21501 = ~n54132 & n16696;
  assign n21502 = ~n54163 & n54886;
  assign n21503 = ~n21501 & ~n21502;
  assign n21504 = ~n21500 & ~n21502;
  assign n21505 = ~n21501 & n21504;
  assign n21506 = ~n21500 & n21503;
  assign n21507 = ~n21499 & n55731;
  assign n21508 = pi17  & ~n21507;
  assign n21509 = ~n21507 & ~n21508;
  assign n21510 = ~pi17  & ~n21507;
  assign n21511 = pi17  & ~n21508;
  assign n21512 = pi17  & n21507;
  assign n21513 = ~n55732 & ~n55733;
  assign n21514 = n21062 & n55640;
  assign n21515 = ~n21062 & ~n21070;
  assign n21516 = ~n55640 & ~n21070;
  assign n21517 = ~n21515 & ~n21516;
  assign n21518 = ~n21070 & ~n21514;
  assign n21519 = ~n21513 & ~n55734;
  assign n21520 = n16079 & n17072;
  assign n21521 = ~n54154 & n16696;
  assign n21522 = ~n54183 & n54886;
  assign n21523 = ~n54163 & n16676;
  assign n21524 = ~n21522 & ~n21523;
  assign n21525 = ~n21521 & n21524;
  assign n21526 = ~n21520 & n21525;
  assign n21527 = pi17  & ~n21526;
  assign n21528 = ~n21526 & ~n21527;
  assign n21529 = ~pi17  & ~n21526;
  assign n21530 = pi17  & ~n21527;
  assign n21531 = pi17  & n21526;
  assign n21532 = ~n55735 & ~n55736;
  assign n21533 = n21053 & n55637;
  assign n21534 = ~n21053 & ~n21061;
  assign n21535 = ~n21053 & n55637;
  assign n21536 = ~n55637 & ~n21061;
  assign n21537 = n21053 & ~n55637;
  assign n21538 = ~n55737 & ~n55738;
  assign n21539 = ~n21061 & ~n21533;
  assign n21540 = ~n21532 & ~n55739;
  assign n21541 = n21044 & n55634;
  assign n21542 = ~n21052 & ~n21541;
  assign n21543 = n16079 & n17524;
  assign n21544 = ~n54183 & n16676;
  assign n21545 = ~n54194 & n54886;
  assign n21546 = ~n54163 & n16696;
  assign n21547 = ~n21545 & ~n21546;
  assign n21548 = ~n21544 & ~n21545;
  assign n21549 = ~n21546 & n21548;
  assign n21550 = ~n21544 & n21547;
  assign n21551 = ~n16079 & n55740;
  assign n21552 = ~n17524 & n55740;
  assign n21553 = ~n21551 & ~n21552;
  assign n21554 = ~n21543 & n55740;
  assign n21555 = pi17  & ~n55741;
  assign n21556 = ~pi17  & n55741;
  assign n21557 = ~n21555 & ~n21556;
  assign n21558 = n21542 & ~n21557;
  assign n21559 = n21040 & ~n21042;
  assign n21560 = ~n21043 & ~n21559;
  assign n21561 = n16079 & n17544;
  assign n21562 = ~n54212 & n54886;
  assign n21563 = ~n54183 & n16696;
  assign n21564 = ~n54194 & n16676;
  assign n21565 = ~n21563 & ~n21564;
  assign n21566 = ~n21562 & ~n21564;
  assign n21567 = ~n21563 & n21566;
  assign n21568 = ~n21562 & n21565;
  assign n21569 = ~n16079 & n55742;
  assign n21570 = ~n17544 & n55742;
  assign n21571 = ~n21569 & ~n21570;
  assign n21572 = ~n21561 & n55742;
  assign n21573 = pi17  & ~n55743;
  assign n21574 = ~pi17  & n55743;
  assign n21575 = ~n21573 & ~n21574;
  assign n21576 = n21560 & ~n21575;
  assign n21577 = n21031 & n55631;
  assign n21578 = ~n21039 & ~n21577;
  assign n21579 = n16079 & n17041;
  assign n21580 = ~n54212 & n16676;
  assign n21581 = ~n54194 & n16696;
  assign n21582 = ~n54240 & n54886;
  assign n21583 = ~n21581 & ~n21582;
  assign n21584 = ~n21580 & ~n21582;
  assign n21585 = ~n21581 & n21584;
  assign n21586 = ~n21580 & n21583;
  assign n21587 = ~n16079 & n55744;
  assign n21588 = ~n17041 & n55744;
  assign n21589 = ~n21587 & ~n21588;
  assign n21590 = ~n21579 & n55744;
  assign n21591 = pi17  & ~n55745;
  assign n21592 = ~pi17  & n55745;
  assign n21593 = ~n21591 & ~n21592;
  assign n21594 = n21578 & ~n21593;
  assign n21595 = n16079 & n17660;
  assign n21596 = ~n54254 & n54886;
  assign n21597 = ~n54212 & n16696;
  assign n21598 = ~n54240 & n16676;
  assign n21599 = ~n21597 & ~n21598;
  assign n21600 = ~n21596 & ~n21598;
  assign n21601 = ~n21597 & n21600;
  assign n21602 = ~n21596 & n21599;
  assign n21603 = ~n21595 & n55746;
  assign n21604 = pi17  & ~n21603;
  assign n21605 = ~n21603 & ~n21604;
  assign n21606 = ~pi17  & ~n21603;
  assign n21607 = pi17  & ~n21604;
  assign n21608 = pi17  & n21603;
  assign n21609 = ~n55747 & ~n55748;
  assign n21610 = n21027 & ~n21029;
  assign n21611 = ~n21030 & ~n21610;
  assign n21612 = ~n21609 & n21611;
  assign n21613 = n16079 & n17804;
  assign n21614 = ~n54254 & n16676;
  assign n21615 = ~n54240 & n16696;
  assign n21616 = ~n54269 & n54886;
  assign n21617 = ~n21615 & ~n21616;
  assign n21618 = ~n21614 & ~n21616;
  assign n21619 = ~n21615 & n21618;
  assign n21620 = ~n21614 & n21617;
  assign n21621 = ~n16079 & n55749;
  assign n21622 = ~n17804 & n55749;
  assign n21623 = ~n21621 & ~n21622;
  assign n21624 = ~n21613 & n55749;
  assign n21625 = pi17  & ~n55750;
  assign n21626 = ~pi17  & n55750;
  assign n21627 = ~n21625 & ~n21626;
  assign n21628 = n21018 & n55628;
  assign n21629 = ~n55628 & ~n21026;
  assign n21630 = ~n21018 & ~n21026;
  assign n21631 = ~n21629 & ~n21630;
  assign n21632 = ~n21026 & ~n21628;
  assign n21633 = ~n21627 & ~n55751;
  assign n21634 = n16079 & n17939;
  assign n21635 = ~n54254 & n16696;
  assign n21636 = ~n54277 & n54886;
  assign n21637 = ~n54269 & n16676;
  assign n21638 = ~n21636 & ~n21637;
  assign n21639 = ~n21635 & n21638;
  assign n21640 = ~n21634 & n21639;
  assign n21641 = pi17  & ~n21640;
  assign n21642 = ~n21640 & ~n21641;
  assign n21643 = ~pi17  & ~n21640;
  assign n21644 = pi17  & ~n21641;
  assign n21645 = pi17  & n21640;
  assign n21646 = ~n55752 & ~n55753;
  assign n21647 = pi20  & ~n55620;
  assign n21648 = ~n55621 & ~n21647;
  assign n21649 = n55621 & n21647;
  assign n21650 = ~n55620 & n21000;
  assign n21651 = ~n55622 & ~n21650;
  assign n21652 = ~n21648 & ~n21649;
  assign n21653 = ~n21646 & n55754;
  assign n21654 = n16079 & n18056;
  assign n21655 = ~n54305 & n54886;
  assign n21656 = ~n54277 & n16676;
  assign n21657 = ~n54269 & n16696;
  assign n21658 = ~n21656 & ~n21657;
  assign n21659 = ~n21655 & ~n21656;
  assign n21660 = ~n21657 & n21659;
  assign n21661 = ~n21655 & n21658;
  assign n21662 = ~n16079 & n55755;
  assign n21663 = ~n18056 & n55755;
  assign n21664 = ~n21662 & ~n21663;
  assign n21665 = ~n21654 & n55755;
  assign n21666 = pi17  & ~n55756;
  assign n21667 = ~pi17  & n55756;
  assign n21668 = ~n21666 & ~n21667;
  assign n21669 = pi20  & n20980;
  assign n21670 = ~n20979 & n21669;
  assign n21671 = n20979 & ~n21669;
  assign n21672 = ~n20981 & n20985;
  assign n21673 = ~n55620 & ~n21672;
  assign n21674 = ~n21670 & ~n21671;
  assign n21675 = ~n21668 & n55757;
  assign n21676 = n16079 & ~n19275;
  assign n21677 = ~n54325 & n16676;
  assign n21678 = ~n54344 & n16696;
  assign n21679 = ~n21677 & ~n21678;
  assign n21680 = ~n21676 & n21679;
  assign n21681 = ~n54325 & n54883;
  assign n21682 = pi17  & ~n21681;
  assign n21683 = pi17  & ~n21680;
  assign n21684 = pi17  & ~n21683;
  assign n21685 = ~n21680 & ~n21683;
  assign n21686 = ~n21684 & ~n21685;
  assign n21687 = n21682 & ~n21686;
  assign n21688 = n21680 & n21682;
  assign n21689 = n16079 & n18156;
  assign n21690 = ~n54305 & n16696;
  assign n21691 = ~n54325 & n54886;
  assign n21692 = ~n54344 & n16676;
  assign n21693 = ~n21691 & ~n21692;
  assign n21694 = ~n21690 & n21693;
  assign n21695 = ~n16079 & n21694;
  assign n21696 = ~n18156 & n21694;
  assign n21697 = ~n21695 & ~n21696;
  assign n21698 = ~n21689 & n21694;
  assign n21699 = pi17  & ~n55759;
  assign n21700 = ~pi17  & n55759;
  assign n21701 = ~n21699 & ~n21700;
  assign n21702 = n55758 & ~n21701;
  assign n21703 = n55758 & ~n55759;
  assign n21704 = n20980 & n55760;
  assign n21705 = n16079 & n18336;
  assign n21706 = ~n54305 & n16676;
  assign n21707 = ~n54277 & n16696;
  assign n21708 = ~n54344 & n54886;
  assign n21709 = ~n21707 & ~n21708;
  assign n21710 = ~n21706 & ~n21708;
  assign n21711 = ~n21707 & n21710;
  assign n21712 = ~n21706 & n21709;
  assign n21713 = ~n21705 & n55761;
  assign n21714 = pi17  & ~n21713;
  assign n21715 = pi17  & ~n21714;
  assign n21716 = pi17  & n21713;
  assign n21717 = ~n21713 & ~n21714;
  assign n21718 = ~pi17  & ~n21713;
  assign n21719 = ~n55762 & ~n55763;
  assign n21720 = ~n20980 & ~n55760;
  assign n21721 = n55760 & ~n21704;
  assign n21722 = ~n20980 & n55760;
  assign n21723 = n20980 & ~n21704;
  assign n21724 = n20980 & ~n55760;
  assign n21725 = ~n55764 & ~n55765;
  assign n21726 = ~n21704 & ~n21720;
  assign n21727 = ~n21719 & ~n55766;
  assign n21728 = ~n21704 & ~n21727;
  assign n21729 = n21668 & ~n55757;
  assign n21730 = ~n21675 & ~n21729;
  assign n21731 = ~n21728 & n21730;
  assign n21732 = ~n21675 & ~n21731;
  assign n21733 = n21646 & ~n55754;
  assign n21734 = ~n21646 & ~n21653;
  assign n21735 = ~n21646 & ~n55754;
  assign n21736 = n55754 & ~n21653;
  assign n21737 = n21646 & n55754;
  assign n21738 = ~n55767 & ~n55768;
  assign n21739 = ~n21653 & ~n21733;
  assign n21740 = ~n21732 & ~n55769;
  assign n21741 = ~n21653 & ~n21740;
  assign n21742 = n21627 & n55751;
  assign n21743 = ~n21633 & ~n21742;
  assign n21744 = ~n21741 & n21743;
  assign n21745 = ~n21633 & ~n21744;
  assign n21746 = n21609 & ~n21611;
  assign n21747 = ~n21609 & ~n21612;
  assign n21748 = ~n21609 & ~n21611;
  assign n21749 = n21611 & ~n21612;
  assign n21750 = n21609 & n21611;
  assign n21751 = ~n55770 & ~n55771;
  assign n21752 = ~n21612 & ~n21746;
  assign n21753 = ~n21745 & ~n55772;
  assign n21754 = ~n21612 & ~n21753;
  assign n21755 = ~n21578 & n21593;
  assign n21756 = n21578 & ~n21594;
  assign n21757 = n21578 & n21593;
  assign n21758 = ~n21593 & ~n21594;
  assign n21759 = ~n21578 & ~n21593;
  assign n21760 = ~n55773 & ~n55774;
  assign n21761 = ~n21594 & ~n21755;
  assign n21762 = ~n21754 & ~n55775;
  assign n21763 = ~n21594 & ~n21762;
  assign n21764 = ~n21560 & n21575;
  assign n21765 = n21560 & ~n21576;
  assign n21766 = n21560 & n21575;
  assign n21767 = ~n21575 & ~n21576;
  assign n21768 = ~n21560 & ~n21575;
  assign n21769 = ~n55776 & ~n55777;
  assign n21770 = ~n21576 & ~n21764;
  assign n21771 = ~n21763 & ~n55778;
  assign n21772 = ~n21576 & ~n21771;
  assign n21773 = ~n21542 & n21557;
  assign n21774 = ~n21558 & ~n21773;
  assign n21775 = ~n21772 & n21774;
  assign n21776 = ~n21558 & ~n21775;
  assign n21777 = n21532 & n55739;
  assign n21778 = ~n21532 & ~n21540;
  assign n21779 = ~n55739 & ~n21540;
  assign n21780 = ~n21778 & ~n21779;
  assign n21781 = ~n21540 & ~n21777;
  assign n21782 = ~n21776 & ~n55779;
  assign n21783 = ~n21540 & ~n21782;
  assign n21784 = n21513 & n55734;
  assign n21785 = ~n21513 & ~n21519;
  assign n21786 = ~n21513 & n55734;
  assign n21787 = ~n55734 & ~n21519;
  assign n21788 = n21513 & ~n55734;
  assign n21789 = ~n55780 & ~n55781;
  assign n21790 = ~n21519 & ~n21784;
  assign n21791 = ~n21783 & ~n55782;
  assign n21792 = ~n21519 & ~n21791;
  assign n21793 = n21495 & ~n21497;
  assign n21794 = ~n21495 & ~n21498;
  assign n21795 = ~n21495 & ~n21497;
  assign n21796 = n21497 & ~n21498;
  assign n21797 = n21495 & n21497;
  assign n21798 = ~n55783 & ~n55784;
  assign n21799 = ~n21498 & ~n21793;
  assign n21800 = ~n21792 & ~n55785;
  assign n21801 = ~n21498 & ~n21800;
  assign n21802 = ~n21464 & n21479;
  assign n21803 = n21464 & ~n21480;
  assign n21804 = n21464 & n21479;
  assign n21805 = ~n21479 & ~n21480;
  assign n21806 = ~n21464 & ~n21479;
  assign n21807 = ~n55786 & ~n55787;
  assign n21808 = ~n21480 & ~n21802;
  assign n21809 = ~n21801 & ~n55788;
  assign n21810 = ~n21480 & ~n21809;
  assign n21811 = ~n21444 & n21461;
  assign n21812 = ~n21462 & ~n21811;
  assign n21813 = ~n21810 & n21812;
  assign n21814 = ~n21462 & ~n21813;
  assign n21815 = n21436 & n55723;
  assign n21816 = ~n21436 & ~n21442;
  assign n21817 = ~n21436 & n55723;
  assign n21818 = ~n55723 & ~n21442;
  assign n21819 = n21436 & ~n55723;
  assign n21820 = ~n55789 & ~n55790;
  assign n21821 = ~n21442 & ~n21815;
  assign n21822 = ~n21814 & ~n55791;
  assign n21823 = ~n21442 & ~n21822;
  assign n21824 = n21413 & n55719;
  assign n21825 = ~n21413 & ~n21421;
  assign n21826 = ~n55719 & ~n21421;
  assign n21827 = ~n21825 & ~n21826;
  assign n21828 = ~n21421 & ~n21824;
  assign n21829 = ~n21823 & ~n55792;
  assign n21830 = ~n21421 & ~n21829;
  assign n21831 = n21390 & n55713;
  assign n21832 = ~n21390 & ~n21398;
  assign n21833 = ~n55713 & ~n21398;
  assign n21834 = ~n21832 & ~n21833;
  assign n21835 = ~n21398 & ~n21831;
  assign n21836 = ~n21830 & ~n55793;
  assign n21837 = ~n21398 & ~n21836;
  assign n21838 = n21369 & n55707;
  assign n21839 = ~n21369 & ~n21375;
  assign n21840 = ~n21369 & n55707;
  assign n21841 = ~n55707 & ~n21375;
  assign n21842 = n21369 & ~n55707;
  assign n21843 = ~n55794 & ~n55795;
  assign n21844 = ~n21375 & ~n21838;
  assign n21845 = ~n21837 & ~n55796;
  assign n21846 = ~n21375 & ~n21845;
  assign n21847 = n21348 & n55703;
  assign n21848 = ~n21348 & ~n21354;
  assign n21849 = ~n21348 & n55703;
  assign n21850 = ~n55703 & ~n21354;
  assign n21851 = n21348 & ~n55703;
  assign n21852 = ~n55797 & ~n55798;
  assign n21853 = ~n21354 & ~n21847;
  assign n21854 = ~n21846 & ~n55799;
  assign n21855 = ~n21354 & ~n21854;
  assign n21856 = n21325 & n55699;
  assign n21857 = ~n21325 & ~n21333;
  assign n21858 = ~n55699 & ~n21333;
  assign n21859 = ~n21857 & ~n21858;
  assign n21860 = ~n21333 & ~n21856;
  assign n21861 = ~n21855 & ~n55800;
  assign n21862 = ~n21333 & ~n21861;
  assign n21863 = n21302 & n55693;
  assign n21864 = ~n21302 & ~n21310;
  assign n21865 = ~n55693 & ~n21310;
  assign n21866 = ~n21864 & ~n21865;
  assign n21867 = ~n21310 & ~n21863;
  assign n21868 = ~n21862 & ~n55801;
  assign n21869 = ~n21310 & ~n21868;
  assign n21870 = n21172 & ~n21174;
  assign n21871 = ~n21175 & ~n21870;
  assign n21872 = ~n21869 & n21871;
  assign n21873 = n12938 & n17265;
  assign n21874 = ~n53819 & n18588;
  assign n21875 = ~n53860 & n55041;
  assign n21876 = ~n53845 & n18556;
  assign n21877 = ~n21875 & ~n21876;
  assign n21878 = ~n21874 & ~n21875;
  assign n21879 = ~n21876 & n21878;
  assign n21880 = ~n21874 & n21877;
  assign n21881 = ~n21873 & n55802;
  assign n21882 = pi14  & ~n21881;
  assign n21883 = ~n21881 & ~n21882;
  assign n21884 = ~pi14  & ~n21881;
  assign n21885 = pi14  & ~n21882;
  assign n21886 = pi14  & n21881;
  assign n21887 = ~n55803 & ~n55804;
  assign n21888 = n21869 & ~n21871;
  assign n21889 = ~n21872 & ~n21888;
  assign n21890 = ~n21887 & n21889;
  assign n21891 = ~n21872 & ~n21890;
  assign n21892 = n21200 & ~n21202;
  assign n21893 = n21202 & ~n21203;
  assign n21894 = ~n21200 & ~n21203;
  assign n21895 = ~n21893 & ~n21894;
  assign n21896 = ~n21203 & ~n21892;
  assign n21897 = ~n21891 & ~n55805;
  assign n21898 = n21891 & n55805;
  assign n21899 = n11889 & n18846;
  assign n21900 = ~n53712 & n19541;
  assign n21901 = ~n53774 & n55247;
  assign n21902 = ~n53741 & n19509;
  assign n21903 = ~n21901 & ~n21902;
  assign n21904 = ~n21900 & ~n21901;
  assign n21905 = ~n21902 & n21904;
  assign n21906 = ~n21900 & n21903;
  assign n21907 = ~n21899 & n55806;
  assign n21908 = pi11  & ~n21907;
  assign n21909 = pi11  & ~n21908;
  assign n21910 = pi11  & n21907;
  assign n21911 = ~n21907 & ~n21908;
  assign n21912 = ~pi11  & ~n21907;
  assign n21913 = ~n55807 & ~n55808;
  assign n21914 = ~n21898 & ~n21913;
  assign n21915 = ~n21897 & ~n21898;
  assign n21916 = ~n21913 & n21915;
  assign n21917 = ~n21897 & ~n21916;
  assign n21918 = ~n21897 & ~n21914;
  assign n21919 = ~n55687 & ~n55809;
  assign n21920 = n55687 & n55809;
  assign n21921 = n11286 & n20085;
  assign n21922 = ~n53650 & n21237;
  assign n21923 = ~n53657 & n55472;
  assign n21924 = ~n53634 & n21269;
  assign n21925 = ~n21923 & ~n21924;
  assign n21926 = ~n21922 & ~n21923;
  assign n21927 = ~n21924 & n21926;
  assign n21928 = ~n21922 & n21925;
  assign n21929 = ~n21921 & n55810;
  assign n21930 = pi8  & ~n21929;
  assign n21931 = pi8  & ~n21930;
  assign n21932 = pi8  & n21929;
  assign n21933 = ~n21929 & ~n21930;
  assign n21934 = ~pi8  & ~n21929;
  assign n21935 = ~n55811 & ~n55812;
  assign n21936 = ~n21920 & ~n21935;
  assign n21937 = ~n21919 & ~n21920;
  assign n21938 = ~n21935 & n21937;
  assign n21939 = ~n21919 & ~n21938;
  assign n21940 = ~n21919 & ~n21936;
  assign n21941 = ~n21282 & ~n55813;
  assign n21942 = ~n21230 & ~n21232;
  assign n21943 = ~n21233 & ~n21942;
  assign n21944 = n21282 & n55813;
  assign n21945 = ~n55813 & ~n21941;
  assign n21946 = n21282 & ~n55813;
  assign n21947 = ~n21282 & ~n21941;
  assign n21948 = ~n21282 & n55813;
  assign n21949 = ~n55814 & ~n55815;
  assign n21950 = ~n21941 & ~n21944;
  assign n21951 = n21943 & ~n55816;
  assign n21952 = ~n21941 & ~n21951;
  assign n21953 = ~n21249 & ~n55683;
  assign n21954 = ~n21257 & ~n21953;
  assign n21955 = ~n21952 & n21954;
  assign n21956 = ~n21943 & ~n55815;
  assign n21957 = ~n55814 & n21956;
  assign n21958 = ~n21943 & ~n55814;
  assign n21959 = ~n55815 & n21958;
  assign n21960 = ~n21943 & n55816;
  assign n21961 = ~n21951 & ~n55817;
  assign n21962 = ~n53439 & n53440;
  assign n21963 = pi3  & ~pi4 ;
  assign n21964 = ~pi3  & pi4 ;
  assign n21965 = ~pi3  & ~pi4 ;
  assign n21966 = pi3  & pi4 ;
  assign n21967 = ~n21965 & ~n21966;
  assign n21968 = ~n21963 & ~n21964;
  assign n21969 = n21962 & ~n55818;
  assign n21970 = n77 & ~n10547;
  assign n21971 = ~n21969 & ~n21970;
  assign n21972 = ~n2325 & n21969;
  assign n21973 = ~n10551 & ~n21972;
  assign n21974 = ~n77 & ~n21972;
  assign n21975 = ~n21973 & ~n21974;
  assign n21976 = ~n2325 & ~n21971;
  assign n21977 = pi5  & ~n55819;
  assign n21978 = ~pi5  & n55819;
  assign n21979 = ~n21977 & ~n21978;
  assign n21980 = n21862 & n55801;
  assign n21981 = ~n21868 & ~n21980;
  assign n21982 = n12918 & n17265;
  assign n21983 = ~n53860 & n18556;
  assign n21984 = ~n53888 & n55041;
  assign n21985 = ~n53845 & n18588;
  assign n21986 = ~n21984 & ~n21985;
  assign n21987 = ~n21983 & ~n21984;
  assign n21988 = ~n21985 & n21987;
  assign n21989 = ~n21983 & n21986;
  assign n21990 = ~n17265 & n55820;
  assign n21991 = ~n12918 & n55820;
  assign n21992 = ~n21990 & ~n21991;
  assign n21993 = ~n21982 & n55820;
  assign n21994 = pi14  & ~n55821;
  assign n21995 = ~pi14  & n55821;
  assign n21996 = ~n21994 & ~n21995;
  assign n21997 = n21981 & ~n21996;
  assign n21998 = n21855 & n55800;
  assign n21999 = ~n21861 & ~n21998;
  assign n22000 = n13336 & n17265;
  assign n22001 = ~n53888 & n18556;
  assign n22002 = ~n53907 & n55041;
  assign n22003 = ~n53860 & n18588;
  assign n22004 = ~n22002 & ~n22003;
  assign n22005 = ~n22001 & ~n22002;
  assign n22006 = ~n22003 & n22005;
  assign n22007 = ~n22001 & n22004;
  assign n22008 = ~n17265 & n55822;
  assign n22009 = ~n13336 & n55822;
  assign n22010 = ~n22008 & ~n22009;
  assign n22011 = ~n22000 & n55822;
  assign n22012 = pi14  & ~n55823;
  assign n22013 = ~pi14  & n55823;
  assign n22014 = ~n22012 & ~n22013;
  assign n22015 = n21999 & ~n22014;
  assign n22016 = n21846 & n55799;
  assign n22017 = ~n21854 & ~n22016;
  assign n22018 = n13360 & n17265;
  assign n22019 = ~n53907 & n18556;
  assign n22020 = ~n53930 & n55041;
  assign n22021 = ~n53888 & n18588;
  assign n22022 = ~n22020 & ~n22021;
  assign n22023 = ~n22019 & ~n22020;
  assign n22024 = ~n22021 & n22023;
  assign n22025 = ~n22019 & n22022;
  assign n22026 = ~n17265 & n55824;
  assign n22027 = ~n13360 & n55824;
  assign n22028 = ~n22026 & ~n22027;
  assign n22029 = ~n22018 & n55824;
  assign n22030 = pi14  & ~n55825;
  assign n22031 = ~pi14  & n55825;
  assign n22032 = ~n22030 & ~n22031;
  assign n22033 = n22017 & ~n22032;
  assign n22034 = n21837 & n55796;
  assign n22035 = ~n21845 & ~n22034;
  assign n22036 = n14263 & n17265;
  assign n22037 = ~n53930 & n18556;
  assign n22038 = ~n53962 & n55041;
  assign n22039 = ~n53907 & n18588;
  assign n22040 = ~n22038 & ~n22039;
  assign n22041 = ~n22037 & ~n22038;
  assign n22042 = ~n22039 & n22041;
  assign n22043 = ~n22037 & n22040;
  assign n22044 = ~n17265 & n55826;
  assign n22045 = ~n14263 & n55826;
  assign n22046 = ~n22044 & ~n22045;
  assign n22047 = ~n22036 & n55826;
  assign n22048 = pi14  & ~n55827;
  assign n22049 = ~pi14  & n55827;
  assign n22050 = ~n22048 & ~n22049;
  assign n22051 = n22035 & ~n22050;
  assign n22052 = n21830 & n55793;
  assign n22053 = ~n21836 & ~n22052;
  assign n22054 = n14020 & n17265;
  assign n22055 = ~n53962 & n18556;
  assign n22056 = ~n53970 & n55041;
  assign n22057 = ~n53930 & n18588;
  assign n22058 = ~n22056 & ~n22057;
  assign n22059 = ~n22055 & ~n22056;
  assign n22060 = ~n22057 & n22059;
  assign n22061 = ~n22055 & n22058;
  assign n22062 = ~n17265 & n55828;
  assign n22063 = ~n14020 & n55828;
  assign n22064 = ~n22062 & ~n22063;
  assign n22065 = ~n22054 & n55828;
  assign n22066 = pi14  & ~n55829;
  assign n22067 = ~pi14  & n55829;
  assign n22068 = ~n22066 & ~n22067;
  assign n22069 = n22053 & ~n22068;
  assign n22070 = n21823 & n55792;
  assign n22071 = ~n21829 & ~n22070;
  assign n22072 = n14708 & n17265;
  assign n22073 = ~n54005 & n55041;
  assign n22074 = ~n53970 & n18556;
  assign n22075 = ~n53962 & n18588;
  assign n22076 = ~n22074 & ~n22075;
  assign n22077 = ~n22073 & ~n22074;
  assign n22078 = ~n22075 & n22077;
  assign n22079 = ~n22073 & n22076;
  assign n22080 = ~n17265 & n55830;
  assign n22081 = ~n14708 & n55830;
  assign n22082 = ~n22080 & ~n22081;
  assign n22083 = ~n22072 & n55830;
  assign n22084 = pi14  & ~n55831;
  assign n22085 = ~pi14  & n55831;
  assign n22086 = ~n22084 & ~n22085;
  assign n22087 = n22071 & ~n22086;
  assign n22088 = n21814 & n55791;
  assign n22089 = ~n21822 & ~n22088;
  assign n22090 = n14688 & n17265;
  assign n22091 = ~n54005 & n18556;
  assign n22092 = ~n54034 & n55041;
  assign n22093 = ~n53970 & n18588;
  assign n22094 = ~n22092 & ~n22093;
  assign n22095 = ~n22091 & ~n22092;
  assign n22096 = ~n22093 & n22095;
  assign n22097 = ~n22091 & n22094;
  assign n22098 = ~n17265 & n55832;
  assign n22099 = ~n14688 & n55832;
  assign n22100 = ~n22098 & ~n22099;
  assign n22101 = ~n22090 & n55832;
  assign n22102 = pi14  & ~n55833;
  assign n22103 = ~pi14  & n55833;
  assign n22104 = ~n22102 & ~n22103;
  assign n22105 = n22089 & ~n22104;
  assign n22106 = n15195 & n17265;
  assign n22107 = ~n54050 & n55041;
  assign n22108 = ~n54005 & n18588;
  assign n22109 = ~n54034 & n18556;
  assign n22110 = ~n22108 & ~n22109;
  assign n22111 = ~n22107 & ~n22109;
  assign n22112 = ~n22108 & n22111;
  assign n22113 = ~n22107 & n22110;
  assign n22114 = ~n22106 & n55834;
  assign n22115 = pi14  & ~n22114;
  assign n22116 = ~n22114 & ~n22115;
  assign n22117 = ~pi14  & ~n22114;
  assign n22118 = pi14  & ~n22115;
  assign n22119 = pi14  & n22114;
  assign n22120 = ~n55835 & ~n55836;
  assign n22121 = n21810 & ~n21812;
  assign n22122 = ~n21813 & ~n22121;
  assign n22123 = ~n22120 & n22122;
  assign n22124 = n15219 & n17265;
  assign n22125 = ~n54050 & n18556;
  assign n22126 = ~n54034 & n18588;
  assign n22127 = ~n54073 & n55041;
  assign n22128 = ~n22126 & ~n22127;
  assign n22129 = ~n22125 & ~n22127;
  assign n22130 = ~n22126 & n22129;
  assign n22131 = ~n22125 & n22128;
  assign n22132 = ~n22124 & n55837;
  assign n22133 = pi14  & ~n22132;
  assign n22134 = ~n22132 & ~n22133;
  assign n22135 = ~pi14  & ~n22132;
  assign n22136 = pi14  & ~n22133;
  assign n22137 = pi14  & n22132;
  assign n22138 = ~n55838 & ~n55839;
  assign n22139 = n21801 & n55788;
  assign n22140 = ~n21801 & ~n21809;
  assign n22141 = ~n55788 & ~n21809;
  assign n22142 = ~n22140 & ~n22141;
  assign n22143 = ~n21809 & ~n22139;
  assign n22144 = ~n22138 & ~n55840;
  assign n22145 = n21792 & n55785;
  assign n22146 = ~n21800 & ~n22145;
  assign n22147 = n16138 & n17265;
  assign n22148 = ~n54098 & n55041;
  assign n22149 = ~n54050 & n18588;
  assign n22150 = ~n54073 & n18556;
  assign n22151 = ~n22149 & ~n22150;
  assign n22152 = ~n22148 & ~n22150;
  assign n22153 = ~n22149 & n22152;
  assign n22154 = ~n22148 & n22151;
  assign n22155 = ~n17265 & n55841;
  assign n22156 = ~n16138 & n55841;
  assign n22157 = ~n22155 & ~n22156;
  assign n22158 = ~n22147 & n55841;
  assign n22159 = pi14  & ~n55842;
  assign n22160 = ~pi14  & n55842;
  assign n22161 = ~n22159 & ~n22160;
  assign n22162 = n22146 & ~n22161;
  assign n22163 = n21783 & n55782;
  assign n22164 = ~n21791 & ~n22163;
  assign n22165 = n15779 & n17265;
  assign n22166 = ~n54098 & n18556;
  assign n22167 = ~n54119 & n55041;
  assign n22168 = ~n54073 & n18588;
  assign n22169 = ~n22167 & ~n22168;
  assign n22170 = ~n22166 & ~n22167;
  assign n22171 = ~n22168 & n22170;
  assign n22172 = ~n22166 & ~n22168;
  assign n22173 = ~n22167 & n22172;
  assign n22174 = ~n22166 & n22169;
  assign n22175 = ~n17265 & n55843;
  assign n22176 = ~n15779 & n55843;
  assign n22177 = ~n22175 & ~n22176;
  assign n22178 = ~n22165 & n55843;
  assign n22179 = pi14  & ~n55844;
  assign n22180 = ~pi14  & n55844;
  assign n22181 = ~n22179 & ~n22180;
  assign n22182 = n22164 & ~n22181;
  assign n22183 = n21776 & n55779;
  assign n22184 = ~n21782 & ~n22183;
  assign n22185 = n16547 & n17265;
  assign n22186 = ~n54119 & n18556;
  assign n22187 = ~n54098 & n18588;
  assign n22188 = ~n54132 & n55041;
  assign n22189 = ~n22187 & ~n22188;
  assign n22190 = ~n22186 & ~n22188;
  assign n22191 = ~n22187 & n22190;
  assign n22192 = ~n22186 & n22189;
  assign n22193 = ~n17265 & n55845;
  assign n22194 = ~n16547 & n55845;
  assign n22195 = ~n22193 & ~n22194;
  assign n22196 = ~n22185 & n55845;
  assign n22197 = pi14  & ~n55846;
  assign n22198 = ~pi14  & n55846;
  assign n22199 = ~n22197 & ~n22198;
  assign n22200 = n22184 & ~n22199;
  assign n22201 = n16772 & n17265;
  assign n22202 = ~n54154 & n55041;
  assign n22203 = ~n54119 & n18588;
  assign n22204 = ~n54132 & n18556;
  assign n22205 = ~n22203 & ~n22204;
  assign n22206 = ~n22202 & ~n22204;
  assign n22207 = ~n22203 & n22206;
  assign n22208 = ~n22202 & n22205;
  assign n22209 = ~n22201 & n55847;
  assign n22210 = pi14  & ~n22209;
  assign n22211 = ~n22209 & ~n22210;
  assign n22212 = ~pi14  & ~n22209;
  assign n22213 = pi14  & ~n22210;
  assign n22214 = pi14  & n22209;
  assign n22215 = ~n55848 & ~n55849;
  assign n22216 = n21772 & ~n21774;
  assign n22217 = ~n21775 & ~n22216;
  assign n22218 = ~n22215 & n22217;
  assign n22219 = n16522 & n17265;
  assign n22220 = ~n54154 & n18556;
  assign n22221 = ~n54132 & n18588;
  assign n22222 = ~n54163 & n55041;
  assign n22223 = ~n22221 & ~n22222;
  assign n22224 = ~n22220 & ~n22222;
  assign n22225 = ~n22221 & n22224;
  assign n22226 = ~n22220 & n22223;
  assign n22227 = ~n22219 & n55850;
  assign n22228 = pi14  & ~n22227;
  assign n22229 = ~n22227 & ~n22228;
  assign n22230 = ~pi14  & ~n22227;
  assign n22231 = pi14  & ~n22228;
  assign n22232 = pi14  & n22227;
  assign n22233 = ~n55851 & ~n55852;
  assign n22234 = n21763 & n55778;
  assign n22235 = ~n21763 & ~n21771;
  assign n22236 = ~n55778 & ~n21771;
  assign n22237 = ~n22235 & ~n22236;
  assign n22238 = ~n21771 & ~n22234;
  assign n22239 = ~n22233 & ~n55853;
  assign n22240 = n17072 & n17265;
  assign n22241 = ~n54154 & n18588;
  assign n22242 = ~n54183 & n55041;
  assign n22243 = ~n54163 & n18556;
  assign n22244 = ~n22242 & ~n22243;
  assign n22245 = ~n22241 & n22244;
  assign n22246 = ~n22240 & n22245;
  assign n22247 = pi14  & ~n22246;
  assign n22248 = ~n22246 & ~n22247;
  assign n22249 = ~pi14  & ~n22246;
  assign n22250 = pi14  & ~n22247;
  assign n22251 = pi14  & n22246;
  assign n22252 = ~n55854 & ~n55855;
  assign n22253 = n21754 & n55775;
  assign n22254 = ~n21754 & ~n21762;
  assign n22255 = ~n21754 & n55775;
  assign n22256 = ~n55775 & ~n21762;
  assign n22257 = n21754 & ~n55775;
  assign n22258 = ~n55856 & ~n55857;
  assign n22259 = ~n21762 & ~n22253;
  assign n22260 = ~n22252 & ~n55858;
  assign n22261 = n21745 & n55772;
  assign n22262 = ~n21753 & ~n22261;
  assign n22263 = n17265 & n17524;
  assign n22264 = ~n54183 & n18556;
  assign n22265 = ~n54194 & n55041;
  assign n22266 = ~n54163 & n18588;
  assign n22267 = ~n22265 & ~n22266;
  assign n22268 = ~n22264 & ~n22265;
  assign n22269 = ~n22266 & n22268;
  assign n22270 = ~n22264 & n22267;
  assign n22271 = ~n17265 & n55859;
  assign n22272 = ~n17524 & n55859;
  assign n22273 = ~n22271 & ~n22272;
  assign n22274 = ~n22263 & n55859;
  assign n22275 = pi14  & ~n55860;
  assign n22276 = ~pi14  & n55860;
  assign n22277 = ~n22275 & ~n22276;
  assign n22278 = n22262 & ~n22277;
  assign n22279 = n21741 & ~n21743;
  assign n22280 = ~n21744 & ~n22279;
  assign n22281 = n17265 & n17544;
  assign n22282 = ~n54212 & n55041;
  assign n22283 = ~n54183 & n18588;
  assign n22284 = ~n54194 & n18556;
  assign n22285 = ~n22283 & ~n22284;
  assign n22286 = ~n22282 & ~n22284;
  assign n22287 = ~n22283 & n22286;
  assign n22288 = ~n22282 & n22285;
  assign n22289 = ~n17265 & n55861;
  assign n22290 = ~n17544 & n55861;
  assign n22291 = ~n22289 & ~n22290;
  assign n22292 = ~n22281 & n55861;
  assign n22293 = pi14  & ~n55862;
  assign n22294 = ~pi14  & n55862;
  assign n22295 = ~n22293 & ~n22294;
  assign n22296 = n22280 & ~n22295;
  assign n22297 = n21732 & n55769;
  assign n22298 = ~n21740 & ~n22297;
  assign n22299 = n17041 & n17265;
  assign n22300 = ~n54212 & n18556;
  assign n22301 = ~n54194 & n18588;
  assign n22302 = ~n54240 & n55041;
  assign n22303 = ~n22301 & ~n22302;
  assign n22304 = ~n22300 & ~n22302;
  assign n22305 = ~n22301 & n22304;
  assign n22306 = ~n22300 & n22303;
  assign n22307 = ~n17265 & n55863;
  assign n22308 = ~n17041 & n55863;
  assign n22309 = ~n22307 & ~n22308;
  assign n22310 = ~n22299 & n55863;
  assign n22311 = pi14  & ~n55864;
  assign n22312 = ~pi14  & n55864;
  assign n22313 = ~n22311 & ~n22312;
  assign n22314 = n22298 & ~n22313;
  assign n22315 = n17265 & n17660;
  assign n22316 = ~n54254 & n55041;
  assign n22317 = ~n54212 & n18588;
  assign n22318 = ~n54240 & n18556;
  assign n22319 = ~n22317 & ~n22318;
  assign n22320 = ~n22316 & ~n22318;
  assign n22321 = ~n22317 & n22320;
  assign n22322 = ~n22316 & n22319;
  assign n22323 = ~n22315 & n55865;
  assign n22324 = pi14  & ~n22323;
  assign n22325 = ~n22323 & ~n22324;
  assign n22326 = ~pi14  & ~n22323;
  assign n22327 = pi14  & ~n22324;
  assign n22328 = pi14  & n22323;
  assign n22329 = ~n55866 & ~n55867;
  assign n22330 = n21728 & ~n21730;
  assign n22331 = ~n21731 & ~n22330;
  assign n22332 = ~n22329 & n22331;
  assign n22333 = n17265 & n17804;
  assign n22334 = ~n54254 & n18556;
  assign n22335 = ~n54240 & n18588;
  assign n22336 = ~n54269 & n55041;
  assign n22337 = ~n22335 & ~n22336;
  assign n22338 = ~n22334 & ~n22336;
  assign n22339 = ~n22335 & n22338;
  assign n22340 = ~n22334 & n22337;
  assign n22341 = ~n17265 & n55868;
  assign n22342 = ~n17804 & n55868;
  assign n22343 = ~n22341 & ~n22342;
  assign n22344 = ~n22333 & n55868;
  assign n22345 = pi14  & ~n55869;
  assign n22346 = ~pi14  & n55869;
  assign n22347 = ~n22345 & ~n22346;
  assign n22348 = n21719 & n55766;
  assign n22349 = ~n55766 & ~n21727;
  assign n22350 = ~n21719 & ~n21727;
  assign n22351 = ~n22349 & ~n22350;
  assign n22352 = ~n21727 & ~n22348;
  assign n22353 = ~n22347 & ~n55870;
  assign n22354 = n17265 & n17939;
  assign n22355 = ~n54254 & n18588;
  assign n22356 = ~n54277 & n55041;
  assign n22357 = ~n54269 & n18556;
  assign n22358 = ~n22356 & ~n22357;
  assign n22359 = ~n22355 & n22358;
  assign n22360 = ~n22354 & n22359;
  assign n22361 = pi14  & ~n22360;
  assign n22362 = ~n22360 & ~n22361;
  assign n22363 = ~pi14  & ~n22360;
  assign n22364 = pi14  & ~n22361;
  assign n22365 = pi14  & n22360;
  assign n22366 = ~n55871 & ~n55872;
  assign n22367 = pi17  & ~n55758;
  assign n22368 = ~n55759 & ~n22367;
  assign n22369 = n55759 & n22367;
  assign n22370 = ~n55758 & n21701;
  assign n22371 = ~n55760 & ~n22370;
  assign n22372 = ~n22368 & ~n22369;
  assign n22373 = ~n22366 & n55873;
  assign n22374 = n17265 & n18056;
  assign n22375 = ~n54305 & n55041;
  assign n22376 = ~n54277 & n18556;
  assign n22377 = ~n54269 & n18588;
  assign n22378 = ~n22376 & ~n22377;
  assign n22379 = ~n22375 & ~n22376;
  assign n22380 = ~n22377 & n22379;
  assign n22381 = ~n22375 & n22378;
  assign n22382 = ~n17265 & n55874;
  assign n22383 = ~n18056 & n55874;
  assign n22384 = ~n22382 & ~n22383;
  assign n22385 = ~n22374 & n55874;
  assign n22386 = pi14  & ~n55875;
  assign n22387 = ~pi14  & n55875;
  assign n22388 = ~n22386 & ~n22387;
  assign n22389 = pi17  & n21681;
  assign n22390 = ~n21680 & n22389;
  assign n22391 = n21680 & ~n22389;
  assign n22392 = ~n21682 & n21686;
  assign n22393 = ~n55758 & ~n22392;
  assign n22394 = ~n22390 & ~n22391;
  assign n22395 = ~n22388 & n55876;
  assign n22396 = n17265 & ~n19275;
  assign n22397 = ~n54325 & n18556;
  assign n22398 = ~n54344 & n18588;
  assign n22399 = ~n22397 & ~n22398;
  assign n22400 = ~n22396 & n22399;
  assign n22401 = ~n54325 & n55039;
  assign n22402 = pi14  & ~n22401;
  assign n22403 = pi14  & ~n22400;
  assign n22404 = pi14  & ~n22403;
  assign n22405 = ~n22400 & ~n22403;
  assign n22406 = ~n22404 & ~n22405;
  assign n22407 = n22402 & ~n22406;
  assign n22408 = n22400 & n22402;
  assign n22409 = n17265 & n18156;
  assign n22410 = ~n54305 & n18588;
  assign n22411 = ~n54325 & n55041;
  assign n22412 = ~n54344 & n18556;
  assign n22413 = ~n22411 & ~n22412;
  assign n22414 = ~n22410 & n22413;
  assign n22415 = ~n17265 & n22414;
  assign n22416 = ~n18156 & n22414;
  assign n22417 = ~n22415 & ~n22416;
  assign n22418 = ~n22409 & n22414;
  assign n22419 = pi14  & ~n55878;
  assign n22420 = ~pi14  & n55878;
  assign n22421 = ~n22419 & ~n22420;
  assign n22422 = n55877 & ~n22421;
  assign n22423 = n55877 & ~n55878;
  assign n22424 = n21681 & n55879;
  assign n22425 = n17265 & n18336;
  assign n22426 = ~n54305 & n18556;
  assign n22427 = ~n54277 & n18588;
  assign n22428 = ~n54344 & n55041;
  assign n22429 = ~n22427 & ~n22428;
  assign n22430 = ~n22426 & ~n22428;
  assign n22431 = ~n22427 & n22430;
  assign n22432 = ~n22426 & n22429;
  assign n22433 = ~n22425 & n55880;
  assign n22434 = pi14  & ~n22433;
  assign n22435 = pi14  & ~n22434;
  assign n22436 = pi14  & n22433;
  assign n22437 = ~n22433 & ~n22434;
  assign n22438 = ~pi14  & ~n22433;
  assign n22439 = ~n55881 & ~n55882;
  assign n22440 = ~n21681 & ~n55879;
  assign n22441 = n55879 & ~n22424;
  assign n22442 = ~n21681 & n55879;
  assign n22443 = n21681 & ~n22424;
  assign n22444 = n21681 & ~n55879;
  assign n22445 = ~n55883 & ~n55884;
  assign n22446 = ~n22424 & ~n22440;
  assign n22447 = ~n22439 & ~n55885;
  assign n22448 = ~n22424 & ~n22447;
  assign n22449 = n22388 & ~n55876;
  assign n22450 = ~n22395 & ~n22449;
  assign n22451 = ~n22448 & n22450;
  assign n22452 = ~n22395 & ~n22451;
  assign n22453 = n22366 & ~n55873;
  assign n22454 = ~n22366 & ~n22373;
  assign n22455 = ~n22366 & ~n55873;
  assign n22456 = n55873 & ~n22373;
  assign n22457 = n22366 & n55873;
  assign n22458 = ~n55886 & ~n55887;
  assign n22459 = ~n22373 & ~n22453;
  assign n22460 = ~n22452 & ~n55888;
  assign n22461 = ~n22373 & ~n22460;
  assign n22462 = n22347 & n55870;
  assign n22463 = ~n22353 & ~n22462;
  assign n22464 = ~n22461 & n22463;
  assign n22465 = ~n22353 & ~n22464;
  assign n22466 = n22329 & ~n22331;
  assign n22467 = ~n22329 & ~n22332;
  assign n22468 = ~n22329 & ~n22331;
  assign n22469 = n22331 & ~n22332;
  assign n22470 = n22329 & n22331;
  assign n22471 = ~n55889 & ~n55890;
  assign n22472 = ~n22332 & ~n22466;
  assign n22473 = ~n22465 & ~n55891;
  assign n22474 = ~n22332 & ~n22473;
  assign n22475 = ~n22298 & n22313;
  assign n22476 = n22298 & ~n22314;
  assign n22477 = n22298 & n22313;
  assign n22478 = ~n22313 & ~n22314;
  assign n22479 = ~n22298 & ~n22313;
  assign n22480 = ~n55892 & ~n55893;
  assign n22481 = ~n22314 & ~n22475;
  assign n22482 = ~n22474 & ~n55894;
  assign n22483 = ~n22314 & ~n22482;
  assign n22484 = ~n22280 & n22295;
  assign n22485 = n22280 & ~n22296;
  assign n22486 = n22280 & n22295;
  assign n22487 = ~n22295 & ~n22296;
  assign n22488 = ~n22280 & ~n22295;
  assign n22489 = ~n55895 & ~n55896;
  assign n22490 = ~n22296 & ~n22484;
  assign n22491 = ~n22483 & ~n55897;
  assign n22492 = ~n22296 & ~n22491;
  assign n22493 = ~n22262 & n22277;
  assign n22494 = ~n22278 & ~n22493;
  assign n22495 = ~n22492 & n22494;
  assign n22496 = ~n22278 & ~n22495;
  assign n22497 = n22252 & n55858;
  assign n22498 = ~n22252 & ~n22260;
  assign n22499 = ~n55858 & ~n22260;
  assign n22500 = ~n22498 & ~n22499;
  assign n22501 = ~n22260 & ~n22497;
  assign n22502 = ~n22496 & ~n55898;
  assign n22503 = ~n22260 & ~n22502;
  assign n22504 = n22233 & n55853;
  assign n22505 = ~n22233 & ~n22239;
  assign n22506 = ~n22233 & n55853;
  assign n22507 = ~n55853 & ~n22239;
  assign n22508 = n22233 & ~n55853;
  assign n22509 = ~n55899 & ~n55900;
  assign n22510 = ~n22239 & ~n22504;
  assign n22511 = ~n22503 & ~n55901;
  assign n22512 = ~n22239 & ~n22511;
  assign n22513 = n22215 & ~n22217;
  assign n22514 = ~n22215 & ~n22218;
  assign n22515 = ~n22215 & ~n22217;
  assign n22516 = n22217 & ~n22218;
  assign n22517 = n22215 & n22217;
  assign n22518 = ~n55902 & ~n55903;
  assign n22519 = ~n22218 & ~n22513;
  assign n22520 = ~n22512 & ~n55904;
  assign n22521 = ~n22218 & ~n22520;
  assign n22522 = ~n22184 & n22199;
  assign n22523 = n22184 & ~n22200;
  assign n22524 = n22184 & n22199;
  assign n22525 = ~n22199 & ~n22200;
  assign n22526 = ~n22184 & ~n22199;
  assign n22527 = ~n55905 & ~n55906;
  assign n22528 = ~n22200 & ~n22522;
  assign n22529 = ~n22521 & ~n55907;
  assign n22530 = ~n22200 & ~n22529;
  assign n22531 = ~n22164 & n22181;
  assign n22532 = n22164 & ~n22182;
  assign n22533 = n22164 & n22181;
  assign n22534 = ~n22181 & ~n22182;
  assign n22535 = ~n22164 & ~n22181;
  assign n22536 = ~n55908 & ~n55909;
  assign n22537 = ~n22182 & ~n22531;
  assign n22538 = ~n22530 & ~n55910;
  assign n22539 = ~n22182 & ~n22538;
  assign n22540 = ~n22146 & n22161;
  assign n22541 = ~n22162 & ~n22540;
  assign n22542 = ~n22539 & n22541;
  assign n22543 = ~n22162 & ~n22542;
  assign n22544 = n22138 & n55840;
  assign n22545 = ~n22138 & ~n22144;
  assign n22546 = ~n22138 & n55840;
  assign n22547 = ~n55840 & ~n22144;
  assign n22548 = n22138 & ~n55840;
  assign n22549 = ~n55911 & ~n55912;
  assign n22550 = ~n22144 & ~n22544;
  assign n22551 = ~n22543 & ~n55913;
  assign n22552 = ~n22144 & ~n22551;
  assign n22553 = n22120 & ~n22122;
  assign n22554 = ~n22120 & ~n22123;
  assign n22555 = ~n22120 & ~n22122;
  assign n22556 = n22122 & ~n22123;
  assign n22557 = n22120 & n22122;
  assign n22558 = ~n55914 & ~n55915;
  assign n22559 = ~n22123 & ~n22553;
  assign n22560 = ~n22552 & ~n55916;
  assign n22561 = ~n22123 & ~n22560;
  assign n22562 = ~n22089 & n22104;
  assign n22563 = n22089 & ~n22105;
  assign n22564 = n22089 & n22104;
  assign n22565 = ~n22104 & ~n22105;
  assign n22566 = ~n22089 & ~n22104;
  assign n22567 = ~n55917 & ~n55918;
  assign n22568 = ~n22105 & ~n22562;
  assign n22569 = ~n22561 & ~n55919;
  assign n22570 = ~n22105 & ~n22569;
  assign n22571 = ~n22071 & n22086;
  assign n22572 = n22071 & ~n22087;
  assign n22573 = n22071 & n22086;
  assign n22574 = ~n22086 & ~n22087;
  assign n22575 = ~n22071 & ~n22086;
  assign n22576 = ~n55920 & ~n55921;
  assign n22577 = ~n22087 & ~n22571;
  assign n22578 = ~n22570 & ~n55922;
  assign n22579 = ~n22087 & ~n22578;
  assign n22580 = ~n22053 & n22068;
  assign n22581 = n22053 & ~n22069;
  assign n22582 = n22053 & n22068;
  assign n22583 = ~n22068 & ~n22069;
  assign n22584 = ~n22053 & ~n22068;
  assign n22585 = ~n55923 & ~n55924;
  assign n22586 = ~n22069 & ~n22580;
  assign n22587 = ~n22579 & ~n55925;
  assign n22588 = ~n22069 & ~n22587;
  assign n22589 = ~n22035 & n22050;
  assign n22590 = n22035 & ~n22051;
  assign n22591 = n22035 & n22050;
  assign n22592 = ~n22050 & ~n22051;
  assign n22593 = ~n22035 & ~n22050;
  assign n22594 = ~n55926 & ~n55927;
  assign n22595 = ~n22051 & ~n22589;
  assign n22596 = ~n22588 & ~n55928;
  assign n22597 = ~n22051 & ~n22596;
  assign n22598 = ~n22017 & n22032;
  assign n22599 = n22017 & ~n22033;
  assign n22600 = n22017 & n22032;
  assign n22601 = ~n22032 & ~n22033;
  assign n22602 = ~n22017 & ~n22032;
  assign n22603 = ~n55929 & ~n55930;
  assign n22604 = ~n22033 & ~n22598;
  assign n22605 = ~n22597 & ~n55931;
  assign n22606 = ~n22033 & ~n22605;
  assign n22607 = ~n21999 & n22014;
  assign n22608 = n21999 & ~n22015;
  assign n22609 = n21999 & n22014;
  assign n22610 = ~n22014 & ~n22015;
  assign n22611 = ~n21999 & ~n22014;
  assign n22612 = ~n55932 & ~n55933;
  assign n22613 = ~n22015 & ~n22607;
  assign n22614 = ~n22606 & ~n55934;
  assign n22615 = ~n22015 & ~n22614;
  assign n22616 = ~n21981 & n21996;
  assign n22617 = n21981 & ~n21997;
  assign n22618 = n21981 & n21996;
  assign n22619 = ~n21996 & ~n21997;
  assign n22620 = ~n21981 & ~n21996;
  assign n22621 = ~n55935 & ~n55936;
  assign n22622 = ~n21997 & ~n22616;
  assign n22623 = ~n22615 & ~n55937;
  assign n22624 = ~n21997 & ~n22623;
  assign n22625 = n21887 & ~n21889;
  assign n22626 = ~n21890 & ~n22625;
  assign n22627 = ~n22624 & n22626;
  assign n22628 = n11913 & n18846;
  assign n22629 = ~n53774 & n19509;
  assign n22630 = ~n53799 & n55247;
  assign n22631 = ~n53741 & n19541;
  assign n22632 = ~n22630 & ~n22631;
  assign n22633 = ~n22629 & ~n22630;
  assign n22634 = ~n22631 & n22633;
  assign n22635 = ~n22629 & n22632;
  assign n22636 = ~n22628 & n55938;
  assign n22637 = pi11  & ~n22636;
  assign n22638 = ~n22636 & ~n22637;
  assign n22639 = ~pi11  & ~n22636;
  assign n22640 = pi11  & ~n22637;
  assign n22641 = pi11  & n22636;
  assign n22642 = ~n55939 & ~n55940;
  assign n22643 = n22624 & ~n22626;
  assign n22644 = ~n22627 & ~n22643;
  assign n22645 = ~n22642 & n22644;
  assign n22646 = ~n22627 & ~n22645;
  assign n22647 = n21915 & ~n21916;
  assign n22648 = n21913 & n21915;
  assign n22649 = ~n21913 & ~n21916;
  assign n22650 = ~n21913 & ~n21915;
  assign n22651 = n21913 & ~n21915;
  assign n22652 = ~n21916 & ~n22651;
  assign n22653 = ~n55941 & ~n55942;
  assign n22654 = ~n22646 & n55943;
  assign n22655 = n22646 & ~n55943;
  assign n22656 = n11213 & n20085;
  assign n22657 = ~n53650 & n21269;
  assign n22658 = ~n53685 & n55472;
  assign n22659 = ~n53657 & n21237;
  assign n22660 = ~n22658 & ~n22659;
  assign n22661 = ~n22657 & n22660;
  assign n22662 = ~n22656 & n22661;
  assign n22663 = pi8  & ~n22662;
  assign n22664 = pi8  & ~n22663;
  assign n22665 = pi8  & n22662;
  assign n22666 = ~n22662 & ~n22663;
  assign n22667 = ~pi8  & ~n22662;
  assign n22668 = ~n55944 & ~n55945;
  assign n22669 = ~n22655 & ~n22668;
  assign n22670 = ~n22654 & ~n22655;
  assign n22671 = ~n22668 & n22670;
  assign n22672 = ~n22654 & ~n22671;
  assign n22673 = ~n22654 & ~n22669;
  assign n22674 = ~n21979 & ~n55946;
  assign n22675 = n21979 & n55946;
  assign n22676 = n21935 & ~n21937;
  assign n22677 = n21937 & ~n21938;
  assign n22678 = ~n21935 & ~n21938;
  assign n22679 = ~n22677 & ~n22678;
  assign n22680 = ~n21938 & ~n22676;
  assign n22681 = ~n22675 & ~n55947;
  assign n22682 = ~n22674 & ~n22675;
  assign n22683 = ~n55947 & n22682;
  assign n22684 = ~n22674 & ~n22683;
  assign n22685 = ~n22674 & ~n22681;
  assign n22686 = n21961 & ~n55948;
  assign n22687 = n12690 & n18846;
  assign n22688 = ~n53774 & n19541;
  assign n22689 = ~n53819 & n55247;
  assign n22690 = ~n53799 & n19509;
  assign n22691 = ~n22689 & ~n22690;
  assign n22692 = ~n22688 & ~n22689;
  assign n22693 = ~n22690 & n22692;
  assign n22694 = ~n22688 & n22691;
  assign n22695 = ~n22687 & n55949;
  assign n22696 = pi11  & ~n22695;
  assign n22697 = ~n22695 & ~n22696;
  assign n22698 = ~pi11  & ~n22695;
  assign n22699 = pi11  & ~n22696;
  assign n22700 = pi11  & n22695;
  assign n22701 = ~n55950 & ~n55951;
  assign n22702 = n22615 & n55937;
  assign n22703 = ~n22615 & ~n22623;
  assign n22704 = ~n55937 & ~n22623;
  assign n22705 = ~n22703 & ~n22704;
  assign n22706 = ~n22623 & ~n22702;
  assign n22707 = ~n22701 & ~n55952;
  assign n22708 = n12550 & n18846;
  assign n22709 = ~n53819 & n19509;
  assign n22710 = ~n53845 & n55247;
  assign n22711 = ~n53799 & n19541;
  assign n22712 = ~n22710 & ~n22711;
  assign n22713 = ~n22709 & ~n22710;
  assign n22714 = ~n22711 & n22713;
  assign n22715 = ~n22709 & n22712;
  assign n22716 = ~n22708 & n55953;
  assign n22717 = pi11  & ~n22716;
  assign n22718 = ~n22716 & ~n22717;
  assign n22719 = ~pi11  & ~n22716;
  assign n22720 = pi11  & ~n22717;
  assign n22721 = pi11  & n22716;
  assign n22722 = ~n55954 & ~n55955;
  assign n22723 = n22606 & n55934;
  assign n22724 = ~n22606 & ~n22614;
  assign n22725 = ~n55934 & ~n22614;
  assign n22726 = ~n22724 & ~n22725;
  assign n22727 = ~n22614 & ~n22723;
  assign n22728 = ~n22722 & ~n55956;
  assign n22729 = n12938 & n18846;
  assign n22730 = ~n53819 & n19541;
  assign n22731 = ~n53860 & n55247;
  assign n22732 = ~n53845 & n19509;
  assign n22733 = ~n22731 & ~n22732;
  assign n22734 = ~n22730 & ~n22731;
  assign n22735 = ~n22732 & n22734;
  assign n22736 = ~n22730 & n22733;
  assign n22737 = ~n22729 & n55957;
  assign n22738 = pi11  & ~n22737;
  assign n22739 = ~n22737 & ~n22738;
  assign n22740 = ~pi11  & ~n22737;
  assign n22741 = pi11  & ~n22738;
  assign n22742 = pi11  & n22737;
  assign n22743 = ~n55958 & ~n55959;
  assign n22744 = n22597 & n55931;
  assign n22745 = ~n22597 & ~n22605;
  assign n22746 = ~n22597 & n55931;
  assign n22747 = ~n55931 & ~n22605;
  assign n22748 = n22597 & ~n55931;
  assign n22749 = ~n55960 & ~n55961;
  assign n22750 = ~n22605 & ~n22744;
  assign n22751 = ~n22743 & ~n55962;
  assign n22752 = n12918 & n18846;
  assign n22753 = ~n53860 & n19509;
  assign n22754 = ~n53888 & n55247;
  assign n22755 = ~n53845 & n19541;
  assign n22756 = ~n22754 & ~n22755;
  assign n22757 = ~n22753 & ~n22754;
  assign n22758 = ~n22755 & n22757;
  assign n22759 = ~n22753 & n22756;
  assign n22760 = ~n22752 & n55963;
  assign n22761 = pi11  & ~n22760;
  assign n22762 = ~n22760 & ~n22761;
  assign n22763 = ~pi11  & ~n22760;
  assign n22764 = pi11  & ~n22761;
  assign n22765 = pi11  & n22760;
  assign n22766 = ~n55964 & ~n55965;
  assign n22767 = n22588 & n55928;
  assign n22768 = ~n22588 & ~n22596;
  assign n22769 = ~n22588 & n55928;
  assign n22770 = ~n55928 & ~n22596;
  assign n22771 = n22588 & ~n55928;
  assign n22772 = ~n55966 & ~n55967;
  assign n22773 = ~n22596 & ~n22767;
  assign n22774 = ~n22766 & ~n55968;
  assign n22775 = n13336 & n18846;
  assign n22776 = ~n53888 & n19509;
  assign n22777 = ~n53907 & n55247;
  assign n22778 = ~n53860 & n19541;
  assign n22779 = ~n22777 & ~n22778;
  assign n22780 = ~n22776 & ~n22777;
  assign n22781 = ~n22778 & n22780;
  assign n22782 = ~n22776 & n22779;
  assign n22783 = ~n22775 & n55969;
  assign n22784 = pi11  & ~n22783;
  assign n22785 = ~n22783 & ~n22784;
  assign n22786 = ~pi11  & ~n22783;
  assign n22787 = pi11  & ~n22784;
  assign n22788 = pi11  & n22783;
  assign n22789 = ~n55970 & ~n55971;
  assign n22790 = n22579 & n55925;
  assign n22791 = ~n22579 & ~n22587;
  assign n22792 = ~n55925 & ~n22587;
  assign n22793 = ~n22791 & ~n22792;
  assign n22794 = ~n22587 & ~n22790;
  assign n22795 = ~n22789 & ~n55972;
  assign n22796 = n13360 & n18846;
  assign n22797 = ~n53907 & n19509;
  assign n22798 = ~n53930 & n55247;
  assign n22799 = ~n53888 & n19541;
  assign n22800 = ~n22798 & ~n22799;
  assign n22801 = ~n22797 & ~n22798;
  assign n22802 = ~n22799 & n22801;
  assign n22803 = ~n22797 & n22800;
  assign n22804 = ~n22796 & n55973;
  assign n22805 = pi11  & ~n22804;
  assign n22806 = ~n22804 & ~n22805;
  assign n22807 = ~pi11  & ~n22804;
  assign n22808 = pi11  & ~n22805;
  assign n22809 = pi11  & n22804;
  assign n22810 = ~n55974 & ~n55975;
  assign n22811 = n22570 & n55922;
  assign n22812 = ~n22570 & ~n22578;
  assign n22813 = ~n55922 & ~n22578;
  assign n22814 = ~n22812 & ~n22813;
  assign n22815 = ~n22578 & ~n22811;
  assign n22816 = ~n22810 & ~n55976;
  assign n22817 = n14263 & n18846;
  assign n22818 = ~n53930 & n19509;
  assign n22819 = ~n53962 & n55247;
  assign n22820 = ~n53907 & n19541;
  assign n22821 = ~n22819 & ~n22820;
  assign n22822 = ~n22818 & ~n22819;
  assign n22823 = ~n22820 & n22822;
  assign n22824 = ~n22818 & n22821;
  assign n22825 = ~n22817 & n55977;
  assign n22826 = pi11  & ~n22825;
  assign n22827 = ~n22825 & ~n22826;
  assign n22828 = ~pi11  & ~n22825;
  assign n22829 = pi11  & ~n22826;
  assign n22830 = pi11  & n22825;
  assign n22831 = ~n55978 & ~n55979;
  assign n22832 = n22561 & n55919;
  assign n22833 = ~n22561 & ~n22569;
  assign n22834 = ~n22561 & n55919;
  assign n22835 = ~n55919 & ~n22569;
  assign n22836 = n22561 & ~n55919;
  assign n22837 = ~n55980 & ~n55981;
  assign n22838 = ~n22569 & ~n22832;
  assign n22839 = ~n22831 & ~n55982;
  assign n22840 = n22552 & n55916;
  assign n22841 = ~n22560 & ~n22840;
  assign n22842 = n14020 & n18846;
  assign n22843 = ~n53962 & n19509;
  assign n22844 = ~n53970 & n55247;
  assign n22845 = ~n53930 & n19541;
  assign n22846 = ~n22844 & ~n22845;
  assign n22847 = ~n22843 & ~n22844;
  assign n22848 = ~n22845 & n22847;
  assign n22849 = ~n22843 & n22846;
  assign n22850 = ~n18846 & n55983;
  assign n22851 = ~n14020 & n55983;
  assign n22852 = ~n22850 & ~n22851;
  assign n22853 = ~n22842 & n55983;
  assign n22854 = pi11  & ~n55984;
  assign n22855 = ~pi11  & n55984;
  assign n22856 = ~n22854 & ~n22855;
  assign n22857 = n22841 & ~n22856;
  assign n22858 = n22543 & n55913;
  assign n22859 = ~n22551 & ~n22858;
  assign n22860 = n14708 & n18846;
  assign n22861 = ~n54005 & n55247;
  assign n22862 = ~n53970 & n19509;
  assign n22863 = ~n53962 & n19541;
  assign n22864 = ~n22862 & ~n22863;
  assign n22865 = ~n22861 & ~n22862;
  assign n22866 = ~n22863 & n22865;
  assign n22867 = ~n22861 & n22864;
  assign n22868 = ~n18846 & n55985;
  assign n22869 = ~n14708 & n55985;
  assign n22870 = ~n22868 & ~n22869;
  assign n22871 = ~n22860 & n55985;
  assign n22872 = pi11  & ~n55986;
  assign n22873 = ~pi11  & n55986;
  assign n22874 = ~n22872 & ~n22873;
  assign n22875 = n22859 & ~n22874;
  assign n22876 = n14688 & n18846;
  assign n22877 = ~n54005 & n19509;
  assign n22878 = ~n54034 & n55247;
  assign n22879 = ~n53970 & n19541;
  assign n22880 = ~n22878 & ~n22879;
  assign n22881 = ~n22877 & ~n22878;
  assign n22882 = ~n22879 & n22881;
  assign n22883 = ~n22877 & n22880;
  assign n22884 = ~n22876 & n55987;
  assign n22885 = pi11  & ~n22884;
  assign n22886 = ~n22884 & ~n22885;
  assign n22887 = ~pi11  & ~n22884;
  assign n22888 = pi11  & ~n22885;
  assign n22889 = pi11  & n22884;
  assign n22890 = ~n55988 & ~n55989;
  assign n22891 = n22539 & ~n22541;
  assign n22892 = ~n22542 & ~n22891;
  assign n22893 = ~n22890 & n22892;
  assign n22894 = n15195 & n18846;
  assign n22895 = ~n54050 & n55247;
  assign n22896 = ~n54005 & n19541;
  assign n22897 = ~n54034 & n19509;
  assign n22898 = ~n22896 & ~n22897;
  assign n22899 = ~n22895 & ~n22897;
  assign n22900 = ~n22896 & n22899;
  assign n22901 = ~n22895 & n22898;
  assign n22902 = ~n22894 & n55990;
  assign n22903 = pi11  & ~n22902;
  assign n22904 = ~n22902 & ~n22903;
  assign n22905 = ~pi11  & ~n22902;
  assign n22906 = pi11  & ~n22903;
  assign n22907 = pi11  & n22902;
  assign n22908 = ~n55991 & ~n55992;
  assign n22909 = n22530 & n55910;
  assign n22910 = ~n22530 & ~n22538;
  assign n22911 = ~n22530 & n55910;
  assign n22912 = ~n55910 & ~n22538;
  assign n22913 = n22530 & ~n55910;
  assign n22914 = ~n55993 & ~n55994;
  assign n22915 = ~n22538 & ~n22909;
  assign n22916 = ~n22908 & ~n55995;
  assign n22917 = n15219 & n18846;
  assign n22918 = ~n54050 & n19509;
  assign n22919 = ~n54034 & n19541;
  assign n22920 = ~n54073 & n55247;
  assign n22921 = ~n22919 & ~n22920;
  assign n22922 = ~n22918 & ~n22920;
  assign n22923 = ~n22919 & n22922;
  assign n22924 = ~n22918 & n22921;
  assign n22925 = ~n22917 & n55996;
  assign n22926 = pi11  & ~n22925;
  assign n22927 = ~n22925 & ~n22926;
  assign n22928 = ~pi11  & ~n22925;
  assign n22929 = pi11  & ~n22926;
  assign n22930 = pi11  & n22925;
  assign n22931 = ~n55997 & ~n55998;
  assign n22932 = n22521 & n55907;
  assign n22933 = ~n22521 & ~n22529;
  assign n22934 = ~n55907 & ~n22529;
  assign n22935 = ~n22933 & ~n22934;
  assign n22936 = ~n22529 & ~n22932;
  assign n22937 = ~n22931 & ~n55999;
  assign n22938 = n22512 & n55904;
  assign n22939 = ~n22520 & ~n22938;
  assign n22940 = n16138 & n18846;
  assign n22941 = ~n54098 & n55247;
  assign n22942 = ~n54050 & n19541;
  assign n22943 = ~n54073 & n19509;
  assign n22944 = ~n22942 & ~n22943;
  assign n22945 = ~n22941 & ~n22943;
  assign n22946 = ~n22942 & n22945;
  assign n22947 = ~n22941 & n22944;
  assign n22948 = ~n18846 & n56000;
  assign n22949 = ~n16138 & n56000;
  assign n22950 = ~n22948 & ~n22949;
  assign n22951 = ~n22940 & n56000;
  assign n22952 = pi11  & ~n56001;
  assign n22953 = ~pi11  & n56001;
  assign n22954 = ~n22952 & ~n22953;
  assign n22955 = n22939 & ~n22954;
  assign n22956 = n22503 & n55901;
  assign n22957 = ~n22511 & ~n22956;
  assign n22958 = n15779 & n18846;
  assign n22959 = ~n54098 & n19509;
  assign n22960 = ~n54119 & n55247;
  assign n22961 = ~n54073 & n19541;
  assign n22962 = ~n22960 & ~n22961;
  assign n22963 = ~n22959 & ~n22960;
  assign n22964 = ~n22961 & n22963;
  assign n22965 = ~n22959 & ~n22961;
  assign n22966 = ~n22960 & n22965;
  assign n22967 = ~n22959 & n22962;
  assign n22968 = ~n18846 & n56002;
  assign n22969 = ~n15779 & n56002;
  assign n22970 = ~n22968 & ~n22969;
  assign n22971 = ~n22958 & n56002;
  assign n22972 = pi11  & ~n56003;
  assign n22973 = ~pi11  & n56003;
  assign n22974 = ~n22972 & ~n22973;
  assign n22975 = n22957 & ~n22974;
  assign n22976 = n22496 & n55898;
  assign n22977 = ~n22502 & ~n22976;
  assign n22978 = n16547 & n18846;
  assign n22979 = ~n54119 & n19509;
  assign n22980 = ~n54098 & n19541;
  assign n22981 = ~n54132 & n55247;
  assign n22982 = ~n22980 & ~n22981;
  assign n22983 = ~n22979 & ~n22981;
  assign n22984 = ~n22980 & n22983;
  assign n22985 = ~n22979 & n22982;
  assign n22986 = ~n18846 & n56004;
  assign n22987 = ~n16547 & n56004;
  assign n22988 = ~n22986 & ~n22987;
  assign n22989 = ~n22978 & n56004;
  assign n22990 = pi11  & ~n56005;
  assign n22991 = ~pi11  & n56005;
  assign n22992 = ~n22990 & ~n22991;
  assign n22993 = n22977 & ~n22992;
  assign n22994 = n16772 & n18846;
  assign n22995 = ~n54154 & n55247;
  assign n22996 = ~n54119 & n19541;
  assign n22997 = ~n54132 & n19509;
  assign n22998 = ~n22996 & ~n22997;
  assign n22999 = ~n22995 & ~n22997;
  assign n23000 = ~n22996 & n22999;
  assign n23001 = ~n22995 & n22998;
  assign n23002 = ~n22994 & n56006;
  assign n23003 = pi11  & ~n23002;
  assign n23004 = ~n23002 & ~n23003;
  assign n23005 = ~pi11  & ~n23002;
  assign n23006 = pi11  & ~n23003;
  assign n23007 = pi11  & n23002;
  assign n23008 = ~n56007 & ~n56008;
  assign n23009 = n22492 & ~n22494;
  assign n23010 = ~n22495 & ~n23009;
  assign n23011 = ~n23008 & n23010;
  assign n23012 = n16522 & n18846;
  assign n23013 = ~n54154 & n19509;
  assign n23014 = ~n54132 & n19541;
  assign n23015 = ~n54163 & n55247;
  assign n23016 = ~n23014 & ~n23015;
  assign n23017 = ~n23013 & ~n23015;
  assign n23018 = ~n23014 & n23017;
  assign n23019 = ~n23013 & n23016;
  assign n23020 = ~n23012 & n56009;
  assign n23021 = pi11  & ~n23020;
  assign n23022 = ~n23020 & ~n23021;
  assign n23023 = ~pi11  & ~n23020;
  assign n23024 = pi11  & ~n23021;
  assign n23025 = pi11  & n23020;
  assign n23026 = ~n56010 & ~n56011;
  assign n23027 = n22483 & n55897;
  assign n23028 = ~n22483 & ~n22491;
  assign n23029 = ~n55897 & ~n22491;
  assign n23030 = ~n23028 & ~n23029;
  assign n23031 = ~n22491 & ~n23027;
  assign n23032 = ~n23026 & ~n56012;
  assign n23033 = n17072 & n18846;
  assign n23034 = ~n54154 & n19541;
  assign n23035 = ~n54183 & n55247;
  assign n23036 = ~n54163 & n19509;
  assign n23037 = ~n23035 & ~n23036;
  assign n23038 = ~n23034 & n23037;
  assign n23039 = ~n23033 & n23038;
  assign n23040 = pi11  & ~n23039;
  assign n23041 = ~n23039 & ~n23040;
  assign n23042 = ~pi11  & ~n23039;
  assign n23043 = pi11  & ~n23040;
  assign n23044 = pi11  & n23039;
  assign n23045 = ~n56013 & ~n56014;
  assign n23046 = n22474 & n55894;
  assign n23047 = ~n22474 & ~n22482;
  assign n23048 = ~n22474 & n55894;
  assign n23049 = ~n55894 & ~n22482;
  assign n23050 = n22474 & ~n55894;
  assign n23051 = ~n56015 & ~n56016;
  assign n23052 = ~n22482 & ~n23046;
  assign n23053 = ~n23045 & ~n56017;
  assign n23054 = n22465 & n55891;
  assign n23055 = ~n22473 & ~n23054;
  assign n23056 = n17524 & n18846;
  assign n23057 = ~n54183 & n19509;
  assign n23058 = ~n54194 & n55247;
  assign n23059 = ~n54163 & n19541;
  assign n23060 = ~n23058 & ~n23059;
  assign n23061 = ~n23057 & ~n23058;
  assign n23062 = ~n23059 & n23061;
  assign n23063 = ~n23057 & n23060;
  assign n23064 = ~n18846 & n56018;
  assign n23065 = ~n17524 & n56018;
  assign n23066 = ~n23064 & ~n23065;
  assign n23067 = ~n23056 & n56018;
  assign n23068 = pi11  & ~n56019;
  assign n23069 = ~pi11  & n56019;
  assign n23070 = ~n23068 & ~n23069;
  assign n23071 = n23055 & ~n23070;
  assign n23072 = n22461 & ~n22463;
  assign n23073 = ~n22464 & ~n23072;
  assign n23074 = n17544 & n18846;
  assign n23075 = ~n54212 & n55247;
  assign n23076 = ~n54183 & n19541;
  assign n23077 = ~n54194 & n19509;
  assign n23078 = ~n23076 & ~n23077;
  assign n23079 = ~n23075 & ~n23077;
  assign n23080 = ~n23076 & n23079;
  assign n23081 = ~n23075 & n23078;
  assign n23082 = ~n18846 & n56020;
  assign n23083 = ~n17544 & n56020;
  assign n23084 = ~n23082 & ~n23083;
  assign n23085 = ~n23074 & n56020;
  assign n23086 = pi11  & ~n56021;
  assign n23087 = ~pi11  & n56021;
  assign n23088 = ~n23086 & ~n23087;
  assign n23089 = n23073 & ~n23088;
  assign n23090 = n22452 & n55888;
  assign n23091 = ~n22460 & ~n23090;
  assign n23092 = n17041 & n18846;
  assign n23093 = ~n54212 & n19509;
  assign n23094 = ~n54194 & n19541;
  assign n23095 = ~n54240 & n55247;
  assign n23096 = ~n23094 & ~n23095;
  assign n23097 = ~n23093 & ~n23095;
  assign n23098 = ~n23094 & n23097;
  assign n23099 = ~n23093 & n23096;
  assign n23100 = ~n18846 & n56022;
  assign n23101 = ~n17041 & n56022;
  assign n23102 = ~n23100 & ~n23101;
  assign n23103 = ~n23092 & n56022;
  assign n23104 = pi11  & ~n56023;
  assign n23105 = ~pi11  & n56023;
  assign n23106 = ~n23104 & ~n23105;
  assign n23107 = n23091 & ~n23106;
  assign n23108 = n17660 & n18846;
  assign n23109 = ~n54254 & n55247;
  assign n23110 = ~n54212 & n19541;
  assign n23111 = ~n54240 & n19509;
  assign n23112 = ~n23110 & ~n23111;
  assign n23113 = ~n23109 & ~n23111;
  assign n23114 = ~n23110 & n23113;
  assign n23115 = ~n23109 & n23112;
  assign n23116 = ~n23108 & n56024;
  assign n23117 = pi11  & ~n23116;
  assign n23118 = ~n23116 & ~n23117;
  assign n23119 = ~pi11  & ~n23116;
  assign n23120 = pi11  & ~n23117;
  assign n23121 = pi11  & n23116;
  assign n23122 = ~n56025 & ~n56026;
  assign n23123 = n22448 & ~n22450;
  assign n23124 = ~n22451 & ~n23123;
  assign n23125 = ~n23122 & n23124;
  assign n23126 = n17804 & n18846;
  assign n23127 = ~n54254 & n19509;
  assign n23128 = ~n54240 & n19541;
  assign n23129 = ~n54269 & n55247;
  assign n23130 = ~n23128 & ~n23129;
  assign n23131 = ~n23127 & ~n23129;
  assign n23132 = ~n23128 & n23131;
  assign n23133 = ~n23127 & n23130;
  assign n23134 = ~n18846 & n56027;
  assign n23135 = ~n17804 & n56027;
  assign n23136 = ~n23134 & ~n23135;
  assign n23137 = ~n23126 & n56027;
  assign n23138 = pi11  & ~n56028;
  assign n23139 = ~pi11  & n56028;
  assign n23140 = ~n23138 & ~n23139;
  assign n23141 = n22439 & n55885;
  assign n23142 = ~n55885 & ~n22447;
  assign n23143 = ~n22439 & ~n22447;
  assign n23144 = ~n23142 & ~n23143;
  assign n23145 = ~n22447 & ~n23141;
  assign n23146 = ~n23140 & ~n56029;
  assign n23147 = n17939 & n18846;
  assign n23148 = ~n54254 & n19541;
  assign n23149 = ~n54277 & n55247;
  assign n23150 = ~n54269 & n19509;
  assign n23151 = ~n23149 & ~n23150;
  assign n23152 = ~n23148 & n23151;
  assign n23153 = ~n23147 & n23152;
  assign n23154 = pi11  & ~n23153;
  assign n23155 = ~n23153 & ~n23154;
  assign n23156 = ~pi11  & ~n23153;
  assign n23157 = pi11  & ~n23154;
  assign n23158 = pi11  & n23153;
  assign n23159 = ~n56030 & ~n56031;
  assign n23160 = pi14  & ~n55877;
  assign n23161 = ~n55878 & ~n23160;
  assign n23162 = n55878 & n23160;
  assign n23163 = ~n55877 & n22421;
  assign n23164 = ~n55879 & ~n23163;
  assign n23165 = ~n23161 & ~n23162;
  assign n23166 = ~n23159 & n56032;
  assign n23167 = n18056 & n18846;
  assign n23168 = ~n54305 & n55247;
  assign n23169 = ~n54277 & n19509;
  assign n23170 = ~n54269 & n19541;
  assign n23171 = ~n23169 & ~n23170;
  assign n23172 = ~n23168 & ~n23169;
  assign n23173 = ~n23170 & n23172;
  assign n23174 = ~n23168 & n23171;
  assign n23175 = ~n18846 & n56033;
  assign n23176 = ~n18056 & n56033;
  assign n23177 = ~n23175 & ~n23176;
  assign n23178 = ~n23167 & n56033;
  assign n23179 = pi11  & ~n56034;
  assign n23180 = ~pi11  & n56034;
  assign n23181 = ~n23179 & ~n23180;
  assign n23182 = pi14  & n22401;
  assign n23183 = ~n22400 & n23182;
  assign n23184 = n22400 & ~n23182;
  assign n23185 = ~n22402 & n22406;
  assign n23186 = ~n55877 & ~n23185;
  assign n23187 = ~n23183 & ~n23184;
  assign n23188 = ~n23181 & n56035;
  assign n23189 = n18846 & ~n19275;
  assign n23190 = ~n54325 & n19509;
  assign n23191 = ~n54344 & n19541;
  assign n23192 = ~n23190 & ~n23191;
  assign n23193 = ~n23189 & n23192;
  assign n23194 = ~n54325 & n55244;
  assign n23195 = pi11  & ~n23194;
  assign n23196 = pi11  & ~n23193;
  assign n23197 = pi11  & ~n23196;
  assign n23198 = ~n23193 & ~n23196;
  assign n23199 = ~n23197 & ~n23198;
  assign n23200 = n23195 & ~n23199;
  assign n23201 = n23193 & n23195;
  assign n23202 = n18156 & n18846;
  assign n23203 = ~n54305 & n19541;
  assign n23204 = ~n54325 & n55247;
  assign n23205 = ~n54344 & n19509;
  assign n23206 = ~n23204 & ~n23205;
  assign n23207 = ~n23203 & n23206;
  assign n23208 = ~n18846 & n23207;
  assign n23209 = ~n18156 & n23207;
  assign n23210 = ~n23208 & ~n23209;
  assign n23211 = ~n23202 & n23207;
  assign n23212 = pi11  & ~n56037;
  assign n23213 = ~pi11  & n56037;
  assign n23214 = ~n23212 & ~n23213;
  assign n23215 = n56036 & ~n23214;
  assign n23216 = n56036 & ~n56037;
  assign n23217 = n22401 & n56038;
  assign n23218 = n18336 & n18846;
  assign n23219 = ~n54305 & n19509;
  assign n23220 = ~n54277 & n19541;
  assign n23221 = ~n54344 & n55247;
  assign n23222 = ~n23220 & ~n23221;
  assign n23223 = ~n23219 & ~n23221;
  assign n23224 = ~n23220 & n23223;
  assign n23225 = ~n23219 & n23222;
  assign n23226 = ~n23218 & n56039;
  assign n23227 = pi11  & ~n23226;
  assign n23228 = pi11  & ~n23227;
  assign n23229 = pi11  & n23226;
  assign n23230 = ~n23226 & ~n23227;
  assign n23231 = ~pi11  & ~n23226;
  assign n23232 = ~n56040 & ~n56041;
  assign n23233 = ~n22401 & ~n56038;
  assign n23234 = n56038 & ~n23217;
  assign n23235 = ~n22401 & n56038;
  assign n23236 = n22401 & ~n23217;
  assign n23237 = n22401 & ~n56038;
  assign n23238 = ~n56042 & ~n56043;
  assign n23239 = ~n23217 & ~n23233;
  assign n23240 = ~n23232 & ~n56044;
  assign n23241 = ~n23217 & ~n23240;
  assign n23242 = n23181 & ~n56035;
  assign n23243 = ~n23188 & ~n23242;
  assign n23244 = ~n23241 & n23243;
  assign n23245 = ~n23188 & ~n23244;
  assign n23246 = n23159 & ~n56032;
  assign n23247 = ~n23159 & ~n23166;
  assign n23248 = ~n23159 & ~n56032;
  assign n23249 = n56032 & ~n23166;
  assign n23250 = n23159 & n56032;
  assign n23251 = ~n56045 & ~n56046;
  assign n23252 = ~n23166 & ~n23246;
  assign n23253 = ~n23245 & ~n56047;
  assign n23254 = ~n23166 & ~n23253;
  assign n23255 = n23140 & n56029;
  assign n23256 = ~n23146 & ~n23255;
  assign n23257 = ~n23254 & n23256;
  assign n23258 = ~n23146 & ~n23257;
  assign n23259 = n23122 & ~n23124;
  assign n23260 = ~n23122 & ~n23125;
  assign n23261 = ~n23122 & ~n23124;
  assign n23262 = n23124 & ~n23125;
  assign n23263 = n23122 & n23124;
  assign n23264 = ~n56048 & ~n56049;
  assign n23265 = ~n23125 & ~n23259;
  assign n23266 = ~n23258 & ~n56050;
  assign n23267 = ~n23125 & ~n23266;
  assign n23268 = ~n23091 & n23106;
  assign n23269 = n23091 & ~n23107;
  assign n23270 = n23091 & n23106;
  assign n23271 = ~n23106 & ~n23107;
  assign n23272 = ~n23091 & ~n23106;
  assign n23273 = ~n56051 & ~n56052;
  assign n23274 = ~n23107 & ~n23268;
  assign n23275 = ~n23267 & ~n56053;
  assign n23276 = ~n23107 & ~n23275;
  assign n23277 = ~n23073 & n23088;
  assign n23278 = n23073 & ~n23089;
  assign n23279 = n23073 & n23088;
  assign n23280 = ~n23088 & ~n23089;
  assign n23281 = ~n23073 & ~n23088;
  assign n23282 = ~n56054 & ~n56055;
  assign n23283 = ~n23089 & ~n23277;
  assign n23284 = ~n23276 & ~n56056;
  assign n23285 = ~n23089 & ~n23284;
  assign n23286 = ~n23055 & n23070;
  assign n23287 = ~n23071 & ~n23286;
  assign n23288 = ~n23285 & n23287;
  assign n23289 = ~n23071 & ~n23288;
  assign n23290 = n23045 & n56017;
  assign n23291 = ~n23045 & ~n23053;
  assign n23292 = ~n56017 & ~n23053;
  assign n23293 = ~n23291 & ~n23292;
  assign n23294 = ~n23053 & ~n23290;
  assign n23295 = ~n23289 & ~n56057;
  assign n23296 = ~n23053 & ~n23295;
  assign n23297 = n23026 & n56012;
  assign n23298 = ~n23026 & ~n23032;
  assign n23299 = ~n23026 & n56012;
  assign n23300 = ~n56012 & ~n23032;
  assign n23301 = n23026 & ~n56012;
  assign n23302 = ~n56058 & ~n56059;
  assign n23303 = ~n23032 & ~n23297;
  assign n23304 = ~n23296 & ~n56060;
  assign n23305 = ~n23032 & ~n23304;
  assign n23306 = n23008 & ~n23010;
  assign n23307 = ~n23008 & ~n23011;
  assign n23308 = ~n23008 & ~n23010;
  assign n23309 = n23010 & ~n23011;
  assign n23310 = n23008 & n23010;
  assign n23311 = ~n56061 & ~n56062;
  assign n23312 = ~n23011 & ~n23306;
  assign n23313 = ~n23305 & ~n56063;
  assign n23314 = ~n23011 & ~n23313;
  assign n23315 = ~n22977 & n22992;
  assign n23316 = n22977 & ~n22993;
  assign n23317 = n22977 & n22992;
  assign n23318 = ~n22992 & ~n22993;
  assign n23319 = ~n22977 & ~n22992;
  assign n23320 = ~n56064 & ~n56065;
  assign n23321 = ~n22993 & ~n23315;
  assign n23322 = ~n23314 & ~n56066;
  assign n23323 = ~n22993 & ~n23322;
  assign n23324 = ~n22957 & n22974;
  assign n23325 = n22957 & ~n22975;
  assign n23326 = n22957 & n22974;
  assign n23327 = ~n22974 & ~n22975;
  assign n23328 = ~n22957 & ~n22974;
  assign n23329 = ~n56067 & ~n56068;
  assign n23330 = ~n22975 & ~n23324;
  assign n23331 = ~n23323 & ~n56069;
  assign n23332 = ~n22975 & ~n23331;
  assign n23333 = ~n22939 & n22954;
  assign n23334 = ~n22955 & ~n23333;
  assign n23335 = ~n23332 & n23334;
  assign n23336 = ~n22955 & ~n23335;
  assign n23337 = n22931 & n55999;
  assign n23338 = ~n22931 & ~n22937;
  assign n23339 = ~n22931 & n55999;
  assign n23340 = ~n55999 & ~n22937;
  assign n23341 = n22931 & ~n55999;
  assign n23342 = ~n56070 & ~n56071;
  assign n23343 = ~n22937 & ~n23337;
  assign n23344 = ~n23336 & ~n56072;
  assign n23345 = ~n22937 & ~n23344;
  assign n23346 = n22908 & n55995;
  assign n23347 = ~n22908 & ~n22916;
  assign n23348 = ~n55995 & ~n22916;
  assign n23349 = ~n23347 & ~n23348;
  assign n23350 = ~n22916 & ~n23346;
  assign n23351 = ~n23345 & ~n56073;
  assign n23352 = ~n22916 & ~n23351;
  assign n23353 = n22890 & ~n22892;
  assign n23354 = ~n22890 & ~n22893;
  assign n23355 = ~n22890 & ~n22892;
  assign n23356 = n22892 & ~n22893;
  assign n23357 = n22890 & n22892;
  assign n23358 = ~n56074 & ~n56075;
  assign n23359 = ~n22893 & ~n23353;
  assign n23360 = ~n23352 & ~n56076;
  assign n23361 = ~n22893 & ~n23360;
  assign n23362 = ~n22859 & n22874;
  assign n23363 = n22859 & ~n22875;
  assign n23364 = n22859 & n22874;
  assign n23365 = ~n22874 & ~n22875;
  assign n23366 = ~n22859 & ~n22874;
  assign n23367 = ~n56077 & ~n56078;
  assign n23368 = ~n22875 & ~n23362;
  assign n23369 = ~n23361 & ~n56079;
  assign n23370 = ~n22875 & ~n23369;
  assign n23371 = ~n22841 & n22856;
  assign n23372 = ~n22857 & ~n23371;
  assign n23373 = ~n23370 & n23372;
  assign n23374 = ~n22857 & ~n23373;
  assign n23375 = n22831 & n55982;
  assign n23376 = ~n22831 & ~n22839;
  assign n23377 = ~n55982 & ~n22839;
  assign n23378 = ~n23376 & ~n23377;
  assign n23379 = ~n22839 & ~n23375;
  assign n23380 = ~n23374 & ~n56080;
  assign n23381 = ~n22839 & ~n23380;
  assign n23382 = n22810 & n55976;
  assign n23383 = ~n22810 & ~n22816;
  assign n23384 = ~n22810 & n55976;
  assign n23385 = ~n55976 & ~n22816;
  assign n23386 = n22810 & ~n55976;
  assign n23387 = ~n56081 & ~n56082;
  assign n23388 = ~n22816 & ~n23382;
  assign n23389 = ~n23381 & ~n56083;
  assign n23390 = ~n22816 & ~n23389;
  assign n23391 = n22789 & n55972;
  assign n23392 = ~n22789 & ~n22795;
  assign n23393 = ~n22789 & n55972;
  assign n23394 = ~n55972 & ~n22795;
  assign n23395 = n22789 & ~n55972;
  assign n23396 = ~n56084 & ~n56085;
  assign n23397 = ~n22795 & ~n23391;
  assign n23398 = ~n23390 & ~n56086;
  assign n23399 = ~n22795 & ~n23398;
  assign n23400 = n22766 & n55968;
  assign n23401 = ~n22766 & ~n22774;
  assign n23402 = ~n55968 & ~n22774;
  assign n23403 = ~n23401 & ~n23402;
  assign n23404 = ~n22774 & ~n23400;
  assign n23405 = ~n23399 & ~n56087;
  assign n23406 = ~n22774 & ~n23405;
  assign n23407 = n22743 & n55962;
  assign n23408 = ~n22743 & ~n22751;
  assign n23409 = ~n55962 & ~n22751;
  assign n23410 = ~n23408 & ~n23409;
  assign n23411 = ~n22751 & ~n23407;
  assign n23412 = ~n23406 & ~n56088;
  assign n23413 = ~n22751 & ~n23412;
  assign n23414 = n22722 & n55956;
  assign n23415 = ~n22722 & ~n22728;
  assign n23416 = ~n22722 & n55956;
  assign n23417 = ~n55956 & ~n22728;
  assign n23418 = n22722 & ~n55956;
  assign n23419 = ~n56089 & ~n56090;
  assign n23420 = ~n22728 & ~n23414;
  assign n23421 = ~n23413 & ~n56091;
  assign n23422 = ~n22728 & ~n23421;
  assign n23423 = n22701 & n55952;
  assign n23424 = ~n22701 & ~n22707;
  assign n23425 = ~n22701 & n55952;
  assign n23426 = ~n55952 & ~n22707;
  assign n23427 = n22701 & ~n55952;
  assign n23428 = ~n56092 & ~n56093;
  assign n23429 = ~n22707 & ~n23423;
  assign n23430 = ~n23422 & ~n56094;
  assign n23431 = ~n22707 & ~n23430;
  assign n23432 = n22642 & ~n22644;
  assign n23433 = ~n22645 & ~n23432;
  assign n23434 = ~n23431 & n23433;
  assign n23435 = n11380 & n20085;
  assign n23436 = ~n53685 & n21237;
  assign n23437 = ~n53657 & n21269;
  assign n23438 = ~n53712 & n55472;
  assign n23439 = ~n23437 & ~n23438;
  assign n23440 = ~n23436 & ~n23438;
  assign n23441 = ~n23437 & n23440;
  assign n23442 = ~n23436 & n23439;
  assign n23443 = ~n23435 & n56095;
  assign n23444 = pi8  & ~n23443;
  assign n23445 = ~n23443 & ~n23444;
  assign n23446 = ~pi8  & ~n23443;
  assign n23447 = pi8  & ~n23444;
  assign n23448 = pi8  & n23443;
  assign n23449 = ~n56096 & ~n56097;
  assign n23450 = n23431 & ~n23433;
  assign n23451 = ~n23431 & ~n23434;
  assign n23452 = n23433 & ~n23434;
  assign n23453 = ~n23451 & ~n23452;
  assign n23454 = ~n23434 & ~n23450;
  assign n23455 = ~n23449 & ~n56098;
  assign n23456 = ~n23434 & ~n23455;
  assign n23457 = n77 & n54351;
  assign n23458 = ~n53634 & n21969;
  assign n23459 = ~n53439 & n55818;
  assign n23460 = ~n2325 & n23459;
  assign n23461 = ~n23458 & ~n23460;
  assign n23462 = ~n77 & n23461;
  assign n23463 = ~n54351 & n23461;
  assign n23464 = ~n23462 & ~n23463;
  assign n23465 = ~n23457 & n23461;
  assign n23466 = pi5  & ~n56099;
  assign n23467 = ~pi5  & n56099;
  assign n23468 = ~n23466 & ~n23467;
  assign n23469 = ~n23456 & ~n23468;
  assign n23470 = n23456 & n23468;
  assign n23471 = ~n23469 & ~n23470;
  assign n23472 = n22668 & ~n22670;
  assign n23473 = n22670 & ~n22671;
  assign n23474 = ~n22668 & ~n22671;
  assign n23475 = ~n23473 & ~n23474;
  assign n23476 = ~n22671 & ~n23472;
  assign n23477 = n23471 & ~n56100;
  assign n23478 = ~n23469 & ~n23477;
  assign n23479 = n55947 & ~n22682;
  assign n23480 = ~n55947 & ~n22683;
  assign n23481 = n22682 & ~n22683;
  assign n23482 = ~n23480 & ~n23481;
  assign n23483 = ~n22683 & ~n23479;
  assign n23484 = ~n23478 & ~n56101;
  assign n23485 = n23478 & n56101;
  assign n23486 = ~n23484 & ~n23485;
  assign n23487 = n23422 & n56094;
  assign n23488 = ~n23430 & ~n23487;
  assign n23489 = n11360 & n20085;
  assign n23490 = ~n53685 & n21269;
  assign n23491 = ~n53741 & n55472;
  assign n23492 = ~n53712 & n21237;
  assign n23493 = ~n23491 & ~n23492;
  assign n23494 = ~n23490 & ~n23491;
  assign n23495 = ~n23492 & n23494;
  assign n23496 = ~n23490 & n23493;
  assign n23497 = ~n20085 & n56102;
  assign n23498 = ~n11360 & n56102;
  assign n23499 = ~n23497 & ~n23498;
  assign n23500 = ~n23489 & n56102;
  assign n23501 = pi8  & ~n56103;
  assign n23502 = ~pi8  & n56103;
  assign n23503 = ~n23501 & ~n23502;
  assign n23504 = n23488 & ~n23503;
  assign n23505 = n23413 & n56091;
  assign n23506 = ~n23421 & ~n23505;
  assign n23507 = n11889 & n20085;
  assign n23508 = ~n53712 & n21269;
  assign n23509 = ~n53774 & n55472;
  assign n23510 = ~n53741 & n21237;
  assign n23511 = ~n23509 & ~n23510;
  assign n23512 = ~n23508 & ~n23509;
  assign n23513 = ~n23510 & n23512;
  assign n23514 = ~n23508 & n23511;
  assign n23515 = ~n20085 & n56104;
  assign n23516 = ~n11889 & n56104;
  assign n23517 = ~n23515 & ~n23516;
  assign n23518 = ~n23507 & n56104;
  assign n23519 = pi8  & ~n56105;
  assign n23520 = ~pi8  & n56105;
  assign n23521 = ~n23519 & ~n23520;
  assign n23522 = n23506 & ~n23521;
  assign n23523 = n23406 & n56088;
  assign n23524 = ~n23412 & ~n23523;
  assign n23525 = n11913 & n20085;
  assign n23526 = ~n53774 & n21237;
  assign n23527 = ~n53799 & n55472;
  assign n23528 = ~n53741 & n21269;
  assign n23529 = ~n23527 & ~n23528;
  assign n23530 = ~n23526 & ~n23527;
  assign n23531 = ~n23528 & n23530;
  assign n23532 = ~n23526 & n23529;
  assign n23533 = ~n20085 & n56106;
  assign n23534 = ~n11913 & n56106;
  assign n23535 = ~n23533 & ~n23534;
  assign n23536 = ~n23525 & n56106;
  assign n23537 = pi8  & ~n56107;
  assign n23538 = ~pi8  & n56107;
  assign n23539 = ~n23537 & ~n23538;
  assign n23540 = n23524 & ~n23539;
  assign n23541 = n23399 & n56087;
  assign n23542 = ~n23405 & ~n23541;
  assign n23543 = n12690 & n20085;
  assign n23544 = ~n53774 & n21269;
  assign n23545 = ~n53819 & n55472;
  assign n23546 = ~n53799 & n21237;
  assign n23547 = ~n23545 & ~n23546;
  assign n23548 = ~n23544 & ~n23545;
  assign n23549 = ~n23546 & n23548;
  assign n23550 = ~n23544 & n23547;
  assign n23551 = ~n20085 & n56108;
  assign n23552 = ~n12690 & n56108;
  assign n23553 = ~n23551 & ~n23552;
  assign n23554 = ~n23543 & n56108;
  assign n23555 = pi8  & ~n56109;
  assign n23556 = ~pi8  & n56109;
  assign n23557 = ~n23555 & ~n23556;
  assign n23558 = n23542 & ~n23557;
  assign n23559 = n23390 & n56086;
  assign n23560 = ~n23398 & ~n23559;
  assign n23561 = n12550 & n20085;
  assign n23562 = ~n53819 & n21237;
  assign n23563 = ~n53845 & n55472;
  assign n23564 = ~n53799 & n21269;
  assign n23565 = ~n23563 & ~n23564;
  assign n23566 = ~n23562 & ~n23563;
  assign n23567 = ~n23564 & n23566;
  assign n23568 = ~n23562 & n23565;
  assign n23569 = ~n20085 & n56110;
  assign n23570 = ~n12550 & n56110;
  assign n23571 = ~n23569 & ~n23570;
  assign n23572 = ~n23561 & n56110;
  assign n23573 = pi8  & ~n56111;
  assign n23574 = ~pi8  & n56111;
  assign n23575 = ~n23573 & ~n23574;
  assign n23576 = n23560 & ~n23575;
  assign n23577 = n23381 & n56083;
  assign n23578 = ~n23389 & ~n23577;
  assign n23579 = n12938 & n20085;
  assign n23580 = ~n53819 & n21269;
  assign n23581 = ~n53860 & n55472;
  assign n23582 = ~n53845 & n21237;
  assign n23583 = ~n23581 & ~n23582;
  assign n23584 = ~n23580 & ~n23581;
  assign n23585 = ~n23582 & n23584;
  assign n23586 = ~n23580 & n23583;
  assign n23587 = ~n20085 & n56112;
  assign n23588 = ~n12938 & n56112;
  assign n23589 = ~n23587 & ~n23588;
  assign n23590 = ~n23579 & n56112;
  assign n23591 = pi8  & ~n56113;
  assign n23592 = ~pi8  & n56113;
  assign n23593 = ~n23591 & ~n23592;
  assign n23594 = n23578 & ~n23593;
  assign n23595 = n23374 & n56080;
  assign n23596 = ~n23380 & ~n23595;
  assign n23597 = n12918 & n20085;
  assign n23598 = ~n53860 & n21237;
  assign n23599 = ~n53888 & n55472;
  assign n23600 = ~n53845 & n21269;
  assign n23601 = ~n23599 & ~n23600;
  assign n23602 = ~n23598 & ~n23599;
  assign n23603 = ~n23600 & n23602;
  assign n23604 = ~n23598 & n23601;
  assign n23605 = ~n20085 & n56114;
  assign n23606 = ~n12918 & n56114;
  assign n23607 = ~n23605 & ~n23606;
  assign n23608 = ~n23597 & n56114;
  assign n23609 = pi8  & ~n56115;
  assign n23610 = ~pi8  & n56115;
  assign n23611 = ~n23609 & ~n23610;
  assign n23612 = n23596 & ~n23611;
  assign n23613 = n13336 & n20085;
  assign n23614 = ~n53888 & n21237;
  assign n23615 = ~n53907 & n55472;
  assign n23616 = ~n53860 & n21269;
  assign n23617 = ~n23615 & ~n23616;
  assign n23618 = ~n23614 & ~n23615;
  assign n23619 = ~n23616 & n23618;
  assign n23620 = ~n23614 & n23617;
  assign n23621 = ~n23613 & n56116;
  assign n23622 = pi8  & ~n23621;
  assign n23623 = ~n23621 & ~n23622;
  assign n23624 = ~pi8  & ~n23621;
  assign n23625 = pi8  & ~n23622;
  assign n23626 = pi8  & n23621;
  assign n23627 = ~n56117 & ~n56118;
  assign n23628 = n23370 & ~n23372;
  assign n23629 = ~n23373 & ~n23628;
  assign n23630 = ~n23627 & n23629;
  assign n23631 = n13360 & n20085;
  assign n23632 = ~n53907 & n21237;
  assign n23633 = ~n53930 & n55472;
  assign n23634 = ~n53888 & n21269;
  assign n23635 = ~n23633 & ~n23634;
  assign n23636 = ~n23632 & ~n23633;
  assign n23637 = ~n23634 & n23636;
  assign n23638 = ~n23632 & n23635;
  assign n23639 = ~n23631 & n56119;
  assign n23640 = pi8  & ~n23639;
  assign n23641 = ~n23639 & ~n23640;
  assign n23642 = ~pi8  & ~n23639;
  assign n23643 = pi8  & ~n23640;
  assign n23644 = pi8  & n23639;
  assign n23645 = ~n56120 & ~n56121;
  assign n23646 = n23361 & n56079;
  assign n23647 = ~n23361 & ~n23369;
  assign n23648 = ~n23361 & n56079;
  assign n23649 = ~n56079 & ~n23369;
  assign n23650 = n23361 & ~n56079;
  assign n23651 = ~n56122 & ~n56123;
  assign n23652 = ~n23369 & ~n23646;
  assign n23653 = ~n23645 & ~n56124;
  assign n23654 = n23352 & n56076;
  assign n23655 = ~n23360 & ~n23654;
  assign n23656 = n14263 & n20085;
  assign n23657 = ~n53930 & n21237;
  assign n23658 = ~n53962 & n55472;
  assign n23659 = ~n53907 & n21269;
  assign n23660 = ~n23658 & ~n23659;
  assign n23661 = ~n23657 & ~n23658;
  assign n23662 = ~n23659 & n23661;
  assign n23663 = ~n23657 & n23660;
  assign n23664 = ~n20085 & n56125;
  assign n23665 = ~n14263 & n56125;
  assign n23666 = ~n23664 & ~n23665;
  assign n23667 = ~n23656 & n56125;
  assign n23668 = pi8  & ~n56126;
  assign n23669 = ~pi8  & n56126;
  assign n23670 = ~n23668 & ~n23669;
  assign n23671 = n23655 & ~n23670;
  assign n23672 = n23345 & n56073;
  assign n23673 = ~n23351 & ~n23672;
  assign n23674 = n14020 & n20085;
  assign n23675 = ~n53962 & n21237;
  assign n23676 = ~n53970 & n55472;
  assign n23677 = ~n53930 & n21269;
  assign n23678 = ~n23676 & ~n23677;
  assign n23679 = ~n23675 & ~n23676;
  assign n23680 = ~n23677 & n23679;
  assign n23681 = ~n23675 & n23678;
  assign n23682 = ~n20085 & n56127;
  assign n23683 = ~n14020 & n56127;
  assign n23684 = ~n23682 & ~n23683;
  assign n23685 = ~n23674 & n56127;
  assign n23686 = pi8  & ~n56128;
  assign n23687 = ~pi8  & n56128;
  assign n23688 = ~n23686 & ~n23687;
  assign n23689 = n23673 & ~n23688;
  assign n23690 = n23336 & n56072;
  assign n23691 = ~n23344 & ~n23690;
  assign n23692 = n14708 & n20085;
  assign n23693 = ~n54005 & n55472;
  assign n23694 = ~n53970 & n21237;
  assign n23695 = ~n53962 & n21269;
  assign n23696 = ~n23694 & ~n23695;
  assign n23697 = ~n23693 & ~n23694;
  assign n23698 = ~n23695 & n23697;
  assign n23699 = ~n23693 & n23696;
  assign n23700 = ~n20085 & n56129;
  assign n23701 = ~n14708 & n56129;
  assign n23702 = ~n23700 & ~n23701;
  assign n23703 = ~n23692 & n56129;
  assign n23704 = pi8  & ~n56130;
  assign n23705 = ~pi8  & n56130;
  assign n23706 = ~n23704 & ~n23705;
  assign n23707 = n23691 & ~n23706;
  assign n23708 = n14688 & n20085;
  assign n23709 = ~n54005 & n21237;
  assign n23710 = ~n54034 & n55472;
  assign n23711 = ~n53970 & n21269;
  assign n23712 = ~n23710 & ~n23711;
  assign n23713 = ~n23709 & ~n23710;
  assign n23714 = ~n23711 & n23713;
  assign n23715 = ~n23709 & n23712;
  assign n23716 = ~n23708 & n56131;
  assign n23717 = pi8  & ~n23716;
  assign n23718 = ~n23716 & ~n23717;
  assign n23719 = ~pi8  & ~n23716;
  assign n23720 = pi8  & ~n23717;
  assign n23721 = pi8  & n23716;
  assign n23722 = ~n56132 & ~n56133;
  assign n23723 = n23332 & ~n23334;
  assign n23724 = ~n23335 & ~n23723;
  assign n23725 = ~n23722 & n23724;
  assign n23726 = n15195 & n20085;
  assign n23727 = ~n54050 & n55472;
  assign n23728 = ~n54005 & n21269;
  assign n23729 = ~n54034 & n21237;
  assign n23730 = ~n23728 & ~n23729;
  assign n23731 = ~n23727 & ~n23729;
  assign n23732 = ~n23728 & n23731;
  assign n23733 = ~n23727 & n23730;
  assign n23734 = ~n23726 & n56134;
  assign n23735 = pi8  & ~n23734;
  assign n23736 = ~n23734 & ~n23735;
  assign n23737 = ~pi8  & ~n23734;
  assign n23738 = pi8  & ~n23735;
  assign n23739 = pi8  & n23734;
  assign n23740 = ~n56135 & ~n56136;
  assign n23741 = n23323 & n56069;
  assign n23742 = ~n23323 & ~n23331;
  assign n23743 = ~n23323 & n56069;
  assign n23744 = ~n56069 & ~n23331;
  assign n23745 = n23323 & ~n56069;
  assign n23746 = ~n56137 & ~n56138;
  assign n23747 = ~n23331 & ~n23741;
  assign n23748 = ~n23740 & ~n56139;
  assign n23749 = n15219 & n20085;
  assign n23750 = ~n54050 & n21237;
  assign n23751 = ~n54034 & n21269;
  assign n23752 = ~n54073 & n55472;
  assign n23753 = ~n23751 & ~n23752;
  assign n23754 = ~n23750 & ~n23752;
  assign n23755 = ~n23751 & n23754;
  assign n23756 = ~n23750 & n23753;
  assign n23757 = ~n23749 & n56140;
  assign n23758 = pi8  & ~n23757;
  assign n23759 = ~n23757 & ~n23758;
  assign n23760 = ~pi8  & ~n23757;
  assign n23761 = pi8  & ~n23758;
  assign n23762 = pi8  & n23757;
  assign n23763 = ~n56141 & ~n56142;
  assign n23764 = n23314 & n56066;
  assign n23765 = ~n23314 & ~n23322;
  assign n23766 = ~n56066 & ~n23322;
  assign n23767 = ~n23765 & ~n23766;
  assign n23768 = ~n23322 & ~n23764;
  assign n23769 = ~n23763 & ~n56143;
  assign n23770 = n23305 & n56063;
  assign n23771 = ~n23313 & ~n23770;
  assign n23772 = n16138 & n20085;
  assign n23773 = ~n54098 & n55472;
  assign n23774 = ~n54050 & n21269;
  assign n23775 = ~n54073 & n21237;
  assign n23776 = ~n23774 & ~n23775;
  assign n23777 = ~n23773 & ~n23775;
  assign n23778 = ~n23774 & n23777;
  assign n23779 = ~n23773 & n23776;
  assign n23780 = ~n20085 & n56144;
  assign n23781 = ~n16138 & n56144;
  assign n23782 = ~n23780 & ~n23781;
  assign n23783 = ~n23772 & n56144;
  assign n23784 = pi8  & ~n56145;
  assign n23785 = ~pi8  & n56145;
  assign n23786 = ~n23784 & ~n23785;
  assign n23787 = n23771 & ~n23786;
  assign n23788 = n23296 & n56060;
  assign n23789 = ~n23304 & ~n23788;
  assign n23790 = n15779 & n20085;
  assign n23791 = ~n54098 & n21237;
  assign n23792 = ~n54119 & n55472;
  assign n23793 = ~n54073 & n21269;
  assign n23794 = ~n23792 & ~n23793;
  assign n23795 = ~n23791 & ~n23792;
  assign n23796 = ~n23793 & n23795;
  assign n23797 = ~n23791 & ~n23793;
  assign n23798 = ~n23792 & n23797;
  assign n23799 = ~n23791 & n23794;
  assign n23800 = ~n20085 & n56146;
  assign n23801 = ~n15779 & n56146;
  assign n23802 = ~n23800 & ~n23801;
  assign n23803 = ~n23790 & n56146;
  assign n23804 = pi8  & ~n56147;
  assign n23805 = ~pi8  & n56147;
  assign n23806 = ~n23804 & ~n23805;
  assign n23807 = n23789 & ~n23806;
  assign n23808 = n23289 & n56057;
  assign n23809 = ~n23295 & ~n23808;
  assign n23810 = n16547 & n20085;
  assign n23811 = ~n54119 & n21237;
  assign n23812 = ~n54098 & n21269;
  assign n23813 = ~n54132 & n55472;
  assign n23814 = ~n23812 & ~n23813;
  assign n23815 = ~n23811 & ~n23813;
  assign n23816 = ~n23812 & n23815;
  assign n23817 = ~n23811 & n23814;
  assign n23818 = ~n20085 & n56148;
  assign n23819 = ~n16547 & n56148;
  assign n23820 = ~n23818 & ~n23819;
  assign n23821 = ~n23810 & n56148;
  assign n23822 = pi8  & ~n56149;
  assign n23823 = ~pi8  & n56149;
  assign n23824 = ~n23822 & ~n23823;
  assign n23825 = n23809 & ~n23824;
  assign n23826 = n16772 & n20085;
  assign n23827 = ~n54154 & n55472;
  assign n23828 = ~n54119 & n21269;
  assign n23829 = ~n54132 & n21237;
  assign n23830 = ~n23828 & ~n23829;
  assign n23831 = ~n23827 & ~n23829;
  assign n23832 = ~n23828 & n23831;
  assign n23833 = ~n23827 & n23830;
  assign n23834 = ~n23826 & n56150;
  assign n23835 = pi8  & ~n23834;
  assign n23836 = ~n23834 & ~n23835;
  assign n23837 = ~pi8  & ~n23834;
  assign n23838 = pi8  & ~n23835;
  assign n23839 = pi8  & n23834;
  assign n23840 = ~n56151 & ~n56152;
  assign n23841 = n23285 & ~n23287;
  assign n23842 = ~n23288 & ~n23841;
  assign n23843 = ~n23840 & n23842;
  assign n23844 = n16522 & n20085;
  assign n23845 = ~n54154 & n21237;
  assign n23846 = ~n54132 & n21269;
  assign n23847 = ~n54163 & n55472;
  assign n23848 = ~n23846 & ~n23847;
  assign n23849 = ~n23845 & ~n23847;
  assign n23850 = ~n23846 & n23849;
  assign n23851 = ~n23845 & n23848;
  assign n23852 = ~n23844 & n56153;
  assign n23853 = pi8  & ~n23852;
  assign n23854 = ~n23852 & ~n23853;
  assign n23855 = ~pi8  & ~n23852;
  assign n23856 = pi8  & ~n23853;
  assign n23857 = pi8  & n23852;
  assign n23858 = ~n56154 & ~n56155;
  assign n23859 = n23276 & n56056;
  assign n23860 = ~n23276 & ~n23284;
  assign n23861 = ~n56056 & ~n23284;
  assign n23862 = ~n23860 & ~n23861;
  assign n23863 = ~n23284 & ~n23859;
  assign n23864 = ~n23858 & ~n56156;
  assign n23865 = n17072 & n20085;
  assign n23866 = ~n54154 & n21269;
  assign n23867 = ~n54183 & n55472;
  assign n23868 = ~n54163 & n21237;
  assign n23869 = ~n23867 & ~n23868;
  assign n23870 = ~n23866 & n23869;
  assign n23871 = ~n23865 & n23870;
  assign n23872 = pi8  & ~n23871;
  assign n23873 = ~n23871 & ~n23872;
  assign n23874 = ~pi8  & ~n23871;
  assign n23875 = pi8  & ~n23872;
  assign n23876 = pi8  & n23871;
  assign n23877 = ~n56157 & ~n56158;
  assign n23878 = n23267 & n56053;
  assign n23879 = ~n23267 & ~n23275;
  assign n23880 = ~n23267 & n56053;
  assign n23881 = ~n56053 & ~n23275;
  assign n23882 = n23267 & ~n56053;
  assign n23883 = ~n56159 & ~n56160;
  assign n23884 = ~n23275 & ~n23878;
  assign n23885 = ~n23877 & ~n56161;
  assign n23886 = n23258 & n56050;
  assign n23887 = ~n23266 & ~n23886;
  assign n23888 = n17524 & n20085;
  assign n23889 = ~n54183 & n21237;
  assign n23890 = ~n54194 & n55472;
  assign n23891 = ~n54163 & n21269;
  assign n23892 = ~n23890 & ~n23891;
  assign n23893 = ~n23889 & ~n23890;
  assign n23894 = ~n23891 & n23893;
  assign n23895 = ~n23889 & n23892;
  assign n23896 = ~n20085 & n56162;
  assign n23897 = ~n17524 & n56162;
  assign n23898 = ~n23896 & ~n23897;
  assign n23899 = ~n23888 & n56162;
  assign n23900 = pi8  & ~n56163;
  assign n23901 = ~pi8  & n56163;
  assign n23902 = ~n23900 & ~n23901;
  assign n23903 = n23887 & ~n23902;
  assign n23904 = n23254 & ~n23256;
  assign n23905 = ~n23257 & ~n23904;
  assign n23906 = n17544 & n20085;
  assign n23907 = ~n54212 & n55472;
  assign n23908 = ~n54183 & n21269;
  assign n23909 = ~n54194 & n21237;
  assign n23910 = ~n23908 & ~n23909;
  assign n23911 = ~n23907 & ~n23909;
  assign n23912 = ~n23908 & n23911;
  assign n23913 = ~n23907 & n23910;
  assign n23914 = ~n20085 & n56164;
  assign n23915 = ~n17544 & n56164;
  assign n23916 = ~n23914 & ~n23915;
  assign n23917 = ~n23906 & n56164;
  assign n23918 = pi8  & ~n56165;
  assign n23919 = ~pi8  & n56165;
  assign n23920 = ~n23918 & ~n23919;
  assign n23921 = n23905 & ~n23920;
  assign n23922 = n23245 & n56047;
  assign n23923 = ~n23253 & ~n23922;
  assign n23924 = n17041 & n20085;
  assign n23925 = ~n54212 & n21237;
  assign n23926 = ~n54194 & n21269;
  assign n23927 = ~n54240 & n55472;
  assign n23928 = ~n23926 & ~n23927;
  assign n23929 = ~n23925 & ~n23927;
  assign n23930 = ~n23926 & n23929;
  assign n23931 = ~n23925 & n23928;
  assign n23932 = ~n20085 & n56166;
  assign n23933 = ~n17041 & n56166;
  assign n23934 = ~n23932 & ~n23933;
  assign n23935 = ~n23924 & n56166;
  assign n23936 = pi8  & ~n56167;
  assign n23937 = ~pi8  & n56167;
  assign n23938 = ~n23936 & ~n23937;
  assign n23939 = n23923 & ~n23938;
  assign n23940 = n17660 & n20085;
  assign n23941 = ~n54254 & n55472;
  assign n23942 = ~n54212 & n21269;
  assign n23943 = ~n54240 & n21237;
  assign n23944 = ~n23942 & ~n23943;
  assign n23945 = ~n23941 & ~n23943;
  assign n23946 = ~n23942 & n23945;
  assign n23947 = ~n23941 & n23944;
  assign n23948 = ~n23940 & n56168;
  assign n23949 = pi8  & ~n23948;
  assign n23950 = ~n23948 & ~n23949;
  assign n23951 = ~pi8  & ~n23948;
  assign n23952 = pi8  & ~n23949;
  assign n23953 = pi8  & n23948;
  assign n23954 = ~n56169 & ~n56170;
  assign n23955 = n23241 & ~n23243;
  assign n23956 = ~n23244 & ~n23955;
  assign n23957 = ~n23954 & n23956;
  assign n23958 = n17804 & n20085;
  assign n23959 = ~n54254 & n21237;
  assign n23960 = ~n54240 & n21269;
  assign n23961 = ~n54269 & n55472;
  assign n23962 = ~n23960 & ~n23961;
  assign n23963 = ~n23959 & ~n23961;
  assign n23964 = ~n23960 & n23963;
  assign n23965 = ~n23959 & n23962;
  assign n23966 = ~n20085 & n56171;
  assign n23967 = ~n17804 & n56171;
  assign n23968 = ~n23966 & ~n23967;
  assign n23969 = ~n23958 & n56171;
  assign n23970 = pi8  & ~n56172;
  assign n23971 = ~pi8  & n56172;
  assign n23972 = ~n23970 & ~n23971;
  assign n23973 = n23232 & n56044;
  assign n23974 = ~n56044 & ~n23240;
  assign n23975 = ~n23232 & ~n23240;
  assign n23976 = ~n23974 & ~n23975;
  assign n23977 = ~n23240 & ~n23973;
  assign n23978 = ~n23972 & ~n56173;
  assign n23979 = n17939 & n20085;
  assign n23980 = ~n54254 & n21269;
  assign n23981 = ~n54277 & n55472;
  assign n23982 = ~n54269 & n21237;
  assign n23983 = ~n23981 & ~n23982;
  assign n23984 = ~n23980 & n23983;
  assign n23985 = ~n23979 & n23984;
  assign n23986 = pi8  & ~n23985;
  assign n23987 = ~n23985 & ~n23986;
  assign n23988 = ~pi8  & ~n23985;
  assign n23989 = pi8  & ~n23986;
  assign n23990 = pi8  & n23985;
  assign n23991 = ~n56174 & ~n56175;
  assign n23992 = pi11  & ~n56036;
  assign n23993 = ~n56037 & ~n23992;
  assign n23994 = n56037 & n23992;
  assign n23995 = ~n56036 & n23214;
  assign n23996 = ~n56038 & ~n23995;
  assign n23997 = ~n23993 & ~n23994;
  assign n23998 = ~n23991 & n56176;
  assign n23999 = n18056 & n20085;
  assign n24000 = ~n54305 & n55472;
  assign n24001 = ~n54277 & n21237;
  assign n24002 = ~n54269 & n21269;
  assign n24003 = ~n24001 & ~n24002;
  assign n24004 = ~n24000 & ~n24001;
  assign n24005 = ~n24002 & n24004;
  assign n24006 = ~n24000 & n24003;
  assign n24007 = ~n20085 & n56177;
  assign n24008 = ~n18056 & n56177;
  assign n24009 = ~n24007 & ~n24008;
  assign n24010 = ~n23999 & n56177;
  assign n24011 = pi8  & ~n56178;
  assign n24012 = ~pi8  & n56178;
  assign n24013 = ~n24011 & ~n24012;
  assign n24014 = pi11  & n23194;
  assign n24015 = ~n23193 & n24014;
  assign n24016 = n23193 & ~n24014;
  assign n24017 = ~n23195 & n23199;
  assign n24018 = ~n56036 & ~n24017;
  assign n24019 = ~n24015 & ~n24016;
  assign n24020 = ~n24013 & n56179;
  assign n24021 = ~n19275 & n20085;
  assign n24022 = ~n54325 & n21237;
  assign n24023 = ~n54344 & n21269;
  assign n24024 = ~n24022 & ~n24023;
  assign n24025 = ~n24021 & n24024;
  assign n24026 = ~n54325 & n55469;
  assign n24027 = pi8  & ~n24026;
  assign n24028 = pi8  & ~n24025;
  assign n24029 = pi8  & ~n24028;
  assign n24030 = ~n24025 & ~n24028;
  assign n24031 = ~n24029 & ~n24030;
  assign n24032 = n24027 & ~n24031;
  assign n24033 = n24025 & n24027;
  assign n24034 = n18156 & n20085;
  assign n24035 = ~n54305 & n21269;
  assign n24036 = ~n54325 & n55472;
  assign n24037 = ~n54344 & n21237;
  assign n24038 = ~n24036 & ~n24037;
  assign n24039 = ~n24035 & n24038;
  assign n24040 = ~n20085 & n24039;
  assign n24041 = ~n18156 & n24039;
  assign n24042 = ~n24040 & ~n24041;
  assign n24043 = ~n24034 & n24039;
  assign n24044 = pi8  & ~n56181;
  assign n24045 = ~pi8  & n56181;
  assign n24046 = ~n24044 & ~n24045;
  assign n24047 = n56180 & ~n24046;
  assign n24048 = n56180 & ~n56181;
  assign n24049 = n23194 & n56182;
  assign n24050 = n18336 & n20085;
  assign n24051 = ~n54305 & n21237;
  assign n24052 = ~n54277 & n21269;
  assign n24053 = ~n54344 & n55472;
  assign n24054 = ~n24052 & ~n24053;
  assign n24055 = ~n24051 & ~n24053;
  assign n24056 = ~n24052 & n24055;
  assign n24057 = ~n24051 & n24054;
  assign n24058 = ~n24050 & n56183;
  assign n24059 = pi8  & ~n24058;
  assign n24060 = pi8  & ~n24059;
  assign n24061 = pi8  & n24058;
  assign n24062 = ~n24058 & ~n24059;
  assign n24063 = ~pi8  & ~n24058;
  assign n24064 = ~n56184 & ~n56185;
  assign n24065 = ~n23194 & ~n56182;
  assign n24066 = n56182 & ~n24049;
  assign n24067 = ~n23194 & n56182;
  assign n24068 = n23194 & ~n24049;
  assign n24069 = n23194 & ~n56182;
  assign n24070 = ~n56186 & ~n56187;
  assign n24071 = ~n24049 & ~n24065;
  assign n24072 = ~n24064 & ~n56188;
  assign n24073 = ~n24049 & ~n24072;
  assign n24074 = n24013 & ~n56179;
  assign n24075 = ~n24020 & ~n24074;
  assign n24076 = ~n24073 & n24075;
  assign n24077 = ~n24020 & ~n24076;
  assign n24078 = n23991 & ~n56176;
  assign n24079 = ~n23991 & ~n23998;
  assign n24080 = ~n23991 & ~n56176;
  assign n24081 = n56176 & ~n23998;
  assign n24082 = n23991 & n56176;
  assign n24083 = ~n56189 & ~n56190;
  assign n24084 = ~n23998 & ~n24078;
  assign n24085 = ~n24077 & ~n56191;
  assign n24086 = ~n23998 & ~n24085;
  assign n24087 = n23972 & n56173;
  assign n24088 = ~n23978 & ~n24087;
  assign n24089 = ~n24086 & n24088;
  assign n24090 = ~n23978 & ~n24089;
  assign n24091 = n23954 & ~n23956;
  assign n24092 = ~n23954 & ~n23957;
  assign n24093 = ~n23954 & ~n23956;
  assign n24094 = n23956 & ~n23957;
  assign n24095 = n23954 & n23956;
  assign n24096 = ~n56192 & ~n56193;
  assign n24097 = ~n23957 & ~n24091;
  assign n24098 = ~n24090 & ~n56194;
  assign n24099 = ~n23957 & ~n24098;
  assign n24100 = ~n23923 & n23938;
  assign n24101 = n23923 & ~n23939;
  assign n24102 = n23923 & n23938;
  assign n24103 = ~n23938 & ~n23939;
  assign n24104 = ~n23923 & ~n23938;
  assign n24105 = ~n56195 & ~n56196;
  assign n24106 = ~n23939 & ~n24100;
  assign n24107 = ~n24099 & ~n56197;
  assign n24108 = ~n23939 & ~n24107;
  assign n24109 = ~n23905 & n23920;
  assign n24110 = n23905 & ~n23921;
  assign n24111 = n23905 & n23920;
  assign n24112 = ~n23920 & ~n23921;
  assign n24113 = ~n23905 & ~n23920;
  assign n24114 = ~n56198 & ~n56199;
  assign n24115 = ~n23921 & ~n24109;
  assign n24116 = ~n24108 & ~n56200;
  assign n24117 = ~n23921 & ~n24116;
  assign n24118 = ~n23887 & n23902;
  assign n24119 = ~n23903 & ~n24118;
  assign n24120 = ~n24117 & n24119;
  assign n24121 = ~n23903 & ~n24120;
  assign n24122 = n23877 & n56161;
  assign n24123 = ~n23877 & ~n23885;
  assign n24124 = ~n56161 & ~n23885;
  assign n24125 = ~n24123 & ~n24124;
  assign n24126 = ~n23885 & ~n24122;
  assign n24127 = ~n24121 & ~n56201;
  assign n24128 = ~n23885 & ~n24127;
  assign n24129 = n23858 & n56156;
  assign n24130 = ~n23858 & ~n23864;
  assign n24131 = ~n23858 & n56156;
  assign n24132 = ~n56156 & ~n23864;
  assign n24133 = n23858 & ~n56156;
  assign n24134 = ~n56202 & ~n56203;
  assign n24135 = ~n23864 & ~n24129;
  assign n24136 = ~n24128 & ~n56204;
  assign n24137 = ~n23864 & ~n24136;
  assign n24138 = n23840 & ~n23842;
  assign n24139 = ~n23840 & ~n23843;
  assign n24140 = ~n23840 & ~n23842;
  assign n24141 = n23842 & ~n23843;
  assign n24142 = n23840 & n23842;
  assign n24143 = ~n56205 & ~n56206;
  assign n24144 = ~n23843 & ~n24138;
  assign n24145 = ~n24137 & ~n56207;
  assign n24146 = ~n23843 & ~n24145;
  assign n24147 = ~n23809 & n23824;
  assign n24148 = n23809 & ~n23825;
  assign n24149 = n23809 & n23824;
  assign n24150 = ~n23824 & ~n23825;
  assign n24151 = ~n23809 & ~n23824;
  assign n24152 = ~n56208 & ~n56209;
  assign n24153 = ~n23825 & ~n24147;
  assign n24154 = ~n24146 & ~n56210;
  assign n24155 = ~n23825 & ~n24154;
  assign n24156 = ~n23789 & n23806;
  assign n24157 = n23789 & ~n23807;
  assign n24158 = n23789 & n23806;
  assign n24159 = ~n23806 & ~n23807;
  assign n24160 = ~n23789 & ~n23806;
  assign n24161 = ~n56211 & ~n56212;
  assign n24162 = ~n23807 & ~n24156;
  assign n24163 = ~n24155 & ~n56213;
  assign n24164 = ~n23807 & ~n24163;
  assign n24165 = ~n23771 & n23786;
  assign n24166 = ~n23787 & ~n24165;
  assign n24167 = ~n24164 & n24166;
  assign n24168 = ~n23787 & ~n24167;
  assign n24169 = n23763 & n56143;
  assign n24170 = ~n23763 & ~n23769;
  assign n24171 = ~n23763 & n56143;
  assign n24172 = ~n56143 & ~n23769;
  assign n24173 = n23763 & ~n56143;
  assign n24174 = ~n56214 & ~n56215;
  assign n24175 = ~n23769 & ~n24169;
  assign n24176 = ~n24168 & ~n56216;
  assign n24177 = ~n23769 & ~n24176;
  assign n24178 = n23740 & n56139;
  assign n24179 = ~n23740 & ~n23748;
  assign n24180 = ~n56139 & ~n23748;
  assign n24181 = ~n24179 & ~n24180;
  assign n24182 = ~n23748 & ~n24178;
  assign n24183 = ~n24177 & ~n56217;
  assign n24184 = ~n23748 & ~n24183;
  assign n24185 = n23722 & ~n23724;
  assign n24186 = ~n23722 & ~n23725;
  assign n24187 = ~n23722 & ~n23724;
  assign n24188 = n23724 & ~n23725;
  assign n24189 = n23722 & n23724;
  assign n24190 = ~n56218 & ~n56219;
  assign n24191 = ~n23725 & ~n24185;
  assign n24192 = ~n24184 & ~n56220;
  assign n24193 = ~n23725 & ~n24192;
  assign n24194 = ~n23691 & n23706;
  assign n24195 = n23691 & ~n23707;
  assign n24196 = n23691 & n23706;
  assign n24197 = ~n23706 & ~n23707;
  assign n24198 = ~n23691 & ~n23706;
  assign n24199 = ~n56221 & ~n56222;
  assign n24200 = ~n23707 & ~n24194;
  assign n24201 = ~n24193 & ~n56223;
  assign n24202 = ~n23707 & ~n24201;
  assign n24203 = ~n23673 & n23688;
  assign n24204 = n23673 & ~n23689;
  assign n24205 = n23673 & n23688;
  assign n24206 = ~n23688 & ~n23689;
  assign n24207 = ~n23673 & ~n23688;
  assign n24208 = ~n56224 & ~n56225;
  assign n24209 = ~n23689 & ~n24203;
  assign n24210 = ~n24202 & ~n56226;
  assign n24211 = ~n23689 & ~n24210;
  assign n24212 = ~n23655 & n23670;
  assign n24213 = ~n23671 & ~n24212;
  assign n24214 = ~n24211 & n24213;
  assign n24215 = ~n23671 & ~n24214;
  assign n24216 = n23645 & n56124;
  assign n24217 = ~n23645 & ~n23653;
  assign n24218 = ~n56124 & ~n23653;
  assign n24219 = ~n24217 & ~n24218;
  assign n24220 = ~n23653 & ~n24216;
  assign n24221 = ~n24215 & ~n56227;
  assign n24222 = ~n23653 & ~n24221;
  assign n24223 = n23627 & ~n23629;
  assign n24224 = ~n23627 & ~n23630;
  assign n24225 = ~n23627 & ~n23629;
  assign n24226 = n23629 & ~n23630;
  assign n24227 = n23627 & n23629;
  assign n24228 = ~n56228 & ~n56229;
  assign n24229 = ~n23630 & ~n24223;
  assign n24230 = ~n24222 & ~n56230;
  assign n24231 = ~n23630 & ~n24230;
  assign n24232 = ~n23596 & n23611;
  assign n24233 = n23596 & ~n23612;
  assign n24234 = n23596 & n23611;
  assign n24235 = ~n23611 & ~n23612;
  assign n24236 = ~n23596 & ~n23611;
  assign n24237 = ~n56231 & ~n56232;
  assign n24238 = ~n23612 & ~n24232;
  assign n24239 = ~n24231 & ~n56233;
  assign n24240 = ~n23612 & ~n24239;
  assign n24241 = ~n23578 & n23593;
  assign n24242 = n23578 & ~n23594;
  assign n24243 = n23578 & n23593;
  assign n24244 = ~n23593 & ~n23594;
  assign n24245 = ~n23578 & ~n23593;
  assign n24246 = ~n56234 & ~n56235;
  assign n24247 = ~n23594 & ~n24241;
  assign n24248 = ~n24240 & ~n56236;
  assign n24249 = ~n23594 & ~n24248;
  assign n24250 = ~n23560 & n23575;
  assign n24251 = n23560 & ~n23576;
  assign n24252 = n23560 & n23575;
  assign n24253 = ~n23575 & ~n23576;
  assign n24254 = ~n23560 & ~n23575;
  assign n24255 = ~n56237 & ~n56238;
  assign n24256 = ~n23576 & ~n24250;
  assign n24257 = ~n24249 & ~n56239;
  assign n24258 = ~n23576 & ~n24257;
  assign n24259 = ~n23542 & n23557;
  assign n24260 = n23542 & ~n23558;
  assign n24261 = n23542 & n23557;
  assign n24262 = ~n23557 & ~n23558;
  assign n24263 = ~n23542 & ~n23557;
  assign n24264 = ~n56240 & ~n56241;
  assign n24265 = ~n23558 & ~n24259;
  assign n24266 = ~n24258 & ~n56242;
  assign n24267 = ~n23558 & ~n24266;
  assign n24268 = ~n23524 & n23539;
  assign n24269 = n23524 & ~n23540;
  assign n24270 = n23524 & n23539;
  assign n24271 = ~n23539 & ~n23540;
  assign n24272 = ~n23524 & ~n23539;
  assign n24273 = ~n56243 & ~n56244;
  assign n24274 = ~n23540 & ~n24268;
  assign n24275 = ~n24267 & ~n56245;
  assign n24276 = ~n23540 & ~n24275;
  assign n24277 = ~n23506 & n23521;
  assign n24278 = n23506 & ~n23522;
  assign n24279 = n23506 & n23521;
  assign n24280 = ~n23521 & ~n23522;
  assign n24281 = ~n23506 & ~n23521;
  assign n24282 = ~n56246 & ~n56247;
  assign n24283 = ~n23522 & ~n24277;
  assign n24284 = ~n24276 & ~n56248;
  assign n24285 = ~n23522 & ~n24284;
  assign n24286 = ~n23488 & n23503;
  assign n24287 = n23488 & ~n23504;
  assign n24288 = n23488 & n23503;
  assign n24289 = ~n23503 & ~n23504;
  assign n24290 = ~n23488 & ~n23503;
  assign n24291 = ~n56249 & ~n56250;
  assign n24292 = ~n23504 & ~n24286;
  assign n24293 = ~n24285 & ~n56251;
  assign n24294 = ~n23504 & ~n24293;
  assign n24295 = n23449 & ~n23452;
  assign n24296 = ~n23451 & n24295;
  assign n24297 = n23449 & n56098;
  assign n24298 = ~n23455 & ~n56252;
  assign n24299 = ~n24294 & n24298;
  assign n24300 = n77 & n11242;
  assign n24301 = ~n53650 & n21969;
  assign n24302 = n53439 & ~n53440;
  assign n24303 = ~n2325 & n24302;
  assign n24304 = ~n53634 & n23459;
  assign n24305 = ~n24303 & ~n24304;
  assign n24306 = ~n24301 & ~n24304;
  assign n24307 = ~n24303 & n24306;
  assign n24308 = ~n24301 & n24305;
  assign n24309 = ~n24300 & n56253;
  assign n24310 = pi5  & ~n24309;
  assign n24311 = ~n24309 & ~n24310;
  assign n24312 = ~pi5  & ~n24309;
  assign n24313 = pi5  & ~n24310;
  assign n24314 = pi5  & n24309;
  assign n24315 = ~n56254 & ~n56255;
  assign n24316 = n24294 & ~n24298;
  assign n24317 = ~n24294 & ~n24299;
  assign n24318 = n24298 & ~n24299;
  assign n24319 = ~n24317 & ~n24318;
  assign n24320 = ~n24299 & ~n24316;
  assign n24321 = ~n24315 & ~n56256;
  assign n24322 = ~n24299 & ~n24321;
  assign n24323 = ~n23471 & n56100;
  assign n24324 = ~n23477 & ~n24323;
  assign n24325 = ~n24322 & n24324;
  assign n24326 = n24315 & ~n24318;
  assign n24327 = ~n24317 & n24326;
  assign n24328 = n24315 & n56256;
  assign n24329 = ~n24321 & ~n56257;
  assign n24330 = ~pi0  & ~pi1 ;
  assign n24331 = pi1  & ~pi2 ;
  assign n24332 = ~pi1  & pi2 ;
  assign n24333 = ~pi1  & ~pi2 ;
  assign n24334 = pi1  & pi2 ;
  assign n24335 = ~n24333 & ~n24334;
  assign n24336 = ~n24331 & ~n24332;
  assign n24337 = n24330 & n56258;
  assign n24338 = pi0  & n56258;
  assign n24339 = ~n10547 & n24338;
  assign n24340 = ~n24337 & ~n24339;
  assign n24341 = ~n2325 & n24337;
  assign n24342 = n10551 & n24338;
  assign n24343 = ~n24341 & ~n24342;
  assign n24344 = ~n2325 & ~n24340;
  assign n24345 = pi2  & ~n56259;
  assign n24346 = ~n56259 & ~n24345;
  assign n24347 = ~pi2  & ~n56259;
  assign n24348 = pi2  & ~n24345;
  assign n24349 = pi2  & n56259;
  assign n24350 = ~n56260 & ~n56261;
  assign n24351 = n77 & n11286;
  assign n24352 = ~n53650 & n23459;
  assign n24353 = ~n53657 & n21969;
  assign n24354 = ~n53634 & n24302;
  assign n24355 = ~n24353 & ~n24354;
  assign n24356 = ~n24352 & ~n24353;
  assign n24357 = ~n24354 & n24356;
  assign n24358 = ~n24352 & n24355;
  assign n24359 = ~n24351 & n56262;
  assign n24360 = pi5  & ~n24359;
  assign n24361 = pi5  & ~n24360;
  assign n24362 = pi5  & n24359;
  assign n24363 = ~n24359 & ~n24360;
  assign n24364 = ~pi5  & ~n24359;
  assign n24365 = ~n56263 & ~n56264;
  assign n24366 = ~n24350 & ~n24365;
  assign n24367 = n24350 & n24365;
  assign n24368 = n24285 & n56251;
  assign n24369 = ~n24285 & ~n24293;
  assign n24370 = ~n24285 & n56251;
  assign n24371 = ~n56251 & ~n24293;
  assign n24372 = n24285 & ~n56251;
  assign n24373 = ~n56265 & ~n56266;
  assign n24374 = ~n24293 & ~n24368;
  assign n24375 = ~n24367 & ~n56267;
  assign n24376 = ~n24350 & ~n24366;
  assign n24377 = ~n24365 & ~n24366;
  assign n24378 = ~n24376 & ~n24377;
  assign n24379 = ~n24366 & ~n24367;
  assign n24380 = ~n56267 & ~n56268;
  assign n24381 = ~n24366 & ~n24380;
  assign n24382 = ~n24366 & ~n24375;
  assign n24383 = n24329 & ~n56269;
  assign n24384 = n77 & n11213;
  assign n24385 = ~n53650 & n24302;
  assign n24386 = ~n53685 & n21969;
  assign n24387 = ~n53657 & n23459;
  assign n24388 = ~n24386 & ~n24387;
  assign n24389 = ~n24385 & n24388;
  assign n24390 = ~n24384 & n24389;
  assign n24391 = pi5  & ~n24390;
  assign n24392 = ~n24390 & ~n24391;
  assign n24393 = ~pi5  & ~n24390;
  assign n24394 = pi5  & ~n24391;
  assign n24395 = pi5  & n24390;
  assign n24396 = ~n56270 & ~n56271;
  assign n24397 = n24276 & n56248;
  assign n24398 = ~n24276 & ~n24284;
  assign n24399 = ~n24276 & n56248;
  assign n24400 = ~n56248 & ~n24284;
  assign n24401 = n24276 & ~n56248;
  assign n24402 = ~n56272 & ~n56273;
  assign n24403 = ~n24284 & ~n24397;
  assign n24404 = ~n24396 & ~n56274;
  assign n24405 = n77 & n11380;
  assign n24406 = ~n53685 & n23459;
  assign n24407 = ~n53657 & n24302;
  assign n24408 = ~n53712 & n21969;
  assign n24409 = ~n24407 & ~n24408;
  assign n24410 = ~n24406 & ~n24408;
  assign n24411 = ~n24407 & n24410;
  assign n24412 = ~n24406 & n24409;
  assign n24413 = ~n24405 & n56275;
  assign n24414 = pi5  & ~n24413;
  assign n24415 = ~n24413 & ~n24414;
  assign n24416 = ~pi5  & ~n24413;
  assign n24417 = pi5  & ~n24414;
  assign n24418 = pi5  & n24413;
  assign n24419 = ~n56276 & ~n56277;
  assign n24420 = n24267 & n56245;
  assign n24421 = ~n24267 & ~n24275;
  assign n24422 = ~n56245 & ~n24275;
  assign n24423 = ~n24421 & ~n24422;
  assign n24424 = ~n24275 & ~n24420;
  assign n24425 = ~n24419 & ~n56278;
  assign n24426 = n77 & n11360;
  assign n24427 = ~n53685 & n24302;
  assign n24428 = ~n53741 & n21969;
  assign n24429 = ~n53712 & n23459;
  assign n24430 = ~n24428 & ~n24429;
  assign n24431 = ~n24427 & ~n24428;
  assign n24432 = ~n24429 & n24431;
  assign n24433 = ~n24427 & n24430;
  assign n24434 = ~n24426 & n56279;
  assign n24435 = pi5  & ~n24434;
  assign n24436 = ~n24434 & ~n24435;
  assign n24437 = ~pi5  & ~n24434;
  assign n24438 = pi5  & ~n24435;
  assign n24439 = pi5  & n24434;
  assign n24440 = ~n56280 & ~n56281;
  assign n24441 = n24258 & n56242;
  assign n24442 = ~n24258 & ~n24266;
  assign n24443 = ~n56242 & ~n24266;
  assign n24444 = ~n24442 & ~n24443;
  assign n24445 = ~n24266 & ~n24441;
  assign n24446 = ~n24440 & ~n56282;
  assign n24447 = n77 & n11889;
  assign n24448 = ~n53712 & n24302;
  assign n24449 = ~n53774 & n21969;
  assign n24450 = ~n53741 & n23459;
  assign n24451 = ~n24449 & ~n24450;
  assign n24452 = ~n24448 & ~n24449;
  assign n24453 = ~n24450 & n24452;
  assign n24454 = ~n24448 & n24451;
  assign n24455 = ~n24447 & n56283;
  assign n24456 = pi5  & ~n24455;
  assign n24457 = ~n24455 & ~n24456;
  assign n24458 = ~pi5  & ~n24455;
  assign n24459 = pi5  & ~n24456;
  assign n24460 = pi5  & n24455;
  assign n24461 = ~n56284 & ~n56285;
  assign n24462 = n24249 & n56239;
  assign n24463 = ~n24249 & ~n24257;
  assign n24464 = ~n24249 & n56239;
  assign n24465 = ~n56239 & ~n24257;
  assign n24466 = n24249 & ~n56239;
  assign n24467 = ~n56286 & ~n56287;
  assign n24468 = ~n24257 & ~n24462;
  assign n24469 = ~n24461 & ~n56288;
  assign n24470 = n77 & n11913;
  assign n24471 = ~n53774 & n23459;
  assign n24472 = ~n53799 & n21969;
  assign n24473 = ~n53741 & n24302;
  assign n24474 = ~n24472 & ~n24473;
  assign n24475 = ~n24471 & ~n24472;
  assign n24476 = ~n24473 & n24475;
  assign n24477 = ~n24471 & n24474;
  assign n24478 = ~n24470 & n56289;
  assign n24479 = pi5  & ~n24478;
  assign n24480 = ~n24478 & ~n24479;
  assign n24481 = ~pi5  & ~n24478;
  assign n24482 = pi5  & ~n24479;
  assign n24483 = pi5  & n24478;
  assign n24484 = ~n56290 & ~n56291;
  assign n24485 = n24240 & n56236;
  assign n24486 = ~n24240 & ~n24248;
  assign n24487 = ~n24240 & n56236;
  assign n24488 = ~n56236 & ~n24248;
  assign n24489 = n24240 & ~n56236;
  assign n24490 = ~n56292 & ~n56293;
  assign n24491 = ~n24248 & ~n24485;
  assign n24492 = ~n24484 & ~n56294;
  assign n24493 = n77 & n12690;
  assign n24494 = ~n53774 & n24302;
  assign n24495 = ~n53819 & n21969;
  assign n24496 = ~n53799 & n23459;
  assign n24497 = ~n24495 & ~n24496;
  assign n24498 = ~n24494 & ~n24495;
  assign n24499 = ~n24496 & n24498;
  assign n24500 = ~n24494 & n24497;
  assign n24501 = ~n24493 & n56295;
  assign n24502 = pi5  & ~n24501;
  assign n24503 = ~n24501 & ~n24502;
  assign n24504 = ~pi5  & ~n24501;
  assign n24505 = pi5  & ~n24502;
  assign n24506 = pi5  & n24501;
  assign n24507 = ~n56296 & ~n56297;
  assign n24508 = n24231 & n56233;
  assign n24509 = ~n24231 & ~n24239;
  assign n24510 = ~n56233 & ~n24239;
  assign n24511 = ~n24509 & ~n24510;
  assign n24512 = ~n24239 & ~n24508;
  assign n24513 = ~n24507 & ~n56298;
  assign n24514 = n24222 & n56230;
  assign n24515 = ~n24230 & ~n24514;
  assign n24516 = n77 & n12550;
  assign n24517 = ~n53819 & n23459;
  assign n24518 = ~n53845 & n21969;
  assign n24519 = ~n53799 & n24302;
  assign n24520 = ~n24518 & ~n24519;
  assign n24521 = ~n24517 & ~n24518;
  assign n24522 = ~n24519 & n24521;
  assign n24523 = ~n24517 & n24520;
  assign n24524 = ~n77 & n56299;
  assign n24525 = ~n12550 & n56299;
  assign n24526 = ~n24524 & ~n24525;
  assign n24527 = ~n24516 & n56299;
  assign n24528 = pi5  & ~n56300;
  assign n24529 = ~pi5  & n56300;
  assign n24530 = ~n24528 & ~n24529;
  assign n24531 = n24515 & ~n24530;
  assign n24532 = n24215 & n56227;
  assign n24533 = ~n24221 & ~n24532;
  assign n24534 = n77 & n12938;
  assign n24535 = ~n53819 & n24302;
  assign n24536 = ~n53860 & n21969;
  assign n24537 = ~n53845 & n23459;
  assign n24538 = ~n24536 & ~n24537;
  assign n24539 = ~n24535 & ~n24536;
  assign n24540 = ~n24537 & n24539;
  assign n24541 = ~n24535 & n24538;
  assign n24542 = ~n77 & n56301;
  assign n24543 = ~n12938 & n56301;
  assign n24544 = ~n24542 & ~n24543;
  assign n24545 = ~n24534 & n56301;
  assign n24546 = pi5  & ~n56302;
  assign n24547 = ~pi5  & n56302;
  assign n24548 = ~n24546 & ~n24547;
  assign n24549 = n24533 & ~n24548;
  assign n24550 = n77 & n12918;
  assign n24551 = ~n53860 & n23459;
  assign n24552 = ~n53888 & n21969;
  assign n24553 = ~n53845 & n24302;
  assign n24554 = ~n24552 & ~n24553;
  assign n24555 = ~n24551 & ~n24552;
  assign n24556 = ~n24553 & n24555;
  assign n24557 = ~n24551 & n24554;
  assign n24558 = ~n24550 & n56303;
  assign n24559 = pi5  & ~n24558;
  assign n24560 = ~n24558 & ~n24559;
  assign n24561 = ~pi5  & ~n24558;
  assign n24562 = pi5  & ~n24559;
  assign n24563 = pi5  & n24558;
  assign n24564 = ~n56304 & ~n56305;
  assign n24565 = n24211 & ~n24213;
  assign n24566 = ~n24214 & ~n24565;
  assign n24567 = ~n24564 & n24566;
  assign n24568 = n77 & n13336;
  assign n24569 = ~n53888 & n23459;
  assign n24570 = ~n53907 & n21969;
  assign n24571 = ~n53860 & n24302;
  assign n24572 = ~n24570 & ~n24571;
  assign n24573 = ~n24569 & ~n24570;
  assign n24574 = ~n24571 & n24573;
  assign n24575 = ~n24569 & n24572;
  assign n24576 = ~n24568 & n56306;
  assign n24577 = pi5  & ~n24576;
  assign n24578 = ~n24576 & ~n24577;
  assign n24579 = ~pi5  & ~n24576;
  assign n24580 = pi5  & ~n24577;
  assign n24581 = pi5  & n24576;
  assign n24582 = ~n56307 & ~n56308;
  assign n24583 = n24202 & n56226;
  assign n24584 = ~n24202 & ~n24210;
  assign n24585 = ~n56226 & ~n24210;
  assign n24586 = ~n24584 & ~n24585;
  assign n24587 = ~n24210 & ~n24583;
  assign n24588 = ~n24582 & ~n56309;
  assign n24589 = n77 & n13360;
  assign n24590 = ~n53907 & n23459;
  assign n24591 = ~n53930 & n21969;
  assign n24592 = ~n53888 & n24302;
  assign n24593 = ~n24591 & ~n24592;
  assign n24594 = ~n24590 & ~n24591;
  assign n24595 = ~n24592 & n24594;
  assign n24596 = ~n24590 & n24593;
  assign n24597 = ~n24589 & n56310;
  assign n24598 = pi5  & ~n24597;
  assign n24599 = ~n24597 & ~n24598;
  assign n24600 = ~pi5  & ~n24597;
  assign n24601 = pi5  & ~n24598;
  assign n24602 = pi5  & n24597;
  assign n24603 = ~n56311 & ~n56312;
  assign n24604 = n24193 & n56223;
  assign n24605 = ~n24193 & ~n24201;
  assign n24606 = ~n24193 & n56223;
  assign n24607 = ~n56223 & ~n24201;
  assign n24608 = n24193 & ~n56223;
  assign n24609 = ~n56313 & ~n56314;
  assign n24610 = ~n24201 & ~n24604;
  assign n24611 = ~n24603 & ~n56315;
  assign n24612 = n24184 & n56220;
  assign n24613 = ~n24192 & ~n24612;
  assign n24614 = n77 & n14263;
  assign n24615 = ~n53930 & n23459;
  assign n24616 = ~n53962 & n21969;
  assign n24617 = ~n53907 & n24302;
  assign n24618 = ~n24616 & ~n24617;
  assign n24619 = ~n24615 & ~n24616;
  assign n24620 = ~n24617 & n24619;
  assign n24621 = ~n24615 & n24618;
  assign n24622 = ~n77 & n56316;
  assign n24623 = ~n14263 & n56316;
  assign n24624 = ~n24622 & ~n24623;
  assign n24625 = ~n24614 & n56316;
  assign n24626 = pi5  & ~n56317;
  assign n24627 = ~pi5  & n56317;
  assign n24628 = ~n24626 & ~n24627;
  assign n24629 = n24613 & ~n24628;
  assign n24630 = n24177 & n56217;
  assign n24631 = ~n24183 & ~n24630;
  assign n24632 = n77 & n14020;
  assign n24633 = ~n53962 & n23459;
  assign n24634 = ~n53970 & n21969;
  assign n24635 = ~n53930 & n24302;
  assign n24636 = ~n24634 & ~n24635;
  assign n24637 = ~n24633 & ~n24634;
  assign n24638 = ~n24635 & n24637;
  assign n24639 = ~n24633 & n24636;
  assign n24640 = ~n77 & n56318;
  assign n24641 = ~n14020 & n56318;
  assign n24642 = ~n24640 & ~n24641;
  assign n24643 = ~n24632 & n56318;
  assign n24644 = pi5  & ~n56319;
  assign n24645 = ~pi5  & n56319;
  assign n24646 = ~n24644 & ~n24645;
  assign n24647 = n24631 & ~n24646;
  assign n24648 = n24168 & n56216;
  assign n24649 = ~n24176 & ~n24648;
  assign n24650 = n77 & n14708;
  assign n24651 = ~n54005 & n21969;
  assign n24652 = ~n53970 & n23459;
  assign n24653 = ~n53962 & n24302;
  assign n24654 = ~n24652 & ~n24653;
  assign n24655 = ~n24651 & ~n24652;
  assign n24656 = ~n24653 & n24655;
  assign n24657 = ~n24651 & n24654;
  assign n24658 = ~n77 & n56320;
  assign n24659 = ~n14708 & n56320;
  assign n24660 = ~n24658 & ~n24659;
  assign n24661 = ~n24650 & n56320;
  assign n24662 = pi5  & ~n56321;
  assign n24663 = ~pi5  & n56321;
  assign n24664 = ~n24662 & ~n24663;
  assign n24665 = n24649 & ~n24664;
  assign n24666 = n77 & n14688;
  assign n24667 = ~n54005 & n23459;
  assign n24668 = ~n54034 & n21969;
  assign n24669 = ~n53970 & n24302;
  assign n24670 = ~n24668 & ~n24669;
  assign n24671 = ~n24667 & ~n24668;
  assign n24672 = ~n24669 & n24671;
  assign n24673 = ~n24667 & n24670;
  assign n24674 = ~n24666 & n56322;
  assign n24675 = pi5  & ~n24674;
  assign n24676 = ~n24674 & ~n24675;
  assign n24677 = ~pi5  & ~n24674;
  assign n24678 = pi5  & ~n24675;
  assign n24679 = pi5  & n24674;
  assign n24680 = ~n56323 & ~n56324;
  assign n24681 = n24164 & ~n24166;
  assign n24682 = ~n24167 & ~n24681;
  assign n24683 = ~n24680 & n24682;
  assign n24684 = n77 & n15195;
  assign n24685 = ~n54050 & n21969;
  assign n24686 = ~n54005 & n24302;
  assign n24687 = ~n54034 & n23459;
  assign n24688 = ~n24686 & ~n24687;
  assign n24689 = ~n24685 & ~n24687;
  assign n24690 = ~n24686 & n24689;
  assign n24691 = ~n24685 & n24688;
  assign n24692 = ~n24684 & n56325;
  assign n24693 = pi5  & ~n24692;
  assign n24694 = ~n24692 & ~n24693;
  assign n24695 = ~pi5  & ~n24692;
  assign n24696 = pi5  & ~n24693;
  assign n24697 = pi5  & n24692;
  assign n24698 = ~n56326 & ~n56327;
  assign n24699 = n24155 & n56213;
  assign n24700 = ~n24155 & ~n24163;
  assign n24701 = ~n24155 & n56213;
  assign n24702 = ~n56213 & ~n24163;
  assign n24703 = n24155 & ~n56213;
  assign n24704 = ~n56328 & ~n56329;
  assign n24705 = ~n24163 & ~n24699;
  assign n24706 = ~n24698 & ~n56330;
  assign n24707 = n77 & n15219;
  assign n24708 = ~n54050 & n23459;
  assign n24709 = ~n54034 & n24302;
  assign n24710 = ~n54073 & n21969;
  assign n24711 = ~n24709 & ~n24710;
  assign n24712 = ~n24708 & ~n24710;
  assign n24713 = ~n24709 & n24712;
  assign n24714 = ~n24708 & n24711;
  assign n24715 = ~n24707 & n56331;
  assign n24716 = pi5  & ~n24715;
  assign n24717 = ~n24715 & ~n24716;
  assign n24718 = ~pi5  & ~n24715;
  assign n24719 = pi5  & ~n24716;
  assign n24720 = pi5  & n24715;
  assign n24721 = ~n56332 & ~n56333;
  assign n24722 = n24146 & n56210;
  assign n24723 = ~n24146 & ~n24154;
  assign n24724 = ~n56210 & ~n24154;
  assign n24725 = ~n24723 & ~n24724;
  assign n24726 = ~n24154 & ~n24722;
  assign n24727 = ~n24721 & ~n56334;
  assign n24728 = n24137 & n56207;
  assign n24729 = ~n24145 & ~n24728;
  assign n24730 = n77 & n16138;
  assign n24731 = ~n54098 & n21969;
  assign n24732 = ~n54050 & n24302;
  assign n24733 = ~n54073 & n23459;
  assign n24734 = ~n24732 & ~n24733;
  assign n24735 = ~n24731 & ~n24733;
  assign n24736 = ~n24732 & n24735;
  assign n24737 = ~n24731 & n24734;
  assign n24738 = ~n77 & n56335;
  assign n24739 = ~n16138 & n56335;
  assign n24740 = ~n24738 & ~n24739;
  assign n24741 = ~n24730 & n56335;
  assign n24742 = pi5  & ~n56336;
  assign n24743 = ~pi5  & n56336;
  assign n24744 = ~n24742 & ~n24743;
  assign n24745 = n24729 & ~n24744;
  assign n24746 = n24128 & n56204;
  assign n24747 = ~n24136 & ~n24746;
  assign n24748 = n77 & n15779;
  assign n24749 = ~n54098 & n23459;
  assign n24750 = ~n54119 & n21969;
  assign n24751 = ~n54073 & n24302;
  assign n24752 = ~n24750 & ~n24751;
  assign n24753 = ~n24749 & ~n24750;
  assign n24754 = ~n24751 & n24753;
  assign n24755 = ~n24749 & ~n24751;
  assign n24756 = ~n24750 & n24755;
  assign n24757 = ~n24749 & n24752;
  assign n24758 = ~n77 & n56337;
  assign n24759 = ~n15779 & n56337;
  assign n24760 = ~n24758 & ~n24759;
  assign n24761 = ~n24748 & n56337;
  assign n24762 = pi5  & ~n56338;
  assign n24763 = ~pi5  & n56338;
  assign n24764 = ~n24762 & ~n24763;
  assign n24765 = n24747 & ~n24764;
  assign n24766 = n24121 & n56201;
  assign n24767 = ~n24127 & ~n24766;
  assign n24768 = n77 & n16547;
  assign n24769 = ~n54119 & n23459;
  assign n24770 = ~n54098 & n24302;
  assign n24771 = ~n54132 & n21969;
  assign n24772 = ~n24770 & ~n24771;
  assign n24773 = ~n24769 & ~n24771;
  assign n24774 = ~n24770 & n24773;
  assign n24775 = ~n24769 & n24772;
  assign n24776 = ~n77 & n56339;
  assign n24777 = ~n16547 & n56339;
  assign n24778 = ~n24776 & ~n24777;
  assign n24779 = ~n24768 & n56339;
  assign n24780 = pi5  & ~n56340;
  assign n24781 = ~pi5  & n56340;
  assign n24782 = ~n24780 & ~n24781;
  assign n24783 = n24767 & ~n24782;
  assign n24784 = n77 & n16772;
  assign n24785 = ~n54154 & n21969;
  assign n24786 = ~n54119 & n24302;
  assign n24787 = ~n54132 & n23459;
  assign n24788 = ~n24786 & ~n24787;
  assign n24789 = ~n24785 & ~n24787;
  assign n24790 = ~n24786 & n24789;
  assign n24791 = ~n24785 & n24788;
  assign n24792 = ~n24784 & n56341;
  assign n24793 = pi5  & ~n24792;
  assign n24794 = ~n24792 & ~n24793;
  assign n24795 = ~pi5  & ~n24792;
  assign n24796 = pi5  & ~n24793;
  assign n24797 = pi5  & n24792;
  assign n24798 = ~n56342 & ~n56343;
  assign n24799 = n24117 & ~n24119;
  assign n24800 = ~n24120 & ~n24799;
  assign n24801 = ~n24798 & n24800;
  assign n24802 = n77 & n16522;
  assign n24803 = ~n54154 & n23459;
  assign n24804 = ~n54132 & n24302;
  assign n24805 = ~n54163 & n21969;
  assign n24806 = ~n24804 & ~n24805;
  assign n24807 = ~n24803 & ~n24805;
  assign n24808 = ~n24804 & n24807;
  assign n24809 = ~n24803 & n24806;
  assign n24810 = ~n24802 & n56344;
  assign n24811 = pi5  & ~n24810;
  assign n24812 = ~n24810 & ~n24811;
  assign n24813 = ~pi5  & ~n24810;
  assign n24814 = pi5  & ~n24811;
  assign n24815 = pi5  & n24810;
  assign n24816 = ~n56345 & ~n56346;
  assign n24817 = n24108 & n56200;
  assign n24818 = ~n24108 & ~n24116;
  assign n24819 = ~n56200 & ~n24116;
  assign n24820 = ~n24818 & ~n24819;
  assign n24821 = ~n24116 & ~n24817;
  assign n24822 = ~n24816 & ~n56347;
  assign n24823 = n77 & n17072;
  assign n24824 = ~n54154 & n24302;
  assign n24825 = ~n54183 & n21969;
  assign n24826 = ~n54163 & n23459;
  assign n24827 = ~n24825 & ~n24826;
  assign n24828 = ~n24824 & n24827;
  assign n24829 = ~n24823 & n24828;
  assign n24830 = pi5  & ~n24829;
  assign n24831 = ~n24829 & ~n24830;
  assign n24832 = ~pi5  & ~n24829;
  assign n24833 = pi5  & ~n24830;
  assign n24834 = pi5  & n24829;
  assign n24835 = ~n56348 & ~n56349;
  assign n24836 = n24099 & n56197;
  assign n24837 = ~n24099 & ~n24107;
  assign n24838 = ~n24099 & n56197;
  assign n24839 = ~n56197 & ~n24107;
  assign n24840 = n24099 & ~n56197;
  assign n24841 = ~n56350 & ~n56351;
  assign n24842 = ~n24107 & ~n24836;
  assign n24843 = ~n24835 & ~n56352;
  assign n24844 = n24090 & n56194;
  assign n24845 = ~n24098 & ~n24844;
  assign n24846 = n77 & n17524;
  assign n24847 = ~n54183 & n23459;
  assign n24848 = ~n54194 & n21969;
  assign n24849 = ~n54163 & n24302;
  assign n24850 = ~n24848 & ~n24849;
  assign n24851 = ~n24847 & ~n24848;
  assign n24852 = ~n24849 & n24851;
  assign n24853 = ~n24847 & n24850;
  assign n24854 = ~n77 & n56353;
  assign n24855 = ~n17524 & n56353;
  assign n24856 = ~n24854 & ~n24855;
  assign n24857 = ~n24846 & n56353;
  assign n24858 = pi5  & ~n56354;
  assign n24859 = ~pi5  & n56354;
  assign n24860 = ~n24858 & ~n24859;
  assign n24861 = n24845 & ~n24860;
  assign n24862 = n24086 & ~n24088;
  assign n24863 = ~n24089 & ~n24862;
  assign n24864 = n77 & n17544;
  assign n24865 = ~n54212 & n21969;
  assign n24866 = ~n54183 & n24302;
  assign n24867 = ~n54194 & n23459;
  assign n24868 = ~n24866 & ~n24867;
  assign n24869 = ~n24865 & ~n24867;
  assign n24870 = ~n24866 & n24869;
  assign n24871 = ~n24865 & n24868;
  assign n24872 = ~n77 & n56355;
  assign n24873 = ~n17544 & n56355;
  assign n24874 = ~n24872 & ~n24873;
  assign n24875 = ~n24864 & n56355;
  assign n24876 = pi5  & ~n56356;
  assign n24877 = ~pi5  & n56356;
  assign n24878 = ~n24876 & ~n24877;
  assign n24879 = n24863 & ~n24878;
  assign n24880 = n24077 & n56191;
  assign n24881 = ~n24085 & ~n24880;
  assign n24882 = n77 & n17041;
  assign n24883 = ~n54212 & n23459;
  assign n24884 = ~n54194 & n24302;
  assign n24885 = ~n54240 & n21969;
  assign n24886 = ~n24884 & ~n24885;
  assign n24887 = ~n24883 & ~n24885;
  assign n24888 = ~n24884 & n24887;
  assign n24889 = ~n24883 & n24886;
  assign n24890 = ~n77 & n56357;
  assign n24891 = ~n17041 & n56357;
  assign n24892 = ~n24890 & ~n24891;
  assign n24893 = ~n24882 & n56357;
  assign n24894 = pi5  & ~n56358;
  assign n24895 = ~pi5  & n56358;
  assign n24896 = ~n24894 & ~n24895;
  assign n24897 = n24881 & ~n24896;
  assign n24898 = n77 & n17660;
  assign n24899 = ~n54254 & n21969;
  assign n24900 = ~n54212 & n24302;
  assign n24901 = ~n54240 & n23459;
  assign n24902 = ~n24900 & ~n24901;
  assign n24903 = ~n24899 & ~n24901;
  assign n24904 = ~n24900 & n24903;
  assign n24905 = ~n24899 & n24902;
  assign n24906 = ~n24898 & n56359;
  assign n24907 = pi5  & ~n24906;
  assign n24908 = ~n24906 & ~n24907;
  assign n24909 = ~pi5  & ~n24906;
  assign n24910 = pi5  & ~n24907;
  assign n24911 = pi5  & n24906;
  assign n24912 = ~n56360 & ~n56361;
  assign n24913 = n24073 & ~n24075;
  assign n24914 = ~n24076 & ~n24913;
  assign n24915 = ~n24912 & n24914;
  assign n24916 = n77 & n17804;
  assign n24917 = ~n54254 & n23459;
  assign n24918 = ~n54240 & n24302;
  assign n24919 = ~n54269 & n21969;
  assign n24920 = ~n24918 & ~n24919;
  assign n24921 = ~n24917 & ~n24919;
  assign n24922 = ~n24918 & n24921;
  assign n24923 = ~n24917 & n24920;
  assign n24924 = ~n77 & n56362;
  assign n24925 = ~n17804 & n56362;
  assign n24926 = ~n24924 & ~n24925;
  assign n24927 = ~n24916 & n56362;
  assign n24928 = pi5  & ~n56363;
  assign n24929 = ~pi5  & n56363;
  assign n24930 = ~n24928 & ~n24929;
  assign n24931 = n24064 & n56188;
  assign n24932 = ~n56188 & ~n24072;
  assign n24933 = ~n24064 & ~n24072;
  assign n24934 = ~n24932 & ~n24933;
  assign n24935 = ~n24072 & ~n24931;
  assign n24936 = ~n24930 & ~n56364;
  assign n24937 = n77 & n17939;
  assign n24938 = ~n54254 & n24302;
  assign n24939 = ~n54277 & n21969;
  assign n24940 = ~n54269 & n23459;
  assign n24941 = ~n24939 & ~n24940;
  assign n24942 = ~n24938 & n24941;
  assign n24943 = ~n24937 & n24942;
  assign n24944 = pi5  & ~n24943;
  assign n24945 = ~n24943 & ~n24944;
  assign n24946 = ~pi5  & ~n24943;
  assign n24947 = pi5  & ~n24944;
  assign n24948 = pi5  & n24943;
  assign n24949 = ~n56365 & ~n56366;
  assign n24950 = pi8  & ~n56180;
  assign n24951 = ~n56181 & ~n24950;
  assign n24952 = n56181 & n24950;
  assign n24953 = ~n56180 & n24046;
  assign n24954 = ~n56182 & ~n24953;
  assign n24955 = ~n24951 & ~n24952;
  assign n24956 = ~n24949 & n56367;
  assign n24957 = n77 & n18056;
  assign n24958 = ~n54305 & n21969;
  assign n24959 = ~n54277 & n23459;
  assign n24960 = ~n54269 & n24302;
  assign n24961 = ~n24959 & ~n24960;
  assign n24962 = ~n24958 & ~n24959;
  assign n24963 = ~n24960 & n24962;
  assign n24964 = ~n24958 & n24961;
  assign n24965 = ~n77 & n56368;
  assign n24966 = ~n18056 & n56368;
  assign n24967 = ~n24965 & ~n24966;
  assign n24968 = ~n24957 & n56368;
  assign n24969 = pi5  & ~n56369;
  assign n24970 = ~pi5  & n56369;
  assign n24971 = ~n24969 & ~n24970;
  assign n24972 = pi8  & n24026;
  assign n24973 = ~n24025 & n24972;
  assign n24974 = n24025 & ~n24972;
  assign n24975 = ~n24027 & n24031;
  assign n24976 = ~n56180 & ~n24975;
  assign n24977 = ~n24973 & ~n24974;
  assign n24978 = ~n24971 & n56370;
  assign n24979 = n77 & ~n19275;
  assign n24980 = ~n54325 & n23459;
  assign n24981 = ~n54344 & n24302;
  assign n24982 = ~n24980 & ~n24981;
  assign n24983 = ~n24979 & n24982;
  assign n24984 = n53439 & ~n54325;
  assign n24985 = pi5  & ~n24984;
  assign n24986 = pi5  & ~n24983;
  assign n24987 = pi5  & ~n24986;
  assign n24988 = ~n24983 & ~n24986;
  assign n24989 = ~n24987 & ~n24988;
  assign n24990 = n24985 & ~n24989;
  assign n24991 = n24983 & n24985;
  assign n24992 = n77 & n18156;
  assign n24993 = ~n54305 & n24302;
  assign n24994 = ~n54325 & n21969;
  assign n24995 = ~n54344 & n23459;
  assign n24996 = ~n24994 & ~n24995;
  assign n24997 = ~n24993 & n24996;
  assign n24998 = ~n77 & n24997;
  assign n24999 = ~n18156 & n24997;
  assign n25000 = ~n24998 & ~n24999;
  assign n25001 = ~n24992 & n24997;
  assign n25002 = pi5  & ~n56372;
  assign n25003 = ~pi5  & n56372;
  assign n25004 = ~n25002 & ~n25003;
  assign n25005 = n56371 & ~n25004;
  assign n25006 = n56371 & ~n56372;
  assign n25007 = n24026 & n56373;
  assign n25008 = n77 & n18336;
  assign n25009 = ~n54305 & n23459;
  assign n25010 = ~n54277 & n24302;
  assign n25011 = ~n54344 & n21969;
  assign n25012 = ~n25010 & ~n25011;
  assign n25013 = ~n25009 & ~n25011;
  assign n25014 = ~n25010 & n25013;
  assign n25015 = ~n25009 & n25012;
  assign n25016 = ~n25008 & n56374;
  assign n25017 = pi5  & ~n25016;
  assign n25018 = pi5  & ~n25017;
  assign n25019 = pi5  & n25016;
  assign n25020 = ~n25016 & ~n25017;
  assign n25021 = ~pi5  & ~n25016;
  assign n25022 = ~n56375 & ~n56376;
  assign n25023 = ~n24026 & ~n56373;
  assign n25024 = n56373 & ~n25007;
  assign n25025 = ~n24026 & n56373;
  assign n25026 = n24026 & ~n25007;
  assign n25027 = n24026 & ~n56373;
  assign n25028 = ~n56377 & ~n56378;
  assign n25029 = ~n25007 & ~n25023;
  assign n25030 = ~n25022 & ~n56379;
  assign n25031 = ~n25007 & ~n25030;
  assign n25032 = n24971 & ~n56370;
  assign n25033 = ~n24978 & ~n25032;
  assign n25034 = ~n25031 & n25033;
  assign n25035 = ~n24978 & ~n25034;
  assign n25036 = n24949 & ~n56367;
  assign n25037 = ~n24949 & ~n24956;
  assign n25038 = ~n24949 & ~n56367;
  assign n25039 = n56367 & ~n24956;
  assign n25040 = n24949 & n56367;
  assign n25041 = ~n56380 & ~n56381;
  assign n25042 = ~n24956 & ~n25036;
  assign n25043 = ~n25035 & ~n56382;
  assign n25044 = ~n24956 & ~n25043;
  assign n25045 = n24930 & n56364;
  assign n25046 = ~n24936 & ~n25045;
  assign n25047 = ~n25044 & n25046;
  assign n25048 = ~n24936 & ~n25047;
  assign n25049 = n24912 & ~n24914;
  assign n25050 = ~n24912 & ~n24915;
  assign n25051 = ~n24912 & ~n24914;
  assign n25052 = n24914 & ~n24915;
  assign n25053 = n24912 & n24914;
  assign n25054 = ~n56383 & ~n56384;
  assign n25055 = ~n24915 & ~n25049;
  assign n25056 = ~n25048 & ~n56385;
  assign n25057 = ~n24915 & ~n25056;
  assign n25058 = ~n24881 & n24896;
  assign n25059 = n24881 & ~n24897;
  assign n25060 = n24881 & n24896;
  assign n25061 = ~n24896 & ~n24897;
  assign n25062 = ~n24881 & ~n24896;
  assign n25063 = ~n56386 & ~n56387;
  assign n25064 = ~n24897 & ~n25058;
  assign n25065 = ~n25057 & ~n56388;
  assign n25066 = ~n24897 & ~n25065;
  assign n25067 = ~n24863 & n24878;
  assign n25068 = n24863 & ~n24879;
  assign n25069 = n24863 & n24878;
  assign n25070 = ~n24878 & ~n24879;
  assign n25071 = ~n24863 & ~n24878;
  assign n25072 = ~n56389 & ~n56390;
  assign n25073 = ~n24879 & ~n25067;
  assign n25074 = ~n25066 & ~n56391;
  assign n25075 = ~n24879 & ~n25074;
  assign n25076 = ~n24845 & n24860;
  assign n25077 = ~n24861 & ~n25076;
  assign n25078 = ~n25075 & n25077;
  assign n25079 = ~n24861 & ~n25078;
  assign n25080 = n24835 & n56352;
  assign n25081 = ~n24835 & ~n24843;
  assign n25082 = ~n56352 & ~n24843;
  assign n25083 = ~n25081 & ~n25082;
  assign n25084 = ~n24843 & ~n25080;
  assign n25085 = ~n25079 & ~n56392;
  assign n25086 = ~n24843 & ~n25085;
  assign n25087 = n24816 & n56347;
  assign n25088 = ~n24816 & ~n24822;
  assign n25089 = ~n24816 & n56347;
  assign n25090 = ~n56347 & ~n24822;
  assign n25091 = n24816 & ~n56347;
  assign n25092 = ~n56393 & ~n56394;
  assign n25093 = ~n24822 & ~n25087;
  assign n25094 = ~n25086 & ~n56395;
  assign n25095 = ~n24822 & ~n25094;
  assign n25096 = n24798 & ~n24800;
  assign n25097 = ~n24798 & ~n24801;
  assign n25098 = ~n24798 & ~n24800;
  assign n25099 = n24800 & ~n24801;
  assign n25100 = n24798 & n24800;
  assign n25101 = ~n56396 & ~n56397;
  assign n25102 = ~n24801 & ~n25096;
  assign n25103 = ~n25095 & ~n56398;
  assign n25104 = ~n24801 & ~n25103;
  assign n25105 = ~n24767 & n24782;
  assign n25106 = n24767 & ~n24783;
  assign n25107 = n24767 & n24782;
  assign n25108 = ~n24782 & ~n24783;
  assign n25109 = ~n24767 & ~n24782;
  assign n25110 = ~n56399 & ~n56400;
  assign n25111 = ~n24783 & ~n25105;
  assign n25112 = ~n25104 & ~n56401;
  assign n25113 = ~n24783 & ~n25112;
  assign n25114 = ~n24747 & n24764;
  assign n25115 = n24747 & ~n24765;
  assign n25116 = n24747 & n24764;
  assign n25117 = ~n24764 & ~n24765;
  assign n25118 = ~n24747 & ~n24764;
  assign n25119 = ~n56402 & ~n56403;
  assign n25120 = ~n24765 & ~n25114;
  assign n25121 = ~n25113 & ~n56404;
  assign n25122 = ~n24765 & ~n25121;
  assign n25123 = ~n24729 & n24744;
  assign n25124 = ~n24745 & ~n25123;
  assign n25125 = ~n25122 & n25124;
  assign n25126 = ~n24745 & ~n25125;
  assign n25127 = n24721 & n56334;
  assign n25128 = ~n24721 & ~n24727;
  assign n25129 = ~n24721 & n56334;
  assign n25130 = ~n56334 & ~n24727;
  assign n25131 = n24721 & ~n56334;
  assign n25132 = ~n56405 & ~n56406;
  assign n25133 = ~n24727 & ~n25127;
  assign n25134 = ~n25126 & ~n56407;
  assign n25135 = ~n24727 & ~n25134;
  assign n25136 = n24698 & n56330;
  assign n25137 = ~n24698 & ~n24706;
  assign n25138 = ~n56330 & ~n24706;
  assign n25139 = ~n25137 & ~n25138;
  assign n25140 = ~n24706 & ~n25136;
  assign n25141 = ~n25135 & ~n56408;
  assign n25142 = ~n24706 & ~n25141;
  assign n25143 = n24680 & ~n24682;
  assign n25144 = ~n24680 & ~n24683;
  assign n25145 = ~n24680 & ~n24682;
  assign n25146 = n24682 & ~n24683;
  assign n25147 = n24680 & n24682;
  assign n25148 = ~n56409 & ~n56410;
  assign n25149 = ~n24683 & ~n25143;
  assign n25150 = ~n25142 & ~n56411;
  assign n25151 = ~n24683 & ~n25150;
  assign n25152 = ~n24649 & n24664;
  assign n25153 = n24649 & ~n24665;
  assign n25154 = n24649 & n24664;
  assign n25155 = ~n24664 & ~n24665;
  assign n25156 = ~n24649 & ~n24664;
  assign n25157 = ~n56412 & ~n56413;
  assign n25158 = ~n24665 & ~n25152;
  assign n25159 = ~n25151 & ~n56414;
  assign n25160 = ~n24665 & ~n25159;
  assign n25161 = ~n24631 & n24646;
  assign n25162 = n24631 & ~n24647;
  assign n25163 = n24631 & n24646;
  assign n25164 = ~n24646 & ~n24647;
  assign n25165 = ~n24631 & ~n24646;
  assign n25166 = ~n56415 & ~n56416;
  assign n25167 = ~n24647 & ~n25161;
  assign n25168 = ~n25160 & ~n56417;
  assign n25169 = ~n24647 & ~n25168;
  assign n25170 = ~n24613 & n24628;
  assign n25171 = ~n24629 & ~n25170;
  assign n25172 = ~n25169 & n25171;
  assign n25173 = ~n24629 & ~n25172;
  assign n25174 = n24603 & n56315;
  assign n25175 = ~n24603 & ~n24611;
  assign n25176 = ~n56315 & ~n24611;
  assign n25177 = ~n25175 & ~n25176;
  assign n25178 = ~n24611 & ~n25174;
  assign n25179 = ~n25173 & ~n56418;
  assign n25180 = ~n24611 & ~n25179;
  assign n25181 = n24582 & n56309;
  assign n25182 = ~n24582 & ~n24588;
  assign n25183 = ~n24582 & n56309;
  assign n25184 = ~n56309 & ~n24588;
  assign n25185 = n24582 & ~n56309;
  assign n25186 = ~n56419 & ~n56420;
  assign n25187 = ~n24588 & ~n25181;
  assign n25188 = ~n25180 & ~n56421;
  assign n25189 = ~n24588 & ~n25188;
  assign n25190 = n24564 & ~n24566;
  assign n25191 = ~n24564 & ~n24567;
  assign n25192 = ~n24564 & ~n24566;
  assign n25193 = n24566 & ~n24567;
  assign n25194 = n24564 & n24566;
  assign n25195 = ~n56422 & ~n56423;
  assign n25196 = ~n24567 & ~n25190;
  assign n25197 = ~n25189 & ~n56424;
  assign n25198 = ~n24567 & ~n25197;
  assign n25199 = ~n24533 & n24548;
  assign n25200 = n24533 & ~n24549;
  assign n25201 = n24533 & n24548;
  assign n25202 = ~n24548 & ~n24549;
  assign n25203 = ~n24533 & ~n24548;
  assign n25204 = ~n56425 & ~n56426;
  assign n25205 = ~n24549 & ~n25199;
  assign n25206 = ~n25198 & ~n56427;
  assign n25207 = ~n24549 & ~n25206;
  assign n25208 = ~n24515 & n24530;
  assign n25209 = ~n24531 & ~n25208;
  assign n25210 = ~n25207 & n25209;
  assign n25211 = ~n24531 & ~n25210;
  assign n25212 = n24507 & n56298;
  assign n25213 = ~n24507 & ~n24513;
  assign n25214 = ~n24507 & n56298;
  assign n25215 = ~n56298 & ~n24513;
  assign n25216 = n24507 & ~n56298;
  assign n25217 = ~n56428 & ~n56429;
  assign n25218 = ~n24513 & ~n25212;
  assign n25219 = ~n25211 & ~n56430;
  assign n25220 = ~n24513 & ~n25219;
  assign n25221 = n24484 & n56294;
  assign n25222 = ~n24484 & ~n24492;
  assign n25223 = ~n56294 & ~n24492;
  assign n25224 = ~n25222 & ~n25223;
  assign n25225 = ~n24492 & ~n25221;
  assign n25226 = ~n25220 & ~n56431;
  assign n25227 = ~n24492 & ~n25226;
  assign n25228 = n24461 & n56288;
  assign n25229 = ~n24461 & ~n24469;
  assign n25230 = ~n56288 & ~n24469;
  assign n25231 = ~n25229 & ~n25230;
  assign n25232 = ~n24469 & ~n25228;
  assign n25233 = ~n25227 & ~n56432;
  assign n25234 = ~n24469 & ~n25233;
  assign n25235 = n24440 & n56282;
  assign n25236 = ~n24440 & ~n24446;
  assign n25237 = ~n24440 & n56282;
  assign n25238 = ~n56282 & ~n24446;
  assign n25239 = n24440 & ~n56282;
  assign n25240 = ~n56433 & ~n56434;
  assign n25241 = ~n24446 & ~n25235;
  assign n25242 = ~n25234 & ~n56435;
  assign n25243 = ~n24446 & ~n25242;
  assign n25244 = n24419 & n56278;
  assign n25245 = ~n24419 & ~n24425;
  assign n25246 = ~n24419 & n56278;
  assign n25247 = ~n56278 & ~n24425;
  assign n25248 = n24419 & ~n56278;
  assign n25249 = ~n56436 & ~n56437;
  assign n25250 = ~n24425 & ~n25244;
  assign n25251 = ~n25243 & ~n56438;
  assign n25252 = ~n24425 & ~n25251;
  assign n25253 = n24396 & n56274;
  assign n25254 = ~n24396 & ~n24404;
  assign n25255 = ~n56274 & ~n24404;
  assign n25256 = ~n25254 & ~n25255;
  assign n25257 = ~n24404 & ~n25253;
  assign n25258 = ~n25252 & ~n56439;
  assign n25259 = ~n24404 & ~n25258;
  assign n25260 = n56267 & n56268;
  assign n25261 = ~n56268 & ~n24380;
  assign n25262 = ~n56267 & ~n24380;
  assign n25263 = ~n25261 & ~n25262;
  assign n25264 = ~n24380 & ~n25260;
  assign n25265 = ~n25259 & ~n56440;
  assign n25266 = n25259 & n56440;
  assign n25267 = ~n25265 & ~n25266;
  assign n25268 = n25252 & n56439;
  assign n25269 = ~n25258 & ~n25268;
  assign n25270 = n54351 & n24338;
  assign n25271 = ~n53634 & n24337;
  assign n25272 = ~pi0  & pi1 ;
  assign n25273 = ~n2325 & n25272;
  assign n25274 = ~n25271 & ~n25273;
  assign n25275 = ~n24338 & n25274;
  assign n25276 = ~n54351 & n25274;
  assign n25277 = ~n25275 & ~n25276;
  assign n25278 = ~n25270 & n25274;
  assign n25279 = pi2  & ~n56441;
  assign n25280 = ~pi2  & n56441;
  assign n25281 = ~n25279 & ~n25280;
  assign n25282 = n25269 & ~n25281;
  assign n25283 = n25243 & n56438;
  assign n25284 = ~n25251 & ~n25283;
  assign n25285 = n11242 & n24338;
  assign n25286 = ~n53650 & n24337;
  assign n25287 = pi0  & ~n56258;
  assign n25288 = ~n2325 & n25287;
  assign n25289 = ~n53634 & n25272;
  assign n25290 = ~n25288 & ~n25289;
  assign n25291 = ~n25286 & ~n25289;
  assign n25292 = ~n25288 & n25291;
  assign n25293 = ~n25286 & n25290;
  assign n25294 = ~n24338 & n56442;
  assign n25295 = ~n11242 & n56442;
  assign n25296 = ~n25294 & ~n25295;
  assign n25297 = ~n25285 & n56442;
  assign n25298 = pi2  & ~n56443;
  assign n25299 = ~pi2  & n56443;
  assign n25300 = ~n25298 & ~n25299;
  assign n25301 = n25284 & ~n25300;
  assign n25302 = n25234 & n56435;
  assign n25303 = ~n25242 & ~n25302;
  assign n25304 = n11286 & n24338;
  assign n25305 = ~n53650 & n25272;
  assign n25306 = ~n53657 & n24337;
  assign n25307 = ~n53634 & n25287;
  assign n25308 = ~n25306 & ~n25307;
  assign n25309 = ~n25305 & ~n25306;
  assign n25310 = ~n25307 & n25309;
  assign n25311 = ~n25305 & n25308;
  assign n25312 = ~n24338 & n56444;
  assign n25313 = ~n11286 & n56444;
  assign n25314 = ~n25312 & ~n25313;
  assign n25315 = ~n25304 & n56444;
  assign n25316 = pi2  & ~n56445;
  assign n25317 = ~pi2  & n56445;
  assign n25318 = ~n25316 & ~n25317;
  assign n25319 = n25303 & ~n25318;
  assign n25320 = n25227 & n56432;
  assign n25321 = ~n25233 & ~n25320;
  assign n25322 = n11213 & n24338;
  assign n25323 = ~n53650 & n25287;
  assign n25324 = ~n53685 & n24337;
  assign n25325 = ~n53657 & n25272;
  assign n25326 = ~n25324 & ~n25325;
  assign n25327 = ~n25323 & n25326;
  assign n25328 = ~n24338 & n25327;
  assign n25329 = ~n11213 & n25327;
  assign n25330 = ~n25328 & ~n25329;
  assign n25331 = ~n25322 & n25327;
  assign n25332 = pi2  & ~n56446;
  assign n25333 = ~pi2  & n56446;
  assign n25334 = ~n25332 & ~n25333;
  assign n25335 = n25321 & ~n25334;
  assign n25336 = n25220 & n56431;
  assign n25337 = ~n25226 & ~n25336;
  assign n25338 = n11380 & n24338;
  assign n25339 = ~n53685 & n25272;
  assign n25340 = ~n53657 & n25287;
  assign n25341 = ~n53712 & n24337;
  assign n25342 = ~n25340 & ~n25341;
  assign n25343 = ~n25339 & ~n25341;
  assign n25344 = ~n25340 & n25343;
  assign n25345 = ~n25339 & n25342;
  assign n25346 = ~n24338 & n56447;
  assign n25347 = ~n11380 & n56447;
  assign n25348 = ~n25346 & ~n25347;
  assign n25349 = ~n25338 & n56447;
  assign n25350 = pi2  & ~n56448;
  assign n25351 = ~pi2  & n56448;
  assign n25352 = ~n25350 & ~n25351;
  assign n25353 = n25337 & ~n25352;
  assign n25354 = n11360 & n24338;
  assign n25355 = ~n53685 & n25287;
  assign n25356 = ~n53741 & n24337;
  assign n25357 = ~n53712 & n25272;
  assign n25358 = ~n25356 & ~n25357;
  assign n25359 = ~n25355 & ~n25356;
  assign n25360 = ~n25357 & n25359;
  assign n25361 = ~n25355 & n25358;
  assign n25362 = ~n24338 & n56449;
  assign n25363 = ~n11360 & n56449;
  assign n25364 = ~n25362 & ~n25363;
  assign n25365 = ~n25354 & n56449;
  assign n25366 = pi2  & ~n56450;
  assign n25367 = ~pi2  & n56450;
  assign n25368 = ~n25366 & ~n25367;
  assign n25369 = n25211 & n56430;
  assign n25370 = ~n25219 & ~n25369;
  assign n25371 = n25368 & ~n25370;
  assign n25372 = n25207 & ~n25209;
  assign n25373 = ~n25210 & ~n25372;
  assign n25374 = n25198 & ~n56426;
  assign n25375 = ~n56425 & n25374;
  assign n25376 = n25198 & n56427;
  assign n25377 = ~n25206 & ~n56451;
  assign n25378 = n25189 & n56424;
  assign n25379 = ~n25197 & ~n25378;
  assign n25380 = n25180 & n56421;
  assign n25381 = ~n25188 & ~n25380;
  assign n25382 = n12938 & n24338;
  assign n25383 = ~n53819 & n25287;
  assign n25384 = ~n53860 & n24337;
  assign n25385 = ~n53845 & n25272;
  assign n25386 = ~n25384 & ~n25385;
  assign n25387 = ~n25383 & ~n25384;
  assign n25388 = ~n25385 & n25387;
  assign n25389 = ~n25383 & n25386;
  assign n25390 = ~n24338 & n56452;
  assign n25391 = ~n12938 & n56452;
  assign n25392 = ~n25390 & ~n25391;
  assign n25393 = ~n25382 & n56452;
  assign n25394 = pi2  & ~n56453;
  assign n25395 = ~pi2  & n56453;
  assign n25396 = ~n25394 & ~n25395;
  assign n25397 = n25173 & n56418;
  assign n25398 = ~n25179 & ~n25397;
  assign n25399 = n25396 & ~n25398;
  assign n25400 = n25169 & ~n25171;
  assign n25401 = ~n25172 & ~n25400;
  assign n25402 = n25160 & ~n56416;
  assign n25403 = ~n56415 & n25402;
  assign n25404 = n25160 & n56417;
  assign n25405 = ~n25168 & ~n56454;
  assign n25406 = n25151 & ~n56413;
  assign n25407 = ~n56412 & n25406;
  assign n25408 = n25151 & n56414;
  assign n25409 = ~n25159 & ~n56455;
  assign n25410 = n25142 & n56411;
  assign n25411 = ~n25150 & ~n25410;
  assign n25412 = n25135 & n56408;
  assign n25413 = ~n25141 & ~n25412;
  assign n25414 = n14708 & n24338;
  assign n25415 = ~n54005 & n24337;
  assign n25416 = ~n53970 & n25272;
  assign n25417 = ~n53962 & n25287;
  assign n25418 = ~n25416 & ~n25417;
  assign n25419 = ~n25415 & ~n25416;
  assign n25420 = ~n25417 & n25419;
  assign n25421 = ~n25415 & n25418;
  assign n25422 = ~n24338 & n56456;
  assign n25423 = ~n14708 & n56456;
  assign n25424 = ~n25422 & ~n25423;
  assign n25425 = ~n25414 & n56456;
  assign n25426 = pi2  & ~n56457;
  assign n25427 = ~pi2  & n56457;
  assign n25428 = ~n25426 & ~n25427;
  assign n25429 = n25126 & n56407;
  assign n25430 = ~n25134 & ~n25429;
  assign n25431 = n25428 & ~n25430;
  assign n25432 = n25122 & ~n25124;
  assign n25433 = ~n25125 & ~n25432;
  assign n25434 = n25113 & ~n56403;
  assign n25435 = ~n56402 & n25434;
  assign n25436 = n25113 & n56404;
  assign n25437 = ~n25121 & ~n56458;
  assign n25438 = n25104 & ~n56400;
  assign n25439 = ~n56399 & n25438;
  assign n25440 = n25104 & n56401;
  assign n25441 = ~n25112 & ~n56459;
  assign n25442 = n25095 & n56398;
  assign n25443 = ~n25103 & ~n25442;
  assign n25444 = n25086 & n56395;
  assign n25445 = ~n25094 & ~n25444;
  assign n25446 = n16547 & n24338;
  assign n25447 = ~n54119 & n25272;
  assign n25448 = ~n54098 & n25287;
  assign n25449 = ~n54132 & n24337;
  assign n25450 = ~n25448 & ~n25449;
  assign n25451 = ~n25447 & ~n25449;
  assign n25452 = ~n25448 & n25451;
  assign n25453 = ~n25447 & n25450;
  assign n25454 = ~n24338 & n56460;
  assign n25455 = ~n16547 & n56460;
  assign n25456 = ~n25454 & ~n25455;
  assign n25457 = ~n25446 & n56460;
  assign n25458 = pi2  & ~n56461;
  assign n25459 = ~pi2  & n56461;
  assign n25460 = ~n25458 & ~n25459;
  assign n25461 = n25079 & n56392;
  assign n25462 = ~n25085 & ~n25461;
  assign n25463 = n25460 & ~n25462;
  assign n25464 = n25075 & ~n25077;
  assign n25465 = ~n25078 & ~n25464;
  assign n25466 = n25066 & ~n56390;
  assign n25467 = ~n56389 & n25466;
  assign n25468 = n25066 & n56391;
  assign n25469 = ~n25074 & ~n56462;
  assign n25470 = n25057 & ~n56387;
  assign n25471 = ~n56386 & n25470;
  assign n25472 = n25057 & n56388;
  assign n25473 = ~n25065 & ~n56463;
  assign n25474 = n25048 & n56385;
  assign n25475 = ~n25056 & ~n25474;
  assign n25476 = n25044 & ~n25046;
  assign n25477 = ~n25047 & ~n25476;
  assign n25478 = n17041 & n24338;
  assign n25479 = ~n54212 & n25272;
  assign n25480 = ~n54194 & n25287;
  assign n25481 = ~n54240 & n24337;
  assign n25482 = ~n25480 & ~n25481;
  assign n25483 = ~n25479 & ~n25481;
  assign n25484 = ~n25480 & n25483;
  assign n25485 = ~n25479 & n25482;
  assign n25486 = ~n24338 & n56464;
  assign n25487 = ~n17041 & n56464;
  assign n25488 = ~n25486 & ~n25487;
  assign n25489 = ~n25478 & n56464;
  assign n25490 = pi2  & ~n56465;
  assign n25491 = ~pi2  & n56465;
  assign n25492 = ~n25490 & ~n25491;
  assign n25493 = n25035 & n56382;
  assign n25494 = ~n25043 & ~n25493;
  assign n25495 = n25492 & ~n25494;
  assign n25496 = n25031 & ~n25033;
  assign n25497 = ~n25034 & ~n25496;
  assign n25498 = n17939 & n24338;
  assign n25499 = ~n54254 & n25287;
  assign n25500 = ~n54277 & n24337;
  assign n25501 = ~n54269 & n25272;
  assign n25502 = ~n25500 & ~n25501;
  assign n25503 = ~n25499 & n25502;
  assign n25504 = ~n25498 & n25503;
  assign n25505 = ~pi2  & ~n25504;
  assign n25506 = pi2  & n25504;
  assign n25507 = pi2  & ~n25504;
  assign n25508 = ~pi2  & n25504;
  assign n25509 = ~n25507 & ~n25508;
  assign n25510 = ~n25505 & ~n25506;
  assign n25511 = pi5  & ~n56371;
  assign n25512 = n56372 & ~n25511;
  assign n25513 = ~n56372 & n25511;
  assign n25514 = ~n56372 & ~n25511;
  assign n25515 = n56372 & n25511;
  assign n25516 = ~n25514 & ~n25515;
  assign n25517 = ~n56371 & n25004;
  assign n25518 = ~n56373 & ~n25517;
  assign n25519 = ~n25512 & ~n25513;
  assign n25520 = n56466 & n56467;
  assign n25521 = n18056 & n24338;
  assign n25522 = ~n54305 & n24337;
  assign n25523 = ~n54269 & n25287;
  assign n25524 = ~n54277 & n25272;
  assign n25525 = ~n25523 & ~n25524;
  assign n25526 = ~n25522 & ~n25524;
  assign n25527 = ~n25523 & n25526;
  assign n25528 = ~n25522 & n25525;
  assign n25529 = ~n24338 & n56468;
  assign n25530 = ~n18056 & n56468;
  assign n25531 = ~n25529 & ~n25530;
  assign n25532 = ~n25521 & n56468;
  assign n25533 = pi2  & ~n56469;
  assign n25534 = ~pi2  & n56469;
  assign n25535 = ~n25533 & ~n25534;
  assign n25536 = n18336 & n24338;
  assign n25537 = ~n54305 & n25272;
  assign n25538 = ~n54277 & n25287;
  assign n25539 = ~n54344 & n24337;
  assign n25540 = ~n25538 & ~n25539;
  assign n25541 = ~n25537 & ~n25539;
  assign n25542 = ~n25538 & n25541;
  assign n25543 = ~n25537 & n25540;
  assign n25544 = ~n25536 & n56470;
  assign n25545 = n24984 & n25544;
  assign n25546 = pi0  & ~n54305;
  assign n25547 = n54344 & ~n25546;
  assign n25548 = ~n24330 & ~n25547;
  assign n25549 = n54325 & ~n25548;
  assign n25550 = pi2  & ~n25549;
  assign n25551 = ~n25545 & n25550;
  assign n25552 = ~pi2  & n25544;
  assign n25553 = ~n24984 & ~n25544;
  assign n25554 = pi2  & n25544;
  assign n25555 = n24984 & ~n25544;
  assign n25556 = ~n25554 & ~n25555;
  assign n25557 = ~n25552 & ~n25553;
  assign n25558 = pi2  & n24338;
  assign n25559 = n18156 & n25558;
  assign n25560 = ~n54305 & n25287;
  assign n25561 = ~n54325 & n24337;
  assign n25562 = ~n54344 & n25272;
  assign n25563 = ~n25561 & ~n25562;
  assign n25564 = ~n25560 & n25563;
  assign n25565 = pi2  & ~n25564;
  assign n25566 = ~n19275 & n25558;
  assign n25567 = pi0  & ~n54325;
  assign n25568 = pi2  & ~n25567;
  assign n25569 = pi2  & n25272;
  assign n25570 = ~n54325 & n25569;
  assign n25571 = pi2  & n25287;
  assign n25572 = ~n54344 & n25571;
  assign n25573 = ~n25570 & ~n25572;
  assign n25574 = ~pi0  & ~n25569;
  assign n25575 = ~n54325 & ~n25574;
  assign n25576 = ~n54344 & n25287;
  assign n25577 = pi2  & ~n25572;
  assign n25578 = pi2  & ~n25576;
  assign n25579 = ~n25575 & n56472;
  assign n25580 = n25568 & n25573;
  assign n25581 = ~n25566 & n56473;
  assign n25582 = ~n25565 & n25581;
  assign n25583 = ~n25570 & n56472;
  assign n25584 = ~n25566 & n25583;
  assign n25585 = ~n25565 & n25584;
  assign n25586 = ~n25559 & n25585;
  assign n25587 = ~n25567 & n25586;
  assign n25588 = n18153 & ~n19274;
  assign n25589 = n25558 & ~n25588;
  assign n25590 = ~n25565 & n56473;
  assign n25591 = ~n25589 & n25590;
  assign n25592 = ~n25559 & n25582;
  assign n25593 = ~n24984 & ~n56474;
  assign n25594 = ~pi2  & ~n25544;
  assign n25595 = pi2  & ~n25544;
  assign n25596 = ~n25552 & ~n25595;
  assign n25597 = ~n25554 & ~n25594;
  assign n25598 = ~n25593 & n56475;
  assign n25599 = ~n25551 & ~n56471;
  assign n25600 = ~n25535 & n56476;
  assign n25601 = n25535 & ~n56476;
  assign n25602 = pi5  & n24984;
  assign n25603 = n24983 & ~n25602;
  assign n25604 = ~n24983 & n25602;
  assign n25605 = ~n24985 & n24989;
  assign n25606 = ~n56371 & ~n25605;
  assign n25607 = ~n25603 & ~n25604;
  assign n25608 = ~n25601 & n56477;
  assign n25609 = ~n25600 & ~n25608;
  assign n25610 = ~n25520 & n25609;
  assign n25611 = ~n56466 & ~n56467;
  assign n25612 = ~n56467 & n25609;
  assign n25613 = n56467 & ~n25609;
  assign n25614 = ~n56466 & ~n25613;
  assign n25615 = ~n25612 & ~n25614;
  assign n25616 = n56466 & ~n25612;
  assign n25617 = ~n25613 & ~n25616;
  assign n25618 = ~n25610 & ~n25611;
  assign n25619 = n25022 & n56379;
  assign n25620 = ~n25030 & ~n25619;
  assign n25621 = n17804 & n24338;
  assign n25622 = ~n54254 & n25272;
  assign n25623 = ~n54240 & n25287;
  assign n25624 = ~n54269 & n24337;
  assign n25625 = ~n25623 & ~n25624;
  assign n25626 = ~n25622 & ~n25624;
  assign n25627 = ~n25623 & n25626;
  assign n25628 = ~n25622 & n25625;
  assign n25629 = ~n24338 & n56479;
  assign n25630 = ~n17804 & n56479;
  assign n25631 = ~n25629 & ~n25630;
  assign n25632 = ~n25621 & n56479;
  assign n25633 = pi2  & ~n56480;
  assign n25634 = ~pi2  & n56480;
  assign n25635 = ~n25633 & ~n25634;
  assign n25636 = n25620 & ~n25635;
  assign n25637 = ~n56478 & ~n25636;
  assign n25638 = ~n25620 & n25635;
  assign n25639 = n56478 & n25620;
  assign n25640 = n25635 & ~n25639;
  assign n25641 = ~n56478 & ~n25620;
  assign n25642 = ~n25640 & ~n25641;
  assign n25643 = n56478 & ~n25635;
  assign n25644 = ~n56478 & n25635;
  assign n25645 = n25620 & ~n25644;
  assign n25646 = ~n25643 & ~n25645;
  assign n25647 = ~n25637 & ~n25638;
  assign n25648 = ~n25497 & ~n56481;
  assign n25649 = n17660 & n24338;
  assign n25650 = ~n54254 & n24337;
  assign n25651 = ~n54212 & n25287;
  assign n25652 = ~n54240 & n25272;
  assign n25653 = ~n25651 & ~n25652;
  assign n25654 = ~n25650 & ~n25652;
  assign n25655 = ~n25651 & n25654;
  assign n25656 = ~n25650 & n25653;
  assign n25657 = ~n25649 & n56482;
  assign n25658 = pi2  & ~n25657;
  assign n25659 = ~pi2  & n25657;
  assign n25660 = ~pi2  & ~n25657;
  assign n25661 = pi2  & n25657;
  assign n25662 = ~n25660 & ~n25661;
  assign n25663 = ~n25658 & ~n25659;
  assign n25664 = ~n25648 & ~n56483;
  assign n25665 = n25497 & n56481;
  assign n25666 = ~n25492 & n25494;
  assign n25667 = ~n25665 & ~n25666;
  assign n25668 = ~n25664 & n25667;
  assign n25669 = ~n25664 & ~n25665;
  assign n25670 = n25492 & n25669;
  assign n25671 = n25494 & ~n25670;
  assign n25672 = ~n25492 & ~n25669;
  assign n25673 = ~n25671 & ~n25672;
  assign n25674 = ~n25495 & ~n25668;
  assign n25675 = ~n25477 & n56484;
  assign n25676 = n25477 & ~n56484;
  assign n25677 = n17544 & n24338;
  assign n25678 = ~n54212 & n24337;
  assign n25679 = ~n54183 & n25287;
  assign n25680 = ~n54194 & n25272;
  assign n25681 = ~n25679 & ~n25680;
  assign n25682 = ~n25678 & ~n25680;
  assign n25683 = ~n25679 & n25682;
  assign n25684 = ~n25678 & n25681;
  assign n25685 = ~n24338 & n56485;
  assign n25686 = ~n17544 & n56485;
  assign n25687 = ~n25685 & ~n25686;
  assign n25688 = ~n25677 & n56485;
  assign n25689 = ~pi2  & n56486;
  assign n25690 = pi2  & ~n56486;
  assign n25691 = ~n25689 & ~n25690;
  assign n25692 = ~n25676 & n25691;
  assign n25693 = n56484 & n25691;
  assign n25694 = n25477 & ~n25693;
  assign n25695 = ~n56484 & ~n25691;
  assign n25696 = ~n25694 & ~n25695;
  assign n25697 = ~n25675 & ~n25692;
  assign n25698 = ~n25475 & n56487;
  assign n25699 = n25475 & ~n56487;
  assign n25700 = n17524 & n24338;
  assign n25701 = ~n54183 & n25272;
  assign n25702 = ~n54194 & n24337;
  assign n25703 = ~n54163 & n25287;
  assign n25704 = ~n25702 & ~n25703;
  assign n25705 = ~n25701 & ~n25702;
  assign n25706 = ~n25703 & n25705;
  assign n25707 = ~n25701 & n25704;
  assign n25708 = ~n24338 & n56488;
  assign n25709 = ~n17524 & n56488;
  assign n25710 = ~n25708 & ~n25709;
  assign n25711 = ~n25700 & n56488;
  assign n25712 = ~pi2  & n56489;
  assign n25713 = pi2  & ~n56489;
  assign n25714 = ~n25712 & ~n25713;
  assign n25715 = ~n25699 & n25714;
  assign n25716 = n56487 & n25714;
  assign n25717 = n25475 & ~n25716;
  assign n25718 = ~n56487 & ~n25714;
  assign n25719 = ~n25717 & ~n25718;
  assign n25720 = ~n25698 & ~n25715;
  assign n25721 = n25473 & ~n56490;
  assign n25722 = ~n25473 & n56490;
  assign n25723 = n17072 & n24338;
  assign n25724 = ~n54154 & n25287;
  assign n25725 = ~n54183 & n24337;
  assign n25726 = ~n54163 & n25272;
  assign n25727 = ~n25725 & ~n25726;
  assign n25728 = ~n25724 & n25727;
  assign n25729 = ~n25723 & n25728;
  assign n25730 = pi2  & ~n25729;
  assign n25731 = ~pi2  & n25729;
  assign n25732 = ~pi2  & ~n25729;
  assign n25733 = pi2  & n25729;
  assign n25734 = ~n25732 & ~n25733;
  assign n25735 = ~n25730 & ~n25731;
  assign n25736 = ~n25722 & ~n56491;
  assign n25737 = ~n25721 & ~n25736;
  assign n25738 = n25469 & ~n25737;
  assign n25739 = ~n25469 & n25737;
  assign n25740 = n16522 & n24338;
  assign n25741 = ~n54154 & n25272;
  assign n25742 = ~n54132 & n25287;
  assign n25743 = ~n54163 & n24337;
  assign n25744 = ~n25742 & ~n25743;
  assign n25745 = ~n25741 & ~n25743;
  assign n25746 = ~n25742 & n25745;
  assign n25747 = ~n25741 & n25744;
  assign n25748 = ~n25740 & n56492;
  assign n25749 = pi2  & ~n25748;
  assign n25750 = ~pi2  & n25748;
  assign n25751 = ~pi2  & ~n25748;
  assign n25752 = pi2  & n25748;
  assign n25753 = ~n25751 & ~n25752;
  assign n25754 = ~n25749 & ~n25750;
  assign n25755 = ~n25739 & ~n56493;
  assign n25756 = ~n25738 & ~n25755;
  assign n25757 = ~n25465 & n25756;
  assign n25758 = n16772 & n24338;
  assign n25759 = ~n54154 & n24337;
  assign n25760 = ~n54119 & n25287;
  assign n25761 = ~n54132 & n25272;
  assign n25762 = ~n25760 & ~n25761;
  assign n25763 = ~n25759 & ~n25761;
  assign n25764 = ~n25760 & n25763;
  assign n25765 = ~n25759 & n25762;
  assign n25766 = ~n25758 & n56494;
  assign n25767 = pi2  & ~n25766;
  assign n25768 = ~pi2  & n25766;
  assign n25769 = ~pi2  & ~n25766;
  assign n25770 = pi2  & n25766;
  assign n25771 = ~n25769 & ~n25770;
  assign n25772 = ~n25767 & ~n25768;
  assign n25773 = ~n25757 & ~n56495;
  assign n25774 = n25465 & ~n25756;
  assign n25775 = ~n25460 & n25462;
  assign n25776 = ~n25774 & ~n25775;
  assign n25777 = ~n25773 & n25776;
  assign n25778 = ~n25773 & ~n25774;
  assign n25779 = n25460 & n25778;
  assign n25780 = n25462 & ~n25779;
  assign n25781 = ~n25460 & ~n25778;
  assign n25782 = ~n25780 & ~n25781;
  assign n25783 = ~n25463 & ~n25777;
  assign n25784 = ~n25445 & n56496;
  assign n25785 = n25445 & ~n56496;
  assign n25786 = n15779 & n24338;
  assign n25787 = ~n54098 & n25272;
  assign n25788 = ~n54119 & n24337;
  assign n25789 = ~n54073 & n25287;
  assign n25790 = ~n25788 & ~n25789;
  assign n25791 = ~n25787 & ~n25788;
  assign n25792 = ~n25789 & n25791;
  assign n25793 = ~n25787 & ~n25789;
  assign n25794 = ~n25788 & n25793;
  assign n25795 = ~n25787 & n25790;
  assign n25796 = ~n24338 & n56497;
  assign n25797 = ~n15779 & n56497;
  assign n25798 = ~n25796 & ~n25797;
  assign n25799 = ~n25786 & n56497;
  assign n25800 = ~pi2  & n56498;
  assign n25801 = pi2  & ~n56498;
  assign n25802 = ~n25800 & ~n25801;
  assign n25803 = ~n25785 & n25802;
  assign n25804 = n56496 & n25802;
  assign n25805 = n25445 & ~n25804;
  assign n25806 = ~n56496 & ~n25802;
  assign n25807 = ~n25805 & ~n25806;
  assign n25808 = ~n25784 & ~n25803;
  assign n25809 = ~n25443 & n56499;
  assign n25810 = n25443 & ~n56499;
  assign n25811 = n16138 & n24338;
  assign n25812 = ~n54098 & n24337;
  assign n25813 = ~n54050 & n25287;
  assign n25814 = ~n54073 & n25272;
  assign n25815 = ~n25813 & ~n25814;
  assign n25816 = ~n25812 & ~n25814;
  assign n25817 = ~n25813 & n25816;
  assign n25818 = ~n25812 & n25815;
  assign n25819 = ~n24338 & n56500;
  assign n25820 = ~n16138 & n56500;
  assign n25821 = ~n25819 & ~n25820;
  assign n25822 = ~n25811 & n56500;
  assign n25823 = ~pi2  & n56501;
  assign n25824 = pi2  & ~n56501;
  assign n25825 = ~n25823 & ~n25824;
  assign n25826 = ~n25810 & n25825;
  assign n25827 = n56499 & n25825;
  assign n25828 = n25443 & ~n25827;
  assign n25829 = ~n56499 & ~n25825;
  assign n25830 = ~n25828 & ~n25829;
  assign n25831 = ~n25809 & ~n25826;
  assign n25832 = n25441 & ~n56502;
  assign n25833 = ~n25441 & n56502;
  assign n25834 = n15219 & n24338;
  assign n25835 = ~n54050 & n25272;
  assign n25836 = ~n54034 & n25287;
  assign n25837 = ~n54073 & n24337;
  assign n25838 = ~n25836 & ~n25837;
  assign n25839 = ~n25835 & ~n25837;
  assign n25840 = ~n25836 & n25839;
  assign n25841 = ~n25835 & n25838;
  assign n25842 = ~n25834 & n56503;
  assign n25843 = pi2  & ~n25842;
  assign n25844 = ~pi2  & n25842;
  assign n25845 = ~pi2  & ~n25842;
  assign n25846 = pi2  & n25842;
  assign n25847 = ~n25845 & ~n25846;
  assign n25848 = ~n25843 & ~n25844;
  assign n25849 = ~n25833 & ~n56504;
  assign n25850 = ~n25832 & ~n25849;
  assign n25851 = n25437 & ~n25850;
  assign n25852 = ~n25437 & n25850;
  assign n25853 = n15195 & n24338;
  assign n25854 = ~n54050 & n24337;
  assign n25855 = ~n54005 & n25287;
  assign n25856 = ~n54034 & n25272;
  assign n25857 = ~n25855 & ~n25856;
  assign n25858 = ~n25854 & ~n25856;
  assign n25859 = ~n25855 & n25858;
  assign n25860 = ~n25854 & n25857;
  assign n25861 = ~n25853 & n56505;
  assign n25862 = pi2  & ~n25861;
  assign n25863 = ~pi2  & n25861;
  assign n25864 = ~pi2  & ~n25861;
  assign n25865 = pi2  & n25861;
  assign n25866 = ~n25864 & ~n25865;
  assign n25867 = ~n25862 & ~n25863;
  assign n25868 = ~n25852 & ~n56506;
  assign n25869 = ~n25851 & ~n25868;
  assign n25870 = ~n25433 & n25869;
  assign n25871 = n14688 & n24338;
  assign n25872 = ~n54005 & n25272;
  assign n25873 = ~n54034 & n24337;
  assign n25874 = ~n53970 & n25287;
  assign n25875 = ~n25873 & ~n25874;
  assign n25876 = ~n25872 & ~n25873;
  assign n25877 = ~n25874 & n25876;
  assign n25878 = ~n25872 & n25875;
  assign n25879 = ~n25871 & n56507;
  assign n25880 = pi2  & ~n25879;
  assign n25881 = ~pi2  & n25879;
  assign n25882 = ~pi2  & ~n25879;
  assign n25883 = pi2  & n25879;
  assign n25884 = ~n25882 & ~n25883;
  assign n25885 = ~n25880 & ~n25881;
  assign n25886 = ~n25870 & ~n56508;
  assign n25887 = n25433 & ~n25869;
  assign n25888 = ~n25428 & n25430;
  assign n25889 = ~n25887 & ~n25888;
  assign n25890 = ~n25886 & n25889;
  assign n25891 = ~n25886 & ~n25887;
  assign n25892 = n25428 & n25891;
  assign n25893 = n25430 & ~n25892;
  assign n25894 = ~n25428 & ~n25891;
  assign n25895 = ~n25893 & ~n25894;
  assign n25896 = ~n25431 & ~n25890;
  assign n25897 = ~n25413 & n56509;
  assign n25898 = n25413 & ~n56509;
  assign n25899 = n14020 & n24338;
  assign n25900 = ~n53962 & n25272;
  assign n25901 = ~n53970 & n24337;
  assign n25902 = ~n53930 & n25287;
  assign n25903 = ~n25901 & ~n25902;
  assign n25904 = ~n25900 & ~n25901;
  assign n25905 = ~n25902 & n25904;
  assign n25906 = ~n25900 & n25903;
  assign n25907 = ~n24338 & n56510;
  assign n25908 = ~n14020 & n56510;
  assign n25909 = ~n25907 & ~n25908;
  assign n25910 = ~n25899 & n56510;
  assign n25911 = ~pi2  & n56511;
  assign n25912 = pi2  & ~n56511;
  assign n25913 = ~n25911 & ~n25912;
  assign n25914 = ~n25898 & n25913;
  assign n25915 = n56509 & n25913;
  assign n25916 = n25413 & ~n25915;
  assign n25917 = ~n56509 & ~n25913;
  assign n25918 = ~n25916 & ~n25917;
  assign n25919 = ~n25897 & ~n25914;
  assign n25920 = ~n25411 & n56512;
  assign n25921 = n25411 & ~n56512;
  assign n25922 = n14263 & n24338;
  assign n25923 = ~n53930 & n25272;
  assign n25924 = ~n53962 & n24337;
  assign n25925 = ~n53907 & n25287;
  assign n25926 = ~n25924 & ~n25925;
  assign n25927 = ~n25923 & ~n25924;
  assign n25928 = ~n25925 & n25927;
  assign n25929 = ~n25923 & n25926;
  assign n25930 = ~n24338 & n56513;
  assign n25931 = ~n14263 & n56513;
  assign n25932 = ~n25930 & ~n25931;
  assign n25933 = ~n25922 & n56513;
  assign n25934 = ~pi2  & n56514;
  assign n25935 = pi2  & ~n56514;
  assign n25936 = ~n25934 & ~n25935;
  assign n25937 = ~n25921 & n25936;
  assign n25938 = n56512 & n25936;
  assign n25939 = n25411 & ~n25938;
  assign n25940 = ~n56512 & ~n25936;
  assign n25941 = ~n25939 & ~n25940;
  assign n25942 = ~n25920 & ~n25937;
  assign n25943 = n25409 & ~n56515;
  assign n25944 = ~n25409 & n56515;
  assign n25945 = n13360 & n24338;
  assign n25946 = ~n53907 & n25272;
  assign n25947 = ~n53930 & n24337;
  assign n25948 = ~n53888 & n25287;
  assign n25949 = ~n25947 & ~n25948;
  assign n25950 = ~n25946 & ~n25947;
  assign n25951 = ~n25948 & n25950;
  assign n25952 = ~n25946 & n25949;
  assign n25953 = ~n25945 & n56516;
  assign n25954 = pi2  & ~n25953;
  assign n25955 = ~pi2  & n25953;
  assign n25956 = ~pi2  & ~n25953;
  assign n25957 = pi2  & n25953;
  assign n25958 = ~n25956 & ~n25957;
  assign n25959 = ~n25954 & ~n25955;
  assign n25960 = ~n25944 & ~n56517;
  assign n25961 = ~n25943 & ~n25960;
  assign n25962 = n25405 & ~n25961;
  assign n25963 = ~n25405 & n25961;
  assign n25964 = n13336 & n24338;
  assign n25965 = ~n53888 & n25272;
  assign n25966 = ~n53907 & n24337;
  assign n25967 = ~n53860 & n25287;
  assign n25968 = ~n25966 & ~n25967;
  assign n25969 = ~n25965 & ~n25966;
  assign n25970 = ~n25967 & n25969;
  assign n25971 = ~n25965 & n25968;
  assign n25972 = ~n25964 & n56518;
  assign n25973 = pi2  & ~n25972;
  assign n25974 = ~pi2  & n25972;
  assign n25975 = ~pi2  & ~n25972;
  assign n25976 = pi2  & n25972;
  assign n25977 = ~n25975 & ~n25976;
  assign n25978 = ~n25973 & ~n25974;
  assign n25979 = ~n25963 & ~n56519;
  assign n25980 = ~n25962 & ~n25979;
  assign n25981 = ~n25401 & n25980;
  assign n25982 = n12918 & n24338;
  assign n25983 = ~n53860 & n25272;
  assign n25984 = ~n53888 & n24337;
  assign n25985 = ~n53845 & n25287;
  assign n25986 = ~n25984 & ~n25985;
  assign n25987 = ~n25983 & ~n25984;
  assign n25988 = ~n25985 & n25987;
  assign n25989 = ~n25983 & n25986;
  assign n25990 = ~n25982 & n56520;
  assign n25991 = pi2  & ~n25990;
  assign n25992 = ~pi2  & n25990;
  assign n25993 = ~pi2  & ~n25990;
  assign n25994 = pi2  & n25990;
  assign n25995 = ~n25993 & ~n25994;
  assign n25996 = ~n25991 & ~n25992;
  assign n25997 = ~n25981 & ~n56521;
  assign n25998 = n25401 & ~n25980;
  assign n25999 = ~n25396 & n25398;
  assign n26000 = ~n25998 & ~n25999;
  assign n26001 = ~n25997 & n26000;
  assign n26002 = ~n25997 & ~n25998;
  assign n26003 = n25396 & n26002;
  assign n26004 = n25398 & ~n26003;
  assign n26005 = ~n25396 & ~n26002;
  assign n26006 = ~n26004 & ~n26005;
  assign n26007 = ~n25399 & ~n26001;
  assign n26008 = ~n25381 & n56522;
  assign n26009 = n25381 & ~n56522;
  assign n26010 = n12550 & n24338;
  assign n26011 = ~n53819 & n25272;
  assign n26012 = ~n53845 & n24337;
  assign n26013 = ~n53799 & n25287;
  assign n26014 = ~n26012 & ~n26013;
  assign n26015 = ~n26011 & ~n26012;
  assign n26016 = ~n26013 & n26015;
  assign n26017 = ~n26011 & n26014;
  assign n26018 = ~n24338 & n56523;
  assign n26019 = ~n12550 & n56523;
  assign n26020 = ~n26018 & ~n26019;
  assign n26021 = ~n26010 & n56523;
  assign n26022 = ~pi2  & n56524;
  assign n26023 = pi2  & ~n56524;
  assign n26024 = ~n26022 & ~n26023;
  assign n26025 = ~n26009 & n26024;
  assign n26026 = n56522 & n26024;
  assign n26027 = n25381 & ~n26026;
  assign n26028 = ~n56522 & ~n26024;
  assign n26029 = ~n26027 & ~n26028;
  assign n26030 = ~n26008 & ~n26025;
  assign n26031 = ~n25379 & n56525;
  assign n26032 = n25379 & ~n56525;
  assign n26033 = n12690 & n24338;
  assign n26034 = ~n53774 & n25287;
  assign n26035 = ~n53819 & n24337;
  assign n26036 = ~n53799 & n25272;
  assign n26037 = ~n26035 & ~n26036;
  assign n26038 = ~n26034 & ~n26035;
  assign n26039 = ~n26036 & n26038;
  assign n26040 = ~n26034 & n26037;
  assign n26041 = ~n24338 & n56526;
  assign n26042 = ~n12690 & n56526;
  assign n26043 = ~n26041 & ~n26042;
  assign n26044 = ~n26033 & n56526;
  assign n26045 = ~pi2  & n56527;
  assign n26046 = pi2  & ~n56527;
  assign n26047 = ~n26045 & ~n26046;
  assign n26048 = ~n26032 & n26047;
  assign n26049 = n56525 & n26047;
  assign n26050 = n25379 & ~n26049;
  assign n26051 = ~n56525 & ~n26047;
  assign n26052 = ~n26050 & ~n26051;
  assign n26053 = ~n26031 & ~n26048;
  assign n26054 = n25377 & ~n56528;
  assign n26055 = ~n25377 & n56528;
  assign n26056 = n11913 & n24338;
  assign n26057 = ~n53774 & n25272;
  assign n26058 = ~n53799 & n24337;
  assign n26059 = ~n53741 & n25287;
  assign n26060 = ~n26058 & ~n26059;
  assign n26061 = ~n26057 & ~n26058;
  assign n26062 = ~n26059 & n26061;
  assign n26063 = ~n26057 & n26060;
  assign n26064 = ~n26056 & n56529;
  assign n26065 = pi2  & ~n26064;
  assign n26066 = ~pi2  & n26064;
  assign n26067 = ~pi2  & ~n26064;
  assign n26068 = pi2  & n26064;
  assign n26069 = ~n26067 & ~n26068;
  assign n26070 = ~n26065 & ~n26066;
  assign n26071 = ~n26055 & ~n56530;
  assign n26072 = ~n26054 & ~n26071;
  assign n26073 = ~n25373 & n26072;
  assign n26074 = n11889 & n24338;
  assign n26075 = ~n53712 & n25287;
  assign n26076 = ~n53774 & n24337;
  assign n26077 = ~n53741 & n25272;
  assign n26078 = ~n26076 & ~n26077;
  assign n26079 = ~n26075 & ~n26076;
  assign n26080 = ~n26077 & n26079;
  assign n26081 = ~n26075 & n26078;
  assign n26082 = ~n26074 & n56531;
  assign n26083 = pi2  & ~n26082;
  assign n26084 = ~pi2  & n26082;
  assign n26085 = ~pi2  & ~n26082;
  assign n26086 = pi2  & n26082;
  assign n26087 = ~n26085 & ~n26086;
  assign n26088 = ~n26083 & ~n26084;
  assign n26089 = ~n26073 & ~n56532;
  assign n26090 = n25373 & ~n26072;
  assign n26091 = ~n25368 & n25370;
  assign n26092 = ~n26090 & ~n26091;
  assign n26093 = ~n26089 & n26092;
  assign n26094 = ~n26089 & ~n26090;
  assign n26095 = n25368 & n26094;
  assign n26096 = n25370 & ~n26095;
  assign n26097 = ~n25368 & ~n26094;
  assign n26098 = ~n26096 & ~n26097;
  assign n26099 = ~n25371 & ~n26093;
  assign n26100 = ~n25337 & n25352;
  assign n26101 = n25337 & ~n25353;
  assign n26102 = n25337 & n25352;
  assign n26103 = ~n25352 & ~n25353;
  assign n26104 = ~n25337 & ~n25352;
  assign n26105 = ~n56534 & ~n56535;
  assign n26106 = ~n25353 & ~n26100;
  assign n26107 = ~n56533 & ~n56536;
  assign n26108 = ~n25353 & ~n26107;
  assign n26109 = ~n25321 & n25334;
  assign n26110 = ~n25335 & ~n26109;
  assign n26111 = ~n26108 & n26110;
  assign n26112 = ~n25335 & ~n26111;
  assign n26113 = ~n25303 & n25318;
  assign n26114 = ~n25319 & ~n26113;
  assign n26115 = ~n26112 & n26114;
  assign n26116 = ~n25319 & ~n26115;
  assign n26117 = ~n25284 & n25300;
  assign n26118 = ~n25301 & ~n26117;
  assign n26119 = ~n26116 & n26118;
  assign n26120 = ~n25301 & ~n26119;
  assign n26121 = ~n25269 & n25281;
  assign n26122 = ~n25282 & ~n26121;
  assign n26123 = ~n26120 & n26122;
  assign n26124 = ~n25282 & ~n26123;
  assign n26125 = n25267 & ~n26124;
  assign n26126 = ~n25265 & ~n26125;
  assign n26127 = ~n24329 & n56269;
  assign n26128 = ~n24383 & ~n26127;
  assign n26129 = ~n26126 & n26128;
  assign n26130 = ~n24383 & ~n26129;
  assign n26131 = n24322 & ~n24324;
  assign n26132 = ~n24325 & ~n26131;
  assign n26133 = ~n26130 & n26132;
  assign n26134 = ~n24325 & ~n26133;
  assign n26135 = n23486 & ~n26134;
  assign n26136 = ~n23484 & ~n26135;
  assign n26137 = ~n21961 & n55948;
  assign n26138 = ~n22686 & ~n26137;
  assign n26139 = ~n26136 & n26138;
  assign n26140 = ~n22686 & ~n26139;
  assign n26141 = n21952 & ~n21954;
  assign n26142 = ~n21955 & ~n26141;
  assign n26143 = ~n26140 & n26142;
  assign n26144 = ~n21955 & ~n26143;
  assign n26145 = n21266 & ~n26144;
  assign n26146 = ~n21264 & ~n26145;
  assign n26147 = n20652 & ~n26146;
  assign n26148 = ~n20650 & ~n26147;
  assign n26149 = ~n19538 & n55467;
  assign n26150 = ~n20055 & ~n26149;
  assign n26151 = ~n26148 & n26150;
  assign n26152 = ~n20055 & ~n26151;
  assign n26153 = n19536 & ~n26152;
  assign n26154 = ~n19534 & ~n26153;
  assign n26155 = ~n18821 & n55292;
  assign n26156 = ~n19077 & ~n26155;
  assign n26157 = ~n26154 & n26156;
  assign n26158 = ~n19077 & ~n26157;
  assign n26159 = n18812 & ~n18814;
  assign n26160 = ~n18815 & ~n26159;
  assign n26161 = ~n26158 & n26160;
  assign n26162 = ~n18815 & ~n26161;
  assign n26163 = n18585 & ~n26162;
  assign n26164 = ~n18583 & ~n26163;
  assign n26165 = n17455 & ~n26164;
  assign n26166 = ~n17453 & ~n26165;
  assign n26167 = n17240 & ~n26166;
  assign n26168 = ~n17238 & ~n26167;
  assign n26169 = n16693 & ~n26168;
  assign n26170 = ~n16691 & ~n26169;
  assign n26171 = ~n16066 & n54922;
  assign n26172 = ~n16283 & ~n26171;
  assign n26173 = ~n26170 & n26172;
  assign n26174 = ~n16283 & ~n26173;
  assign n26175 = n16064 & ~n26174;
  assign n26176 = ~n16062 & ~n26175;
  assign n26177 = n15918 & ~n26176;
  assign n26178 = ~n15916 & ~n26177;
  assign n26179 = n14816 & ~n26178;
  assign n26180 = ~n14814 & ~n26179;
  assign n26181 = ~n14233 & n54714;
  assign n26182 = ~n14383 & ~n26181;
  assign n26183 = ~n26180 & n26182;
  assign n26184 = ~n14383 & ~n26183;
  assign n26185 = n14231 & ~n26184;
  assign n26186 = ~n14229 & ~n26185;
  assign n26187 = ~n13115 & n54671;
  assign n26188 = ~n14136 & ~n26187;
  assign n26189 = ~n26186 & n26188;
  assign n26190 = ~n14136 & ~n26189;
  assign n26191 = n13104 & ~n13108;
  assign n26192 = ~n13109 & ~n26191;
  assign n26193 = ~n26190 & n26192;
  assign n26194 = ~n13109 & ~n26193;
  assign n26195 = n13029 & ~n13031;
  assign n26196 = ~n13032 & ~n26195;
  assign n26197 = ~n26194 & n26196;
  assign n26198 = ~n13032 & ~n26197;
  assign n26199 = n12675 & n54536;
  assign n26200 = ~n54536 & ~n12681;
  assign n26201 = ~n12675 & ~n12681;
  assign n26202 = ~n26200 & ~n26201;
  assign n26203 = ~n12681 & ~n26199;
  assign n26204 = ~n26198 & ~n56537;
  assign n26205 = ~n12681 & ~n26204;
  assign n26206 = n12638 & ~n26205;
  assign n26207 = ~n12636 & ~n26206;
  assign n26208 = n54428 & n11420;
  assign n26209 = ~n11421 & ~n26208;
  assign n26210 = ~n26207 & n26209;
  assign n26211 = ~n11421 & ~n26210;
  assign n26212 = ~n11259 & n54415;
  assign n26213 = ~n11311 & ~n26212;
  assign n26214 = ~n26211 & n26213;
  assign n26215 = ~n11311 & ~n26214;
  assign n26216 = n11257 & ~n26215;
  assign n26217 = ~n11255 & ~n26216;
  assign n26218 = n10576 & ~n26217;
  assign n26219 = ~n10574 & ~n26218;
  assign n26220 = n407 & n53484;
  assign n26221 = ~n443 & ~n630;
  assign n26222 = ~n630 & ~n1081;
  assign n26223 = ~n443 & n26222;
  assign n26224 = ~n1081 & n26221;
  assign n26225 = n798 & n56538;
  assign n26226 = n804 & n7093;
  assign n26227 = n26220 & n56539;
  assign n26228 = n53630 & n26227;
  assign n26229 = n798 & n53641;
  assign n26230 = n26220 & n26229;
  assign n26231 = n53630 & n26230;
  assign n26232 = ~n1081 & n26231;
  assign n26233 = ~n630 & n26232;
  assign n26234 = ~n443 & n26233;
  assign n26235 = n53641 & n26228;
  assign n26236 = n53487 & n56540;
  assign n26237 = ~n53487 & ~n56540;
  assign n26238 = ~n26236 & ~n26237;
  assign n26239 = ~n875 & ~n26238;
  assign n26240 = ~n26219 & n26239;
  assign n26241 = n26219 & ~n26239;
  assign n26242 = ~n26240 & ~n26241;
  assign n26243 = ~n10576 & n26217;
  assign n26244 = ~n26218 & ~n26243;
  assign n26245 = n26242 & n26244;
  assign n26246 = ~n11257 & n26215;
  assign n26247 = ~n26216 & ~n26246;
  assign n26248 = n26244 & n26247;
  assign n26249 = n26211 & ~n26213;
  assign n26250 = ~n26214 & ~n26249;
  assign n26251 = n26247 & n26250;
  assign n26252 = n26207 & ~n26209;
  assign n26253 = ~n26210 & ~n26252;
  assign n26254 = n26250 & n26253;
  assign n26255 = ~n12638 & n26205;
  assign n26256 = ~n26206 & ~n26255;
  assign n26257 = n26253 & n26256;
  assign n26258 = n26198 & n56537;
  assign n26259 = ~n26204 & ~n26258;
  assign n26260 = n26256 & n26259;
  assign n26261 = n26194 & ~n26196;
  assign n26262 = ~n26197 & ~n26261;
  assign n26263 = n26259 & n26262;
  assign n26264 = n26190 & ~n26192;
  assign n26265 = ~n26193 & ~n26264;
  assign n26266 = n26262 & n26265;
  assign n26267 = n26186 & ~n26188;
  assign n26268 = ~n26189 & ~n26267;
  assign n26269 = n26265 & n26268;
  assign n26270 = ~n14231 & n26184;
  assign n26271 = ~n26185 & ~n26270;
  assign n26272 = n26268 & n26271;
  assign n26273 = n26180 & ~n26182;
  assign n26274 = ~n26183 & ~n26273;
  assign n26275 = n26271 & n26274;
  assign n26276 = ~n14816 & n26178;
  assign n26277 = ~n26179 & ~n26276;
  assign n26278 = n26274 & n26277;
  assign n26279 = ~n15918 & n26176;
  assign n26280 = ~n26177 & ~n26279;
  assign n26281 = n26277 & n26280;
  assign n26282 = ~n16064 & n26174;
  assign n26283 = ~n26175 & ~n26282;
  assign n26284 = n26280 & n26283;
  assign n26285 = n26170 & ~n26172;
  assign n26286 = ~n26173 & ~n26285;
  assign n26287 = n26283 & n26286;
  assign n26288 = ~n16693 & n26168;
  assign n26289 = ~n26169 & ~n26288;
  assign n26290 = n26286 & n26289;
  assign n26291 = ~n17240 & n26166;
  assign n26292 = ~n26167 & ~n26291;
  assign n26293 = n26289 & n26292;
  assign n26294 = ~n17455 & n26164;
  assign n26295 = ~n26165 & ~n26294;
  assign n26296 = n26292 & n26295;
  assign n26297 = ~n18585 & n26162;
  assign n26298 = ~n26163 & ~n26297;
  assign n26299 = n26295 & n26298;
  assign n26300 = n26158 & ~n26160;
  assign n26301 = ~n26161 & ~n26300;
  assign n26302 = n26298 & n26301;
  assign n26303 = n26154 & ~n26156;
  assign n26304 = ~n26157 & ~n26303;
  assign n26305 = n26301 & n26304;
  assign n26306 = ~n19536 & n26152;
  assign n26307 = ~n26153 & ~n26306;
  assign n26308 = n26304 & n26307;
  assign n26309 = n26148 & ~n26150;
  assign n26310 = ~n26151 & ~n26309;
  assign n26311 = n26307 & n26310;
  assign n26312 = ~n20652 & n26146;
  assign n26313 = ~n26147 & ~n26312;
  assign n26314 = n26310 & n26313;
  assign n26315 = ~n21266 & n26144;
  assign n26316 = ~n26145 & ~n26315;
  assign n26317 = n26313 & n26316;
  assign n26318 = n26140 & ~n26142;
  assign n26319 = ~n26143 & ~n26318;
  assign n26320 = n26316 & n26319;
  assign n26321 = n26136 & ~n26138;
  assign n26322 = ~n26139 & ~n26321;
  assign n26323 = n26319 & n26322;
  assign n26324 = ~n23486 & n26134;
  assign n26325 = ~n26135 & ~n26324;
  assign n26326 = n26322 & n26325;
  assign n26327 = n26130 & ~n26132;
  assign n26328 = ~n26133 & ~n26327;
  assign n26329 = n26325 & n26328;
  assign n26330 = n26126 & ~n26128;
  assign n26331 = ~n26129 & ~n26330;
  assign n26332 = n26328 & n26331;
  assign n26333 = ~n25267 & n26124;
  assign n26334 = ~n26125 & ~n26333;
  assign n26335 = n26331 & n26334;
  assign n26336 = n26120 & ~n26122;
  assign n26337 = ~n26123 & ~n26336;
  assign n26338 = n26334 & n26337;
  assign n26339 = n26116 & ~n26118;
  assign n26340 = ~n26119 & ~n26339;
  assign n26341 = n26337 & n26340;
  assign n26342 = n26112 & ~n26114;
  assign n26343 = ~n26115 & ~n26342;
  assign n26344 = n26340 & n26343;
  assign n26345 = ~n26340 & ~n26343;
  assign n26346 = ~n26344 & ~n26345;
  assign n26347 = n26108 & ~n26110;
  assign n26348 = ~n26111 & ~n26347;
  assign n26349 = n56533 & n56536;
  assign n26350 = ~n56533 & ~n26107;
  assign n26351 = ~n56533 & n56536;
  assign n26352 = ~n56536 & ~n26107;
  assign n26353 = n56533 & ~n56536;
  assign n26354 = ~n56541 & ~n56542;
  assign n26355 = ~n26107 & ~n26349;
  assign n26356 = ~n26343 & n56543;
  assign n26357 = n26343 & n26348;
  assign n26358 = n26348 & ~n56543;
  assign n26359 = ~n26343 & n26358;
  assign n26360 = ~n26357 & ~n26359;
  assign n26361 = n26348 & ~n26356;
  assign n26362 = n26346 & ~n56544;
  assign n26363 = ~n26344 & ~n26362;
  assign n26364 = ~n26337 & ~n26340;
  assign n26365 = ~n26341 & ~n26364;
  assign n26366 = ~n26363 & n26365;
  assign n26367 = ~n26341 & ~n26366;
  assign n26368 = ~n26334 & ~n26337;
  assign n26369 = ~n26338 & ~n26368;
  assign n26370 = ~n26338 & ~n26367;
  assign n26371 = ~n26368 & n26370;
  assign n26372 = ~n26367 & n26369;
  assign n26373 = ~n26338 & ~n56545;
  assign n26374 = ~n26331 & ~n26334;
  assign n26375 = ~n26335 & ~n26374;
  assign n26376 = ~n26373 & ~n26374;
  assign n26377 = ~n26335 & n26376;
  assign n26378 = ~n26373 & n26375;
  assign n26379 = ~n26335 & ~n56546;
  assign n26380 = ~n26328 & ~n26331;
  assign n26381 = ~n26332 & ~n26380;
  assign n26382 = ~n26379 & n26381;
  assign n26383 = ~n26332 & ~n26382;
  assign n26384 = ~n26325 & ~n26328;
  assign n26385 = ~n26329 & ~n26384;
  assign n26386 = ~n26383 & ~n26384;
  assign n26387 = ~n26329 & n26386;
  assign n26388 = ~n26383 & n26385;
  assign n26389 = ~n26329 & ~n56547;
  assign n26390 = ~n26322 & ~n26325;
  assign n26391 = ~n26326 & ~n26390;
  assign n26392 = ~n26389 & ~n26390;
  assign n26393 = ~n26326 & n26392;
  assign n26394 = ~n26389 & n26391;
  assign n26395 = ~n26326 & ~n56548;
  assign n26396 = ~n26319 & ~n26322;
  assign n26397 = ~n26323 & ~n26396;
  assign n26398 = ~n26395 & n26397;
  assign n26399 = ~n26323 & ~n26398;
  assign n26400 = ~n26316 & ~n26319;
  assign n26401 = ~n26320 & ~n26400;
  assign n26402 = ~n26399 & ~n26400;
  assign n26403 = ~n26320 & n26402;
  assign n26404 = ~n26399 & n26401;
  assign n26405 = ~n26320 & ~n56549;
  assign n26406 = ~n26313 & ~n26316;
  assign n26407 = ~n26317 & ~n26406;
  assign n26408 = ~n26405 & n26407;
  assign n26409 = ~n26317 & ~n26408;
  assign n26410 = ~n26310 & ~n26313;
  assign n26411 = ~n26314 & ~n26410;
  assign n26412 = ~n26409 & ~n26410;
  assign n26413 = ~n26314 & n26412;
  assign n26414 = ~n26409 & n26411;
  assign n26415 = ~n26314 & ~n56550;
  assign n26416 = ~n26307 & ~n26310;
  assign n26417 = ~n26311 & ~n26416;
  assign n26418 = ~n26415 & ~n26416;
  assign n26419 = ~n26311 & n26418;
  assign n26420 = ~n26415 & n26417;
  assign n26421 = ~n26311 & ~n56551;
  assign n26422 = ~n26304 & ~n26307;
  assign n26423 = ~n26308 & ~n26422;
  assign n26424 = ~n26421 & ~n26422;
  assign n26425 = ~n26308 & n26424;
  assign n26426 = ~n26421 & n26423;
  assign n26427 = ~n26308 & ~n56552;
  assign n26428 = ~n26301 & ~n26304;
  assign n26429 = ~n26305 & ~n26428;
  assign n26430 = ~n26427 & n26429;
  assign n26431 = ~n26305 & ~n26430;
  assign n26432 = ~n26298 & ~n26301;
  assign n26433 = ~n26302 & ~n26432;
  assign n26434 = ~n26431 & ~n26432;
  assign n26435 = ~n26302 & n26434;
  assign n26436 = ~n26431 & n26433;
  assign n26437 = ~n26302 & ~n56553;
  assign n26438 = ~n26295 & ~n26298;
  assign n26439 = ~n26299 & ~n26438;
  assign n26440 = ~n26437 & n26439;
  assign n26441 = ~n26299 & ~n26440;
  assign n26442 = ~n26292 & ~n26295;
  assign n26443 = ~n26296 & ~n26442;
  assign n26444 = ~n26441 & n26443;
  assign n26445 = ~n26296 & ~n26444;
  assign n26446 = ~n26289 & ~n26292;
  assign n26447 = ~n26293 & ~n26446;
  assign n26448 = ~n26445 & n26447;
  assign n26449 = ~n26293 & ~n26448;
  assign n26450 = ~n26286 & ~n26289;
  assign n26451 = ~n26290 & ~n26450;
  assign n26452 = ~n26449 & ~n26450;
  assign n26453 = ~n26290 & n26452;
  assign n26454 = ~n26449 & n26451;
  assign n26455 = ~n26290 & ~n56554;
  assign n26456 = ~n26283 & ~n26286;
  assign n26457 = ~n26287 & ~n26456;
  assign n26458 = ~n26455 & ~n26456;
  assign n26459 = ~n26287 & n26458;
  assign n26460 = ~n26455 & n26457;
  assign n26461 = ~n26287 & ~n56555;
  assign n26462 = ~n26280 & ~n26283;
  assign n26463 = ~n26284 & ~n26462;
  assign n26464 = ~n26461 & n26463;
  assign n26465 = ~n26284 & ~n26464;
  assign n26466 = ~n26277 & ~n26280;
  assign n26467 = ~n26281 & ~n26466;
  assign n26468 = ~n26465 & n26467;
  assign n26469 = ~n26281 & ~n26468;
  assign n26470 = ~n26274 & ~n26277;
  assign n26471 = ~n26278 & ~n26470;
  assign n26472 = ~n26469 & ~n26470;
  assign n26473 = ~n26278 & n26472;
  assign n26474 = ~n26469 & n26471;
  assign n26475 = ~n26278 & ~n56556;
  assign n26476 = ~n26271 & ~n26274;
  assign n26477 = ~n26275 & ~n26476;
  assign n26478 = ~n26475 & ~n26476;
  assign n26479 = ~n26275 & n26478;
  assign n26480 = ~n26475 & n26477;
  assign n26481 = ~n26275 & ~n56557;
  assign n26482 = ~n26268 & ~n26271;
  assign n26483 = ~n26272 & ~n26482;
  assign n26484 = ~n26481 & ~n26482;
  assign n26485 = ~n26272 & n26484;
  assign n26486 = ~n26481 & n26483;
  assign n26487 = ~n26272 & ~n56558;
  assign n26488 = ~n26265 & ~n26268;
  assign n26489 = ~n26269 & ~n26488;
  assign n26490 = ~n26487 & n26489;
  assign n26491 = ~n26269 & ~n26490;
  assign n26492 = ~n26262 & ~n26265;
  assign n26493 = ~n26266 & ~n26492;
  assign n26494 = ~n26491 & n26493;
  assign n26495 = ~n26266 & ~n26494;
  assign n26496 = ~n26259 & ~n26262;
  assign n26497 = ~n26263 & ~n26496;
  assign n26498 = ~n26495 & ~n26496;
  assign n26499 = ~n26263 & n26498;
  assign n26500 = ~n26495 & n26497;
  assign n26501 = ~n26263 & ~n56559;
  assign n26502 = ~n26256 & ~n26259;
  assign n26503 = ~n26260 & ~n26502;
  assign n26504 = ~n26501 & n26503;
  assign n26505 = ~n26260 & ~n26504;
  assign n26506 = ~n26253 & ~n26256;
  assign n26507 = ~n26257 & ~n26506;
  assign n26508 = ~n26505 & ~n26506;
  assign n26509 = ~n26257 & n26508;
  assign n26510 = ~n26505 & n26507;
  assign n26511 = ~n26257 & ~n56560;
  assign n26512 = ~n26250 & ~n26253;
  assign n26513 = ~n26254 & ~n26512;
  assign n26514 = ~n26511 & n26513;
  assign n26515 = ~n26254 & ~n26514;
  assign n26516 = ~n26247 & ~n26250;
  assign n26517 = ~n26251 & ~n26516;
  assign n26518 = ~n26515 & ~n26516;
  assign n26519 = ~n26251 & n26518;
  assign n26520 = ~n26515 & n26517;
  assign n26521 = ~n26251 & ~n56561;
  assign n26522 = ~n26244 & ~n26247;
  assign n26523 = ~n26248 & ~n26522;
  assign n26524 = ~n26521 & n26523;
  assign n26525 = ~n26248 & ~n26524;
  assign n26526 = ~n26242 & ~n26244;
  assign n26527 = ~n26245 & ~n26526;
  assign n26528 = ~n26525 & n26527;
  assign n26529 = ~n26245 & ~n26528;
  assign n26530 = ~n875 & ~n26240;
  assign n26531 = n1642 & ~n1658;
  assign n26532 = n53623 & n26531;
  assign n26533 = n1657 & ~n1658;
  assign n26534 = n53622 & n56562;
  assign n26535 = ~n1658 & n53569;
  assign n26536 = ~n26236 & ~n56563;
  assign n26537 = n26530 & ~n26536;
  assign n26538 = n26242 & ~n26537;
  assign n26539 = ~n26529 & ~n26538;
  assign n26540 = n26529 & n26538;
  assign n26541 = ~n26538 & ~n26539;
  assign n26542 = ~n26529 & ~n26539;
  assign n26543 = ~n26541 & ~n26542;
  assign n26544 = ~n26539 & ~n26540;
  assign n26545 = n90 & ~n56564;
  assign n26546 = n14236 & ~n26537;
  assign n26547 = n54667 & n26244;
  assign n26548 = n14210 & n26242;
  assign n26549 = ~n26547 & ~n26548;
  assign n26550 = ~n26546 & n26549;
  assign n26551 = ~n26545 & n26550;
  assign n26552 = pi23  & ~n26551;
  assign n26553 = pi23  & ~n26552;
  assign n26554 = pi23  & n26551;
  assign n26555 = ~n26551 & ~n26552;
  assign n26556 = ~pi23  & ~n26551;
  assign n26557 = ~n56565 & ~n56566;
  assign n26558 = n26515 & ~n26517;
  assign n26559 = ~n26515 & ~n56561;
  assign n26560 = ~n26516 & n26521;
  assign n26561 = ~n26559 & ~n26560;
  assign n26562 = ~n56561 & ~n26558;
  assign n26563 = n123 & ~n56567;
  assign n26564 = n128 & n26247;
  assign n26565 = n53444 & n26253;
  assign n26566 = n127 & n26250;
  assign n26567 = ~n26565 & ~n26566;
  assign n26568 = ~n26564 & n26567;
  assign n26569 = ~n26563 & n26568;
  assign n26570 = pi26  & ~n26569;
  assign n26571 = pi26  & ~n26570;
  assign n26572 = pi26  & n26569;
  assign n26573 = ~n26569 & ~n26570;
  assign n26574 = ~pi26  & ~n26569;
  assign n26575 = ~n56568 & ~n56569;
  assign n26576 = n7646 & n8091;
  assign n26577 = n7646 & n13230;
  assign n26578 = n8091 & n26577;
  assign n26579 = n13230 & n26576;
  assign n26580 = ~n250 & ~n567;
  assign n26581 = ~n414 & ~n1065;
  assign n26582 = ~n567 & ~n1065;
  assign n26583 = ~n250 & ~n414;
  assign n26584 = n26582 & n26583;
  assign n26585 = n26580 & n26581;
  assign n26586 = n55089 & n56571;
  assign n26587 = n8091 & n55089;
  assign n26588 = n7646 & n26587;
  assign n26589 = ~n1065 & n26588;
  assign n26590 = ~n414 & n26589;
  assign n26591 = ~n567 & n26590;
  assign n26592 = ~n250 & n26591;
  assign n26593 = ~n553 & n26592;
  assign n26594 = ~n788 & n26593;
  assign n26595 = n56570 & n26586;
  assign n26596 = n752 & ~n1125;
  assign n26597 = ~n1125 & n1711;
  assign n26598 = n752 & n26597;
  assign n26599 = n1711 & n26596;
  assign n26600 = n9331 & n56573;
  assign n26601 = ~n584 & n1534;
  assign n26602 = ~n215 & ~n1234;
  assign n26603 = n2193 & n26602;
  assign n26604 = ~n215 & n8268;
  assign n26605 = ~n584 & n26604;
  assign n26606 = ~n852 & n26605;
  assign n26607 = ~n443 & n26606;
  assign n26608 = ~n753 & n26607;
  assign n26609 = ~n584 & ~n852;
  assign n26610 = ~n215 & n26609;
  assign n26611 = n1534 & n8268;
  assign n26612 = n26610 & n26611;
  assign n26613 = n26601 & n26603;
  assign n26614 = n54769 & n56574;
  assign n26615 = n26600 & n26614;
  assign n26616 = n1711 & n54769;
  assign n26617 = n56572 & n26616;
  assign n26618 = n56574 & n26617;
  assign n26619 = n9331 & n26618;
  assign n26620 = ~n1125 & n26619;
  assign n26621 = ~n751 & n26620;
  assign n26622 = ~n750 & n26621;
  assign n26623 = n56572 & n26615;
  assign n26624 = ~n272 & ~n568;
  assign n26625 = ~n464 & ~n1466;
  assign n26626 = ~n568 & ~n1466;
  assign n26627 = ~n272 & ~n464;
  assign n26628 = n26626 & n26627;
  assign n26629 = n26624 & n26625;
  assign n26630 = n1702 & n4020;
  assign n26631 = n56576 & n26630;
  assign n26632 = n13598 & n26631;
  assign n26633 = ~n259 & ~n319;
  assign n26634 = ~n1090 & ~n1471;
  assign n26635 = n26633 & n26634;
  assign n26636 = ~n295 & ~n617;
  assign n26637 = ~n174 & ~n1641;
  assign n26638 = n26636 & n26637;
  assign n26639 = ~n174 & ~n1090;
  assign n26640 = ~n295 & ~n1471;
  assign n26641 = ~n1090 & n26640;
  assign n26642 = ~n174 & n26641;
  assign n26643 = n26639 & n26640;
  assign n26644 = ~n259 & n56577;
  assign n26645 = ~n319 & n26644;
  assign n26646 = ~n1641 & n26645;
  assign n26647 = ~n617 & n26646;
  assign n26648 = ~n319 & ~n1641;
  assign n26649 = n26636 & n26648;
  assign n26650 = ~n259 & ~n1090;
  assign n26651 = ~n174 & ~n1471;
  assign n26652 = n26650 & n26651;
  assign n26653 = n26649 & n26652;
  assign n26654 = ~n617 & ~n1641;
  assign n26655 = n26633 & n26654;
  assign n26656 = n56577 & n26655;
  assign n26657 = n26635 & n26638;
  assign n26658 = n1542 & n5874;
  assign n26659 = n9510 & n26658;
  assign n26660 = n56578 & n26659;
  assign n26661 = n4020 & n5874;
  assign n26662 = n56576 & n26661;
  assign n26663 = n13598 & n26662;
  assign n26664 = n1542 & n1702;
  assign n26665 = n9510 & n26664;
  assign n26666 = n56578 & n26665;
  assign n26667 = n26663 & n26666;
  assign n26668 = n5874 & n9510;
  assign n26669 = n56576 & n26668;
  assign n26670 = n13598 & n26669;
  assign n26671 = n1542 & n26630;
  assign n26672 = n4020 & n26664;
  assign n26673 = n56578 & n56580;
  assign n26674 = n26670 & n26673;
  assign n26675 = n26632 & n26660;
  assign n26676 = ~n513 & n4317;
  assign n26677 = ~n647 & n26676;
  assign n26678 = n4317 & n11562;
  assign n26679 = n54630 & n56581;
  assign n26680 = ~n340 & ~n773;
  assign n26681 = ~n218 & ~n258;
  assign n26682 = n26680 & n26681;
  assign n26683 = ~n614 & ~n2042;
  assign n26684 = n7045 & n26683;
  assign n26685 = ~n258 & ~n773;
  assign n26686 = ~n218 & ~n614;
  assign n26687 = n26685 & n26686;
  assign n26688 = ~n340 & ~n2042;
  assign n26689 = n7045 & n26688;
  assign n26690 = n26687 & n26689;
  assign n26691 = n26682 & n26684;
  assign n26692 = ~n614 & ~n773;
  assign n26693 = ~n218 & ~n340;
  assign n26694 = ~n2042 & n26693;
  assign n26695 = n26692 & n26694;
  assign n26696 = ~n258 & n7045;
  assign n26697 = n7045 & n54630;
  assign n26698 = n56581 & n26697;
  assign n26699 = ~n258 & n26698;
  assign n26700 = n54630 & n26696;
  assign n26701 = n56581 & n26700;
  assign n26702 = n26679 & n26696;
  assign n26703 = n26695 & n56583;
  assign n26704 = ~n218 & n56583;
  assign n26705 = ~n340 & n26704;
  assign n26706 = ~n773 & n26705;
  assign n26707 = ~n614 & n26706;
  assign n26708 = ~n2042 & n26707;
  assign n26709 = n26679 & n56582;
  assign n26710 = ~n628 & ~n957;
  assign n26711 = ~n957 & ~n1196;
  assign n26712 = ~n628 & n26711;
  assign n26713 = ~n1196 & n26710;
  assign n26714 = ~n353 & n4262;
  assign n26715 = ~n353 & n6482;
  assign n26716 = n4262 & n26715;
  assign n26717 = n6482 & n26714;
  assign n26718 = n4262 & n56585;
  assign n26719 = n6482 & n26718;
  assign n26720 = ~n353 & n26719;
  assign n26721 = n56585 & n56586;
  assign n26722 = n56584 & n56587;
  assign n26723 = n56579 & n56587;
  assign n26724 = n56584 & n26723;
  assign n26725 = n56579 & n26722;
  assign n26726 = n56575 & n56588;
  assign n26727 = n9510 & n56580;
  assign n26728 = n56587 & n26727;
  assign n26729 = n56575 & n26728;
  assign n26730 = n54290 & n26729;
  assign n26731 = n56584 & n26730;
  assign n26732 = n56578 & n26731;
  assign n26733 = n5874 & n26732;
  assign n26734 = n13598 & n26733;
  assign n26735 = ~n464 & n26734;
  assign n26736 = ~n1466 & n26735;
  assign n26737 = ~n272 & n26736;
  assign n26738 = ~n568 & n26737;
  assign n26739 = n54290 & n26726;
  assign n26740 = ~n822 & ~n1059;
  assign n26741 = n3877 & n26740;
  assign n26742 = n6563 & n10182;
  assign n26743 = ~n881 & n10182;
  assign n26744 = ~n894 & n26743;
  assign n26745 = ~n2103 & n26744;
  assign n26746 = ~n311 & n26745;
  assign n26747 = ~n1059 & n26746;
  assign n26748 = ~n822 & n26747;
  assign n26749 = ~n822 & ~n881;
  assign n26750 = ~n311 & ~n2103;
  assign n26751 = n26749 & n26750;
  assign n26752 = ~n894 & ~n1059;
  assign n26753 = n10182 & n26752;
  assign n26754 = n26751 & n26753;
  assign n26755 = n26741 & n26742;
  assign n26756 = n903 & n1184;
  assign n26757 = ~n172 & ~n464;
  assign n26758 = n10901 & n26757;
  assign n26759 = n26756 & n26758;
  assign n26760 = ~n177 & ~n357;
  assign n26761 = n347 & n26760;
  assign n26762 = n1277 & n3522;
  assign n26763 = n26761 & n26762;
  assign n26764 = n26759 & n26763;
  assign n26765 = n56590 & n26764;
  assign n26766 = ~n419 & ~n422;
  assign n26767 = ~n1280 & ~n1476;
  assign n26768 = n26766 & n26767;
  assign n26769 = n54010 & n26768;
  assign n26770 = n54256 & n26769;
  assign n26771 = n54825 & n26770;
  assign n26772 = n347 & n903;
  assign n26773 = n424 & n26757;
  assign n26774 = n26772 & n26773;
  assign n26775 = ~n177 & ~n419;
  assign n26776 = n10901 & n26775;
  assign n26777 = n26762 & n26776;
  assign n26778 = n26774 & n26777;
  assign n26779 = n56590 & n26778;
  assign n26780 = ~n788 & ~n1280;
  assign n26781 = ~n357 & ~n1476;
  assign n26782 = n26780 & n26781;
  assign n26783 = n54010 & n26782;
  assign n26784 = n54256 & n26783;
  assign n26785 = n54825 & n26784;
  assign n26786 = n26779 & n26785;
  assign n26787 = n903 & n3522;
  assign n26788 = n26758 & n26787;
  assign n26789 = n424 & n26780;
  assign n26790 = n347 & n1277;
  assign n26791 = n26789 & n26790;
  assign n26792 = n26788 & n26791;
  assign n26793 = n56590 & n26792;
  assign n26794 = n26775 & n26781;
  assign n26795 = n54010 & n26794;
  assign n26796 = n54256 & n26795;
  assign n26797 = n54825 & n26796;
  assign n26798 = n26793 & n26797;
  assign n26799 = n26765 & n26771;
  assign n26800 = n54227 & n56591;
  assign n26801 = n3522 & n54010;
  assign n26802 = n54256 & n26801;
  assign n26803 = n54227 & n26802;
  assign n26804 = n56590 & n26803;
  assign n26805 = n347 & n26804;
  assign n26806 = n54487 & n26805;
  assign n26807 = n54825 & n26806;
  assign n26808 = n10901 & n26807;
  assign n26809 = n1277 & n26808;
  assign n26810 = n424 & n26809;
  assign n26811 = n903 & n26810;
  assign n26812 = ~n1476 & n26811;
  assign n26813 = n26757 & n26812;
  assign n26814 = ~n177 & n26813;
  assign n26815 = ~n1280 & n26814;
  assign n26816 = ~n419 & n26815;
  assign n26817 = ~n357 & n26816;
  assign n26818 = ~n788 & n26817;
  assign n26819 = n54487 & n26800;
  assign n26820 = ~n361 & ~n404;
  assign n26821 = n318 & ~n404;
  assign n26822 = ~n361 & n26821;
  assign n26823 = n318 & n26820;
  assign n26824 = ~n177 & ~n776;
  assign n26825 = ~n112 & ~n177;
  assign n26826 = ~n824 & n26825;
  assign n26827 = ~n776 & n26826;
  assign n26828 = n5322 & n26824;
  assign n26829 = n55125 & n56594;
  assign n26830 = n55125 & n56593;
  assign n26831 = n56594 & n26830;
  assign n26832 = n56593 & n26829;
  assign n26833 = n421 & n1803;
  assign n26834 = n7144 & n9337;
  assign n26835 = n421 & n9337;
  assign n26836 = n1803 & n7144;
  assign n26837 = n26835 & n26836;
  assign n26838 = n26833 & n26834;
  assign n26839 = ~n491 & ~n567;
  assign n26840 = ~n1125 & ~n1881;
  assign n26841 = ~n567 & ~n1125;
  assign n26842 = ~n491 & ~n1881;
  assign n26843 = n26841 & n26842;
  assign n26844 = n26839 & n26840;
  assign n26845 = n10078 & n56597;
  assign n26846 = n56596 & n26845;
  assign n26847 = n56595 & n26846;
  assign n26848 = n54282 & n26847;
  assign n26849 = n56584 & n26847;
  assign n26850 = n54282 & n26849;
  assign n26851 = n56584 & n26848;
  assign n26852 = n53536 & n54736;
  assign n26853 = n10078 & n56593;
  assign n26854 = n55125 & n26853;
  assign n26855 = n53536 & n26854;
  assign n26856 = n56594 & n26855;
  assign n26857 = n56584 & n26856;
  assign n26858 = n54736 & n26857;
  assign n26859 = n54282 & n26858;
  assign n26860 = n7144 & n26859;
  assign n26861 = n9337 & n26860;
  assign n26862 = n421 & n26861;
  assign n26863 = n1803 & n26862;
  assign n26864 = ~n1125 & n26863;
  assign n26865 = ~n567 & n26864;
  assign n26866 = ~n491 & n26865;
  assign n26867 = ~n1881 & n26866;
  assign n26868 = n56598 & n26852;
  assign n26869 = ~n56592 & ~n56599;
  assign n26870 = ~n16676 & ~n16696;
  assign n26871 = ~n54884 & n26870;
  assign n26872 = ~n16079 & ~n54886;
  assign n26873 = n26870 & n26872;
  assign n26874 = ~n54886 & n26870;
  assign n26875 = ~n16079 & n26874;
  assign n26876 = ~n54884 & n16087;
  assign n26877 = pi17  & n56600;
  assign n26878 = ~pi17  & ~n56600;
  assign n26879 = ~n26877 & ~n26878;
  assign n26880 = n56592 & n56599;
  assign n26881 = ~n26869 & ~n26880;
  assign n26882 = n26879 & n26881;
  assign n26883 = ~n26869 & ~n26882;
  assign n26884 = n56589 & ~n26883;
  assign n26885 = ~n56589 & n26883;
  assign n26886 = ~n26884 & ~n26885;
  assign n26887 = n26481 & ~n26483;
  assign n26888 = ~n26481 & ~n56558;
  assign n26889 = ~n26482 & n26487;
  assign n26890 = ~n26888 & ~n26889;
  assign n26891 = ~n56558 & ~n26887;
  assign n26892 = n1576 & ~n56601;
  assign n26893 = n11215 & n26268;
  assign n26894 = n10564 & n26271;
  assign n26895 = n54403 & n26274;
  assign n26896 = ~n26894 & ~n26895;
  assign n26897 = ~n26893 & n26896;
  assign n26898 = ~n26892 & ~n26895;
  assign n26899 = ~n26894 & n26898;
  assign n26900 = ~n26893 & n26899;
  assign n26901 = ~n26892 & n26897;
  assign n26902 = n26886 & ~n56602;
  assign n26903 = ~n26884 & ~n26902;
  assign n26904 = ~n353 & ~n507;
  assign n26905 = ~n911 & n26904;
  assign n26906 = ~n414 & ~n662;
  assign n26907 = n248 & n26906;
  assign n26908 = ~n911 & n26906;
  assign n26909 = n248 & n26904;
  assign n26910 = n26908 & n26909;
  assign n26911 = n26905 & n26907;
  assign n26912 = n12331 & n54633;
  assign n26913 = n56603 & n26912;
  assign n26914 = ~n977 & n4752;
  assign n26915 = ~n977 & ~n1469;
  assign n26916 = ~n1476 & n26915;
  assign n26917 = ~n161 & n26916;
  assign n26918 = ~n1769 & n26917;
  assign n26919 = n7850 & n26914;
  assign n26920 = n1265 & n3606;
  assign n26921 = n6806 & n10685;
  assign n26922 = n26920 & n26921;
  assign n26923 = n53965 & n26922;
  assign n26924 = n56604 & n26923;
  assign n26925 = ~n507 & ~n662;
  assign n26926 = n6806 & n26925;
  assign n26927 = n4026 & n10685;
  assign n26928 = n26926 & n26927;
  assign n26929 = ~n414 & ~n911;
  assign n26930 = ~n353 & n26929;
  assign n26931 = n54633 & n26930;
  assign n26932 = n26928 & n26931;
  assign n26933 = n248 & n905;
  assign n26934 = n26920 & n26933;
  assign n26935 = n53965 & n26934;
  assign n26936 = n56604 & n26935;
  assign n26937 = n26932 & n26936;
  assign n26938 = ~n353 & ~n414;
  assign n26939 = n3606 & n26938;
  assign n26940 = n905 & n10685;
  assign n26941 = n26939 & n26940;
  assign n26942 = ~n507 & ~n911;
  assign n26943 = ~n662 & n26942;
  assign n26944 = n54633 & n26943;
  assign n26945 = n26941 & n26944;
  assign n26946 = n1265 & n4026;
  assign n26947 = n248 & n6806;
  assign n26948 = n26946 & n26947;
  assign n26949 = n53965 & n26948;
  assign n26950 = n56604 & n26949;
  assign n26951 = n26945 & n26950;
  assign n26952 = n26913 & n26924;
  assign n26953 = n54145 & n56605;
  assign n26954 = ~n733 & ~n771;
  assign n26955 = ~n894 & n26954;
  assign n26956 = n53765 & n26955;
  assign n26957 = n10239 & n26956;
  assign n26958 = n976 & n5199;
  assign n26959 = n1957 & n26958;
  assign n26960 = ~n292 & ~n349;
  assign n26961 = ~n493 & ~n503;
  assign n26962 = n26960 & n26961;
  assign n26963 = ~n258 & ~n659;
  assign n26964 = n3083 & n26963;
  assign n26965 = n26962 & n26964;
  assign n26966 = n26959 & n26965;
  assign n26967 = n976 & n1957;
  assign n26968 = n1186 & n5199;
  assign n26969 = n26967 & n26968;
  assign n26970 = ~n733 & ~n894;
  assign n26971 = ~n292 & ~n503;
  assign n26972 = n26970 & n26971;
  assign n26973 = n2338 & n3083;
  assign n26974 = n26972 & n26973;
  assign n26975 = ~n258 & ~n349;
  assign n26976 = ~n493 & ~n659;
  assign n26977 = n26975 & n26976;
  assign n26978 = n10239 & n26977;
  assign n26979 = ~n349 & ~n493;
  assign n26980 = ~n503 & ~n659;
  assign n26981 = n26979 & n26980;
  assign n26982 = n26973 & n26981;
  assign n26983 = ~n258 & ~n292;
  assign n26984 = n26970 & n26983;
  assign n26985 = n10239 & n26984;
  assign n26986 = n26982 & n26985;
  assign n26987 = n26974 & n26978;
  assign n26988 = n26969 & n56606;
  assign n26989 = n2338 & n5199;
  assign n26990 = n1186 & n3083;
  assign n26991 = n26989 & n26990;
  assign n26992 = ~n258 & ~n894;
  assign n26993 = ~n503 & ~n733;
  assign n26994 = n26992 & n26993;
  assign n26995 = n26967 & n26994;
  assign n26996 = ~n292 & ~n659;
  assign n26997 = n26979 & n26996;
  assign n26998 = n10239 & n26997;
  assign n26999 = n26995 & n26998;
  assign n27000 = n26991 & n26999;
  assign n27001 = n26957 & n26966;
  assign n27002 = n3083 & n10239;
  assign n27003 = n1186 & n27002;
  assign n27004 = n54149 & n27003;
  assign n27005 = n5199 & n27004;
  assign n27006 = n2338 & n27005;
  assign n27007 = n1957 & n27006;
  assign n27008 = n976 & n27007;
  assign n27009 = ~n894 & n27008;
  assign n27010 = ~n659 & n27009;
  assign n27011 = ~n258 & n27010;
  assign n27012 = ~n292 & n27011;
  assign n27013 = ~n493 & n27012;
  assign n27014 = ~n503 & n27013;
  assign n27015 = ~n733 & n27014;
  assign n27016 = ~n349 & n27015;
  assign n27017 = n54149 & n56607;
  assign n27018 = n54818 & n56608;
  assign n27019 = n248 & n54633;
  assign n27020 = n56604 & n27019;
  assign n27021 = n53965 & n27020;
  assign n27022 = n54818 & n27021;
  assign n27023 = n54145 & n27022;
  assign n27024 = n56608 & n27023;
  assign n27025 = n6806 & n27024;
  assign n27026 = n1265 & n27025;
  assign n27027 = n4026 & n27026;
  assign n27028 = n905 & n27027;
  assign n27029 = ~n414 & n27028;
  assign n27030 = ~n957 & n27029;
  assign n27031 = ~n662 & n27030;
  assign n27032 = ~n911 & n27031;
  assign n27033 = n10685 & n27032;
  assign n27034 = ~n507 & n27033;
  assign n27035 = ~n649 & n27034;
  assign n27036 = ~n353 & n27035;
  assign n27037 = n26953 & n27018;
  assign n27038 = n56589 & ~n56609;
  assign n27039 = ~n56589 & n56609;
  assign n27040 = ~n27038 & ~n27039;
  assign n27041 = n26487 & ~n26489;
  assign n27042 = ~n26490 & ~n27041;
  assign n27043 = n1576 & n27042;
  assign n27044 = n11215 & n26265;
  assign n27045 = n54403 & n26271;
  assign n27046 = n10564 & n26268;
  assign n27047 = ~n27045 & ~n27046;
  assign n27048 = ~n27044 & n27047;
  assign n27049 = ~n27043 & n27048;
  assign n27050 = ~n27038 & ~n27049;
  assign n27051 = ~n27039 & n27050;
  assign n27052 = n27040 & ~n27049;
  assign n27053 = ~n27040 & n27049;
  assign n27054 = ~n27049 & ~n56610;
  assign n27055 = ~n27038 & ~n56610;
  assign n27056 = ~n27039 & n27055;
  assign n27057 = ~n27054 & ~n27056;
  assign n27058 = ~n56610 & ~n27053;
  assign n27059 = ~n26903 & ~n56611;
  assign n27060 = n26903 & n56611;
  assign n27061 = ~n27059 & ~n27060;
  assign n27062 = ~n26879 & ~n26881;
  assign n27063 = ~n26882 & ~n27062;
  assign n27064 = n26475 & ~n26477;
  assign n27065 = ~n26475 & ~n56557;
  assign n27066 = ~n26476 & n26481;
  assign n27067 = ~n27065 & ~n27066;
  assign n27068 = ~n56557 & ~n27064;
  assign n27069 = n1576 & ~n56612;
  assign n27070 = n11215 & n26271;
  assign n27071 = n54403 & n26277;
  assign n27072 = n10564 & n26274;
  assign n27073 = ~n27071 & ~n27072;
  assign n27074 = ~n27070 & n27073;
  assign n27075 = ~n27069 & n27074;
  assign n27076 = n27063 & ~n27075;
  assign n27077 = ~n440 & ~n504;
  assign n27078 = n12286 & n14519;
  assign n27079 = n27077 & n27078;
  assign n27080 = ~n271 & ~n647;
  assign n27081 = ~n141 & ~n1192;
  assign n27082 = ~n647 & ~n1192;
  assign n27083 = ~n141 & ~n271;
  assign n27084 = n27082 & n27083;
  assign n27085 = n27080 & n27081;
  assign n27086 = n906 & n10298;
  assign n27087 = n56613 & n27086;
  assign n27088 = n906 & n12286;
  assign n27089 = n27077 & n27088;
  assign n27090 = n10298 & n27081;
  assign n27091 = n14519 & n27080;
  assign n27092 = n27090 & n27091;
  assign n27093 = n27089 & n27092;
  assign n27094 = n27079 & n27087;
  assign n27095 = ~n296 & ~n956;
  assign n27096 = ~n922 & ~n1490;
  assign n27097 = n27095 & n27096;
  assign n27098 = ~n902 & ~n922;
  assign n27099 = ~n296 & n27098;
  assign n27100 = ~n1490 & n27099;
  assign n27101 = ~n956 & n27100;
  assign n27102 = ~n447 & n27101;
  assign n27103 = ~n447 & ~n1490;
  assign n27104 = ~n902 & ~n956;
  assign n27105 = ~n296 & ~n922;
  assign n27106 = n27104 & n27105;
  assign n27107 = n27103 & n27106;
  assign n27108 = n1360 & n27097;
  assign n27109 = n54987 & n56615;
  assign n27110 = n56614 & n27109;
  assign n27111 = n12286 & n27077;
  assign n27112 = n56615 & n27111;
  assign n27113 = n54628 & n27112;
  assign n27114 = n54987 & n27113;
  assign n27115 = n906 & n27114;
  assign n27116 = ~n295 & n27115;
  assign n27117 = ~n1192 & n27116;
  assign n27118 = ~n662 & n27117;
  assign n27119 = ~n271 & n27118;
  assign n27120 = ~n141 & n27119;
  assign n27121 = ~n568 & n27120;
  assign n27122 = ~n647 & n27121;
  assign n27123 = ~n751 & n27122;
  assign n27124 = n54628 & n27110;
  assign n27125 = ~n2109 & n7277;
  assign n27126 = ~n1472 & n10238;
  assign n27127 = n10238 & n56616;
  assign n27128 = ~n1472 & n27127;
  assign n27129 = n56616 & n56617;
  assign n27130 = n1032 & n3878;
  assign n27131 = n6150 & n9453;
  assign n27132 = n3878 & n6150;
  assign n27133 = n1032 & n9453;
  assign n27134 = n27132 & n27133;
  assign n27135 = n27130 & n27131;
  assign n27136 = ~n1465 & n4478;
  assign n27137 = ~n215 & ~n788;
  assign n27138 = n180 & n27137;
  assign n27139 = ~n215 & ~n1088;
  assign n27140 = ~n1478 & n27139;
  assign n27141 = n180 & n1697;
  assign n27142 = n27140 & n27141;
  assign n27143 = n27136 & n27138;
  assign n27144 = n180 & n6150;
  assign n27145 = n3878 & n27144;
  assign n27146 = n1032 & n27145;
  assign n27147 = n27130 & n27144;
  assign n27148 = ~n1088 & n56621;
  assign n27149 = ~n1465 & n27148;
  assign n27150 = ~n1478 & n27149;
  assign n27151 = ~n215 & n27150;
  assign n27152 = ~n206 & n27151;
  assign n27153 = ~n364 & n27152;
  assign n27154 = ~n788 & n27153;
  assign n27155 = ~n206 & ~n1478;
  assign n27156 = ~n1088 & n27155;
  assign n27157 = ~n364 & ~n1465;
  assign n27158 = n27137 & n27157;
  assign n27159 = n27156 & n27158;
  assign n27160 = n56621 & n27159;
  assign n27161 = n56619 & n56620;
  assign n27162 = ~n443 & ~n451;
  assign n27163 = ~n1127 & n27162;
  assign n27164 = n53992 & n27163;
  assign n27165 = n7144 & n9477;
  assign n27166 = n54137 & n27165;
  assign n27167 = n27164 & n27166;
  assign n27168 = n976 & n2476;
  assign n27169 = ~n416 & ~n465;
  assign n27170 = n13427 & n27169;
  assign n27171 = n2476 & n13427;
  assign n27172 = n976 & n27169;
  assign n27173 = n27171 & n27172;
  assign n27174 = n27168 & n27170;
  assign n27175 = n54376 & n56623;
  assign n27176 = ~n451 & ~n879;
  assign n27177 = ~n1127 & n27176;
  assign n27178 = ~n404 & ~n443;
  assign n27179 = n27169 & n27178;
  assign n27180 = n27177 & n27179;
  assign n27181 = n53992 & n54137;
  assign n27182 = n27180 & n27181;
  assign n27183 = n27165 & n27168;
  assign n27184 = n54376 & n27183;
  assign n27185 = n27182 & n27184;
  assign n27186 = n27167 & n27175;
  assign n27187 = n56622 & n56624;
  assign n27188 = n54312 & n27187;
  assign n27189 = n53992 & n56618;
  assign n27190 = n54137 & n27189;
  assign n27191 = n54376 & n27190;
  assign n27192 = n54312 & n27191;
  assign n27193 = n56622 & n27192;
  assign n27194 = n7144 & n27193;
  assign n27195 = n9477 & n27194;
  assign n27196 = n2476 & n27195;
  assign n27197 = n976 & n27196;
  assign n27198 = ~n416 & n27197;
  assign n27199 = ~n1127 & n27198;
  assign n27200 = ~n879 & n27199;
  assign n27201 = ~n404 & n27200;
  assign n27202 = ~n443 & n27201;
  assign n27203 = ~n465 & n27202;
  assign n27204 = ~n451 & n27203;
  assign n27205 = n56618 & n27188;
  assign n27206 = n56592 & ~n56625;
  assign n27207 = ~n247 & ~n1125;
  assign n27208 = ~n1125 & n54787;
  assign n27209 = ~n247 & n27208;
  assign n27210 = n54787 & n27207;
  assign n27211 = n2627 & n11134;
  assign n27212 = ~n770 & ~n1490;
  assign n27213 = ~n408 & ~n851;
  assign n27214 = n27212 & n27213;
  assign n27215 = n27211 & n27214;
  assign n27216 = ~n207 & ~n353;
  assign n27217 = n1266 & n27216;
  assign n27218 = n54826 & n27217;
  assign n27219 = n1266 & n2627;
  assign n27220 = n27214 & n27219;
  assign n27221 = n11134 & n27216;
  assign n27222 = n54826 & n27221;
  assign n27223 = n27220 & n27222;
  assign n27224 = n2627 & n27213;
  assign n27225 = n1266 & n11134;
  assign n27226 = n27224 & n27225;
  assign n27227 = ~n353 & ~n1490;
  assign n27228 = ~n207 & ~n770;
  assign n27229 = n27227 & n27228;
  assign n27230 = n54826 & n27229;
  assign n27231 = n27226 & n27230;
  assign n27232 = n27215 & n27218;
  assign n27233 = n53958 & n56627;
  assign n27234 = n54338 & n27233;
  assign n27235 = n53764 & n27234;
  assign n27236 = n54826 & n56626;
  assign n27237 = n1266 & n27236;
  assign n27238 = n54338 & n27237;
  assign n27239 = n53764 & n27238;
  assign n27240 = n11134 & n27239;
  assign n27241 = n53958 & n27240;
  assign n27242 = ~n408 & n27241;
  assign n27243 = ~n1490 & n27242;
  assign n27244 = ~n207 & n27243;
  assign n27245 = n2627 & n27244;
  assign n27246 = ~n851 & n27245;
  assign n27247 = ~n353 & n27246;
  assign n27248 = ~n770 & n27247;
  assign n27249 = n56626 & n27235;
  assign n27250 = ~n441 & ~n560;
  assign n27251 = ~n441 & ~n1192;
  assign n27252 = ~n560 & n27251;
  assign n27253 = ~n1192 & n27250;
  assign n27254 = ~n292 & ~n401;
  assign n27255 = n1850 & n27254;
  assign n27256 = n56629 & n27255;
  assign n27257 = n53820 & n27256;
  assign n27258 = ~n274 & ~n2109;
  assign n27259 = n4530 & n27258;
  assign n27260 = ~n507 & ~n1195;
  assign n27261 = n906 & n27260;
  assign n27262 = n906 & n4530;
  assign n27263 = ~n1195 & n27262;
  assign n27264 = ~n274 & n27263;
  assign n27265 = ~n507 & n27264;
  assign n27266 = ~n2109 & n27265;
  assign n27267 = n906 & n27258;
  assign n27268 = n4530 & n27260;
  assign n27269 = n27267 & n27268;
  assign n27270 = ~n274 & ~n507;
  assign n27271 = ~n1195 & ~n2109;
  assign n27272 = n27270 & n27271;
  assign n27273 = n27262 & n27272;
  assign n27274 = n27259 & n27261;
  assign n27275 = n54473 & n56630;
  assign n27276 = n27257 & n27275;
  assign n27277 = n1091 & n2974;
  assign n27278 = n54624 & n13955;
  assign n27279 = n27277 & n27278;
  assign n27280 = n54100 & n27279;
  assign n27281 = ~n401 & ~n560;
  assign n27282 = ~n292 & ~n441;
  assign n27283 = n27281 & n27282;
  assign n27284 = n13955 & n27283;
  assign n27285 = n53820 & n27284;
  assign n27286 = n27275 & n27285;
  assign n27287 = ~n771 & ~n1192;
  assign n27288 = ~n354 & n27287;
  assign n27289 = n54624 & n27288;
  assign n27290 = n27277 & n27289;
  assign n27291 = n54100 & n27290;
  assign n27292 = n27286 & n27291;
  assign n27293 = n27276 & n27280;
  assign n27294 = n54112 & n56631;
  assign n27295 = n6481 & n27277;
  assign n27296 = n54624 & n27295;
  assign n27297 = n54473 & n27296;
  assign n27298 = n53820 & n27297;
  assign n27299 = n56630 & n27298;
  assign n27300 = n54112 & n27299;
  assign n27301 = n55100 & n27300;
  assign n27302 = n1078 & n27301;
  assign n27303 = n54100 & n27302;
  assign n27304 = ~n1192 & n27303;
  assign n27305 = ~n292 & n27304;
  assign n27306 = ~n560 & n27305;
  assign n27307 = ~n401 & n27306;
  assign n27308 = ~n441 & n27307;
  assign n27309 = ~n354 & n27308;
  assign n27310 = ~n771 & n27309;
  assign n27311 = n55100 & n27294;
  assign n27312 = ~n56628 & ~n56632;
  assign n27313 = ~n18556 & ~n18588;
  assign n27314 = ~n55041 & ~n17265;
  assign n27315 = n27313 & n27314;
  assign n27316 = ~n55041 & n27313;
  assign n27317 = ~n17265 & n27316;
  assign n27318 = n17255 & ~n55040;
  assign n27319 = pi14  & n56633;
  assign n27320 = ~pi14  & ~n56633;
  assign n27321 = ~n27319 & ~n27320;
  assign n27322 = n56628 & n56632;
  assign n27323 = ~n27312 & ~n27322;
  assign n27324 = n27321 & n27323;
  assign n27325 = ~n27312 & ~n27324;
  assign n27326 = n56625 & ~n27325;
  assign n27327 = ~n56625 & n27325;
  assign n27328 = ~n27326 & ~n27327;
  assign n27329 = n26465 & ~n26467;
  assign n27330 = ~n26468 & ~n27329;
  assign n27331 = n1576 & n27330;
  assign n27332 = n11215 & n26277;
  assign n27333 = n10564 & n26280;
  assign n27334 = n54403 & n26283;
  assign n27335 = ~n27333 & ~n27334;
  assign n27336 = ~n27332 & n27335;
  assign n27337 = ~n27331 & ~n27334;
  assign n27338 = ~n27333 & n27337;
  assign n27339 = ~n27332 & n27338;
  assign n27340 = ~n27331 & n27336;
  assign n27341 = n27328 & ~n56634;
  assign n27342 = ~n27326 & ~n27341;
  assign n27343 = ~n56592 & n56625;
  assign n27344 = ~n27206 & ~n27343;
  assign n27345 = ~n27342 & ~n27343;
  assign n27346 = ~n27206 & n27345;
  assign n27347 = ~n27342 & n27344;
  assign n27348 = ~n27206 & ~n56635;
  assign n27349 = ~n27063 & n27075;
  assign n27350 = n27063 & ~n27076;
  assign n27351 = n27063 & n27075;
  assign n27352 = ~n27075 & ~n27076;
  assign n27353 = ~n27063 & ~n27075;
  assign n27354 = ~n56636 & ~n56637;
  assign n27355 = ~n27076 & ~n27349;
  assign n27356 = ~n27348 & ~n56638;
  assign n27357 = ~n27076 & ~n27356;
  assign n27358 = ~n26886 & n56602;
  assign n27359 = ~n26902 & ~n27358;
  assign n27360 = ~n27357 & n27359;
  assign n27361 = n27357 & ~n27359;
  assign n27362 = ~n27360 & ~n27361;
  assign n27363 = n26495 & ~n26497;
  assign n27364 = ~n26495 & ~n56559;
  assign n27365 = ~n26496 & n26501;
  assign n27366 = ~n27364 & ~n27365;
  assign n27367 = ~n56559 & ~n27363;
  assign n27368 = n11279 & ~n56639;
  assign n27369 = n12584 & n26259;
  assign n27370 = n54410 & n26265;
  assign n27371 = n11267 & n26262;
  assign n27372 = ~n27370 & ~n27371;
  assign n27373 = ~n27369 & n27372;
  assign n27374 = ~n11279 & n27373;
  assign n27375 = n56639 & n27373;
  assign n27376 = ~n27374 & ~n27375;
  assign n27377 = ~n27368 & n27373;
  assign n27378 = pi29  & ~n56640;
  assign n27379 = ~pi29  & n56640;
  assign n27380 = ~n27378 & ~n27379;
  assign n27381 = n27362 & ~n27380;
  assign n27382 = ~n27360 & ~n27381;
  assign n27383 = n27061 & ~n27382;
  assign n27384 = ~n27061 & n27382;
  assign n27385 = ~n27383 & ~n27384;
  assign n27386 = n26501 & ~n26503;
  assign n27387 = ~n26504 & ~n27386;
  assign n27388 = n11279 & n27387;
  assign n27389 = n12584 & n26256;
  assign n27390 = n54410 & n26262;
  assign n27391 = n11267 & n26259;
  assign n27392 = ~n27390 & ~n27391;
  assign n27393 = ~n27389 & n27392;
  assign n27394 = ~n27388 & n27393;
  assign n27395 = pi29  & ~n27394;
  assign n27396 = pi29  & ~n27395;
  assign n27397 = pi29  & n27394;
  assign n27398 = ~n27394 & ~n27395;
  assign n27399 = ~pi29  & ~n27394;
  assign n27400 = ~n56641 & ~n56642;
  assign n27401 = n27385 & ~n27400;
  assign n27402 = ~n27385 & n27400;
  assign n27403 = n27385 & ~n27401;
  assign n27404 = n27385 & n27400;
  assign n27405 = ~n27400 & ~n27401;
  assign n27406 = ~n27385 & ~n27400;
  assign n27407 = ~n56643 & ~n56644;
  assign n27408 = ~n27401 & ~n27402;
  assign n27409 = ~n26575 & ~n56645;
  assign n27410 = n26575 & n56645;
  assign n27411 = ~n56645 & ~n27409;
  assign n27412 = ~n26575 & ~n27409;
  assign n27413 = ~n27411 & ~n27412;
  assign n27414 = ~n27409 & ~n27410;
  assign n27415 = ~n27362 & n27380;
  assign n27416 = ~n27381 & ~n27415;
  assign n27417 = n27342 & ~n27344;
  assign n27418 = ~n27342 & ~n56635;
  assign n27419 = ~n27343 & n27348;
  assign n27420 = ~n27418 & ~n27419;
  assign n27421 = ~n56635 & ~n27417;
  assign n27422 = n26469 & ~n26471;
  assign n27423 = ~n26469 & ~n56556;
  assign n27424 = ~n26470 & n26475;
  assign n27425 = ~n27423 & ~n27424;
  assign n27426 = ~n56556 & ~n27422;
  assign n27427 = n1576 & ~n56648;
  assign n27428 = n11215 & n26274;
  assign n27429 = n54403 & n26280;
  assign n27430 = n10564 & n26277;
  assign n27431 = ~n27429 & ~n27430;
  assign n27432 = ~n27428 & n27431;
  assign n27433 = ~n27427 & n27432;
  assign n27434 = ~n56647 & ~n27433;
  assign n27435 = n11279 & n27042;
  assign n27436 = n12584 & n26265;
  assign n27437 = n54410 & n26271;
  assign n27438 = n11267 & n26268;
  assign n27439 = ~n27437 & ~n27438;
  assign n27440 = ~n27436 & n27439;
  assign n27441 = ~n11279 & n27440;
  assign n27442 = ~n27042 & n27440;
  assign n27443 = ~n27441 & ~n27442;
  assign n27444 = ~n27435 & n27440;
  assign n27445 = pi29  & ~n56649;
  assign n27446 = ~pi29  & n56649;
  assign n27447 = ~n27445 & ~n27446;
  assign n27448 = n56647 & n27433;
  assign n27449 = ~n56647 & ~n27434;
  assign n27450 = ~n56647 & n27433;
  assign n27451 = ~n27433 & ~n27434;
  assign n27452 = n56647 & ~n27433;
  assign n27453 = ~n56650 & ~n56651;
  assign n27454 = ~n27434 & ~n27448;
  assign n27455 = ~n27447 & ~n56652;
  assign n27456 = ~n27434 & ~n27455;
  assign n27457 = n27348 & n56638;
  assign n27458 = ~n56638 & ~n27356;
  assign n27459 = n27348 & ~n56638;
  assign n27460 = ~n27348 & ~n27356;
  assign n27461 = ~n27348 & n56638;
  assign n27462 = ~n56653 & ~n56654;
  assign n27463 = ~n27356 & ~n27457;
  assign n27464 = ~n27456 & ~n56655;
  assign n27465 = n26491 & ~n26493;
  assign n27466 = ~n26494 & ~n27465;
  assign n27467 = n11279 & n27466;
  assign n27468 = n12584 & n26262;
  assign n27469 = n54410 & n26268;
  assign n27470 = n11267 & n26265;
  assign n27471 = ~n27469 & ~n27470;
  assign n27472 = ~n27468 & n27471;
  assign n27473 = ~n27467 & n27472;
  assign n27474 = pi29  & ~n27473;
  assign n27475 = pi29  & ~n27474;
  assign n27476 = pi29  & n27473;
  assign n27477 = ~n27473 & ~n27474;
  assign n27478 = ~pi29  & ~n27473;
  assign n27479 = ~n56656 & ~n56657;
  assign n27480 = n27456 & n56655;
  assign n27481 = ~n27479 & ~n27480;
  assign n27482 = ~n27456 & ~n27464;
  assign n27483 = ~n56655 & ~n27464;
  assign n27484 = ~n27482 & ~n27483;
  assign n27485 = ~n27464 & ~n27480;
  assign n27486 = ~n27479 & ~n56658;
  assign n27487 = ~n27464 & ~n27486;
  assign n27488 = ~n27464 & ~n27481;
  assign n27489 = n27416 & ~n56659;
  assign n27490 = n26511 & ~n26513;
  assign n27491 = ~n26514 & ~n27490;
  assign n27492 = n123 & n27491;
  assign n27493 = n128 & n26250;
  assign n27494 = n53444 & n26256;
  assign n27495 = n127 & n26253;
  assign n27496 = ~n27494 & ~n27495;
  assign n27497 = ~n27493 & n27496;
  assign n27498 = ~n27492 & n27497;
  assign n27499 = pi26  & ~n27498;
  assign n27500 = pi26  & ~n27499;
  assign n27501 = pi26  & n27498;
  assign n27502 = ~n27498 & ~n27499;
  assign n27503 = ~pi26  & ~n27498;
  assign n27504 = ~n56660 & ~n56661;
  assign n27505 = ~n27416 & n56659;
  assign n27506 = ~n27504 & ~n27505;
  assign n27507 = ~n27489 & ~n27505;
  assign n27508 = ~n27504 & n27507;
  assign n27509 = ~n27489 & ~n27508;
  assign n27510 = ~n27489 & ~n27506;
  assign n27511 = ~n56646 & ~n56662;
  assign n27512 = n56646 & n56662;
  assign n27513 = ~n27511 & ~n27512;
  assign n27514 = ~n26557 & n27513;
  assign n27515 = ~n26557 & ~n27514;
  assign n27516 = ~n26557 & ~n27513;
  assign n27517 = n27513 & ~n27514;
  assign n27518 = n26557 & n27513;
  assign n27519 = n26557 & ~n27513;
  assign n27520 = ~n27514 & ~n27519;
  assign n27521 = ~n56663 & ~n56664;
  assign n27522 = ~n15901 & ~n15921;
  assign n27523 = ~n14407 & ~n14413;
  assign n27524 = ~n54719 & n56666;
  assign n27525 = ~n14413 & n27524;
  assign n27526 = ~n54719 & ~n14413;
  assign n27527 = n56666 & n27526;
  assign n27528 = ~n54716 & n14407;
  assign n27529 = pi20  & n56667;
  assign n27530 = ~pi20  & ~n56667;
  assign n27531 = ~n27529 & ~n27530;
  assign n27532 = n26505 & ~n26507;
  assign n27533 = ~n26505 & ~n56560;
  assign n27534 = ~n26506 & n26511;
  assign n27535 = ~n27533 & ~n27534;
  assign n27536 = ~n56560 & ~n27532;
  assign n27537 = n123 & ~n56668;
  assign n27538 = n128 & n26253;
  assign n27539 = n53444 & n26259;
  assign n27540 = n127 & n26256;
  assign n27541 = ~n27539 & ~n27540;
  assign n27542 = ~n27538 & n27541;
  assign n27543 = ~n27537 & n27542;
  assign n27544 = pi26  & ~n27543;
  assign n27545 = pi26  & ~n27544;
  assign n27546 = pi26  & n27543;
  assign n27547 = ~n27543 & ~n27544;
  assign n27548 = ~pi26  & ~n27543;
  assign n27549 = ~n56669 & ~n56670;
  assign n27550 = ~n27479 & ~n27486;
  assign n27551 = ~n27479 & n56658;
  assign n27552 = ~n56658 & ~n27486;
  assign n27553 = n27479 & ~n56658;
  assign n27554 = n27479 & n56658;
  assign n27555 = ~n27486 & ~n27554;
  assign n27556 = ~n56671 & ~n56672;
  assign n27557 = ~n27549 & n56673;
  assign n27558 = n27549 & ~n56673;
  assign n27559 = n56673 & ~n27557;
  assign n27560 = n27549 & n56673;
  assign n27561 = ~n27549 & ~n27557;
  assign n27562 = ~n27549 & ~n56673;
  assign n27563 = ~n56674 & ~n56675;
  assign n27564 = ~n27557 & ~n27558;
  assign n27565 = ~n27328 & n56634;
  assign n27566 = ~n27341 & ~n27565;
  assign n27567 = n53771 & n5749;
  assign n27568 = n1712 & n2340;
  assign n27569 = n54372 & n27568;
  assign n27570 = n27567 & n27569;
  assign n27571 = ~n168 & ~n349;
  assign n27572 = ~n440 & ~n498;
  assign n27573 = ~n168 & ~n498;
  assign n27574 = ~n349 & ~n440;
  assign n27575 = n27573 & n27574;
  assign n27576 = n27571 & n27572;
  assign n27577 = ~n168 & ~n1634;
  assign n27578 = ~n1641 & n27577;
  assign n27579 = ~n498 & n27578;
  assign n27580 = ~n440 & n27579;
  assign n27581 = ~n349 & n27580;
  assign n27582 = ~n440 & ~n1634;
  assign n27583 = ~n349 & ~n1641;
  assign n27584 = n27582 & n27583;
  assign n27585 = n27573 & n27584;
  assign n27586 = n5587 & n56677;
  assign n27587 = n1078 & n5378;
  assign n27588 = n2175 & n27587;
  assign n27589 = ~n249 & ~n585;
  assign n27590 = n3639 & n27589;
  assign n27591 = n53673 & n27590;
  assign n27592 = n27588 & n27591;
  assign n27593 = n56678 & n27592;
  assign n27594 = n54372 & n27567;
  assign n27595 = n56678 & n27594;
  assign n27596 = n3639 & n27595;
  assign n27597 = n1712 & n27596;
  assign n27598 = n5378 & n27597;
  assign n27599 = n1078 & n27598;
  assign n27600 = n53673 & n27599;
  assign n27601 = n2340 & n27600;
  assign n27602 = ~n922 & n27601;
  assign n27603 = ~n249 & n27602;
  assign n27604 = ~n409 & n27603;
  assign n27605 = ~n585 & n27604;
  assign n27606 = n53673 & n53771;
  assign n27607 = n5749 & n27568;
  assign n27608 = n27606 & n27607;
  assign n27609 = n54372 & n27590;
  assign n27610 = n27588 & n27609;
  assign n27611 = n56678 & n27610;
  assign n27612 = n27608 & n27611;
  assign n27613 = n53673 & n5749;
  assign n27614 = n53771 & n54372;
  assign n27615 = n27613 & n27614;
  assign n27616 = n3639 & n27587;
  assign n27617 = ~n249 & ~n409;
  assign n27618 = ~n585 & ~n922;
  assign n27619 = n27617 & n27618;
  assign n27620 = n27568 & n27619;
  assign n27621 = n27616 & n27620;
  assign n27622 = n56678 & n27621;
  assign n27623 = n27615 & n27622;
  assign n27624 = n27570 & n27593;
  assign n27625 = n1035 & n1541;
  assign n27626 = n4538 & n27625;
  assign n27627 = n54232 & n27626;
  assign n27628 = n54436 & n27627;
  assign n27629 = n1267 & n1709;
  assign n27630 = n5485 & n7646;
  assign n27631 = n1709 & n7646;
  assign n27632 = n1267 & n5485;
  assign n27633 = n27631 & n27632;
  assign n27634 = n27629 & n27630;
  assign n27635 = ~n617 & ~n628;
  assign n27636 = ~n495 & ~n894;
  assign n27637 = ~n495 & ~n617;
  assign n27638 = ~n628 & ~n894;
  assign n27639 = n27637 & n27638;
  assign n27640 = ~n617 & ~n894;
  assign n27641 = ~n495 & ~n628;
  assign n27642 = n27640 & n27641;
  assign n27643 = n27635 & n27636;
  assign n27644 = n54497 & n56681;
  assign n27645 = n1709 & n54497;
  assign n27646 = n1267 & n27645;
  assign n27647 = n5485 & n27646;
  assign n27648 = n7646 & n27647;
  assign n27649 = ~n628 & n27648;
  assign n27650 = ~n894 & n27649;
  assign n27651 = ~n495 & n27650;
  assign n27652 = ~n617 & n27651;
  assign n27653 = n56680 & n27644;
  assign n27654 = ~n735 & ~n914;
  assign n27655 = ~n1125 & ~n1535;
  assign n27656 = n27654 & n27655;
  assign n27657 = ~n184 & ~n401;
  assign n27658 = ~n364 & ~n419;
  assign n27659 = ~n184 & ~n364;
  assign n27660 = ~n401 & ~n419;
  assign n27661 = n27659 & n27660;
  assign n27662 = n27657 & n27658;
  assign n27663 = n27656 & n56683;
  assign n27664 = n3776 & n13164;
  assign n27665 = n53836 & n27664;
  assign n27666 = n27663 & n27665;
  assign n27667 = n56682 & n27666;
  assign n27668 = n1541 & n4538;
  assign n27669 = n13164 & n27668;
  assign n27670 = n54232 & n27669;
  assign n27671 = n54436 & n27670;
  assign n27672 = ~n184 & ~n419;
  assign n27673 = n27655 & n27672;
  assign n27674 = n1035 & n3776;
  assign n27675 = n27673 & n27674;
  assign n27676 = ~n364 & ~n401;
  assign n27677 = n27654 & n27676;
  assign n27678 = n53836 & n27677;
  assign n27679 = n27675 & n27678;
  assign n27680 = n56682 & n27679;
  assign n27681 = n27671 & n27680;
  assign n27682 = n1541 & n3776;
  assign n27683 = n13164 & n27682;
  assign n27684 = n54232 & n27683;
  assign n27685 = n54436 & n27684;
  assign n27686 = ~n364 & ~n1125;
  assign n27687 = ~n401 & ~n1535;
  assign n27688 = n27686 & n27687;
  assign n27689 = n1035 & n4538;
  assign n27690 = n27688 & n27689;
  assign n27691 = ~n419 & ~n735;
  assign n27692 = ~n184 & ~n914;
  assign n27693 = n27691 & n27692;
  assign n27694 = n53836 & n27693;
  assign n27695 = n27690 & n27694;
  assign n27696 = n56682 & n27695;
  assign n27697 = n27685 & n27696;
  assign n27698 = n27628 & n27667;
  assign n27699 = n54182 & n56684;
  assign n27700 = n53836 & n56682;
  assign n27701 = n54436 & n27700;
  assign n27702 = n54232 & n27701;
  assign n27703 = n56679 & n27702;
  assign n27704 = n1541 & n27703;
  assign n27705 = n4538 & n27704;
  assign n27706 = n1035 & n27705;
  assign n27707 = n54182 & n27706;
  assign n27708 = n13164 & n27707;
  assign n27709 = n3776 & n27708;
  assign n27710 = ~n1125 & n27709;
  assign n27711 = ~n184 & n27710;
  assign n27712 = ~n401 & n27711;
  assign n27713 = ~n1535 & n27712;
  assign n27714 = ~n914 & n27713;
  assign n27715 = ~n419 & n27714;
  assign n27716 = ~n364 & n27715;
  assign n27717 = ~n735 & n27716;
  assign n27718 = n56679 & n27699;
  assign n27719 = n56628 & ~n56685;
  assign n27720 = ~n56628 & n56685;
  assign n27721 = ~n27719 & ~n27720;
  assign n27722 = n26455 & ~n26457;
  assign n27723 = ~n26455 & ~n56555;
  assign n27724 = ~n26456 & n26461;
  assign n27725 = ~n27723 & ~n27724;
  assign n27726 = ~n56555 & ~n27722;
  assign n27727 = n1576 & ~n56686;
  assign n27728 = n11215 & n26283;
  assign n27729 = n54403 & n26289;
  assign n27730 = n10564 & n26286;
  assign n27731 = ~n27729 & ~n27730;
  assign n27732 = ~n27728 & n27731;
  assign n27733 = ~n27727 & n27732;
  assign n27734 = ~n27719 & ~n27733;
  assign n27735 = ~n27720 & n27734;
  assign n27736 = n27721 & ~n27733;
  assign n27737 = ~n27719 & ~n56687;
  assign n27738 = ~n27321 & ~n27323;
  assign n27739 = ~n27324 & ~n27738;
  assign n27740 = ~n27737 & n27739;
  assign n27741 = n27737 & ~n27739;
  assign n27742 = n26461 & ~n26463;
  assign n27743 = ~n26464 & ~n27742;
  assign n27744 = n1576 & n27743;
  assign n27745 = n11215 & n26280;
  assign n27746 = n54403 & n26286;
  assign n27747 = n10564 & n26283;
  assign n27748 = ~n27746 & ~n27747;
  assign n27749 = ~n27745 & n27748;
  assign n27750 = ~n27744 & n27749;
  assign n27751 = ~n27741 & ~n27750;
  assign n27752 = ~n27740 & ~n27741;
  assign n27753 = ~n27750 & n27752;
  assign n27754 = ~n27740 & ~n27753;
  assign n27755 = ~n27740 & ~n27751;
  assign n27756 = n27566 & ~n56688;
  assign n27757 = ~n27566 & n56688;
  assign n27758 = ~n27756 & ~n27757;
  assign n27759 = n11279 & ~n56601;
  assign n27760 = n12584 & n26268;
  assign n27761 = n54410 & n26274;
  assign n27762 = n11267 & n26271;
  assign n27763 = ~n27761 & ~n27762;
  assign n27764 = ~n27760 & n27763;
  assign n27765 = ~n11279 & n27764;
  assign n27766 = n56601 & n27764;
  assign n27767 = ~n27765 & ~n27766;
  assign n27768 = ~n27759 & n27764;
  assign n27769 = pi29  & ~n56689;
  assign n27770 = ~pi29  & n56689;
  assign n27771 = ~n27769 & ~n27770;
  assign n27772 = n27758 & ~n27771;
  assign n27773 = ~n27756 & ~n27772;
  assign n27774 = n27447 & n56652;
  assign n27775 = ~n27455 & ~n27774;
  assign n27776 = ~n27773 & n27775;
  assign n27777 = n27773 & ~n27775;
  assign n27778 = n123 & n27387;
  assign n27779 = n128 & n26256;
  assign n27780 = n53444 & n26262;
  assign n27781 = n127 & n26259;
  assign n27782 = ~n27780 & ~n27781;
  assign n27783 = ~n27779 & n27782;
  assign n27784 = ~n27778 & n27783;
  assign n27785 = pi26  & ~n27784;
  assign n27786 = pi26  & ~n27785;
  assign n27787 = pi26  & n27784;
  assign n27788 = ~n27784 & ~n27785;
  assign n27789 = ~pi26  & ~n27784;
  assign n27790 = ~n56690 & ~n56691;
  assign n27791 = ~n27777 & ~n27790;
  assign n27792 = ~n27776 & ~n27777;
  assign n27793 = ~n27790 & n27792;
  assign n27794 = ~n27776 & ~n27793;
  assign n27795 = ~n27776 & ~n27791;
  assign n27796 = ~n56676 & ~n56692;
  assign n27797 = ~n27557 & ~n27796;
  assign n27798 = ~n27504 & ~n27508;
  assign n27799 = ~n27504 & ~n27507;
  assign n27800 = n27507 & ~n27508;
  assign n27801 = n27504 & n27507;
  assign n27802 = n27504 & ~n27507;
  assign n27803 = ~n27508 & ~n27802;
  assign n27804 = ~n56693 & ~n56694;
  assign n27805 = ~n27797 & n56695;
  assign n27806 = n27797 & ~n56695;
  assign n27807 = n26525 & ~n26527;
  assign n27808 = ~n26528 & ~n27807;
  assign n27809 = n90 & n27808;
  assign n27810 = n14236 & n26242;
  assign n27811 = n54667 & n26247;
  assign n27812 = n14210 & n26244;
  assign n27813 = ~n27811 & ~n27812;
  assign n27814 = ~n27810 & n27813;
  assign n27815 = ~n27809 & n27814;
  assign n27816 = pi23  & ~n27815;
  assign n27817 = pi23  & ~n27816;
  assign n27818 = pi23  & n27815;
  assign n27819 = ~n27815 & ~n27816;
  assign n27820 = ~pi23  & ~n27815;
  assign n27821 = ~n56696 & ~n56697;
  assign n27822 = ~n27806 & ~n27821;
  assign n27823 = ~n27805 & ~n27806;
  assign n27824 = ~n27821 & n27823;
  assign n27825 = ~n27805 & ~n27824;
  assign n27826 = ~n27805 & ~n27822;
  assign n27827 = ~n27531 & ~n56698;
  assign n27828 = n27531 & n56698;
  assign n27829 = ~n27827 & ~n27828;
  assign n27830 = n56665 & n27829;
  assign n27831 = ~n56665 & ~n27829;
  assign n27832 = n56665 & ~n27830;
  assign n27833 = n27829 & ~n27830;
  assign n27834 = ~n27832 & ~n27833;
  assign n27835 = ~n27830 & ~n27831;
  assign n27836 = n56676 & n56692;
  assign n27837 = ~n27796 & ~n27836;
  assign n27838 = n26521 & ~n26523;
  assign n27839 = ~n26524 & ~n27838;
  assign n27840 = n90 & n27839;
  assign n27841 = n14236 & n26244;
  assign n27842 = n54667 & n26250;
  assign n27843 = n14210 & n26247;
  assign n27844 = ~n27842 & ~n27843;
  assign n27845 = ~n27841 & n27844;
  assign n27846 = ~n27840 & n27845;
  assign n27847 = pi23  & ~n27846;
  assign n27848 = pi23  & ~n27847;
  assign n27849 = pi23  & n27846;
  assign n27850 = ~n27846 & ~n27847;
  assign n27851 = ~pi23  & ~n27846;
  assign n27852 = ~n56700 & ~n56701;
  assign n27853 = n27837 & ~n27852;
  assign n27854 = ~n27837 & n27852;
  assign n27855 = n27837 & ~n27853;
  assign n27856 = n27837 & n27852;
  assign n27857 = ~n27852 & ~n27853;
  assign n27858 = ~n27837 & ~n27852;
  assign n27859 = ~n56702 & ~n56703;
  assign n27860 = ~n27853 & ~n27854;
  assign n27861 = n27790 & ~n27792;
  assign n27862 = n27792 & ~n27793;
  assign n27863 = ~n27790 & ~n27793;
  assign n27864 = ~n27862 & ~n27863;
  assign n27865 = ~n27793 & ~n27861;
  assign n27866 = n11279 & ~n56612;
  assign n27867 = n12584 & n26271;
  assign n27868 = n54410 & n26277;
  assign n27869 = n11267 & n26274;
  assign n27870 = ~n27868 & ~n27869;
  assign n27871 = ~n27867 & n27870;
  assign n27872 = ~n27866 & n27871;
  assign n27873 = pi29  & ~n27872;
  assign n27874 = pi29  & ~n27873;
  assign n27875 = pi29  & n27872;
  assign n27876 = ~n27872 & ~n27873;
  assign n27877 = ~pi29  & ~n27872;
  assign n27878 = ~n56706 & ~n56707;
  assign n27879 = n27750 & ~n27752;
  assign n27880 = n27752 & ~n27753;
  assign n27881 = ~n27750 & ~n27753;
  assign n27882 = ~n27880 & ~n27881;
  assign n27883 = ~n27753 & ~n27879;
  assign n27884 = ~n27878 & ~n56708;
  assign n27885 = ~n249 & ~n356;
  assign n27886 = ~n1455 & n27885;
  assign n27887 = ~n733 & ~n1079;
  assign n27888 = n1683 & n27887;
  assign n27889 = ~n1079 & n1456;
  assign n27890 = ~n141 & n27889;
  assign n27891 = ~n249 & n27890;
  assign n27892 = ~n748 & n27891;
  assign n27893 = ~n356 & n27892;
  assign n27894 = ~n1079 & n27885;
  assign n27895 = n1456 & n1683;
  assign n27896 = n27894 & n27895;
  assign n27897 = ~n1079 & n1683;
  assign n27898 = n1456 & n27885;
  assign n27899 = n27897 & n27898;
  assign n27900 = n27886 & n27888;
  assign n27901 = ~n647 & ~n650;
  assign n27902 = n462 & n27901;
  assign n27903 = n424 & n13597;
  assign n27904 = n27902 & n27903;
  assign n27905 = n54601 & n27904;
  assign n27906 = n56709 & n27905;
  assign n27907 = ~n268 & ~n663;
  assign n27908 = n2537 & n27907;
  assign n27909 = n7016 & n14605;
  assign n27910 = n27908 & n27909;
  assign n27911 = ~n108 & ~n182;
  assign n27912 = ~n401 & ~n984;
  assign n27913 = n27911 & n27912;
  assign n27914 = n53977 & n27913;
  assign n27915 = n53977 & n7016;
  assign n27916 = n2537 & n27915;
  assign n27917 = ~n984 & n27916;
  assign n27918 = ~n2103 & n27917;
  assign n27919 = ~n108 & n27918;
  assign n27920 = ~n182 & n27919;
  assign n27921 = ~n663 & n27920;
  assign n27922 = ~n401 & n27921;
  assign n27923 = ~n975 & n27922;
  assign n27924 = ~n268 & n27923;
  assign n27925 = ~n401 & ~n663;
  assign n27926 = n2537 & n27925;
  assign n27927 = n27909 & n27926;
  assign n27928 = ~n268 & ~n984;
  assign n27929 = n27911 & n27928;
  assign n27930 = n53977 & n27929;
  assign n27931 = n27927 & n27930;
  assign n27932 = ~n182 & ~n401;
  assign n27933 = n27928 & n27932;
  assign n27934 = n2537 & n7016;
  assign n27935 = n27933 & n27934;
  assign n27936 = ~n108 & ~n975;
  assign n27937 = ~n663 & ~n2103;
  assign n27938 = n27936 & n27937;
  assign n27939 = n53977 & n27938;
  assign n27940 = n27935 & n27939;
  assign n27941 = n27910 & n27914;
  assign n27942 = ~n316 & ~n410;
  assign n27943 = ~n491 & ~n977;
  assign n27944 = ~n316 & ~n491;
  assign n27945 = ~n410 & ~n977;
  assign n27946 = n27944 & n27945;
  assign n27947 = n27942 & n27943;
  assign n27948 = n54156 & n56711;
  assign n27949 = n164 & n3639;
  assign n27950 = n53512 & n27949;
  assign n27951 = n27948 & n27950;
  assign n27952 = n56710 & n27951;
  assign n27953 = ~n491 & ~n647;
  assign n27954 = n462 & n27953;
  assign n27955 = n27903 & n27954;
  assign n27956 = n54601 & n27955;
  assign n27957 = n56709 & n27956;
  assign n27958 = ~n316 & ~n650;
  assign n27959 = n27945 & n27958;
  assign n27960 = n54156 & n27959;
  assign n27961 = n27950 & n27960;
  assign n27962 = n56710 & n27961;
  assign n27963 = n27957 & n27962;
  assign n27964 = n27903 & n27949;
  assign n27965 = n54601 & n27964;
  assign n27966 = n56709 & n27965;
  assign n27967 = n53512 & n54156;
  assign n27968 = ~n316 & ~n977;
  assign n27969 = ~n410 & ~n647;
  assign n27970 = n27968 & n27969;
  assign n27971 = ~n491 & ~n650;
  assign n27972 = n462 & n27971;
  assign n27973 = n27970 & n27972;
  assign n27974 = n27967 & n27973;
  assign n27975 = n56710 & n27974;
  assign n27976 = n27966 & n27975;
  assign n27977 = n424 & n462;
  assign n27978 = n27949 & n27977;
  assign n27979 = n54601 & n27978;
  assign n27980 = n56709 & n27979;
  assign n27981 = n13597 & n27901;
  assign n27982 = n56711 & n27981;
  assign n27983 = n27967 & n27982;
  assign n27984 = n56710 & n27983;
  assign n27985 = n27980 & n27984;
  assign n27986 = n27906 & n27952;
  assign n27987 = n54318 & n56712;
  assign n27988 = n54601 & n27967;
  assign n27989 = n3639 & n27988;
  assign n27990 = n56709 & n27989;
  assign n27991 = n54318 & n27990;
  assign n27992 = n54999 & n27991;
  assign n27993 = n56710 & n27992;
  assign n27994 = n424 & n27993;
  assign n27995 = n462 & n27994;
  assign n27996 = n164 & n27995;
  assign n27997 = ~n316 & n27996;
  assign n27998 = ~n977 & n27997;
  assign n27999 = n13597 & n27998;
  assign n28000 = ~n491 & n27999;
  assign n28001 = ~n647 & n28000;
  assign n28002 = ~n410 & n28001;
  assign n28003 = ~n650 & n28002;
  assign n28004 = n54999 & n27987;
  assign n28005 = n53814 & n53934;
  assign n28006 = n54933 & n28005;
  assign n28007 = ~n506 & ~n659;
  assign n28008 = ~n770 & n8824;
  assign n28009 = ~n770 & n28007;
  assign n28010 = n8824 & n28009;
  assign n28011 = n28007 & n28008;
  assign n28012 = n5848 & n8824;
  assign n28013 = ~n659 & n28012;
  assign n28014 = ~n506 & n28013;
  assign n28015 = ~n770 & n28014;
  assign n28016 = n5848 & n56714;
  assign n28017 = n53760 & n54215;
  assign n28018 = n13598 & n28017;
  assign n28019 = ~n256 & ~n402;
  assign n28020 = n897 & n5390;
  assign n28021 = n28019 & n28020;
  assign n28022 = ~n824 & ~n1472;
  assign n28023 = n472 & n28022;
  assign n28024 = n2628 & n28023;
  assign n28025 = n472 & n897;
  assign n28026 = n28019 & n28025;
  assign n28027 = n5390 & n28022;
  assign n28028 = n2628 & n28027;
  assign n28029 = n28026 & n28028;
  assign n28030 = n472 & n5390;
  assign n28031 = n28019 & n28030;
  assign n28032 = n897 & n28022;
  assign n28033 = n2628 & n28032;
  assign n28034 = n28031 & n28033;
  assign n28035 = n28021 & n28024;
  assign n28036 = n2628 & n54215;
  assign n28037 = n53760 & n28036;
  assign n28038 = n897 & n28030;
  assign n28039 = n28019 & n28022;
  assign n28040 = n13598 & n28039;
  assign n28041 = n28038 & n28040;
  assign n28042 = n28037 & n28041;
  assign n28043 = n28018 & n56716;
  assign n28044 = n56715 & n56717;
  assign n28045 = n53693 & n28044;
  assign n28046 = n897 & n28036;
  assign n28047 = n472 & n28046;
  assign n28048 = n54933 & n28047;
  assign n28049 = n53934 & n28048;
  assign n28050 = n53814 & n28049;
  assign n28051 = n53693 & n28050;
  assign n28052 = n53760 & n28051;
  assign n28053 = n56715 & n28052;
  assign n28054 = n5390 & n28053;
  assign n28055 = n13598 & n28054;
  assign n28056 = ~n1472 & n28055;
  assign n28057 = ~n256 & n28056;
  assign n28058 = ~n402 & n28057;
  assign n28059 = ~n824 & n28058;
  assign n28060 = n28006 & n28045;
  assign n28061 = ~n56713 & ~n56718;
  assign n28062 = ~n19509 & ~n19541;
  assign n28063 = ~n18834 & ~n18846;
  assign n28064 = ~n55247 & ~n18846;
  assign n28065 = n56719 & n28064;
  assign n28066 = ~n55247 & n56719;
  assign n28067 = ~n18846 & n28066;
  assign n28068 = n18834 & ~n55246;
  assign n28069 = pi11  & n56720;
  assign n28070 = ~pi11  & ~n56720;
  assign n28071 = ~n28069 & ~n28070;
  assign n28072 = n56713 & n56718;
  assign n28073 = ~n28061 & ~n28072;
  assign n28074 = n28071 & n28073;
  assign n28075 = ~n28061 & ~n28074;
  assign n28076 = n56628 & ~n28075;
  assign n28077 = ~n56628 & n28075;
  assign n28078 = ~n28076 & ~n28077;
  assign n28079 = n26449 & ~n26451;
  assign n28080 = ~n26449 & ~n56554;
  assign n28081 = ~n26450 & n26455;
  assign n28082 = ~n28080 & ~n28081;
  assign n28083 = ~n56554 & ~n28079;
  assign n28084 = n1576 & ~n56721;
  assign n28085 = n11215 & n26286;
  assign n28086 = n10564 & n26289;
  assign n28087 = n54403 & n26292;
  assign n28088 = ~n28086 & ~n28087;
  assign n28089 = ~n28085 & n28088;
  assign n28090 = ~n28084 & ~n28087;
  assign n28091 = ~n28086 & n28090;
  assign n28092 = ~n28085 & n28091;
  assign n28093 = ~n28084 & n28089;
  assign n28094 = n28078 & ~n56722;
  assign n28095 = ~n28076 & ~n28094;
  assign n28096 = ~n27721 & n27733;
  assign n28097 = ~n27733 & ~n56687;
  assign n28098 = ~n27720 & n27737;
  assign n28099 = ~n28097 & ~n28098;
  assign n28100 = ~n56687 & ~n28096;
  assign n28101 = ~n28095 & ~n56723;
  assign n28102 = n28095 & n56723;
  assign n28103 = ~n28101 & ~n28102;
  assign n28104 = ~n28071 & ~n28073;
  assign n28105 = ~n28074 & ~n28104;
  assign n28106 = n26445 & ~n26447;
  assign n28107 = ~n26448 & ~n28106;
  assign n28108 = n1576 & n28107;
  assign n28109 = n11215 & n26289;
  assign n28110 = n54403 & n26295;
  assign n28111 = n10564 & n26292;
  assign n28112 = ~n28110 & ~n28111;
  assign n28113 = ~n28109 & n28112;
  assign n28114 = ~n28108 & n28113;
  assign n28115 = n28105 & ~n28114;
  assign n28116 = ~n112 & ~n848;
  assign n28117 = ~n112 & ~n1059;
  assign n28118 = ~n848 & n28117;
  assign n28119 = ~n848 & ~n1059;
  assign n28120 = ~n112 & n28119;
  assign n28121 = ~n1059 & n28116;
  assign n28122 = ~n112 & n4584;
  assign n28123 = ~n1059 & n28122;
  assign n28124 = ~n848 & n28123;
  assign n28125 = n4584 & n56724;
  assign n28126 = n54303 & n54642;
  assign n28127 = n56725 & n28126;
  assign n28128 = ~n174 & ~n747;
  assign n28129 = ~n852 & ~n1881;
  assign n28130 = ~n174 & ~n852;
  assign n28131 = ~n747 & n28130;
  assign n28132 = ~n1881 & n28131;
  assign n28133 = ~n747 & ~n1881;
  assign n28134 = n28130 & n28133;
  assign n28135 = n28128 & n28129;
  assign n28136 = ~n770 & ~n1079;
  assign n28137 = ~n770 & ~n883;
  assign n28138 = ~n1079 & n28137;
  assign n28139 = ~n883 & n28136;
  assign n28140 = ~n415 & ~n741;
  assign n28141 = n1488 & n28140;
  assign n28142 = ~n415 & ~n883;
  assign n28143 = ~n1079 & n28142;
  assign n28144 = ~n741 & ~n770;
  assign n28145 = n1488 & n28144;
  assign n28146 = n28143 & n28145;
  assign n28147 = n56727 & n28141;
  assign n28148 = n56726 & n56728;
  assign n28149 = n3474 & n3536;
  assign n28150 = n1531 & n1803;
  assign n28151 = n28149 & n28150;
  assign n28152 = n53730 & n28151;
  assign n28153 = n28148 & n28152;
  assign n28154 = n54642 & n56726;
  assign n28155 = n56728 & n28154;
  assign n28156 = n54303 & n56725;
  assign n28157 = n28152 & n28156;
  assign n28158 = n28155 & n28157;
  assign n28159 = n355 & n28140;
  assign n28160 = n1488 & n3536;
  assign n28161 = n28159 & n28160;
  assign n28162 = n56726 & n56727;
  assign n28163 = n28161 & n28162;
  assign n28164 = n1803 & n3214;
  assign n28165 = n1531 & n3474;
  assign n28166 = n28164 & n28165;
  assign n28167 = n53730 & n28166;
  assign n28168 = n28156 & n28167;
  assign n28169 = n28163 & n28168;
  assign n28170 = n28127 & n28153;
  assign n28171 = n54303 & n28165;
  assign n28172 = n56725 & n28171;
  assign n28173 = n53730 & n28172;
  assign n28174 = n54136 & n28173;
  assign n28175 = n56726 & n28174;
  assign n28176 = n1488 & n28175;
  assign n28177 = n3214 & n28176;
  assign n28178 = n355 & n28177;
  assign n28179 = n1803 & n28178;
  assign n28180 = n3536 & n28179;
  assign n28181 = ~n883 & n28180;
  assign n28182 = ~n415 & n28181;
  assign n28183 = ~n1079 & n28182;
  assign n28184 = ~n741 & n28183;
  assign n28185 = ~n770 & n28184;
  assign n28186 = n54136 & n56729;
  assign n28187 = n14937 & n15061;
  assign n28188 = n26636 & n28187;
  assign n28189 = ~n663 & n846;
  assign n28190 = n2172 & n2477;
  assign n28191 = n28189 & n28190;
  assign n28192 = n846 & n2477;
  assign n28193 = n846 & n28190;
  assign n28194 = n2172 & n28192;
  assign n28195 = ~n902 & n56731;
  assign n28196 = ~n291 & n28195;
  assign n28197 = ~n295 & n28196;
  assign n28198 = ~n218 & n28197;
  assign n28199 = ~n663 & n28198;
  assign n28200 = ~n552 & n28199;
  assign n28201 = ~n617 & n28200;
  assign n28202 = n2172 & n14937;
  assign n28203 = n15061 & n28202;
  assign n28204 = ~n663 & n26636;
  assign n28205 = n28192 & n28204;
  assign n28206 = n28203 & n28205;
  assign n28207 = ~n663 & n15061;
  assign n28208 = n14937 & n26636;
  assign n28209 = n28207 & n28208;
  assign n28210 = n56731 & n28209;
  assign n28211 = n28188 & n28191;
  assign n28212 = ~n141 & ~n649;
  assign n28213 = ~n777 & ~n1703;
  assign n28214 = ~n649 & ~n1703;
  assign n28215 = ~n141 & ~n777;
  assign n28216 = n28214 & n28215;
  assign n28217 = n28212 & n28213;
  assign n28218 = n3370 & n56733;
  assign n28219 = n27568 & n28218;
  assign n28220 = n180 & n248;
  assign n28221 = n3165 & n11546;
  assign n28222 = n180 & n3165;
  assign n28223 = n248 & n11546;
  assign n28224 = n28222 & n28223;
  assign n28225 = n28220 & n28221;
  assign n28226 = n54070 & n56734;
  assign n28227 = n27568 & n28222;
  assign n28228 = ~n416 & ~n1703;
  assign n28229 = n248 & n28228;
  assign n28230 = n3370 & n28229;
  assign n28231 = ~n554 & ~n777;
  assign n28232 = n28212 & n28231;
  assign n28233 = n54070 & n28232;
  assign n28234 = n28230 & n28233;
  assign n28235 = n28227 & n28234;
  assign n28236 = n28219 & n28226;
  assign n28237 = n56732 & n56735;
  assign n28238 = n54614 & n28237;
  assign n28239 = n3165 & n54070;
  assign n28240 = n248 & n28239;
  assign n28241 = n3369 & n28240;
  assign n28242 = n56730 & n28241;
  assign n28243 = n54614 & n28242;
  assign n28244 = n56732 & n28243;
  assign n28245 = n1712 & n28244;
  assign n28246 = n180 & n28245;
  assign n28247 = n2476 & n28246;
  assign n28248 = n2340 & n28247;
  assign n28249 = ~n416 & n28248;
  assign n28250 = ~n1703 & n28249;
  assign n28251 = ~n141 & n28250;
  assign n28252 = ~n554 & n28251;
  assign n28253 = ~n649 & n28252;
  assign n28254 = ~n777 & n28253;
  assign n28255 = n56730 & n28238;
  assign n28256 = n56713 & ~n56736;
  assign n28257 = n1265 & n3950;
  assign n28258 = n8196 & n28257;
  assign n28259 = ~n179 & ~n770;
  assign n28260 = ~n770 & ~n1033;
  assign n28261 = ~n179 & n28260;
  assign n28262 = ~n1033 & n28259;
  assign n28263 = n749 & n2340;
  assign n28264 = n56737 & n28263;
  assign n28265 = n8196 & n28263;
  assign n28266 = n28257 & n56737;
  assign n28267 = n28265 & n28266;
  assign n28268 = n28258 & n28264;
  assign n28269 = n54493 & n56738;
  assign n28270 = n613 & n3670;
  assign n28271 = n1818 & n3670;
  assign n28272 = n613 & n28271;
  assign n28273 = n1818 & n28270;
  assign n28274 = ~n294 & ~n830;
  assign n28275 = ~n294 & n1659;
  assign n28276 = ~n830 & n28275;
  assign n28277 = n1659 & n28274;
  assign n28278 = ~n108 & ~n211;
  assign n28279 = ~n211 & ~n1881;
  assign n28280 = ~n108 & n28279;
  assign n28281 = ~n1881 & n28278;
  assign n28282 = n56740 & n56741;
  assign n28283 = n613 & n56740;
  assign n28284 = n3670 & n28283;
  assign n28285 = ~n108 & n28284;
  assign n28286 = ~n211 & n28285;
  assign n28287 = ~n617 & n28286;
  assign n28288 = ~n450 & n28287;
  assign n28289 = ~n1881 & n28288;
  assign n28290 = n56739 & n28282;
  assign n28291 = n53753 & n53797;
  assign n28292 = n53753 & n9331;
  assign n28293 = n53797 & n28292;
  assign n28294 = n53797 & n9331;
  assign n28295 = n53753 & n28294;
  assign n28296 = n9331 & n28291;
  assign n28297 = n56742 & n56743;
  assign n28298 = n28269 & n28297;
  assign n28299 = n4538 & n8320;
  assign n28300 = n8754 & n28299;
  assign n28301 = ~n513 & ~n649;
  assign n28302 = ~n1487 & n28301;
  assign n28303 = n4319 & n4751;
  assign n28304 = n28302 & n28303;
  assign n28305 = n6327 & n54598;
  assign n28306 = n28304 & n28305;
  assign n28307 = n4751 & n6327;
  assign n28308 = n54598 & n28307;
  assign n28309 = n8754 & n28308;
  assign n28310 = n4538 & n28309;
  assign n28311 = n4319 & n28310;
  assign n28312 = ~n1487 & n28311;
  assign n28313 = ~n271 & n28312;
  assign n28314 = ~n161 & n28313;
  assign n28315 = ~n513 & n28314;
  assign n28316 = ~n649 & n28315;
  assign n28317 = n4751 & n8320;
  assign n28318 = n8754 & n28317;
  assign n28319 = n4319 & n4538;
  assign n28320 = n28302 & n28319;
  assign n28321 = n28305 & n28320;
  assign n28322 = n28318 & n28321;
  assign n28323 = n4538 & n4751;
  assign n28324 = n8320 & n28323;
  assign n28325 = n4319 & n8754;
  assign n28326 = n28302 & n28325;
  assign n28327 = n28305 & n28326;
  assign n28328 = n28324 & n28327;
  assign n28329 = n8754 & n28323;
  assign n28330 = ~n161 & ~n649;
  assign n28331 = ~n1487 & n28330;
  assign n28332 = ~n271 & ~n513;
  assign n28333 = n4319 & n28332;
  assign n28334 = n28331 & n28333;
  assign n28335 = n28305 & n28334;
  assign n28336 = n28329 & n28335;
  assign n28337 = n28300 & n28306;
  assign n28338 = n1467 & n5955;
  assign n28339 = n16984 & n28338;
  assign n28340 = ~n112 & ~n184;
  assign n28341 = ~n495 & ~n851;
  assign n28342 = ~n112 & ~n495;
  assign n28343 = ~n184 & ~n851;
  assign n28344 = n28342 & n28343;
  assign n28345 = n28340 & n28341;
  assign n28346 = n53804 & n56745;
  assign n28347 = n56593 & n28346;
  assign n28348 = n53804 & n56593;
  assign n28349 = n5955 & n28348;
  assign n28350 = n1467 & n28349;
  assign n28351 = ~n184 & n28350;
  assign n28352 = ~n112 & n28351;
  assign n28353 = ~n495 & n28352;
  assign n28354 = ~n849 & n28353;
  assign n28355 = ~n851 & n28354;
  assign n28356 = ~n651 & n28355;
  assign n28357 = n1467 & n28340;
  assign n28358 = n5955 & n28357;
  assign n28359 = n16984 & n28341;
  assign n28360 = n53804 & n28359;
  assign n28361 = n56593 & n28360;
  assign n28362 = n28358 & n28361;
  assign n28363 = ~n849 & ~n851;
  assign n28364 = n5955 & n28363;
  assign n28365 = n1467 & n28364;
  assign n28366 = ~n112 & ~n651;
  assign n28367 = ~n184 & ~n495;
  assign n28368 = n28366 & n28367;
  assign n28369 = n53804 & n28368;
  assign n28370 = n56593 & n28369;
  assign n28371 = n28365 & n28370;
  assign n28372 = n28339 & n28347;
  assign n28373 = n56744 & n56746;
  assign n28374 = n28298 & n28373;
  assign n28375 = n53797 & n8196;
  assign n28376 = n53753 & n28375;
  assign n28377 = n54239 & n28376;
  assign n28378 = n54493 & n28377;
  assign n28379 = n56744 & n28378;
  assign n28380 = n56746 & n28379;
  assign n28381 = n56742 & n28380;
  assign n28382 = n1265 & n28381;
  assign n28383 = n9331 & n28382;
  assign n28384 = n749 & n28383;
  assign n28385 = n2340 & n28384;
  assign n28386 = n3950 & n28385;
  assign n28387 = ~n1033 & n28386;
  assign n28388 = ~n179 & n28387;
  assign n28389 = ~n770 & n28388;
  assign n28390 = n54239 & n28374;
  assign n28391 = ~n647 & ~n1189;
  assign n28392 = n3062 & n28391;
  assign n28393 = n7016 & n7094;
  assign n28394 = ~n647 & ~n1195;
  assign n28395 = ~n956 & ~n1189;
  assign n28396 = n28394 & n28395;
  assign n28397 = n3062 & n7016;
  assign n28398 = n28396 & n28397;
  assign n28399 = n28392 & n28393;
  assign n28400 = n54077 & n56748;
  assign n28401 = n54077 & n54158;
  assign n28402 = n7016 & n28401;
  assign n28403 = n3062 & n28402;
  assign n28404 = ~n1195 & n28403;
  assign n28405 = ~n956 & n28404;
  assign n28406 = ~n1189 & n28405;
  assign n28407 = ~n647 & n28406;
  assign n28408 = n54158 & n28400;
  assign n28409 = ~n402 & ~n499;
  assign n28410 = ~n883 & ~n1088;
  assign n28411 = n28409 & n28410;
  assign n28412 = n2854 & n3561;
  assign n28413 = n28411 & n28412;
  assign n28414 = n53858 & n54772;
  assign n28415 = n28413 & n28414;
  assign n28416 = ~n211 & ~n495;
  assign n28417 = ~n211 & ~n1455;
  assign n28418 = ~n495 & n28417;
  assign n28419 = ~n1455 & n28416;
  assign n28420 = ~n216 & ~n419;
  assign n28421 = ~n415 & ~n419;
  assign n28422 = ~n216 & ~n1191;
  assign n28423 = n28421 & n28422;
  assign n28424 = n13941 & n28420;
  assign n28425 = ~n415 & n56750;
  assign n28426 = ~n1191 & n28425;
  assign n28427 = ~n216 & n28426;
  assign n28428 = ~n419 & n28427;
  assign n28429 = n56750 & n56751;
  assign n28430 = n4261 & n7275;
  assign n28431 = n12112 & n28430;
  assign n28432 = n54120 & n28431;
  assign n28433 = n56752 & n28432;
  assign n28434 = ~n402 & ~n460;
  assign n28435 = ~n499 & ~n1088;
  assign n28436 = n28434 & n28435;
  assign n28437 = ~n883 & ~n1337;
  assign n28438 = n3561 & n28437;
  assign n28439 = n28436 & n28438;
  assign n28440 = n28414 & n28439;
  assign n28441 = n2854 & n4261;
  assign n28442 = n7275 & n28441;
  assign n28443 = n54120 & n28442;
  assign n28444 = n56752 & n28443;
  assign n28445 = n28440 & n28444;
  assign n28446 = n4261 & n28437;
  assign n28447 = n28436 & n28446;
  assign n28448 = n28414 & n28447;
  assign n28449 = n3561 & n7275;
  assign n28450 = n2854 & n28449;
  assign n28451 = n54120 & n28450;
  assign n28452 = n56752 & n28451;
  assign n28453 = n28448 & n28452;
  assign n28454 = n28415 & n28433;
  assign n28455 = n56749 & n56753;
  assign n28456 = n53961 & n54391;
  assign n28457 = n2854 & n54120;
  assign n28458 = n53858 & n28457;
  assign n28459 = n54772 & n28458;
  assign n28460 = n7275 & n28459;
  assign n28461 = n54391 & n28460;
  assign n28462 = n56749 & n28461;
  assign n28463 = n53961 & n28462;
  assign n28464 = n4261 & n28463;
  assign n28465 = n56752 & n28464;
  assign n28466 = n3561 & n28465;
  assign n28467 = ~n1088 & n28466;
  assign n28468 = ~n883 & n28467;
  assign n28469 = ~n402 & n28468;
  assign n28470 = ~n1337 & n28469;
  assign n28471 = ~n460 & n28470;
  assign n28472 = ~n499 & n28471;
  assign n28473 = n28455 & n28456;
  assign n28474 = ~n56747 & ~n56754;
  assign n28475 = ~n21237 & ~n21269;
  assign n28476 = ~n20073 & ~n20085;
  assign n28477 = ~n55472 & ~n20085;
  assign n28478 = n56755 & n28477;
  assign n28479 = ~n55472 & n56755;
  assign n28480 = ~n20085 & n28479;
  assign n28481 = n20073 & ~n55471;
  assign n28482 = pi8  & n56756;
  assign n28483 = ~pi8  & ~n56756;
  assign n28484 = ~n28482 & ~n28483;
  assign n28485 = n56747 & n56754;
  assign n28486 = ~n28474 & ~n28485;
  assign n28487 = n28484 & n28486;
  assign n28488 = ~n28474 & ~n28487;
  assign n28489 = n56713 & ~n28488;
  assign n28490 = ~n56713 & n28488;
  assign n28491 = ~n28489 & ~n28490;
  assign n28492 = n26437 & ~n26439;
  assign n28493 = ~n26440 & ~n28492;
  assign n28494 = n1576 & n28493;
  assign n28495 = n11215 & n26295;
  assign n28496 = n10564 & n26298;
  assign n28497 = n54403 & n26301;
  assign n28498 = ~n28496 & ~n28497;
  assign n28499 = ~n28495 & n28498;
  assign n28500 = ~n28494 & ~n28497;
  assign n28501 = ~n28496 & n28500;
  assign n28502 = ~n28495 & n28501;
  assign n28503 = ~n28494 & n28499;
  assign n28504 = n28491 & ~n56757;
  assign n28505 = ~n28489 & ~n28504;
  assign n28506 = ~n56713 & n56736;
  assign n28507 = ~n28256 & ~n28506;
  assign n28508 = ~n28256 & ~n28505;
  assign n28509 = ~n28506 & n28508;
  assign n28510 = ~n28505 & n28507;
  assign n28511 = ~n28256 & ~n56758;
  assign n28512 = ~n28105 & n28114;
  assign n28513 = n28105 & ~n28115;
  assign n28514 = n28105 & n28114;
  assign n28515 = ~n28114 & ~n28115;
  assign n28516 = ~n28105 & ~n28114;
  assign n28517 = ~n56759 & ~n56760;
  assign n28518 = ~n28115 & ~n28512;
  assign n28519 = ~n28511 & ~n56761;
  assign n28520 = ~n28115 & ~n28519;
  assign n28521 = ~n28078 & n56722;
  assign n28522 = ~n28094 & ~n28521;
  assign n28523 = ~n28520 & n28522;
  assign n28524 = n28520 & ~n28522;
  assign n28525 = ~n28523 & ~n28524;
  assign n28526 = n11279 & n27330;
  assign n28527 = n12584 & n26277;
  assign n28528 = n54410 & n26283;
  assign n28529 = n11267 & n26280;
  assign n28530 = ~n28528 & ~n28529;
  assign n28531 = ~n28527 & n28530;
  assign n28532 = ~n11279 & n28531;
  assign n28533 = ~n27330 & n28531;
  assign n28534 = ~n28532 & ~n28533;
  assign n28535 = ~n28526 & n28531;
  assign n28536 = pi29  & ~n56762;
  assign n28537 = ~pi29  & n56762;
  assign n28538 = ~n28536 & ~n28537;
  assign n28539 = n28525 & ~n28538;
  assign n28540 = ~n28523 & ~n28539;
  assign n28541 = n28103 & ~n28540;
  assign n28542 = ~n28101 & ~n28541;
  assign n28543 = n27878 & n56708;
  assign n28544 = ~n56708 & ~n27884;
  assign n28545 = ~n27878 & ~n27884;
  assign n28546 = ~n28544 & ~n28545;
  assign n28547 = ~n27884 & ~n28543;
  assign n28548 = ~n28542 & ~n56763;
  assign n28549 = ~n27884 & ~n28548;
  assign n28550 = ~n27758 & n27771;
  assign n28551 = ~n27772 & ~n28550;
  assign n28552 = ~n28549 & n28551;
  assign n28553 = n28549 & ~n28551;
  assign n28554 = n123 & ~n56639;
  assign n28555 = n128 & n26259;
  assign n28556 = n53444 & n26265;
  assign n28557 = n127 & n26262;
  assign n28558 = ~n28556 & ~n28557;
  assign n28559 = ~n28555 & n28558;
  assign n28560 = ~n28554 & n28559;
  assign n28561 = pi26  & ~n28560;
  assign n28562 = pi26  & ~n28561;
  assign n28563 = pi26  & n28560;
  assign n28564 = ~n28560 & ~n28561;
  assign n28565 = ~pi26  & ~n28560;
  assign n28566 = ~n56764 & ~n56765;
  assign n28567 = ~n28553 & ~n28566;
  assign n28568 = ~n28552 & ~n28553;
  assign n28569 = ~n28566 & n28568;
  assign n28570 = ~n28552 & ~n28569;
  assign n28571 = ~n28552 & ~n28567;
  assign n28572 = ~n56705 & ~n56766;
  assign n28573 = n56705 & n56766;
  assign n28574 = n90 & ~n56567;
  assign n28575 = n14236 & n26247;
  assign n28576 = n54667 & n26253;
  assign n28577 = n14210 & n26250;
  assign n28578 = ~n28576 & ~n28577;
  assign n28579 = ~n28575 & n28578;
  assign n28580 = ~n28574 & n28579;
  assign n28581 = pi23  & ~n28580;
  assign n28582 = pi23  & ~n28581;
  assign n28583 = pi23  & n28580;
  assign n28584 = ~n28580 & ~n28581;
  assign n28585 = ~pi23  & ~n28580;
  assign n28586 = ~n56767 & ~n56768;
  assign n28587 = ~n28573 & ~n28586;
  assign n28588 = ~n28572 & ~n28573;
  assign n28589 = ~n28586 & n28588;
  assign n28590 = ~n28572 & ~n28589;
  assign n28591 = ~n28572 & ~n28587;
  assign n28592 = ~n56704 & ~n56769;
  assign n28593 = ~n27853 & ~n28592;
  assign n28594 = n27821 & ~n27823;
  assign n28595 = n27823 & ~n27824;
  assign n28596 = n27821 & n27823;
  assign n28597 = ~n27821 & ~n27824;
  assign n28598 = ~n27821 & ~n27823;
  assign n28599 = ~n56770 & ~n56771;
  assign n28600 = ~n27824 & ~n28594;
  assign n28601 = ~n28593 & ~n56772;
  assign n28602 = n28593 & n56772;
  assign n28603 = n54719 & ~n26537;
  assign n28604 = ~n15901 & ~n28603;
  assign n28605 = ~n15921 & n28604;
  assign n28606 = ~n15921 & ~n28603;
  assign n28607 = ~n15901 & n28606;
  assign n28608 = n56666 & ~n28603;
  assign n28609 = ~n14413 & n56773;
  assign n28610 = pi20  & ~n28609;
  assign n28611 = pi20  & ~n28610;
  assign n28612 = pi20  & n28609;
  assign n28613 = ~n28609 & ~n28610;
  assign n28614 = ~pi20  & ~n28609;
  assign n28615 = ~n56774 & ~n56775;
  assign n28616 = ~n28602 & ~n28615;
  assign n28617 = ~n28601 & ~n28602;
  assign n28618 = ~n28615 & n28617;
  assign n28619 = ~n28601 & ~n28618;
  assign n28620 = ~n28601 & ~n28616;
  assign n28621 = ~n56699 & ~n56776;
  assign n28622 = n56699 & n56776;
  assign n28623 = ~n28621 & ~n28622;
  assign n28624 = ~n26537 & ~n26541;
  assign n28625 = n14413 & n28624;
  assign n28626 = n15901 & ~n26537;
  assign n28627 = n54719 & n26242;
  assign n28628 = ~n15921 & ~n28627;
  assign n28629 = ~n28626 & ~n28627;
  assign n28630 = ~n15921 & n28629;
  assign n28631 = ~n28626 & n28628;
  assign n28632 = ~n28625 & n56777;
  assign n28633 = pi20  & ~n28632;
  assign n28634 = pi20  & ~n28633;
  assign n28635 = pi20  & n28632;
  assign n28636 = ~n28632 & ~n28633;
  assign n28637 = ~pi20  & ~n28632;
  assign n28638 = ~n56778 & ~n56779;
  assign n28639 = n28586 & ~n28588;
  assign n28640 = n28588 & ~n28589;
  assign n28641 = ~n28586 & ~n28589;
  assign n28642 = ~n28640 & ~n28641;
  assign n28643 = ~n28589 & ~n28639;
  assign n28644 = n28542 & n56763;
  assign n28645 = ~n28548 & ~n28644;
  assign n28646 = n123 & n27466;
  assign n28647 = n128 & n26262;
  assign n28648 = n53444 & n26268;
  assign n28649 = n127 & n26265;
  assign n28650 = ~n28648 & ~n28649;
  assign n28651 = ~n28647 & n28650;
  assign n28652 = ~n28646 & n28651;
  assign n28653 = pi26  & ~n28652;
  assign n28654 = pi26  & ~n28653;
  assign n28655 = pi26  & n28652;
  assign n28656 = ~n28652 & ~n28653;
  assign n28657 = ~pi26  & ~n28652;
  assign n28658 = ~n56781 & ~n56782;
  assign n28659 = n28645 & ~n28658;
  assign n28660 = ~n28103 & n28540;
  assign n28661 = ~n28541 & ~n28660;
  assign n28662 = n11279 & ~n56648;
  assign n28663 = n12584 & n26274;
  assign n28664 = n54410 & n26280;
  assign n28665 = n11267 & n26277;
  assign n28666 = ~n28664 & ~n28665;
  assign n28667 = ~n28663 & n28666;
  assign n28668 = ~n28662 & n28667;
  assign n28669 = pi29  & ~n28668;
  assign n28670 = pi29  & ~n28669;
  assign n28671 = pi29  & n28668;
  assign n28672 = ~n28668 & ~n28669;
  assign n28673 = ~pi29  & ~n28668;
  assign n28674 = ~n56783 & ~n56784;
  assign n28675 = n28661 & ~n28674;
  assign n28676 = n123 & n27042;
  assign n28677 = n128 & n26265;
  assign n28678 = n53444 & n26271;
  assign n28679 = n127 & n26268;
  assign n28680 = ~n28678 & ~n28679;
  assign n28681 = ~n28677 & n28680;
  assign n28682 = ~n28676 & n28681;
  assign n28683 = pi26  & ~n28682;
  assign n28684 = pi26  & ~n28683;
  assign n28685 = pi26  & n28682;
  assign n28686 = ~n28682 & ~n28683;
  assign n28687 = ~pi26  & ~n28682;
  assign n28688 = ~n56785 & ~n56786;
  assign n28689 = ~n28661 & n28674;
  assign n28690 = n28661 & ~n28675;
  assign n28691 = n28661 & n28674;
  assign n28692 = ~n28674 & ~n28675;
  assign n28693 = ~n28661 & ~n28674;
  assign n28694 = ~n56787 & ~n56788;
  assign n28695 = ~n28675 & ~n28689;
  assign n28696 = ~n28688 & ~n56789;
  assign n28697 = ~n28675 & ~n28696;
  assign n28698 = ~n28645 & n28658;
  assign n28699 = n28645 & ~n28659;
  assign n28700 = n28645 & n28658;
  assign n28701 = ~n28658 & ~n28659;
  assign n28702 = ~n28645 & ~n28658;
  assign n28703 = ~n56790 & ~n56791;
  assign n28704 = ~n28659 & ~n28698;
  assign n28705 = ~n28697 & ~n56792;
  assign n28706 = ~n28659 & ~n28705;
  assign n28707 = n28566 & ~n28568;
  assign n28708 = n28568 & ~n28569;
  assign n28709 = ~n28566 & ~n28569;
  assign n28710 = ~n28708 & ~n28709;
  assign n28711 = ~n28569 & ~n28707;
  assign n28712 = ~n28706 & ~n56793;
  assign n28713 = n28706 & n56793;
  assign n28714 = n90 & n27491;
  assign n28715 = n14236 & n26250;
  assign n28716 = n54667 & n26256;
  assign n28717 = n14210 & n26253;
  assign n28718 = ~n28716 & ~n28717;
  assign n28719 = ~n28715 & n28718;
  assign n28720 = ~n28714 & n28719;
  assign n28721 = pi23  & ~n28720;
  assign n28722 = pi23  & ~n28721;
  assign n28723 = pi23  & n28720;
  assign n28724 = ~n28720 & ~n28721;
  assign n28725 = ~pi23  & ~n28720;
  assign n28726 = ~n56794 & ~n56795;
  assign n28727 = ~n28713 & ~n28726;
  assign n28728 = ~n28712 & ~n28713;
  assign n28729 = ~n28726 & n28728;
  assign n28730 = ~n28712 & ~n28729;
  assign n28731 = ~n28712 & ~n28727;
  assign n28732 = ~n56780 & ~n56796;
  assign n28733 = n56780 & n56796;
  assign n28734 = n14413 & ~n56564;
  assign n28735 = n15921 & ~n26537;
  assign n28736 = n54719 & n26244;
  assign n28737 = n15901 & n26242;
  assign n28738 = ~n28736 & ~n28737;
  assign n28739 = ~n28735 & n28738;
  assign n28740 = ~n28734 & n28739;
  assign n28741 = pi20  & ~n28740;
  assign n28742 = pi20  & ~n28741;
  assign n28743 = pi20  & n28740;
  assign n28744 = ~n28740 & ~n28741;
  assign n28745 = ~pi20  & ~n28740;
  assign n28746 = ~n56797 & ~n56798;
  assign n28747 = ~n28733 & ~n28746;
  assign n28748 = ~n28732 & ~n28733;
  assign n28749 = ~n28746 & n28748;
  assign n28750 = ~n28732 & ~n28749;
  assign n28751 = ~n28732 & ~n28747;
  assign n28752 = ~n28638 & ~n56799;
  assign n28753 = n56704 & n56769;
  assign n28754 = ~n28592 & ~n28753;
  assign n28755 = n28638 & n56799;
  assign n28756 = ~n56799 & ~n28752;
  assign n28757 = n28638 & ~n56799;
  assign n28758 = ~n28638 & ~n28752;
  assign n28759 = ~n28638 & n56799;
  assign n28760 = ~n56800 & ~n56801;
  assign n28761 = ~n28752 & ~n28755;
  assign n28762 = n28754 & ~n56802;
  assign n28763 = ~n28752 & ~n28762;
  assign n28764 = n28615 & ~n28617;
  assign n28765 = n28617 & ~n28618;
  assign n28766 = ~n28615 & ~n28618;
  assign n28767 = ~n28765 & ~n28766;
  assign n28768 = ~n28618 & ~n28764;
  assign n28769 = ~n28763 & ~n56803;
  assign n28770 = ~n28754 & n56802;
  assign n28771 = ~n28762 & ~n28770;
  assign n28772 = n28697 & n56792;
  assign n28773 = ~n28705 & ~n28772;
  assign n28774 = n90 & ~n56668;
  assign n28775 = n14236 & n26253;
  assign n28776 = n54667 & n26259;
  assign n28777 = n14210 & n26256;
  assign n28778 = ~n28776 & ~n28777;
  assign n28779 = ~n28775 & n28778;
  assign n28780 = ~n28774 & n28779;
  assign n28781 = pi23  & ~n28780;
  assign n28782 = pi23  & ~n28781;
  assign n28783 = pi23  & n28780;
  assign n28784 = ~n28780 & ~n28781;
  assign n28785 = ~pi23  & ~n28780;
  assign n28786 = ~n56804 & ~n56805;
  assign n28787 = n28773 & ~n28786;
  assign n28788 = ~n28773 & n28786;
  assign n28789 = n28773 & ~n28787;
  assign n28790 = n28773 & n28786;
  assign n28791 = ~n28786 & ~n28787;
  assign n28792 = ~n28773 & ~n28786;
  assign n28793 = ~n56806 & ~n56807;
  assign n28794 = ~n28787 & ~n28788;
  assign n28795 = n28688 & n56789;
  assign n28796 = ~n56789 & ~n28696;
  assign n28797 = ~n28688 & ~n28696;
  assign n28798 = ~n28796 & ~n28797;
  assign n28799 = ~n28696 & ~n28795;
  assign n28800 = ~n28525 & n28538;
  assign n28801 = ~n28539 & ~n28800;
  assign n28802 = n28505 & ~n28507;
  assign n28803 = ~n28505 & ~n56758;
  assign n28804 = ~n28506 & n28511;
  assign n28805 = ~n28803 & ~n28804;
  assign n28806 = ~n56758 & ~n28802;
  assign n28807 = n26441 & ~n26443;
  assign n28808 = ~n26444 & ~n28807;
  assign n28809 = n1576 & n28808;
  assign n28810 = n11215 & n26292;
  assign n28811 = n54403 & n26298;
  assign n28812 = n10564 & n26295;
  assign n28813 = ~n28811 & ~n28812;
  assign n28814 = ~n28810 & n28813;
  assign n28815 = ~n28809 & n28814;
  assign n28816 = ~n56810 & ~n28815;
  assign n28817 = n11279 & ~n56686;
  assign n28818 = n12584 & n26283;
  assign n28819 = n54410 & n26289;
  assign n28820 = n11267 & n26286;
  assign n28821 = ~n28819 & ~n28820;
  assign n28822 = ~n28818 & n28821;
  assign n28823 = ~n11279 & n28822;
  assign n28824 = n56686 & n28822;
  assign n28825 = ~n28823 & ~n28824;
  assign n28826 = ~n28817 & n28822;
  assign n28827 = pi29  & ~n56811;
  assign n28828 = ~pi29  & n56811;
  assign n28829 = ~n28827 & ~n28828;
  assign n28830 = n56810 & n28815;
  assign n28831 = ~n56810 & ~n28816;
  assign n28832 = ~n56810 & n28815;
  assign n28833 = ~n28815 & ~n28816;
  assign n28834 = n56810 & ~n28815;
  assign n28835 = ~n56812 & ~n56813;
  assign n28836 = ~n28816 & ~n28830;
  assign n28837 = ~n28829 & ~n56814;
  assign n28838 = ~n28816 & ~n28837;
  assign n28839 = n28511 & n56761;
  assign n28840 = ~n56761 & ~n28519;
  assign n28841 = n28511 & ~n56761;
  assign n28842 = ~n28511 & ~n28519;
  assign n28843 = ~n28511 & n56761;
  assign n28844 = ~n56815 & ~n56816;
  assign n28845 = ~n28519 & ~n28839;
  assign n28846 = ~n28838 & ~n56817;
  assign n28847 = n28838 & n56817;
  assign n28848 = n11279 & n27743;
  assign n28849 = n12584 & n26280;
  assign n28850 = n54410 & n26286;
  assign n28851 = n11267 & n26283;
  assign n28852 = ~n28850 & ~n28851;
  assign n28853 = ~n28849 & n28852;
  assign n28854 = ~n28848 & n28853;
  assign n28855 = pi29  & ~n28854;
  assign n28856 = pi29  & ~n28855;
  assign n28857 = pi29  & n28854;
  assign n28858 = ~n28854 & ~n28855;
  assign n28859 = ~pi29  & ~n28854;
  assign n28860 = ~n56818 & ~n56819;
  assign n28861 = ~n28847 & ~n28860;
  assign n28862 = ~n28838 & ~n28846;
  assign n28863 = ~n56817 & ~n28846;
  assign n28864 = ~n28862 & ~n28863;
  assign n28865 = ~n28846 & ~n28847;
  assign n28866 = ~n28860 & ~n56820;
  assign n28867 = ~n28846 & ~n28866;
  assign n28868 = ~n28846 & ~n28861;
  assign n28869 = n28801 & ~n56821;
  assign n28870 = ~n28801 & n56821;
  assign n28871 = n123 & ~n56601;
  assign n28872 = n128 & n26268;
  assign n28873 = n53444 & n26274;
  assign n28874 = n127 & n26271;
  assign n28875 = ~n28873 & ~n28874;
  assign n28876 = ~n28872 & n28875;
  assign n28877 = ~n28871 & n28876;
  assign n28878 = pi26  & ~n28877;
  assign n28879 = pi26  & ~n28878;
  assign n28880 = pi26  & n28877;
  assign n28881 = ~n28877 & ~n28878;
  assign n28882 = ~pi26  & ~n28877;
  assign n28883 = ~n56822 & ~n56823;
  assign n28884 = ~n28870 & ~n28883;
  assign n28885 = ~n28869 & ~n28870;
  assign n28886 = ~n28883 & n28885;
  assign n28887 = ~n28869 & ~n28886;
  assign n28888 = ~n28869 & ~n28884;
  assign n28889 = ~n56809 & ~n56824;
  assign n28890 = n56809 & n56824;
  assign n28891 = n90 & n27387;
  assign n28892 = n14236 & n26256;
  assign n28893 = n54667 & n26262;
  assign n28894 = n14210 & n26259;
  assign n28895 = ~n28893 & ~n28894;
  assign n28896 = ~n28892 & n28895;
  assign n28897 = ~n28891 & n28896;
  assign n28898 = pi23  & ~n28897;
  assign n28899 = pi23  & ~n28898;
  assign n28900 = pi23  & n28897;
  assign n28901 = ~n28897 & ~n28898;
  assign n28902 = ~pi23  & ~n28897;
  assign n28903 = ~n56825 & ~n56826;
  assign n28904 = ~n28890 & ~n28903;
  assign n28905 = ~n28889 & ~n28890;
  assign n28906 = ~n28903 & n28905;
  assign n28907 = ~n28889 & ~n28906;
  assign n28908 = ~n28889 & ~n28904;
  assign n28909 = ~n56808 & ~n56827;
  assign n28910 = ~n28787 & ~n28909;
  assign n28911 = n28728 & ~n28729;
  assign n28912 = n28726 & n28728;
  assign n28913 = ~n28726 & ~n28729;
  assign n28914 = ~n28726 & ~n28728;
  assign n28915 = n28726 & ~n28728;
  assign n28916 = ~n28729 & ~n28915;
  assign n28917 = ~n56828 & ~n56829;
  assign n28918 = ~n28910 & n56830;
  assign n28919 = n28910 & ~n56830;
  assign n28920 = n14413 & n27808;
  assign n28921 = n15921 & n26242;
  assign n28922 = n54719 & n26247;
  assign n28923 = n15901 & n26244;
  assign n28924 = ~n28922 & ~n28923;
  assign n28925 = ~n28921 & n28924;
  assign n28926 = ~n28920 & n28925;
  assign n28927 = pi20  & ~n28926;
  assign n28928 = pi20  & ~n28927;
  assign n28929 = pi20  & n28926;
  assign n28930 = ~n28926 & ~n28927;
  assign n28931 = ~pi20  & ~n28926;
  assign n28932 = ~n56831 & ~n56832;
  assign n28933 = ~n28919 & ~n28932;
  assign n28934 = ~n28918 & ~n28919;
  assign n28935 = ~n28932 & n28934;
  assign n28936 = ~n28918 & ~n28935;
  assign n28937 = ~n28918 & ~n28933;
  assign n28938 = ~n26879 & ~n56833;
  assign n28939 = n26879 & n56833;
  assign n28940 = n28746 & ~n28748;
  assign n28941 = n28748 & ~n28749;
  assign n28942 = ~n28746 & ~n28749;
  assign n28943 = ~n28941 & ~n28942;
  assign n28944 = ~n28749 & ~n28940;
  assign n28945 = ~n28939 & ~n56834;
  assign n28946 = ~n28938 & ~n28939;
  assign n28947 = ~n56834 & n28946;
  assign n28948 = ~n28938 & ~n28947;
  assign n28949 = ~n28938 & ~n28945;
  assign n28950 = n28771 & ~n56835;
  assign n28951 = n56834 & ~n28946;
  assign n28952 = ~n56834 & ~n28947;
  assign n28953 = n28946 & ~n28947;
  assign n28954 = ~n28952 & ~n28953;
  assign n28955 = ~n28947 & ~n28951;
  assign n28956 = n56808 & n56827;
  assign n28957 = ~n28909 & ~n28956;
  assign n28958 = n14413 & n27839;
  assign n28959 = n15921 & n26244;
  assign n28960 = n54719 & n26250;
  assign n28961 = n15901 & n26247;
  assign n28962 = ~n28960 & ~n28961;
  assign n28963 = ~n28959 & n28962;
  assign n28964 = ~n28958 & n28963;
  assign n28965 = pi20  & ~n28964;
  assign n28966 = pi20  & ~n28965;
  assign n28967 = pi20  & n28964;
  assign n28968 = ~n28964 & ~n28965;
  assign n28969 = ~pi20  & ~n28964;
  assign n28970 = ~n56837 & ~n56838;
  assign n28971 = n28957 & ~n28970;
  assign n28972 = ~n28957 & n28970;
  assign n28973 = n28957 & ~n28971;
  assign n28974 = n28957 & n28970;
  assign n28975 = ~n28970 & ~n28971;
  assign n28976 = ~n28957 & ~n28970;
  assign n28977 = ~n56839 & ~n56840;
  assign n28978 = ~n28971 & ~n28972;
  assign n28979 = n28903 & ~n28905;
  assign n28980 = n28905 & ~n28906;
  assign n28981 = ~n28903 & ~n28906;
  assign n28982 = ~n28980 & ~n28981;
  assign n28983 = ~n28906 & ~n28979;
  assign n28984 = n123 & ~n56612;
  assign n28985 = n128 & n26271;
  assign n28986 = n53444 & n26277;
  assign n28987 = n127 & n26274;
  assign n28988 = ~n28986 & ~n28987;
  assign n28989 = ~n28985 & n28988;
  assign n28990 = ~n28984 & n28989;
  assign n28991 = pi26  & ~n28990;
  assign n28992 = pi26  & ~n28991;
  assign n28993 = pi26  & n28990;
  assign n28994 = ~n28990 & ~n28991;
  assign n28995 = ~pi26  & ~n28990;
  assign n28996 = ~n56843 & ~n56844;
  assign n28997 = n28860 & n56820;
  assign n28998 = ~n56820 & ~n28866;
  assign n28999 = ~n28860 & ~n28866;
  assign n29000 = ~n28998 & ~n28999;
  assign n29001 = ~n28866 & ~n28997;
  assign n29002 = ~n28996 & ~n56845;
  assign n29003 = n28996 & n56845;
  assign n29004 = ~n56845 & ~n29002;
  assign n29005 = n28996 & ~n56845;
  assign n29006 = ~n28996 & ~n29002;
  assign n29007 = ~n28996 & n56845;
  assign n29008 = ~n56846 & ~n56847;
  assign n29009 = ~n29002 & ~n29003;
  assign n29010 = ~n28491 & n56757;
  assign n29011 = ~n28504 & ~n29010;
  assign n29012 = ~n419 & ~n649;
  assign n29013 = ~n977 & ~n1088;
  assign n29014 = n29012 & n29013;
  assign n29015 = n358 & n417;
  assign n29016 = n29014 & n29015;
  assign n29017 = ~n295 & ~n751;
  assign n29018 = ~n295 & n1672;
  assign n29019 = ~n751 & n29018;
  assign n29020 = n1672 & n29017;
  assign n29021 = n54804 & n56849;
  assign n29022 = n29016 & n29021;
  assign n29023 = n494 & n2327;
  assign n29024 = n4320 & n8267;
  assign n29025 = n29023 & n29024;
  assign n29026 = n53716 & n29025;
  assign n29027 = n358 & n494;
  assign n29028 = n29014 & n29027;
  assign n29029 = n29021 & n29028;
  assign n29030 = n417 & n2327;
  assign n29031 = n29024 & n29030;
  assign n29032 = n53716 & n29031;
  assign n29033 = n29029 & n29032;
  assign n29034 = ~n419 & ~n977;
  assign n29035 = ~n1088 & ~n1191;
  assign n29036 = n29034 & n29035;
  assign n29037 = ~n649 & ~n2103;
  assign n29038 = n4320 & n29037;
  assign n29039 = n29036 & n29038;
  assign n29040 = n29021 & n29039;
  assign n29041 = n358 & n8267;
  assign n29042 = n417 & n494;
  assign n29043 = n29041 & n29042;
  assign n29044 = n53716 & n29043;
  assign n29045 = n29040 & n29044;
  assign n29046 = n29022 & n29026;
  assign n29047 = n53726 & n56850;
  assign n29048 = n54104 & n29047;
  assign n29049 = n4320 & n54804;
  assign n29050 = n56849 & n29049;
  assign n29051 = n8267 & n29050;
  assign n29052 = n54144 & n29051;
  assign n29053 = n53716 & n29052;
  assign n29054 = n417 & n29053;
  assign n29055 = n53726 & n29054;
  assign n29056 = n494 & n29055;
  assign n29057 = n358 & n29056;
  assign n29058 = n54104 & n29057;
  assign n29059 = ~n1088 & n29058;
  assign n29060 = ~n1191 & n29059;
  assign n29061 = ~n977 & n29060;
  assign n29062 = ~n2103 & n29061;
  assign n29063 = ~n649 & n29062;
  assign n29064 = ~n419 & n29063;
  assign n29065 = n54144 & n29048;
  assign n29066 = n56747 & ~n56851;
  assign n29067 = ~n25272 & ~n25287;
  assign n29068 = ~n24330 & ~n24338;
  assign n29069 = ~n24337 & n56852;
  assign n29070 = ~n24338 & n29069;
  assign n29071 = n24330 & ~n56258;
  assign n29072 = n24337 & ~n26537;
  assign n29073 = ~n25272 & ~n29072;
  assign n29074 = ~n25287 & n29073;
  assign n29075 = ~n25287 & ~n29072;
  assign n29076 = ~n25272 & n29075;
  assign n29077 = n56852 & ~n29072;
  assign n29078 = ~n24338 & n56854;
  assign n29079 = ~pi2  & ~n29078;
  assign n29080 = ~pi2  & ~n56853;
  assign n29081 = ~n218 & ~n776;
  assign n29082 = ~n1472 & n29081;
  assign n29083 = n3636 & n4070;
  assign n29084 = n4470 & n5955;
  assign n29085 = n29083 & n29084;
  assign n29086 = n29082 & n29085;
  assign n29087 = n7350 & n9396;
  assign n29088 = n11155 & n29087;
  assign n29089 = n53736 & n29088;
  assign n29090 = n5955 & n7350;
  assign n29091 = n7350 & n11155;
  assign n29092 = n5955 & n29091;
  assign n29093 = n11155 & n29090;
  assign n29094 = n53736 & n56856;
  assign n29095 = n4470 & n29094;
  assign n29096 = n4070 & n29095;
  assign n29097 = ~n1472 & n29096;
  assign n29098 = ~n218 & n29097;
  assign n29099 = ~n612 & n29098;
  assign n29100 = ~n460 & n29099;
  assign n29101 = ~n450 & n29100;
  assign n29102 = ~n776 & n29101;
  assign n29103 = ~n346 & n29102;
  assign n29104 = ~n218 & ~n612;
  assign n29105 = ~n460 & n29104;
  assign n29106 = ~n776 & ~n1472;
  assign n29107 = n4470 & n29106;
  assign n29108 = n4070 & n11155;
  assign n29109 = n29107 & n29108;
  assign n29110 = n29105 & n29109;
  assign n29111 = n9396 & n29090;
  assign n29112 = n53736 & n29111;
  assign n29113 = n29110 & n29112;
  assign n29114 = ~n346 & ~n612;
  assign n29115 = ~n460 & n29114;
  assign n29116 = ~n218 & ~n450;
  assign n29117 = n29106 & n29116;
  assign n29118 = n4070 & n4470;
  assign n29119 = n29117 & n29118;
  assign n29120 = n29115 & n29119;
  assign n29121 = n29094 & n29120;
  assign n29122 = n29086 & n29089;
  assign n29123 = ~n416 & ~n1124;
  assign n29124 = n3780 & n29123;
  assign n29125 = n3780 & n56726;
  assign n29126 = ~n1124 & n29125;
  assign n29127 = ~n416 & n29126;
  assign n29128 = n56726 & n29124;
  assign n29129 = n586 & n53807;
  assign n29130 = n53609 & n29129;
  assign n29131 = n56858 & n29130;
  assign n29132 = n5482 & n8680;
  assign n29133 = n54501 & n27277;
  assign n29134 = n29132 & n29133;
  assign n29135 = n54285 & n29134;
  assign n29136 = n586 & n8680;
  assign n29137 = n53609 & n29136;
  assign n29138 = n56858 & n29137;
  assign n29139 = n53807 & n5482;
  assign n29140 = n29133 & n29139;
  assign n29141 = n54285 & n29140;
  assign n29142 = n29138 & n29141;
  assign n29143 = n29131 & n29135;
  assign n29144 = n53807 & n29133;
  assign n29145 = n8679 & n29144;
  assign n29146 = n56858 & n29145;
  assign n29147 = n53609 & n29146;
  assign n29148 = n54285 & n29147;
  assign n29149 = n4376 & n29148;
  assign n29150 = n586 & n29149;
  assign n29151 = n56857 & n29150;
  assign n29152 = n164 & n29151;
  assign n29153 = ~n311 & n29152;
  assign n29154 = n56857 & n56859;
  assign n29155 = n4206 & n6806;
  assign n29156 = n9767 & n11428;
  assign n29157 = n29155 & n29156;
  assign n29158 = ~n447 & ~n1703;
  assign n29159 = n3085 & n29158;
  assign n29160 = n12339 & n29159;
  assign n29161 = n3085 & n4206;
  assign n29162 = n29156 & n29161;
  assign n29163 = n6806 & n29158;
  assign n29164 = n12339 & n29163;
  assign n29165 = n29162 & n29164;
  assign n29166 = n3085 & n11428;
  assign n29167 = n29155 & n29166;
  assign n29168 = n9767 & n29158;
  assign n29169 = n12339 & n29168;
  assign n29170 = n29167 & n29169;
  assign n29171 = n29157 & n29160;
  assign n29172 = n55000 & n55126;
  assign n29173 = n56861 & n29172;
  assign n29174 = n54457 & n56710;
  assign n29175 = n29173 & n29174;
  assign n29176 = n4206 & n12339;
  assign n29177 = n55000 & n29176;
  assign n29178 = n55126 & n29177;
  assign n29179 = n56710 & n29178;
  assign n29180 = n54457 & n29179;
  assign n29181 = n56860 & n29180;
  assign n29182 = n6806 & n29181;
  assign n29183 = n3085 & n29182;
  assign n29184 = n11428 & n29183;
  assign n29185 = ~n1703 & n29184;
  assign n29186 = ~n172 & n29185;
  assign n29187 = ~n294 & n29186;
  assign n29188 = ~n447 & n29187;
  assign n29189 = n56860 & n29175;
  assign n29190 = ~n56855 & ~n56862;
  assign n29191 = ~n23459 & ~n24302;
  assign n29192 = ~n77 & ~n21969;
  assign n29193 = n29191 & n29192;
  assign n29194 = ~n21969 & n29191;
  assign n29195 = ~n21962 & n29191;
  assign n29196 = ~n77 & n56864;
  assign n29197 = ~n53440 & n29191;
  assign n29198 = ~pi5  & ~n56863;
  assign n29199 = pi5  & n56863;
  assign n29200 = ~n29198 & ~n29199;
  assign n29201 = n56855 & n56862;
  assign n29202 = ~n56855 & n56862;
  assign n29203 = n56855 & ~n56862;
  assign n29204 = ~n29202 & ~n29203;
  assign n29205 = ~n29190 & ~n29201;
  assign n29206 = ~n29199 & ~n56865;
  assign n29207 = ~n29198 & n29206;
  assign n29208 = n29200 & ~n56865;
  assign n29209 = ~n29190 & ~n56866;
  assign n29210 = n56747 & ~n29209;
  assign n29211 = ~n56747 & n29209;
  assign n29212 = ~n29210 & ~n29211;
  assign n29213 = n26421 & ~n26423;
  assign n29214 = ~n26421 & ~n56552;
  assign n29215 = ~n26422 & n26427;
  assign n29216 = ~n29214 & ~n29215;
  assign n29217 = ~n56552 & ~n29213;
  assign n29218 = n1576 & ~n56867;
  assign n29219 = n11215 & n26304;
  assign n29220 = n10564 & n26307;
  assign n29221 = n54403 & n26310;
  assign n29222 = ~n29220 & ~n29221;
  assign n29223 = ~n29219 & n29222;
  assign n29224 = ~n29218 & ~n29221;
  assign n29225 = ~n29220 & n29224;
  assign n29226 = ~n29219 & n29225;
  assign n29227 = ~n29218 & n29223;
  assign n29228 = n29212 & ~n56868;
  assign n29229 = ~n29210 & ~n29228;
  assign n29230 = ~n56747 & n56851;
  assign n29231 = ~n29066 & ~n29230;
  assign n29232 = ~n29066 & ~n29229;
  assign n29233 = ~n29230 & n29232;
  assign n29234 = ~n29229 & n29231;
  assign n29235 = ~n29066 & ~n56869;
  assign n29236 = ~n28484 & ~n28486;
  assign n29237 = ~n28487 & ~n29236;
  assign n29238 = ~n29235 & n29237;
  assign n29239 = n29235 & ~n29237;
  assign n29240 = n26431 & ~n26433;
  assign n29241 = ~n26431 & ~n56553;
  assign n29242 = ~n26432 & n26437;
  assign n29243 = ~n29241 & ~n29242;
  assign n29244 = ~n56553 & ~n29240;
  assign n29245 = n1576 & ~n56870;
  assign n29246 = n11215 & n26298;
  assign n29247 = n54403 & n26304;
  assign n29248 = n10564 & n26301;
  assign n29249 = ~n29247 & ~n29248;
  assign n29250 = ~n29246 & n29249;
  assign n29251 = ~n29245 & n29250;
  assign n29252 = ~n29239 & ~n29251;
  assign n29253 = ~n29238 & ~n29239;
  assign n29254 = ~n29251 & n29253;
  assign n29255 = ~n29238 & ~n29254;
  assign n29256 = ~n29238 & ~n29252;
  assign n29257 = n29011 & ~n56871;
  assign n29258 = ~n29011 & n56871;
  assign n29259 = ~n29257 & ~n29258;
  assign n29260 = n11279 & ~n56721;
  assign n29261 = n12584 & n26286;
  assign n29262 = n54410 & n26292;
  assign n29263 = n11267 & n26289;
  assign n29264 = ~n29262 & ~n29263;
  assign n29265 = ~n29261 & n29264;
  assign n29266 = ~n11279 & n29265;
  assign n29267 = n56721 & n29265;
  assign n29268 = ~n29266 & ~n29267;
  assign n29269 = ~n29260 & n29265;
  assign n29270 = pi29  & ~n56872;
  assign n29271 = ~pi29  & n56872;
  assign n29272 = ~n29270 & ~n29271;
  assign n29273 = n29259 & ~n29272;
  assign n29274 = ~n29257 & ~n29273;
  assign n29275 = n28829 & n56814;
  assign n29276 = ~n28837 & ~n29275;
  assign n29277 = ~n29274 & n29276;
  assign n29278 = n29274 & ~n29276;
  assign n29279 = n123 & ~n56648;
  assign n29280 = n128 & n26274;
  assign n29281 = n53444 & n26280;
  assign n29282 = n127 & n26277;
  assign n29283 = ~n29281 & ~n29282;
  assign n29284 = ~n29280 & n29283;
  assign n29285 = ~n29279 & n29284;
  assign n29286 = pi26  & ~n29285;
  assign n29287 = pi26  & ~n29286;
  assign n29288 = pi26  & n29285;
  assign n29289 = ~n29285 & ~n29286;
  assign n29290 = ~pi26  & ~n29285;
  assign n29291 = ~n56873 & ~n56874;
  assign n29292 = ~n29278 & ~n29291;
  assign n29293 = ~n29277 & ~n29278;
  assign n29294 = ~n29291 & n29293;
  assign n29295 = ~n29277 & ~n29294;
  assign n29296 = ~n29277 & ~n29292;
  assign n29297 = ~n56848 & ~n56875;
  assign n29298 = ~n29002 & ~n29297;
  assign n29299 = n28883 & ~n28885;
  assign n29300 = n28885 & ~n28886;
  assign n29301 = ~n28883 & ~n28886;
  assign n29302 = ~n29300 & ~n29301;
  assign n29303 = ~n28886 & ~n29299;
  assign n29304 = ~n29298 & ~n56876;
  assign n29305 = n29298 & n56876;
  assign n29306 = n90 & ~n56639;
  assign n29307 = n14236 & n26259;
  assign n29308 = n54667 & n26265;
  assign n29309 = n14210 & n26262;
  assign n29310 = ~n29308 & ~n29309;
  assign n29311 = ~n29307 & n29310;
  assign n29312 = ~n29306 & n29311;
  assign n29313 = pi23  & ~n29312;
  assign n29314 = pi23  & ~n29313;
  assign n29315 = pi23  & n29312;
  assign n29316 = ~n29312 & ~n29313;
  assign n29317 = ~pi23  & ~n29312;
  assign n29318 = ~n56877 & ~n56878;
  assign n29319 = ~n29305 & ~n29318;
  assign n29320 = ~n29304 & ~n29305;
  assign n29321 = ~n29318 & n29320;
  assign n29322 = ~n29304 & ~n29321;
  assign n29323 = ~n29304 & ~n29319;
  assign n29324 = ~n56842 & ~n56879;
  assign n29325 = n56842 & n56879;
  assign n29326 = n14413 & ~n56567;
  assign n29327 = n15921 & n26247;
  assign n29328 = n54719 & n26253;
  assign n29329 = n15901 & n26250;
  assign n29330 = ~n29328 & ~n29329;
  assign n29331 = ~n29327 & n29330;
  assign n29332 = ~n29326 & n29331;
  assign n29333 = pi20  & ~n29332;
  assign n29334 = pi20  & ~n29333;
  assign n29335 = pi20  & n29332;
  assign n29336 = ~n29332 & ~n29333;
  assign n29337 = ~pi20  & ~n29332;
  assign n29338 = ~n56880 & ~n56881;
  assign n29339 = ~n29325 & ~n29338;
  assign n29340 = ~n29324 & ~n29325;
  assign n29341 = ~n29338 & n29340;
  assign n29342 = ~n29324 & ~n29341;
  assign n29343 = ~n29324 & ~n29339;
  assign n29344 = ~n56841 & ~n56882;
  assign n29345 = ~n28971 & ~n29344;
  assign n29346 = n28932 & ~n28934;
  assign n29347 = n28934 & ~n28935;
  assign n29348 = ~n28932 & ~n28935;
  assign n29349 = ~n29347 & ~n29348;
  assign n29350 = ~n28935 & ~n29346;
  assign n29351 = ~n29345 & ~n56883;
  assign n29352 = n29345 & n56883;
  assign n29353 = n54886 & ~n26537;
  assign n29354 = ~n16676 & ~n29353;
  assign n29355 = ~n16696 & n29354;
  assign n29356 = ~n16696 & ~n29353;
  assign n29357 = ~n16676 & n29356;
  assign n29358 = n26870 & ~n29353;
  assign n29359 = ~n16079 & n56884;
  assign n29360 = pi17  & ~n29359;
  assign n29361 = pi17  & ~n29360;
  assign n29362 = pi17  & n29359;
  assign n29363 = ~n29359 & ~n29360;
  assign n29364 = ~pi17  & ~n29359;
  assign n29365 = ~n56885 & ~n56886;
  assign n29366 = ~n29352 & ~n29365;
  assign n29367 = ~n29351 & ~n29352;
  assign n29368 = ~n29365 & n29367;
  assign n29369 = ~n29351 & ~n29368;
  assign n29370 = ~n29351 & ~n29366;
  assign n29371 = ~n56836 & ~n56887;
  assign n29372 = n56836 & n56887;
  assign n29373 = ~n29371 & ~n29372;
  assign n29374 = n16079 & n28624;
  assign n29375 = n16676 & ~n26537;
  assign n29376 = n54886 & n26242;
  assign n29377 = ~n16696 & ~n29376;
  assign n29378 = ~n29375 & ~n29376;
  assign n29379 = ~n16696 & n29378;
  assign n29380 = ~n29375 & n29377;
  assign n29381 = ~n29374 & n56888;
  assign n29382 = pi17  & ~n29381;
  assign n29383 = pi17  & ~n29382;
  assign n29384 = pi17  & n29381;
  assign n29385 = ~n29381 & ~n29382;
  assign n29386 = ~pi17  & ~n29381;
  assign n29387 = ~n56889 & ~n56890;
  assign n29388 = n29338 & ~n29340;
  assign n29389 = n29340 & ~n29341;
  assign n29390 = ~n29338 & ~n29341;
  assign n29391 = ~n29389 & ~n29390;
  assign n29392 = ~n29341 & ~n29388;
  assign n29393 = n56848 & n56875;
  assign n29394 = ~n29297 & ~n29393;
  assign n29395 = n90 & n27466;
  assign n29396 = n14236 & n26262;
  assign n29397 = n54667 & n26268;
  assign n29398 = n14210 & n26265;
  assign n29399 = ~n29397 & ~n29398;
  assign n29400 = ~n29396 & n29399;
  assign n29401 = ~n29395 & n29400;
  assign n29402 = pi23  & ~n29401;
  assign n29403 = pi23  & ~n29402;
  assign n29404 = pi23  & n29401;
  assign n29405 = ~n29401 & ~n29402;
  assign n29406 = ~pi23  & ~n29401;
  assign n29407 = ~n56892 & ~n56893;
  assign n29408 = n29394 & ~n29407;
  assign n29409 = ~n29394 & n29407;
  assign n29410 = n29394 & ~n29408;
  assign n29411 = n29394 & n29407;
  assign n29412 = ~n29407 & ~n29408;
  assign n29413 = ~n29394 & ~n29407;
  assign n29414 = ~n56894 & ~n56895;
  assign n29415 = ~n29408 & ~n29409;
  assign n29416 = n29291 & ~n29293;
  assign n29417 = n29293 & ~n29294;
  assign n29418 = ~n29291 & ~n29294;
  assign n29419 = ~n29417 & ~n29418;
  assign n29420 = ~n29294 & ~n29416;
  assign n29421 = n11279 & n28107;
  assign n29422 = n12584 & n26289;
  assign n29423 = n54410 & n26295;
  assign n29424 = n11267 & n26292;
  assign n29425 = ~n29423 & ~n29424;
  assign n29426 = ~n29422 & n29425;
  assign n29427 = ~n29421 & n29426;
  assign n29428 = pi29  & ~n29427;
  assign n29429 = pi29  & ~n29428;
  assign n29430 = pi29  & n29427;
  assign n29431 = ~n29427 & ~n29428;
  assign n29432 = ~pi29  & ~n29427;
  assign n29433 = ~n56898 & ~n56899;
  assign n29434 = n29251 & ~n29253;
  assign n29435 = n29253 & ~n29254;
  assign n29436 = ~n29251 & ~n29254;
  assign n29437 = ~n29435 & ~n29436;
  assign n29438 = ~n29254 & ~n29434;
  assign n29439 = ~n29433 & ~n56900;
  assign n29440 = n29229 & ~n29231;
  assign n29441 = ~n29229 & ~n56869;
  assign n29442 = ~n29230 & n29235;
  assign n29443 = ~n29441 & ~n29442;
  assign n29444 = ~n56869 & ~n29440;
  assign n29445 = n26427 & ~n26429;
  assign n29446 = ~n26430 & ~n29445;
  assign n29447 = n1576 & n29446;
  assign n29448 = n11215 & n26301;
  assign n29449 = n54403 & n26307;
  assign n29450 = n10564 & n26304;
  assign n29451 = ~n29449 & ~n29450;
  assign n29452 = ~n29448 & n29451;
  assign n29453 = ~n29447 & n29452;
  assign n29454 = ~n56901 & ~n29453;
  assign n29455 = n8265 & n8860;
  assign n29456 = n12275 & n13217;
  assign n29457 = n29455 & n29456;
  assign n29458 = ~n354 & ~n361;
  assign n29459 = ~n506 & ~n948;
  assign n29460 = n29458 & n29459;
  assign n29461 = n3950 & n7755;
  assign n29462 = n29460 & n29461;
  assign n29463 = n7755 & n8265;
  assign n29464 = n8860 & n13217;
  assign n29465 = n29463 & n29464;
  assign n29466 = ~n354 & ~n441;
  assign n29467 = ~n182 & ~n506;
  assign n29468 = n29466 & n29467;
  assign n29469 = ~n361 & ~n948;
  assign n29470 = n3950 & n29469;
  assign n29471 = n29468 & n29470;
  assign n29472 = n29465 & n29471;
  assign n29473 = ~n174 & ~n948;
  assign n29474 = n8860 & n29473;
  assign n29475 = n29461 & n29474;
  assign n29476 = ~n361 & ~n506;
  assign n29477 = n29466 & n29476;
  assign n29478 = ~n182 & ~n340;
  assign n29479 = n8265 & n29478;
  assign n29480 = n29477 & n29479;
  assign n29481 = n29475 & n29480;
  assign n29482 = n29457 & n29462;
  assign n29483 = n53523 & n54307;
  assign n29484 = n56902 & n29483;
  assign n29485 = n54374 & n29484;
  assign n29486 = n53662 & n29485;
  assign n29487 = n53523 & n8860;
  assign n29488 = n7755 & n29487;
  assign n29489 = n53662 & n29488;
  assign n29490 = n54435 & n29489;
  assign n29491 = n54374 & n29490;
  assign n29492 = n54307 & n29491;
  assign n29493 = n3950 & n29492;
  assign n29494 = ~n948 & n29493;
  assign n29495 = ~n174 & n29494;
  assign n29496 = ~n182 & n29495;
  assign n29497 = ~n441 & n29496;
  assign n29498 = ~n268 & n29497;
  assign n29499 = ~n506 & n29498;
  assign n29500 = ~n340 & n29499;
  assign n29501 = ~n361 & n29500;
  assign n29502 = ~n354 & n29501;
  assign n29503 = ~n646 & n29502;
  assign n29504 = n54435 & n29486;
  assign n29505 = n56855 & ~n56903;
  assign n29506 = ~n1081 & n1716;
  assign n29507 = n1716 & n27077;
  assign n29508 = ~n1081 & n29507;
  assign n29509 = n27077 & n29506;
  assign n29510 = n7307 & n8052;
  assign n29511 = n13164 & n26692;
  assign n29512 = n29510 & n29511;
  assign n29513 = n53598 & n29512;
  assign n29514 = n56904 & n29513;
  assign n29515 = ~n751 & ~n1535;
  assign n29516 = n421 & n29515;
  assign n29517 = n4378 & n6310;
  assign n29518 = n29516 & n29517;
  assign n29519 = n323 & n7955;
  assign n29520 = n29518 & n29519;
  assign n29521 = n53844 & n29520;
  assign n29522 = n53516 & n29521;
  assign n29523 = n8052 & n13164;
  assign n29524 = n6310 & n7307;
  assign n29525 = n29523 & n29524;
  assign n29526 = n53598 & n29525;
  assign n29527 = n56904 & n29526;
  assign n29528 = n4378 & n29515;
  assign n29529 = n421 & n26692;
  assign n29530 = n29528 & n29529;
  assign n29531 = n29519 & n29530;
  assign n29532 = n53844 & n29531;
  assign n29533 = n53516 & n29532;
  assign n29534 = n29527 & n29533;
  assign n29535 = n322 & n7307;
  assign n29536 = n29523 & n29535;
  assign n29537 = n53598 & n29536;
  assign n29538 = n56904 & n29537;
  assign n29539 = n421 & n4378;
  assign n29540 = n7955 & n29539;
  assign n29541 = ~n1535 & n6310;
  assign n29542 = ~n319 & ~n614;
  assign n29543 = ~n751 & ~n773;
  assign n29544 = n29542 & n29543;
  assign n29545 = n29541 & n29544;
  assign n29546 = n29540 & n29545;
  assign n29547 = n53844 & n29546;
  assign n29548 = n53516 & n29547;
  assign n29549 = n29538 & n29548;
  assign n29550 = n29514 & n29522;
  assign n29551 = n53598 & n56904;
  assign n29552 = n7307 & n29551;
  assign n29553 = n56860 & n29552;
  assign n29554 = n53844 & n29553;
  assign n29555 = n4585 & n29554;
  assign n29556 = n8052 & n29555;
  assign n29557 = n1067 & n29556;
  assign n29558 = n4378 & n29557;
  assign n29559 = n53516 & n29558;
  assign n29560 = n322 & n29559;
  assign n29561 = n421 & n29560;
  assign n29562 = n13164 & n29561;
  assign n29563 = ~n1044 & n29562;
  assign n29564 = ~n215 & n29563;
  assign n29565 = ~n1535 & n29564;
  assign n29566 = ~n319 & n29565;
  assign n29567 = ~n773 & n29566;
  assign n29568 = ~n751 & n29567;
  assign n29569 = ~n614 & n29568;
  assign n29570 = n56860 & n56905;
  assign n29571 = n56855 & ~n56906;
  assign n29572 = ~n56855 & n56906;
  assign n29573 = ~n29571 & ~n29572;
  assign n29574 = n6309 & n9510;
  assign n29575 = n11547 & n29574;
  assign n29576 = ~n423 & ~n1034;
  assign n29577 = ~n1034 & ~n1195;
  assign n29578 = ~n423 & n29577;
  assign n29579 = ~n1195 & n29576;
  assign n29580 = n1578 & n4259;
  assign n29581 = n56907 & n29580;
  assign n29582 = n53519 & n54458;
  assign n29583 = n29581 & n29582;
  assign n29584 = n4259 & n6309;
  assign n29585 = n1578 & n29584;
  assign n29586 = ~n310 & n29577;
  assign n29587 = ~n423 & ~n510;
  assign n29588 = n9510 & n29587;
  assign n29589 = n29586 & n29588;
  assign n29590 = n29582 & n29589;
  assign n29591 = n29585 & n29590;
  assign n29592 = n29575 & n29583;
  assign n29593 = ~n316 & ~n789;
  assign n29594 = ~n1079 & n29593;
  assign n29595 = ~n271 & ~n591;
  assign n29596 = n6860 & n29595;
  assign n29597 = n8823 & n29596;
  assign n29598 = ~n316 & ~n1079;
  assign n29599 = n6860 & n29598;
  assign n29600 = n6860 & n8823;
  assign n29601 = ~n316 & n29600;
  assign n29602 = ~n1079 & n29601;
  assign n29603 = n8823 & n29599;
  assign n29604 = ~n271 & n56909;
  assign n29605 = ~n591 & n29604;
  assign n29606 = ~n789 & n29605;
  assign n29607 = ~n591 & ~n789;
  assign n29608 = ~n1079 & n29607;
  assign n29609 = ~n271 & ~n316;
  assign n29610 = n6860 & n29609;
  assign n29611 = n8823 & n29610;
  assign n29612 = n29608 & n29611;
  assign n29613 = ~n271 & ~n789;
  assign n29614 = ~n591 & n29613;
  assign n29615 = n56909 & n29614;
  assign n29616 = n29594 & n29597;
  assign n29617 = n54092 & n56910;
  assign n29618 = n9510 & n29584;
  assign n29619 = n54458 & n29618;
  assign n29620 = n53519 & n29619;
  assign n29621 = n54092 & n29620;
  assign n29622 = n56910 & n29621;
  assign n29623 = n1578 & n29622;
  assign n29624 = ~n1195 & n29623;
  assign n29625 = ~n310 & n29624;
  assign n29626 = ~n1034 & n29625;
  assign n29627 = ~n510 & n29626;
  assign n29628 = ~n423 & n29627;
  assign n29629 = n56908 & n29617;
  assign n29630 = ~n340 & ~n447;
  assign n29631 = ~n340 & ~n1472;
  assign n29632 = ~n447 & n29631;
  assign n29633 = ~n1472 & n29630;
  assign n29634 = n1802 & n7275;
  assign n29635 = ~n447 & ~n1062;
  assign n29636 = ~n1457 & n29635;
  assign n29637 = n7275 & n29631;
  assign n29638 = n29636 & n29637;
  assign n29639 = n56912 & n29634;
  assign n29640 = n7275 & n56911;
  assign n29641 = ~n1062 & n29640;
  assign n29642 = ~n1472 & n29641;
  assign n29643 = ~n1457 & n29642;
  assign n29644 = ~n340 & n29643;
  assign n29645 = ~n447 & n29644;
  assign n29646 = n56911 & n56913;
  assign n29647 = ~n163 & ~n1646;
  assign n29648 = ~n1044 & n29647;
  assign n29649 = n11830 & n17873;
  assign n29650 = ~n496 & ~n1192;
  assign n29651 = ~n922 & n29650;
  assign n29652 = ~n1044 & ~n1646;
  assign n29653 = ~n163 & ~n1681;
  assign n29654 = n29652 & n29653;
  assign n29655 = n29651 & n29654;
  assign n29656 = n29648 & n29649;
  assign n29657 = ~n922 & n53686;
  assign n29658 = ~n1044 & n29657;
  assign n29659 = ~n1192 & n29658;
  assign n29660 = ~n1681 & n29659;
  assign n29661 = ~n163 & n29660;
  assign n29662 = ~n1646 & n29661;
  assign n29663 = ~n496 & n29662;
  assign n29664 = n53686 & n56915;
  assign n29665 = ~n294 & ~n361;
  assign n29666 = ~n1065 & n29665;
  assign n29667 = ~n108 & ~n166;
  assign n29668 = n4529 & n29667;
  assign n29669 = ~n1065 & n29667;
  assign n29670 = n4529 & n29665;
  assign n29671 = n29669 & n29670;
  assign n29672 = n29666 & n29668;
  assign n29673 = n54035 & n56726;
  assign n29674 = n56917 & n29673;
  assign n29675 = ~n956 & ~n1492;
  assign n29676 = n6482 & n10182;
  assign n29677 = n29675 & n29676;
  assign n29678 = n54096 & n29677;
  assign n29679 = ~n108 & ~n294;
  assign n29680 = ~n166 & n29679;
  assign n29681 = ~n361 & ~n1065;
  assign n29682 = n6482 & n29681;
  assign n29683 = n29680 & n29682;
  assign n29684 = n29673 & n29683;
  assign n29685 = n4529 & n10182;
  assign n29686 = n29675 & n29685;
  assign n29687 = n54096 & n29686;
  assign n29688 = n29684 & n29687;
  assign n29689 = ~n166 & ~n1492;
  assign n29690 = ~n956 & n29689;
  assign n29691 = ~n294 & ~n1065;
  assign n29692 = ~n108 & ~n361;
  assign n29693 = n29691 & n29692;
  assign n29694 = n29690 & n29693;
  assign n29695 = n29673 & n29694;
  assign n29696 = n4529 & n6482;
  assign n29697 = n10182 & n29696;
  assign n29698 = n54096 & n29697;
  assign n29699 = n29695 & n29698;
  assign n29700 = n29674 & n29678;
  assign n29701 = n56916 & n56918;
  assign n29702 = n56608 & n29701;
  assign n29703 = n4529 & n54035;
  assign n29704 = n10182 & n29703;
  assign n29705 = n54096 & n29704;
  assign n29706 = n56916 & n29705;
  assign n29707 = n56608 & n29706;
  assign n29708 = n56914 & n29707;
  assign n29709 = n56726 & n29708;
  assign n29710 = n6482 & n29709;
  assign n29711 = ~n1065 & n29710;
  assign n29712 = ~n1492 & n29711;
  assign n29713 = ~n108 & n29712;
  assign n29714 = ~n294 & n29713;
  assign n29715 = ~n166 & n29714;
  assign n29716 = ~n956 & n29715;
  assign n29717 = ~n361 & n29716;
  assign n29718 = n56914 & n29702;
  assign n29719 = n56855 & ~n56919;
  assign n29720 = ~n56855 & n56919;
  assign n29721 = n26399 & ~n26401;
  assign n29722 = ~n26399 & ~n56549;
  assign n29723 = ~n26400 & n26405;
  assign n29724 = ~n29722 & ~n29723;
  assign n29725 = ~n56549 & ~n29721;
  assign n29726 = n1576 & ~n56920;
  assign n29727 = n11215 & n26316;
  assign n29728 = n54403 & n26322;
  assign n29729 = n10564 & n26319;
  assign n29730 = ~n29728 & ~n29729;
  assign n29731 = ~n29727 & n29730;
  assign n29732 = ~n29726 & n29731;
  assign n29733 = ~n29720 & ~n29732;
  assign n29734 = ~n29719 & ~n29720;
  assign n29735 = ~n29719 & n29733;
  assign n29736 = ~n29719 & ~n29732;
  assign n29737 = ~n29720 & n29736;
  assign n29738 = ~n29732 & n29734;
  assign n29739 = ~n29719 & ~n56921;
  assign n29740 = ~n29719 & ~n29733;
  assign n29741 = ~n29572 & ~n56922;
  assign n29742 = ~n29571 & n29741;
  assign n29743 = n29573 & ~n56922;
  assign n29744 = ~n29571 & ~n56923;
  assign n29745 = ~n56855 & n56903;
  assign n29746 = ~n29505 & ~n29745;
  assign n29747 = ~n29744 & ~n29745;
  assign n29748 = ~n29505 & n29747;
  assign n29749 = ~n29744 & n29746;
  assign n29750 = ~n29505 & ~n56924;
  assign n29751 = ~n29200 & n56865;
  assign n29752 = ~n56865 & ~n56866;
  assign n29753 = ~n29199 & ~n56866;
  assign n29754 = ~n29198 & n29753;
  assign n29755 = n29200 & ~n56866;
  assign n29756 = ~n29752 & ~n56925;
  assign n29757 = ~n56866 & ~n29751;
  assign n29758 = ~n29750 & ~n56926;
  assign n29759 = n29750 & n56926;
  assign n29760 = ~n29750 & n56926;
  assign n29761 = n29750 & ~n56926;
  assign n29762 = ~n29760 & ~n29761;
  assign n29763 = ~n29758 & ~n29759;
  assign n29764 = n26415 & ~n26417;
  assign n29765 = ~n26415 & ~n56551;
  assign n29766 = ~n26416 & n26421;
  assign n29767 = ~n29765 & ~n29766;
  assign n29768 = ~n56551 & ~n29764;
  assign n29769 = n1576 & ~n56928;
  assign n29770 = n11215 & n26307;
  assign n29771 = n54403 & n26313;
  assign n29772 = n10564 & n26310;
  assign n29773 = ~n29771 & ~n29772;
  assign n29774 = ~n29770 & n29773;
  assign n29775 = ~n29769 & n29774;
  assign n29776 = ~n56927 & ~n29775;
  assign n29777 = ~n29758 & ~n29776;
  assign n29778 = ~n29212 & n56868;
  assign n29779 = ~n29228 & ~n29778;
  assign n29780 = ~n29777 & n29779;
  assign n29781 = n29777 & ~n29779;
  assign n29782 = ~n29780 & ~n29781;
  assign n29783 = n11279 & n28493;
  assign n29784 = n12584 & n26295;
  assign n29785 = n54410 & n26301;
  assign n29786 = n11267 & n26298;
  assign n29787 = ~n29785 & ~n29786;
  assign n29788 = ~n29784 & n29787;
  assign n29789 = ~n11279 & n29788;
  assign n29790 = ~n28493 & n29788;
  assign n29791 = ~n29789 & ~n29790;
  assign n29792 = ~n29783 & n29788;
  assign n29793 = pi29  & ~n56929;
  assign n29794 = ~pi29  & n56929;
  assign n29795 = ~n29793 & ~n29794;
  assign n29796 = n29782 & ~n29795;
  assign n29797 = ~n29780 & ~n29796;
  assign n29798 = n56901 & n29453;
  assign n29799 = ~n56901 & ~n29454;
  assign n29800 = ~n56901 & n29453;
  assign n29801 = ~n29453 & ~n29454;
  assign n29802 = n56901 & ~n29453;
  assign n29803 = ~n56930 & ~n56931;
  assign n29804 = ~n29454 & ~n29798;
  assign n29805 = ~n29797 & ~n56932;
  assign n29806 = ~n29454 & ~n29805;
  assign n29807 = n29433 & n56900;
  assign n29808 = ~n56900 & ~n29439;
  assign n29809 = ~n29433 & ~n29439;
  assign n29810 = ~n29808 & ~n29809;
  assign n29811 = ~n29439 & ~n29807;
  assign n29812 = ~n29806 & ~n56933;
  assign n29813 = ~n29439 & ~n29812;
  assign n29814 = ~n29259 & n29272;
  assign n29815 = ~n29273 & ~n29814;
  assign n29816 = ~n29813 & n29815;
  assign n29817 = n29813 & ~n29815;
  assign n29818 = n123 & n27330;
  assign n29819 = n128 & n26277;
  assign n29820 = n53444 & n26283;
  assign n29821 = n127 & n26280;
  assign n29822 = ~n29820 & ~n29821;
  assign n29823 = ~n29819 & n29822;
  assign n29824 = ~n29818 & n29823;
  assign n29825 = pi26  & ~n29824;
  assign n29826 = pi26  & ~n29825;
  assign n29827 = pi26  & n29824;
  assign n29828 = ~n29824 & ~n29825;
  assign n29829 = ~pi26  & ~n29824;
  assign n29830 = ~n56934 & ~n56935;
  assign n29831 = ~n29817 & ~n29830;
  assign n29832 = ~n29816 & ~n29817;
  assign n29833 = ~n29830 & n29832;
  assign n29834 = ~n29816 & ~n29833;
  assign n29835 = ~n29816 & ~n29831;
  assign n29836 = ~n56897 & ~n56936;
  assign n29837 = n56897 & n56936;
  assign n29838 = n90 & n27042;
  assign n29839 = n14236 & n26265;
  assign n29840 = n54667 & n26271;
  assign n29841 = n14210 & n26268;
  assign n29842 = ~n29840 & ~n29841;
  assign n29843 = ~n29839 & n29842;
  assign n29844 = ~n29838 & n29843;
  assign n29845 = pi23  & ~n29844;
  assign n29846 = pi23  & ~n29845;
  assign n29847 = pi23  & n29844;
  assign n29848 = ~n29844 & ~n29845;
  assign n29849 = ~pi23  & ~n29844;
  assign n29850 = ~n56937 & ~n56938;
  assign n29851 = ~n29837 & ~n29850;
  assign n29852 = ~n29836 & ~n29837;
  assign n29853 = ~n29850 & n29852;
  assign n29854 = ~n29836 & ~n29853;
  assign n29855 = ~n29836 & ~n29851;
  assign n29856 = ~n56896 & ~n56939;
  assign n29857 = ~n29408 & ~n29856;
  assign n29858 = n29320 & ~n29321;
  assign n29859 = n29318 & n29320;
  assign n29860 = ~n29318 & ~n29321;
  assign n29861 = ~n29318 & ~n29320;
  assign n29862 = n29318 & ~n29320;
  assign n29863 = ~n29321 & ~n29862;
  assign n29864 = ~n56940 & ~n56941;
  assign n29865 = ~n29857 & n56942;
  assign n29866 = n29857 & ~n56942;
  assign n29867 = n14413 & n27491;
  assign n29868 = n15921 & n26250;
  assign n29869 = n54719 & n26256;
  assign n29870 = n15901 & n26253;
  assign n29871 = ~n29869 & ~n29870;
  assign n29872 = ~n29868 & n29871;
  assign n29873 = ~n29867 & n29872;
  assign n29874 = pi20  & ~n29873;
  assign n29875 = pi20  & ~n29874;
  assign n29876 = pi20  & n29873;
  assign n29877 = ~n29873 & ~n29874;
  assign n29878 = ~pi20  & ~n29873;
  assign n29879 = ~n56943 & ~n56944;
  assign n29880 = ~n29866 & ~n29879;
  assign n29881 = ~n29865 & ~n29866;
  assign n29882 = ~n29879 & n29881;
  assign n29883 = ~n29865 & ~n29882;
  assign n29884 = ~n29865 & ~n29880;
  assign n29885 = ~n56891 & ~n56945;
  assign n29886 = n56891 & n56945;
  assign n29887 = n16079 & ~n56564;
  assign n29888 = n16696 & ~n26537;
  assign n29889 = n54886 & n26244;
  assign n29890 = n16676 & n26242;
  assign n29891 = ~n29889 & ~n29890;
  assign n29892 = ~n29888 & n29891;
  assign n29893 = ~n29887 & n29892;
  assign n29894 = pi17  & ~n29893;
  assign n29895 = pi17  & ~n29894;
  assign n29896 = pi17  & n29893;
  assign n29897 = ~n29893 & ~n29894;
  assign n29898 = ~pi17  & ~n29893;
  assign n29899 = ~n56946 & ~n56947;
  assign n29900 = ~n29886 & ~n29899;
  assign n29901 = ~n29885 & ~n29886;
  assign n29902 = ~n29899 & n29901;
  assign n29903 = ~n29885 & ~n29902;
  assign n29904 = ~n29885 & ~n29900;
  assign n29905 = ~n29387 & ~n56948;
  assign n29906 = n56841 & n56882;
  assign n29907 = ~n29344 & ~n29906;
  assign n29908 = n29387 & n56948;
  assign n29909 = ~n56948 & ~n29905;
  assign n29910 = n29387 & ~n56948;
  assign n29911 = ~n29387 & ~n29905;
  assign n29912 = ~n29387 & n56948;
  assign n29913 = ~n56949 & ~n56950;
  assign n29914 = ~n29905 & ~n29908;
  assign n29915 = n29907 & ~n56951;
  assign n29916 = ~n29905 & ~n29915;
  assign n29917 = n29367 & ~n29368;
  assign n29918 = n29365 & n29367;
  assign n29919 = ~n29365 & ~n29368;
  assign n29920 = ~n29365 & ~n29367;
  assign n29921 = n29365 & ~n29367;
  assign n29922 = ~n29368 & ~n29921;
  assign n29923 = ~n56952 & ~n56953;
  assign n29924 = ~n29916 & n56954;
  assign n29925 = ~n29907 & n56951;
  assign n29926 = ~n29915 & ~n29925;
  assign n29927 = n56896 & n56939;
  assign n29928 = ~n29856 & ~n29927;
  assign n29929 = n14413 & ~n56668;
  assign n29930 = n15921 & n26253;
  assign n29931 = n54719 & n26259;
  assign n29932 = n15901 & n26256;
  assign n29933 = ~n29931 & ~n29932;
  assign n29934 = ~n29930 & n29933;
  assign n29935 = ~n29929 & n29934;
  assign n29936 = pi20  & ~n29935;
  assign n29937 = pi20  & ~n29936;
  assign n29938 = pi20  & n29935;
  assign n29939 = ~n29935 & ~n29936;
  assign n29940 = ~pi20  & ~n29935;
  assign n29941 = ~n56955 & ~n56956;
  assign n29942 = n29928 & ~n29941;
  assign n29943 = ~n29928 & n29941;
  assign n29944 = n29928 & ~n29942;
  assign n29945 = n29928 & n29941;
  assign n29946 = ~n29941 & ~n29942;
  assign n29947 = ~n29928 & ~n29941;
  assign n29948 = ~n56957 & ~n56958;
  assign n29949 = ~n29942 & ~n29943;
  assign n29950 = n29850 & ~n29852;
  assign n29951 = n29852 & ~n29853;
  assign n29952 = ~n29850 & ~n29853;
  assign n29953 = ~n29951 & ~n29952;
  assign n29954 = ~n29853 & ~n29950;
  assign n29955 = n29806 & n56933;
  assign n29956 = ~n29812 & ~n29955;
  assign n29957 = n123 & n27743;
  assign n29958 = n128 & n26280;
  assign n29959 = n53444 & n26286;
  assign n29960 = n127 & n26283;
  assign n29961 = ~n29959 & ~n29960;
  assign n29962 = ~n29958 & n29961;
  assign n29963 = ~n29957 & n29962;
  assign n29964 = pi26  & ~n29963;
  assign n29965 = pi26  & ~n29964;
  assign n29966 = pi26  & n29963;
  assign n29967 = ~n29963 & ~n29964;
  assign n29968 = ~pi26  & ~n29963;
  assign n29969 = ~n56961 & ~n56962;
  assign n29970 = n29956 & ~n29969;
  assign n29971 = n29797 & n56932;
  assign n29972 = ~n29805 & ~n29971;
  assign n29973 = n11279 & n28808;
  assign n29974 = n12584 & n26292;
  assign n29975 = n54410 & n26298;
  assign n29976 = n11267 & n26295;
  assign n29977 = ~n29975 & ~n29976;
  assign n29978 = ~n29974 & n29977;
  assign n29979 = ~n29973 & n29978;
  assign n29980 = pi29  & ~n29979;
  assign n29981 = pi29  & ~n29980;
  assign n29982 = pi29  & n29979;
  assign n29983 = ~n29979 & ~n29980;
  assign n29984 = ~pi29  & ~n29979;
  assign n29985 = ~n56963 & ~n56964;
  assign n29986 = n29972 & ~n29985;
  assign n29987 = n123 & ~n56686;
  assign n29988 = n128 & n26283;
  assign n29989 = n53444 & n26289;
  assign n29990 = n127 & n26286;
  assign n29991 = ~n29989 & ~n29990;
  assign n29992 = ~n29988 & n29991;
  assign n29993 = ~n29987 & n29992;
  assign n29994 = pi26  & ~n29993;
  assign n29995 = pi26  & ~n29994;
  assign n29996 = pi26  & n29993;
  assign n29997 = ~n29993 & ~n29994;
  assign n29998 = ~pi26  & ~n29993;
  assign n29999 = ~n56965 & ~n56966;
  assign n30000 = ~n29972 & n29985;
  assign n30001 = n29972 & ~n29986;
  assign n30002 = n29972 & n29985;
  assign n30003 = ~n29985 & ~n29986;
  assign n30004 = ~n29972 & ~n29985;
  assign n30005 = ~n56967 & ~n56968;
  assign n30006 = ~n29986 & ~n30000;
  assign n30007 = ~n29999 & ~n56969;
  assign n30008 = ~n29986 & ~n30007;
  assign n30009 = ~n29956 & n29969;
  assign n30010 = n29956 & ~n29970;
  assign n30011 = n29956 & n29969;
  assign n30012 = ~n29969 & ~n29970;
  assign n30013 = ~n29956 & ~n29969;
  assign n30014 = ~n56970 & ~n56971;
  assign n30015 = ~n29970 & ~n30009;
  assign n30016 = ~n30008 & ~n56972;
  assign n30017 = ~n29970 & ~n30016;
  assign n30018 = n29830 & ~n29832;
  assign n30019 = n29832 & ~n29833;
  assign n30020 = ~n29830 & ~n29833;
  assign n30021 = ~n30019 & ~n30020;
  assign n30022 = ~n29833 & ~n30018;
  assign n30023 = ~n30017 & ~n56973;
  assign n30024 = n30017 & n56973;
  assign n30025 = n90 & ~n56601;
  assign n30026 = n14236 & n26268;
  assign n30027 = n54667 & n26274;
  assign n30028 = n14210 & n26271;
  assign n30029 = ~n30027 & ~n30028;
  assign n30030 = ~n30026 & n30029;
  assign n30031 = ~n30025 & n30030;
  assign n30032 = pi23  & ~n30031;
  assign n30033 = pi23  & ~n30032;
  assign n30034 = pi23  & n30031;
  assign n30035 = ~n30031 & ~n30032;
  assign n30036 = ~pi23  & ~n30031;
  assign n30037 = ~n56974 & ~n56975;
  assign n30038 = ~n30024 & ~n30037;
  assign n30039 = ~n30023 & ~n30024;
  assign n30040 = ~n30037 & n30039;
  assign n30041 = ~n30023 & ~n30040;
  assign n30042 = ~n30023 & ~n30038;
  assign n30043 = ~n56960 & ~n56976;
  assign n30044 = n56960 & n56976;
  assign n30045 = n14413 & n27387;
  assign n30046 = n15921 & n26256;
  assign n30047 = n54719 & n26262;
  assign n30048 = n15901 & n26259;
  assign n30049 = ~n30047 & ~n30048;
  assign n30050 = ~n30046 & n30049;
  assign n30051 = ~n30045 & n30050;
  assign n30052 = pi20  & ~n30051;
  assign n30053 = pi20  & ~n30052;
  assign n30054 = pi20  & n30051;
  assign n30055 = ~n30051 & ~n30052;
  assign n30056 = ~pi20  & ~n30051;
  assign n30057 = ~n56977 & ~n56978;
  assign n30058 = ~n30044 & ~n30057;
  assign n30059 = ~n30043 & ~n30044;
  assign n30060 = ~n30057 & n30059;
  assign n30061 = ~n30043 & ~n30060;
  assign n30062 = ~n30043 & ~n30058;
  assign n30063 = ~n56959 & ~n56979;
  assign n30064 = ~n29942 & ~n30063;
  assign n30065 = n29879 & ~n29881;
  assign n30066 = n29881 & ~n29882;
  assign n30067 = ~n29879 & ~n29882;
  assign n30068 = ~n30066 & ~n30067;
  assign n30069 = ~n29882 & ~n30065;
  assign n30070 = ~n30064 & ~n56980;
  assign n30071 = n30064 & n56980;
  assign n30072 = n16079 & n27808;
  assign n30073 = n16696 & n26242;
  assign n30074 = n54886 & n26247;
  assign n30075 = n16676 & n26244;
  assign n30076 = ~n30074 & ~n30075;
  assign n30077 = ~n30073 & n30076;
  assign n30078 = ~n30072 & n30077;
  assign n30079 = pi17  & ~n30078;
  assign n30080 = pi17  & ~n30079;
  assign n30081 = pi17  & n30078;
  assign n30082 = ~n30078 & ~n30079;
  assign n30083 = ~pi17  & ~n30078;
  assign n30084 = ~n56981 & ~n56982;
  assign n30085 = ~n30071 & ~n30084;
  assign n30086 = ~n30070 & ~n30071;
  assign n30087 = ~n30084 & n30086;
  assign n30088 = ~n30070 & ~n30087;
  assign n30089 = ~n30070 & ~n30085;
  assign n30090 = ~n27321 & ~n56983;
  assign n30091 = n27321 & n56983;
  assign n30092 = n29899 & ~n29901;
  assign n30093 = n29901 & ~n29902;
  assign n30094 = ~n29899 & ~n29902;
  assign n30095 = ~n30093 & ~n30094;
  assign n30096 = ~n29902 & ~n30092;
  assign n30097 = ~n30091 & ~n56984;
  assign n30098 = ~n30090 & ~n30091;
  assign n30099 = ~n56984 & n30098;
  assign n30100 = ~n30090 & ~n30099;
  assign n30101 = ~n30090 & ~n30097;
  assign n30102 = n29926 & ~n56985;
  assign n30103 = n56984 & ~n30098;
  assign n30104 = ~n56984 & ~n30099;
  assign n30105 = n30098 & ~n30099;
  assign n30106 = ~n30104 & ~n30105;
  assign n30107 = ~n30099 & ~n30103;
  assign n30108 = n56959 & n56979;
  assign n30109 = ~n30063 & ~n30108;
  assign n30110 = n16079 & n27839;
  assign n30111 = n16696 & n26244;
  assign n30112 = n54886 & n26250;
  assign n30113 = n16676 & n26247;
  assign n30114 = ~n30112 & ~n30113;
  assign n30115 = ~n30111 & n30114;
  assign n30116 = ~n30110 & n30115;
  assign n30117 = pi17  & ~n30116;
  assign n30118 = pi17  & ~n30117;
  assign n30119 = pi17  & n30116;
  assign n30120 = ~n30116 & ~n30117;
  assign n30121 = ~pi17  & ~n30116;
  assign n30122 = ~n56987 & ~n56988;
  assign n30123 = n30109 & ~n30122;
  assign n30124 = ~n30109 & n30122;
  assign n30125 = n30109 & ~n30123;
  assign n30126 = n30109 & n30122;
  assign n30127 = ~n30122 & ~n30123;
  assign n30128 = ~n30109 & ~n30122;
  assign n30129 = ~n56989 & ~n56990;
  assign n30130 = ~n30123 & ~n30124;
  assign n30131 = n30057 & ~n30059;
  assign n30132 = n30059 & ~n30060;
  assign n30133 = ~n30057 & ~n30060;
  assign n30134 = ~n30132 & ~n30133;
  assign n30135 = ~n30060 & ~n30131;
  assign n30136 = n30008 & n56972;
  assign n30137 = ~n30016 & ~n30136;
  assign n30138 = n90 & ~n56612;
  assign n30139 = n14236 & n26271;
  assign n30140 = n54667 & n26277;
  assign n30141 = n14210 & n26274;
  assign n30142 = ~n30140 & ~n30141;
  assign n30143 = ~n30139 & n30142;
  assign n30144 = ~n30138 & n30143;
  assign n30145 = pi23  & ~n30144;
  assign n30146 = pi23  & ~n30145;
  assign n30147 = pi23  & n30144;
  assign n30148 = ~n30144 & ~n30145;
  assign n30149 = ~pi23  & ~n30144;
  assign n30150 = ~n56993 & ~n56994;
  assign n30151 = n30137 & ~n30150;
  assign n30152 = ~n30137 & n30150;
  assign n30153 = n30137 & ~n30151;
  assign n30154 = n30137 & n30150;
  assign n30155 = ~n30150 & ~n30151;
  assign n30156 = ~n30137 & ~n30150;
  assign n30157 = ~n56995 & ~n56996;
  assign n30158 = ~n30151 & ~n30152;
  assign n30159 = n29999 & n56969;
  assign n30160 = ~n56969 & ~n30007;
  assign n30161 = n29999 & ~n56969;
  assign n30162 = ~n29999 & ~n30007;
  assign n30163 = ~n29999 & n56969;
  assign n30164 = ~n56998 & ~n56999;
  assign n30165 = ~n30007 & ~n30159;
  assign n30166 = ~n29782 & n29795;
  assign n30167 = ~n29796 & ~n30166;
  assign n30168 = n29744 & ~n29746;
  assign n30169 = ~n29744 & ~n56924;
  assign n30170 = ~n29745 & n29750;
  assign n30171 = ~n30169 & ~n30170;
  assign n30172 = ~n56924 & ~n30168;
  assign n30173 = n26409 & ~n26411;
  assign n30174 = ~n26409 & ~n56550;
  assign n30175 = ~n26410 & n26415;
  assign n30176 = ~n30174 & ~n30175;
  assign n30177 = ~n56550 & ~n30173;
  assign n30178 = n1576 & ~n57002;
  assign n30179 = n11215 & n26310;
  assign n30180 = n54403 & n26316;
  assign n30181 = n10564 & n26313;
  assign n30182 = ~n30180 & ~n30181;
  assign n30183 = ~n30179 & n30182;
  assign n30184 = ~n30178 & n30183;
  assign n30185 = ~n57001 & ~n30184;
  assign n30186 = ~n29573 & n56922;
  assign n30187 = ~n56922 & ~n56923;
  assign n30188 = ~n29572 & n29744;
  assign n30189 = ~n30187 & ~n30188;
  assign n30190 = ~n56923 & ~n30186;
  assign n30191 = n26405 & ~n26407;
  assign n30192 = ~n26408 & ~n30191;
  assign n30193 = n1576 & n30192;
  assign n30194 = n11215 & n26313;
  assign n30195 = n54403 & n26319;
  assign n30196 = n10564 & n26316;
  assign n30197 = ~n30195 & ~n30196;
  assign n30198 = ~n30194 & n30197;
  assign n30199 = ~n30193 & n30198;
  assign n30200 = ~n57003 & ~n30199;
  assign n30201 = n3715 & n4002;
  assign n30202 = n3937 & n10183;
  assign n30203 = n30201 & n30202;
  assign n30204 = n54208 & n30203;
  assign n30205 = n56709 & n30204;
  assign n30206 = ~n553 & ~n1881;
  assign n30207 = ~n1191 & n30206;
  assign n30208 = ~n513 & ~n1881;
  assign n30209 = ~n514 & ~n553;
  assign n30210 = ~n1191 & n30209;
  assign n30211 = n30208 & n30210;
  assign n30212 = ~n513 & ~n553;
  assign n30213 = ~n514 & ~n1881;
  assign n30214 = ~n1191 & n30213;
  assign n30215 = n30212 & n30214;
  assign n30216 = n515 & n30207;
  assign n30217 = ~n1191 & n54417;
  assign n30218 = ~n553 & n30217;
  assign n30219 = ~n514 & n30218;
  assign n30220 = ~n513 & n30219;
  assign n30221 = ~n1881 & n30220;
  assign n30222 = n54417 & n57004;
  assign n30223 = ~n259 & ~n649;
  assign n30224 = ~n1234 & n30223;
  assign n30225 = n54306 & n30224;
  assign n30226 = n10950 & n54496;
  assign n30227 = n54306 & n54496;
  assign n30228 = n10950 & n30224;
  assign n30229 = n30227 & n30228;
  assign n30230 = n30225 & n30226;
  assign n30231 = n57005 & n57006;
  assign n30232 = n2340 & n4002;
  assign n30233 = n3715 & n10183;
  assign n30234 = n30232 & n30233;
  assign n30235 = n54208 & n30234;
  assign n30236 = n56709 & n30235;
  assign n30237 = ~n587 & ~n649;
  assign n30238 = ~n219 & n30237;
  assign n30239 = ~n259 & ~n1234;
  assign n30240 = n3014 & n30239;
  assign n30241 = n30238 & n30240;
  assign n30242 = n30227 & n30241;
  assign n30243 = n57005 & n30242;
  assign n30244 = n30236 & n30243;
  assign n30245 = n30205 & n30231;
  assign n30246 = n53853 & n57007;
  assign n30247 = n10183 & n30227;
  assign n30248 = n54208 & n30247;
  assign n30249 = n3715 & n30248;
  assign n30250 = n53853 & n30249;
  assign n30251 = n54736 & n30250;
  assign n30252 = n56709 & n30251;
  assign n30253 = n57005 & n30252;
  assign n30254 = n4002 & n30253;
  assign n30255 = n2340 & n30254;
  assign n30256 = n3014 & n30255;
  assign n30257 = ~n219 & n30256;
  assign n30258 = ~n259 & n30257;
  assign n30259 = ~n1234 & n30258;
  assign n30260 = ~n587 & n30259;
  assign n30261 = ~n649 & n30260;
  assign n30262 = n54736 & n30246;
  assign n30263 = n26395 & ~n26397;
  assign n30264 = ~n26398 & ~n30263;
  assign n30265 = n1576 & n30264;
  assign n30266 = n11215 & n26319;
  assign n30267 = n10564 & n26322;
  assign n30268 = n54403 & n26325;
  assign n30269 = ~n30267 & ~n30268;
  assign n30270 = ~n30266 & n30269;
  assign n30271 = ~n30265 & ~n30268;
  assign n30272 = ~n30267 & n30271;
  assign n30273 = ~n30266 & n30272;
  assign n30274 = ~n30265 & n30270;
  assign n30275 = ~n57008 & ~n57009;
  assign n30276 = ~n587 & ~n1455;
  assign n30277 = ~n1124 & ~n2201;
  assign n30278 = n30276 & n30277;
  assign n30279 = n1659 & n3252;
  assign n30280 = n4317 & n5952;
  assign n30281 = n30279 & n30280;
  assign n30282 = n3252 & n30277;
  assign n30283 = n1659 & n30276;
  assign n30284 = n30280 & n30283;
  assign n30285 = n30282 & n30284;
  assign n30286 = ~n788 & ~n1124;
  assign n30287 = n30276 & n30286;
  assign n30288 = ~n174 & ~n2201;
  assign n30289 = n4317 & n30288;
  assign n30290 = n1659 & n5952;
  assign n30291 = n30289 & n30290;
  assign n30292 = n30287 & n30291;
  assign n30293 = n30278 & n30281;
  assign n30294 = n10184 & n10301;
  assign n30295 = n12008 & n30294;
  assign n30296 = n54245 & n30295;
  assign n30297 = n57010 & n30296;
  assign n30298 = n54368 & n54990;
  assign n30299 = n30297 & n30298;
  assign n30300 = n53837 & n30299;
  assign n30301 = n5952 & n12008;
  assign n30302 = n10301 & n30301;
  assign n30303 = n10184 & n30302;
  assign n30304 = n54245 & n30303;
  assign n30305 = n54368 & n30304;
  assign n30306 = n54990 & n30305;
  assign n30307 = n53921 & n30306;
  assign n30308 = n53837 & n30307;
  assign n30309 = n4317 & n30308;
  assign n30310 = n1659 & n30309;
  assign n30311 = ~n1124 & n30310;
  assign n30312 = ~n174 & n30311;
  assign n30313 = ~n1455 & n30312;
  assign n30314 = ~n587 & n30313;
  assign n30315 = ~n788 & n30314;
  assign n30316 = ~n2201 & n30315;
  assign n30317 = n53921 & n30300;
  assign n30318 = n26389 & ~n26391;
  assign n30319 = ~n26389 & ~n56548;
  assign n30320 = ~n26390 & n26395;
  assign n30321 = ~n30319 & ~n30320;
  assign n30322 = ~n56548 & ~n30318;
  assign n30323 = n1576 & ~n57012;
  assign n30324 = n11215 & n26322;
  assign n30325 = n10564 & n26325;
  assign n30326 = n54403 & n26328;
  assign n30327 = ~n30325 & ~n30326;
  assign n30328 = ~n30324 & n30327;
  assign n30329 = ~n30323 & ~n30326;
  assign n30330 = ~n30325 & n30329;
  assign n30331 = ~n30324 & n30330;
  assign n30332 = ~n30323 & n30328;
  assign n30333 = ~n57011 & ~n57013;
  assign n30334 = n54042 & n54286;
  assign n30335 = n13598 & n30334;
  assign n30336 = ~n346 & ~n364;
  assign n30337 = n5378 & n30336;
  assign n30338 = n5639 & n7004;
  assign n30339 = n30337 & n30338;
  assign n30340 = ~n460 & ~n977;
  assign n30341 = ~n1491 & n30340;
  assign n30342 = n53454 & n30341;
  assign n30343 = ~n364 & ~n460;
  assign n30344 = n5378 & n30343;
  assign n30345 = n30338 & n30344;
  assign n30346 = ~n346 & ~n977;
  assign n30347 = ~n1491 & n30346;
  assign n30348 = n53454 & n30347;
  assign n30349 = n30345 & n30348;
  assign n30350 = n30339 & n30342;
  assign n30351 = n53454 & n54286;
  assign n30352 = n13598 & n30351;
  assign n30353 = ~n364 & ~n977;
  assign n30354 = n5639 & n30353;
  assign n30355 = n5378 & n7004;
  assign n30356 = n30354 & n30355;
  assign n30357 = ~n346 & ~n1491;
  assign n30358 = ~n460 & n30357;
  assign n30359 = n54042 & n30358;
  assign n30360 = n30356 & n30359;
  assign n30361 = n30352 & n30360;
  assign n30362 = n53454 & n30334;
  assign n30363 = ~n364 & ~n1491;
  assign n30364 = n5378 & n30363;
  assign n30365 = n30338 & n30364;
  assign n30366 = ~n460 & n30346;
  assign n30367 = n13598 & n30366;
  assign n30368 = n30365 & n30367;
  assign n30369 = n30362 & n30368;
  assign n30370 = n30335 & n57014;
  assign n30371 = n54271 & n57015;
  assign n30372 = n54087 & n30371;
  assign n30373 = n7004 & n30351;
  assign n30374 = n54087 & n30373;
  assign n30375 = n54271 & n30374;
  assign n30376 = n56914 & n30375;
  assign n30377 = n5378 & n30376;
  assign n30378 = n54042 & n30377;
  assign n30379 = n13598 & n30378;
  assign n30380 = n5639 & n30379;
  assign n30381 = ~n977 & n30380;
  assign n30382 = ~n1491 & n30381;
  assign n30383 = ~n460 & n30382;
  assign n30384 = ~n364 & n30383;
  assign n30385 = ~n346 & n30384;
  assign n30386 = n56914 & n30372;
  assign n30387 = n26383 & ~n26385;
  assign n30388 = ~n26383 & ~n56547;
  assign n30389 = ~n26384 & n26389;
  assign n30390 = ~n30388 & ~n30389;
  assign n30391 = ~n56547 & ~n30387;
  assign n30392 = n1576 & ~n57017;
  assign n30393 = n11215 & n26325;
  assign n30394 = n10564 & n26328;
  assign n30395 = n54403 & n26331;
  assign n30396 = ~n30394 & ~n30395;
  assign n30397 = ~n30393 & n30396;
  assign n30398 = ~n30392 & ~n30395;
  assign n30399 = ~n30394 & n30398;
  assign n30400 = ~n30393 & n30399;
  assign n30401 = ~n30392 & n30397;
  assign n30402 = ~n57016 & ~n57018;
  assign n30403 = ~n161 & ~n587;
  assign n30404 = ~n172 & ~n422;
  assign n30405 = ~n161 & ~n172;
  assign n30406 = ~n422 & ~n587;
  assign n30407 = n30405 & n30406;
  assign n30408 = ~n161 & ~n422;
  assign n30409 = ~n172 & ~n587;
  assign n30410 = n30408 & n30409;
  assign n30411 = n30403 & n30404;
  assign n30412 = n217 & n755;
  assign n30413 = n57019 & n30412;
  assign n30414 = n54042 & n10686;
  assign n30415 = n30413 & n30414;
  assign n30416 = ~n105 & ~n499;
  assign n30417 = ~n733 & ~n1085;
  assign n30418 = ~n105 & ~n733;
  assign n30419 = ~n499 & ~n1085;
  assign n30420 = n30418 & n30419;
  assign n30421 = ~n105 & ~n1085;
  assign n30422 = ~n499 & ~n733;
  assign n30423 = n30421 & n30422;
  assign n30424 = n30416 & n30417;
  assign n30425 = n421 & n5362;
  assign n30426 = ~n1085 & n30425;
  assign n30427 = ~n105 & n30426;
  assign n30428 = ~n499 & n30427;
  assign n30429 = ~n733 & n30428;
  assign n30430 = n57020 & n30425;
  assign n30431 = n3819 & n6205;
  assign n30432 = n13738 & n30431;
  assign n30433 = n57021 & n30432;
  assign n30434 = n755 & n3819;
  assign n30435 = n57019 & n30434;
  assign n30436 = n30414 & n30435;
  assign n30437 = n217 & n6205;
  assign n30438 = n13738 & n30437;
  assign n30439 = n57021 & n30438;
  assign n30440 = n30436 & n30439;
  assign n30441 = n13738 & n30403;
  assign n30442 = n6205 & n30404;
  assign n30443 = n30441 & n30442;
  assign n30444 = n30414 & n30443;
  assign n30445 = n217 & n30434;
  assign n30446 = n57021 & n30445;
  assign n30447 = n30444 & n30446;
  assign n30448 = n30415 & n30433;
  assign n30449 = n53698 & n54509;
  assign n30450 = n57022 & n30449;
  assign n30451 = n54451 & n30431;
  assign n30452 = n54509 & n30451;
  assign n30453 = n53698 & n30452;
  assign n30454 = n54448 & n30453;
  assign n30455 = n10686 & n30454;
  assign n30456 = n217 & n30455;
  assign n30457 = n54042 & n30456;
  assign n30458 = n755 & n30457;
  assign n30459 = n57021 & n30458;
  assign n30460 = ~n422 & n30459;
  assign n30461 = ~n172 & n30460;
  assign n30462 = ~n161 & n30461;
  assign n30463 = ~n849 & n30462;
  assign n30464 = ~n587 & n30463;
  assign n30465 = ~n360 & n30464;
  assign n30466 = n54448 & n30450;
  assign n30467 = n54451 & n30466;
  assign n30468 = n11761 & n30450;
  assign n30469 = n26379 & ~n26381;
  assign n30470 = ~n26382 & ~n30469;
  assign n30471 = n1576 & n30470;
  assign n30472 = n11215 & n26328;
  assign n30473 = n10564 & n26331;
  assign n30474 = n54403 & n26334;
  assign n30475 = ~n30473 & ~n30474;
  assign n30476 = ~n30472 & n30475;
  assign n30477 = ~n30471 & ~n30474;
  assign n30478 = ~n30473 & n30477;
  assign n30479 = ~n30472 & n30478;
  assign n30480 = ~n30471 & n30476;
  assign n30481 = ~n57023 & ~n57024;
  assign n30482 = n10686 & n54800;
  assign n30483 = n1035 & n1642;
  assign n30484 = n56740 & n30483;
  assign n30485 = n30482 & n30484;
  assign n30486 = n3672 & n8823;
  assign n30487 = n27213 & n30486;
  assign n30488 = ~n750 & ~n771;
  assign n30489 = n775 & n30488;
  assign n30490 = n53460 & n30489;
  assign n30491 = n30487 & n30490;
  assign n30492 = n53455 & n30491;
  assign n30493 = n8823 & n56740;
  assign n30494 = n53460 & n30493;
  assign n30495 = n54800 & n30494;
  assign n30496 = n10686 & n30495;
  assign n30497 = n53455 & n30496;
  assign n30498 = n775 & n30497;
  assign n30499 = n1035 & n30498;
  assign n30500 = n1642 & n30499;
  assign n30501 = n3672 & n30500;
  assign n30502 = ~n408 & n30501;
  assign n30503 = ~n851 & n30502;
  assign n30504 = ~n771 & n30503;
  assign n30505 = ~n750 & n30504;
  assign n30506 = n53460 & n54800;
  assign n30507 = n30484 & n30506;
  assign n30508 = n10686 & n30489;
  assign n30509 = n30487 & n30508;
  assign n30510 = n53455 & n30509;
  assign n30511 = n30507 & n30510;
  assign n30512 = n10686 & n56740;
  assign n30513 = n30506 & n30512;
  assign n30514 = n1035 & n8823;
  assign n30515 = n775 & n30514;
  assign n30516 = n27213 & n30488;
  assign n30517 = n1642 & n3672;
  assign n30518 = n30516 & n30517;
  assign n30519 = n30515 & n30518;
  assign n30520 = n53455 & n30519;
  assign n30521 = n30513 & n30520;
  assign n30522 = n30485 & n30492;
  assign n30523 = ~n354 & ~n565;
  assign n30524 = ~n1490 & n30523;
  assign n30525 = n54017 & n30524;
  assign n30526 = ~n510 & ~n552;
  assign n30527 = ~n552 & ~n1337;
  assign n30528 = ~n510 & n30527;
  assign n30529 = ~n510 & ~n1337;
  assign n30530 = ~n552 & n30529;
  assign n30531 = ~n1337 & n30526;
  assign n30532 = n27664 & n57026;
  assign n30533 = n30525 & n30532;
  assign n30534 = ~n588 & ~n615;
  assign n30535 = n4892 & n30534;
  assign n30536 = n26602 & n30535;
  assign n30537 = n54498 & n30536;
  assign n30538 = ~n565 & ~n588;
  assign n30539 = ~n1490 & n30538;
  assign n30540 = n54017 & n30539;
  assign n30541 = n30532 & n30540;
  assign n30542 = ~n354 & ~n615;
  assign n30543 = n4892 & n30542;
  assign n30544 = n26602 & n30543;
  assign n30545 = n54498 & n30544;
  assign n30546 = n30541 & n30545;
  assign n30547 = n54017 & n57026;
  assign n30548 = ~n354 & ~n588;
  assign n30549 = ~n615 & n30548;
  assign n30550 = ~n565 & ~n1490;
  assign n30551 = n3776 & n30550;
  assign n30552 = n30549 & n30551;
  assign n30553 = n30547 & n30552;
  assign n30554 = n4892 & n13164;
  assign n30555 = n26602 & n30554;
  assign n30556 = n54498 & n30555;
  assign n30557 = n30553 & n30556;
  assign n30558 = ~n565 & n30548;
  assign n30559 = ~n215 & ~n615;
  assign n30560 = ~n1234 & ~n1490;
  assign n30561 = n30559 & n30560;
  assign n30562 = n30558 & n30561;
  assign n30563 = n30547 & n30562;
  assign n30564 = n3776 & n4892;
  assign n30565 = n13164 & n30564;
  assign n30566 = n54498 & n30565;
  assign n30567 = n30563 & n30566;
  assign n30568 = n30533 & n30537;
  assign n30569 = n4892 & n30547;
  assign n30570 = n13164 & n30569;
  assign n30571 = n54498 & n30570;
  assign n30572 = n55115 & n30571;
  assign n30573 = n3776 & n30572;
  assign n30574 = ~n1490 & n30573;
  assign n30575 = ~n215 & n30574;
  assign n30576 = ~n565 & n30575;
  assign n30577 = ~n1234 & n30576;
  assign n30578 = ~n615 & n30577;
  assign n30579 = ~n354 & n30578;
  assign n30580 = ~n588 & n30579;
  assign n30581 = n55115 & n57027;
  assign n30582 = n5874 & n8052;
  assign n30583 = n27260 & n30582;
  assign n30584 = ~n650 & ~n662;
  assign n30585 = ~n340 & ~n879;
  assign n30586 = ~n340 & ~n662;
  assign n30587 = ~n650 & ~n879;
  assign n30588 = n30586 & n30587;
  assign n30589 = ~n662 & ~n879;
  assign n30590 = ~n340 & ~n650;
  assign n30591 = n30589 & n30590;
  assign n30592 = n30584 & n30585;
  assign n30593 = n425 & n57029;
  assign n30594 = n424 & n8052;
  assign n30595 = n27260 & n30594;
  assign n30596 = n421 & n5874;
  assign n30597 = n57029 & n30596;
  assign n30598 = n30595 & n30597;
  assign n30599 = n425 & n8052;
  assign n30600 = ~n507 & ~n650;
  assign n30601 = ~n662 & ~n1195;
  assign n30602 = n30600 & n30601;
  assign n30603 = n5874 & n30585;
  assign n30604 = n30602 & n30603;
  assign n30605 = n30599 & n30604;
  assign n30606 = n30583 & n30593;
  assign n30607 = n53448 & n55091;
  assign n30608 = n57030 & n30607;
  assign n30609 = ~n448 & ~n664;
  assign n30610 = ~n664 & n10951;
  assign n30611 = ~n448 & n30610;
  assign n30612 = n10951 & n30609;
  assign n30613 = n53976 & n54314;
  assign n30614 = n57031 & n30613;
  assign n30615 = n56682 & n30614;
  assign n30616 = n30608 & n30615;
  assign n30617 = n57028 & n30616;
  assign n30618 = n55091 & n30614;
  assign n30619 = n56682 & n30618;
  assign n30620 = n53448 & n30619;
  assign n30621 = n57025 & n30620;
  assign n30622 = n8052 & n30621;
  assign n30623 = n5874 & n30622;
  assign n30624 = n424 & n30623;
  assign n30625 = n421 & n30624;
  assign n30626 = n57028 & n30625;
  assign n30627 = ~n879 & n30626;
  assign n30628 = ~n1195 & n30627;
  assign n30629 = ~n662 & n30628;
  assign n30630 = ~n507 & n30629;
  assign n30631 = ~n340 & n30630;
  assign n30632 = ~n650 & n30631;
  assign n30633 = n57025 & n30616;
  assign n30634 = n57028 & n30633;
  assign n30635 = n57025 & n30617;
  assign n30636 = n26373 & ~n26375;
  assign n30637 = ~n26373 & ~n56546;
  assign n30638 = ~n26374 & n26379;
  assign n30639 = ~n30637 & ~n30638;
  assign n30640 = ~n56546 & ~n30636;
  assign n30641 = n1576 & ~n57033;
  assign n30642 = n11215 & n26331;
  assign n30643 = n10564 & n26334;
  assign n30644 = n54403 & n26337;
  assign n30645 = ~n30643 & ~n30644;
  assign n30646 = ~n30642 & n30645;
  assign n30647 = ~n30641 & ~n30644;
  assign n30648 = ~n30643 & n30647;
  assign n30649 = ~n30642 & n30648;
  assign n30650 = ~n30641 & n30646;
  assign n30651 = ~n57032 & ~n57034;
  assign n30652 = ~n503 & ~n849;
  assign n30653 = ~n957 & ~n1644;
  assign n30654 = ~n503 & ~n957;
  assign n30655 = ~n849 & ~n1644;
  assign n30656 = n30654 & n30655;
  assign n30657 = ~n503 & ~n1644;
  assign n30658 = ~n849 & ~n957;
  assign n30659 = n30657 & n30658;
  assign n30660 = n30652 & n30653;
  assign n30661 = n54388 & n57035;
  assign n30662 = n53615 & n57035;
  assign n30663 = n54388 & n30662;
  assign n30664 = n53615 & n30661;
  assign n30665 = n586 & n1067;
  assign n30666 = n9511 & n30665;
  assign n30667 = n1716 & n3085;
  assign n30668 = n1712 & n5943;
  assign n30669 = n30667 & n30668;
  assign n30670 = n586 & n5943;
  assign n30671 = n9511 & n30670;
  assign n30672 = n1067 & n3085;
  assign n30673 = n1712 & n1716;
  assign n30674 = n30672 & n30673;
  assign n30675 = n30671 & n30674;
  assign n30676 = n30666 & n30669;
  assign n30677 = n57036 & n57037;
  assign n30678 = n53971 & n30677;
  assign n30679 = n53615 & n54388;
  assign n30680 = n56749 & n30679;
  assign n30681 = n3085 & n30680;
  assign n30682 = n1712 & n30681;
  assign n30683 = n53971 & n30682;
  assign n30684 = n1067 & n30683;
  assign n30685 = n5943 & n30684;
  assign n30686 = n586 & n30685;
  assign n30687 = n9511 & n30686;
  assign n30688 = n1716 & n30687;
  assign n30689 = ~n957 & n30688;
  assign n30690 = ~n849 & n30689;
  assign n30691 = ~n1644 & n30690;
  assign n30692 = ~n503 & n30691;
  assign n30693 = n56749 & n30678;
  assign n30694 = n8368 & n9330;
  assign n30695 = n10910 & n16475;
  assign n30696 = n30694 & n30695;
  assign n30697 = n406 & ~n415;
  assign n30698 = n3639 & n5021;
  assign n30699 = n30697 & n30698;
  assign n30700 = n8368 & n16475;
  assign n30701 = n30698 & n30700;
  assign n30702 = ~n415 & n10910;
  assign n30703 = n406 & n9330;
  assign n30704 = n30702 & n30703;
  assign n30705 = n30701 & n30704;
  assign n30706 = n5021 & n9330;
  assign n30707 = n406 & n3639;
  assign n30708 = n30706 & n30707;
  assign n30709 = ~n256 & ~n1490;
  assign n30710 = ~n460 & n30709;
  assign n30711 = ~n274 & ~n415;
  assign n30712 = ~n1031 & ~n1535;
  assign n30713 = n30711 & n30712;
  assign n30714 = n30710 & n30713;
  assign n30715 = n30708 & n30714;
  assign n30716 = n30696 & n30699;
  assign n30717 = n54108 & n57039;
  assign n30718 = n53607 & n30717;
  assign n30719 = n53603 & n30717;
  assign n30720 = n53607 & n30719;
  assign n30721 = n53603 & n30718;
  assign n30722 = n54108 & n9330;
  assign n30723 = n3639 & n30722;
  assign n30724 = n53607 & n30723;
  assign n30725 = n53603 & n30724;
  assign n30726 = n57038 & n30725;
  assign n30727 = n5021 & n30726;
  assign n30728 = n406 & n30727;
  assign n30729 = ~n1031 & n30728;
  assign n30730 = ~n415 & n30729;
  assign n30731 = ~n1490 & n30730;
  assign n30732 = ~n256 & n30731;
  assign n30733 = ~n1535 & n30732;
  assign n30734 = ~n274 & n30733;
  assign n30735 = ~n460 & n30734;
  assign n30736 = n57038 & n57040;
  assign n30737 = n26367 & ~n26369;
  assign n30738 = ~n26367 & ~n56545;
  assign n30739 = ~n26368 & n26373;
  assign n30740 = ~n30738 & ~n30739;
  assign n30741 = ~n56545 & ~n30737;
  assign n30742 = n1576 & ~n57042;
  assign n30743 = n11215 & n26334;
  assign n30744 = n10564 & n26337;
  assign n30745 = n54403 & n26340;
  assign n30746 = ~n30744 & ~n30745;
  assign n30747 = ~n30743 & n30746;
  assign n30748 = ~n30742 & ~n30745;
  assign n30749 = ~n30744 & n30748;
  assign n30750 = ~n30743 & n30749;
  assign n30751 = ~n30742 & n30747;
  assign n30752 = ~n57041 & ~n57043;
  assign n30753 = ~n423 & ~n459;
  assign n30754 = ~n832 & ~n1044;
  assign n30755 = n30753 & n30754;
  assign n30756 = n359 & n30755;
  assign n30757 = n9331 & n30756;
  assign n30758 = ~n514 & n5106;
  assign n30759 = ~n307 & n26757;
  assign n30760 = ~n584 & n30759;
  assign n30761 = ~n514 & n30760;
  assign n30762 = n26757 & n30758;
  assign n30763 = ~n320 & ~n622;
  assign n30764 = n4083 & n30763;
  assign n30765 = n27254 & n30764;
  assign n30766 = n57044 & n30765;
  assign n30767 = ~n320 & ~n423;
  assign n30768 = n30754 & n30767;
  assign n30769 = n359 & n30768;
  assign n30770 = n9331 & n30769;
  assign n30771 = ~n459 & ~n622;
  assign n30772 = n4083 & n30771;
  assign n30773 = n27254 & n30772;
  assign n30774 = n57044 & n30773;
  assign n30775 = n30770 & n30774;
  assign n30776 = ~n423 & ~n622;
  assign n30777 = ~n459 & ~n1044;
  assign n30778 = n30776 & n30777;
  assign n30779 = n9331 & n30778;
  assign n30780 = n359 & n30779;
  assign n30781 = ~n320 & ~n832;
  assign n30782 = n4083 & n30781;
  assign n30783 = n27254 & n30782;
  assign n30784 = n57044 & n30783;
  assign n30785 = n30780 & n30784;
  assign n30786 = ~n292 & ~n832;
  assign n30787 = ~n320 & ~n1044;
  assign n30788 = n30786 & n30787;
  assign n30789 = ~n401 & ~n423;
  assign n30790 = n30771 & n30789;
  assign n30791 = n30788 & n30790;
  assign n30792 = n9331 & n30791;
  assign n30793 = n359 & n4083;
  assign n30794 = n57044 & n30793;
  assign n30795 = n30792 & n30794;
  assign n30796 = n30757 & n30766;
  assign n30797 = ~n628 & ~n1280;
  assign n30798 = ~n1280 & ~n1472;
  assign n30799 = ~n628 & n30798;
  assign n30800 = ~n1472 & n30797;
  assign n30801 = n12286 & n57046;
  assign n30802 = n53689 & n12286;
  assign n30803 = ~n628 & n30802;
  assign n30804 = ~n1472 & n30803;
  assign n30805 = ~n1280 & n30804;
  assign n30806 = n53689 & n30801;
  assign n30807 = n56732 & n57047;
  assign n30808 = n56732 & n57044;
  assign n30809 = n57047 & n30808;
  assign n30810 = n358 & n30809;
  assign n30811 = n4083 & n30810;
  assign n30812 = n9331 & n30811;
  assign n30813 = n355 & n30812;
  assign n30814 = ~n1044 & n30813;
  assign n30815 = ~n320 & n30814;
  assign n30816 = ~n292 & n30815;
  assign n30817 = ~n401 & n30816;
  assign n30818 = ~n459 & n30817;
  assign n30819 = ~n832 & n30818;
  assign n30820 = ~n423 & n30819;
  assign n30821 = ~n622 & n30820;
  assign n30822 = n57045 & n30807;
  assign n30823 = ~n1189 & ~n1680;
  assign n30824 = ~n1491 & ~n1680;
  assign n30825 = ~n1189 & n30824;
  assign n30826 = ~n1491 & n30823;
  assign n30827 = ~n311 & ~n823;
  assign n30828 = n497 & n30827;
  assign n30829 = n57049 & n30828;
  assign n30830 = n53944 & n30829;
  assign n30831 = n1956 & n6150;
  assign n30832 = n8754 & n30831;
  assign n30833 = n53827 & n30832;
  assign n30834 = n54724 & n30833;
  assign n30835 = ~n311 & ~n1189;
  assign n30836 = ~n823 & n30835;
  assign n30837 = n6150 & n30824;
  assign n30838 = n6150 & n30827;
  assign n30839 = n57049 & n30838;
  assign n30840 = n30836 & n30837;
  assign n30841 = n53944 & n57050;
  assign n30842 = n497 & n1956;
  assign n30843 = n497 & n8754;
  assign n30844 = n1956 & n30843;
  assign n30845 = n8754 & n30842;
  assign n30846 = n53827 & n57051;
  assign n30847 = n54724 & n57051;
  assign n30848 = n53827 & n30847;
  assign n30849 = n54724 & n30846;
  assign n30850 = n30841 & n57052;
  assign n30851 = n30830 & n30834;
  assign n30852 = n54214 & n57053;
  assign n30853 = n57048 & n30852;
  assign n30854 = n54040 & n57052;
  assign n30855 = n54214 & n30854;
  assign n30856 = n53944 & n30855;
  assign n30857 = n57048 & n30856;
  assign n30858 = n6150 & n30857;
  assign n30859 = ~n1680 & n30858;
  assign n30860 = ~n1491 & n30859;
  assign n30861 = ~n311 & n30860;
  assign n30862 = ~n1189 & n30861;
  assign n30863 = ~n823 & n30862;
  assign n30864 = n54040 & n30853;
  assign n30865 = n26363 & ~n26365;
  assign n30866 = ~n26366 & ~n30865;
  assign n30867 = n1576 & n30866;
  assign n30868 = n11215 & n26337;
  assign n30869 = n10564 & n26340;
  assign n30870 = n54403 & n26343;
  assign n30871 = ~n30869 & ~n30870;
  assign n30872 = ~n30868 & n30871;
  assign n30873 = ~n30867 & ~n30870;
  assign n30874 = ~n30869 & n30873;
  assign n30875 = ~n30868 & n30874;
  assign n30876 = ~n30867 & n30872;
  assign n30877 = ~n57054 & ~n57055;
  assign n30878 = n53543 & n54295;
  assign n30879 = n55104 & n30878;
  assign n30880 = n217 & n293;
  assign n30881 = n217 & n4884;
  assign n30882 = n293 & n30881;
  assign n30883 = n4884 & n30880;
  assign n30884 = ~n611 & ~n618;
  assign n30885 = ~n1455 & ~n1492;
  assign n30886 = ~n618 & ~n1455;
  assign n30887 = ~n611 & ~n1492;
  assign n30888 = n30886 & n30887;
  assign n30889 = ~n611 & ~n1455;
  assign n30890 = ~n618 & ~n1492;
  assign n30891 = n30889 & n30890;
  assign n30892 = n30884 & n30885;
  assign n30893 = n54510 & n57057;
  assign n30894 = n57056 & n30893;
  assign n30895 = n54831 & n30894;
  assign n30896 = n30879 & n30895;
  assign n30897 = n53534 & n54361;
  assign n30898 = n30896 & n30897;
  assign n30899 = n54295 & n54510;
  assign n30900 = n4884 & n30899;
  assign n30901 = n55104 & n30900;
  assign n30902 = n54831 & n30901;
  assign n30903 = n54507 & n30902;
  assign n30904 = n54361 & n30903;
  assign n30905 = n53534 & n30904;
  assign n30906 = n53543 & n30905;
  assign n30907 = n217 & n30906;
  assign n30908 = n293 & n30907;
  assign n30909 = ~n1492 & n30908;
  assign n30910 = ~n618 & n30909;
  assign n30911 = ~n1455 & n30910;
  assign n30912 = ~n611 & n30911;
  assign n30913 = n54507 & n30898;
  assign n30914 = ~n26346 & n56544;
  assign n30915 = ~n26362 & ~n30914;
  assign n30916 = n1576 & n30915;
  assign n30917 = n11215 & n26340;
  assign n30918 = n10564 & n26343;
  assign n30919 = n54403 & n26348;
  assign n30920 = ~n30918 & ~n30919;
  assign n30921 = ~n30917 & n30920;
  assign n30922 = ~n30916 & ~n30919;
  assign n30923 = ~n30918 & n30922;
  assign n30924 = ~n30917 & n30923;
  assign n30925 = ~n30916 & n30921;
  assign n30926 = ~n57058 & ~n57059;
  assign n30927 = n53540 & n54399;
  assign n30928 = n57021 & n30927;
  assign n30929 = ~n215 & ~n296;
  assign n30930 = ~n215 & ~n1658;
  assign n30931 = ~n296 & n30930;
  assign n30932 = ~n1658 & n30929;
  assign n30933 = ~n207 & ~n409;
  assign n30934 = n8753 & n30933;
  assign n30935 = ~n207 & ~n1658;
  assign n30936 = ~n296 & n30935;
  assign n30937 = ~n215 & ~n409;
  assign n30938 = n8753 & n30937;
  assign n30939 = n30936 & n30938;
  assign n30940 = n57060 & n30934;
  assign n30941 = n53939 & n8753;
  assign n30942 = ~n296 & n30941;
  assign n30943 = ~n215 & n30942;
  assign n30944 = ~n207 & n30943;
  assign n30945 = ~n1658 & n30944;
  assign n30946 = ~n409 & n30945;
  assign n30947 = n53939 & n57061;
  assign n30948 = n355 & n2093;
  assign n30949 = n3273 & n3463;
  assign n30950 = n2093 & n3273;
  assign n30951 = n355 & n3463;
  assign n30952 = n30950 & n30951;
  assign n30953 = n30948 & n30949;
  assign n30954 = ~n166 & ~n405;
  assign n30955 = ~n448 & ~n1769;
  assign n30956 = ~n166 & ~n448;
  assign n30957 = ~n405 & ~n1769;
  assign n30958 = n30956 & n30957;
  assign n30959 = ~n405 & ~n448;
  assign n30960 = ~n166 & ~n1769;
  assign n30961 = n30959 & n30960;
  assign n30962 = n30954 & n30955;
  assign n30963 = n2404 & n57064;
  assign n30964 = n57063 & n30963;
  assign n30965 = n57062 & n30964;
  assign n30966 = n2404 & n3463;
  assign n30967 = n54399 & n30966;
  assign n30968 = n53540 & n30967;
  assign n30969 = n3273 & n30968;
  assign n30970 = n57021 & n30969;
  assign n30971 = n57062 & n30970;
  assign n30972 = n2093 & n30971;
  assign n30973 = n355 & n30972;
  assign n30974 = ~n166 & n30973;
  assign n30975 = ~n405 & n30974;
  assign n30976 = ~n448 & n30975;
  assign n30977 = ~n1769 & n30976;
  assign n30978 = n30928 & n30965;
  assign n30979 = ~n444 & ~n514;
  assign n30980 = ~n514 & ~n1044;
  assign n30981 = ~n444 & n30980;
  assign n30982 = ~n1044 & n30979;
  assign n30983 = n1578 & n6733;
  assign n30984 = n7130 & n8971;
  assign n30985 = n6733 & n8971;
  assign n30986 = n1578 & n7130;
  assign n30987 = n30985 & n30986;
  assign n30988 = n30983 & n30984;
  assign n30989 = n57066 & n57067;
  assign n30990 = n53676 & n54171;
  assign n30991 = n54175 & n54190;
  assign n30992 = n53676 & n54175;
  assign n30993 = n54171 & n54190;
  assign n30994 = n30992 & n30993;
  assign n30995 = n54171 & n54175;
  assign n30996 = n53676 & n54190;
  assign n30997 = n30995 & n30996;
  assign n30998 = n30990 & n30991;
  assign n30999 = n30989 & n57068;
  assign n31000 = n55123 & n30999;
  assign n31001 = n57065 & n31000;
  assign n31002 = n6733 & n7130;
  assign n31003 = n54248 & n31002;
  assign n31004 = n54190 & n31003;
  assign n31005 = n53676 & n31004;
  assign n31006 = n54175 & n31005;
  assign n31007 = n55123 & n31006;
  assign n31008 = n54171 & n31007;
  assign n31009 = n1578 & n31008;
  assign n31010 = n57065 & n31009;
  assign n31011 = ~n1044 & n31010;
  assign n31012 = ~n272 & n31011;
  assign n31013 = ~n1535 & n31012;
  assign n31014 = ~n514 & n31013;
  assign n31015 = ~n444 & n31014;
  assign n31016 = n54248 & n31001;
  assign n31017 = n26348 & n56543;
  assign n31018 = ~n26348 & ~n56543;
  assign n31019 = ~n31017 & ~n31018;
  assign n31020 = n1576 & ~n31019;
  assign n31021 = n11215 & n26348;
  assign n31022 = n10564 & ~n56543;
  assign n31023 = ~n31021 & ~n31022;
  assign n31024 = ~n31020 & ~n31022;
  assign n31025 = ~n31021 & n31024;
  assign n31026 = ~n31020 & n31023;
  assign n31027 = ~n57069 & ~n57070;
  assign n31028 = n5362 & n5733;
  assign n31029 = n814 & n6733;
  assign n31030 = n31028 & n31029;
  assign n31031 = ~n914 & ~n2201;
  assign n31032 = n4697 & n31031;
  assign n31033 = n53877 & n31032;
  assign n31034 = ~n591 & ~n1997;
  assign n31035 = ~n1492 & ~n1997;
  assign n31036 = ~n591 & n31035;
  assign n31037 = ~n1492 & n31034;
  assign n31038 = n12340 & n57071;
  assign n31039 = ~n914 & n26582;
  assign n31040 = ~n753 & ~n2201;
  assign n31041 = n5021 & n31040;
  assign n31042 = n31039 & n31041;
  assign n31043 = n53877 & n57071;
  assign n31044 = n31042 & n31043;
  assign n31045 = n31033 & n31038;
  assign n31046 = n6733 & n57071;
  assign n31047 = n5733 & n31046;
  assign n31048 = n5362 & n31047;
  assign n31049 = n53877 & n31048;
  assign n31050 = n814 & n31049;
  assign n31051 = n5021 & n31050;
  assign n31052 = ~n1065 & n31051;
  assign n31053 = ~n567 & n31052;
  assign n31054 = ~n914 & n31053;
  assign n31055 = ~n753 & n31054;
  assign n31056 = ~n2201 & n31055;
  assign n31057 = n5733 & n6733;
  assign n31058 = n11141 & n11841;
  assign n31059 = n31057 & n31058;
  assign n31060 = n814 & ~n914;
  assign n31061 = n4697 & n5362;
  assign n31062 = n31060 & n31061;
  assign n31063 = n31043 & n31062;
  assign n31064 = n31059 & n31063;
  assign n31065 = n6733 & n11841;
  assign n31066 = n31028 & n31065;
  assign n31067 = ~n914 & n11141;
  assign n31068 = n814 & n4697;
  assign n31069 = n31067 & n31068;
  assign n31070 = n31043 & n31069;
  assign n31071 = n31066 & n31070;
  assign n31072 = n31030 & n57072;
  assign n31073 = ~n1081 & ~n1455;
  assign n31074 = ~n2109 & n31073;
  assign n31075 = n53796 & n31074;
  assign n31076 = n53519 & n53577;
  assign n31077 = n31075 & n31076;
  assign n31078 = n3742 & n4799;
  assign n31079 = n2094 & n31078;
  assign n31080 = ~n272 & ~n553;
  assign n31081 = ~n182 & ~n444;
  assign n31082 = ~n272 & ~n444;
  assign n31083 = ~n182 & ~n553;
  assign n31084 = n31082 & n31083;
  assign n31085 = n31080 & n31081;
  assign n31086 = n1467 & n2694;
  assign n31087 = n57074 & n31086;
  assign n31088 = n31079 & n31087;
  assign n31089 = ~n182 & n31080;
  assign n31090 = n53796 & n31089;
  assign n31091 = n31076 & n31090;
  assign n31092 = n2094 & n4799;
  assign n31093 = n1467 & n4799;
  assign n31094 = n2094 & n31093;
  assign n31095 = n1467 & n31092;
  assign n31096 = ~n444 & ~n2109;
  assign n31097 = n31073 & n31096;
  assign n31098 = n2694 & n3742;
  assign n31099 = n31097 & n31098;
  assign n31100 = n57075 & n31099;
  assign n31101 = n31091 & n31100;
  assign n31102 = ~n1081 & ~n1468;
  assign n31103 = ~n444 & n31102;
  assign n31104 = n53796 & n31103;
  assign n31105 = n31076 & n31104;
  assign n31106 = ~n250 & ~n553;
  assign n31107 = ~n1455 & ~n2109;
  assign n31108 = n31106 & n31107;
  assign n31109 = ~n182 & ~n272;
  assign n31110 = n3742 & n31109;
  assign n31111 = n31108 & n31110;
  assign n31112 = n57075 & n31111;
  assign n31113 = n31105 & n31112;
  assign n31114 = n31077 & n31088;
  assign n31115 = n56916 & n57076;
  assign n31116 = n57073 & n31115;
  assign n31117 = n53577 & n53796;
  assign n31118 = n4799 & n31117;
  assign n31119 = n1467 & n31118;
  assign n31120 = n57073 & n31119;
  assign n31121 = n56730 & n31120;
  assign n31122 = n56916 & n31121;
  assign n31123 = n53519 & n31122;
  assign n31124 = n2094 & n31123;
  assign n31125 = n3742 & n31124;
  assign n31126 = ~n1081 & n31125;
  assign n31127 = ~n1468 & n31126;
  assign n31128 = ~n250 & n31127;
  assign n31129 = ~n272 & n31128;
  assign n31130 = ~n182 & n31129;
  assign n31131 = ~n553 & n31130;
  assign n31132 = ~n1455 & n31131;
  assign n31133 = ~n444 & n31132;
  assign n31134 = ~n2109 & n31133;
  assign n31135 = n56730 & n31116;
  assign n31136 = n31027 & ~n57077;
  assign n31137 = ~n31027 & n57077;
  assign n31138 = n26343 & ~n31017;
  assign n31139 = ~n26343 & n31017;
  assign n31140 = ~n31138 & ~n31139;
  assign n31141 = n1576 & ~n31140;
  assign n31142 = n11215 & n26343;
  assign n31143 = n54403 & ~n56543;
  assign n31144 = n10564 & n26348;
  assign n31145 = ~n31143 & ~n31144;
  assign n31146 = ~n31142 & n31145;
  assign n31147 = ~n31141 & n31146;
  assign n31148 = ~n31137 & ~n31147;
  assign n31149 = ~n31136 & ~n31137;
  assign n31150 = ~n31147 & n31149;
  assign n31151 = ~n31136 & ~n31150;
  assign n31152 = ~n31136 & ~n31148;
  assign n31153 = n57058 & n57059;
  assign n31154 = ~n57058 & ~n30926;
  assign n31155 = ~n57058 & n57059;
  assign n31156 = ~n57059 & ~n30926;
  assign n31157 = n57058 & ~n57059;
  assign n31158 = ~n57079 & ~n57080;
  assign n31159 = ~n30926 & ~n31153;
  assign n31160 = ~n57078 & ~n57081;
  assign n31161 = ~n30926 & ~n31160;
  assign n31162 = n57054 & n57055;
  assign n31163 = ~n57054 & ~n30877;
  assign n31164 = ~n57054 & n57055;
  assign n31165 = ~n57055 & ~n30877;
  assign n31166 = n57054 & ~n57055;
  assign n31167 = ~n57082 & ~n57083;
  assign n31168 = ~n30877 & ~n31162;
  assign n31169 = ~n31161 & ~n57084;
  assign n31170 = ~n30877 & ~n31169;
  assign n31171 = n57041 & n57043;
  assign n31172 = ~n57041 & ~n30752;
  assign n31173 = ~n57041 & n57043;
  assign n31174 = ~n57043 & ~n30752;
  assign n31175 = n57041 & ~n57043;
  assign n31176 = ~n57085 & ~n57086;
  assign n31177 = ~n30752 & ~n31171;
  assign n31178 = ~n31170 & ~n57087;
  assign n31179 = ~n30752 & ~n31178;
  assign n31180 = n57032 & n57034;
  assign n31181 = ~n57032 & ~n30651;
  assign n31182 = ~n57032 & n57034;
  assign n31183 = ~n57034 & ~n30651;
  assign n31184 = n57032 & ~n57034;
  assign n31185 = ~n57088 & ~n57089;
  assign n31186 = ~n30651 & ~n31180;
  assign n31187 = ~n31179 & ~n57090;
  assign n31188 = ~n30651 & ~n31187;
  assign n31189 = n57023 & n57024;
  assign n31190 = ~n57023 & ~n30481;
  assign n31191 = ~n57023 & n57024;
  assign n31192 = ~n57024 & ~n30481;
  assign n31193 = n57023 & ~n57024;
  assign n31194 = ~n57091 & ~n57092;
  assign n31195 = ~n30481 & ~n31189;
  assign n31196 = ~n31188 & ~n57093;
  assign n31197 = ~n30481 & ~n31196;
  assign n31198 = n57016 & n57018;
  assign n31199 = ~n57016 & ~n30402;
  assign n31200 = ~n57016 & n57018;
  assign n31201 = ~n57018 & ~n30402;
  assign n31202 = n57016 & ~n57018;
  assign n31203 = ~n57094 & ~n57095;
  assign n31204 = ~n30402 & ~n31198;
  assign n31205 = ~n31197 & ~n57096;
  assign n31206 = ~n30402 & ~n31205;
  assign n31207 = n57011 & n57013;
  assign n31208 = ~n57011 & ~n30333;
  assign n31209 = ~n57011 & n57013;
  assign n31210 = ~n57013 & ~n30333;
  assign n31211 = n57011 & ~n57013;
  assign n31212 = ~n57097 & ~n57098;
  assign n31213 = ~n30333 & ~n31207;
  assign n31214 = ~n31206 & ~n57099;
  assign n31215 = ~n30333 & ~n31214;
  assign n31216 = n57008 & n57009;
  assign n31217 = ~n57008 & ~n30275;
  assign n31218 = ~n57008 & n57009;
  assign n31219 = ~n57009 & ~n30275;
  assign n31220 = n57008 & ~n57009;
  assign n31221 = ~n57100 & ~n57101;
  assign n31222 = ~n30275 & ~n31216;
  assign n31223 = ~n31215 & ~n57102;
  assign n31224 = ~n30275 & ~n31223;
  assign n31225 = n29732 & ~n29734;
  assign n31226 = ~n29732 & ~n56921;
  assign n31227 = ~n29720 & n56922;
  assign n31228 = ~n31226 & ~n31227;
  assign n31229 = ~n56921 & ~n31225;
  assign n31230 = ~n31224 & ~n57103;
  assign n31231 = n31224 & n57103;
  assign n31232 = ~n31230 & ~n31231;
  assign n31233 = n11279 & ~n56928;
  assign n31234 = n12584 & n26307;
  assign n31235 = n54410 & n26313;
  assign n31236 = n11267 & n26310;
  assign n31237 = ~n31235 & ~n31236;
  assign n31238 = ~n31234 & n31237;
  assign n31239 = ~n11279 & n31238;
  assign n31240 = n56928 & n31238;
  assign n31241 = ~n31239 & ~n31240;
  assign n31242 = ~n31233 & n31238;
  assign n31243 = pi29  & ~n57104;
  assign n31244 = ~pi29  & n57104;
  assign n31245 = ~n31243 & ~n31244;
  assign n31246 = n31232 & ~n31245;
  assign n31247 = ~n31230 & ~n31246;
  assign n31248 = n57003 & n30199;
  assign n31249 = ~n57003 & ~n30200;
  assign n31250 = ~n57003 & n30199;
  assign n31251 = ~n30199 & ~n30200;
  assign n31252 = n57003 & ~n30199;
  assign n31253 = ~n57105 & ~n57106;
  assign n31254 = ~n30200 & ~n31248;
  assign n31255 = ~n31247 & ~n57107;
  assign n31256 = ~n30200 & ~n31255;
  assign n31257 = n57001 & n30184;
  assign n31258 = ~n57001 & ~n30185;
  assign n31259 = ~n57001 & n30184;
  assign n31260 = ~n30184 & ~n30185;
  assign n31261 = n57001 & ~n30184;
  assign n31262 = ~n57108 & ~n57109;
  assign n31263 = ~n30185 & ~n31257;
  assign n31264 = ~n31256 & ~n57110;
  assign n31265 = ~n30185 & ~n31264;
  assign n31266 = n56927 & n29775;
  assign n31267 = ~n29776 & ~n31266;
  assign n31268 = ~n31265 & n31267;
  assign n31269 = n31265 & ~n31267;
  assign n31270 = n11279 & ~n56870;
  assign n31271 = n12584 & n26298;
  assign n31272 = n54410 & n26304;
  assign n31273 = n11267 & n26301;
  assign n31274 = ~n31272 & ~n31273;
  assign n31275 = ~n31271 & n31274;
  assign n31276 = ~n31270 & n31275;
  assign n31277 = pi29  & ~n31276;
  assign n31278 = pi29  & ~n31277;
  assign n31279 = pi29  & n31276;
  assign n31280 = ~n31276 & ~n31277;
  assign n31281 = ~pi29  & ~n31276;
  assign n31282 = ~n57111 & ~n57112;
  assign n31283 = ~n31269 & ~n31282;
  assign n31284 = ~n31268 & ~n31269;
  assign n31285 = ~n31282 & n31284;
  assign n31286 = ~n31268 & ~n31285;
  assign n31287 = ~n31268 & ~n31283;
  assign n31288 = n30167 & ~n57113;
  assign n31289 = ~n30167 & n57113;
  assign n31290 = n123 & ~n56721;
  assign n31291 = n128 & n26286;
  assign n31292 = n53444 & n26292;
  assign n31293 = n127 & n26289;
  assign n31294 = ~n31292 & ~n31293;
  assign n31295 = ~n31291 & n31294;
  assign n31296 = ~n31290 & n31295;
  assign n31297 = pi26  & ~n31296;
  assign n31298 = pi26  & ~n31297;
  assign n31299 = pi26  & n31296;
  assign n31300 = ~n31296 & ~n31297;
  assign n31301 = ~pi26  & ~n31296;
  assign n31302 = ~n57114 & ~n57115;
  assign n31303 = ~n31289 & ~n31302;
  assign n31304 = ~n31288 & ~n31289;
  assign n31305 = ~n31302 & n31304;
  assign n31306 = ~n31288 & ~n31305;
  assign n31307 = ~n31288 & ~n31303;
  assign n31308 = ~n57000 & ~n57116;
  assign n31309 = n57000 & n57116;
  assign n31310 = n90 & ~n56648;
  assign n31311 = n14236 & n26274;
  assign n31312 = n54667 & n26280;
  assign n31313 = n14210 & n26277;
  assign n31314 = ~n31312 & ~n31313;
  assign n31315 = ~n31311 & n31314;
  assign n31316 = ~n31310 & n31315;
  assign n31317 = pi23  & ~n31316;
  assign n31318 = pi23  & ~n31317;
  assign n31319 = pi23  & n31316;
  assign n31320 = ~n31316 & ~n31317;
  assign n31321 = ~pi23  & ~n31316;
  assign n31322 = ~n57117 & ~n57118;
  assign n31323 = ~n31309 & ~n31322;
  assign n31324 = ~n31308 & ~n31309;
  assign n31325 = ~n31322 & n31324;
  assign n31326 = ~n31308 & ~n31325;
  assign n31327 = ~n31308 & ~n31323;
  assign n31328 = ~n56997 & ~n57119;
  assign n31329 = ~n30151 & ~n31328;
  assign n31330 = n30039 & ~n30040;
  assign n31331 = n30037 & n30039;
  assign n31332 = ~n30037 & ~n30040;
  assign n31333 = ~n30037 & ~n30039;
  assign n31334 = n30037 & ~n30039;
  assign n31335 = ~n30040 & ~n31334;
  assign n31336 = ~n57120 & ~n57121;
  assign n31337 = ~n31329 & n57122;
  assign n31338 = n31329 & ~n57122;
  assign n31339 = n14413 & ~n56639;
  assign n31340 = n15921 & n26259;
  assign n31341 = n54719 & n26265;
  assign n31342 = n15901 & n26262;
  assign n31343 = ~n31341 & ~n31342;
  assign n31344 = ~n31340 & n31343;
  assign n31345 = ~n31339 & n31344;
  assign n31346 = pi20  & ~n31345;
  assign n31347 = pi20  & ~n31346;
  assign n31348 = pi20  & n31345;
  assign n31349 = ~n31345 & ~n31346;
  assign n31350 = ~pi20  & ~n31345;
  assign n31351 = ~n57123 & ~n57124;
  assign n31352 = ~n31338 & ~n31351;
  assign n31353 = ~n31337 & ~n31338;
  assign n31354 = ~n31351 & n31353;
  assign n31355 = ~n31337 & ~n31354;
  assign n31356 = ~n31337 & ~n31352;
  assign n31357 = ~n56992 & ~n57125;
  assign n31358 = n56992 & n57125;
  assign n31359 = n16079 & ~n56567;
  assign n31360 = n16696 & n26247;
  assign n31361 = n54886 & n26253;
  assign n31362 = n16676 & n26250;
  assign n31363 = ~n31361 & ~n31362;
  assign n31364 = ~n31360 & n31363;
  assign n31365 = ~n31359 & n31364;
  assign n31366 = pi17  & ~n31365;
  assign n31367 = pi17  & ~n31366;
  assign n31368 = pi17  & n31365;
  assign n31369 = ~n31365 & ~n31366;
  assign n31370 = ~pi17  & ~n31365;
  assign n31371 = ~n57126 & ~n57127;
  assign n31372 = ~n31358 & ~n31371;
  assign n31373 = ~n31357 & ~n31358;
  assign n31374 = ~n31371 & n31373;
  assign n31375 = ~n31357 & ~n31374;
  assign n31376 = ~n31357 & ~n31372;
  assign n31377 = ~n56991 & ~n57128;
  assign n31378 = ~n30123 & ~n31377;
  assign n31379 = n30086 & ~n30087;
  assign n31380 = n30084 & n30086;
  assign n31381 = ~n30084 & ~n30087;
  assign n31382 = ~n30084 & ~n30086;
  assign n31383 = n30084 & ~n30086;
  assign n31384 = ~n30087 & ~n31383;
  assign n31385 = ~n57129 & ~n57130;
  assign n31386 = ~n31378 & n57131;
  assign n31387 = n31378 & ~n57131;
  assign n31388 = n55041 & ~n26537;
  assign n31389 = ~n18556 & ~n31388;
  assign n31390 = ~n18588 & n31389;
  assign n31391 = ~n18588 & ~n31388;
  assign n31392 = ~n18556 & n31391;
  assign n31393 = n27313 & ~n31388;
  assign n31394 = ~n17265 & n57132;
  assign n31395 = pi14  & ~n31394;
  assign n31396 = pi14  & ~n31395;
  assign n31397 = pi14  & n31394;
  assign n31398 = ~n31394 & ~n31395;
  assign n31399 = ~pi14  & ~n31394;
  assign n31400 = ~n57133 & ~n57134;
  assign n31401 = ~n31387 & ~n31400;
  assign n31402 = ~n31386 & ~n31387;
  assign n31403 = ~n31400 & n31402;
  assign n31404 = ~n31386 & ~n31403;
  assign n31405 = ~n31386 & ~n31401;
  assign n31406 = ~n56986 & ~n57135;
  assign n31407 = n56986 & n57135;
  assign n31408 = ~n31406 & ~n31407;
  assign n31409 = n17265 & n28624;
  assign n31410 = n18556 & ~n26537;
  assign n31411 = n55041 & n26242;
  assign n31412 = ~n18588 & ~n31411;
  assign n31413 = ~n31410 & ~n31411;
  assign n31414 = ~n18588 & n31413;
  assign n31415 = ~n31410 & n31412;
  assign n31416 = ~n31409 & n57136;
  assign n31417 = pi14  & ~n31416;
  assign n31418 = pi14  & ~n31417;
  assign n31419 = pi14  & n31416;
  assign n31420 = ~n31416 & ~n31417;
  assign n31421 = ~pi14  & ~n31416;
  assign n31422 = ~n57137 & ~n57138;
  assign n31423 = n31371 & ~n31373;
  assign n31424 = n31373 & ~n31374;
  assign n31425 = ~n31371 & ~n31374;
  assign n31426 = ~n31424 & ~n31425;
  assign n31427 = ~n31374 & ~n31423;
  assign n31428 = n56997 & n57119;
  assign n31429 = ~n31328 & ~n31428;
  assign n31430 = n14413 & n27466;
  assign n31431 = n15921 & n26262;
  assign n31432 = n54719 & n26268;
  assign n31433 = n15901 & n26265;
  assign n31434 = ~n31432 & ~n31433;
  assign n31435 = ~n31431 & n31434;
  assign n31436 = ~n31430 & n31435;
  assign n31437 = pi20  & ~n31436;
  assign n31438 = pi20  & ~n31437;
  assign n31439 = pi20  & n31436;
  assign n31440 = ~n31436 & ~n31437;
  assign n31441 = ~pi20  & ~n31436;
  assign n31442 = ~n57140 & ~n57141;
  assign n31443 = n31429 & ~n31442;
  assign n31444 = ~n31429 & n31442;
  assign n31445 = n31429 & ~n31443;
  assign n31446 = n31429 & n31442;
  assign n31447 = ~n31442 & ~n31443;
  assign n31448 = ~n31429 & ~n31442;
  assign n31449 = ~n57142 & ~n57143;
  assign n31450 = ~n31443 & ~n31444;
  assign n31451 = n31322 & ~n31324;
  assign n31452 = n31324 & ~n31325;
  assign n31453 = ~n31322 & ~n31325;
  assign n31454 = ~n31452 & ~n31453;
  assign n31455 = ~n31325 & ~n31451;
  assign n31456 = n123 & n28107;
  assign n31457 = n128 & n26289;
  assign n31458 = n53444 & n26295;
  assign n31459 = n127 & n26292;
  assign n31460 = ~n31458 & ~n31459;
  assign n31461 = ~n31457 & n31460;
  assign n31462 = ~n31456 & n31461;
  assign n31463 = pi26  & ~n31462;
  assign n31464 = pi26  & ~n31463;
  assign n31465 = pi26  & n31462;
  assign n31466 = ~n31462 & ~n31463;
  assign n31467 = ~pi26  & ~n31462;
  assign n31468 = ~n57146 & ~n57147;
  assign n31469 = n31282 & ~n31284;
  assign n31470 = n31284 & ~n31285;
  assign n31471 = ~n31282 & ~n31285;
  assign n31472 = ~n31470 & ~n31471;
  assign n31473 = ~n31285 & ~n31469;
  assign n31474 = ~n31468 & ~n57148;
  assign n31475 = n31256 & n57110;
  assign n31476 = ~n31264 & ~n31475;
  assign n31477 = n11279 & n29446;
  assign n31478 = n12584 & n26301;
  assign n31479 = n54410 & n26307;
  assign n31480 = n11267 & n26304;
  assign n31481 = ~n31479 & ~n31480;
  assign n31482 = ~n31478 & n31481;
  assign n31483 = ~n31477 & n31482;
  assign n31484 = pi29  & ~n31483;
  assign n31485 = pi29  & ~n31484;
  assign n31486 = pi29  & n31483;
  assign n31487 = ~n31483 & ~n31484;
  assign n31488 = ~pi29  & ~n31483;
  assign n31489 = ~n57149 & ~n57150;
  assign n31490 = n31476 & ~n31489;
  assign n31491 = n123 & n28808;
  assign n31492 = n128 & n26292;
  assign n31493 = n53444 & n26298;
  assign n31494 = n127 & n26295;
  assign n31495 = ~n31493 & ~n31494;
  assign n31496 = ~n31492 & ~n31494;
  assign n31497 = ~n31493 & n31496;
  assign n31498 = ~n31492 & n31495;
  assign n31499 = ~n31491 & n57151;
  assign n31500 = pi26  & ~n31499;
  assign n31501 = pi26  & ~n31500;
  assign n31502 = pi26  & n31499;
  assign n31503 = ~n31499 & ~n31500;
  assign n31504 = ~pi26  & ~n31499;
  assign n31505 = ~n57152 & ~n57153;
  assign n31506 = ~n31476 & n31489;
  assign n31507 = n31476 & ~n31490;
  assign n31508 = n31476 & n31489;
  assign n31509 = ~n31489 & ~n31490;
  assign n31510 = ~n31476 & ~n31489;
  assign n31511 = ~n57154 & ~n57155;
  assign n31512 = ~n31490 & ~n31506;
  assign n31513 = ~n31505 & ~n57156;
  assign n31514 = ~n31490 & ~n31513;
  assign n31515 = n31468 & n57148;
  assign n31516 = ~n57148 & ~n31474;
  assign n31517 = ~n31468 & ~n31474;
  assign n31518 = ~n31516 & ~n31517;
  assign n31519 = ~n31474 & ~n31515;
  assign n31520 = ~n31514 & ~n57157;
  assign n31521 = ~n31474 & ~n31520;
  assign n31522 = n31302 & ~n31304;
  assign n31523 = n31304 & ~n31305;
  assign n31524 = ~n31302 & ~n31305;
  assign n31525 = ~n31523 & ~n31524;
  assign n31526 = ~n31305 & ~n31522;
  assign n31527 = ~n31521 & ~n57158;
  assign n31528 = n31521 & n57158;
  assign n31529 = n90 & n27330;
  assign n31530 = n14236 & n26277;
  assign n31531 = n54667 & n26283;
  assign n31532 = n14210 & n26280;
  assign n31533 = ~n31531 & ~n31532;
  assign n31534 = ~n31530 & n31533;
  assign n31535 = ~n31529 & n31534;
  assign n31536 = pi23  & ~n31535;
  assign n31537 = pi23  & ~n31536;
  assign n31538 = pi23  & n31535;
  assign n31539 = ~n31535 & ~n31536;
  assign n31540 = ~pi23  & ~n31535;
  assign n31541 = ~n57159 & ~n57160;
  assign n31542 = ~n31528 & ~n31541;
  assign n31543 = ~n31527 & ~n31528;
  assign n31544 = ~n31541 & n31543;
  assign n31545 = ~n31527 & ~n31544;
  assign n31546 = ~n31527 & ~n31542;
  assign n31547 = ~n57145 & ~n57161;
  assign n31548 = n57145 & n57161;
  assign n31549 = n14413 & n27042;
  assign n31550 = n15921 & n26265;
  assign n31551 = n54719 & n26271;
  assign n31552 = n15901 & n26268;
  assign n31553 = ~n31551 & ~n31552;
  assign n31554 = ~n31550 & n31553;
  assign n31555 = ~n31549 & n31554;
  assign n31556 = pi20  & ~n31555;
  assign n31557 = pi20  & ~n31556;
  assign n31558 = pi20  & n31555;
  assign n31559 = ~n31555 & ~n31556;
  assign n31560 = ~pi20  & ~n31555;
  assign n31561 = ~n57162 & ~n57163;
  assign n31562 = ~n31548 & ~n31561;
  assign n31563 = ~n31547 & ~n31548;
  assign n31564 = ~n31561 & n31563;
  assign n31565 = ~n31547 & ~n31564;
  assign n31566 = ~n31547 & ~n31562;
  assign n31567 = ~n57144 & ~n57164;
  assign n31568 = ~n31443 & ~n31567;
  assign n31569 = n31351 & ~n31353;
  assign n31570 = n31353 & ~n31354;
  assign n31571 = ~n31351 & ~n31354;
  assign n31572 = ~n31570 & ~n31571;
  assign n31573 = ~n31354 & ~n31569;
  assign n31574 = ~n31568 & ~n57165;
  assign n31575 = n31568 & n57165;
  assign n31576 = n16079 & n27491;
  assign n31577 = n16696 & n26250;
  assign n31578 = n54886 & n26256;
  assign n31579 = n16676 & n26253;
  assign n31580 = ~n31578 & ~n31579;
  assign n31581 = ~n31577 & n31580;
  assign n31582 = ~n31576 & n31581;
  assign n31583 = pi17  & ~n31582;
  assign n31584 = pi17  & ~n31583;
  assign n31585 = pi17  & n31582;
  assign n31586 = ~n31582 & ~n31583;
  assign n31587 = ~pi17  & ~n31582;
  assign n31588 = ~n57166 & ~n57167;
  assign n31589 = ~n31575 & ~n31588;
  assign n31590 = ~n31574 & ~n31575;
  assign n31591 = ~n31588 & n31590;
  assign n31592 = ~n31574 & ~n31591;
  assign n31593 = ~n31574 & ~n31589;
  assign n31594 = ~n57139 & ~n57168;
  assign n31595 = n57139 & n57168;
  assign n31596 = n17265 & ~n56564;
  assign n31597 = n18588 & ~n26537;
  assign n31598 = n55041 & n26244;
  assign n31599 = n18556 & n26242;
  assign n31600 = ~n31598 & ~n31599;
  assign n31601 = ~n31597 & n31600;
  assign n31602 = ~n31596 & n31601;
  assign n31603 = pi14  & ~n31602;
  assign n31604 = pi14  & ~n31603;
  assign n31605 = pi14  & n31602;
  assign n31606 = ~n31602 & ~n31603;
  assign n31607 = ~pi14  & ~n31602;
  assign n31608 = ~n57169 & ~n57170;
  assign n31609 = ~n31595 & ~n31608;
  assign n31610 = ~n31594 & ~n31595;
  assign n31611 = ~n31608 & n31610;
  assign n31612 = ~n31594 & ~n31611;
  assign n31613 = ~n31594 & ~n31609;
  assign n31614 = ~n31422 & ~n57171;
  assign n31615 = n56991 & n57128;
  assign n31616 = ~n31377 & ~n31615;
  assign n31617 = n31422 & n57171;
  assign n31618 = ~n57171 & ~n31614;
  assign n31619 = n31422 & ~n57171;
  assign n31620 = ~n31422 & ~n31614;
  assign n31621 = ~n31422 & n57171;
  assign n31622 = ~n57172 & ~n57173;
  assign n31623 = ~n31614 & ~n31617;
  assign n31624 = n31616 & ~n57174;
  assign n31625 = ~n31614 & ~n31624;
  assign n31626 = n31400 & ~n31402;
  assign n31627 = n31402 & ~n31403;
  assign n31628 = ~n31400 & ~n31403;
  assign n31629 = ~n31627 & ~n31628;
  assign n31630 = ~n31403 & ~n31626;
  assign n31631 = ~n31625 & ~n57175;
  assign n31632 = ~n31616 & n57174;
  assign n31633 = ~n31624 & ~n31632;
  assign n31634 = n57144 & n57164;
  assign n31635 = ~n31567 & ~n31634;
  assign n31636 = n16079 & ~n56668;
  assign n31637 = n16696 & n26253;
  assign n31638 = n54886 & n26259;
  assign n31639 = n16676 & n26256;
  assign n31640 = ~n31638 & ~n31639;
  assign n31641 = ~n31637 & n31640;
  assign n31642 = ~n31636 & n31641;
  assign n31643 = pi17  & ~n31642;
  assign n31644 = pi17  & ~n31643;
  assign n31645 = pi17  & n31642;
  assign n31646 = ~n31642 & ~n31643;
  assign n31647 = ~pi17  & ~n31642;
  assign n31648 = ~n57176 & ~n57177;
  assign n31649 = n31635 & ~n31648;
  assign n31650 = ~n31635 & n31648;
  assign n31651 = n31635 & ~n31649;
  assign n31652 = n31635 & n31648;
  assign n31653 = ~n31648 & ~n31649;
  assign n31654 = ~n31635 & ~n31648;
  assign n31655 = ~n57178 & ~n57179;
  assign n31656 = ~n31649 & ~n31650;
  assign n31657 = n31561 & ~n31563;
  assign n31658 = n31563 & ~n31564;
  assign n31659 = ~n31561 & ~n31564;
  assign n31660 = ~n31658 & ~n31659;
  assign n31661 = ~n31564 & ~n31657;
  assign n31662 = n31514 & n57157;
  assign n31663 = ~n31520 & ~n31662;
  assign n31664 = n90 & n27743;
  assign n31665 = n14236 & n26280;
  assign n31666 = n54667 & n26286;
  assign n31667 = n14210 & n26283;
  assign n31668 = ~n31666 & ~n31667;
  assign n31669 = ~n31665 & n31668;
  assign n31670 = ~n31664 & n31669;
  assign n31671 = pi23  & ~n31670;
  assign n31672 = pi23  & ~n31671;
  assign n31673 = pi23  & n31670;
  assign n31674 = ~n31670 & ~n31671;
  assign n31675 = ~pi23  & ~n31670;
  assign n31676 = ~n57182 & ~n57183;
  assign n31677 = n31663 & ~n31676;
  assign n31678 = ~n31663 & n31676;
  assign n31679 = n31663 & ~n31677;
  assign n31680 = n31663 & n31676;
  assign n31681 = ~n31676 & ~n31677;
  assign n31682 = ~n31663 & ~n31676;
  assign n31683 = ~n57184 & ~n57185;
  assign n31684 = ~n31677 & ~n31678;
  assign n31685 = n31247 & n57107;
  assign n31686 = ~n31255 & ~n31685;
  assign n31687 = n11279 & ~n56867;
  assign n31688 = n12584 & n26304;
  assign n31689 = n54410 & n26310;
  assign n31690 = n11267 & n26307;
  assign n31691 = ~n31689 & ~n31690;
  assign n31692 = ~n31688 & n31691;
  assign n31693 = ~n31687 & n31692;
  assign n31694 = pi29  & ~n31693;
  assign n31695 = pi29  & ~n31694;
  assign n31696 = pi29  & n31693;
  assign n31697 = ~n31693 & ~n31694;
  assign n31698 = ~pi29  & ~n31693;
  assign n31699 = ~n57187 & ~n57188;
  assign n31700 = n31686 & ~n31699;
  assign n31701 = n123 & n28493;
  assign n31702 = n128 & n26295;
  assign n31703 = n127 & n26298;
  assign n31704 = n53444 & n26301;
  assign n31705 = ~n31703 & ~n31704;
  assign n31706 = ~n31702 & ~n31704;
  assign n31707 = ~n31703 & n31706;
  assign n31708 = ~n31702 & n31705;
  assign n31709 = ~n31701 & n57189;
  assign n31710 = pi26  & ~n31709;
  assign n31711 = pi26  & ~n31710;
  assign n31712 = pi26  & n31709;
  assign n31713 = ~n31709 & ~n31710;
  assign n31714 = ~pi26  & ~n31709;
  assign n31715 = ~n57190 & ~n57191;
  assign n31716 = ~n31686 & n31699;
  assign n31717 = n31686 & ~n31700;
  assign n31718 = n31686 & n31699;
  assign n31719 = ~n31699 & ~n31700;
  assign n31720 = ~n31686 & ~n31699;
  assign n31721 = ~n57192 & ~n57193;
  assign n31722 = ~n31700 & ~n31716;
  assign n31723 = ~n31715 & ~n57194;
  assign n31724 = ~n31700 & ~n31723;
  assign n31725 = n31505 & n57156;
  assign n31726 = ~n57156 & ~n31513;
  assign n31727 = n31505 & ~n57156;
  assign n31728 = ~n31505 & ~n31513;
  assign n31729 = ~n31505 & n57156;
  assign n31730 = ~n57195 & ~n57196;
  assign n31731 = ~n31513 & ~n31725;
  assign n31732 = ~n31724 & ~n57197;
  assign n31733 = n31724 & n57197;
  assign n31734 = n90 & ~n56686;
  assign n31735 = n14236 & n26283;
  assign n31736 = n54667 & n26289;
  assign n31737 = n14210 & n26286;
  assign n31738 = ~n31736 & ~n31737;
  assign n31739 = ~n31735 & n31738;
  assign n31740 = ~n31734 & n31739;
  assign n31741 = pi23  & ~n31740;
  assign n31742 = pi23  & ~n31741;
  assign n31743 = pi23  & n31740;
  assign n31744 = ~n31740 & ~n31741;
  assign n31745 = ~pi23  & ~n31740;
  assign n31746 = ~n57198 & ~n57199;
  assign n31747 = ~n31733 & ~n31746;
  assign n31748 = ~n31732 & ~n31733;
  assign n31749 = ~n31746 & n31748;
  assign n31750 = ~n31732 & ~n31749;
  assign n31751 = ~n31732 & ~n31747;
  assign n31752 = ~n57186 & ~n57200;
  assign n31753 = ~n31677 & ~n31752;
  assign n31754 = n31543 & ~n31544;
  assign n31755 = n31541 & n31543;
  assign n31756 = ~n31541 & ~n31544;
  assign n31757 = ~n31541 & ~n31543;
  assign n31758 = n31541 & ~n31543;
  assign n31759 = ~n31544 & ~n31758;
  assign n31760 = ~n57201 & ~n57202;
  assign n31761 = ~n31753 & n57203;
  assign n31762 = n31753 & ~n57203;
  assign n31763 = n14413 & ~n56601;
  assign n31764 = n15921 & n26268;
  assign n31765 = n54719 & n26274;
  assign n31766 = n15901 & n26271;
  assign n31767 = ~n31765 & ~n31766;
  assign n31768 = ~n31764 & n31767;
  assign n31769 = ~n31763 & n31768;
  assign n31770 = pi20  & ~n31769;
  assign n31771 = pi20  & ~n31770;
  assign n31772 = pi20  & n31769;
  assign n31773 = ~n31769 & ~n31770;
  assign n31774 = ~pi20  & ~n31769;
  assign n31775 = ~n57204 & ~n57205;
  assign n31776 = ~n31762 & ~n31775;
  assign n31777 = ~n31761 & ~n31762;
  assign n31778 = ~n31775 & n31777;
  assign n31779 = ~n31761 & ~n31778;
  assign n31780 = ~n31761 & ~n31776;
  assign n31781 = ~n57181 & ~n57206;
  assign n31782 = n57181 & n57206;
  assign n31783 = n16079 & n27387;
  assign n31784 = n16696 & n26256;
  assign n31785 = n54886 & n26262;
  assign n31786 = n16676 & n26259;
  assign n31787 = ~n31785 & ~n31786;
  assign n31788 = ~n31784 & n31787;
  assign n31789 = ~n31783 & n31788;
  assign n31790 = pi17  & ~n31789;
  assign n31791 = pi17  & ~n31790;
  assign n31792 = pi17  & n31789;
  assign n31793 = ~n31789 & ~n31790;
  assign n31794 = ~pi17  & ~n31789;
  assign n31795 = ~n57207 & ~n57208;
  assign n31796 = ~n31782 & ~n31795;
  assign n31797 = ~n31781 & ~n31782;
  assign n31798 = ~n31795 & n31797;
  assign n31799 = ~n31781 & ~n31798;
  assign n31800 = ~n31781 & ~n31796;
  assign n31801 = ~n57180 & ~n57209;
  assign n31802 = ~n31649 & ~n31801;
  assign n31803 = n31590 & ~n31591;
  assign n31804 = n31588 & n31590;
  assign n31805 = ~n31588 & ~n31591;
  assign n31806 = ~n31588 & ~n31590;
  assign n31807 = n31588 & ~n31590;
  assign n31808 = ~n31591 & ~n31807;
  assign n31809 = ~n57210 & ~n57211;
  assign n31810 = ~n31802 & n57212;
  assign n31811 = n31802 & ~n57212;
  assign n31812 = n17265 & n27808;
  assign n31813 = n18588 & n26242;
  assign n31814 = n55041 & n26247;
  assign n31815 = n18556 & n26244;
  assign n31816 = ~n31814 & ~n31815;
  assign n31817 = ~n31813 & n31816;
  assign n31818 = ~n31812 & n31817;
  assign n31819 = pi14  & ~n31818;
  assign n31820 = pi14  & ~n31819;
  assign n31821 = pi14  & n31818;
  assign n31822 = ~n31818 & ~n31819;
  assign n31823 = ~pi14  & ~n31818;
  assign n31824 = ~n57213 & ~n57214;
  assign n31825 = ~n31811 & ~n31824;
  assign n31826 = ~n31810 & ~n31811;
  assign n31827 = ~n31824 & n31826;
  assign n31828 = ~n31810 & ~n31827;
  assign n31829 = ~n31810 & ~n31825;
  assign n31830 = ~n28071 & ~n57215;
  assign n31831 = n28071 & n57215;
  assign n31832 = n31608 & ~n31610;
  assign n31833 = n31610 & ~n31611;
  assign n31834 = ~n31608 & ~n31611;
  assign n31835 = ~n31833 & ~n31834;
  assign n31836 = ~n31611 & ~n31832;
  assign n31837 = ~n31831 & ~n57216;
  assign n31838 = ~n31830 & ~n31831;
  assign n31839 = ~n57216 & n31838;
  assign n31840 = ~n31830 & ~n31839;
  assign n31841 = ~n31830 & ~n31837;
  assign n31842 = n31633 & ~n57217;
  assign n31843 = n57216 & ~n31838;
  assign n31844 = ~n57216 & ~n31839;
  assign n31845 = n31838 & ~n31839;
  assign n31846 = ~n31844 & ~n31845;
  assign n31847 = ~n31839 & ~n31843;
  assign n31848 = n57180 & n57209;
  assign n31849 = ~n31801 & ~n31848;
  assign n31850 = n17265 & n27839;
  assign n31851 = n18588 & n26244;
  assign n31852 = n55041 & n26250;
  assign n31853 = n18556 & n26247;
  assign n31854 = ~n31852 & ~n31853;
  assign n31855 = ~n31851 & n31854;
  assign n31856 = ~n31850 & n31855;
  assign n31857 = pi14  & ~n31856;
  assign n31858 = pi14  & ~n31857;
  assign n31859 = pi14  & n31856;
  assign n31860 = ~n31856 & ~n31857;
  assign n31861 = ~pi14  & ~n31856;
  assign n31862 = ~n57219 & ~n57220;
  assign n31863 = n31849 & ~n31862;
  assign n31864 = ~n31849 & n31862;
  assign n31865 = n31849 & ~n31863;
  assign n31866 = n31849 & n31862;
  assign n31867 = ~n31862 & ~n31863;
  assign n31868 = ~n31849 & ~n31862;
  assign n31869 = ~n57221 & ~n57222;
  assign n31870 = ~n31863 & ~n31864;
  assign n31871 = n31795 & ~n31797;
  assign n31872 = n31797 & ~n31798;
  assign n31873 = ~n31795 & ~n31798;
  assign n31874 = ~n31872 & ~n31873;
  assign n31875 = ~n31798 & ~n31871;
  assign n31876 = n57186 & n57200;
  assign n31877 = ~n31752 & ~n31876;
  assign n31878 = n14413 & ~n56612;
  assign n31879 = n15921 & n26271;
  assign n31880 = n54719 & n26277;
  assign n31881 = n15901 & n26274;
  assign n31882 = ~n31880 & ~n31881;
  assign n31883 = ~n31879 & n31882;
  assign n31884 = ~n31878 & n31883;
  assign n31885 = pi20  & ~n31884;
  assign n31886 = pi20  & ~n31885;
  assign n31887 = pi20  & n31884;
  assign n31888 = ~n31884 & ~n31885;
  assign n31889 = ~pi20  & ~n31884;
  assign n31890 = ~n57225 & ~n57226;
  assign n31891 = n31877 & ~n31890;
  assign n31892 = ~n31877 & n31890;
  assign n31893 = n31877 & ~n31891;
  assign n31894 = n31877 & n31890;
  assign n31895 = ~n31890 & ~n31891;
  assign n31896 = ~n31877 & ~n31890;
  assign n31897 = ~n57227 & ~n57228;
  assign n31898 = ~n31891 & ~n31892;
  assign n31899 = n31746 & ~n31748;
  assign n31900 = n31748 & ~n31749;
  assign n31901 = ~n31746 & ~n31749;
  assign n31902 = ~n31900 & ~n31901;
  assign n31903 = ~n31749 & ~n31899;
  assign n31904 = n31715 & n57194;
  assign n31905 = ~n57194 & ~n31723;
  assign n31906 = n31715 & ~n57194;
  assign n31907 = ~n31715 & ~n31723;
  assign n31908 = ~n31715 & n57194;
  assign n31909 = ~n57231 & ~n57232;
  assign n31910 = ~n31723 & ~n31904;
  assign n31911 = n11279 & ~n57002;
  assign n31912 = n12584 & n26310;
  assign n31913 = n54410 & n26316;
  assign n31914 = n11267 & n26313;
  assign n31915 = ~n31913 & ~n31914;
  assign n31916 = ~n31912 & n31915;
  assign n31917 = ~n11279 & n31916;
  assign n31918 = n57002 & n31916;
  assign n31919 = ~n31917 & ~n31918;
  assign n31920 = ~n31911 & n31916;
  assign n31921 = pi29  & ~n57234;
  assign n31922 = ~pi29  & n57234;
  assign n31923 = ~n31921 & ~n31922;
  assign n31924 = n31215 & n57102;
  assign n31925 = ~n31215 & ~n31223;
  assign n31926 = ~n57102 & ~n31223;
  assign n31927 = ~n31925 & ~n31926;
  assign n31928 = ~n31223 & ~n31924;
  assign n31929 = ~n31923 & ~n57235;
  assign n31930 = n11279 & n30192;
  assign n31931 = n12584 & n26313;
  assign n31932 = n54410 & n26319;
  assign n31933 = n11267 & n26316;
  assign n31934 = ~n31932 & ~n31933;
  assign n31935 = ~n31931 & n31934;
  assign n31936 = ~n11279 & n31935;
  assign n31937 = ~n30192 & n31935;
  assign n31938 = ~n31936 & ~n31937;
  assign n31939 = ~n31930 & n31935;
  assign n31940 = pi29  & ~n57236;
  assign n31941 = ~pi29  & n57236;
  assign n31942 = ~n31940 & ~n31941;
  assign n31943 = n31206 & n57099;
  assign n31944 = ~n31206 & ~n31214;
  assign n31945 = ~n57099 & ~n31214;
  assign n31946 = ~n31944 & ~n31945;
  assign n31947 = ~n31214 & ~n31943;
  assign n31948 = ~n31942 & ~n57237;
  assign n31949 = n11279 & ~n56920;
  assign n31950 = n12584 & n26316;
  assign n31951 = n54410 & n26322;
  assign n31952 = n11267 & n26319;
  assign n31953 = ~n31951 & ~n31952;
  assign n31954 = ~n31950 & n31953;
  assign n31955 = ~n11279 & n31954;
  assign n31956 = n56920 & n31954;
  assign n31957 = ~n31955 & ~n31956;
  assign n31958 = ~n31949 & n31954;
  assign n31959 = pi29  & ~n57238;
  assign n31960 = ~pi29  & n57238;
  assign n31961 = ~n31959 & ~n31960;
  assign n31962 = n31197 & n57096;
  assign n31963 = ~n31197 & ~n31205;
  assign n31964 = ~n57096 & ~n31205;
  assign n31965 = ~n31963 & ~n31964;
  assign n31966 = ~n31205 & ~n31962;
  assign n31967 = ~n31961 & ~n57239;
  assign n31968 = n11279 & n30264;
  assign n31969 = n12584 & n26319;
  assign n31970 = n54410 & n26325;
  assign n31971 = n11267 & n26322;
  assign n31972 = ~n31970 & ~n31971;
  assign n31973 = ~n31969 & n31972;
  assign n31974 = ~n11279 & n31973;
  assign n31975 = ~n30264 & n31973;
  assign n31976 = ~n31974 & ~n31975;
  assign n31977 = ~n31968 & n31973;
  assign n31978 = pi29  & ~n57240;
  assign n31979 = ~pi29  & n57240;
  assign n31980 = ~n31978 & ~n31979;
  assign n31981 = n31188 & n57093;
  assign n31982 = ~n31188 & ~n31196;
  assign n31983 = ~n57093 & ~n31196;
  assign n31984 = ~n31982 & ~n31983;
  assign n31985 = ~n31196 & ~n31981;
  assign n31986 = ~n31980 & ~n57241;
  assign n31987 = n11279 & ~n57012;
  assign n31988 = n12584 & n26322;
  assign n31989 = n54410 & n26328;
  assign n31990 = n11267 & n26325;
  assign n31991 = ~n31989 & ~n31990;
  assign n31992 = ~n31988 & n31991;
  assign n31993 = ~n11279 & n31992;
  assign n31994 = n57012 & n31992;
  assign n31995 = ~n31993 & ~n31994;
  assign n31996 = ~n31987 & n31992;
  assign n31997 = pi29  & ~n57242;
  assign n31998 = ~pi29  & n57242;
  assign n31999 = ~n31997 & ~n31998;
  assign n32000 = n31179 & n57090;
  assign n32001 = ~n31179 & ~n31187;
  assign n32002 = ~n57090 & ~n31187;
  assign n32003 = ~n32001 & ~n32002;
  assign n32004 = ~n31187 & ~n32000;
  assign n32005 = ~n31999 & ~n57243;
  assign n32006 = n11279 & ~n57017;
  assign n32007 = n12584 & n26325;
  assign n32008 = n54410 & n26331;
  assign n32009 = n11267 & n26328;
  assign n32010 = ~n32008 & ~n32009;
  assign n32011 = ~n32007 & n32010;
  assign n32012 = ~n32006 & n32011;
  assign n32013 = pi29  & ~n32012;
  assign n32014 = ~n32012 & ~n32013;
  assign n32015 = ~pi29  & ~n32012;
  assign n32016 = pi29  & ~n32013;
  assign n32017 = pi29  & n32012;
  assign n32018 = ~n57244 & ~n57245;
  assign n32019 = n31170 & n57087;
  assign n32020 = ~n31170 & ~n31178;
  assign n32021 = ~n57087 & ~n31178;
  assign n32022 = ~n32020 & ~n32021;
  assign n32023 = ~n31178 & ~n32019;
  assign n32024 = ~n32018 & ~n57246;
  assign n32025 = n11279 & n30470;
  assign n32026 = n12584 & n26328;
  assign n32027 = n54410 & n26334;
  assign n32028 = n11267 & n26331;
  assign n32029 = ~n32027 & ~n32028;
  assign n32030 = ~n32026 & n32029;
  assign n32031 = ~n32025 & n32030;
  assign n32032 = pi29  & ~n32031;
  assign n32033 = ~n32031 & ~n32032;
  assign n32034 = ~pi29  & ~n32031;
  assign n32035 = pi29  & ~n32032;
  assign n32036 = pi29  & n32031;
  assign n32037 = ~n57247 & ~n57248;
  assign n32038 = n31161 & n57084;
  assign n32039 = ~n31161 & ~n31169;
  assign n32040 = ~n57084 & ~n31169;
  assign n32041 = ~n32039 & ~n32040;
  assign n32042 = ~n31169 & ~n32038;
  assign n32043 = ~n32037 & ~n57249;
  assign n32044 = n11279 & ~n57033;
  assign n32045 = n12584 & n26331;
  assign n32046 = n54410 & n26337;
  assign n32047 = n11267 & n26334;
  assign n32048 = ~n32046 & ~n32047;
  assign n32049 = ~n32045 & n32048;
  assign n32050 = ~n32044 & n32049;
  assign n32051 = pi29  & ~n32050;
  assign n32052 = ~n32050 & ~n32051;
  assign n32053 = ~pi29  & ~n32050;
  assign n32054 = pi29  & ~n32051;
  assign n32055 = pi29  & n32050;
  assign n32056 = ~n57250 & ~n57251;
  assign n32057 = n57078 & n57081;
  assign n32058 = ~n57078 & ~n31160;
  assign n32059 = ~n57081 & ~n31160;
  assign n32060 = ~n32058 & ~n32059;
  assign n32061 = ~n31160 & ~n32057;
  assign n32062 = ~n32056 & ~n57252;
  assign n32063 = n11279 & ~n57042;
  assign n32064 = n12584 & n26334;
  assign n32065 = n54410 & n26340;
  assign n32066 = n11267 & n26337;
  assign n32067 = ~n32065 & ~n32066;
  assign n32068 = ~n32064 & n32067;
  assign n32069 = ~n32063 & n32068;
  assign n32070 = pi29  & ~n32069;
  assign n32071 = ~n32069 & ~n32070;
  assign n32072 = ~pi29  & ~n32069;
  assign n32073 = pi29  & ~n32070;
  assign n32074 = pi29  & n32069;
  assign n32075 = ~n57253 & ~n57254;
  assign n32076 = n31147 & ~n31149;
  assign n32077 = ~n31147 & ~n31150;
  assign n32078 = n31149 & ~n31150;
  assign n32079 = ~n32077 & ~n32078;
  assign n32080 = ~n31150 & ~n32076;
  assign n32081 = ~n32075 & ~n57255;
  assign n32082 = n11279 & n30866;
  assign n32083 = n12584 & n26337;
  assign n32084 = n54410 & n26343;
  assign n32085 = n11267 & n26340;
  assign n32086 = ~n32084 & ~n32085;
  assign n32087 = ~n32083 & n32086;
  assign n32088 = ~n32082 & n32087;
  assign n32089 = pi29  & ~n32088;
  assign n32090 = ~n32088 & ~n32089;
  assign n32091 = ~pi29  & ~n32088;
  assign n32092 = pi29  & ~n32089;
  assign n32093 = pi29  & n32088;
  assign n32094 = ~n57256 & ~n57257;
  assign n32095 = n57069 & n57070;
  assign n32096 = ~n57069 & ~n31027;
  assign n32097 = ~n57069 & n57070;
  assign n32098 = ~n57070 & ~n31027;
  assign n32099 = n57069 & ~n57070;
  assign n32100 = ~n57258 & ~n57259;
  assign n32101 = ~n31027 & ~n32095;
  assign n32102 = ~n32094 & ~n57260;
  assign n32103 = ~n94 & ~n56543;
  assign n32104 = n11279 & ~n31019;
  assign n32105 = n11267 & ~n56543;
  assign n32106 = n12584 & n26348;
  assign n32107 = ~n32105 & ~n32106;
  assign n32108 = ~n32104 & n32107;
  assign n32109 = n54407 & ~n56543;
  assign n32110 = pi29  & ~n32109;
  assign n32111 = pi29  & ~n32108;
  assign n32112 = pi29  & ~n32111;
  assign n32113 = ~n32108 & ~n32111;
  assign n32114 = ~n32112 & ~n32113;
  assign n32115 = n32110 & ~n32114;
  assign n32116 = n32108 & n32110;
  assign n32117 = n11279 & ~n31140;
  assign n32118 = n12584 & n26343;
  assign n32119 = n54410 & ~n56543;
  assign n32120 = n11267 & n26348;
  assign n32121 = ~n32119 & ~n32120;
  assign n32122 = ~n32118 & n32121;
  assign n32123 = ~n11279 & n32122;
  assign n32124 = n31140 & n32122;
  assign n32125 = ~n32123 & ~n32124;
  assign n32126 = ~n32117 & n32122;
  assign n32127 = pi29  & ~n57262;
  assign n32128 = ~pi29  & n57262;
  assign n32129 = ~n32127 & ~n32128;
  assign n32130 = n57261 & ~n32129;
  assign n32131 = n57261 & ~n57262;
  assign n32132 = n32103 & n57263;
  assign n32133 = n11279 & n30915;
  assign n32134 = n12584 & n26340;
  assign n32135 = n54410 & n26348;
  assign n32136 = n11267 & n26343;
  assign n32137 = ~n32135 & ~n32136;
  assign n32138 = ~n32134 & n32137;
  assign n32139 = ~n32133 & n32138;
  assign n32140 = pi29  & ~n32139;
  assign n32141 = ~n32139 & ~n32140;
  assign n32142 = ~pi29  & ~n32139;
  assign n32143 = pi29  & ~n32140;
  assign n32144 = pi29  & n32139;
  assign n32145 = ~n57264 & ~n57265;
  assign n32146 = ~n32103 & ~n57263;
  assign n32147 = ~n32103 & n57263;
  assign n32148 = n32103 & ~n57263;
  assign n32149 = ~n32147 & ~n32148;
  assign n32150 = ~n32132 & ~n32146;
  assign n32151 = ~n32145 & ~n57266;
  assign n32152 = ~n32132 & ~n32151;
  assign n32153 = n32094 & n57260;
  assign n32154 = ~n32094 & ~n32102;
  assign n32155 = ~n57260 & ~n32102;
  assign n32156 = ~n32154 & ~n32155;
  assign n32157 = ~n32102 & ~n32153;
  assign n32158 = ~n32152 & ~n57267;
  assign n32159 = ~n32102 & ~n32158;
  assign n32160 = n32075 & n57255;
  assign n32161 = ~n32075 & ~n32081;
  assign n32162 = ~n57255 & ~n32081;
  assign n32163 = ~n32161 & ~n32162;
  assign n32164 = ~n32081 & ~n32160;
  assign n32165 = ~n32159 & ~n57268;
  assign n32166 = ~n32081 & ~n32165;
  assign n32167 = n32056 & n57252;
  assign n32168 = ~n32056 & ~n32062;
  assign n32169 = ~n32056 & n57252;
  assign n32170 = ~n57252 & ~n32062;
  assign n32171 = n32056 & ~n57252;
  assign n32172 = ~n57269 & ~n57270;
  assign n32173 = ~n32062 & ~n32167;
  assign n32174 = ~n32166 & ~n57271;
  assign n32175 = ~n32062 & ~n32174;
  assign n32176 = n32037 & n57249;
  assign n32177 = ~n32037 & ~n32043;
  assign n32178 = ~n32037 & n57249;
  assign n32179 = ~n57249 & ~n32043;
  assign n32180 = n32037 & ~n57249;
  assign n32181 = ~n57272 & ~n57273;
  assign n32182 = ~n32043 & ~n32176;
  assign n32183 = ~n32175 & ~n57274;
  assign n32184 = ~n32043 & ~n32183;
  assign n32185 = n32018 & n57246;
  assign n32186 = ~n32018 & ~n32024;
  assign n32187 = ~n32018 & n57246;
  assign n32188 = ~n57246 & ~n32024;
  assign n32189 = n32018 & ~n57246;
  assign n32190 = ~n57275 & ~n57276;
  assign n32191 = ~n32024 & ~n32185;
  assign n32192 = ~n32184 & ~n57277;
  assign n32193 = ~n32024 & ~n32192;
  assign n32194 = n31999 & n57243;
  assign n32195 = ~n32005 & ~n32194;
  assign n32196 = ~n32193 & n32195;
  assign n32197 = ~n32005 & ~n32196;
  assign n32198 = n31980 & n57241;
  assign n32199 = ~n31986 & ~n32198;
  assign n32200 = ~n32197 & n32199;
  assign n32201 = ~n31986 & ~n32200;
  assign n32202 = n31961 & n57239;
  assign n32203 = ~n31967 & ~n32202;
  assign n32204 = ~n32201 & n32203;
  assign n32205 = ~n31967 & ~n32204;
  assign n32206 = n31942 & n57237;
  assign n32207 = ~n31948 & ~n32206;
  assign n32208 = ~n32205 & n32207;
  assign n32209 = ~n31948 & ~n32208;
  assign n32210 = n31923 & n57235;
  assign n32211 = ~n31929 & ~n32210;
  assign n32212 = ~n32209 & n32211;
  assign n32213 = ~n31929 & ~n32212;
  assign n32214 = ~n31232 & n31245;
  assign n32215 = ~n31246 & ~n32214;
  assign n32216 = ~n32213 & n32215;
  assign n32217 = n32213 & ~n32215;
  assign n32218 = n123 & ~n56870;
  assign n32219 = n128 & n26298;
  assign n32220 = n53444 & n26304;
  assign n32221 = n127 & n26301;
  assign n32222 = ~n32220 & ~n32221;
  assign n32223 = ~n32219 & n32222;
  assign n32224 = ~n32218 & n32223;
  assign n32225 = pi26  & ~n32224;
  assign n32226 = pi26  & ~n32225;
  assign n32227 = pi26  & n32224;
  assign n32228 = ~n32224 & ~n32225;
  assign n32229 = ~pi26  & ~n32224;
  assign n32230 = ~n57278 & ~n57279;
  assign n32231 = ~n32217 & ~n32230;
  assign n32232 = ~n32216 & ~n32217;
  assign n32233 = ~n32230 & n32232;
  assign n32234 = ~n32216 & ~n32233;
  assign n32235 = ~n32216 & ~n32231;
  assign n32236 = ~n57233 & ~n57280;
  assign n32237 = n57233 & n57280;
  assign n32238 = n90 & ~n56721;
  assign n32239 = n14236 & n26286;
  assign n32240 = n54667 & n26292;
  assign n32241 = n14210 & n26289;
  assign n32242 = ~n32240 & ~n32241;
  assign n32243 = ~n32239 & n32242;
  assign n32244 = ~n32238 & n32243;
  assign n32245 = pi23  & ~n32244;
  assign n32246 = pi23  & ~n32245;
  assign n32247 = pi23  & n32244;
  assign n32248 = ~n32244 & ~n32245;
  assign n32249 = ~pi23  & ~n32244;
  assign n32250 = ~n57281 & ~n57282;
  assign n32251 = ~n32237 & ~n32250;
  assign n32252 = ~n32236 & ~n32237;
  assign n32253 = ~n32250 & n32252;
  assign n32254 = ~n32236 & ~n32253;
  assign n32255 = ~n32236 & ~n32251;
  assign n32256 = ~n57230 & ~n57283;
  assign n32257 = n57230 & n57283;
  assign n32258 = n14413 & ~n56648;
  assign n32259 = n15921 & n26274;
  assign n32260 = n54719 & n26280;
  assign n32261 = n15901 & n26277;
  assign n32262 = ~n32260 & ~n32261;
  assign n32263 = ~n32259 & n32262;
  assign n32264 = ~n32258 & n32263;
  assign n32265 = pi20  & ~n32264;
  assign n32266 = pi20  & ~n32265;
  assign n32267 = pi20  & n32264;
  assign n32268 = ~n32264 & ~n32265;
  assign n32269 = ~pi20  & ~n32264;
  assign n32270 = ~n57284 & ~n57285;
  assign n32271 = ~n32257 & ~n32270;
  assign n32272 = ~n32256 & ~n32257;
  assign n32273 = ~n32270 & n32272;
  assign n32274 = ~n32256 & ~n32273;
  assign n32275 = ~n32256 & ~n32271;
  assign n32276 = ~n57229 & ~n57286;
  assign n32277 = ~n31891 & ~n32276;
  assign n32278 = n31775 & ~n31777;
  assign n32279 = n31777 & ~n31778;
  assign n32280 = ~n31775 & ~n31778;
  assign n32281 = ~n32279 & ~n32280;
  assign n32282 = ~n31778 & ~n32278;
  assign n32283 = ~n32277 & ~n57287;
  assign n32284 = n32277 & n57287;
  assign n32285 = n16079 & ~n56639;
  assign n32286 = n16696 & n26259;
  assign n32287 = n54886 & n26265;
  assign n32288 = n16676 & n26262;
  assign n32289 = ~n32287 & ~n32288;
  assign n32290 = ~n32286 & n32289;
  assign n32291 = ~n32285 & n32290;
  assign n32292 = pi17  & ~n32291;
  assign n32293 = pi17  & ~n32292;
  assign n32294 = pi17  & n32291;
  assign n32295 = ~n32291 & ~n32292;
  assign n32296 = ~pi17  & ~n32291;
  assign n32297 = ~n57288 & ~n57289;
  assign n32298 = ~n32284 & ~n32297;
  assign n32299 = ~n32283 & ~n32284;
  assign n32300 = ~n32297 & n32299;
  assign n32301 = ~n32283 & ~n32300;
  assign n32302 = ~n32283 & ~n32298;
  assign n32303 = ~n57224 & ~n57290;
  assign n32304 = n57224 & n57290;
  assign n32305 = n17265 & ~n56567;
  assign n32306 = n18588 & n26247;
  assign n32307 = n55041 & n26253;
  assign n32308 = n18556 & n26250;
  assign n32309 = ~n32307 & ~n32308;
  assign n32310 = ~n32306 & n32309;
  assign n32311 = ~n32305 & n32310;
  assign n32312 = pi14  & ~n32311;
  assign n32313 = pi14  & ~n32312;
  assign n32314 = pi14  & n32311;
  assign n32315 = ~n32311 & ~n32312;
  assign n32316 = ~pi14  & ~n32311;
  assign n32317 = ~n57291 & ~n57292;
  assign n32318 = ~n32304 & ~n32317;
  assign n32319 = ~n32303 & ~n32304;
  assign n32320 = ~n32317 & n32319;
  assign n32321 = ~n32303 & ~n32320;
  assign n32322 = ~n32303 & ~n32318;
  assign n32323 = ~n57223 & ~n57293;
  assign n32324 = ~n31863 & ~n32323;
  assign n32325 = n31824 & ~n31826;
  assign n32326 = n31826 & ~n31827;
  assign n32327 = ~n31824 & ~n31827;
  assign n32328 = ~n32326 & ~n32327;
  assign n32329 = ~n31827 & ~n32325;
  assign n32330 = ~n32324 & ~n57294;
  assign n32331 = n32324 & n57294;
  assign n32332 = n55247 & ~n26537;
  assign n32333 = ~n19509 & ~n32332;
  assign n32334 = ~n19541 & n32333;
  assign n32335 = ~n19541 & ~n32332;
  assign n32336 = ~n19509 & n32335;
  assign n32337 = n56719 & ~n32332;
  assign n32338 = ~n18846 & n57295;
  assign n32339 = pi11  & ~n32338;
  assign n32340 = pi11  & ~n32339;
  assign n32341 = pi11  & n32338;
  assign n32342 = ~n32338 & ~n32339;
  assign n32343 = ~pi11  & ~n32338;
  assign n32344 = ~n57296 & ~n57297;
  assign n32345 = ~n32331 & ~n32344;
  assign n32346 = ~n32330 & ~n32331;
  assign n32347 = ~n32344 & n32346;
  assign n32348 = ~n32330 & ~n32347;
  assign n32349 = ~n32330 & ~n32345;
  assign n32350 = ~n57218 & ~n57298;
  assign n32351 = n57218 & n57298;
  assign n32352 = ~n32350 & ~n32351;
  assign n32353 = n18846 & n28624;
  assign n32354 = n19509 & ~n26537;
  assign n32355 = n55247 & n26242;
  assign n32356 = ~n19541 & ~n32355;
  assign n32357 = ~n32354 & ~n32355;
  assign n32358 = ~n19541 & n32357;
  assign n32359 = ~n32354 & n32356;
  assign n32360 = ~n32353 & n57299;
  assign n32361 = pi11  & ~n32360;
  assign n32362 = pi11  & ~n32361;
  assign n32363 = pi11  & n32360;
  assign n32364 = ~n32360 & ~n32361;
  assign n32365 = ~pi11  & ~n32360;
  assign n32366 = ~n57300 & ~n57301;
  assign n32367 = n32317 & ~n32319;
  assign n32368 = n32319 & ~n32320;
  assign n32369 = ~n32317 & ~n32320;
  assign n32370 = ~n32368 & ~n32369;
  assign n32371 = ~n32320 & ~n32367;
  assign n32372 = n57229 & n57286;
  assign n32373 = ~n32276 & ~n32372;
  assign n32374 = n16079 & n27466;
  assign n32375 = n16696 & n26262;
  assign n32376 = n54886 & n26268;
  assign n32377 = n16676 & n26265;
  assign n32378 = ~n32376 & ~n32377;
  assign n32379 = ~n32375 & n32378;
  assign n32380 = ~n32374 & n32379;
  assign n32381 = pi17  & ~n32380;
  assign n32382 = pi17  & ~n32381;
  assign n32383 = pi17  & n32380;
  assign n32384 = ~n32380 & ~n32381;
  assign n32385 = ~pi17  & ~n32380;
  assign n32386 = ~n57303 & ~n57304;
  assign n32387 = n32373 & ~n32386;
  assign n32388 = ~n32373 & n32386;
  assign n32389 = n32373 & ~n32387;
  assign n32390 = n32373 & n32386;
  assign n32391 = ~n32386 & ~n32387;
  assign n32392 = ~n32373 & ~n32386;
  assign n32393 = ~n57305 & ~n57306;
  assign n32394 = ~n32387 & ~n32388;
  assign n32395 = n32270 & ~n32272;
  assign n32396 = n32272 & ~n32273;
  assign n32397 = ~n32270 & ~n32273;
  assign n32398 = ~n32396 & ~n32397;
  assign n32399 = ~n32273 & ~n32395;
  assign n32400 = n32250 & ~n32252;
  assign n32401 = n32252 & ~n32253;
  assign n32402 = ~n32250 & ~n32253;
  assign n32403 = ~n32401 & ~n32402;
  assign n32404 = ~n32253 & ~n32400;
  assign n32405 = n32209 & ~n32211;
  assign n32406 = ~n32212 & ~n32405;
  assign n32407 = n123 & n29446;
  assign n32408 = n128 & n26301;
  assign n32409 = n53444 & n26307;
  assign n32410 = n127 & n26304;
  assign n32411 = ~n32409 & ~n32410;
  assign n32412 = ~n32408 & n32411;
  assign n32413 = ~n123 & n32412;
  assign n32414 = ~n29446 & n32412;
  assign n32415 = ~n32413 & ~n32414;
  assign n32416 = ~n32407 & n32412;
  assign n32417 = pi26  & ~n57310;
  assign n32418 = ~pi26  & n57310;
  assign n32419 = ~n32417 & ~n32418;
  assign n32420 = n32406 & ~n32419;
  assign n32421 = n32205 & ~n32207;
  assign n32422 = ~n32208 & ~n32421;
  assign n32423 = n123 & ~n56867;
  assign n32424 = n128 & n26304;
  assign n32425 = n53444 & n26310;
  assign n32426 = n127 & n26307;
  assign n32427 = ~n32425 & ~n32426;
  assign n32428 = ~n32424 & n32427;
  assign n32429 = ~n123 & n32428;
  assign n32430 = n56867 & n32428;
  assign n32431 = ~n32429 & ~n32430;
  assign n32432 = ~n32423 & n32428;
  assign n32433 = pi26  & ~n57311;
  assign n32434 = ~pi26  & n57311;
  assign n32435 = ~n32433 & ~n32434;
  assign n32436 = n32422 & ~n32435;
  assign n32437 = n32201 & ~n32203;
  assign n32438 = ~n32204 & ~n32437;
  assign n32439 = n123 & ~n56928;
  assign n32440 = n128 & n26307;
  assign n32441 = n53444 & n26313;
  assign n32442 = n127 & n26310;
  assign n32443 = ~n32441 & ~n32442;
  assign n32444 = ~n32440 & n32443;
  assign n32445 = ~n123 & n32444;
  assign n32446 = n56928 & n32444;
  assign n32447 = ~n32445 & ~n32446;
  assign n32448 = ~n32439 & n32444;
  assign n32449 = pi26  & ~n57312;
  assign n32450 = ~pi26  & n57312;
  assign n32451 = ~n32449 & ~n32450;
  assign n32452 = n32438 & ~n32451;
  assign n32453 = n32197 & ~n32199;
  assign n32454 = ~n32200 & ~n32453;
  assign n32455 = n123 & ~n57002;
  assign n32456 = n128 & n26310;
  assign n32457 = n53444 & n26316;
  assign n32458 = n127 & n26313;
  assign n32459 = ~n32457 & ~n32458;
  assign n32460 = ~n32456 & n32459;
  assign n32461 = ~n123 & n32460;
  assign n32462 = n57002 & n32460;
  assign n32463 = ~n32461 & ~n32462;
  assign n32464 = ~n32455 & n32460;
  assign n32465 = pi26  & ~n57313;
  assign n32466 = ~pi26  & n57313;
  assign n32467 = ~n32465 & ~n32466;
  assign n32468 = n32454 & ~n32467;
  assign n32469 = n32193 & ~n32195;
  assign n32470 = ~n32196 & ~n32469;
  assign n32471 = n123 & n30192;
  assign n32472 = n128 & n26313;
  assign n32473 = n53444 & n26319;
  assign n32474 = n127 & n26316;
  assign n32475 = ~n32473 & ~n32474;
  assign n32476 = ~n32472 & n32475;
  assign n32477 = ~n123 & n32476;
  assign n32478 = ~n30192 & n32476;
  assign n32479 = ~n32477 & ~n32478;
  assign n32480 = ~n32471 & n32476;
  assign n32481 = pi26  & ~n57314;
  assign n32482 = ~pi26  & n57314;
  assign n32483 = ~n32481 & ~n32482;
  assign n32484 = n32470 & ~n32483;
  assign n32485 = n32184 & n57277;
  assign n32486 = ~n32192 & ~n32485;
  assign n32487 = n123 & ~n56920;
  assign n32488 = n128 & n26316;
  assign n32489 = n53444 & n26322;
  assign n32490 = n127 & n26319;
  assign n32491 = ~n32489 & ~n32490;
  assign n32492 = ~n32488 & n32491;
  assign n32493 = ~n123 & n32492;
  assign n32494 = n56920 & n32492;
  assign n32495 = ~n32493 & ~n32494;
  assign n32496 = ~n32487 & n32492;
  assign n32497 = pi26  & ~n57315;
  assign n32498 = ~pi26  & n57315;
  assign n32499 = ~n32497 & ~n32498;
  assign n32500 = n32486 & ~n32499;
  assign n32501 = n32175 & n57274;
  assign n32502 = ~n32183 & ~n32501;
  assign n32503 = n123 & n30264;
  assign n32504 = n128 & n26319;
  assign n32505 = n53444 & n26325;
  assign n32506 = n127 & n26322;
  assign n32507 = ~n32505 & ~n32506;
  assign n32508 = ~n32504 & ~n32506;
  assign n32509 = ~n32505 & n32508;
  assign n32510 = ~n32504 & n32507;
  assign n32511 = ~n123 & n57316;
  assign n32512 = ~n30264 & n57316;
  assign n32513 = ~n32511 & ~n32512;
  assign n32514 = ~n32503 & n57316;
  assign n32515 = pi26  & ~n57317;
  assign n32516 = ~pi26  & n57317;
  assign n32517 = ~n32515 & ~n32516;
  assign n32518 = n32502 & ~n32517;
  assign n32519 = n32166 & n57271;
  assign n32520 = ~n32174 & ~n32519;
  assign n32521 = n123 & ~n57012;
  assign n32522 = n128 & n26322;
  assign n32523 = n53444 & n26328;
  assign n32524 = n127 & n26325;
  assign n32525 = ~n32523 & ~n32524;
  assign n32526 = ~n32522 & ~n32524;
  assign n32527 = ~n32523 & n32526;
  assign n32528 = ~n32522 & n32525;
  assign n32529 = ~n123 & n57318;
  assign n32530 = n57012 & n57318;
  assign n32531 = ~n32529 & ~n32530;
  assign n32532 = ~n32521 & n57318;
  assign n32533 = pi26  & ~n57319;
  assign n32534 = ~pi26  & n57319;
  assign n32535 = ~n32533 & ~n32534;
  assign n32536 = n32520 & ~n32535;
  assign n32537 = n32159 & n57268;
  assign n32538 = ~n32165 & ~n32537;
  assign n32539 = n123 & ~n57017;
  assign n32540 = n128 & n26325;
  assign n32541 = n127 & n26328;
  assign n32542 = n53444 & n26331;
  assign n32543 = ~n32541 & ~n32542;
  assign n32544 = ~n32540 & ~n32542;
  assign n32545 = ~n32541 & n32544;
  assign n32546 = ~n32540 & n32543;
  assign n32547 = ~n123 & n57320;
  assign n32548 = n57017 & n57320;
  assign n32549 = ~n32547 & ~n32548;
  assign n32550 = ~n32539 & n57320;
  assign n32551 = pi26  & ~n57321;
  assign n32552 = ~pi26  & n57321;
  assign n32553 = ~n32551 & ~n32552;
  assign n32554 = n32538 & ~n32553;
  assign n32555 = n123 & n30470;
  assign n32556 = n128 & n26328;
  assign n32557 = n53444 & n26334;
  assign n32558 = n127 & n26331;
  assign n32559 = ~n32557 & ~n32558;
  assign n32560 = ~n32556 & ~n32558;
  assign n32561 = ~n32557 & n32560;
  assign n32562 = ~n32556 & n32559;
  assign n32563 = ~n123 & n57322;
  assign n32564 = ~n30470 & n57322;
  assign n32565 = ~n32563 & ~n32564;
  assign n32566 = ~n32555 & n57322;
  assign n32567 = pi26  & ~n57323;
  assign n32568 = ~pi26  & n57323;
  assign n32569 = ~n32567 & ~n32568;
  assign n32570 = n32152 & n57267;
  assign n32571 = ~n57267 & ~n32158;
  assign n32572 = ~n32152 & ~n32158;
  assign n32573 = ~n32571 & ~n32572;
  assign n32574 = ~n32158 & ~n32570;
  assign n32575 = ~n32569 & ~n57324;
  assign n32576 = n123 & ~n57033;
  assign n32577 = n128 & n26331;
  assign n32578 = n127 & n26334;
  assign n32579 = n53444 & n26337;
  assign n32580 = ~n32578 & ~n32579;
  assign n32581 = ~n32577 & ~n32579;
  assign n32582 = ~n32578 & n32581;
  assign n32583 = ~n32577 & n32580;
  assign n32584 = ~n32576 & n57325;
  assign n32585 = pi26  & ~n32584;
  assign n32586 = ~n32584 & ~n32585;
  assign n32587 = ~pi26  & ~n32584;
  assign n32588 = pi26  & ~n32585;
  assign n32589 = pi26  & n32584;
  assign n32590 = ~n57326 & ~n57327;
  assign n32591 = n32145 & n57266;
  assign n32592 = ~n32151 & ~n32591;
  assign n32593 = ~n32590 & n32592;
  assign n32594 = n123 & ~n57042;
  assign n32595 = n128 & n26334;
  assign n32596 = n53444 & n26340;
  assign n32597 = n127 & n26337;
  assign n32598 = ~n32596 & ~n32597;
  assign n32599 = ~n32595 & ~n32597;
  assign n32600 = ~n32596 & n32599;
  assign n32601 = ~n32595 & n32598;
  assign n32602 = ~n32594 & n57328;
  assign n32603 = pi26  & ~n32602;
  assign n32604 = ~n32602 & ~n32603;
  assign n32605 = ~pi26  & ~n32602;
  assign n32606 = pi26  & ~n32603;
  assign n32607 = pi26  & n32602;
  assign n32608 = ~n57329 & ~n57330;
  assign n32609 = pi29  & ~n57261;
  assign n32610 = ~n57262 & ~n32609;
  assign n32611 = n57262 & n32609;
  assign n32612 = ~n57261 & n32129;
  assign n32613 = ~n57263 & ~n32612;
  assign n32614 = ~n32610 & ~n32611;
  assign n32615 = ~n32608 & n57331;
  assign n32616 = n123 & n30866;
  assign n32617 = n128 & n26337;
  assign n32618 = n53444 & n26343;
  assign n32619 = n127 & n26340;
  assign n32620 = ~n32618 & ~n32619;
  assign n32621 = ~n32617 & ~n32619;
  assign n32622 = ~n32618 & n32621;
  assign n32623 = ~n32617 & n32620;
  assign n32624 = ~n123 & n57332;
  assign n32625 = ~n30866 & n57332;
  assign n32626 = ~n32624 & ~n32625;
  assign n32627 = ~n32616 & n57332;
  assign n32628 = pi26  & ~n57333;
  assign n32629 = ~pi26  & n57333;
  assign n32630 = ~n32628 & ~n32629;
  assign n32631 = pi29  & n32109;
  assign n32632 = ~n32108 & n32631;
  assign n32633 = n32108 & ~n32631;
  assign n32634 = ~n32110 & n32114;
  assign n32635 = ~n57261 & ~n32634;
  assign n32636 = ~n32632 & ~n32633;
  assign n32637 = ~n32630 & n57334;
  assign n32638 = n123 & ~n31019;
  assign n32639 = n128 & n26348;
  assign n32640 = n127 & ~n56543;
  assign n32641 = ~n32639 & ~n32640;
  assign n32642 = ~n32638 & n32641;
  assign n32643 = ~n120 & ~n56543;
  assign n32644 = pi26  & ~n32643;
  assign n32645 = pi26  & ~n32642;
  assign n32646 = pi26  & ~n32645;
  assign n32647 = ~n32642 & ~n32645;
  assign n32648 = ~n32646 & ~n32647;
  assign n32649 = n32644 & ~n32648;
  assign n32650 = n32642 & n32644;
  assign n32651 = n123 & ~n31140;
  assign n32652 = n128 & n26343;
  assign n32653 = n53444 & ~n56543;
  assign n32654 = n127 & n26348;
  assign n32655 = ~n32653 & ~n32654;
  assign n32656 = ~n32652 & ~n32654;
  assign n32657 = ~n32653 & n32656;
  assign n32658 = ~n32652 & n32655;
  assign n32659 = ~n123 & n57336;
  assign n32660 = n31140 & n57336;
  assign n32661 = ~n32659 & ~n32660;
  assign n32662 = ~n32651 & n57336;
  assign n32663 = pi26  & ~n57337;
  assign n32664 = ~pi26  & n57337;
  assign n32665 = ~n32663 & ~n32664;
  assign n32666 = n57335 & ~n32665;
  assign n32667 = n57335 & ~n57337;
  assign n32668 = n32109 & n57338;
  assign n32669 = n123 & n30915;
  assign n32670 = n128 & n26340;
  assign n32671 = n53444 & n26348;
  assign n32672 = n127 & n26343;
  assign n32673 = ~n32671 & ~n32672;
  assign n32674 = ~n32670 & ~n32672;
  assign n32675 = ~n32671 & n32674;
  assign n32676 = ~n32670 & n32673;
  assign n32677 = ~n32669 & n57339;
  assign n32678 = pi26  & ~n32677;
  assign n32679 = pi26  & ~n32678;
  assign n32680 = pi26  & n32677;
  assign n32681 = ~n32677 & ~n32678;
  assign n32682 = ~pi26  & ~n32677;
  assign n32683 = ~n57340 & ~n57341;
  assign n32684 = ~n32109 & ~n57338;
  assign n32685 = n57338 & ~n32668;
  assign n32686 = ~n32109 & n57338;
  assign n32687 = n32109 & ~n32668;
  assign n32688 = n32109 & ~n57338;
  assign n32689 = ~n57342 & ~n57343;
  assign n32690 = ~n32668 & ~n32684;
  assign n32691 = ~n32683 & ~n57344;
  assign n32692 = ~n32668 & ~n32691;
  assign n32693 = n32630 & ~n57334;
  assign n32694 = ~n32637 & ~n32693;
  assign n32695 = ~n32692 & n32694;
  assign n32696 = ~n32637 & ~n32695;
  assign n32697 = n32608 & ~n57331;
  assign n32698 = ~n32608 & ~n32615;
  assign n32699 = ~n32608 & ~n57331;
  assign n32700 = n57331 & ~n32615;
  assign n32701 = n32608 & n57331;
  assign n32702 = ~n57345 & ~n57346;
  assign n32703 = ~n32615 & ~n32697;
  assign n32704 = ~n32696 & ~n57347;
  assign n32705 = ~n32615 & ~n32704;
  assign n32706 = n32590 & ~n32592;
  assign n32707 = ~n32590 & ~n32593;
  assign n32708 = ~n32590 & ~n32592;
  assign n32709 = n32592 & ~n32593;
  assign n32710 = n32590 & n32592;
  assign n32711 = ~n57348 & ~n57349;
  assign n32712 = ~n32593 & ~n32706;
  assign n32713 = ~n32705 & ~n57350;
  assign n32714 = ~n32593 & ~n32713;
  assign n32715 = n32569 & n57324;
  assign n32716 = ~n57324 & ~n32575;
  assign n32717 = n32569 & ~n57324;
  assign n32718 = ~n32569 & ~n32575;
  assign n32719 = ~n32569 & n57324;
  assign n32720 = ~n57351 & ~n57352;
  assign n32721 = ~n32575 & ~n32715;
  assign n32722 = ~n32714 & ~n57353;
  assign n32723 = ~n32575 & ~n32722;
  assign n32724 = ~n32538 & n32553;
  assign n32725 = n32538 & ~n32554;
  assign n32726 = n32538 & n32553;
  assign n32727 = ~n32553 & ~n32554;
  assign n32728 = ~n32538 & ~n32553;
  assign n32729 = ~n57354 & ~n57355;
  assign n32730 = ~n32554 & ~n32724;
  assign n32731 = ~n32723 & ~n57356;
  assign n32732 = ~n32554 & ~n32731;
  assign n32733 = ~n32520 & n32535;
  assign n32734 = n32520 & ~n32536;
  assign n32735 = n32520 & n32535;
  assign n32736 = ~n32535 & ~n32536;
  assign n32737 = ~n32520 & ~n32535;
  assign n32738 = ~n57357 & ~n57358;
  assign n32739 = ~n32536 & ~n32733;
  assign n32740 = ~n32732 & ~n57359;
  assign n32741 = ~n32536 & ~n32740;
  assign n32742 = ~n32502 & n32517;
  assign n32743 = n32502 & ~n32518;
  assign n32744 = n32502 & n32517;
  assign n32745 = ~n32517 & ~n32518;
  assign n32746 = ~n32502 & ~n32517;
  assign n32747 = ~n57360 & ~n57361;
  assign n32748 = ~n32518 & ~n32742;
  assign n32749 = ~n32741 & ~n57362;
  assign n32750 = ~n32518 & ~n32749;
  assign n32751 = ~n32486 & n32499;
  assign n32752 = n32486 & ~n32500;
  assign n32753 = n32486 & n32499;
  assign n32754 = ~n32499 & ~n32500;
  assign n32755 = ~n32486 & ~n32499;
  assign n32756 = ~n57363 & ~n57364;
  assign n32757 = ~n32500 & ~n32751;
  assign n32758 = ~n32750 & ~n57365;
  assign n32759 = ~n32500 & ~n32758;
  assign n32760 = ~n32470 & n32483;
  assign n32761 = n32470 & ~n32484;
  assign n32762 = n32470 & n32483;
  assign n32763 = ~n32483 & ~n32484;
  assign n32764 = ~n32470 & ~n32483;
  assign n32765 = ~n57366 & ~n57367;
  assign n32766 = ~n32484 & ~n32760;
  assign n32767 = ~n32759 & ~n57368;
  assign n32768 = ~n32484 & ~n32767;
  assign n32769 = ~n32454 & n32467;
  assign n32770 = n32454 & ~n32468;
  assign n32771 = n32454 & n32467;
  assign n32772 = ~n32467 & ~n32468;
  assign n32773 = ~n32454 & ~n32467;
  assign n32774 = ~n57369 & ~n57370;
  assign n32775 = ~n32468 & ~n32769;
  assign n32776 = ~n32768 & ~n57371;
  assign n32777 = ~n32468 & ~n32776;
  assign n32778 = ~n32438 & n32451;
  assign n32779 = n32438 & ~n32452;
  assign n32780 = n32438 & n32451;
  assign n32781 = ~n32451 & ~n32452;
  assign n32782 = ~n32438 & ~n32451;
  assign n32783 = ~n57372 & ~n57373;
  assign n32784 = ~n32452 & ~n32778;
  assign n32785 = ~n32777 & ~n57374;
  assign n32786 = ~n32452 & ~n32785;
  assign n32787 = ~n32422 & n32435;
  assign n32788 = n32422 & ~n32436;
  assign n32789 = n32422 & n32435;
  assign n32790 = ~n32435 & ~n32436;
  assign n32791 = ~n32422 & ~n32435;
  assign n32792 = ~n57375 & ~n57376;
  assign n32793 = ~n32436 & ~n32787;
  assign n32794 = ~n32786 & ~n57377;
  assign n32795 = ~n32436 & ~n32794;
  assign n32796 = ~n32406 & n32419;
  assign n32797 = ~n32420 & ~n32796;
  assign n32798 = ~n32795 & n32797;
  assign n32799 = ~n32420 & ~n32798;
  assign n32800 = n32230 & ~n32232;
  assign n32801 = n32232 & ~n32233;
  assign n32802 = ~n32230 & ~n32233;
  assign n32803 = ~n32801 & ~n32802;
  assign n32804 = ~n32233 & ~n32800;
  assign n32805 = ~n32799 & ~n57378;
  assign n32806 = n32799 & n57378;
  assign n32807 = n90 & n28107;
  assign n32808 = n14236 & n26289;
  assign n32809 = n54667 & n26295;
  assign n32810 = n14210 & n26292;
  assign n32811 = ~n32809 & ~n32810;
  assign n32812 = ~n32808 & n32811;
  assign n32813 = ~n32807 & n32812;
  assign n32814 = pi23  & ~n32813;
  assign n32815 = pi23  & ~n32814;
  assign n32816 = pi23  & n32813;
  assign n32817 = ~n32813 & ~n32814;
  assign n32818 = ~pi23  & ~n32813;
  assign n32819 = ~n57379 & ~n57380;
  assign n32820 = ~n32806 & ~n32819;
  assign n32821 = ~n32805 & ~n32806;
  assign n32822 = ~n32819 & n32821;
  assign n32823 = ~n32805 & ~n32822;
  assign n32824 = ~n32805 & ~n32820;
  assign n32825 = ~n57309 & ~n57381;
  assign n32826 = n57309 & n57381;
  assign n32827 = n14413 & n27330;
  assign n32828 = n15921 & n26277;
  assign n32829 = n54719 & n26283;
  assign n32830 = n15901 & n26280;
  assign n32831 = ~n32829 & ~n32830;
  assign n32832 = ~n32828 & n32831;
  assign n32833 = ~n32827 & n32832;
  assign n32834 = pi20  & ~n32833;
  assign n32835 = pi20  & ~n32834;
  assign n32836 = pi20  & n32833;
  assign n32837 = ~n32833 & ~n32834;
  assign n32838 = ~pi20  & ~n32833;
  assign n32839 = ~n57382 & ~n57383;
  assign n32840 = ~n32826 & ~n32839;
  assign n32841 = ~n32825 & ~n32826;
  assign n32842 = ~n32839 & n32841;
  assign n32843 = ~n32825 & ~n32842;
  assign n32844 = ~n32825 & ~n32840;
  assign n32845 = ~n57308 & ~n57384;
  assign n32846 = n57308 & n57384;
  assign n32847 = n16079 & n27042;
  assign n32848 = n16696 & n26265;
  assign n32849 = n54886 & n26271;
  assign n32850 = n16676 & n26268;
  assign n32851 = ~n32849 & ~n32850;
  assign n32852 = ~n32848 & n32851;
  assign n32853 = ~n32847 & n32852;
  assign n32854 = pi17  & ~n32853;
  assign n32855 = pi17  & ~n32854;
  assign n32856 = pi17  & n32853;
  assign n32857 = ~n32853 & ~n32854;
  assign n32858 = ~pi17  & ~n32853;
  assign n32859 = ~n57385 & ~n57386;
  assign n32860 = ~n32846 & ~n32859;
  assign n32861 = ~n32845 & ~n32846;
  assign n32862 = ~n32859 & n32861;
  assign n32863 = ~n32845 & ~n32862;
  assign n32864 = ~n32845 & ~n32860;
  assign n32865 = ~n57307 & ~n57387;
  assign n32866 = ~n32387 & ~n32865;
  assign n32867 = n32299 & ~n32300;
  assign n32868 = n32297 & n32299;
  assign n32869 = ~n32297 & ~n32300;
  assign n32870 = ~n32297 & ~n32299;
  assign n32871 = n32297 & ~n32299;
  assign n32872 = ~n32300 & ~n32871;
  assign n32873 = ~n57388 & ~n57389;
  assign n32874 = ~n32866 & n57390;
  assign n32875 = n32866 & ~n57390;
  assign n32876 = n17265 & n27491;
  assign n32877 = n18588 & n26250;
  assign n32878 = n55041 & n26256;
  assign n32879 = n18556 & n26253;
  assign n32880 = ~n32878 & ~n32879;
  assign n32881 = ~n32877 & n32880;
  assign n32882 = ~n32876 & n32881;
  assign n32883 = pi14  & ~n32882;
  assign n32884 = pi14  & ~n32883;
  assign n32885 = pi14  & n32882;
  assign n32886 = ~n32882 & ~n32883;
  assign n32887 = ~pi14  & ~n32882;
  assign n32888 = ~n57391 & ~n57392;
  assign n32889 = ~n32875 & ~n32888;
  assign n32890 = ~n32874 & ~n32875;
  assign n32891 = ~n32888 & n32890;
  assign n32892 = ~n32874 & ~n32891;
  assign n32893 = ~n32874 & ~n32889;
  assign n32894 = ~n57302 & ~n57393;
  assign n32895 = n57302 & n57393;
  assign n32896 = n18846 & ~n56564;
  assign n32897 = n19541 & ~n26537;
  assign n32898 = n55247 & n26244;
  assign n32899 = n19509 & n26242;
  assign n32900 = ~n32898 & ~n32899;
  assign n32901 = ~n32897 & n32900;
  assign n32902 = ~n32896 & n32901;
  assign n32903 = pi11  & ~n32902;
  assign n32904 = pi11  & ~n32903;
  assign n32905 = pi11  & n32902;
  assign n32906 = ~n32902 & ~n32903;
  assign n32907 = ~pi11  & ~n32902;
  assign n32908 = ~n57394 & ~n57395;
  assign n32909 = ~n32895 & ~n32908;
  assign n32910 = ~n32894 & ~n32895;
  assign n32911 = ~n32908 & n32910;
  assign n32912 = ~n32894 & ~n32911;
  assign n32913 = ~n32894 & ~n32909;
  assign n32914 = ~n32366 & ~n57396;
  assign n32915 = n57223 & n57293;
  assign n32916 = ~n32323 & ~n32915;
  assign n32917 = n32366 & n57396;
  assign n32918 = ~n57396 & ~n32914;
  assign n32919 = n32366 & ~n57396;
  assign n32920 = ~n32366 & ~n32914;
  assign n32921 = ~n32366 & n57396;
  assign n32922 = ~n57397 & ~n57398;
  assign n32923 = ~n32914 & ~n32917;
  assign n32924 = n32916 & ~n57399;
  assign n32925 = ~n32914 & ~n32924;
  assign n32926 = n32346 & ~n32347;
  assign n32927 = n32344 & n32346;
  assign n32928 = ~n32344 & ~n32347;
  assign n32929 = ~n32344 & ~n32346;
  assign n32930 = n32344 & ~n32346;
  assign n32931 = ~n32347 & ~n32930;
  assign n32932 = ~n57400 & ~n57401;
  assign n32933 = ~n32925 & n57402;
  assign n32934 = ~n32916 & n57399;
  assign n32935 = ~n32924 & ~n32934;
  assign n32936 = n57307 & n57387;
  assign n32937 = ~n32865 & ~n32936;
  assign n32938 = n17265 & ~n56668;
  assign n32939 = n18588 & n26253;
  assign n32940 = n55041 & n26259;
  assign n32941 = n18556 & n26256;
  assign n32942 = ~n32940 & ~n32941;
  assign n32943 = ~n32939 & n32942;
  assign n32944 = ~n32938 & n32943;
  assign n32945 = pi14  & ~n32944;
  assign n32946 = pi14  & ~n32945;
  assign n32947 = pi14  & n32944;
  assign n32948 = ~n32944 & ~n32945;
  assign n32949 = ~pi14  & ~n32944;
  assign n32950 = ~n57403 & ~n57404;
  assign n32951 = n32937 & ~n32950;
  assign n32952 = ~n32937 & n32950;
  assign n32953 = n32937 & ~n32951;
  assign n32954 = n32937 & n32950;
  assign n32955 = ~n32950 & ~n32951;
  assign n32956 = ~n32937 & ~n32950;
  assign n32957 = ~n57405 & ~n57406;
  assign n32958 = ~n32951 & ~n32952;
  assign n32959 = n32859 & ~n32861;
  assign n32960 = n32861 & ~n32862;
  assign n32961 = ~n32859 & ~n32862;
  assign n32962 = ~n32960 & ~n32961;
  assign n32963 = ~n32862 & ~n32959;
  assign n32964 = n32839 & ~n32841;
  assign n32965 = n32841 & ~n32842;
  assign n32966 = ~n32839 & ~n32842;
  assign n32967 = ~n32965 & ~n32966;
  assign n32968 = ~n32842 & ~n32964;
  assign n32969 = n90 & n28808;
  assign n32970 = n14236 & n26292;
  assign n32971 = n54667 & n26298;
  assign n32972 = n14210 & n26295;
  assign n32973 = ~n32971 & ~n32972;
  assign n32974 = ~n32970 & n32973;
  assign n32975 = ~n32969 & n32974;
  assign n32976 = pi23  & ~n32975;
  assign n32977 = ~n32975 & ~n32976;
  assign n32978 = ~pi23  & ~n32975;
  assign n32979 = pi23  & ~n32976;
  assign n32980 = pi23  & n32975;
  assign n32981 = ~n57410 & ~n57411;
  assign n32982 = n32795 & ~n32797;
  assign n32983 = ~n32798 & ~n32982;
  assign n32984 = ~n32981 & n32983;
  assign n32985 = n90 & n28493;
  assign n32986 = n14236 & n26295;
  assign n32987 = n54667 & n26301;
  assign n32988 = n14210 & n26298;
  assign n32989 = ~n32987 & ~n32988;
  assign n32990 = ~n32986 & n32989;
  assign n32991 = ~n32985 & n32990;
  assign n32992 = pi23  & ~n32991;
  assign n32993 = ~n32991 & ~n32992;
  assign n32994 = ~pi23  & ~n32991;
  assign n32995 = pi23  & ~n32992;
  assign n32996 = pi23  & n32991;
  assign n32997 = ~n57412 & ~n57413;
  assign n32998 = n32786 & n57377;
  assign n32999 = ~n32786 & ~n32794;
  assign n33000 = ~n57377 & ~n32794;
  assign n33001 = ~n32999 & ~n33000;
  assign n33002 = ~n32794 & ~n32998;
  assign n33003 = ~n32997 & ~n57414;
  assign n33004 = n90 & ~n56870;
  assign n33005 = n14236 & n26298;
  assign n33006 = n54667 & n26304;
  assign n33007 = n14210 & n26301;
  assign n33008 = ~n33006 & ~n33007;
  assign n33009 = ~n33005 & n33008;
  assign n33010 = ~n33004 & n33009;
  assign n33011 = pi23  & ~n33010;
  assign n33012 = ~n33010 & ~n33011;
  assign n33013 = ~pi23  & ~n33010;
  assign n33014 = pi23  & ~n33011;
  assign n33015 = pi23  & n33010;
  assign n33016 = ~n57415 & ~n57416;
  assign n33017 = n32777 & n57374;
  assign n33018 = ~n32777 & ~n32785;
  assign n33019 = ~n57374 & ~n32785;
  assign n33020 = ~n33018 & ~n33019;
  assign n33021 = ~n32785 & ~n33017;
  assign n33022 = ~n33016 & ~n57417;
  assign n33023 = n90 & n29446;
  assign n33024 = n14236 & n26301;
  assign n33025 = n54667 & n26307;
  assign n33026 = n14210 & n26304;
  assign n33027 = ~n33025 & ~n33026;
  assign n33028 = ~n33024 & n33027;
  assign n33029 = ~n33023 & n33028;
  assign n33030 = pi23  & ~n33029;
  assign n33031 = ~n33029 & ~n33030;
  assign n33032 = ~pi23  & ~n33029;
  assign n33033 = pi23  & ~n33030;
  assign n33034 = pi23  & n33029;
  assign n33035 = ~n57418 & ~n57419;
  assign n33036 = n32768 & n57371;
  assign n33037 = ~n32768 & ~n32776;
  assign n33038 = ~n57371 & ~n32776;
  assign n33039 = ~n33037 & ~n33038;
  assign n33040 = ~n32776 & ~n33036;
  assign n33041 = ~n33035 & ~n57420;
  assign n33042 = n90 & ~n56867;
  assign n33043 = n14236 & n26304;
  assign n33044 = n54667 & n26310;
  assign n33045 = n14210 & n26307;
  assign n33046 = ~n33044 & ~n33045;
  assign n33047 = ~n33043 & n33046;
  assign n33048 = ~n33042 & n33047;
  assign n33049 = pi23  & ~n33048;
  assign n33050 = ~n33048 & ~n33049;
  assign n33051 = ~pi23  & ~n33048;
  assign n33052 = pi23  & ~n33049;
  assign n33053 = pi23  & n33048;
  assign n33054 = ~n57421 & ~n57422;
  assign n33055 = n32759 & n57368;
  assign n33056 = ~n32759 & ~n32767;
  assign n33057 = ~n57368 & ~n32767;
  assign n33058 = ~n33056 & ~n33057;
  assign n33059 = ~n32767 & ~n33055;
  assign n33060 = ~n33054 & ~n57423;
  assign n33061 = n90 & ~n56928;
  assign n33062 = n14236 & n26307;
  assign n33063 = n54667 & n26313;
  assign n33064 = n14210 & n26310;
  assign n33065 = ~n33063 & ~n33064;
  assign n33066 = ~n33062 & n33065;
  assign n33067 = ~n33061 & n33066;
  assign n33068 = pi23  & ~n33067;
  assign n33069 = ~n33067 & ~n33068;
  assign n33070 = ~pi23  & ~n33067;
  assign n33071 = pi23  & ~n33068;
  assign n33072 = pi23  & n33067;
  assign n33073 = ~n57424 & ~n57425;
  assign n33074 = n32750 & n57365;
  assign n33075 = ~n32750 & ~n32758;
  assign n33076 = ~n32750 & n57365;
  assign n33077 = ~n57365 & ~n32758;
  assign n33078 = n32750 & ~n57365;
  assign n33079 = ~n57426 & ~n57427;
  assign n33080 = ~n32758 & ~n33074;
  assign n33081 = ~n33073 & ~n57428;
  assign n33082 = n90 & ~n57002;
  assign n33083 = n14236 & n26310;
  assign n33084 = n54667 & n26316;
  assign n33085 = n14210 & n26313;
  assign n33086 = ~n33084 & ~n33085;
  assign n33087 = ~n33083 & n33086;
  assign n33088 = ~n33082 & n33087;
  assign n33089 = pi23  & ~n33088;
  assign n33090 = ~n33088 & ~n33089;
  assign n33091 = ~pi23  & ~n33088;
  assign n33092 = pi23  & ~n33089;
  assign n33093 = pi23  & n33088;
  assign n33094 = ~n57429 & ~n57430;
  assign n33095 = n32741 & n57362;
  assign n33096 = ~n32741 & ~n32749;
  assign n33097 = ~n32741 & n57362;
  assign n33098 = ~n57362 & ~n32749;
  assign n33099 = n32741 & ~n57362;
  assign n33100 = ~n57431 & ~n57432;
  assign n33101 = ~n32749 & ~n33095;
  assign n33102 = ~n33094 & ~n57433;
  assign n33103 = n90 & n30192;
  assign n33104 = n14236 & n26313;
  assign n33105 = n54667 & n26319;
  assign n33106 = n14210 & n26316;
  assign n33107 = ~n33105 & ~n33106;
  assign n33108 = ~n33104 & n33107;
  assign n33109 = ~n33103 & n33108;
  assign n33110 = pi23  & ~n33109;
  assign n33111 = ~n33109 & ~n33110;
  assign n33112 = ~pi23  & ~n33109;
  assign n33113 = pi23  & ~n33110;
  assign n33114 = pi23  & n33109;
  assign n33115 = ~n57434 & ~n57435;
  assign n33116 = n32732 & n57359;
  assign n33117 = ~n32732 & ~n32740;
  assign n33118 = ~n32732 & n57359;
  assign n33119 = ~n57359 & ~n32740;
  assign n33120 = n32732 & ~n57359;
  assign n33121 = ~n57436 & ~n57437;
  assign n33122 = ~n32740 & ~n33116;
  assign n33123 = ~n33115 & ~n57438;
  assign n33124 = n90 & ~n56920;
  assign n33125 = n14236 & n26316;
  assign n33126 = n54667 & n26322;
  assign n33127 = n14210 & n26319;
  assign n33128 = ~n33126 & ~n33127;
  assign n33129 = ~n33125 & n33128;
  assign n33130 = ~n33124 & n33129;
  assign n33131 = pi23  & ~n33130;
  assign n33132 = ~n33130 & ~n33131;
  assign n33133 = ~pi23  & ~n33130;
  assign n33134 = pi23  & ~n33131;
  assign n33135 = pi23  & n33130;
  assign n33136 = ~n57439 & ~n57440;
  assign n33137 = n32723 & n57356;
  assign n33138 = ~n32723 & ~n32731;
  assign n33139 = ~n57356 & ~n32731;
  assign n33140 = ~n33138 & ~n33139;
  assign n33141 = ~n32731 & ~n33137;
  assign n33142 = ~n33136 & ~n57441;
  assign n33143 = n90 & n30264;
  assign n33144 = n14236 & n26319;
  assign n33145 = n54667 & n26325;
  assign n33146 = n14210 & n26322;
  assign n33147 = ~n33145 & ~n33146;
  assign n33148 = ~n33144 & n33147;
  assign n33149 = ~n33143 & n33148;
  assign n33150 = pi23  & ~n33149;
  assign n33151 = ~n33149 & ~n33150;
  assign n33152 = ~pi23  & ~n33149;
  assign n33153 = pi23  & ~n33150;
  assign n33154 = pi23  & n33149;
  assign n33155 = ~n57442 & ~n57443;
  assign n33156 = n32714 & n57353;
  assign n33157 = ~n32714 & ~n32722;
  assign n33158 = ~n57353 & ~n32722;
  assign n33159 = ~n33157 & ~n33158;
  assign n33160 = ~n32722 & ~n33156;
  assign n33161 = ~n33155 & ~n57444;
  assign n33162 = n32705 & n57350;
  assign n33163 = ~n32713 & ~n33162;
  assign n33164 = n90 & ~n57012;
  assign n33165 = n14236 & n26322;
  assign n33166 = n54667 & n26328;
  assign n33167 = n14210 & n26325;
  assign n33168 = ~n33166 & ~n33167;
  assign n33169 = ~n33165 & n33168;
  assign n33170 = ~n90 & n33169;
  assign n33171 = n57012 & n33169;
  assign n33172 = ~n33170 & ~n33171;
  assign n33173 = ~n33164 & n33169;
  assign n33174 = pi23  & ~n57445;
  assign n33175 = ~pi23  & n57445;
  assign n33176 = ~n33174 & ~n33175;
  assign n33177 = n33163 & ~n33176;
  assign n33178 = n32696 & n57347;
  assign n33179 = ~n32704 & ~n33178;
  assign n33180 = n90 & ~n57017;
  assign n33181 = n14236 & n26325;
  assign n33182 = n54667 & n26331;
  assign n33183 = n14210 & n26328;
  assign n33184 = ~n33182 & ~n33183;
  assign n33185 = ~n33181 & n33184;
  assign n33186 = ~n90 & n33185;
  assign n33187 = n57017 & n33185;
  assign n33188 = ~n33186 & ~n33187;
  assign n33189 = ~n33180 & n33185;
  assign n33190 = pi23  & ~n57446;
  assign n33191 = ~pi23  & n57446;
  assign n33192 = ~n33190 & ~n33191;
  assign n33193 = n33179 & ~n33192;
  assign n33194 = n90 & n30470;
  assign n33195 = n14236 & n26328;
  assign n33196 = n54667 & n26334;
  assign n33197 = n14210 & n26331;
  assign n33198 = ~n33196 & ~n33197;
  assign n33199 = ~n33195 & n33198;
  assign n33200 = ~n33194 & n33199;
  assign n33201 = pi23  & ~n33200;
  assign n33202 = ~n33200 & ~n33201;
  assign n33203 = ~pi23  & ~n33200;
  assign n33204 = pi23  & ~n33201;
  assign n33205 = pi23  & n33200;
  assign n33206 = ~n57447 & ~n57448;
  assign n33207 = n32692 & ~n32694;
  assign n33208 = ~n32695 & ~n33207;
  assign n33209 = ~n33206 & n33208;
  assign n33210 = n90 & ~n57033;
  assign n33211 = n14236 & n26331;
  assign n33212 = n54667 & n26337;
  assign n33213 = n14210 & n26334;
  assign n33214 = ~n33212 & ~n33213;
  assign n33215 = ~n33211 & n33214;
  assign n33216 = ~n90 & n33215;
  assign n33217 = n57033 & n33215;
  assign n33218 = ~n33216 & ~n33217;
  assign n33219 = ~n33210 & n33215;
  assign n33220 = pi23  & ~n57449;
  assign n33221 = ~pi23  & n57449;
  assign n33222 = ~n33220 & ~n33221;
  assign n33223 = n32683 & n57344;
  assign n33224 = ~n57344 & ~n32691;
  assign n33225 = ~n32683 & ~n32691;
  assign n33226 = ~n33224 & ~n33225;
  assign n33227 = ~n32691 & ~n33223;
  assign n33228 = ~n33222 & ~n57450;
  assign n33229 = n90 & ~n57042;
  assign n33230 = n14236 & n26334;
  assign n33231 = n54667 & n26340;
  assign n33232 = n14210 & n26337;
  assign n33233 = ~n33231 & ~n33232;
  assign n33234 = ~n33230 & n33233;
  assign n33235 = ~n33229 & n33234;
  assign n33236 = pi23  & ~n33235;
  assign n33237 = ~n33235 & ~n33236;
  assign n33238 = ~pi23  & ~n33235;
  assign n33239 = pi23  & ~n33236;
  assign n33240 = pi23  & n33235;
  assign n33241 = ~n57451 & ~n57452;
  assign n33242 = pi26  & ~n57335;
  assign n33243 = ~n57337 & ~n33242;
  assign n33244 = n57337 & n33242;
  assign n33245 = ~n57335 & n32665;
  assign n33246 = ~n57338 & ~n33245;
  assign n33247 = ~n33243 & ~n33244;
  assign n33248 = ~n33241 & n57453;
  assign n33249 = n90 & n30866;
  assign n33250 = n14236 & n26337;
  assign n33251 = n54667 & n26343;
  assign n33252 = n14210 & n26340;
  assign n33253 = ~n33251 & ~n33252;
  assign n33254 = ~n33250 & n33253;
  assign n33255 = ~n90 & n33254;
  assign n33256 = ~n30866 & n33254;
  assign n33257 = ~n33255 & ~n33256;
  assign n33258 = ~n33249 & n33254;
  assign n33259 = pi23  & ~n57454;
  assign n33260 = ~pi23  & n57454;
  assign n33261 = ~n33259 & ~n33260;
  assign n33262 = pi26  & n32643;
  assign n33263 = ~n32642 & n33262;
  assign n33264 = n32642 & ~n33262;
  assign n33265 = ~n32644 & n32648;
  assign n33266 = ~n57335 & ~n33265;
  assign n33267 = ~n33263 & ~n33264;
  assign n33268 = ~n33261 & n57455;
  assign n33269 = n90 & ~n31019;
  assign n33270 = n14210 & ~n56543;
  assign n33271 = n14236 & n26348;
  assign n33272 = ~n33270 & ~n33271;
  assign n33273 = ~n33269 & n33272;
  assign n33274 = n53441 & ~n56543;
  assign n33275 = pi23  & ~n33274;
  assign n33276 = pi23  & ~n33273;
  assign n33277 = pi23  & ~n33276;
  assign n33278 = ~n33273 & ~n33276;
  assign n33279 = ~n33277 & ~n33278;
  assign n33280 = n33275 & ~n33279;
  assign n33281 = n33273 & n33275;
  assign n33282 = n90 & ~n31140;
  assign n33283 = n14236 & n26343;
  assign n33284 = n54667 & ~n56543;
  assign n33285 = n14210 & n26348;
  assign n33286 = ~n33284 & ~n33285;
  assign n33287 = ~n33283 & n33286;
  assign n33288 = ~n90 & n33287;
  assign n33289 = n31140 & n33287;
  assign n33290 = ~n33288 & ~n33289;
  assign n33291 = ~n33282 & n33287;
  assign n33292 = pi23  & ~n57457;
  assign n33293 = ~pi23  & n57457;
  assign n33294 = ~n33292 & ~n33293;
  assign n33295 = n57456 & ~n33294;
  assign n33296 = n57456 & ~n57457;
  assign n33297 = n32643 & n57458;
  assign n33298 = n90 & n30915;
  assign n33299 = n14236 & n26340;
  assign n33300 = n54667 & n26348;
  assign n33301 = n14210 & n26343;
  assign n33302 = ~n33300 & ~n33301;
  assign n33303 = ~n33299 & n33302;
  assign n33304 = ~n33298 & n33303;
  assign n33305 = pi23  & ~n33304;
  assign n33306 = pi23  & ~n33305;
  assign n33307 = pi23  & n33304;
  assign n33308 = ~n33304 & ~n33305;
  assign n33309 = ~pi23  & ~n33304;
  assign n33310 = ~n57459 & ~n57460;
  assign n33311 = ~n32643 & ~n57458;
  assign n33312 = n57458 & ~n33297;
  assign n33313 = ~n32643 & n57458;
  assign n33314 = n32643 & ~n33297;
  assign n33315 = n32643 & ~n57458;
  assign n33316 = ~n57461 & ~n57462;
  assign n33317 = ~n33297 & ~n33311;
  assign n33318 = ~n33310 & ~n57463;
  assign n33319 = ~n33297 & ~n33318;
  assign n33320 = n33261 & ~n57455;
  assign n33321 = ~n33268 & ~n33320;
  assign n33322 = ~n33319 & n33321;
  assign n33323 = ~n33268 & ~n33322;
  assign n33324 = n33241 & ~n57453;
  assign n33325 = ~n33241 & ~n33248;
  assign n33326 = ~n33241 & ~n57453;
  assign n33327 = n57453 & ~n33248;
  assign n33328 = n33241 & n57453;
  assign n33329 = ~n57464 & ~n57465;
  assign n33330 = ~n33248 & ~n33324;
  assign n33331 = ~n33323 & ~n57466;
  assign n33332 = ~n33248 & ~n33331;
  assign n33333 = n33222 & n57450;
  assign n33334 = ~n33228 & ~n33333;
  assign n33335 = ~n33332 & n33334;
  assign n33336 = ~n33228 & ~n33335;
  assign n33337 = n33206 & ~n33208;
  assign n33338 = ~n33206 & ~n33209;
  assign n33339 = ~n33206 & ~n33208;
  assign n33340 = n33208 & ~n33209;
  assign n33341 = n33206 & n33208;
  assign n33342 = ~n57467 & ~n57468;
  assign n33343 = ~n33209 & ~n33337;
  assign n33344 = ~n33336 & ~n57469;
  assign n33345 = ~n33209 & ~n33344;
  assign n33346 = ~n33179 & n33192;
  assign n33347 = n33179 & ~n33193;
  assign n33348 = n33179 & n33192;
  assign n33349 = ~n33192 & ~n33193;
  assign n33350 = ~n33179 & ~n33192;
  assign n33351 = ~n57470 & ~n57471;
  assign n33352 = ~n33193 & ~n33346;
  assign n33353 = ~n33345 & ~n57472;
  assign n33354 = ~n33193 & ~n33353;
  assign n33355 = ~n33163 & n33176;
  assign n33356 = ~n33177 & ~n33355;
  assign n33357 = ~n33354 & n33356;
  assign n33358 = ~n33177 & ~n33357;
  assign n33359 = n33155 & n57444;
  assign n33360 = ~n33155 & ~n33161;
  assign n33361 = ~n33155 & n57444;
  assign n33362 = ~n57444 & ~n33161;
  assign n33363 = n33155 & ~n57444;
  assign n33364 = ~n57473 & ~n57474;
  assign n33365 = ~n33161 & ~n33359;
  assign n33366 = ~n33358 & ~n57475;
  assign n33367 = ~n33161 & ~n33366;
  assign n33368 = n33136 & n57441;
  assign n33369 = ~n33136 & ~n33142;
  assign n33370 = ~n33136 & n57441;
  assign n33371 = ~n57441 & ~n33142;
  assign n33372 = n33136 & ~n57441;
  assign n33373 = ~n57476 & ~n57477;
  assign n33374 = ~n33142 & ~n33368;
  assign n33375 = ~n33367 & ~n57478;
  assign n33376 = ~n33142 & ~n33375;
  assign n33377 = n33115 & n57438;
  assign n33378 = ~n33115 & ~n33123;
  assign n33379 = ~n57438 & ~n33123;
  assign n33380 = ~n33378 & ~n33379;
  assign n33381 = ~n33123 & ~n33377;
  assign n33382 = ~n33376 & ~n57479;
  assign n33383 = ~n33123 & ~n33382;
  assign n33384 = n33094 & n57433;
  assign n33385 = ~n33094 & ~n33102;
  assign n33386 = ~n57433 & ~n33102;
  assign n33387 = ~n33385 & ~n33386;
  assign n33388 = ~n33102 & ~n33384;
  assign n33389 = ~n33383 & ~n57480;
  assign n33390 = ~n33102 & ~n33389;
  assign n33391 = n33073 & n57428;
  assign n33392 = ~n33073 & ~n33081;
  assign n33393 = ~n57428 & ~n33081;
  assign n33394 = ~n33392 & ~n33393;
  assign n33395 = ~n33081 & ~n33391;
  assign n33396 = ~n33390 & ~n57481;
  assign n33397 = ~n33081 & ~n33396;
  assign n33398 = n33054 & n57423;
  assign n33399 = ~n33054 & ~n33060;
  assign n33400 = ~n33054 & n57423;
  assign n33401 = ~n57423 & ~n33060;
  assign n33402 = n33054 & ~n57423;
  assign n33403 = ~n57482 & ~n57483;
  assign n33404 = ~n33060 & ~n33398;
  assign n33405 = ~n33397 & ~n57484;
  assign n33406 = ~n33060 & ~n33405;
  assign n33407 = n33035 & n57420;
  assign n33408 = ~n33035 & ~n33041;
  assign n33409 = ~n33035 & n57420;
  assign n33410 = ~n57420 & ~n33041;
  assign n33411 = n33035 & ~n57420;
  assign n33412 = ~n57485 & ~n57486;
  assign n33413 = ~n33041 & ~n33407;
  assign n33414 = ~n33406 & ~n57487;
  assign n33415 = ~n33041 & ~n33414;
  assign n33416 = n33016 & n57417;
  assign n33417 = ~n33016 & ~n33022;
  assign n33418 = ~n33016 & n57417;
  assign n33419 = ~n57417 & ~n33022;
  assign n33420 = n33016 & ~n57417;
  assign n33421 = ~n57488 & ~n57489;
  assign n33422 = ~n33022 & ~n33416;
  assign n33423 = ~n33415 & ~n57490;
  assign n33424 = ~n33022 & ~n33423;
  assign n33425 = n32997 & n57414;
  assign n33426 = ~n32997 & ~n33003;
  assign n33427 = ~n32997 & n57414;
  assign n33428 = ~n57414 & ~n33003;
  assign n33429 = n32997 & ~n57414;
  assign n33430 = ~n57491 & ~n57492;
  assign n33431 = ~n33003 & ~n33425;
  assign n33432 = ~n33424 & ~n57493;
  assign n33433 = ~n33003 & ~n33432;
  assign n33434 = n32981 & ~n32983;
  assign n33435 = ~n32981 & ~n32984;
  assign n33436 = ~n32981 & ~n32983;
  assign n33437 = n32983 & ~n32984;
  assign n33438 = n32981 & n32983;
  assign n33439 = ~n57494 & ~n57495;
  assign n33440 = ~n32984 & ~n33434;
  assign n33441 = ~n33433 & ~n57496;
  assign n33442 = ~n32984 & ~n33441;
  assign n33443 = n32821 & ~n32822;
  assign n33444 = n32819 & n32821;
  assign n33445 = ~n32819 & ~n32822;
  assign n33446 = ~n32819 & ~n32821;
  assign n33447 = n32819 & ~n32821;
  assign n33448 = ~n32822 & ~n33447;
  assign n33449 = ~n57497 & ~n57498;
  assign n33450 = ~n33442 & n57499;
  assign n33451 = n33442 & ~n57499;
  assign n33452 = n14413 & n27743;
  assign n33453 = n15921 & n26280;
  assign n33454 = n54719 & n26286;
  assign n33455 = n15901 & n26283;
  assign n33456 = ~n33454 & ~n33455;
  assign n33457 = ~n33453 & n33456;
  assign n33458 = ~n33452 & n33457;
  assign n33459 = pi20  & ~n33458;
  assign n33460 = pi20  & ~n33459;
  assign n33461 = pi20  & n33458;
  assign n33462 = ~n33458 & ~n33459;
  assign n33463 = ~pi20  & ~n33458;
  assign n33464 = ~n57500 & ~n57501;
  assign n33465 = ~n33451 & ~n33464;
  assign n33466 = ~n33450 & ~n33451;
  assign n33467 = ~n33464 & n33466;
  assign n33468 = ~n33450 & ~n33467;
  assign n33469 = ~n33450 & ~n33465;
  assign n33470 = ~n57409 & ~n57502;
  assign n33471 = n57409 & n57502;
  assign n33472 = n16079 & ~n56601;
  assign n33473 = n16696 & n26268;
  assign n33474 = n54886 & n26274;
  assign n33475 = n16676 & n26271;
  assign n33476 = ~n33474 & ~n33475;
  assign n33477 = ~n33473 & n33476;
  assign n33478 = ~n33472 & n33477;
  assign n33479 = pi17  & ~n33478;
  assign n33480 = pi17  & ~n33479;
  assign n33481 = pi17  & n33478;
  assign n33482 = ~n33478 & ~n33479;
  assign n33483 = ~pi17  & ~n33478;
  assign n33484 = ~n57503 & ~n57504;
  assign n33485 = ~n33471 & ~n33484;
  assign n33486 = ~n33470 & ~n33471;
  assign n33487 = ~n33484 & n33486;
  assign n33488 = ~n33470 & ~n33487;
  assign n33489 = ~n33470 & ~n33485;
  assign n33490 = ~n57408 & ~n57505;
  assign n33491 = n57408 & n57505;
  assign n33492 = n17265 & n27387;
  assign n33493 = n18588 & n26256;
  assign n33494 = n55041 & n26262;
  assign n33495 = n18556 & n26259;
  assign n33496 = ~n33494 & ~n33495;
  assign n33497 = ~n33493 & n33496;
  assign n33498 = ~n33492 & n33497;
  assign n33499 = pi14  & ~n33498;
  assign n33500 = pi14  & ~n33499;
  assign n33501 = pi14  & n33498;
  assign n33502 = ~n33498 & ~n33499;
  assign n33503 = ~pi14  & ~n33498;
  assign n33504 = ~n57506 & ~n57507;
  assign n33505 = ~n33491 & ~n33504;
  assign n33506 = ~n33490 & ~n33491;
  assign n33507 = ~n33504 & n33506;
  assign n33508 = ~n33490 & ~n33507;
  assign n33509 = ~n33490 & ~n33505;
  assign n33510 = ~n57407 & ~n57508;
  assign n33511 = ~n32951 & ~n33510;
  assign n33512 = n32888 & ~n32890;
  assign n33513 = n32890 & ~n32891;
  assign n33514 = ~n32888 & ~n32891;
  assign n33515 = ~n33513 & ~n33514;
  assign n33516 = ~n32891 & ~n33512;
  assign n33517 = ~n33511 & ~n57509;
  assign n33518 = n33511 & n57509;
  assign n33519 = n18846 & n27808;
  assign n33520 = n19541 & n26242;
  assign n33521 = n55247 & n26247;
  assign n33522 = n19509 & n26244;
  assign n33523 = ~n33521 & ~n33522;
  assign n33524 = ~n33520 & n33523;
  assign n33525 = ~n33519 & n33524;
  assign n33526 = pi11  & ~n33525;
  assign n33527 = pi11  & ~n33526;
  assign n33528 = pi11  & n33525;
  assign n33529 = ~n33525 & ~n33526;
  assign n33530 = ~pi11  & ~n33525;
  assign n33531 = ~n57510 & ~n57511;
  assign n33532 = ~n33518 & ~n33531;
  assign n33533 = ~n33517 & ~n33518;
  assign n33534 = ~n33531 & n33533;
  assign n33535 = ~n33517 & ~n33534;
  assign n33536 = ~n33517 & ~n33532;
  assign n33537 = ~n28484 & ~n57512;
  assign n33538 = n28484 & n57512;
  assign n33539 = n32908 & ~n32910;
  assign n33540 = n32910 & ~n32911;
  assign n33541 = ~n32908 & ~n32911;
  assign n33542 = ~n33540 & ~n33541;
  assign n33543 = ~n32911 & ~n33539;
  assign n33544 = ~n33538 & ~n57513;
  assign n33545 = ~n33537 & ~n33538;
  assign n33546 = ~n57513 & n33545;
  assign n33547 = ~n33537 & ~n33546;
  assign n33548 = ~n33537 & ~n33544;
  assign n33549 = n32935 & ~n57514;
  assign n33550 = n57513 & ~n33545;
  assign n33551 = ~n57513 & ~n33546;
  assign n33552 = n33545 & ~n33546;
  assign n33553 = ~n33551 & ~n33552;
  assign n33554 = ~n33546 & ~n33550;
  assign n33555 = n57407 & n57508;
  assign n33556 = ~n33510 & ~n33555;
  assign n33557 = n18846 & n27839;
  assign n33558 = n19541 & n26244;
  assign n33559 = n55247 & n26250;
  assign n33560 = n19509 & n26247;
  assign n33561 = ~n33559 & ~n33560;
  assign n33562 = ~n33558 & n33561;
  assign n33563 = ~n33557 & n33562;
  assign n33564 = pi11  & ~n33563;
  assign n33565 = pi11  & ~n33564;
  assign n33566 = pi11  & n33563;
  assign n33567 = ~n33563 & ~n33564;
  assign n33568 = ~pi11  & ~n33563;
  assign n33569 = ~n57516 & ~n57517;
  assign n33570 = n33556 & ~n33569;
  assign n33571 = ~n33556 & n33569;
  assign n33572 = n33556 & ~n33570;
  assign n33573 = n33556 & n33569;
  assign n33574 = ~n33569 & ~n33570;
  assign n33575 = ~n33556 & ~n33569;
  assign n33576 = ~n57518 & ~n57519;
  assign n33577 = ~n33570 & ~n33571;
  assign n33578 = n33504 & ~n33506;
  assign n33579 = n33506 & ~n33507;
  assign n33580 = ~n33504 & ~n33507;
  assign n33581 = ~n33579 & ~n33580;
  assign n33582 = ~n33507 & ~n33578;
  assign n33583 = n33484 & ~n33486;
  assign n33584 = n33486 & ~n33487;
  assign n33585 = ~n33484 & ~n33487;
  assign n33586 = ~n33584 & ~n33585;
  assign n33587 = ~n33487 & ~n33583;
  assign n33588 = n33433 & n57496;
  assign n33589 = ~n33441 & ~n33588;
  assign n33590 = n14413 & ~n56686;
  assign n33591 = n15921 & n26283;
  assign n33592 = n54719 & n26289;
  assign n33593 = n15901 & n26286;
  assign n33594 = ~n33592 & ~n33593;
  assign n33595 = ~n33591 & n33594;
  assign n33596 = ~n14413 & n33595;
  assign n33597 = n56686 & n33595;
  assign n33598 = ~n33596 & ~n33597;
  assign n33599 = ~n33590 & n33595;
  assign n33600 = pi20  & ~n57523;
  assign n33601 = ~pi20  & n57523;
  assign n33602 = ~n33600 & ~n33601;
  assign n33603 = n33589 & ~n33602;
  assign n33604 = n33424 & n57493;
  assign n33605 = ~n33432 & ~n33604;
  assign n33606 = n14413 & ~n56721;
  assign n33607 = n15921 & n26286;
  assign n33608 = n54719 & n26292;
  assign n33609 = n15901 & n26289;
  assign n33610 = ~n33608 & ~n33609;
  assign n33611 = ~n33607 & n33610;
  assign n33612 = ~n14413 & n33611;
  assign n33613 = n56721 & n33611;
  assign n33614 = ~n33612 & ~n33613;
  assign n33615 = ~n33606 & n33611;
  assign n33616 = pi20  & ~n57524;
  assign n33617 = ~pi20  & n57524;
  assign n33618 = ~n33616 & ~n33617;
  assign n33619 = n33605 & ~n33618;
  assign n33620 = n33415 & n57490;
  assign n33621 = ~n33423 & ~n33620;
  assign n33622 = n14413 & n28107;
  assign n33623 = n15921 & n26289;
  assign n33624 = n54719 & n26295;
  assign n33625 = n15901 & n26292;
  assign n33626 = ~n33624 & ~n33625;
  assign n33627 = ~n33623 & n33626;
  assign n33628 = ~n14413 & n33627;
  assign n33629 = ~n28107 & n33627;
  assign n33630 = ~n33628 & ~n33629;
  assign n33631 = ~n33622 & n33627;
  assign n33632 = pi20  & ~n57525;
  assign n33633 = ~pi20  & n57525;
  assign n33634 = ~n33632 & ~n33633;
  assign n33635 = n33621 & ~n33634;
  assign n33636 = n33406 & n57487;
  assign n33637 = ~n33414 & ~n33636;
  assign n33638 = n14413 & n28808;
  assign n33639 = n15921 & n26292;
  assign n33640 = n54719 & n26298;
  assign n33641 = n15901 & n26295;
  assign n33642 = ~n33640 & ~n33641;
  assign n33643 = ~n33639 & n33642;
  assign n33644 = ~n14413 & n33643;
  assign n33645 = ~n28808 & n33643;
  assign n33646 = ~n33644 & ~n33645;
  assign n33647 = ~n33638 & n33643;
  assign n33648 = pi20  & ~n57526;
  assign n33649 = ~pi20  & n57526;
  assign n33650 = ~n33648 & ~n33649;
  assign n33651 = n33637 & ~n33650;
  assign n33652 = n33397 & n57484;
  assign n33653 = ~n33405 & ~n33652;
  assign n33654 = n14413 & n28493;
  assign n33655 = n15921 & n26295;
  assign n33656 = n54719 & n26301;
  assign n33657 = n15901 & n26298;
  assign n33658 = ~n33656 & ~n33657;
  assign n33659 = ~n33655 & n33658;
  assign n33660 = ~n14413 & n33659;
  assign n33661 = ~n28493 & n33659;
  assign n33662 = ~n33660 & ~n33661;
  assign n33663 = ~n33654 & n33659;
  assign n33664 = pi20  & ~n57527;
  assign n33665 = ~pi20  & n57527;
  assign n33666 = ~n33664 & ~n33665;
  assign n33667 = n33653 & ~n33666;
  assign n33668 = n33390 & n57481;
  assign n33669 = ~n33396 & ~n33668;
  assign n33670 = n14413 & ~n56870;
  assign n33671 = n15921 & n26298;
  assign n33672 = n54719 & n26304;
  assign n33673 = n15901 & n26301;
  assign n33674 = ~n33672 & ~n33673;
  assign n33675 = ~n33671 & n33674;
  assign n33676 = ~n14413 & n33675;
  assign n33677 = n56870 & n33675;
  assign n33678 = ~n33676 & ~n33677;
  assign n33679 = ~n33670 & n33675;
  assign n33680 = pi20  & ~n57528;
  assign n33681 = ~pi20  & n57528;
  assign n33682 = ~n33680 & ~n33681;
  assign n33683 = n33669 & ~n33682;
  assign n33684 = n33383 & n57480;
  assign n33685 = ~n33389 & ~n33684;
  assign n33686 = n14413 & n29446;
  assign n33687 = n15921 & n26301;
  assign n33688 = n54719 & n26307;
  assign n33689 = n15901 & n26304;
  assign n33690 = ~n33688 & ~n33689;
  assign n33691 = ~n33687 & n33690;
  assign n33692 = ~n14413 & n33691;
  assign n33693 = ~n29446 & n33691;
  assign n33694 = ~n33692 & ~n33693;
  assign n33695 = ~n33686 & n33691;
  assign n33696 = pi20  & ~n57529;
  assign n33697 = ~pi20  & n57529;
  assign n33698 = ~n33696 & ~n33697;
  assign n33699 = n33685 & ~n33698;
  assign n33700 = n33376 & n57479;
  assign n33701 = ~n33382 & ~n33700;
  assign n33702 = n14413 & ~n56867;
  assign n33703 = n15921 & n26304;
  assign n33704 = n54719 & n26310;
  assign n33705 = n15901 & n26307;
  assign n33706 = ~n33704 & ~n33705;
  assign n33707 = ~n33703 & n33706;
  assign n33708 = ~n14413 & n33707;
  assign n33709 = n56867 & n33707;
  assign n33710 = ~n33708 & ~n33709;
  assign n33711 = ~n33702 & n33707;
  assign n33712 = pi20  & ~n57530;
  assign n33713 = ~pi20  & n57530;
  assign n33714 = ~n33712 & ~n33713;
  assign n33715 = n33701 & ~n33714;
  assign n33716 = n33367 & n57478;
  assign n33717 = ~n33375 & ~n33716;
  assign n33718 = n14413 & ~n56928;
  assign n33719 = n15921 & n26307;
  assign n33720 = n54719 & n26313;
  assign n33721 = n15901 & n26310;
  assign n33722 = ~n33720 & ~n33721;
  assign n33723 = ~n33719 & n33722;
  assign n33724 = ~n14413 & n33723;
  assign n33725 = n56928 & n33723;
  assign n33726 = ~n33724 & ~n33725;
  assign n33727 = ~n33718 & n33723;
  assign n33728 = pi20  & ~n57531;
  assign n33729 = ~pi20  & n57531;
  assign n33730 = ~n33728 & ~n33729;
  assign n33731 = n33717 & ~n33730;
  assign n33732 = n33358 & n57475;
  assign n33733 = ~n33366 & ~n33732;
  assign n33734 = n14413 & ~n57002;
  assign n33735 = n15921 & n26310;
  assign n33736 = n54719 & n26316;
  assign n33737 = n15901 & n26313;
  assign n33738 = ~n33736 & ~n33737;
  assign n33739 = ~n33735 & n33738;
  assign n33740 = ~n14413 & n33739;
  assign n33741 = n57002 & n33739;
  assign n33742 = ~n33740 & ~n33741;
  assign n33743 = ~n33734 & n33739;
  assign n33744 = pi20  & ~n57532;
  assign n33745 = ~pi20  & n57532;
  assign n33746 = ~n33744 & ~n33745;
  assign n33747 = n33733 & ~n33746;
  assign n33748 = n14413 & n30192;
  assign n33749 = n15921 & n26313;
  assign n33750 = n54719 & n26319;
  assign n33751 = n15901 & n26316;
  assign n33752 = ~n33750 & ~n33751;
  assign n33753 = ~n33749 & n33752;
  assign n33754 = ~n33748 & n33753;
  assign n33755 = pi20  & ~n33754;
  assign n33756 = ~n33754 & ~n33755;
  assign n33757 = ~pi20  & ~n33754;
  assign n33758 = pi20  & ~n33755;
  assign n33759 = pi20  & n33754;
  assign n33760 = ~n57533 & ~n57534;
  assign n33761 = n33354 & ~n33356;
  assign n33762 = ~n33357 & ~n33761;
  assign n33763 = ~n33760 & n33762;
  assign n33764 = n14413 & ~n56920;
  assign n33765 = n15921 & n26316;
  assign n33766 = n54719 & n26322;
  assign n33767 = n15901 & n26319;
  assign n33768 = ~n33766 & ~n33767;
  assign n33769 = ~n33765 & n33768;
  assign n33770 = ~n33764 & n33769;
  assign n33771 = pi20  & ~n33770;
  assign n33772 = ~n33770 & ~n33771;
  assign n33773 = ~pi20  & ~n33770;
  assign n33774 = pi20  & ~n33771;
  assign n33775 = pi20  & n33770;
  assign n33776 = ~n57535 & ~n57536;
  assign n33777 = n33345 & n57472;
  assign n33778 = ~n33345 & ~n33353;
  assign n33779 = ~n33345 & n57472;
  assign n33780 = ~n57472 & ~n33353;
  assign n33781 = n33345 & ~n57472;
  assign n33782 = ~n57537 & ~n57538;
  assign n33783 = ~n33353 & ~n33777;
  assign n33784 = ~n33776 & ~n57539;
  assign n33785 = n33336 & n57469;
  assign n33786 = ~n33344 & ~n33785;
  assign n33787 = n14413 & n30264;
  assign n33788 = n15921 & n26319;
  assign n33789 = n54719 & n26325;
  assign n33790 = n15901 & n26322;
  assign n33791 = ~n33789 & ~n33790;
  assign n33792 = ~n33788 & n33791;
  assign n33793 = ~n14413 & n33792;
  assign n33794 = ~n30264 & n33792;
  assign n33795 = ~n33793 & ~n33794;
  assign n33796 = ~n33787 & n33792;
  assign n33797 = pi20  & ~n57540;
  assign n33798 = ~pi20  & n57540;
  assign n33799 = ~n33797 & ~n33798;
  assign n33800 = n33786 & ~n33799;
  assign n33801 = n33332 & ~n33334;
  assign n33802 = ~n33335 & ~n33801;
  assign n33803 = n14413 & ~n57012;
  assign n33804 = n15921 & n26322;
  assign n33805 = n54719 & n26328;
  assign n33806 = n15901 & n26325;
  assign n33807 = ~n33805 & ~n33806;
  assign n33808 = ~n33804 & n33807;
  assign n33809 = ~n14413 & n33808;
  assign n33810 = n57012 & n33808;
  assign n33811 = ~n33809 & ~n33810;
  assign n33812 = ~n33803 & n33808;
  assign n33813 = pi20  & ~n57541;
  assign n33814 = ~pi20  & n57541;
  assign n33815 = ~n33813 & ~n33814;
  assign n33816 = n33802 & ~n33815;
  assign n33817 = n33323 & n57466;
  assign n33818 = ~n33331 & ~n33817;
  assign n33819 = n14413 & ~n57017;
  assign n33820 = n15921 & n26325;
  assign n33821 = n54719 & n26331;
  assign n33822 = n15901 & n26328;
  assign n33823 = ~n33821 & ~n33822;
  assign n33824 = ~n33820 & n33823;
  assign n33825 = ~n14413 & n33824;
  assign n33826 = n57017 & n33824;
  assign n33827 = ~n33825 & ~n33826;
  assign n33828 = ~n33819 & n33824;
  assign n33829 = pi20  & ~n57542;
  assign n33830 = ~pi20  & n57542;
  assign n33831 = ~n33829 & ~n33830;
  assign n33832 = n33818 & ~n33831;
  assign n33833 = n14413 & n30470;
  assign n33834 = n15921 & n26328;
  assign n33835 = n54719 & n26334;
  assign n33836 = n15901 & n26331;
  assign n33837 = ~n33835 & ~n33836;
  assign n33838 = ~n33834 & n33837;
  assign n33839 = ~n33833 & n33838;
  assign n33840 = pi20  & ~n33839;
  assign n33841 = ~n33839 & ~n33840;
  assign n33842 = ~pi20  & ~n33839;
  assign n33843 = pi20  & ~n33840;
  assign n33844 = pi20  & n33839;
  assign n33845 = ~n57543 & ~n57544;
  assign n33846 = n33319 & ~n33321;
  assign n33847 = ~n33322 & ~n33846;
  assign n33848 = ~n33845 & n33847;
  assign n33849 = n14413 & ~n57033;
  assign n33850 = n15921 & n26331;
  assign n33851 = n54719 & n26337;
  assign n33852 = n15901 & n26334;
  assign n33853 = ~n33851 & ~n33852;
  assign n33854 = ~n33850 & n33853;
  assign n33855 = ~n14413 & n33854;
  assign n33856 = n57033 & n33854;
  assign n33857 = ~n33855 & ~n33856;
  assign n33858 = ~n33849 & n33854;
  assign n33859 = pi20  & ~n57545;
  assign n33860 = ~pi20  & n57545;
  assign n33861 = ~n33859 & ~n33860;
  assign n33862 = n33310 & n57463;
  assign n33863 = ~n57463 & ~n33318;
  assign n33864 = ~n33310 & ~n33318;
  assign n33865 = ~n33863 & ~n33864;
  assign n33866 = ~n33318 & ~n33862;
  assign n33867 = ~n33861 & ~n57546;
  assign n33868 = n14413 & ~n57042;
  assign n33869 = n15921 & n26334;
  assign n33870 = n54719 & n26340;
  assign n33871 = n15901 & n26337;
  assign n33872 = ~n33870 & ~n33871;
  assign n33873 = ~n33869 & n33872;
  assign n33874 = ~n33868 & n33873;
  assign n33875 = pi20  & ~n33874;
  assign n33876 = ~n33874 & ~n33875;
  assign n33877 = ~pi20  & ~n33874;
  assign n33878 = pi20  & ~n33875;
  assign n33879 = pi20  & n33874;
  assign n33880 = ~n57547 & ~n57548;
  assign n33881 = pi23  & ~n57456;
  assign n33882 = ~n57457 & ~n33881;
  assign n33883 = n57457 & n33881;
  assign n33884 = ~n57456 & n33294;
  assign n33885 = ~n57458 & ~n33884;
  assign n33886 = ~n33882 & ~n33883;
  assign n33887 = ~n33880 & n57549;
  assign n33888 = n14413 & n30866;
  assign n33889 = n15921 & n26337;
  assign n33890 = n54719 & n26343;
  assign n33891 = n15901 & n26340;
  assign n33892 = ~n33890 & ~n33891;
  assign n33893 = ~n33889 & n33892;
  assign n33894 = ~n14413 & n33893;
  assign n33895 = ~n30866 & n33893;
  assign n33896 = ~n33894 & ~n33895;
  assign n33897 = ~n33888 & n33893;
  assign n33898 = pi20  & ~n57550;
  assign n33899 = ~pi20  & n57550;
  assign n33900 = ~n33898 & ~n33899;
  assign n33901 = pi23  & n33274;
  assign n33902 = ~n33273 & n33901;
  assign n33903 = n33273 & ~n33901;
  assign n33904 = ~n33275 & n33279;
  assign n33905 = ~n57456 & ~n33904;
  assign n33906 = ~n33902 & ~n33903;
  assign n33907 = ~n33900 & n57551;
  assign n33908 = n14413 & ~n31019;
  assign n33909 = n15901 & ~n56543;
  assign n33910 = n15921 & n26348;
  assign n33911 = ~n33909 & ~n33910;
  assign n33912 = ~n33908 & n33911;
  assign n33913 = n54717 & ~n56543;
  assign n33914 = pi20  & ~n33913;
  assign n33915 = pi20  & ~n33912;
  assign n33916 = pi20  & ~n33915;
  assign n33917 = ~n33912 & ~n33915;
  assign n33918 = ~n33916 & ~n33917;
  assign n33919 = n33914 & ~n33918;
  assign n33920 = n33912 & n33914;
  assign n33921 = n14413 & ~n31140;
  assign n33922 = n15921 & n26343;
  assign n33923 = n54719 & ~n56543;
  assign n33924 = n15901 & n26348;
  assign n33925 = ~n33923 & ~n33924;
  assign n33926 = ~n33922 & n33925;
  assign n33927 = ~n14413 & n33926;
  assign n33928 = n31140 & n33926;
  assign n33929 = ~n33927 & ~n33928;
  assign n33930 = ~n33921 & n33926;
  assign n33931 = pi20  & ~n57553;
  assign n33932 = ~pi20  & n57553;
  assign n33933 = ~n33931 & ~n33932;
  assign n33934 = n57552 & ~n33933;
  assign n33935 = n57552 & ~n57553;
  assign n33936 = n33274 & n57554;
  assign n33937 = n14413 & n30915;
  assign n33938 = n15921 & n26340;
  assign n33939 = n54719 & n26348;
  assign n33940 = n15901 & n26343;
  assign n33941 = ~n33939 & ~n33940;
  assign n33942 = ~n33938 & n33941;
  assign n33943 = ~n33937 & n33942;
  assign n33944 = pi20  & ~n33943;
  assign n33945 = pi20  & ~n33944;
  assign n33946 = pi20  & n33943;
  assign n33947 = ~n33943 & ~n33944;
  assign n33948 = ~pi20  & ~n33943;
  assign n33949 = ~n57555 & ~n57556;
  assign n33950 = ~n33274 & ~n57554;
  assign n33951 = n57554 & ~n33936;
  assign n33952 = ~n33274 & n57554;
  assign n33953 = n33274 & ~n33936;
  assign n33954 = n33274 & ~n57554;
  assign n33955 = ~n57557 & ~n57558;
  assign n33956 = ~n33936 & ~n33950;
  assign n33957 = ~n33949 & ~n57559;
  assign n33958 = ~n33936 & ~n33957;
  assign n33959 = n33900 & ~n57551;
  assign n33960 = ~n33907 & ~n33959;
  assign n33961 = ~n33958 & n33960;
  assign n33962 = ~n33907 & ~n33961;
  assign n33963 = n33880 & ~n57549;
  assign n33964 = ~n33880 & ~n33887;
  assign n33965 = ~n33880 & ~n57549;
  assign n33966 = n57549 & ~n33887;
  assign n33967 = n33880 & n57549;
  assign n33968 = ~n57560 & ~n57561;
  assign n33969 = ~n33887 & ~n33963;
  assign n33970 = ~n33962 & ~n57562;
  assign n33971 = ~n33887 & ~n33970;
  assign n33972 = n33861 & n57546;
  assign n33973 = ~n33867 & ~n33972;
  assign n33974 = ~n33971 & n33973;
  assign n33975 = ~n33867 & ~n33974;
  assign n33976 = n33845 & ~n33847;
  assign n33977 = ~n33845 & ~n33848;
  assign n33978 = ~n33845 & ~n33847;
  assign n33979 = n33847 & ~n33848;
  assign n33980 = n33845 & n33847;
  assign n33981 = ~n57563 & ~n57564;
  assign n33982 = ~n33848 & ~n33976;
  assign n33983 = ~n33975 & ~n57565;
  assign n33984 = ~n33848 & ~n33983;
  assign n33985 = ~n33818 & n33831;
  assign n33986 = n33818 & ~n33832;
  assign n33987 = n33818 & n33831;
  assign n33988 = ~n33831 & ~n33832;
  assign n33989 = ~n33818 & ~n33831;
  assign n33990 = ~n57566 & ~n57567;
  assign n33991 = ~n33832 & ~n33985;
  assign n33992 = ~n33984 & ~n57568;
  assign n33993 = ~n33832 & ~n33992;
  assign n33994 = ~n33802 & n33815;
  assign n33995 = n33802 & ~n33816;
  assign n33996 = n33802 & n33815;
  assign n33997 = ~n33815 & ~n33816;
  assign n33998 = ~n33802 & ~n33815;
  assign n33999 = ~n57569 & ~n57570;
  assign n34000 = ~n33816 & ~n33994;
  assign n34001 = ~n33993 & ~n57571;
  assign n34002 = ~n33816 & ~n34001;
  assign n34003 = ~n33786 & n33799;
  assign n34004 = ~n33800 & ~n34003;
  assign n34005 = ~n34002 & n34004;
  assign n34006 = ~n33800 & ~n34005;
  assign n34007 = n33776 & n57539;
  assign n34008 = ~n33776 & ~n33784;
  assign n34009 = ~n57539 & ~n33784;
  assign n34010 = ~n34008 & ~n34009;
  assign n34011 = ~n33784 & ~n34007;
  assign n34012 = ~n34006 & ~n57572;
  assign n34013 = ~n33784 & ~n34012;
  assign n34014 = n33760 & ~n33762;
  assign n34015 = ~n33760 & ~n33763;
  assign n34016 = ~n33760 & ~n33762;
  assign n34017 = n33762 & ~n33763;
  assign n34018 = n33760 & n33762;
  assign n34019 = ~n57573 & ~n57574;
  assign n34020 = ~n33763 & ~n34014;
  assign n34021 = ~n34013 & ~n57575;
  assign n34022 = ~n33763 & ~n34021;
  assign n34023 = ~n33733 & n33746;
  assign n34024 = n33733 & ~n33747;
  assign n34025 = n33733 & n33746;
  assign n34026 = ~n33746 & ~n33747;
  assign n34027 = ~n33733 & ~n33746;
  assign n34028 = ~n57576 & ~n57577;
  assign n34029 = ~n33747 & ~n34023;
  assign n34030 = ~n34022 & ~n57578;
  assign n34031 = ~n33747 & ~n34030;
  assign n34032 = ~n33717 & n33730;
  assign n34033 = n33717 & ~n33731;
  assign n34034 = n33717 & n33730;
  assign n34035 = ~n33730 & ~n33731;
  assign n34036 = ~n33717 & ~n33730;
  assign n34037 = ~n57579 & ~n57580;
  assign n34038 = ~n33731 & ~n34032;
  assign n34039 = ~n34031 & ~n57581;
  assign n34040 = ~n33731 & ~n34039;
  assign n34041 = ~n33701 & n33714;
  assign n34042 = n33701 & ~n33715;
  assign n34043 = n33701 & n33714;
  assign n34044 = ~n33714 & ~n33715;
  assign n34045 = ~n33701 & ~n33714;
  assign n34046 = ~n57582 & ~n57583;
  assign n34047 = ~n33715 & ~n34041;
  assign n34048 = ~n34040 & ~n57584;
  assign n34049 = ~n33715 & ~n34048;
  assign n34050 = ~n33685 & n33698;
  assign n34051 = n33685 & ~n33699;
  assign n34052 = n33685 & n33698;
  assign n34053 = ~n33698 & ~n33699;
  assign n34054 = ~n33685 & ~n33698;
  assign n34055 = ~n57585 & ~n57586;
  assign n34056 = ~n33699 & ~n34050;
  assign n34057 = ~n34049 & ~n57587;
  assign n34058 = ~n33699 & ~n34057;
  assign n34059 = ~n33669 & n33682;
  assign n34060 = n33669 & ~n33683;
  assign n34061 = n33669 & n33682;
  assign n34062 = ~n33682 & ~n33683;
  assign n34063 = ~n33669 & ~n33682;
  assign n34064 = ~n57588 & ~n57589;
  assign n34065 = ~n33683 & ~n34059;
  assign n34066 = ~n34058 & ~n57590;
  assign n34067 = ~n33683 & ~n34066;
  assign n34068 = ~n33653 & n33666;
  assign n34069 = n33653 & ~n33667;
  assign n34070 = n33653 & n33666;
  assign n34071 = ~n33666 & ~n33667;
  assign n34072 = ~n33653 & ~n33666;
  assign n34073 = ~n57591 & ~n57592;
  assign n34074 = ~n33667 & ~n34068;
  assign n34075 = ~n34067 & ~n57593;
  assign n34076 = ~n33667 & ~n34075;
  assign n34077 = ~n33637 & n33650;
  assign n34078 = n33637 & ~n33651;
  assign n34079 = n33637 & n33650;
  assign n34080 = ~n33650 & ~n33651;
  assign n34081 = ~n33637 & ~n33650;
  assign n34082 = ~n57594 & ~n57595;
  assign n34083 = ~n33651 & ~n34077;
  assign n34084 = ~n34076 & ~n57596;
  assign n34085 = ~n33651 & ~n34084;
  assign n34086 = ~n33621 & n33634;
  assign n34087 = n33621 & ~n33635;
  assign n34088 = n33621 & n33634;
  assign n34089 = ~n33634 & ~n33635;
  assign n34090 = ~n33621 & ~n33634;
  assign n34091 = ~n57597 & ~n57598;
  assign n34092 = ~n33635 & ~n34086;
  assign n34093 = ~n34085 & ~n57599;
  assign n34094 = ~n33635 & ~n34093;
  assign n34095 = ~n33605 & n33618;
  assign n34096 = n33605 & ~n33619;
  assign n34097 = n33605 & n33618;
  assign n34098 = ~n33618 & ~n33619;
  assign n34099 = ~n33605 & ~n33618;
  assign n34100 = ~n57600 & ~n57601;
  assign n34101 = ~n33619 & ~n34095;
  assign n34102 = ~n34094 & ~n57602;
  assign n34103 = ~n33619 & ~n34102;
  assign n34104 = ~n33589 & n33602;
  assign n34105 = ~n33603 & ~n34104;
  assign n34106 = ~n34103 & n34105;
  assign n34107 = ~n33603 & ~n34106;
  assign n34108 = n33464 & ~n33466;
  assign n34109 = n33466 & ~n33467;
  assign n34110 = ~n33464 & ~n33467;
  assign n34111 = ~n34109 & ~n34110;
  assign n34112 = ~n33467 & ~n34108;
  assign n34113 = ~n34107 & ~n57603;
  assign n34114 = n34107 & n57603;
  assign n34115 = n16079 & ~n56612;
  assign n34116 = n16696 & n26271;
  assign n34117 = n54886 & n26277;
  assign n34118 = n16676 & n26274;
  assign n34119 = ~n34117 & ~n34118;
  assign n34120 = ~n34116 & n34119;
  assign n34121 = ~n34115 & n34120;
  assign n34122 = pi17  & ~n34121;
  assign n34123 = pi17  & ~n34122;
  assign n34124 = pi17  & n34121;
  assign n34125 = ~n34121 & ~n34122;
  assign n34126 = ~pi17  & ~n34121;
  assign n34127 = ~n57604 & ~n57605;
  assign n34128 = ~n34114 & ~n34127;
  assign n34129 = ~n34113 & ~n34114;
  assign n34130 = ~n34127 & n34129;
  assign n34131 = ~n34113 & ~n34130;
  assign n34132 = ~n34113 & ~n34128;
  assign n34133 = ~n57522 & ~n57606;
  assign n34134 = n57522 & n57606;
  assign n34135 = n17265 & ~n56639;
  assign n34136 = n18588 & n26259;
  assign n34137 = n55041 & n26265;
  assign n34138 = n18556 & n26262;
  assign n34139 = ~n34137 & ~n34138;
  assign n34140 = ~n34136 & n34139;
  assign n34141 = ~n34135 & n34140;
  assign n34142 = pi14  & ~n34141;
  assign n34143 = pi14  & ~n34142;
  assign n34144 = pi14  & n34141;
  assign n34145 = ~n34141 & ~n34142;
  assign n34146 = ~pi14  & ~n34141;
  assign n34147 = ~n57607 & ~n57608;
  assign n34148 = ~n34134 & ~n34147;
  assign n34149 = ~n34133 & ~n34134;
  assign n34150 = ~n34147 & n34149;
  assign n34151 = ~n34133 & ~n34150;
  assign n34152 = ~n34133 & ~n34148;
  assign n34153 = ~n57521 & ~n57609;
  assign n34154 = n57521 & n57609;
  assign n34155 = n18846 & ~n56567;
  assign n34156 = n19541 & n26247;
  assign n34157 = n55247 & n26253;
  assign n34158 = n19509 & n26250;
  assign n34159 = ~n34157 & ~n34158;
  assign n34160 = ~n34156 & n34159;
  assign n34161 = ~n34155 & n34160;
  assign n34162 = pi11  & ~n34161;
  assign n34163 = pi11  & ~n34162;
  assign n34164 = pi11  & n34161;
  assign n34165 = ~n34161 & ~n34162;
  assign n34166 = ~pi11  & ~n34161;
  assign n34167 = ~n57610 & ~n57611;
  assign n34168 = ~n34154 & ~n34167;
  assign n34169 = ~n34153 & ~n34154;
  assign n34170 = ~n34167 & n34169;
  assign n34171 = ~n34153 & ~n34170;
  assign n34172 = ~n34153 & ~n34168;
  assign n34173 = ~n57520 & ~n57612;
  assign n34174 = ~n33570 & ~n34173;
  assign n34175 = n33533 & ~n33534;
  assign n34176 = n33531 & n33533;
  assign n34177 = ~n33531 & ~n33534;
  assign n34178 = ~n33531 & ~n33533;
  assign n34179 = n33531 & ~n33533;
  assign n34180 = ~n33534 & ~n34179;
  assign n34181 = ~n57613 & ~n57614;
  assign n34182 = ~n34174 & n57615;
  assign n34183 = n34174 & ~n57615;
  assign n34184 = n55472 & ~n26537;
  assign n34185 = ~n21237 & ~n34184;
  assign n34186 = ~n21269 & n34185;
  assign n34187 = ~n21269 & ~n34184;
  assign n34188 = ~n21237 & n34187;
  assign n34189 = n56755 & ~n34184;
  assign n34190 = ~n20085 & n57616;
  assign n34191 = pi8  & ~n34190;
  assign n34192 = pi8  & ~n34191;
  assign n34193 = pi8  & n34190;
  assign n34194 = ~n34190 & ~n34191;
  assign n34195 = ~pi8  & ~n34190;
  assign n34196 = ~n57617 & ~n57618;
  assign n34197 = ~n34183 & ~n34196;
  assign n34198 = ~n34182 & ~n34183;
  assign n34199 = ~n34196 & n34198;
  assign n34200 = ~n34182 & ~n34199;
  assign n34201 = ~n34182 & ~n34197;
  assign n34202 = ~n57515 & ~n57619;
  assign n34203 = n57515 & n57619;
  assign n34204 = ~n34202 & ~n34203;
  assign n34205 = n20085 & n28624;
  assign n34206 = n21237 & ~n26537;
  assign n34207 = n55472 & n26242;
  assign n34208 = ~n21269 & ~n34207;
  assign n34209 = ~n34206 & ~n34207;
  assign n34210 = ~n21269 & n34209;
  assign n34211 = ~n34206 & n34208;
  assign n34212 = ~n34205 & n57620;
  assign n34213 = pi8  & ~n34212;
  assign n34214 = pi8  & ~n34213;
  assign n34215 = pi8  & n34212;
  assign n34216 = ~n34212 & ~n34213;
  assign n34217 = ~pi8  & ~n34212;
  assign n34218 = ~n57621 & ~n57622;
  assign n34219 = n34167 & ~n34169;
  assign n34220 = n34169 & ~n34170;
  assign n34221 = ~n34167 & ~n34170;
  assign n34222 = ~n34220 & ~n34221;
  assign n34223 = ~n34170 & ~n34219;
  assign n34224 = n34147 & ~n34149;
  assign n34225 = n34149 & ~n34150;
  assign n34226 = ~n34147 & ~n34150;
  assign n34227 = ~n34225 & ~n34226;
  assign n34228 = ~n34150 & ~n34224;
  assign n34229 = n16079 & ~n56648;
  assign n34230 = n16696 & n26274;
  assign n34231 = n54886 & n26280;
  assign n34232 = n16676 & n26277;
  assign n34233 = ~n34231 & ~n34232;
  assign n34234 = ~n34230 & n34233;
  assign n34235 = ~n34229 & n34234;
  assign n34236 = pi17  & ~n34235;
  assign n34237 = ~n34235 & ~n34236;
  assign n34238 = ~pi17  & ~n34235;
  assign n34239 = pi17  & ~n34236;
  assign n34240 = pi17  & n34235;
  assign n34241 = ~n57625 & ~n57626;
  assign n34242 = n34103 & ~n34105;
  assign n34243 = ~n34106 & ~n34242;
  assign n34244 = ~n34241 & n34243;
  assign n34245 = n16079 & n27330;
  assign n34246 = n16696 & n26277;
  assign n34247 = n54886 & n26283;
  assign n34248 = n16676 & n26280;
  assign n34249 = ~n34247 & ~n34248;
  assign n34250 = ~n34246 & n34249;
  assign n34251 = ~n34245 & n34250;
  assign n34252 = pi17  & ~n34251;
  assign n34253 = ~n34251 & ~n34252;
  assign n34254 = ~pi17  & ~n34251;
  assign n34255 = pi17  & ~n34252;
  assign n34256 = pi17  & n34251;
  assign n34257 = ~n57627 & ~n57628;
  assign n34258 = n34094 & n57602;
  assign n34259 = ~n34094 & ~n34102;
  assign n34260 = ~n34094 & n57602;
  assign n34261 = ~n57602 & ~n34102;
  assign n34262 = n34094 & ~n57602;
  assign n34263 = ~n57629 & ~n57630;
  assign n34264 = ~n34102 & ~n34258;
  assign n34265 = ~n34257 & ~n57631;
  assign n34266 = n16079 & n27743;
  assign n34267 = n16696 & n26280;
  assign n34268 = n54886 & n26286;
  assign n34269 = n16676 & n26283;
  assign n34270 = ~n34268 & ~n34269;
  assign n34271 = ~n34267 & n34270;
  assign n34272 = ~n34266 & n34271;
  assign n34273 = pi17  & ~n34272;
  assign n34274 = ~n34272 & ~n34273;
  assign n34275 = ~pi17  & ~n34272;
  assign n34276 = pi17  & ~n34273;
  assign n34277 = pi17  & n34272;
  assign n34278 = ~n57632 & ~n57633;
  assign n34279 = n34085 & n57599;
  assign n34280 = ~n34085 & ~n34093;
  assign n34281 = ~n34085 & n57599;
  assign n34282 = ~n57599 & ~n34093;
  assign n34283 = n34085 & ~n57599;
  assign n34284 = ~n57634 & ~n57635;
  assign n34285 = ~n34093 & ~n34279;
  assign n34286 = ~n34278 & ~n57636;
  assign n34287 = n16079 & ~n56686;
  assign n34288 = n16696 & n26283;
  assign n34289 = n54886 & n26289;
  assign n34290 = n16676 & n26286;
  assign n34291 = ~n34289 & ~n34290;
  assign n34292 = ~n34288 & n34291;
  assign n34293 = ~n34287 & n34292;
  assign n34294 = pi17  & ~n34293;
  assign n34295 = ~n34293 & ~n34294;
  assign n34296 = ~pi17  & ~n34293;
  assign n34297 = pi17  & ~n34294;
  assign n34298 = pi17  & n34293;
  assign n34299 = ~n57637 & ~n57638;
  assign n34300 = n34076 & n57596;
  assign n34301 = ~n34076 & ~n34084;
  assign n34302 = ~n34076 & n57596;
  assign n34303 = ~n57596 & ~n34084;
  assign n34304 = n34076 & ~n57596;
  assign n34305 = ~n57639 & ~n57640;
  assign n34306 = ~n34084 & ~n34300;
  assign n34307 = ~n34299 & ~n57641;
  assign n34308 = n16079 & ~n56721;
  assign n34309 = n16696 & n26286;
  assign n34310 = n54886 & n26292;
  assign n34311 = n16676 & n26289;
  assign n34312 = ~n34310 & ~n34311;
  assign n34313 = ~n34309 & n34312;
  assign n34314 = ~n34308 & n34313;
  assign n34315 = pi17  & ~n34314;
  assign n34316 = ~n34314 & ~n34315;
  assign n34317 = ~pi17  & ~n34314;
  assign n34318 = pi17  & ~n34315;
  assign n34319 = pi17  & n34314;
  assign n34320 = ~n57642 & ~n57643;
  assign n34321 = n34067 & n57593;
  assign n34322 = ~n34067 & ~n34075;
  assign n34323 = ~n34067 & n57593;
  assign n34324 = ~n57593 & ~n34075;
  assign n34325 = n34067 & ~n57593;
  assign n34326 = ~n57644 & ~n57645;
  assign n34327 = ~n34075 & ~n34321;
  assign n34328 = ~n34320 & ~n57646;
  assign n34329 = n16079 & n28107;
  assign n34330 = n16696 & n26289;
  assign n34331 = n54886 & n26295;
  assign n34332 = n16676 & n26292;
  assign n34333 = ~n34331 & ~n34332;
  assign n34334 = ~n34330 & n34333;
  assign n34335 = ~n34329 & n34334;
  assign n34336 = pi17  & ~n34335;
  assign n34337 = ~n34335 & ~n34336;
  assign n34338 = ~pi17  & ~n34335;
  assign n34339 = pi17  & ~n34336;
  assign n34340 = pi17  & n34335;
  assign n34341 = ~n57647 & ~n57648;
  assign n34342 = n34058 & n57590;
  assign n34343 = ~n34058 & ~n34066;
  assign n34344 = ~n57590 & ~n34066;
  assign n34345 = ~n34343 & ~n34344;
  assign n34346 = ~n34066 & ~n34342;
  assign n34347 = ~n34341 & ~n57649;
  assign n34348 = n16079 & n28808;
  assign n34349 = n16696 & n26292;
  assign n34350 = n54886 & n26298;
  assign n34351 = n16676 & n26295;
  assign n34352 = ~n34350 & ~n34351;
  assign n34353 = ~n34349 & n34352;
  assign n34354 = ~n34348 & n34353;
  assign n34355 = pi17  & ~n34354;
  assign n34356 = ~n34354 & ~n34355;
  assign n34357 = ~pi17  & ~n34354;
  assign n34358 = pi17  & ~n34355;
  assign n34359 = pi17  & n34354;
  assign n34360 = ~n57650 & ~n57651;
  assign n34361 = n34049 & n57587;
  assign n34362 = ~n34049 & ~n34057;
  assign n34363 = ~n57587 & ~n34057;
  assign n34364 = ~n34362 & ~n34363;
  assign n34365 = ~n34057 & ~n34361;
  assign n34366 = ~n34360 & ~n57652;
  assign n34367 = n16079 & n28493;
  assign n34368 = n16696 & n26295;
  assign n34369 = n54886 & n26301;
  assign n34370 = n16676 & n26298;
  assign n34371 = ~n34369 & ~n34370;
  assign n34372 = ~n34368 & n34371;
  assign n34373 = ~n34367 & n34372;
  assign n34374 = pi17  & ~n34373;
  assign n34375 = ~n34373 & ~n34374;
  assign n34376 = ~pi17  & ~n34373;
  assign n34377 = pi17  & ~n34374;
  assign n34378 = pi17  & n34373;
  assign n34379 = ~n57653 & ~n57654;
  assign n34380 = n34040 & n57584;
  assign n34381 = ~n34040 & ~n34048;
  assign n34382 = ~n57584 & ~n34048;
  assign n34383 = ~n34381 & ~n34382;
  assign n34384 = ~n34048 & ~n34380;
  assign n34385 = ~n34379 & ~n57655;
  assign n34386 = n16079 & ~n56870;
  assign n34387 = n16696 & n26298;
  assign n34388 = n54886 & n26304;
  assign n34389 = n16676 & n26301;
  assign n34390 = ~n34388 & ~n34389;
  assign n34391 = ~n34387 & n34390;
  assign n34392 = ~n34386 & n34391;
  assign n34393 = pi17  & ~n34392;
  assign n34394 = ~n34392 & ~n34393;
  assign n34395 = ~pi17  & ~n34392;
  assign n34396 = pi17  & ~n34393;
  assign n34397 = pi17  & n34392;
  assign n34398 = ~n57656 & ~n57657;
  assign n34399 = n34031 & n57581;
  assign n34400 = ~n34031 & ~n34039;
  assign n34401 = ~n34031 & n57581;
  assign n34402 = ~n57581 & ~n34039;
  assign n34403 = n34031 & ~n57581;
  assign n34404 = ~n57658 & ~n57659;
  assign n34405 = ~n34039 & ~n34399;
  assign n34406 = ~n34398 & ~n57660;
  assign n34407 = n16079 & n29446;
  assign n34408 = n16696 & n26301;
  assign n34409 = n54886 & n26307;
  assign n34410 = n16676 & n26304;
  assign n34411 = ~n34409 & ~n34410;
  assign n34412 = ~n34408 & n34411;
  assign n34413 = ~n34407 & n34412;
  assign n34414 = pi17  & ~n34413;
  assign n34415 = ~n34413 & ~n34414;
  assign n34416 = ~pi17  & ~n34413;
  assign n34417 = pi17  & ~n34414;
  assign n34418 = pi17  & n34413;
  assign n34419 = ~n57661 & ~n57662;
  assign n34420 = n34022 & n57578;
  assign n34421 = ~n34022 & ~n34030;
  assign n34422 = ~n34022 & n57578;
  assign n34423 = ~n57578 & ~n34030;
  assign n34424 = n34022 & ~n57578;
  assign n34425 = ~n57663 & ~n57664;
  assign n34426 = ~n34030 & ~n34420;
  assign n34427 = ~n34419 & ~n57665;
  assign n34428 = n34013 & n57575;
  assign n34429 = ~n34021 & ~n34428;
  assign n34430 = n16079 & ~n56867;
  assign n34431 = n16696 & n26304;
  assign n34432 = n54886 & n26310;
  assign n34433 = n16676 & n26307;
  assign n34434 = ~n34432 & ~n34433;
  assign n34435 = ~n34431 & n34434;
  assign n34436 = ~n16079 & n34435;
  assign n34437 = n56867 & n34435;
  assign n34438 = ~n34436 & ~n34437;
  assign n34439 = ~n34430 & n34435;
  assign n34440 = pi17  & ~n57666;
  assign n34441 = ~pi17  & n57666;
  assign n34442 = ~n34440 & ~n34441;
  assign n34443 = n34429 & ~n34442;
  assign n34444 = n34006 & n57572;
  assign n34445 = ~n34012 & ~n34444;
  assign n34446 = n16079 & ~n56928;
  assign n34447 = n16696 & n26307;
  assign n34448 = n54886 & n26313;
  assign n34449 = n16676 & n26310;
  assign n34450 = ~n34448 & ~n34449;
  assign n34451 = ~n34447 & n34450;
  assign n34452 = ~n16079 & n34451;
  assign n34453 = n56928 & n34451;
  assign n34454 = ~n34452 & ~n34453;
  assign n34455 = ~n34446 & n34451;
  assign n34456 = pi17  & ~n57667;
  assign n34457 = ~pi17  & n57667;
  assign n34458 = ~n34456 & ~n34457;
  assign n34459 = n34445 & ~n34458;
  assign n34460 = n16079 & ~n57002;
  assign n34461 = n16696 & n26310;
  assign n34462 = n54886 & n26316;
  assign n34463 = n16676 & n26313;
  assign n34464 = ~n34462 & ~n34463;
  assign n34465 = ~n34461 & n34464;
  assign n34466 = ~n34460 & n34465;
  assign n34467 = pi17  & ~n34466;
  assign n34468 = ~n34466 & ~n34467;
  assign n34469 = ~pi17  & ~n34466;
  assign n34470 = pi17  & ~n34467;
  assign n34471 = pi17  & n34466;
  assign n34472 = ~n57668 & ~n57669;
  assign n34473 = n34002 & ~n34004;
  assign n34474 = ~n34005 & ~n34473;
  assign n34475 = ~n34472 & n34474;
  assign n34476 = n16079 & n30192;
  assign n34477 = n16696 & n26313;
  assign n34478 = n54886 & n26319;
  assign n34479 = n16676 & n26316;
  assign n34480 = ~n34478 & ~n34479;
  assign n34481 = ~n34477 & n34480;
  assign n34482 = ~n34476 & n34481;
  assign n34483 = pi17  & ~n34482;
  assign n34484 = ~n34482 & ~n34483;
  assign n34485 = ~pi17  & ~n34482;
  assign n34486 = pi17  & ~n34483;
  assign n34487 = pi17  & n34482;
  assign n34488 = ~n57670 & ~n57671;
  assign n34489 = n33993 & n57571;
  assign n34490 = ~n33993 & ~n34001;
  assign n34491 = ~n57571 & ~n34001;
  assign n34492 = ~n34490 & ~n34491;
  assign n34493 = ~n34001 & ~n34489;
  assign n34494 = ~n34488 & ~n57672;
  assign n34495 = n16079 & ~n56920;
  assign n34496 = n16696 & n26316;
  assign n34497 = n54886 & n26322;
  assign n34498 = n16676 & n26319;
  assign n34499 = ~n34497 & ~n34498;
  assign n34500 = ~n34496 & n34499;
  assign n34501 = ~n34495 & n34500;
  assign n34502 = pi17  & ~n34501;
  assign n34503 = ~n34501 & ~n34502;
  assign n34504 = ~pi17  & ~n34501;
  assign n34505 = pi17  & ~n34502;
  assign n34506 = pi17  & n34501;
  assign n34507 = ~n57673 & ~n57674;
  assign n34508 = n33984 & n57568;
  assign n34509 = ~n33984 & ~n33992;
  assign n34510 = ~n33984 & n57568;
  assign n34511 = ~n57568 & ~n33992;
  assign n34512 = n33984 & ~n57568;
  assign n34513 = ~n57675 & ~n57676;
  assign n34514 = ~n33992 & ~n34508;
  assign n34515 = ~n34507 & ~n57677;
  assign n34516 = n33975 & n57565;
  assign n34517 = ~n33983 & ~n34516;
  assign n34518 = n16079 & n30264;
  assign n34519 = n16696 & n26319;
  assign n34520 = n54886 & n26325;
  assign n34521 = n16676 & n26322;
  assign n34522 = ~n34520 & ~n34521;
  assign n34523 = ~n34519 & n34522;
  assign n34524 = ~n16079 & n34523;
  assign n34525 = ~n30264 & n34523;
  assign n34526 = ~n34524 & ~n34525;
  assign n34527 = ~n34518 & n34523;
  assign n34528 = pi17  & ~n57678;
  assign n34529 = ~pi17  & n57678;
  assign n34530 = ~n34528 & ~n34529;
  assign n34531 = n34517 & ~n34530;
  assign n34532 = n33971 & ~n33973;
  assign n34533 = ~n33974 & ~n34532;
  assign n34534 = n16079 & ~n57012;
  assign n34535 = n16696 & n26322;
  assign n34536 = n54886 & n26328;
  assign n34537 = n16676 & n26325;
  assign n34538 = ~n34536 & ~n34537;
  assign n34539 = ~n34535 & n34538;
  assign n34540 = ~n16079 & n34539;
  assign n34541 = n57012 & n34539;
  assign n34542 = ~n34540 & ~n34541;
  assign n34543 = ~n34534 & n34539;
  assign n34544 = pi17  & ~n57679;
  assign n34545 = ~pi17  & n57679;
  assign n34546 = ~n34544 & ~n34545;
  assign n34547 = n34533 & ~n34546;
  assign n34548 = n33962 & n57562;
  assign n34549 = ~n33970 & ~n34548;
  assign n34550 = n16079 & ~n57017;
  assign n34551 = n16696 & n26325;
  assign n34552 = n54886 & n26331;
  assign n34553 = n16676 & n26328;
  assign n34554 = ~n34552 & ~n34553;
  assign n34555 = ~n34551 & n34554;
  assign n34556 = ~n16079 & n34555;
  assign n34557 = n57017 & n34555;
  assign n34558 = ~n34556 & ~n34557;
  assign n34559 = ~n34550 & n34555;
  assign n34560 = pi17  & ~n57680;
  assign n34561 = ~pi17  & n57680;
  assign n34562 = ~n34560 & ~n34561;
  assign n34563 = n34549 & ~n34562;
  assign n34564 = n16079 & n30470;
  assign n34565 = n16696 & n26328;
  assign n34566 = n54886 & n26334;
  assign n34567 = n16676 & n26331;
  assign n34568 = ~n34566 & ~n34567;
  assign n34569 = ~n34565 & n34568;
  assign n34570 = ~n34564 & n34569;
  assign n34571 = pi17  & ~n34570;
  assign n34572 = ~n34570 & ~n34571;
  assign n34573 = ~pi17  & ~n34570;
  assign n34574 = pi17  & ~n34571;
  assign n34575 = pi17  & n34570;
  assign n34576 = ~n57681 & ~n57682;
  assign n34577 = n33958 & ~n33960;
  assign n34578 = ~n33961 & ~n34577;
  assign n34579 = ~n34576 & n34578;
  assign n34580 = n16079 & ~n57033;
  assign n34581 = n16696 & n26331;
  assign n34582 = n54886 & n26337;
  assign n34583 = n16676 & n26334;
  assign n34584 = ~n34582 & ~n34583;
  assign n34585 = ~n34581 & n34584;
  assign n34586 = ~n16079 & n34585;
  assign n34587 = n57033 & n34585;
  assign n34588 = ~n34586 & ~n34587;
  assign n34589 = ~n34580 & n34585;
  assign n34590 = pi17  & ~n57683;
  assign n34591 = ~pi17  & n57683;
  assign n34592 = ~n34590 & ~n34591;
  assign n34593 = n33949 & n57559;
  assign n34594 = ~n57559 & ~n33957;
  assign n34595 = ~n33949 & ~n33957;
  assign n34596 = ~n34594 & ~n34595;
  assign n34597 = ~n33957 & ~n34593;
  assign n34598 = ~n34592 & ~n57684;
  assign n34599 = n16079 & ~n57042;
  assign n34600 = n16696 & n26334;
  assign n34601 = n54886 & n26340;
  assign n34602 = n16676 & n26337;
  assign n34603 = ~n34601 & ~n34602;
  assign n34604 = ~n34600 & n34603;
  assign n34605 = ~n34599 & n34604;
  assign n34606 = pi17  & ~n34605;
  assign n34607 = ~n34605 & ~n34606;
  assign n34608 = ~pi17  & ~n34605;
  assign n34609 = pi17  & ~n34606;
  assign n34610 = pi17  & n34605;
  assign n34611 = ~n57685 & ~n57686;
  assign n34612 = pi20  & ~n57552;
  assign n34613 = ~n57553 & ~n34612;
  assign n34614 = n57553 & n34612;
  assign n34615 = ~n57552 & n33933;
  assign n34616 = ~n57554 & ~n34615;
  assign n34617 = ~n34613 & ~n34614;
  assign n34618 = ~n34611 & n57687;
  assign n34619 = n16079 & n30866;
  assign n34620 = n16696 & n26337;
  assign n34621 = n54886 & n26343;
  assign n34622 = n16676 & n26340;
  assign n34623 = ~n34621 & ~n34622;
  assign n34624 = ~n34620 & n34623;
  assign n34625 = ~n16079 & n34624;
  assign n34626 = ~n30866 & n34624;
  assign n34627 = ~n34625 & ~n34626;
  assign n34628 = ~n34619 & n34624;
  assign n34629 = pi17  & ~n57688;
  assign n34630 = ~pi17  & n57688;
  assign n34631 = ~n34629 & ~n34630;
  assign n34632 = pi20  & n33913;
  assign n34633 = ~n33912 & n34632;
  assign n34634 = n33912 & ~n34632;
  assign n34635 = ~n33914 & n33918;
  assign n34636 = ~n57552 & ~n34635;
  assign n34637 = ~n34633 & ~n34634;
  assign n34638 = ~n34631 & n57689;
  assign n34639 = n16079 & ~n31019;
  assign n34640 = n16676 & ~n56543;
  assign n34641 = n16696 & n26348;
  assign n34642 = ~n34640 & ~n34641;
  assign n34643 = ~n34639 & n34642;
  assign n34644 = n54883 & ~n56543;
  assign n34645 = pi17  & ~n34644;
  assign n34646 = pi17  & ~n34643;
  assign n34647 = pi17  & ~n34646;
  assign n34648 = ~n34643 & ~n34646;
  assign n34649 = ~n34647 & ~n34648;
  assign n34650 = n34645 & ~n34649;
  assign n34651 = n34643 & n34645;
  assign n34652 = n16079 & ~n31140;
  assign n34653 = n16696 & n26343;
  assign n34654 = n54886 & ~n56543;
  assign n34655 = n16676 & n26348;
  assign n34656 = ~n34654 & ~n34655;
  assign n34657 = ~n34653 & n34656;
  assign n34658 = ~n16079 & n34657;
  assign n34659 = n31140 & n34657;
  assign n34660 = ~n34658 & ~n34659;
  assign n34661 = ~n34652 & n34657;
  assign n34662 = pi17  & ~n57691;
  assign n34663 = ~pi17  & n57691;
  assign n34664 = ~n34662 & ~n34663;
  assign n34665 = n57690 & ~n34664;
  assign n34666 = n57690 & ~n57691;
  assign n34667 = n33913 & n57692;
  assign n34668 = n16079 & n30915;
  assign n34669 = n16696 & n26340;
  assign n34670 = n54886 & n26348;
  assign n34671 = n16676 & n26343;
  assign n34672 = ~n34670 & ~n34671;
  assign n34673 = ~n34669 & n34672;
  assign n34674 = ~n34668 & n34673;
  assign n34675 = pi17  & ~n34674;
  assign n34676 = pi17  & ~n34675;
  assign n34677 = pi17  & n34674;
  assign n34678 = ~n34674 & ~n34675;
  assign n34679 = ~pi17  & ~n34674;
  assign n34680 = ~n57693 & ~n57694;
  assign n34681 = ~n33913 & ~n57692;
  assign n34682 = n57692 & ~n34667;
  assign n34683 = ~n33913 & n57692;
  assign n34684 = n33913 & ~n34667;
  assign n34685 = n33913 & ~n57692;
  assign n34686 = ~n57695 & ~n57696;
  assign n34687 = ~n34667 & ~n34681;
  assign n34688 = ~n34680 & ~n57697;
  assign n34689 = ~n34667 & ~n34688;
  assign n34690 = n34631 & ~n57689;
  assign n34691 = ~n34638 & ~n34690;
  assign n34692 = ~n34689 & n34691;
  assign n34693 = ~n34638 & ~n34692;
  assign n34694 = n34611 & ~n57687;
  assign n34695 = ~n34611 & ~n34618;
  assign n34696 = ~n34611 & ~n57687;
  assign n34697 = n57687 & ~n34618;
  assign n34698 = n34611 & n57687;
  assign n34699 = ~n57698 & ~n57699;
  assign n34700 = ~n34618 & ~n34694;
  assign n34701 = ~n34693 & ~n57700;
  assign n34702 = ~n34618 & ~n34701;
  assign n34703 = n34592 & n57684;
  assign n34704 = ~n34598 & ~n34703;
  assign n34705 = ~n34702 & n34704;
  assign n34706 = ~n34598 & ~n34705;
  assign n34707 = n34576 & ~n34578;
  assign n34708 = ~n34576 & ~n34579;
  assign n34709 = ~n34576 & ~n34578;
  assign n34710 = n34578 & ~n34579;
  assign n34711 = n34576 & n34578;
  assign n34712 = ~n57701 & ~n57702;
  assign n34713 = ~n34579 & ~n34707;
  assign n34714 = ~n34706 & ~n57703;
  assign n34715 = ~n34579 & ~n34714;
  assign n34716 = ~n34549 & n34562;
  assign n34717 = n34549 & ~n34563;
  assign n34718 = n34549 & n34562;
  assign n34719 = ~n34562 & ~n34563;
  assign n34720 = ~n34549 & ~n34562;
  assign n34721 = ~n57704 & ~n57705;
  assign n34722 = ~n34563 & ~n34716;
  assign n34723 = ~n34715 & ~n57706;
  assign n34724 = ~n34563 & ~n34723;
  assign n34725 = ~n34533 & n34546;
  assign n34726 = n34533 & ~n34547;
  assign n34727 = n34533 & n34546;
  assign n34728 = ~n34546 & ~n34547;
  assign n34729 = ~n34533 & ~n34546;
  assign n34730 = ~n57707 & ~n57708;
  assign n34731 = ~n34547 & ~n34725;
  assign n34732 = ~n34724 & ~n57709;
  assign n34733 = ~n34547 & ~n34732;
  assign n34734 = ~n34517 & n34530;
  assign n34735 = ~n34531 & ~n34734;
  assign n34736 = ~n34733 & n34735;
  assign n34737 = ~n34531 & ~n34736;
  assign n34738 = n34507 & n57677;
  assign n34739 = ~n34507 & ~n34515;
  assign n34740 = ~n57677 & ~n34515;
  assign n34741 = ~n34739 & ~n34740;
  assign n34742 = ~n34515 & ~n34738;
  assign n34743 = ~n34737 & ~n57710;
  assign n34744 = ~n34515 & ~n34743;
  assign n34745 = n34488 & n57672;
  assign n34746 = ~n34488 & ~n34494;
  assign n34747 = ~n34488 & n57672;
  assign n34748 = ~n57672 & ~n34494;
  assign n34749 = n34488 & ~n57672;
  assign n34750 = ~n57711 & ~n57712;
  assign n34751 = ~n34494 & ~n34745;
  assign n34752 = ~n34744 & ~n57713;
  assign n34753 = ~n34494 & ~n34752;
  assign n34754 = n34472 & ~n34474;
  assign n34755 = ~n34472 & ~n34475;
  assign n34756 = ~n34472 & ~n34474;
  assign n34757 = n34474 & ~n34475;
  assign n34758 = n34472 & n34474;
  assign n34759 = ~n57714 & ~n57715;
  assign n34760 = ~n34475 & ~n34754;
  assign n34761 = ~n34753 & ~n57716;
  assign n34762 = ~n34475 & ~n34761;
  assign n34763 = ~n34445 & n34458;
  assign n34764 = n34445 & ~n34459;
  assign n34765 = n34445 & n34458;
  assign n34766 = ~n34458 & ~n34459;
  assign n34767 = ~n34445 & ~n34458;
  assign n34768 = ~n57717 & ~n57718;
  assign n34769 = ~n34459 & ~n34763;
  assign n34770 = ~n34762 & ~n57719;
  assign n34771 = ~n34459 & ~n34770;
  assign n34772 = ~n34429 & n34442;
  assign n34773 = ~n34443 & ~n34772;
  assign n34774 = ~n34771 & n34773;
  assign n34775 = ~n34443 & ~n34774;
  assign n34776 = n34419 & n57665;
  assign n34777 = ~n34419 & ~n34427;
  assign n34778 = ~n57665 & ~n34427;
  assign n34779 = ~n34777 & ~n34778;
  assign n34780 = ~n34427 & ~n34776;
  assign n34781 = ~n34775 & ~n57720;
  assign n34782 = ~n34427 & ~n34781;
  assign n34783 = n34398 & n57660;
  assign n34784 = ~n34398 & ~n34406;
  assign n34785 = ~n57660 & ~n34406;
  assign n34786 = ~n34784 & ~n34785;
  assign n34787 = ~n34406 & ~n34783;
  assign n34788 = ~n34782 & ~n57721;
  assign n34789 = ~n34406 & ~n34788;
  assign n34790 = n34379 & n57655;
  assign n34791 = ~n34379 & ~n34385;
  assign n34792 = ~n34379 & n57655;
  assign n34793 = ~n57655 & ~n34385;
  assign n34794 = n34379 & ~n57655;
  assign n34795 = ~n57722 & ~n57723;
  assign n34796 = ~n34385 & ~n34790;
  assign n34797 = ~n34789 & ~n57724;
  assign n34798 = ~n34385 & ~n34797;
  assign n34799 = n34360 & n57652;
  assign n34800 = ~n34360 & ~n34366;
  assign n34801 = ~n34360 & n57652;
  assign n34802 = ~n57652 & ~n34366;
  assign n34803 = n34360 & ~n57652;
  assign n34804 = ~n57725 & ~n57726;
  assign n34805 = ~n34366 & ~n34799;
  assign n34806 = ~n34798 & ~n57727;
  assign n34807 = ~n34366 & ~n34806;
  assign n34808 = n34341 & n57649;
  assign n34809 = ~n34341 & ~n34347;
  assign n34810 = ~n34341 & n57649;
  assign n34811 = ~n57649 & ~n34347;
  assign n34812 = n34341 & ~n57649;
  assign n34813 = ~n57728 & ~n57729;
  assign n34814 = ~n34347 & ~n34808;
  assign n34815 = ~n34807 & ~n57730;
  assign n34816 = ~n34347 & ~n34815;
  assign n34817 = n34320 & n57646;
  assign n34818 = ~n34320 & ~n34328;
  assign n34819 = ~n57646 & ~n34328;
  assign n34820 = ~n34818 & ~n34819;
  assign n34821 = ~n34328 & ~n34817;
  assign n34822 = ~n34816 & ~n57731;
  assign n34823 = ~n34328 & ~n34822;
  assign n34824 = n34299 & n57641;
  assign n34825 = ~n34299 & ~n34307;
  assign n34826 = ~n57641 & ~n34307;
  assign n34827 = ~n34825 & ~n34826;
  assign n34828 = ~n34307 & ~n34824;
  assign n34829 = ~n34823 & ~n57732;
  assign n34830 = ~n34307 & ~n34829;
  assign n34831 = n34278 & n57636;
  assign n34832 = ~n34278 & ~n34286;
  assign n34833 = ~n57636 & ~n34286;
  assign n34834 = ~n34832 & ~n34833;
  assign n34835 = ~n34286 & ~n34831;
  assign n34836 = ~n34830 & ~n57733;
  assign n34837 = ~n34286 & ~n34836;
  assign n34838 = n34257 & n57631;
  assign n34839 = ~n34257 & ~n34265;
  assign n34840 = ~n57631 & ~n34265;
  assign n34841 = ~n34839 & ~n34840;
  assign n34842 = ~n34265 & ~n34838;
  assign n34843 = ~n34837 & ~n57734;
  assign n34844 = ~n34265 & ~n34843;
  assign n34845 = n34241 & ~n34243;
  assign n34846 = ~n34241 & ~n34244;
  assign n34847 = ~n34241 & ~n34243;
  assign n34848 = n34243 & ~n34244;
  assign n34849 = n34241 & n34243;
  assign n34850 = ~n57735 & ~n57736;
  assign n34851 = ~n34244 & ~n34845;
  assign n34852 = ~n34844 & ~n57737;
  assign n34853 = ~n34244 & ~n34852;
  assign n34854 = n34129 & ~n34130;
  assign n34855 = n34127 & n34129;
  assign n34856 = ~n34127 & ~n34130;
  assign n34857 = ~n34127 & ~n34129;
  assign n34858 = n34127 & ~n34129;
  assign n34859 = ~n34130 & ~n34858;
  assign n34860 = ~n57738 & ~n57739;
  assign n34861 = ~n34853 & n57740;
  assign n34862 = n34853 & ~n57740;
  assign n34863 = n17265 & n27466;
  assign n34864 = n18588 & n26262;
  assign n34865 = n55041 & n26268;
  assign n34866 = n18556 & n26265;
  assign n34867 = ~n34865 & ~n34866;
  assign n34868 = ~n34864 & n34867;
  assign n34869 = ~n34863 & n34868;
  assign n34870 = pi14  & ~n34869;
  assign n34871 = pi14  & ~n34870;
  assign n34872 = pi14  & n34869;
  assign n34873 = ~n34869 & ~n34870;
  assign n34874 = ~pi14  & ~n34869;
  assign n34875 = ~n57741 & ~n57742;
  assign n34876 = ~n34862 & ~n34875;
  assign n34877 = ~n34861 & ~n34862;
  assign n34878 = ~n34875 & n34877;
  assign n34879 = ~n34861 & ~n34878;
  assign n34880 = ~n34861 & ~n34876;
  assign n34881 = ~n57624 & ~n57743;
  assign n34882 = n57624 & n57743;
  assign n34883 = n18846 & n27491;
  assign n34884 = n19541 & n26250;
  assign n34885 = n55247 & n26256;
  assign n34886 = n19509 & n26253;
  assign n34887 = ~n34885 & ~n34886;
  assign n34888 = ~n34884 & n34887;
  assign n34889 = ~n34883 & n34888;
  assign n34890 = pi11  & ~n34889;
  assign n34891 = pi11  & ~n34890;
  assign n34892 = pi11  & n34889;
  assign n34893 = ~n34889 & ~n34890;
  assign n34894 = ~pi11  & ~n34889;
  assign n34895 = ~n57744 & ~n57745;
  assign n34896 = ~n34882 & ~n34895;
  assign n34897 = ~n34881 & ~n34882;
  assign n34898 = ~n34895 & n34897;
  assign n34899 = ~n34881 & ~n34898;
  assign n34900 = ~n34881 & ~n34896;
  assign n34901 = ~n57623 & ~n57746;
  assign n34902 = n57623 & n57746;
  assign n34903 = n20085 & ~n56564;
  assign n34904 = n21269 & ~n26537;
  assign n34905 = n55472 & n26244;
  assign n34906 = n21237 & n26242;
  assign n34907 = ~n34905 & ~n34906;
  assign n34908 = ~n34904 & n34907;
  assign n34909 = ~n34903 & n34908;
  assign n34910 = pi8  & ~n34909;
  assign n34911 = pi8  & ~n34910;
  assign n34912 = pi8  & n34909;
  assign n34913 = ~n34909 & ~n34910;
  assign n34914 = ~pi8  & ~n34909;
  assign n34915 = ~n57747 & ~n57748;
  assign n34916 = ~n34902 & ~n34915;
  assign n34917 = ~n34901 & ~n34902;
  assign n34918 = ~n34915 & n34917;
  assign n34919 = ~n34901 & ~n34918;
  assign n34920 = ~n34901 & ~n34916;
  assign n34921 = ~n34218 & ~n57749;
  assign n34922 = n57520 & n57612;
  assign n34923 = ~n34173 & ~n34922;
  assign n34924 = n34218 & n57749;
  assign n34925 = ~n57749 & ~n34921;
  assign n34926 = n34218 & ~n57749;
  assign n34927 = ~n34218 & ~n34921;
  assign n34928 = ~n34218 & n57749;
  assign n34929 = ~n57750 & ~n57751;
  assign n34930 = ~n34921 & ~n34924;
  assign n34931 = n34923 & ~n57752;
  assign n34932 = ~n34921 & ~n34931;
  assign n34933 = n34196 & ~n34198;
  assign n34934 = n34198 & ~n34199;
  assign n34935 = ~n34196 & ~n34199;
  assign n34936 = ~n34934 & ~n34935;
  assign n34937 = ~n34199 & ~n34933;
  assign n34938 = ~n34932 & ~n57753;
  assign n34939 = ~n34923 & n57752;
  assign n34940 = ~n34931 & ~n34939;
  assign n34941 = n34895 & ~n34897;
  assign n34942 = n34897 & ~n34898;
  assign n34943 = ~n34895 & ~n34898;
  assign n34944 = ~n34942 & ~n34943;
  assign n34945 = ~n34898 & ~n34941;
  assign n34946 = n34844 & n57737;
  assign n34947 = ~n34852 & ~n34946;
  assign n34948 = n17265 & n27042;
  assign n34949 = n18588 & n26265;
  assign n34950 = n55041 & n26271;
  assign n34951 = n18556 & n26268;
  assign n34952 = ~n34950 & ~n34951;
  assign n34953 = ~n34949 & n34952;
  assign n34954 = ~n17265 & n34953;
  assign n34955 = ~n27042 & n34953;
  assign n34956 = ~n34954 & ~n34955;
  assign n34957 = ~n34948 & n34953;
  assign n34958 = pi14  & ~n57755;
  assign n34959 = ~pi14  & n57755;
  assign n34960 = ~n34958 & ~n34959;
  assign n34961 = n34947 & ~n34960;
  assign n34962 = n34837 & n57734;
  assign n34963 = ~n34843 & ~n34962;
  assign n34964 = n17265 & ~n56601;
  assign n34965 = n18588 & n26268;
  assign n34966 = n55041 & n26274;
  assign n34967 = n18556 & n26271;
  assign n34968 = ~n34966 & ~n34967;
  assign n34969 = ~n34965 & n34968;
  assign n34970 = ~n17265 & n34969;
  assign n34971 = n56601 & n34969;
  assign n34972 = ~n34970 & ~n34971;
  assign n34973 = ~n34964 & n34969;
  assign n34974 = pi14  & ~n57756;
  assign n34975 = ~pi14  & n57756;
  assign n34976 = ~n34974 & ~n34975;
  assign n34977 = n34963 & ~n34976;
  assign n34978 = n34830 & n57733;
  assign n34979 = ~n34836 & ~n34978;
  assign n34980 = n17265 & ~n56612;
  assign n34981 = n18588 & n26271;
  assign n34982 = n55041 & n26277;
  assign n34983 = n18556 & n26274;
  assign n34984 = ~n34982 & ~n34983;
  assign n34985 = ~n34981 & n34984;
  assign n34986 = ~n17265 & n34985;
  assign n34987 = n56612 & n34985;
  assign n34988 = ~n34986 & ~n34987;
  assign n34989 = ~n34980 & n34985;
  assign n34990 = pi14  & ~n57757;
  assign n34991 = ~pi14  & n57757;
  assign n34992 = ~n34990 & ~n34991;
  assign n34993 = n34979 & ~n34992;
  assign n34994 = n34823 & n57732;
  assign n34995 = ~n34829 & ~n34994;
  assign n34996 = n17265 & ~n56648;
  assign n34997 = n18588 & n26274;
  assign n34998 = n55041 & n26280;
  assign n34999 = n18556 & n26277;
  assign n35000 = ~n34998 & ~n34999;
  assign n35001 = ~n34997 & n35000;
  assign n35002 = ~n17265 & n35001;
  assign n35003 = n56648 & n35001;
  assign n35004 = ~n35002 & ~n35003;
  assign n35005 = ~n34996 & n35001;
  assign n35006 = pi14  & ~n57758;
  assign n35007 = ~pi14  & n57758;
  assign n35008 = ~n35006 & ~n35007;
  assign n35009 = n34995 & ~n35008;
  assign n35010 = n34816 & n57731;
  assign n35011 = ~n34822 & ~n35010;
  assign n35012 = n17265 & n27330;
  assign n35013 = n18588 & n26277;
  assign n35014 = n55041 & n26283;
  assign n35015 = n18556 & n26280;
  assign n35016 = ~n35014 & ~n35015;
  assign n35017 = ~n35013 & n35016;
  assign n35018 = ~n17265 & n35017;
  assign n35019 = ~n27330 & n35017;
  assign n35020 = ~n35018 & ~n35019;
  assign n35021 = ~n35012 & n35017;
  assign n35022 = pi14  & ~n57759;
  assign n35023 = ~pi14  & n57759;
  assign n35024 = ~n35022 & ~n35023;
  assign n35025 = n35011 & ~n35024;
  assign n35026 = n34807 & n57730;
  assign n35027 = ~n34815 & ~n35026;
  assign n35028 = n17265 & n27743;
  assign n35029 = n18588 & n26280;
  assign n35030 = n55041 & n26286;
  assign n35031 = n18556 & n26283;
  assign n35032 = ~n35030 & ~n35031;
  assign n35033 = ~n35029 & n35032;
  assign n35034 = ~n17265 & n35033;
  assign n35035 = ~n27743 & n35033;
  assign n35036 = ~n35034 & ~n35035;
  assign n35037 = ~n35028 & n35033;
  assign n35038 = pi14  & ~n57760;
  assign n35039 = ~pi14  & n57760;
  assign n35040 = ~n35038 & ~n35039;
  assign n35041 = n35027 & ~n35040;
  assign n35042 = n34798 & n57727;
  assign n35043 = ~n34806 & ~n35042;
  assign n35044 = n17265 & ~n56686;
  assign n35045 = n18588 & n26283;
  assign n35046 = n55041 & n26289;
  assign n35047 = n18556 & n26286;
  assign n35048 = ~n35046 & ~n35047;
  assign n35049 = ~n35045 & n35048;
  assign n35050 = ~n17265 & n35049;
  assign n35051 = n56686 & n35049;
  assign n35052 = ~n35050 & ~n35051;
  assign n35053 = ~n35044 & n35049;
  assign n35054 = pi14  & ~n57761;
  assign n35055 = ~pi14  & n57761;
  assign n35056 = ~n35054 & ~n35055;
  assign n35057 = n35043 & ~n35056;
  assign n35058 = n34789 & n57724;
  assign n35059 = ~n34797 & ~n35058;
  assign n35060 = n17265 & ~n56721;
  assign n35061 = n18588 & n26286;
  assign n35062 = n55041 & n26292;
  assign n35063 = n18556 & n26289;
  assign n35064 = ~n35062 & ~n35063;
  assign n35065 = ~n35061 & n35064;
  assign n35066 = ~n17265 & n35065;
  assign n35067 = n56721 & n35065;
  assign n35068 = ~n35066 & ~n35067;
  assign n35069 = ~n35060 & n35065;
  assign n35070 = pi14  & ~n57762;
  assign n35071 = ~pi14  & n57762;
  assign n35072 = ~n35070 & ~n35071;
  assign n35073 = n35059 & ~n35072;
  assign n35074 = n34782 & n57721;
  assign n35075 = ~n34788 & ~n35074;
  assign n35076 = n17265 & n28107;
  assign n35077 = n18588 & n26289;
  assign n35078 = n55041 & n26295;
  assign n35079 = n18556 & n26292;
  assign n35080 = ~n35078 & ~n35079;
  assign n35081 = ~n35077 & n35080;
  assign n35082 = ~n17265 & n35081;
  assign n35083 = ~n28107 & n35081;
  assign n35084 = ~n35082 & ~n35083;
  assign n35085 = ~n35076 & n35081;
  assign n35086 = pi14  & ~n57763;
  assign n35087 = ~pi14  & n57763;
  assign n35088 = ~n35086 & ~n35087;
  assign n35089 = n35075 & ~n35088;
  assign n35090 = n34775 & n57720;
  assign n35091 = ~n34781 & ~n35090;
  assign n35092 = n17265 & n28808;
  assign n35093 = n18588 & n26292;
  assign n35094 = n55041 & n26298;
  assign n35095 = n18556 & n26295;
  assign n35096 = ~n35094 & ~n35095;
  assign n35097 = ~n35093 & n35096;
  assign n35098 = ~n17265 & n35097;
  assign n35099 = ~n28808 & n35097;
  assign n35100 = ~n35098 & ~n35099;
  assign n35101 = ~n35092 & n35097;
  assign n35102 = pi14  & ~n57764;
  assign n35103 = ~pi14  & n57764;
  assign n35104 = ~n35102 & ~n35103;
  assign n35105 = n35091 & ~n35104;
  assign n35106 = n17265 & n28493;
  assign n35107 = n18588 & n26295;
  assign n35108 = n55041 & n26301;
  assign n35109 = n18556 & n26298;
  assign n35110 = ~n35108 & ~n35109;
  assign n35111 = ~n35107 & n35110;
  assign n35112 = ~n35106 & n35111;
  assign n35113 = pi14  & ~n35112;
  assign n35114 = ~n35112 & ~n35113;
  assign n35115 = ~pi14  & ~n35112;
  assign n35116 = pi14  & ~n35113;
  assign n35117 = pi14  & n35112;
  assign n35118 = ~n57765 & ~n57766;
  assign n35119 = n34771 & ~n34773;
  assign n35120 = ~n34774 & ~n35119;
  assign n35121 = ~n35118 & n35120;
  assign n35122 = n17265 & ~n56870;
  assign n35123 = n18588 & n26298;
  assign n35124 = n55041 & n26304;
  assign n35125 = n18556 & n26301;
  assign n35126 = ~n35124 & ~n35125;
  assign n35127 = ~n35123 & n35126;
  assign n35128 = ~n35122 & n35127;
  assign n35129 = pi14  & ~n35128;
  assign n35130 = ~n35128 & ~n35129;
  assign n35131 = ~pi14  & ~n35128;
  assign n35132 = pi14  & ~n35129;
  assign n35133 = pi14  & n35128;
  assign n35134 = ~n57767 & ~n57768;
  assign n35135 = n34762 & n57719;
  assign n35136 = ~n34762 & ~n34770;
  assign n35137 = ~n57719 & ~n34770;
  assign n35138 = ~n35136 & ~n35137;
  assign n35139 = ~n34770 & ~n35135;
  assign n35140 = ~n35134 & ~n57769;
  assign n35141 = n34753 & n57716;
  assign n35142 = ~n34761 & ~n35141;
  assign n35143 = n17265 & n29446;
  assign n35144 = n18588 & n26301;
  assign n35145 = n55041 & n26307;
  assign n35146 = n18556 & n26304;
  assign n35147 = ~n35145 & ~n35146;
  assign n35148 = ~n35144 & n35147;
  assign n35149 = ~n17265 & n35148;
  assign n35150 = ~n29446 & n35148;
  assign n35151 = ~n35149 & ~n35150;
  assign n35152 = ~n35143 & n35148;
  assign n35153 = pi14  & ~n57770;
  assign n35154 = ~pi14  & n57770;
  assign n35155 = ~n35153 & ~n35154;
  assign n35156 = n35142 & ~n35155;
  assign n35157 = n34744 & n57713;
  assign n35158 = ~n34752 & ~n35157;
  assign n35159 = n17265 & ~n56867;
  assign n35160 = n18588 & n26304;
  assign n35161 = n55041 & n26310;
  assign n35162 = n18556 & n26307;
  assign n35163 = ~n35161 & ~n35162;
  assign n35164 = ~n35160 & n35163;
  assign n35165 = ~n17265 & n35164;
  assign n35166 = n56867 & n35164;
  assign n35167 = ~n35165 & ~n35166;
  assign n35168 = ~n35159 & n35164;
  assign n35169 = pi14  & ~n57771;
  assign n35170 = ~pi14  & n57771;
  assign n35171 = ~n35169 & ~n35170;
  assign n35172 = n35158 & ~n35171;
  assign n35173 = n34737 & n57710;
  assign n35174 = ~n34743 & ~n35173;
  assign n35175 = n17265 & ~n56928;
  assign n35176 = n18588 & n26307;
  assign n35177 = n55041 & n26313;
  assign n35178 = n18556 & n26310;
  assign n35179 = ~n35177 & ~n35178;
  assign n35180 = ~n35176 & n35179;
  assign n35181 = ~n17265 & n35180;
  assign n35182 = n56928 & n35180;
  assign n35183 = ~n35181 & ~n35182;
  assign n35184 = ~n35175 & n35180;
  assign n35185 = pi14  & ~n57772;
  assign n35186 = ~pi14  & n57772;
  assign n35187 = ~n35185 & ~n35186;
  assign n35188 = n35174 & ~n35187;
  assign n35189 = n17265 & ~n57002;
  assign n35190 = n18588 & n26310;
  assign n35191 = n55041 & n26316;
  assign n35192 = n18556 & n26313;
  assign n35193 = ~n35191 & ~n35192;
  assign n35194 = ~n35190 & n35193;
  assign n35195 = ~n35189 & n35194;
  assign n35196 = pi14  & ~n35195;
  assign n35197 = ~n35195 & ~n35196;
  assign n35198 = ~pi14  & ~n35195;
  assign n35199 = pi14  & ~n35196;
  assign n35200 = pi14  & n35195;
  assign n35201 = ~n57773 & ~n57774;
  assign n35202 = n34733 & ~n34735;
  assign n35203 = ~n34736 & ~n35202;
  assign n35204 = ~n35201 & n35203;
  assign n35205 = n17265 & n30192;
  assign n35206 = n18588 & n26313;
  assign n35207 = n55041 & n26319;
  assign n35208 = n18556 & n26316;
  assign n35209 = ~n35207 & ~n35208;
  assign n35210 = ~n35206 & n35209;
  assign n35211 = ~n35205 & n35210;
  assign n35212 = pi14  & ~n35211;
  assign n35213 = ~n35211 & ~n35212;
  assign n35214 = ~pi14  & ~n35211;
  assign n35215 = pi14  & ~n35212;
  assign n35216 = pi14  & n35211;
  assign n35217 = ~n57775 & ~n57776;
  assign n35218 = n34724 & n57709;
  assign n35219 = ~n34724 & ~n34732;
  assign n35220 = ~n57709 & ~n34732;
  assign n35221 = ~n35219 & ~n35220;
  assign n35222 = ~n34732 & ~n35218;
  assign n35223 = ~n35217 & ~n57777;
  assign n35224 = n17265 & ~n56920;
  assign n35225 = n18588 & n26316;
  assign n35226 = n55041 & n26322;
  assign n35227 = n18556 & n26319;
  assign n35228 = ~n35226 & ~n35227;
  assign n35229 = ~n35225 & n35228;
  assign n35230 = ~n35224 & n35229;
  assign n35231 = pi14  & ~n35230;
  assign n35232 = ~n35230 & ~n35231;
  assign n35233 = ~pi14  & ~n35230;
  assign n35234 = pi14  & ~n35231;
  assign n35235 = pi14  & n35230;
  assign n35236 = ~n57778 & ~n57779;
  assign n35237 = n34715 & n57706;
  assign n35238 = ~n34715 & ~n34723;
  assign n35239 = ~n34715 & n57706;
  assign n35240 = ~n57706 & ~n34723;
  assign n35241 = n34715 & ~n57706;
  assign n35242 = ~n57780 & ~n57781;
  assign n35243 = ~n34723 & ~n35237;
  assign n35244 = ~n35236 & ~n57782;
  assign n35245 = n34706 & n57703;
  assign n35246 = ~n34714 & ~n35245;
  assign n35247 = n17265 & n30264;
  assign n35248 = n18588 & n26319;
  assign n35249 = n55041 & n26325;
  assign n35250 = n18556 & n26322;
  assign n35251 = ~n35249 & ~n35250;
  assign n35252 = ~n35248 & n35251;
  assign n35253 = ~n17265 & n35252;
  assign n35254 = ~n30264 & n35252;
  assign n35255 = ~n35253 & ~n35254;
  assign n35256 = ~n35247 & n35252;
  assign n35257 = pi14  & ~n57783;
  assign n35258 = ~pi14  & n57783;
  assign n35259 = ~n35257 & ~n35258;
  assign n35260 = n35246 & ~n35259;
  assign n35261 = n34702 & ~n34704;
  assign n35262 = ~n34705 & ~n35261;
  assign n35263 = n17265 & ~n57012;
  assign n35264 = n18588 & n26322;
  assign n35265 = n55041 & n26328;
  assign n35266 = n18556 & n26325;
  assign n35267 = ~n35265 & ~n35266;
  assign n35268 = ~n35264 & n35267;
  assign n35269 = ~n17265 & n35268;
  assign n35270 = n57012 & n35268;
  assign n35271 = ~n35269 & ~n35270;
  assign n35272 = ~n35263 & n35268;
  assign n35273 = pi14  & ~n57784;
  assign n35274 = ~pi14  & n57784;
  assign n35275 = ~n35273 & ~n35274;
  assign n35276 = n35262 & ~n35275;
  assign n35277 = n34693 & n57700;
  assign n35278 = ~n34701 & ~n35277;
  assign n35279 = n17265 & ~n57017;
  assign n35280 = n18588 & n26325;
  assign n35281 = n55041 & n26331;
  assign n35282 = n18556 & n26328;
  assign n35283 = ~n35281 & ~n35282;
  assign n35284 = ~n35280 & n35283;
  assign n35285 = ~n17265 & n35284;
  assign n35286 = n57017 & n35284;
  assign n35287 = ~n35285 & ~n35286;
  assign n35288 = ~n35279 & n35284;
  assign n35289 = pi14  & ~n57785;
  assign n35290 = ~pi14  & n57785;
  assign n35291 = ~n35289 & ~n35290;
  assign n35292 = n35278 & ~n35291;
  assign n35293 = n17265 & n30470;
  assign n35294 = n18588 & n26328;
  assign n35295 = n55041 & n26334;
  assign n35296 = n18556 & n26331;
  assign n35297 = ~n35295 & ~n35296;
  assign n35298 = ~n35294 & n35297;
  assign n35299 = ~n35293 & n35298;
  assign n35300 = pi14  & ~n35299;
  assign n35301 = ~n35299 & ~n35300;
  assign n35302 = ~pi14  & ~n35299;
  assign n35303 = pi14  & ~n35300;
  assign n35304 = pi14  & n35299;
  assign n35305 = ~n57786 & ~n57787;
  assign n35306 = n34689 & ~n34691;
  assign n35307 = ~n34692 & ~n35306;
  assign n35308 = ~n35305 & n35307;
  assign n35309 = n17265 & ~n57033;
  assign n35310 = n18588 & n26331;
  assign n35311 = n55041 & n26337;
  assign n35312 = n18556 & n26334;
  assign n35313 = ~n35311 & ~n35312;
  assign n35314 = ~n35310 & n35313;
  assign n35315 = ~n17265 & n35314;
  assign n35316 = n57033 & n35314;
  assign n35317 = ~n35315 & ~n35316;
  assign n35318 = ~n35309 & n35314;
  assign n35319 = pi14  & ~n57788;
  assign n35320 = ~pi14  & n57788;
  assign n35321 = ~n35319 & ~n35320;
  assign n35322 = n34680 & n57697;
  assign n35323 = ~n57697 & ~n34688;
  assign n35324 = ~n34680 & ~n34688;
  assign n35325 = ~n35323 & ~n35324;
  assign n35326 = ~n34688 & ~n35322;
  assign n35327 = ~n35321 & ~n57789;
  assign n35328 = n17265 & ~n57042;
  assign n35329 = n18588 & n26334;
  assign n35330 = n55041 & n26340;
  assign n35331 = n18556 & n26337;
  assign n35332 = ~n35330 & ~n35331;
  assign n35333 = ~n35329 & n35332;
  assign n35334 = ~n35328 & n35333;
  assign n35335 = pi14  & ~n35334;
  assign n35336 = ~n35334 & ~n35335;
  assign n35337 = ~pi14  & ~n35334;
  assign n35338 = pi14  & ~n35335;
  assign n35339 = pi14  & n35334;
  assign n35340 = ~n57790 & ~n57791;
  assign n35341 = pi17  & ~n57690;
  assign n35342 = ~n57691 & ~n35341;
  assign n35343 = n57691 & n35341;
  assign n35344 = ~n57690 & n34664;
  assign n35345 = ~n57692 & ~n35344;
  assign n35346 = ~n35342 & ~n35343;
  assign n35347 = ~n35340 & n57792;
  assign n35348 = n17265 & n30866;
  assign n35349 = n18588 & n26337;
  assign n35350 = n55041 & n26343;
  assign n35351 = n18556 & n26340;
  assign n35352 = ~n35350 & ~n35351;
  assign n35353 = ~n35349 & n35352;
  assign n35354 = ~n17265 & n35353;
  assign n35355 = ~n30866 & n35353;
  assign n35356 = ~n35354 & ~n35355;
  assign n35357 = ~n35348 & n35353;
  assign n35358 = pi14  & ~n57793;
  assign n35359 = ~pi14  & n57793;
  assign n35360 = ~n35358 & ~n35359;
  assign n35361 = pi17  & n34644;
  assign n35362 = ~n34643 & n35361;
  assign n35363 = n34643 & ~n35361;
  assign n35364 = ~n34645 & n34649;
  assign n35365 = ~n57690 & ~n35364;
  assign n35366 = ~n35362 & ~n35363;
  assign n35367 = ~n35360 & n57794;
  assign n35368 = n17265 & ~n31019;
  assign n35369 = n18556 & ~n56543;
  assign n35370 = n18588 & n26348;
  assign n35371 = ~n35369 & ~n35370;
  assign n35372 = ~n35368 & n35371;
  assign n35373 = n55039 & ~n56543;
  assign n35374 = pi14  & ~n35373;
  assign n35375 = pi14  & ~n35372;
  assign n35376 = pi14  & ~n35375;
  assign n35377 = ~n35372 & ~n35375;
  assign n35378 = ~n35376 & ~n35377;
  assign n35379 = n35374 & ~n35378;
  assign n35380 = n35372 & n35374;
  assign n35381 = n17265 & ~n31140;
  assign n35382 = n18588 & n26343;
  assign n35383 = n55041 & ~n56543;
  assign n35384 = n18556 & n26348;
  assign n35385 = ~n35383 & ~n35384;
  assign n35386 = ~n35382 & n35385;
  assign n35387 = ~n17265 & n35386;
  assign n35388 = n31140 & n35386;
  assign n35389 = ~n35387 & ~n35388;
  assign n35390 = ~n35381 & n35386;
  assign n35391 = pi14  & ~n57796;
  assign n35392 = ~pi14  & n57796;
  assign n35393 = ~n35391 & ~n35392;
  assign n35394 = n57795 & ~n35393;
  assign n35395 = n57795 & ~n57796;
  assign n35396 = n34644 & n57797;
  assign n35397 = n17265 & n30915;
  assign n35398 = n18588 & n26340;
  assign n35399 = n55041 & n26348;
  assign n35400 = n18556 & n26343;
  assign n35401 = ~n35399 & ~n35400;
  assign n35402 = ~n35398 & n35401;
  assign n35403 = ~n35397 & n35402;
  assign n35404 = pi14  & ~n35403;
  assign n35405 = pi14  & ~n35404;
  assign n35406 = pi14  & n35403;
  assign n35407 = ~n35403 & ~n35404;
  assign n35408 = ~pi14  & ~n35403;
  assign n35409 = ~n57798 & ~n57799;
  assign n35410 = ~n34644 & ~n57797;
  assign n35411 = n57797 & ~n35396;
  assign n35412 = ~n34644 & n57797;
  assign n35413 = n34644 & ~n35396;
  assign n35414 = n34644 & ~n57797;
  assign n35415 = ~n57800 & ~n57801;
  assign n35416 = ~n35396 & ~n35410;
  assign n35417 = ~n35409 & ~n57802;
  assign n35418 = ~n35396 & ~n35417;
  assign n35419 = n35360 & ~n57794;
  assign n35420 = ~n35367 & ~n35419;
  assign n35421 = ~n35418 & n35420;
  assign n35422 = ~n35367 & ~n35421;
  assign n35423 = n35340 & ~n57792;
  assign n35424 = ~n35340 & ~n35347;
  assign n35425 = ~n35340 & ~n57792;
  assign n35426 = n57792 & ~n35347;
  assign n35427 = n35340 & n57792;
  assign n35428 = ~n57803 & ~n57804;
  assign n35429 = ~n35347 & ~n35423;
  assign n35430 = ~n35422 & ~n57805;
  assign n35431 = ~n35347 & ~n35430;
  assign n35432 = n35321 & n57789;
  assign n35433 = ~n35327 & ~n35432;
  assign n35434 = ~n35431 & n35433;
  assign n35435 = ~n35327 & ~n35434;
  assign n35436 = n35305 & ~n35307;
  assign n35437 = ~n35305 & ~n35308;
  assign n35438 = ~n35305 & ~n35307;
  assign n35439 = n35307 & ~n35308;
  assign n35440 = n35305 & n35307;
  assign n35441 = ~n57806 & ~n57807;
  assign n35442 = ~n35308 & ~n35436;
  assign n35443 = ~n35435 & ~n57808;
  assign n35444 = ~n35308 & ~n35443;
  assign n35445 = ~n35278 & n35291;
  assign n35446 = n35278 & ~n35292;
  assign n35447 = n35278 & n35291;
  assign n35448 = ~n35291 & ~n35292;
  assign n35449 = ~n35278 & ~n35291;
  assign n35450 = ~n57809 & ~n57810;
  assign n35451 = ~n35292 & ~n35445;
  assign n35452 = ~n35444 & ~n57811;
  assign n35453 = ~n35292 & ~n35452;
  assign n35454 = ~n35262 & n35275;
  assign n35455 = n35262 & ~n35276;
  assign n35456 = n35262 & n35275;
  assign n35457 = ~n35275 & ~n35276;
  assign n35458 = ~n35262 & ~n35275;
  assign n35459 = ~n57812 & ~n57813;
  assign n35460 = ~n35276 & ~n35454;
  assign n35461 = ~n35453 & ~n57814;
  assign n35462 = ~n35276 & ~n35461;
  assign n35463 = ~n35246 & n35259;
  assign n35464 = ~n35260 & ~n35463;
  assign n35465 = ~n35462 & n35464;
  assign n35466 = ~n35260 & ~n35465;
  assign n35467 = n35236 & n57782;
  assign n35468 = ~n35236 & ~n35244;
  assign n35469 = ~n57782 & ~n35244;
  assign n35470 = ~n35468 & ~n35469;
  assign n35471 = ~n35244 & ~n35467;
  assign n35472 = ~n35466 & ~n57815;
  assign n35473 = ~n35244 & ~n35472;
  assign n35474 = n35217 & n57777;
  assign n35475 = ~n35217 & ~n35223;
  assign n35476 = ~n35217 & n57777;
  assign n35477 = ~n57777 & ~n35223;
  assign n35478 = n35217 & ~n57777;
  assign n35479 = ~n57816 & ~n57817;
  assign n35480 = ~n35223 & ~n35474;
  assign n35481 = ~n35473 & ~n57818;
  assign n35482 = ~n35223 & ~n35481;
  assign n35483 = n35201 & ~n35203;
  assign n35484 = ~n35201 & ~n35204;
  assign n35485 = ~n35201 & ~n35203;
  assign n35486 = n35203 & ~n35204;
  assign n35487 = n35201 & n35203;
  assign n35488 = ~n57819 & ~n57820;
  assign n35489 = ~n35204 & ~n35483;
  assign n35490 = ~n35482 & ~n57821;
  assign n35491 = ~n35204 & ~n35490;
  assign n35492 = ~n35174 & n35187;
  assign n35493 = n35174 & ~n35188;
  assign n35494 = n35174 & n35187;
  assign n35495 = ~n35187 & ~n35188;
  assign n35496 = ~n35174 & ~n35187;
  assign n35497 = ~n57822 & ~n57823;
  assign n35498 = ~n35188 & ~n35492;
  assign n35499 = ~n35491 & ~n57824;
  assign n35500 = ~n35188 & ~n35499;
  assign n35501 = ~n35158 & n35171;
  assign n35502 = n35158 & ~n35172;
  assign n35503 = n35158 & n35171;
  assign n35504 = ~n35171 & ~n35172;
  assign n35505 = ~n35158 & ~n35171;
  assign n35506 = ~n57825 & ~n57826;
  assign n35507 = ~n35172 & ~n35501;
  assign n35508 = ~n35500 & ~n57827;
  assign n35509 = ~n35172 & ~n35508;
  assign n35510 = ~n35142 & n35155;
  assign n35511 = ~n35156 & ~n35510;
  assign n35512 = ~n35509 & n35511;
  assign n35513 = ~n35156 & ~n35512;
  assign n35514 = n35134 & n57769;
  assign n35515 = ~n35134 & ~n35140;
  assign n35516 = ~n35134 & n57769;
  assign n35517 = ~n57769 & ~n35140;
  assign n35518 = n35134 & ~n57769;
  assign n35519 = ~n57828 & ~n57829;
  assign n35520 = ~n35140 & ~n35514;
  assign n35521 = ~n35513 & ~n57830;
  assign n35522 = ~n35140 & ~n35521;
  assign n35523 = n35118 & ~n35120;
  assign n35524 = ~n35118 & ~n35121;
  assign n35525 = ~n35118 & ~n35120;
  assign n35526 = n35120 & ~n35121;
  assign n35527 = n35118 & n35120;
  assign n35528 = ~n57831 & ~n57832;
  assign n35529 = ~n35121 & ~n35523;
  assign n35530 = ~n35522 & ~n57833;
  assign n35531 = ~n35121 & ~n35530;
  assign n35532 = ~n35091 & n35104;
  assign n35533 = n35091 & ~n35105;
  assign n35534 = n35091 & n35104;
  assign n35535 = ~n35104 & ~n35105;
  assign n35536 = ~n35091 & ~n35104;
  assign n35537 = ~n57834 & ~n57835;
  assign n35538 = ~n35105 & ~n35532;
  assign n35539 = ~n35531 & ~n57836;
  assign n35540 = ~n35105 & ~n35539;
  assign n35541 = ~n35075 & n35088;
  assign n35542 = n35075 & ~n35089;
  assign n35543 = n35075 & n35088;
  assign n35544 = ~n35088 & ~n35089;
  assign n35545 = ~n35075 & ~n35088;
  assign n35546 = ~n57837 & ~n57838;
  assign n35547 = ~n35089 & ~n35541;
  assign n35548 = ~n35540 & ~n57839;
  assign n35549 = ~n35089 & ~n35548;
  assign n35550 = ~n35059 & n35072;
  assign n35551 = n35059 & ~n35073;
  assign n35552 = n35059 & n35072;
  assign n35553 = ~n35072 & ~n35073;
  assign n35554 = ~n35059 & ~n35072;
  assign n35555 = ~n57840 & ~n57841;
  assign n35556 = ~n35073 & ~n35550;
  assign n35557 = ~n35549 & ~n57842;
  assign n35558 = ~n35073 & ~n35557;
  assign n35559 = ~n35043 & n35056;
  assign n35560 = n35043 & ~n35057;
  assign n35561 = n35043 & n35056;
  assign n35562 = ~n35056 & ~n35057;
  assign n35563 = ~n35043 & ~n35056;
  assign n35564 = ~n57843 & ~n57844;
  assign n35565 = ~n35057 & ~n35559;
  assign n35566 = ~n35558 & ~n57845;
  assign n35567 = ~n35057 & ~n35566;
  assign n35568 = ~n35027 & n35040;
  assign n35569 = n35027 & ~n35041;
  assign n35570 = n35027 & n35040;
  assign n35571 = ~n35040 & ~n35041;
  assign n35572 = ~n35027 & ~n35040;
  assign n35573 = ~n57846 & ~n57847;
  assign n35574 = ~n35041 & ~n35568;
  assign n35575 = ~n35567 & ~n57848;
  assign n35576 = ~n35041 & ~n35575;
  assign n35577 = ~n35011 & n35024;
  assign n35578 = n35011 & ~n35025;
  assign n35579 = n35011 & n35024;
  assign n35580 = ~n35024 & ~n35025;
  assign n35581 = ~n35011 & ~n35024;
  assign n35582 = ~n57849 & ~n57850;
  assign n35583 = ~n35025 & ~n35577;
  assign n35584 = ~n35576 & ~n57851;
  assign n35585 = ~n35025 & ~n35584;
  assign n35586 = ~n34995 & n35008;
  assign n35587 = n34995 & ~n35009;
  assign n35588 = n34995 & n35008;
  assign n35589 = ~n35008 & ~n35009;
  assign n35590 = ~n34995 & ~n35008;
  assign n35591 = ~n57852 & ~n57853;
  assign n35592 = ~n35009 & ~n35586;
  assign n35593 = ~n35585 & ~n57854;
  assign n35594 = ~n35009 & ~n35593;
  assign n35595 = ~n34979 & n34992;
  assign n35596 = n34979 & ~n34993;
  assign n35597 = n34979 & n34992;
  assign n35598 = ~n34992 & ~n34993;
  assign n35599 = ~n34979 & ~n34992;
  assign n35600 = ~n57855 & ~n57856;
  assign n35601 = ~n34993 & ~n35595;
  assign n35602 = ~n35594 & ~n57857;
  assign n35603 = ~n34993 & ~n35602;
  assign n35604 = ~n34963 & n34976;
  assign n35605 = n34963 & ~n34977;
  assign n35606 = n34963 & n34976;
  assign n35607 = ~n34976 & ~n34977;
  assign n35608 = ~n34963 & ~n34976;
  assign n35609 = ~n57858 & ~n57859;
  assign n35610 = ~n34977 & ~n35604;
  assign n35611 = ~n35603 & ~n57860;
  assign n35612 = ~n34977 & ~n35611;
  assign n35613 = ~n34947 & n34960;
  assign n35614 = ~n34961 & ~n35613;
  assign n35615 = ~n35612 & n35614;
  assign n35616 = ~n34961 & ~n35615;
  assign n35617 = n34875 & ~n34877;
  assign n35618 = n34877 & ~n34878;
  assign n35619 = ~n34875 & ~n34878;
  assign n35620 = ~n35618 & ~n35619;
  assign n35621 = ~n34878 & ~n35617;
  assign n35622 = ~n35616 & ~n57861;
  assign n35623 = n35616 & n57861;
  assign n35624 = n18846 & ~n56668;
  assign n35625 = n19541 & n26253;
  assign n35626 = n55247 & n26259;
  assign n35627 = n19509 & n26256;
  assign n35628 = ~n35626 & ~n35627;
  assign n35629 = ~n35625 & n35628;
  assign n35630 = ~n35624 & n35629;
  assign n35631 = pi11  & ~n35630;
  assign n35632 = pi11  & ~n35631;
  assign n35633 = pi11  & n35630;
  assign n35634 = ~n35630 & ~n35631;
  assign n35635 = ~pi11  & ~n35630;
  assign n35636 = ~n57862 & ~n57863;
  assign n35637 = ~n35623 & ~n35636;
  assign n35638 = ~n35622 & ~n35623;
  assign n35639 = ~n35636 & n35638;
  assign n35640 = ~n35622 & ~n35639;
  assign n35641 = ~n35622 & ~n35637;
  assign n35642 = ~n57754 & ~n57864;
  assign n35643 = n57754 & n57864;
  assign n35644 = n20085 & n27808;
  assign n35645 = n21269 & n26242;
  assign n35646 = n55472 & n26247;
  assign n35647 = n21237 & n26244;
  assign n35648 = ~n35646 & ~n35647;
  assign n35649 = ~n35645 & n35648;
  assign n35650 = ~n35644 & n35649;
  assign n35651 = pi8  & ~n35650;
  assign n35652 = pi8  & ~n35651;
  assign n35653 = pi8  & n35650;
  assign n35654 = ~n35650 & ~n35651;
  assign n35655 = ~pi8  & ~n35650;
  assign n35656 = ~n57865 & ~n57866;
  assign n35657 = ~n35643 & ~n35656;
  assign n35658 = ~n35642 & ~n35643;
  assign n35659 = ~n35656 & n35658;
  assign n35660 = ~n35642 & ~n35659;
  assign n35661 = ~n35642 & ~n35657;
  assign n35662 = ~n29200 & ~n57867;
  assign n35663 = n29200 & n57867;
  assign n35664 = n34915 & ~n34917;
  assign n35665 = n34917 & ~n34918;
  assign n35666 = ~n34915 & ~n34918;
  assign n35667 = ~n35665 & ~n35666;
  assign n35668 = ~n34918 & ~n35664;
  assign n35669 = ~n35663 & ~n57868;
  assign n35670 = ~n35662 & ~n35663;
  assign n35671 = ~n57868 & n35670;
  assign n35672 = ~n35662 & ~n35671;
  assign n35673 = ~n35662 & ~n35669;
  assign n35674 = n34940 & ~n57869;
  assign n35675 = n57868 & ~n35670;
  assign n35676 = ~n57868 & ~n35671;
  assign n35677 = n35670 & ~n35671;
  assign n35678 = ~n35676 & ~n35677;
  assign n35679 = ~n35671 & ~n35675;
  assign n35680 = n35656 & ~n35658;
  assign n35681 = n35658 & ~n35659;
  assign n35682 = ~n35656 & ~n35659;
  assign n35683 = ~n35681 & ~n35682;
  assign n35684 = ~n35659 & ~n35680;
  assign n35685 = n18846 & n27387;
  assign n35686 = n19541 & n26256;
  assign n35687 = n55247 & n26262;
  assign n35688 = n19509 & n26259;
  assign n35689 = ~n35687 & ~n35688;
  assign n35690 = ~n35686 & n35689;
  assign n35691 = ~n35685 & n35690;
  assign n35692 = pi11  & ~n35691;
  assign n35693 = ~n35691 & ~n35692;
  assign n35694 = ~pi11  & ~n35691;
  assign n35695 = pi11  & ~n35692;
  assign n35696 = pi11  & n35691;
  assign n35697 = ~n57872 & ~n57873;
  assign n35698 = n35612 & ~n35614;
  assign n35699 = ~n35615 & ~n35698;
  assign n35700 = ~n35697 & n35699;
  assign n35701 = n18846 & ~n56639;
  assign n35702 = n19541 & n26259;
  assign n35703 = n55247 & n26265;
  assign n35704 = n19509 & n26262;
  assign n35705 = ~n35703 & ~n35704;
  assign n35706 = ~n35702 & n35705;
  assign n35707 = ~n35701 & n35706;
  assign n35708 = pi11  & ~n35707;
  assign n35709 = ~n35707 & ~n35708;
  assign n35710 = ~pi11  & ~n35707;
  assign n35711 = pi11  & ~n35708;
  assign n35712 = pi11  & n35707;
  assign n35713 = ~n57874 & ~n57875;
  assign n35714 = n35603 & n57860;
  assign n35715 = ~n35603 & ~n35611;
  assign n35716 = ~n57860 & ~n35611;
  assign n35717 = ~n35715 & ~n35716;
  assign n35718 = ~n35611 & ~n35714;
  assign n35719 = ~n35713 & ~n57876;
  assign n35720 = n18846 & n27466;
  assign n35721 = n19541 & n26262;
  assign n35722 = n55247 & n26268;
  assign n35723 = n19509 & n26265;
  assign n35724 = ~n35722 & ~n35723;
  assign n35725 = ~n35721 & n35724;
  assign n35726 = ~n35720 & n35725;
  assign n35727 = pi11  & ~n35726;
  assign n35728 = ~n35726 & ~n35727;
  assign n35729 = ~pi11  & ~n35726;
  assign n35730 = pi11  & ~n35727;
  assign n35731 = pi11  & n35726;
  assign n35732 = ~n57877 & ~n57878;
  assign n35733 = n35594 & n57857;
  assign n35734 = ~n35594 & ~n35602;
  assign n35735 = ~n57857 & ~n35602;
  assign n35736 = ~n35734 & ~n35735;
  assign n35737 = ~n35602 & ~n35733;
  assign n35738 = ~n35732 & ~n57879;
  assign n35739 = n18846 & n27042;
  assign n35740 = n19541 & n26265;
  assign n35741 = n55247 & n26271;
  assign n35742 = n19509 & n26268;
  assign n35743 = ~n35741 & ~n35742;
  assign n35744 = ~n35740 & n35743;
  assign n35745 = ~n35739 & n35744;
  assign n35746 = pi11  & ~n35745;
  assign n35747 = ~n35745 & ~n35746;
  assign n35748 = ~pi11  & ~n35745;
  assign n35749 = pi11  & ~n35746;
  assign n35750 = pi11  & n35745;
  assign n35751 = ~n57880 & ~n57881;
  assign n35752 = n35585 & n57854;
  assign n35753 = ~n35585 & ~n35593;
  assign n35754 = ~n57854 & ~n35593;
  assign n35755 = ~n35753 & ~n35754;
  assign n35756 = ~n35593 & ~n35752;
  assign n35757 = ~n35751 & ~n57882;
  assign n35758 = n18846 & ~n56601;
  assign n35759 = n19541 & n26268;
  assign n35760 = n55247 & n26274;
  assign n35761 = n19509 & n26271;
  assign n35762 = ~n35760 & ~n35761;
  assign n35763 = ~n35759 & n35762;
  assign n35764 = ~n35758 & n35763;
  assign n35765 = pi11  & ~n35764;
  assign n35766 = ~n35764 & ~n35765;
  assign n35767 = ~pi11  & ~n35764;
  assign n35768 = pi11  & ~n35765;
  assign n35769 = pi11  & n35764;
  assign n35770 = ~n57883 & ~n57884;
  assign n35771 = n35576 & n57851;
  assign n35772 = ~n35576 & ~n35584;
  assign n35773 = ~n57851 & ~n35584;
  assign n35774 = ~n35772 & ~n35773;
  assign n35775 = ~n35584 & ~n35771;
  assign n35776 = ~n35770 & ~n57885;
  assign n35777 = n18846 & ~n56612;
  assign n35778 = n19541 & n26271;
  assign n35779 = n55247 & n26277;
  assign n35780 = n19509 & n26274;
  assign n35781 = ~n35779 & ~n35780;
  assign n35782 = ~n35778 & n35781;
  assign n35783 = ~n35777 & n35782;
  assign n35784 = pi11  & ~n35783;
  assign n35785 = ~n35783 & ~n35784;
  assign n35786 = ~pi11  & ~n35783;
  assign n35787 = pi11  & ~n35784;
  assign n35788 = pi11  & n35783;
  assign n35789 = ~n57886 & ~n57887;
  assign n35790 = n35567 & n57848;
  assign n35791 = ~n35567 & ~n35575;
  assign n35792 = ~n35567 & n57848;
  assign n35793 = ~n57848 & ~n35575;
  assign n35794 = n35567 & ~n57848;
  assign n35795 = ~n57888 & ~n57889;
  assign n35796 = ~n35575 & ~n35790;
  assign n35797 = ~n35789 & ~n57890;
  assign n35798 = n18846 & ~n56648;
  assign n35799 = n19541 & n26274;
  assign n35800 = n55247 & n26280;
  assign n35801 = n19509 & n26277;
  assign n35802 = ~n35800 & ~n35801;
  assign n35803 = ~n35799 & n35802;
  assign n35804 = ~n35798 & n35803;
  assign n35805 = pi11  & ~n35804;
  assign n35806 = ~n35804 & ~n35805;
  assign n35807 = ~pi11  & ~n35804;
  assign n35808 = pi11  & ~n35805;
  assign n35809 = pi11  & n35804;
  assign n35810 = ~n57891 & ~n57892;
  assign n35811 = n35558 & n57845;
  assign n35812 = ~n35558 & ~n35566;
  assign n35813 = ~n35558 & n57845;
  assign n35814 = ~n57845 & ~n35566;
  assign n35815 = n35558 & ~n57845;
  assign n35816 = ~n57893 & ~n57894;
  assign n35817 = ~n35566 & ~n35811;
  assign n35818 = ~n35810 & ~n57895;
  assign n35819 = n18846 & n27330;
  assign n35820 = n19541 & n26277;
  assign n35821 = n55247 & n26283;
  assign n35822 = n19509 & n26280;
  assign n35823 = ~n35821 & ~n35822;
  assign n35824 = ~n35820 & n35823;
  assign n35825 = ~n35819 & n35824;
  assign n35826 = pi11  & ~n35825;
  assign n35827 = ~n35825 & ~n35826;
  assign n35828 = ~pi11  & ~n35825;
  assign n35829 = pi11  & ~n35826;
  assign n35830 = pi11  & n35825;
  assign n35831 = ~n57896 & ~n57897;
  assign n35832 = n35549 & n57842;
  assign n35833 = ~n35549 & ~n35557;
  assign n35834 = ~n35549 & n57842;
  assign n35835 = ~n57842 & ~n35557;
  assign n35836 = n35549 & ~n57842;
  assign n35837 = ~n57898 & ~n57899;
  assign n35838 = ~n35557 & ~n35832;
  assign n35839 = ~n35831 & ~n57900;
  assign n35840 = n18846 & n27743;
  assign n35841 = n19541 & n26280;
  assign n35842 = n55247 & n26286;
  assign n35843 = n19509 & n26283;
  assign n35844 = ~n35842 & ~n35843;
  assign n35845 = ~n35841 & n35844;
  assign n35846 = ~n35840 & n35845;
  assign n35847 = pi11  & ~n35846;
  assign n35848 = ~n35846 & ~n35847;
  assign n35849 = ~pi11  & ~n35846;
  assign n35850 = pi11  & ~n35847;
  assign n35851 = pi11  & n35846;
  assign n35852 = ~n57901 & ~n57902;
  assign n35853 = n35540 & n57839;
  assign n35854 = ~n35540 & ~n35548;
  assign n35855 = ~n57839 & ~n35548;
  assign n35856 = ~n35854 & ~n35855;
  assign n35857 = ~n35548 & ~n35853;
  assign n35858 = ~n35852 & ~n57903;
  assign n35859 = n18846 & ~n56686;
  assign n35860 = n19541 & n26283;
  assign n35861 = n55247 & n26289;
  assign n35862 = n19509 & n26286;
  assign n35863 = ~n35861 & ~n35862;
  assign n35864 = ~n35860 & n35863;
  assign n35865 = ~n35859 & n35864;
  assign n35866 = pi11  & ~n35865;
  assign n35867 = ~n35865 & ~n35866;
  assign n35868 = ~pi11  & ~n35865;
  assign n35869 = pi11  & ~n35866;
  assign n35870 = pi11  & n35865;
  assign n35871 = ~n57904 & ~n57905;
  assign n35872 = n35531 & n57836;
  assign n35873 = ~n35531 & ~n35539;
  assign n35874 = ~n57836 & ~n35539;
  assign n35875 = ~n35873 & ~n35874;
  assign n35876 = ~n35539 & ~n35872;
  assign n35877 = ~n35871 & ~n57906;
  assign n35878 = n35522 & n57833;
  assign n35879 = ~n35530 & ~n35878;
  assign n35880 = n18846 & ~n56721;
  assign n35881 = n19541 & n26286;
  assign n35882 = n55247 & n26292;
  assign n35883 = n19509 & n26289;
  assign n35884 = ~n35882 & ~n35883;
  assign n35885 = ~n35881 & n35884;
  assign n35886 = ~n18846 & n35885;
  assign n35887 = n56721 & n35885;
  assign n35888 = ~n35886 & ~n35887;
  assign n35889 = ~n35880 & n35885;
  assign n35890 = pi11  & ~n57907;
  assign n35891 = ~pi11  & n57907;
  assign n35892 = ~n35890 & ~n35891;
  assign n35893 = n35879 & ~n35892;
  assign n35894 = n35513 & n57830;
  assign n35895 = ~n35521 & ~n35894;
  assign n35896 = n18846 & n28107;
  assign n35897 = n19541 & n26289;
  assign n35898 = n55247 & n26295;
  assign n35899 = n19509 & n26292;
  assign n35900 = ~n35898 & ~n35899;
  assign n35901 = ~n35897 & n35900;
  assign n35902 = ~n18846 & n35901;
  assign n35903 = ~n28107 & n35901;
  assign n35904 = ~n35902 & ~n35903;
  assign n35905 = ~n35896 & n35901;
  assign n35906 = pi11  & ~n57908;
  assign n35907 = ~pi11  & n57908;
  assign n35908 = ~n35906 & ~n35907;
  assign n35909 = n35895 & ~n35908;
  assign n35910 = n18846 & n28808;
  assign n35911 = n19541 & n26292;
  assign n35912 = n55247 & n26298;
  assign n35913 = n19509 & n26295;
  assign n35914 = ~n35912 & ~n35913;
  assign n35915 = ~n35911 & n35914;
  assign n35916 = ~n35910 & n35915;
  assign n35917 = pi11  & ~n35916;
  assign n35918 = ~n35916 & ~n35917;
  assign n35919 = ~pi11  & ~n35916;
  assign n35920 = pi11  & ~n35917;
  assign n35921 = pi11  & n35916;
  assign n35922 = ~n57909 & ~n57910;
  assign n35923 = n35509 & ~n35511;
  assign n35924 = ~n35512 & ~n35923;
  assign n35925 = ~n35922 & n35924;
  assign n35926 = n18846 & n28493;
  assign n35927 = n19541 & n26295;
  assign n35928 = n55247 & n26301;
  assign n35929 = n19509 & n26298;
  assign n35930 = ~n35928 & ~n35929;
  assign n35931 = ~n35927 & n35930;
  assign n35932 = ~n35926 & n35931;
  assign n35933 = pi11  & ~n35932;
  assign n35934 = ~n35932 & ~n35933;
  assign n35935 = ~pi11  & ~n35932;
  assign n35936 = pi11  & ~n35933;
  assign n35937 = pi11  & n35932;
  assign n35938 = ~n57911 & ~n57912;
  assign n35939 = n35500 & n57827;
  assign n35940 = ~n35500 & ~n35508;
  assign n35941 = ~n35500 & n57827;
  assign n35942 = ~n57827 & ~n35508;
  assign n35943 = n35500 & ~n57827;
  assign n35944 = ~n57913 & ~n57914;
  assign n35945 = ~n35508 & ~n35939;
  assign n35946 = ~n35938 & ~n57915;
  assign n35947 = n18846 & ~n56870;
  assign n35948 = n19541 & n26298;
  assign n35949 = n55247 & n26304;
  assign n35950 = n19509 & n26301;
  assign n35951 = ~n35949 & ~n35950;
  assign n35952 = ~n35948 & n35951;
  assign n35953 = ~n35947 & n35952;
  assign n35954 = pi11  & ~n35953;
  assign n35955 = ~n35953 & ~n35954;
  assign n35956 = ~pi11  & ~n35953;
  assign n35957 = pi11  & ~n35954;
  assign n35958 = pi11  & n35953;
  assign n35959 = ~n57916 & ~n57917;
  assign n35960 = n35491 & n57824;
  assign n35961 = ~n35491 & ~n35499;
  assign n35962 = ~n57824 & ~n35499;
  assign n35963 = ~n35961 & ~n35962;
  assign n35964 = ~n35499 & ~n35960;
  assign n35965 = ~n35959 & ~n57918;
  assign n35966 = n35482 & n57821;
  assign n35967 = ~n35490 & ~n35966;
  assign n35968 = n18846 & n29446;
  assign n35969 = n19541 & n26301;
  assign n35970 = n55247 & n26307;
  assign n35971 = n19509 & n26304;
  assign n35972 = ~n35970 & ~n35971;
  assign n35973 = ~n35969 & n35972;
  assign n35974 = ~n18846 & n35973;
  assign n35975 = ~n29446 & n35973;
  assign n35976 = ~n35974 & ~n35975;
  assign n35977 = ~n35968 & n35973;
  assign n35978 = pi11  & ~n57919;
  assign n35979 = ~pi11  & n57919;
  assign n35980 = ~n35978 & ~n35979;
  assign n35981 = n35967 & ~n35980;
  assign n35982 = n35473 & n57818;
  assign n35983 = ~n35481 & ~n35982;
  assign n35984 = n18846 & ~n56867;
  assign n35985 = n19541 & n26304;
  assign n35986 = n55247 & n26310;
  assign n35987 = n19509 & n26307;
  assign n35988 = ~n35986 & ~n35987;
  assign n35989 = ~n35985 & n35988;
  assign n35990 = ~n18846 & n35989;
  assign n35991 = n56867 & n35989;
  assign n35992 = ~n35990 & ~n35991;
  assign n35993 = ~n35984 & n35989;
  assign n35994 = pi11  & ~n57920;
  assign n35995 = ~pi11  & n57920;
  assign n35996 = ~n35994 & ~n35995;
  assign n35997 = n35983 & ~n35996;
  assign n35998 = n35466 & n57815;
  assign n35999 = ~n35472 & ~n35998;
  assign n36000 = n18846 & ~n56928;
  assign n36001 = n19541 & n26307;
  assign n36002 = n55247 & n26313;
  assign n36003 = n19509 & n26310;
  assign n36004 = ~n36002 & ~n36003;
  assign n36005 = ~n36001 & n36004;
  assign n36006 = ~n18846 & n36005;
  assign n36007 = n56928 & n36005;
  assign n36008 = ~n36006 & ~n36007;
  assign n36009 = ~n36000 & n36005;
  assign n36010 = pi11  & ~n57921;
  assign n36011 = ~pi11  & n57921;
  assign n36012 = ~n36010 & ~n36011;
  assign n36013 = n35999 & ~n36012;
  assign n36014 = n18846 & ~n57002;
  assign n36015 = n19541 & n26310;
  assign n36016 = n55247 & n26316;
  assign n36017 = n19509 & n26313;
  assign n36018 = ~n36016 & ~n36017;
  assign n36019 = ~n36015 & n36018;
  assign n36020 = ~n36014 & n36019;
  assign n36021 = pi11  & ~n36020;
  assign n36022 = ~n36020 & ~n36021;
  assign n36023 = ~pi11  & ~n36020;
  assign n36024 = pi11  & ~n36021;
  assign n36025 = pi11  & n36020;
  assign n36026 = ~n57922 & ~n57923;
  assign n36027 = n35462 & ~n35464;
  assign n36028 = ~n35465 & ~n36027;
  assign n36029 = ~n36026 & n36028;
  assign n36030 = n18846 & n30192;
  assign n36031 = n19541 & n26313;
  assign n36032 = n55247 & n26319;
  assign n36033 = n19509 & n26316;
  assign n36034 = ~n36032 & ~n36033;
  assign n36035 = ~n36031 & n36034;
  assign n36036 = ~n36030 & n36035;
  assign n36037 = pi11  & ~n36036;
  assign n36038 = ~n36036 & ~n36037;
  assign n36039 = ~pi11  & ~n36036;
  assign n36040 = pi11  & ~n36037;
  assign n36041 = pi11  & n36036;
  assign n36042 = ~n57924 & ~n57925;
  assign n36043 = n35453 & n57814;
  assign n36044 = ~n35453 & ~n35461;
  assign n36045 = ~n57814 & ~n35461;
  assign n36046 = ~n36044 & ~n36045;
  assign n36047 = ~n35461 & ~n36043;
  assign n36048 = ~n36042 & ~n57926;
  assign n36049 = n18846 & ~n56920;
  assign n36050 = n19541 & n26316;
  assign n36051 = n55247 & n26322;
  assign n36052 = n19509 & n26319;
  assign n36053 = ~n36051 & ~n36052;
  assign n36054 = ~n36050 & n36053;
  assign n36055 = ~n36049 & n36054;
  assign n36056 = pi11  & ~n36055;
  assign n36057 = ~n36055 & ~n36056;
  assign n36058 = ~pi11  & ~n36055;
  assign n36059 = pi11  & ~n36056;
  assign n36060 = pi11  & n36055;
  assign n36061 = ~n57927 & ~n57928;
  assign n36062 = n35444 & n57811;
  assign n36063 = ~n35444 & ~n35452;
  assign n36064 = ~n35444 & n57811;
  assign n36065 = ~n57811 & ~n35452;
  assign n36066 = n35444 & ~n57811;
  assign n36067 = ~n57929 & ~n57930;
  assign n36068 = ~n35452 & ~n36062;
  assign n36069 = ~n36061 & ~n57931;
  assign n36070 = n35435 & n57808;
  assign n36071 = ~n35443 & ~n36070;
  assign n36072 = n18846 & n30264;
  assign n36073 = n19541 & n26319;
  assign n36074 = n55247 & n26325;
  assign n36075 = n19509 & n26322;
  assign n36076 = ~n36074 & ~n36075;
  assign n36077 = ~n36073 & n36076;
  assign n36078 = ~n18846 & n36077;
  assign n36079 = ~n30264 & n36077;
  assign n36080 = ~n36078 & ~n36079;
  assign n36081 = ~n36072 & n36077;
  assign n36082 = pi11  & ~n57932;
  assign n36083 = ~pi11  & n57932;
  assign n36084 = ~n36082 & ~n36083;
  assign n36085 = n36071 & ~n36084;
  assign n36086 = n35431 & ~n35433;
  assign n36087 = ~n35434 & ~n36086;
  assign n36088 = n18846 & ~n57012;
  assign n36089 = n19541 & n26322;
  assign n36090 = n55247 & n26328;
  assign n36091 = n19509 & n26325;
  assign n36092 = ~n36090 & ~n36091;
  assign n36093 = ~n36089 & n36092;
  assign n36094 = ~n18846 & n36093;
  assign n36095 = n57012 & n36093;
  assign n36096 = ~n36094 & ~n36095;
  assign n36097 = ~n36088 & n36093;
  assign n36098 = pi11  & ~n57933;
  assign n36099 = ~pi11  & n57933;
  assign n36100 = ~n36098 & ~n36099;
  assign n36101 = n36087 & ~n36100;
  assign n36102 = n35422 & n57805;
  assign n36103 = ~n35430 & ~n36102;
  assign n36104 = n18846 & ~n57017;
  assign n36105 = n19541 & n26325;
  assign n36106 = n55247 & n26331;
  assign n36107 = n19509 & n26328;
  assign n36108 = ~n36106 & ~n36107;
  assign n36109 = ~n36105 & n36108;
  assign n36110 = ~n18846 & n36109;
  assign n36111 = n57017 & n36109;
  assign n36112 = ~n36110 & ~n36111;
  assign n36113 = ~n36104 & n36109;
  assign n36114 = pi11  & ~n57934;
  assign n36115 = ~pi11  & n57934;
  assign n36116 = ~n36114 & ~n36115;
  assign n36117 = n36103 & ~n36116;
  assign n36118 = n18846 & n30470;
  assign n36119 = n19541 & n26328;
  assign n36120 = n55247 & n26334;
  assign n36121 = n19509 & n26331;
  assign n36122 = ~n36120 & ~n36121;
  assign n36123 = ~n36119 & n36122;
  assign n36124 = ~n36118 & n36123;
  assign n36125 = pi11  & ~n36124;
  assign n36126 = ~n36124 & ~n36125;
  assign n36127 = ~pi11  & ~n36124;
  assign n36128 = pi11  & ~n36125;
  assign n36129 = pi11  & n36124;
  assign n36130 = ~n57935 & ~n57936;
  assign n36131 = n35418 & ~n35420;
  assign n36132 = ~n35421 & ~n36131;
  assign n36133 = ~n36130 & n36132;
  assign n36134 = n18846 & ~n57033;
  assign n36135 = n19541 & n26331;
  assign n36136 = n55247 & n26337;
  assign n36137 = n19509 & n26334;
  assign n36138 = ~n36136 & ~n36137;
  assign n36139 = ~n36135 & n36138;
  assign n36140 = ~n18846 & n36139;
  assign n36141 = n57033 & n36139;
  assign n36142 = ~n36140 & ~n36141;
  assign n36143 = ~n36134 & n36139;
  assign n36144 = pi11  & ~n57937;
  assign n36145 = ~pi11  & n57937;
  assign n36146 = ~n36144 & ~n36145;
  assign n36147 = n35409 & n57802;
  assign n36148 = ~n57802 & ~n35417;
  assign n36149 = ~n35409 & ~n35417;
  assign n36150 = ~n36148 & ~n36149;
  assign n36151 = ~n35417 & ~n36147;
  assign n36152 = ~n36146 & ~n57938;
  assign n36153 = n18846 & ~n57042;
  assign n36154 = n19541 & n26334;
  assign n36155 = n55247 & n26340;
  assign n36156 = n19509 & n26337;
  assign n36157 = ~n36155 & ~n36156;
  assign n36158 = ~n36154 & n36157;
  assign n36159 = ~n36153 & n36158;
  assign n36160 = pi11  & ~n36159;
  assign n36161 = ~n36159 & ~n36160;
  assign n36162 = ~pi11  & ~n36159;
  assign n36163 = pi11  & ~n36160;
  assign n36164 = pi11  & n36159;
  assign n36165 = ~n57939 & ~n57940;
  assign n36166 = pi14  & ~n57795;
  assign n36167 = ~n57796 & ~n36166;
  assign n36168 = n57796 & n36166;
  assign n36169 = ~n57795 & n35393;
  assign n36170 = ~n57797 & ~n36169;
  assign n36171 = ~n36167 & ~n36168;
  assign n36172 = ~n36165 & n57941;
  assign n36173 = n18846 & n30866;
  assign n36174 = n19541 & n26337;
  assign n36175 = n55247 & n26343;
  assign n36176 = n19509 & n26340;
  assign n36177 = ~n36175 & ~n36176;
  assign n36178 = ~n36174 & n36177;
  assign n36179 = ~n18846 & n36178;
  assign n36180 = ~n30866 & n36178;
  assign n36181 = ~n36179 & ~n36180;
  assign n36182 = ~n36173 & n36178;
  assign n36183 = pi11  & ~n57942;
  assign n36184 = ~pi11  & n57942;
  assign n36185 = ~n36183 & ~n36184;
  assign n36186 = pi14  & n35373;
  assign n36187 = ~n35372 & n36186;
  assign n36188 = n35372 & ~n36186;
  assign n36189 = ~n35374 & n35378;
  assign n36190 = ~n57795 & ~n36189;
  assign n36191 = ~n36187 & ~n36188;
  assign n36192 = ~n36185 & n57943;
  assign n36193 = n18846 & ~n31019;
  assign n36194 = n19509 & ~n56543;
  assign n36195 = n19541 & n26348;
  assign n36196 = ~n36194 & ~n36195;
  assign n36197 = ~n36193 & n36196;
  assign n36198 = n55244 & ~n56543;
  assign n36199 = pi11  & ~n36198;
  assign n36200 = pi11  & ~n36197;
  assign n36201 = pi11  & ~n36200;
  assign n36202 = ~n36197 & ~n36200;
  assign n36203 = ~n36201 & ~n36202;
  assign n36204 = n36199 & ~n36203;
  assign n36205 = n36197 & n36199;
  assign n36206 = n18846 & ~n31140;
  assign n36207 = n19541 & n26343;
  assign n36208 = n55247 & ~n56543;
  assign n36209 = n19509 & n26348;
  assign n36210 = ~n36208 & ~n36209;
  assign n36211 = ~n36207 & n36210;
  assign n36212 = ~n18846 & n36211;
  assign n36213 = n31140 & n36211;
  assign n36214 = ~n36212 & ~n36213;
  assign n36215 = ~n36206 & n36211;
  assign n36216 = pi11  & ~n57945;
  assign n36217 = ~pi11  & n57945;
  assign n36218 = ~n36216 & ~n36217;
  assign n36219 = n57944 & ~n36218;
  assign n36220 = n57944 & ~n57945;
  assign n36221 = n35373 & n57946;
  assign n36222 = n18846 & n30915;
  assign n36223 = n19541 & n26340;
  assign n36224 = n55247 & n26348;
  assign n36225 = n19509 & n26343;
  assign n36226 = ~n36224 & ~n36225;
  assign n36227 = ~n36223 & n36226;
  assign n36228 = ~n36222 & n36227;
  assign n36229 = pi11  & ~n36228;
  assign n36230 = pi11  & ~n36229;
  assign n36231 = pi11  & n36228;
  assign n36232 = ~n36228 & ~n36229;
  assign n36233 = ~pi11  & ~n36228;
  assign n36234 = ~n57947 & ~n57948;
  assign n36235 = ~n35373 & ~n57946;
  assign n36236 = n57946 & ~n36221;
  assign n36237 = ~n35373 & n57946;
  assign n36238 = n35373 & ~n36221;
  assign n36239 = n35373 & ~n57946;
  assign n36240 = ~n57949 & ~n57950;
  assign n36241 = ~n36221 & ~n36235;
  assign n36242 = ~n36234 & ~n57951;
  assign n36243 = ~n36221 & ~n36242;
  assign n36244 = n36185 & ~n57943;
  assign n36245 = ~n36192 & ~n36244;
  assign n36246 = ~n36243 & n36245;
  assign n36247 = ~n36192 & ~n36246;
  assign n36248 = n36165 & ~n57941;
  assign n36249 = ~n36165 & ~n36172;
  assign n36250 = ~n36165 & ~n57941;
  assign n36251 = n57941 & ~n36172;
  assign n36252 = n36165 & n57941;
  assign n36253 = ~n57952 & ~n57953;
  assign n36254 = ~n36172 & ~n36248;
  assign n36255 = ~n36247 & ~n57954;
  assign n36256 = ~n36172 & ~n36255;
  assign n36257 = n36146 & n57938;
  assign n36258 = ~n36152 & ~n36257;
  assign n36259 = ~n36256 & n36258;
  assign n36260 = ~n36152 & ~n36259;
  assign n36261 = n36130 & ~n36132;
  assign n36262 = ~n36130 & ~n36133;
  assign n36263 = ~n36130 & ~n36132;
  assign n36264 = n36132 & ~n36133;
  assign n36265 = n36130 & n36132;
  assign n36266 = ~n57955 & ~n57956;
  assign n36267 = ~n36133 & ~n36261;
  assign n36268 = ~n36260 & ~n57957;
  assign n36269 = ~n36133 & ~n36268;
  assign n36270 = ~n36103 & n36116;
  assign n36271 = n36103 & ~n36117;
  assign n36272 = n36103 & n36116;
  assign n36273 = ~n36116 & ~n36117;
  assign n36274 = ~n36103 & ~n36116;
  assign n36275 = ~n57958 & ~n57959;
  assign n36276 = ~n36117 & ~n36270;
  assign n36277 = ~n36269 & ~n57960;
  assign n36278 = ~n36117 & ~n36277;
  assign n36279 = ~n36087 & n36100;
  assign n36280 = n36087 & ~n36101;
  assign n36281 = n36087 & n36100;
  assign n36282 = ~n36100 & ~n36101;
  assign n36283 = ~n36087 & ~n36100;
  assign n36284 = ~n57961 & ~n57962;
  assign n36285 = ~n36101 & ~n36279;
  assign n36286 = ~n36278 & ~n57963;
  assign n36287 = ~n36101 & ~n36286;
  assign n36288 = ~n36071 & n36084;
  assign n36289 = ~n36085 & ~n36288;
  assign n36290 = ~n36287 & n36289;
  assign n36291 = ~n36085 & ~n36290;
  assign n36292 = n36061 & n57931;
  assign n36293 = ~n36061 & ~n36069;
  assign n36294 = ~n57931 & ~n36069;
  assign n36295 = ~n36293 & ~n36294;
  assign n36296 = ~n36069 & ~n36292;
  assign n36297 = ~n36291 & ~n57964;
  assign n36298 = ~n36069 & ~n36297;
  assign n36299 = n36042 & n57926;
  assign n36300 = ~n36042 & ~n36048;
  assign n36301 = ~n36042 & n57926;
  assign n36302 = ~n57926 & ~n36048;
  assign n36303 = n36042 & ~n57926;
  assign n36304 = ~n57965 & ~n57966;
  assign n36305 = ~n36048 & ~n36299;
  assign n36306 = ~n36298 & ~n57967;
  assign n36307 = ~n36048 & ~n36306;
  assign n36308 = n36026 & ~n36028;
  assign n36309 = ~n36026 & ~n36029;
  assign n36310 = ~n36026 & ~n36028;
  assign n36311 = n36028 & ~n36029;
  assign n36312 = n36026 & n36028;
  assign n36313 = ~n57968 & ~n57969;
  assign n36314 = ~n36029 & ~n36308;
  assign n36315 = ~n36307 & ~n57970;
  assign n36316 = ~n36029 & ~n36315;
  assign n36317 = ~n35999 & n36012;
  assign n36318 = n35999 & ~n36013;
  assign n36319 = n35999 & n36012;
  assign n36320 = ~n36012 & ~n36013;
  assign n36321 = ~n35999 & ~n36012;
  assign n36322 = ~n57971 & ~n57972;
  assign n36323 = ~n36013 & ~n36317;
  assign n36324 = ~n36316 & ~n57973;
  assign n36325 = ~n36013 & ~n36324;
  assign n36326 = ~n35983 & n35996;
  assign n36327 = n35983 & ~n35997;
  assign n36328 = n35983 & n35996;
  assign n36329 = ~n35996 & ~n35997;
  assign n36330 = ~n35983 & ~n35996;
  assign n36331 = ~n57974 & ~n57975;
  assign n36332 = ~n35997 & ~n36326;
  assign n36333 = ~n36325 & ~n57976;
  assign n36334 = ~n35997 & ~n36333;
  assign n36335 = ~n35967 & n35980;
  assign n36336 = ~n35981 & ~n36335;
  assign n36337 = ~n36334 & n36336;
  assign n36338 = ~n35981 & ~n36337;
  assign n36339 = n35959 & n57918;
  assign n36340 = ~n35959 & ~n35965;
  assign n36341 = ~n35959 & n57918;
  assign n36342 = ~n57918 & ~n35965;
  assign n36343 = n35959 & ~n57918;
  assign n36344 = ~n57977 & ~n57978;
  assign n36345 = ~n35965 & ~n36339;
  assign n36346 = ~n36338 & ~n57979;
  assign n36347 = ~n35965 & ~n36346;
  assign n36348 = n35938 & n57915;
  assign n36349 = ~n35938 & ~n35946;
  assign n36350 = ~n57915 & ~n35946;
  assign n36351 = ~n36349 & ~n36350;
  assign n36352 = ~n35946 & ~n36348;
  assign n36353 = ~n36347 & ~n57980;
  assign n36354 = ~n35946 & ~n36353;
  assign n36355 = n35922 & ~n35924;
  assign n36356 = ~n35922 & ~n35925;
  assign n36357 = ~n35922 & ~n35924;
  assign n36358 = n35924 & ~n35925;
  assign n36359 = n35922 & n35924;
  assign n36360 = ~n57981 & ~n57982;
  assign n36361 = ~n35925 & ~n36355;
  assign n36362 = ~n36354 & ~n57983;
  assign n36363 = ~n35925 & ~n36362;
  assign n36364 = ~n35895 & n35908;
  assign n36365 = n35895 & ~n35909;
  assign n36366 = n35895 & n35908;
  assign n36367 = ~n35908 & ~n35909;
  assign n36368 = ~n35895 & ~n35908;
  assign n36369 = ~n57984 & ~n57985;
  assign n36370 = ~n35909 & ~n36364;
  assign n36371 = ~n36363 & ~n57986;
  assign n36372 = ~n35909 & ~n36371;
  assign n36373 = ~n35879 & n35892;
  assign n36374 = ~n35893 & ~n36373;
  assign n36375 = ~n36372 & n36374;
  assign n36376 = ~n35893 & ~n36375;
  assign n36377 = n35871 & n57906;
  assign n36378 = ~n35871 & ~n35877;
  assign n36379 = ~n35871 & n57906;
  assign n36380 = ~n57906 & ~n35877;
  assign n36381 = n35871 & ~n57906;
  assign n36382 = ~n57987 & ~n57988;
  assign n36383 = ~n35877 & ~n36377;
  assign n36384 = ~n36376 & ~n57989;
  assign n36385 = ~n35877 & ~n36384;
  assign n36386 = n35852 & n57903;
  assign n36387 = ~n35852 & ~n35858;
  assign n36388 = ~n35852 & n57903;
  assign n36389 = ~n57903 & ~n35858;
  assign n36390 = n35852 & ~n57903;
  assign n36391 = ~n57990 & ~n57991;
  assign n36392 = ~n35858 & ~n36386;
  assign n36393 = ~n36385 & ~n57992;
  assign n36394 = ~n35858 & ~n36393;
  assign n36395 = n35831 & n57900;
  assign n36396 = ~n35831 & ~n35839;
  assign n36397 = ~n57900 & ~n35839;
  assign n36398 = ~n36396 & ~n36397;
  assign n36399 = ~n35839 & ~n36395;
  assign n36400 = ~n36394 & ~n57993;
  assign n36401 = ~n35839 & ~n36400;
  assign n36402 = n35810 & n57895;
  assign n36403 = ~n35810 & ~n35818;
  assign n36404 = ~n57895 & ~n35818;
  assign n36405 = ~n36403 & ~n36404;
  assign n36406 = ~n35818 & ~n36402;
  assign n36407 = ~n36401 & ~n57994;
  assign n36408 = ~n35818 & ~n36407;
  assign n36409 = n35789 & n57890;
  assign n36410 = ~n35789 & ~n35797;
  assign n36411 = ~n57890 & ~n35797;
  assign n36412 = ~n36410 & ~n36411;
  assign n36413 = ~n35797 & ~n36409;
  assign n36414 = ~n36408 & ~n57995;
  assign n36415 = ~n35797 & ~n36414;
  assign n36416 = n35770 & n57885;
  assign n36417 = ~n35770 & ~n35776;
  assign n36418 = ~n35770 & n57885;
  assign n36419 = ~n57885 & ~n35776;
  assign n36420 = n35770 & ~n57885;
  assign n36421 = ~n57996 & ~n57997;
  assign n36422 = ~n35776 & ~n36416;
  assign n36423 = ~n36415 & ~n57998;
  assign n36424 = ~n35776 & ~n36423;
  assign n36425 = n35751 & n57882;
  assign n36426 = ~n35751 & ~n35757;
  assign n36427 = ~n35751 & n57882;
  assign n36428 = ~n57882 & ~n35757;
  assign n36429 = n35751 & ~n57882;
  assign n36430 = ~n57999 & ~n58000;
  assign n36431 = ~n35757 & ~n36425;
  assign n36432 = ~n36424 & ~n58001;
  assign n36433 = ~n35757 & ~n36432;
  assign n36434 = n35732 & n57879;
  assign n36435 = ~n35732 & ~n35738;
  assign n36436 = ~n35732 & n57879;
  assign n36437 = ~n57879 & ~n35738;
  assign n36438 = n35732 & ~n57879;
  assign n36439 = ~n58002 & ~n58003;
  assign n36440 = ~n35738 & ~n36434;
  assign n36441 = ~n36433 & ~n58004;
  assign n36442 = ~n35738 & ~n36441;
  assign n36443 = n35713 & n57876;
  assign n36444 = ~n35713 & ~n35719;
  assign n36445 = ~n35713 & n57876;
  assign n36446 = ~n57876 & ~n35719;
  assign n36447 = n35713 & ~n57876;
  assign n36448 = ~n58005 & ~n58006;
  assign n36449 = ~n35719 & ~n36443;
  assign n36450 = ~n36442 & ~n58007;
  assign n36451 = ~n35719 & ~n36450;
  assign n36452 = n35697 & ~n35699;
  assign n36453 = ~n35697 & ~n35700;
  assign n36454 = ~n35697 & ~n35699;
  assign n36455 = n35699 & ~n35700;
  assign n36456 = n35697 & n35699;
  assign n36457 = ~n58008 & ~n58009;
  assign n36458 = ~n35700 & ~n36452;
  assign n36459 = ~n36451 & ~n58010;
  assign n36460 = ~n35700 & ~n36459;
  assign n36461 = n35638 & ~n35639;
  assign n36462 = n35636 & n35638;
  assign n36463 = ~n35636 & ~n35639;
  assign n36464 = ~n35636 & ~n35638;
  assign n36465 = n35636 & ~n35638;
  assign n36466 = ~n35639 & ~n36465;
  assign n36467 = ~n58011 & ~n58012;
  assign n36468 = ~n36460 & n58013;
  assign n36469 = n36460 & ~n58013;
  assign n36470 = n20085 & n27839;
  assign n36471 = n21269 & n26244;
  assign n36472 = n55472 & n26250;
  assign n36473 = n21237 & n26247;
  assign n36474 = ~n36472 & ~n36473;
  assign n36475 = ~n36471 & n36474;
  assign n36476 = ~n36470 & n36475;
  assign n36477 = pi8  & ~n36476;
  assign n36478 = pi8  & ~n36477;
  assign n36479 = pi8  & n36476;
  assign n36480 = ~n36476 & ~n36477;
  assign n36481 = ~pi8  & ~n36476;
  assign n36482 = ~n58014 & ~n58015;
  assign n36483 = ~n36469 & ~n36482;
  assign n36484 = ~n36468 & ~n36469;
  assign n36485 = ~n36482 & n36484;
  assign n36486 = ~n36468 & ~n36485;
  assign n36487 = ~n36468 & ~n36483;
  assign n36488 = ~n57871 & ~n58016;
  assign n36489 = n57871 & n58016;
  assign n36490 = n21969 & ~n26537;
  assign n36491 = ~n23459 & ~n36490;
  assign n36492 = ~n24302 & n36491;
  assign n36493 = ~n24302 & ~n36490;
  assign n36494 = ~n23459 & n36493;
  assign n36495 = n29191 & ~n36490;
  assign n36496 = ~n77 & n58017;
  assign n36497 = pi5  & ~n36496;
  assign n36498 = pi5  & ~n36497;
  assign n36499 = pi5  & n36496;
  assign n36500 = ~n36496 & ~n36497;
  assign n36501 = ~pi5  & ~n36496;
  assign n36502 = ~n58018 & ~n58019;
  assign n36503 = ~n36489 & ~n36502;
  assign n36504 = ~n36488 & ~n36489;
  assign n36505 = ~n36502 & n36504;
  assign n36506 = ~n36488 & ~n36505;
  assign n36507 = ~n36488 & ~n36503;
  assign n36508 = ~n57870 & ~n58020;
  assign n36509 = n57870 & n58020;
  assign n36510 = ~n36508 & ~n36509;
  assign n36511 = n36502 & ~n36504;
  assign n36512 = n36504 & ~n36505;
  assign n36513 = ~n36502 & ~n36505;
  assign n36514 = ~n36512 & ~n36513;
  assign n36515 = ~n36505 & ~n36511;
  assign n36516 = n36451 & n58010;
  assign n36517 = ~n36459 & ~n36516;
  assign n36518 = n20085 & ~n56567;
  assign n36519 = n21269 & n26247;
  assign n36520 = n55472 & n26253;
  assign n36521 = n21237 & n26250;
  assign n36522 = ~n36520 & ~n36521;
  assign n36523 = ~n36519 & n36522;
  assign n36524 = ~n20085 & n36523;
  assign n36525 = n56567 & n36523;
  assign n36526 = ~n36524 & ~n36525;
  assign n36527 = ~n36518 & n36523;
  assign n36528 = pi8  & ~n58022;
  assign n36529 = ~pi8  & n58022;
  assign n36530 = ~n36528 & ~n36529;
  assign n36531 = n36517 & ~n36530;
  assign n36532 = n36442 & n58007;
  assign n36533 = ~n36450 & ~n36532;
  assign n36534 = n20085 & n27491;
  assign n36535 = n21269 & n26250;
  assign n36536 = n55472 & n26256;
  assign n36537 = n21237 & n26253;
  assign n36538 = ~n36536 & ~n36537;
  assign n36539 = ~n36535 & n36538;
  assign n36540 = ~n20085 & n36539;
  assign n36541 = ~n27491 & n36539;
  assign n36542 = ~n36540 & ~n36541;
  assign n36543 = ~n36534 & n36539;
  assign n36544 = pi8  & ~n58023;
  assign n36545 = ~pi8  & n58023;
  assign n36546 = ~n36544 & ~n36545;
  assign n36547 = n36533 & ~n36546;
  assign n36548 = n36433 & n58004;
  assign n36549 = ~n36441 & ~n36548;
  assign n36550 = n20085 & ~n56668;
  assign n36551 = n21269 & n26253;
  assign n36552 = n55472 & n26259;
  assign n36553 = n21237 & n26256;
  assign n36554 = ~n36552 & ~n36553;
  assign n36555 = ~n36551 & n36554;
  assign n36556 = ~n20085 & n36555;
  assign n36557 = n56668 & n36555;
  assign n36558 = ~n36556 & ~n36557;
  assign n36559 = ~n36550 & n36555;
  assign n36560 = pi8  & ~n58024;
  assign n36561 = ~pi8  & n58024;
  assign n36562 = ~n36560 & ~n36561;
  assign n36563 = n36549 & ~n36562;
  assign n36564 = n36424 & n58001;
  assign n36565 = ~n36432 & ~n36564;
  assign n36566 = n20085 & n27387;
  assign n36567 = n21269 & n26256;
  assign n36568 = n55472 & n26262;
  assign n36569 = n21237 & n26259;
  assign n36570 = ~n36568 & ~n36569;
  assign n36571 = ~n36567 & n36570;
  assign n36572 = ~n20085 & n36571;
  assign n36573 = ~n27387 & n36571;
  assign n36574 = ~n36572 & ~n36573;
  assign n36575 = ~n36566 & n36571;
  assign n36576 = pi8  & ~n58025;
  assign n36577 = ~pi8  & n58025;
  assign n36578 = ~n36576 & ~n36577;
  assign n36579 = n36565 & ~n36578;
  assign n36580 = n36415 & n57998;
  assign n36581 = ~n36423 & ~n36580;
  assign n36582 = n20085 & ~n56639;
  assign n36583 = n21269 & n26259;
  assign n36584 = n55472 & n26265;
  assign n36585 = n21237 & n26262;
  assign n36586 = ~n36584 & ~n36585;
  assign n36587 = ~n36583 & n36586;
  assign n36588 = ~n20085 & n36587;
  assign n36589 = n56639 & n36587;
  assign n36590 = ~n36588 & ~n36589;
  assign n36591 = ~n36582 & n36587;
  assign n36592 = pi8  & ~n58026;
  assign n36593 = ~pi8  & n58026;
  assign n36594 = ~n36592 & ~n36593;
  assign n36595 = n36581 & ~n36594;
  assign n36596 = n36408 & n57995;
  assign n36597 = ~n36414 & ~n36596;
  assign n36598 = n20085 & n27466;
  assign n36599 = n21269 & n26262;
  assign n36600 = n55472 & n26268;
  assign n36601 = n21237 & n26265;
  assign n36602 = ~n36600 & ~n36601;
  assign n36603 = ~n36599 & n36602;
  assign n36604 = ~n20085 & n36603;
  assign n36605 = ~n27466 & n36603;
  assign n36606 = ~n36604 & ~n36605;
  assign n36607 = ~n36598 & n36603;
  assign n36608 = pi8  & ~n58027;
  assign n36609 = ~pi8  & n58027;
  assign n36610 = ~n36608 & ~n36609;
  assign n36611 = n36597 & ~n36610;
  assign n36612 = n36401 & n57994;
  assign n36613 = ~n36407 & ~n36612;
  assign n36614 = n20085 & n27042;
  assign n36615 = n21269 & n26265;
  assign n36616 = n55472 & n26271;
  assign n36617 = n21237 & n26268;
  assign n36618 = ~n36616 & ~n36617;
  assign n36619 = ~n36615 & n36618;
  assign n36620 = ~n20085 & n36619;
  assign n36621 = ~n27042 & n36619;
  assign n36622 = ~n36620 & ~n36621;
  assign n36623 = ~n36614 & n36619;
  assign n36624 = pi8  & ~n58028;
  assign n36625 = ~pi8  & n58028;
  assign n36626 = ~n36624 & ~n36625;
  assign n36627 = n36613 & ~n36626;
  assign n36628 = n36394 & n57993;
  assign n36629 = ~n36400 & ~n36628;
  assign n36630 = n20085 & ~n56601;
  assign n36631 = n21269 & n26268;
  assign n36632 = n55472 & n26274;
  assign n36633 = n21237 & n26271;
  assign n36634 = ~n36632 & ~n36633;
  assign n36635 = ~n36631 & n36634;
  assign n36636 = ~n20085 & n36635;
  assign n36637 = n56601 & n36635;
  assign n36638 = ~n36636 & ~n36637;
  assign n36639 = ~n36630 & n36635;
  assign n36640 = pi8  & ~n58029;
  assign n36641 = ~pi8  & n58029;
  assign n36642 = ~n36640 & ~n36641;
  assign n36643 = n36629 & ~n36642;
  assign n36644 = n36385 & n57992;
  assign n36645 = ~n36393 & ~n36644;
  assign n36646 = n20085 & ~n56612;
  assign n36647 = n21269 & n26271;
  assign n36648 = n55472 & n26277;
  assign n36649 = n21237 & n26274;
  assign n36650 = ~n36648 & ~n36649;
  assign n36651 = ~n36647 & n36650;
  assign n36652 = ~n20085 & n36651;
  assign n36653 = n56612 & n36651;
  assign n36654 = ~n36652 & ~n36653;
  assign n36655 = ~n36646 & n36651;
  assign n36656 = pi8  & ~n58030;
  assign n36657 = ~pi8  & n58030;
  assign n36658 = ~n36656 & ~n36657;
  assign n36659 = n36645 & ~n36658;
  assign n36660 = n36376 & n57989;
  assign n36661 = ~n36384 & ~n36660;
  assign n36662 = n20085 & ~n56648;
  assign n36663 = n21269 & n26274;
  assign n36664 = n55472 & n26280;
  assign n36665 = n21237 & n26277;
  assign n36666 = ~n36664 & ~n36665;
  assign n36667 = ~n36663 & n36666;
  assign n36668 = ~n20085 & n36667;
  assign n36669 = n56648 & n36667;
  assign n36670 = ~n36668 & ~n36669;
  assign n36671 = ~n36662 & n36667;
  assign n36672 = pi8  & ~n58031;
  assign n36673 = ~pi8  & n58031;
  assign n36674 = ~n36672 & ~n36673;
  assign n36675 = n36661 & ~n36674;
  assign n36676 = n20085 & n27330;
  assign n36677 = n21269 & n26277;
  assign n36678 = n55472 & n26283;
  assign n36679 = n21237 & n26280;
  assign n36680 = ~n36678 & ~n36679;
  assign n36681 = ~n36677 & n36680;
  assign n36682 = ~n36676 & n36681;
  assign n36683 = pi8  & ~n36682;
  assign n36684 = ~n36682 & ~n36683;
  assign n36685 = ~pi8  & ~n36682;
  assign n36686 = pi8  & ~n36683;
  assign n36687 = pi8  & n36682;
  assign n36688 = ~n58032 & ~n58033;
  assign n36689 = n36372 & ~n36374;
  assign n36690 = ~n36375 & ~n36689;
  assign n36691 = ~n36688 & n36690;
  assign n36692 = n20085 & n27743;
  assign n36693 = n21269 & n26280;
  assign n36694 = n55472 & n26286;
  assign n36695 = n21237 & n26283;
  assign n36696 = ~n36694 & ~n36695;
  assign n36697 = ~n36693 & n36696;
  assign n36698 = ~n36692 & n36697;
  assign n36699 = pi8  & ~n36698;
  assign n36700 = ~n36698 & ~n36699;
  assign n36701 = ~pi8  & ~n36698;
  assign n36702 = pi8  & ~n36699;
  assign n36703 = pi8  & n36698;
  assign n36704 = ~n58034 & ~n58035;
  assign n36705 = n36363 & n57986;
  assign n36706 = ~n36363 & ~n36371;
  assign n36707 = ~n36363 & n57986;
  assign n36708 = ~n57986 & ~n36371;
  assign n36709 = n36363 & ~n57986;
  assign n36710 = ~n58036 & ~n58037;
  assign n36711 = ~n36371 & ~n36705;
  assign n36712 = ~n36704 & ~n58038;
  assign n36713 = n36354 & n57983;
  assign n36714 = ~n36362 & ~n36713;
  assign n36715 = n20085 & ~n56686;
  assign n36716 = n21269 & n26283;
  assign n36717 = n55472 & n26289;
  assign n36718 = n21237 & n26286;
  assign n36719 = ~n36717 & ~n36718;
  assign n36720 = ~n36716 & n36719;
  assign n36721 = ~n20085 & n36720;
  assign n36722 = n56686 & n36720;
  assign n36723 = ~n36721 & ~n36722;
  assign n36724 = ~n36715 & n36720;
  assign n36725 = pi8  & ~n58039;
  assign n36726 = ~pi8  & n58039;
  assign n36727 = ~n36725 & ~n36726;
  assign n36728 = n36714 & ~n36727;
  assign n36729 = n36347 & n57980;
  assign n36730 = ~n36353 & ~n36729;
  assign n36731 = n20085 & ~n56721;
  assign n36732 = n21269 & n26286;
  assign n36733 = n55472 & n26292;
  assign n36734 = n21237 & n26289;
  assign n36735 = ~n36733 & ~n36734;
  assign n36736 = ~n36732 & n36735;
  assign n36737 = ~n20085 & n36736;
  assign n36738 = n56721 & n36736;
  assign n36739 = ~n36737 & ~n36738;
  assign n36740 = ~n36731 & n36736;
  assign n36741 = pi8  & ~n58040;
  assign n36742 = ~pi8  & n58040;
  assign n36743 = ~n36741 & ~n36742;
  assign n36744 = n36730 & ~n36743;
  assign n36745 = n36338 & n57979;
  assign n36746 = ~n36346 & ~n36745;
  assign n36747 = n20085 & n28107;
  assign n36748 = n21269 & n26289;
  assign n36749 = n55472 & n26295;
  assign n36750 = n21237 & n26292;
  assign n36751 = ~n36749 & ~n36750;
  assign n36752 = ~n36748 & n36751;
  assign n36753 = ~n20085 & n36752;
  assign n36754 = ~n28107 & n36752;
  assign n36755 = ~n36753 & ~n36754;
  assign n36756 = ~n36747 & n36752;
  assign n36757 = pi8  & ~n58041;
  assign n36758 = ~pi8  & n58041;
  assign n36759 = ~n36757 & ~n36758;
  assign n36760 = n36746 & ~n36759;
  assign n36761 = n20085 & n28808;
  assign n36762 = n21269 & n26292;
  assign n36763 = n55472 & n26298;
  assign n36764 = n21237 & n26295;
  assign n36765 = ~n36763 & ~n36764;
  assign n36766 = ~n36762 & n36765;
  assign n36767 = ~n36761 & n36766;
  assign n36768 = pi8  & ~n36767;
  assign n36769 = ~n36767 & ~n36768;
  assign n36770 = ~pi8  & ~n36767;
  assign n36771 = pi8  & ~n36768;
  assign n36772 = pi8  & n36767;
  assign n36773 = ~n58042 & ~n58043;
  assign n36774 = n36334 & ~n36336;
  assign n36775 = ~n36337 & ~n36774;
  assign n36776 = ~n36773 & n36775;
  assign n36777 = n20085 & n28493;
  assign n36778 = n21269 & n26295;
  assign n36779 = n55472 & n26301;
  assign n36780 = n21237 & n26298;
  assign n36781 = ~n36779 & ~n36780;
  assign n36782 = ~n36778 & n36781;
  assign n36783 = ~n36777 & n36782;
  assign n36784 = pi8  & ~n36783;
  assign n36785 = ~n36783 & ~n36784;
  assign n36786 = ~pi8  & ~n36783;
  assign n36787 = pi8  & ~n36784;
  assign n36788 = pi8  & n36783;
  assign n36789 = ~n58044 & ~n58045;
  assign n36790 = n36325 & n57976;
  assign n36791 = ~n36325 & ~n36333;
  assign n36792 = ~n36325 & n57976;
  assign n36793 = ~n57976 & ~n36333;
  assign n36794 = n36325 & ~n57976;
  assign n36795 = ~n58046 & ~n58047;
  assign n36796 = ~n36333 & ~n36790;
  assign n36797 = ~n36789 & ~n58048;
  assign n36798 = n20085 & ~n56870;
  assign n36799 = n21269 & n26298;
  assign n36800 = n55472 & n26304;
  assign n36801 = n21237 & n26301;
  assign n36802 = ~n36800 & ~n36801;
  assign n36803 = ~n36799 & n36802;
  assign n36804 = ~n36798 & n36803;
  assign n36805 = pi8  & ~n36804;
  assign n36806 = ~n36804 & ~n36805;
  assign n36807 = ~pi8  & ~n36804;
  assign n36808 = pi8  & ~n36805;
  assign n36809 = pi8  & n36804;
  assign n36810 = ~n58049 & ~n58050;
  assign n36811 = n36316 & n57973;
  assign n36812 = ~n36316 & ~n36324;
  assign n36813 = ~n57973 & ~n36324;
  assign n36814 = ~n36812 & ~n36813;
  assign n36815 = ~n36324 & ~n36811;
  assign n36816 = ~n36810 & ~n58051;
  assign n36817 = n36307 & n57970;
  assign n36818 = ~n36315 & ~n36817;
  assign n36819 = n20085 & n29446;
  assign n36820 = n21269 & n26301;
  assign n36821 = n55472 & n26307;
  assign n36822 = n21237 & n26304;
  assign n36823 = ~n36821 & ~n36822;
  assign n36824 = ~n36820 & n36823;
  assign n36825 = ~n20085 & n36824;
  assign n36826 = ~n29446 & n36824;
  assign n36827 = ~n36825 & ~n36826;
  assign n36828 = ~n36819 & n36824;
  assign n36829 = pi8  & ~n58052;
  assign n36830 = ~pi8  & n58052;
  assign n36831 = ~n36829 & ~n36830;
  assign n36832 = n36818 & ~n36831;
  assign n36833 = n36298 & n57967;
  assign n36834 = ~n36306 & ~n36833;
  assign n36835 = n20085 & ~n56867;
  assign n36836 = n21269 & n26304;
  assign n36837 = n55472 & n26310;
  assign n36838 = n21237 & n26307;
  assign n36839 = ~n36837 & ~n36838;
  assign n36840 = ~n36836 & n36839;
  assign n36841 = ~n20085 & n36840;
  assign n36842 = n56867 & n36840;
  assign n36843 = ~n36841 & ~n36842;
  assign n36844 = ~n36835 & n36840;
  assign n36845 = pi8  & ~n58053;
  assign n36846 = ~pi8  & n58053;
  assign n36847 = ~n36845 & ~n36846;
  assign n36848 = n36834 & ~n36847;
  assign n36849 = n36291 & n57964;
  assign n36850 = ~n36297 & ~n36849;
  assign n36851 = n20085 & ~n56928;
  assign n36852 = n21269 & n26307;
  assign n36853 = n55472 & n26313;
  assign n36854 = n21237 & n26310;
  assign n36855 = ~n36853 & ~n36854;
  assign n36856 = ~n36852 & n36855;
  assign n36857 = ~n20085 & n36856;
  assign n36858 = n56928 & n36856;
  assign n36859 = ~n36857 & ~n36858;
  assign n36860 = ~n36851 & n36856;
  assign n36861 = pi8  & ~n58054;
  assign n36862 = ~pi8  & n58054;
  assign n36863 = ~n36861 & ~n36862;
  assign n36864 = n36850 & ~n36863;
  assign n36865 = n20085 & ~n57002;
  assign n36866 = n21269 & n26310;
  assign n36867 = n55472 & n26316;
  assign n36868 = n21237 & n26313;
  assign n36869 = ~n36867 & ~n36868;
  assign n36870 = ~n36866 & n36869;
  assign n36871 = ~n36865 & n36870;
  assign n36872 = pi8  & ~n36871;
  assign n36873 = ~n36871 & ~n36872;
  assign n36874 = ~pi8  & ~n36871;
  assign n36875 = pi8  & ~n36872;
  assign n36876 = pi8  & n36871;
  assign n36877 = ~n58055 & ~n58056;
  assign n36878 = n36287 & ~n36289;
  assign n36879 = ~n36290 & ~n36878;
  assign n36880 = ~n36877 & n36879;
  assign n36881 = n20085 & n30192;
  assign n36882 = n21269 & n26313;
  assign n36883 = n55472 & n26319;
  assign n36884 = n21237 & n26316;
  assign n36885 = ~n36883 & ~n36884;
  assign n36886 = ~n36882 & n36885;
  assign n36887 = ~n36881 & n36886;
  assign n36888 = pi8  & ~n36887;
  assign n36889 = ~n36887 & ~n36888;
  assign n36890 = ~pi8  & ~n36887;
  assign n36891 = pi8  & ~n36888;
  assign n36892 = pi8  & n36887;
  assign n36893 = ~n58057 & ~n58058;
  assign n36894 = n36278 & n57963;
  assign n36895 = ~n36278 & ~n36286;
  assign n36896 = ~n57963 & ~n36286;
  assign n36897 = ~n36895 & ~n36896;
  assign n36898 = ~n36286 & ~n36894;
  assign n36899 = ~n36893 & ~n58059;
  assign n36900 = n20085 & ~n56920;
  assign n36901 = n21269 & n26316;
  assign n36902 = n55472 & n26322;
  assign n36903 = n21237 & n26319;
  assign n36904 = ~n36902 & ~n36903;
  assign n36905 = ~n36901 & n36904;
  assign n36906 = ~n36900 & n36905;
  assign n36907 = pi8  & ~n36906;
  assign n36908 = ~n36906 & ~n36907;
  assign n36909 = ~pi8  & ~n36906;
  assign n36910 = pi8  & ~n36907;
  assign n36911 = pi8  & n36906;
  assign n36912 = ~n58060 & ~n58061;
  assign n36913 = n36269 & n57960;
  assign n36914 = ~n36269 & ~n36277;
  assign n36915 = ~n36269 & n57960;
  assign n36916 = ~n57960 & ~n36277;
  assign n36917 = n36269 & ~n57960;
  assign n36918 = ~n58062 & ~n58063;
  assign n36919 = ~n36277 & ~n36913;
  assign n36920 = ~n36912 & ~n58064;
  assign n36921 = n36260 & n57957;
  assign n36922 = ~n36268 & ~n36921;
  assign n36923 = n20085 & n30264;
  assign n36924 = n21269 & n26319;
  assign n36925 = n55472 & n26325;
  assign n36926 = n21237 & n26322;
  assign n36927 = ~n36925 & ~n36926;
  assign n36928 = ~n36924 & n36927;
  assign n36929 = ~n20085 & n36928;
  assign n36930 = ~n30264 & n36928;
  assign n36931 = ~n36929 & ~n36930;
  assign n36932 = ~n36923 & n36928;
  assign n36933 = pi8  & ~n58065;
  assign n36934 = ~pi8  & n58065;
  assign n36935 = ~n36933 & ~n36934;
  assign n36936 = n36922 & ~n36935;
  assign n36937 = n36256 & ~n36258;
  assign n36938 = ~n36259 & ~n36937;
  assign n36939 = n20085 & ~n57012;
  assign n36940 = n21269 & n26322;
  assign n36941 = n55472 & n26328;
  assign n36942 = n21237 & n26325;
  assign n36943 = ~n36941 & ~n36942;
  assign n36944 = ~n36940 & n36943;
  assign n36945 = ~n20085 & n36944;
  assign n36946 = n57012 & n36944;
  assign n36947 = ~n36945 & ~n36946;
  assign n36948 = ~n36939 & n36944;
  assign n36949 = pi8  & ~n58066;
  assign n36950 = ~pi8  & n58066;
  assign n36951 = ~n36949 & ~n36950;
  assign n36952 = n36938 & ~n36951;
  assign n36953 = n36247 & n57954;
  assign n36954 = ~n36255 & ~n36953;
  assign n36955 = n20085 & ~n57017;
  assign n36956 = n21269 & n26325;
  assign n36957 = n55472 & n26331;
  assign n36958 = n21237 & n26328;
  assign n36959 = ~n36957 & ~n36958;
  assign n36960 = ~n36956 & n36959;
  assign n36961 = ~n20085 & n36960;
  assign n36962 = n57017 & n36960;
  assign n36963 = ~n36961 & ~n36962;
  assign n36964 = ~n36955 & n36960;
  assign n36965 = pi8  & ~n58067;
  assign n36966 = ~pi8  & n58067;
  assign n36967 = ~n36965 & ~n36966;
  assign n36968 = n36954 & ~n36967;
  assign n36969 = n20085 & n30470;
  assign n36970 = n21269 & n26328;
  assign n36971 = n55472 & n26334;
  assign n36972 = n21237 & n26331;
  assign n36973 = ~n36971 & ~n36972;
  assign n36974 = ~n36970 & n36973;
  assign n36975 = ~n36969 & n36974;
  assign n36976 = pi8  & ~n36975;
  assign n36977 = ~n36975 & ~n36976;
  assign n36978 = ~pi8  & ~n36975;
  assign n36979 = pi8  & ~n36976;
  assign n36980 = pi8  & n36975;
  assign n36981 = ~n58068 & ~n58069;
  assign n36982 = n36243 & ~n36245;
  assign n36983 = ~n36246 & ~n36982;
  assign n36984 = ~n36981 & n36983;
  assign n36985 = n20085 & ~n57033;
  assign n36986 = n21269 & n26331;
  assign n36987 = n55472 & n26337;
  assign n36988 = n21237 & n26334;
  assign n36989 = ~n36987 & ~n36988;
  assign n36990 = ~n36986 & n36989;
  assign n36991 = ~n20085 & n36990;
  assign n36992 = n57033 & n36990;
  assign n36993 = ~n36991 & ~n36992;
  assign n36994 = ~n36985 & n36990;
  assign n36995 = pi8  & ~n58070;
  assign n36996 = ~pi8  & n58070;
  assign n36997 = ~n36995 & ~n36996;
  assign n36998 = n36234 & n57951;
  assign n36999 = ~n57951 & ~n36242;
  assign n37000 = ~n36234 & ~n36242;
  assign n37001 = ~n36999 & ~n37000;
  assign n37002 = ~n36242 & ~n36998;
  assign n37003 = ~n36997 & ~n58071;
  assign n37004 = n20085 & ~n57042;
  assign n37005 = n21269 & n26334;
  assign n37006 = n55472 & n26340;
  assign n37007 = n21237 & n26337;
  assign n37008 = ~n37006 & ~n37007;
  assign n37009 = ~n37005 & n37008;
  assign n37010 = ~n37004 & n37009;
  assign n37011 = pi8  & ~n37010;
  assign n37012 = ~n37010 & ~n37011;
  assign n37013 = ~pi8  & ~n37010;
  assign n37014 = pi8  & ~n37011;
  assign n37015 = pi8  & n37010;
  assign n37016 = ~n58072 & ~n58073;
  assign n37017 = pi11  & ~n57944;
  assign n37018 = ~n57945 & ~n37017;
  assign n37019 = n57945 & n37017;
  assign n37020 = ~n57944 & n36218;
  assign n37021 = ~n57946 & ~n37020;
  assign n37022 = ~n37018 & ~n37019;
  assign n37023 = ~n37016 & n58074;
  assign n37024 = n20085 & n30866;
  assign n37025 = n21269 & n26337;
  assign n37026 = n55472 & n26343;
  assign n37027 = n21237 & n26340;
  assign n37028 = ~n37026 & ~n37027;
  assign n37029 = ~n37025 & n37028;
  assign n37030 = ~n20085 & n37029;
  assign n37031 = ~n30866 & n37029;
  assign n37032 = ~n37030 & ~n37031;
  assign n37033 = ~n37024 & n37029;
  assign n37034 = pi8  & ~n58075;
  assign n37035 = ~pi8  & n58075;
  assign n37036 = ~n37034 & ~n37035;
  assign n37037 = pi11  & n36198;
  assign n37038 = ~n36197 & n37037;
  assign n37039 = n36197 & ~n37037;
  assign n37040 = ~n36199 & n36203;
  assign n37041 = ~n57944 & ~n37040;
  assign n37042 = ~n37038 & ~n37039;
  assign n37043 = ~n37036 & n58076;
  assign n37044 = n20085 & ~n31019;
  assign n37045 = n21237 & ~n56543;
  assign n37046 = n21269 & n26348;
  assign n37047 = ~n37045 & ~n37046;
  assign n37048 = ~n37044 & n37047;
  assign n37049 = n55469 & ~n56543;
  assign n37050 = pi8  & ~n37049;
  assign n37051 = pi8  & ~n37048;
  assign n37052 = pi8  & ~n37051;
  assign n37053 = ~n37048 & ~n37051;
  assign n37054 = ~n37052 & ~n37053;
  assign n37055 = n37050 & ~n37054;
  assign n37056 = n37048 & n37050;
  assign n37057 = n20085 & ~n31140;
  assign n37058 = n21269 & n26343;
  assign n37059 = n55472 & ~n56543;
  assign n37060 = n21237 & n26348;
  assign n37061 = ~n37059 & ~n37060;
  assign n37062 = ~n37058 & n37061;
  assign n37063 = ~n20085 & n37062;
  assign n37064 = n31140 & n37062;
  assign n37065 = ~n37063 & ~n37064;
  assign n37066 = ~n37057 & n37062;
  assign n37067 = pi8  & ~n58078;
  assign n37068 = ~pi8  & n58078;
  assign n37069 = ~n37067 & ~n37068;
  assign n37070 = n58077 & ~n37069;
  assign n37071 = n58077 & ~n58078;
  assign n37072 = n36198 & n58079;
  assign n37073 = n20085 & n30915;
  assign n37074 = n21269 & n26340;
  assign n37075 = n55472 & n26348;
  assign n37076 = n21237 & n26343;
  assign n37077 = ~n37075 & ~n37076;
  assign n37078 = ~n37074 & n37077;
  assign n37079 = ~n37073 & n37078;
  assign n37080 = pi8  & ~n37079;
  assign n37081 = pi8  & ~n37080;
  assign n37082 = pi8  & n37079;
  assign n37083 = ~n37079 & ~n37080;
  assign n37084 = ~pi8  & ~n37079;
  assign n37085 = ~n58080 & ~n58081;
  assign n37086 = ~n36198 & ~n58079;
  assign n37087 = n58079 & ~n37072;
  assign n37088 = ~n36198 & n58079;
  assign n37089 = n36198 & ~n37072;
  assign n37090 = n36198 & ~n58079;
  assign n37091 = ~n58082 & ~n58083;
  assign n37092 = ~n37072 & ~n37086;
  assign n37093 = ~n37085 & ~n58084;
  assign n37094 = ~n37072 & ~n37093;
  assign n37095 = n37036 & ~n58076;
  assign n37096 = ~n37043 & ~n37095;
  assign n37097 = ~n37094 & n37096;
  assign n37098 = ~n37043 & ~n37097;
  assign n37099 = n37016 & ~n58074;
  assign n37100 = ~n37016 & ~n37023;
  assign n37101 = ~n37016 & ~n58074;
  assign n37102 = n58074 & ~n37023;
  assign n37103 = n37016 & n58074;
  assign n37104 = ~n58085 & ~n58086;
  assign n37105 = ~n37023 & ~n37099;
  assign n37106 = ~n37098 & ~n58087;
  assign n37107 = ~n37023 & ~n37106;
  assign n37108 = n36997 & n58071;
  assign n37109 = ~n37003 & ~n37108;
  assign n37110 = ~n37107 & n37109;
  assign n37111 = ~n37003 & ~n37110;
  assign n37112 = n36981 & ~n36983;
  assign n37113 = ~n36981 & ~n36984;
  assign n37114 = ~n36981 & ~n36983;
  assign n37115 = n36983 & ~n36984;
  assign n37116 = n36981 & n36983;
  assign n37117 = ~n58088 & ~n58089;
  assign n37118 = ~n36984 & ~n37112;
  assign n37119 = ~n37111 & ~n58090;
  assign n37120 = ~n36984 & ~n37119;
  assign n37121 = ~n36954 & n36967;
  assign n37122 = n36954 & ~n36968;
  assign n37123 = n36954 & n36967;
  assign n37124 = ~n36967 & ~n36968;
  assign n37125 = ~n36954 & ~n36967;
  assign n37126 = ~n58091 & ~n58092;
  assign n37127 = ~n36968 & ~n37121;
  assign n37128 = ~n37120 & ~n58093;
  assign n37129 = ~n36968 & ~n37128;
  assign n37130 = ~n36938 & n36951;
  assign n37131 = n36938 & ~n36952;
  assign n37132 = n36938 & n36951;
  assign n37133 = ~n36951 & ~n36952;
  assign n37134 = ~n36938 & ~n36951;
  assign n37135 = ~n58094 & ~n58095;
  assign n37136 = ~n36952 & ~n37130;
  assign n37137 = ~n37129 & ~n58096;
  assign n37138 = ~n36952 & ~n37137;
  assign n37139 = ~n36922 & n36935;
  assign n37140 = ~n36936 & ~n37139;
  assign n37141 = ~n37138 & n37140;
  assign n37142 = ~n36936 & ~n37141;
  assign n37143 = n36912 & n58064;
  assign n37144 = ~n36912 & ~n36920;
  assign n37145 = ~n58064 & ~n36920;
  assign n37146 = ~n37144 & ~n37145;
  assign n37147 = ~n36920 & ~n37143;
  assign n37148 = ~n37142 & ~n58097;
  assign n37149 = ~n36920 & ~n37148;
  assign n37150 = n36893 & n58059;
  assign n37151 = ~n36893 & ~n36899;
  assign n37152 = ~n36893 & n58059;
  assign n37153 = ~n58059 & ~n36899;
  assign n37154 = n36893 & ~n58059;
  assign n37155 = ~n58098 & ~n58099;
  assign n37156 = ~n36899 & ~n37150;
  assign n37157 = ~n37149 & ~n58100;
  assign n37158 = ~n36899 & ~n37157;
  assign n37159 = n36877 & ~n36879;
  assign n37160 = ~n36877 & ~n36880;
  assign n37161 = ~n36877 & ~n36879;
  assign n37162 = n36879 & ~n36880;
  assign n37163 = n36877 & n36879;
  assign n37164 = ~n58101 & ~n58102;
  assign n37165 = ~n36880 & ~n37159;
  assign n37166 = ~n37158 & ~n58103;
  assign n37167 = ~n36880 & ~n37166;
  assign n37168 = ~n36850 & n36863;
  assign n37169 = n36850 & ~n36864;
  assign n37170 = n36850 & n36863;
  assign n37171 = ~n36863 & ~n36864;
  assign n37172 = ~n36850 & ~n36863;
  assign n37173 = ~n58104 & ~n58105;
  assign n37174 = ~n36864 & ~n37168;
  assign n37175 = ~n37167 & ~n58106;
  assign n37176 = ~n36864 & ~n37175;
  assign n37177 = ~n36834 & n36847;
  assign n37178 = n36834 & ~n36848;
  assign n37179 = n36834 & n36847;
  assign n37180 = ~n36847 & ~n36848;
  assign n37181 = ~n36834 & ~n36847;
  assign n37182 = ~n58107 & ~n58108;
  assign n37183 = ~n36848 & ~n37177;
  assign n37184 = ~n37176 & ~n58109;
  assign n37185 = ~n36848 & ~n37184;
  assign n37186 = ~n36818 & n36831;
  assign n37187 = ~n36832 & ~n37186;
  assign n37188 = ~n37185 & n37187;
  assign n37189 = ~n36832 & ~n37188;
  assign n37190 = n36810 & n58051;
  assign n37191 = ~n36810 & ~n36816;
  assign n37192 = ~n36810 & n58051;
  assign n37193 = ~n58051 & ~n36816;
  assign n37194 = n36810 & ~n58051;
  assign n37195 = ~n58110 & ~n58111;
  assign n37196 = ~n36816 & ~n37190;
  assign n37197 = ~n37189 & ~n58112;
  assign n37198 = ~n36816 & ~n37197;
  assign n37199 = n36789 & n58048;
  assign n37200 = ~n36789 & ~n36797;
  assign n37201 = ~n58048 & ~n36797;
  assign n37202 = ~n37200 & ~n37201;
  assign n37203 = ~n36797 & ~n37199;
  assign n37204 = ~n37198 & ~n58113;
  assign n37205 = ~n36797 & ~n37204;
  assign n37206 = n36773 & ~n36775;
  assign n37207 = ~n36773 & ~n36776;
  assign n37208 = ~n36773 & ~n36775;
  assign n37209 = n36775 & ~n36776;
  assign n37210 = n36773 & n36775;
  assign n37211 = ~n58114 & ~n58115;
  assign n37212 = ~n36776 & ~n37206;
  assign n37213 = ~n37205 & ~n58116;
  assign n37214 = ~n36776 & ~n37213;
  assign n37215 = ~n36746 & n36759;
  assign n37216 = n36746 & ~n36760;
  assign n37217 = n36746 & n36759;
  assign n37218 = ~n36759 & ~n36760;
  assign n37219 = ~n36746 & ~n36759;
  assign n37220 = ~n58117 & ~n58118;
  assign n37221 = ~n36760 & ~n37215;
  assign n37222 = ~n37214 & ~n58119;
  assign n37223 = ~n36760 & ~n37222;
  assign n37224 = ~n36730 & n36743;
  assign n37225 = n36730 & ~n36744;
  assign n37226 = n36730 & n36743;
  assign n37227 = ~n36743 & ~n36744;
  assign n37228 = ~n36730 & ~n36743;
  assign n37229 = ~n58120 & ~n58121;
  assign n37230 = ~n36744 & ~n37224;
  assign n37231 = ~n37223 & ~n58122;
  assign n37232 = ~n36744 & ~n37231;
  assign n37233 = ~n36714 & n36727;
  assign n37234 = ~n36728 & ~n37233;
  assign n37235 = ~n37232 & n37234;
  assign n37236 = ~n36728 & ~n37235;
  assign n37237 = n36704 & n58038;
  assign n37238 = ~n36704 & ~n36712;
  assign n37239 = ~n58038 & ~n36712;
  assign n37240 = ~n37238 & ~n37239;
  assign n37241 = ~n36712 & ~n37237;
  assign n37242 = ~n37236 & ~n58123;
  assign n37243 = ~n36712 & ~n37242;
  assign n37244 = n36688 & ~n36690;
  assign n37245 = ~n36688 & ~n36691;
  assign n37246 = ~n36688 & ~n36690;
  assign n37247 = n36690 & ~n36691;
  assign n37248 = n36688 & n36690;
  assign n37249 = ~n58124 & ~n58125;
  assign n37250 = ~n36691 & ~n37244;
  assign n37251 = ~n37243 & ~n58126;
  assign n37252 = ~n36691 & ~n37251;
  assign n37253 = ~n36661 & n36674;
  assign n37254 = n36661 & ~n36675;
  assign n37255 = n36661 & n36674;
  assign n37256 = ~n36674 & ~n36675;
  assign n37257 = ~n36661 & ~n36674;
  assign n37258 = ~n58127 & ~n58128;
  assign n37259 = ~n36675 & ~n37253;
  assign n37260 = ~n37252 & ~n58129;
  assign n37261 = ~n36675 & ~n37260;
  assign n37262 = ~n36645 & n36658;
  assign n37263 = n36645 & ~n36659;
  assign n37264 = n36645 & n36658;
  assign n37265 = ~n36658 & ~n36659;
  assign n37266 = ~n36645 & ~n36658;
  assign n37267 = ~n58130 & ~n58131;
  assign n37268 = ~n36659 & ~n37262;
  assign n37269 = ~n37261 & ~n58132;
  assign n37270 = ~n36659 & ~n37269;
  assign n37271 = ~n36629 & n36642;
  assign n37272 = n36629 & ~n36643;
  assign n37273 = n36629 & n36642;
  assign n37274 = ~n36642 & ~n36643;
  assign n37275 = ~n36629 & ~n36642;
  assign n37276 = ~n58133 & ~n58134;
  assign n37277 = ~n36643 & ~n37271;
  assign n37278 = ~n37270 & ~n58135;
  assign n37279 = ~n36643 & ~n37278;
  assign n37280 = ~n36613 & n36626;
  assign n37281 = n36613 & ~n36627;
  assign n37282 = n36613 & n36626;
  assign n37283 = ~n36626 & ~n36627;
  assign n37284 = ~n36613 & ~n36626;
  assign n37285 = ~n58136 & ~n58137;
  assign n37286 = ~n36627 & ~n37280;
  assign n37287 = ~n37279 & ~n58138;
  assign n37288 = ~n36627 & ~n37287;
  assign n37289 = ~n36597 & n36610;
  assign n37290 = n36597 & ~n36611;
  assign n37291 = n36597 & n36610;
  assign n37292 = ~n36610 & ~n36611;
  assign n37293 = ~n36597 & ~n36610;
  assign n37294 = ~n58139 & ~n58140;
  assign n37295 = ~n36611 & ~n37289;
  assign n37296 = ~n37288 & ~n58141;
  assign n37297 = ~n36611 & ~n37296;
  assign n37298 = ~n36581 & n36594;
  assign n37299 = n36581 & ~n36595;
  assign n37300 = n36581 & n36594;
  assign n37301 = ~n36594 & ~n36595;
  assign n37302 = ~n36581 & ~n36594;
  assign n37303 = ~n58142 & ~n58143;
  assign n37304 = ~n36595 & ~n37298;
  assign n37305 = ~n37297 & ~n58144;
  assign n37306 = ~n36595 & ~n37305;
  assign n37307 = ~n36565 & n36578;
  assign n37308 = n36565 & ~n36579;
  assign n37309 = n36565 & n36578;
  assign n37310 = ~n36578 & ~n36579;
  assign n37311 = ~n36565 & ~n36578;
  assign n37312 = ~n58145 & ~n58146;
  assign n37313 = ~n36579 & ~n37307;
  assign n37314 = ~n37306 & ~n58147;
  assign n37315 = ~n36579 & ~n37314;
  assign n37316 = ~n36549 & n36562;
  assign n37317 = n36549 & ~n36563;
  assign n37318 = n36549 & n36562;
  assign n37319 = ~n36562 & ~n36563;
  assign n37320 = ~n36549 & ~n36562;
  assign n37321 = ~n58148 & ~n58149;
  assign n37322 = ~n36563 & ~n37316;
  assign n37323 = ~n37315 & ~n58150;
  assign n37324 = ~n36563 & ~n37323;
  assign n37325 = ~n36533 & n36546;
  assign n37326 = n36533 & ~n36547;
  assign n37327 = n36533 & n36546;
  assign n37328 = ~n36546 & ~n36547;
  assign n37329 = ~n36533 & ~n36546;
  assign n37330 = ~n58151 & ~n58152;
  assign n37331 = ~n36547 & ~n37325;
  assign n37332 = ~n37324 & ~n58153;
  assign n37333 = ~n36547 & ~n37332;
  assign n37334 = ~n36517 & n36530;
  assign n37335 = ~n36531 & ~n37334;
  assign n37336 = ~n37333 & n37335;
  assign n37337 = ~n36531 & ~n37336;
  assign n37338 = n36482 & ~n36484;
  assign n37339 = n36484 & ~n36485;
  assign n37340 = ~n36482 & ~n36485;
  assign n37341 = ~n37339 & ~n37340;
  assign n37342 = ~n36485 & ~n37338;
  assign n37343 = ~n37337 & ~n58154;
  assign n37344 = n37337 & n58154;
  assign n37345 = n77 & n28624;
  assign n37346 = n23459 & ~n26537;
  assign n37347 = n21969 & n26242;
  assign n37348 = ~n24302 & ~n37347;
  assign n37349 = ~n37346 & ~n37347;
  assign n37350 = ~n24302 & n37349;
  assign n37351 = ~n37346 & n37348;
  assign n37352 = ~n37345 & n58155;
  assign n37353 = pi5  & ~n37352;
  assign n37354 = pi5  & ~n37353;
  assign n37355 = pi5  & n37352;
  assign n37356 = ~n37352 & ~n37353;
  assign n37357 = ~pi5  & ~n37352;
  assign n37358 = ~n58156 & ~n58157;
  assign n37359 = ~n37344 & ~n37358;
  assign n37360 = ~n37343 & ~n37344;
  assign n37361 = ~n37358 & n37360;
  assign n37362 = ~n37343 & ~n37361;
  assign n37363 = ~n37343 & ~n37359;
  assign n37364 = ~n58021 & ~n58158;
  assign n37365 = n58021 & n58158;
  assign n37366 = ~n37364 & ~n37365;
  assign n37367 = n77 & ~n56564;
  assign n37368 = n24302 & ~n26537;
  assign n37369 = n21969 & n26244;
  assign n37370 = n23459 & n26242;
  assign n37371 = ~n37369 & ~n37370;
  assign n37372 = ~n37368 & n37371;
  assign n37373 = ~n37367 & n37372;
  assign n37374 = pi5  & ~n37373;
  assign n37375 = ~n37373 & ~n37374;
  assign n37376 = ~pi5  & ~n37373;
  assign n37377 = pi5  & ~n37374;
  assign n37378 = pi5  & n37373;
  assign n37379 = ~n58159 & ~n58160;
  assign n37380 = n37333 & ~n37335;
  assign n37381 = ~n37336 & ~n37380;
  assign n37382 = ~n37379 & n37381;
  assign n37383 = n37379 & ~n37381;
  assign n37384 = ~n37379 & ~n37382;
  assign n37385 = ~n37379 & ~n37381;
  assign n37386 = n37381 & ~n37382;
  assign n37387 = n37379 & n37381;
  assign n37388 = ~n58161 & ~n58162;
  assign n37389 = ~n37382 & ~n37383;
  assign n37390 = n56855 & ~n58163;
  assign n37391 = ~n37382 & ~n37390;
  assign n37392 = n37360 & ~n37361;
  assign n37393 = n37358 & n37360;
  assign n37394 = ~n37358 & ~n37361;
  assign n37395 = ~n37358 & ~n37360;
  assign n37396 = n37358 & ~n37360;
  assign n37397 = ~n37361 & ~n37396;
  assign n37398 = ~n58164 & ~n58165;
  assign n37399 = ~n37391 & n58166;
  assign n37400 = n37391 & ~n58166;
  assign n37401 = ~n37399 & ~n37400;
  assign n37402 = n77 & n27808;
  assign n37403 = n24302 & n26242;
  assign n37404 = n21969 & n26247;
  assign n37405 = n23459 & n26244;
  assign n37406 = ~n37404 & ~n37405;
  assign n37407 = ~n37403 & n37406;
  assign n37408 = ~n37402 & n37407;
  assign n37409 = pi5  & ~n37408;
  assign n37410 = ~n37408 & ~n37409;
  assign n37411 = ~pi5  & ~n37408;
  assign n37412 = pi5  & ~n37409;
  assign n37413 = pi5  & n37408;
  assign n37414 = ~n58167 & ~n58168;
  assign n37415 = n37324 & n58153;
  assign n37416 = ~n37324 & ~n37332;
  assign n37417 = ~n37324 & n58153;
  assign n37418 = ~n58153 & ~n37332;
  assign n37419 = n37324 & ~n58153;
  assign n37420 = ~n58169 & ~n58170;
  assign n37421 = ~n37332 & ~n37415;
  assign n37422 = ~n37414 & ~n58171;
  assign n37423 = n77 & n27839;
  assign n37424 = n24302 & n26244;
  assign n37425 = n21969 & n26250;
  assign n37426 = n23459 & n26247;
  assign n37427 = ~n37425 & ~n37426;
  assign n37428 = ~n37424 & n37427;
  assign n37429 = ~n37423 & n37428;
  assign n37430 = pi5  & ~n37429;
  assign n37431 = ~n37429 & ~n37430;
  assign n37432 = ~pi5  & ~n37429;
  assign n37433 = pi5  & ~n37430;
  assign n37434 = pi5  & n37429;
  assign n37435 = ~n58172 & ~n58173;
  assign n37436 = n37315 & n58150;
  assign n37437 = ~n37315 & ~n37323;
  assign n37438 = ~n37315 & n58150;
  assign n37439 = ~n58150 & ~n37323;
  assign n37440 = n37315 & ~n58150;
  assign n37441 = ~n58174 & ~n58175;
  assign n37442 = ~n37323 & ~n37436;
  assign n37443 = ~n37435 & ~n58176;
  assign n37444 = n77 & ~n56567;
  assign n37445 = n24302 & n26247;
  assign n37446 = n21969 & n26253;
  assign n37447 = n23459 & n26250;
  assign n37448 = ~n37446 & ~n37447;
  assign n37449 = ~n37445 & n37448;
  assign n37450 = ~n37444 & n37449;
  assign n37451 = pi5  & ~n37450;
  assign n37452 = ~n37450 & ~n37451;
  assign n37453 = ~pi5  & ~n37450;
  assign n37454 = pi5  & ~n37451;
  assign n37455 = pi5  & n37450;
  assign n37456 = ~n58177 & ~n58178;
  assign n37457 = n37306 & n58147;
  assign n37458 = ~n37306 & ~n37314;
  assign n37459 = ~n37306 & n58147;
  assign n37460 = ~n58147 & ~n37314;
  assign n37461 = n37306 & ~n58147;
  assign n37462 = ~n58179 & ~n58180;
  assign n37463 = ~n37314 & ~n37457;
  assign n37464 = ~n37456 & ~n58181;
  assign n37465 = n77 & n27491;
  assign n37466 = n24302 & n26250;
  assign n37467 = n21969 & n26256;
  assign n37468 = n23459 & n26253;
  assign n37469 = ~n37467 & ~n37468;
  assign n37470 = ~n37466 & n37469;
  assign n37471 = ~n37465 & n37470;
  assign n37472 = pi5  & ~n37471;
  assign n37473 = ~n37471 & ~n37472;
  assign n37474 = ~pi5  & ~n37471;
  assign n37475 = pi5  & ~n37472;
  assign n37476 = pi5  & n37471;
  assign n37477 = ~n58182 & ~n58183;
  assign n37478 = n37297 & n58144;
  assign n37479 = ~n37297 & ~n37305;
  assign n37480 = ~n37297 & n58144;
  assign n37481 = ~n58144 & ~n37305;
  assign n37482 = n37297 & ~n58144;
  assign n37483 = ~n58184 & ~n58185;
  assign n37484 = ~n37305 & ~n37478;
  assign n37485 = ~n37477 & ~n58186;
  assign n37486 = n77 & ~n56668;
  assign n37487 = n24302 & n26253;
  assign n37488 = n21969 & n26259;
  assign n37489 = n23459 & n26256;
  assign n37490 = ~n37488 & ~n37489;
  assign n37491 = ~n37487 & n37490;
  assign n37492 = ~n37486 & n37491;
  assign n37493 = pi5  & ~n37492;
  assign n37494 = ~n37492 & ~n37493;
  assign n37495 = ~pi5  & ~n37492;
  assign n37496 = pi5  & ~n37493;
  assign n37497 = pi5  & n37492;
  assign n37498 = ~n58187 & ~n58188;
  assign n37499 = n37288 & n58141;
  assign n37500 = ~n37288 & ~n37296;
  assign n37501 = ~n58141 & ~n37296;
  assign n37502 = ~n37500 & ~n37501;
  assign n37503 = ~n37296 & ~n37499;
  assign n37504 = ~n37498 & ~n58189;
  assign n37505 = n77 & n27387;
  assign n37506 = n24302 & n26256;
  assign n37507 = n21969 & n26262;
  assign n37508 = n23459 & n26259;
  assign n37509 = ~n37507 & ~n37508;
  assign n37510 = ~n37506 & n37509;
  assign n37511 = ~n37505 & n37510;
  assign n37512 = pi5  & ~n37511;
  assign n37513 = ~n37511 & ~n37512;
  assign n37514 = ~pi5  & ~n37511;
  assign n37515 = pi5  & ~n37512;
  assign n37516 = pi5  & n37511;
  assign n37517 = ~n58190 & ~n58191;
  assign n37518 = n37279 & n58138;
  assign n37519 = ~n37279 & ~n37287;
  assign n37520 = ~n58138 & ~n37287;
  assign n37521 = ~n37519 & ~n37520;
  assign n37522 = ~n37287 & ~n37518;
  assign n37523 = ~n37517 & ~n58192;
  assign n37524 = n77 & ~n56639;
  assign n37525 = n24302 & n26259;
  assign n37526 = n21969 & n26265;
  assign n37527 = n23459 & n26262;
  assign n37528 = ~n37526 & ~n37527;
  assign n37529 = ~n37525 & n37528;
  assign n37530 = ~n37524 & n37529;
  assign n37531 = pi5  & ~n37530;
  assign n37532 = ~n37530 & ~n37531;
  assign n37533 = ~pi5  & ~n37530;
  assign n37534 = pi5  & ~n37531;
  assign n37535 = pi5  & n37530;
  assign n37536 = ~n58193 & ~n58194;
  assign n37537 = n37270 & n58135;
  assign n37538 = ~n37270 & ~n37278;
  assign n37539 = ~n58135 & ~n37278;
  assign n37540 = ~n37538 & ~n37539;
  assign n37541 = ~n37278 & ~n37537;
  assign n37542 = ~n37536 & ~n58195;
  assign n37543 = n77 & n27466;
  assign n37544 = n24302 & n26262;
  assign n37545 = n21969 & n26268;
  assign n37546 = n23459 & n26265;
  assign n37547 = ~n37545 & ~n37546;
  assign n37548 = ~n37544 & n37547;
  assign n37549 = ~n37543 & n37548;
  assign n37550 = pi5  & ~n37549;
  assign n37551 = ~n37549 & ~n37550;
  assign n37552 = ~pi5  & ~n37549;
  assign n37553 = pi5  & ~n37550;
  assign n37554 = pi5  & n37549;
  assign n37555 = ~n58196 & ~n58197;
  assign n37556 = n37261 & n58132;
  assign n37557 = ~n37261 & ~n37269;
  assign n37558 = ~n37261 & n58132;
  assign n37559 = ~n58132 & ~n37269;
  assign n37560 = n37261 & ~n58132;
  assign n37561 = ~n58198 & ~n58199;
  assign n37562 = ~n37269 & ~n37556;
  assign n37563 = ~n37555 & ~n58200;
  assign n37564 = n77 & n27042;
  assign n37565 = n24302 & n26265;
  assign n37566 = n21969 & n26271;
  assign n37567 = n23459 & n26268;
  assign n37568 = ~n37566 & ~n37567;
  assign n37569 = ~n37565 & n37568;
  assign n37570 = ~n37564 & n37569;
  assign n37571 = pi5  & ~n37570;
  assign n37572 = ~n37570 & ~n37571;
  assign n37573 = ~pi5  & ~n37570;
  assign n37574 = pi5  & ~n37571;
  assign n37575 = pi5  & n37570;
  assign n37576 = ~n58201 & ~n58202;
  assign n37577 = n37252 & n58129;
  assign n37578 = ~n37252 & ~n37260;
  assign n37579 = ~n37252 & n58129;
  assign n37580 = ~n58129 & ~n37260;
  assign n37581 = n37252 & ~n58129;
  assign n37582 = ~n58203 & ~n58204;
  assign n37583 = ~n37260 & ~n37577;
  assign n37584 = ~n37576 & ~n58205;
  assign n37585 = n37243 & n58126;
  assign n37586 = ~n37251 & ~n37585;
  assign n37587 = n77 & ~n56601;
  assign n37588 = n24302 & n26268;
  assign n37589 = n21969 & n26274;
  assign n37590 = n23459 & n26271;
  assign n37591 = ~n37589 & ~n37590;
  assign n37592 = ~n37588 & n37591;
  assign n37593 = ~n77 & n37592;
  assign n37594 = n56601 & n37592;
  assign n37595 = ~n37593 & ~n37594;
  assign n37596 = ~n37587 & n37592;
  assign n37597 = pi5  & ~n58206;
  assign n37598 = ~pi5  & n58206;
  assign n37599 = ~n37597 & ~n37598;
  assign n37600 = n37586 & ~n37599;
  assign n37601 = n37236 & n58123;
  assign n37602 = ~n37242 & ~n37601;
  assign n37603 = n77 & ~n56612;
  assign n37604 = n24302 & n26271;
  assign n37605 = n21969 & n26277;
  assign n37606 = n23459 & n26274;
  assign n37607 = ~n37605 & ~n37606;
  assign n37608 = ~n37604 & n37607;
  assign n37609 = ~n77 & n37608;
  assign n37610 = n56612 & n37608;
  assign n37611 = ~n37609 & ~n37610;
  assign n37612 = ~n37603 & n37608;
  assign n37613 = pi5  & ~n58207;
  assign n37614 = ~pi5  & n58207;
  assign n37615 = ~n37613 & ~n37614;
  assign n37616 = n37602 & ~n37615;
  assign n37617 = n77 & ~n56648;
  assign n37618 = n24302 & n26274;
  assign n37619 = n21969 & n26280;
  assign n37620 = n23459 & n26277;
  assign n37621 = ~n37619 & ~n37620;
  assign n37622 = ~n37618 & n37621;
  assign n37623 = ~n37617 & n37622;
  assign n37624 = pi5  & ~n37623;
  assign n37625 = ~n37623 & ~n37624;
  assign n37626 = ~pi5  & ~n37623;
  assign n37627 = pi5  & ~n37624;
  assign n37628 = pi5  & n37623;
  assign n37629 = ~n58208 & ~n58209;
  assign n37630 = n37232 & ~n37234;
  assign n37631 = ~n37235 & ~n37630;
  assign n37632 = ~n37629 & n37631;
  assign n37633 = n77 & n27330;
  assign n37634 = n24302 & n26277;
  assign n37635 = n21969 & n26283;
  assign n37636 = n23459 & n26280;
  assign n37637 = ~n37635 & ~n37636;
  assign n37638 = ~n37634 & n37637;
  assign n37639 = ~n37633 & n37638;
  assign n37640 = pi5  & ~n37639;
  assign n37641 = ~n37639 & ~n37640;
  assign n37642 = ~pi5  & ~n37639;
  assign n37643 = pi5  & ~n37640;
  assign n37644 = pi5  & n37639;
  assign n37645 = ~n58210 & ~n58211;
  assign n37646 = n37223 & n58122;
  assign n37647 = ~n37223 & ~n37231;
  assign n37648 = ~n58122 & ~n37231;
  assign n37649 = ~n37647 & ~n37648;
  assign n37650 = ~n37231 & ~n37646;
  assign n37651 = ~n37645 & ~n58212;
  assign n37652 = n77 & n27743;
  assign n37653 = n24302 & n26280;
  assign n37654 = n21969 & n26286;
  assign n37655 = n23459 & n26283;
  assign n37656 = ~n37654 & ~n37655;
  assign n37657 = ~n37653 & n37656;
  assign n37658 = ~n37652 & n37657;
  assign n37659 = pi5  & ~n37658;
  assign n37660 = ~n37658 & ~n37659;
  assign n37661 = ~pi5  & ~n37658;
  assign n37662 = pi5  & ~n37659;
  assign n37663 = pi5  & n37658;
  assign n37664 = ~n58213 & ~n58214;
  assign n37665 = n37214 & n58119;
  assign n37666 = ~n37214 & ~n37222;
  assign n37667 = ~n37214 & n58119;
  assign n37668 = ~n58119 & ~n37222;
  assign n37669 = n37214 & ~n58119;
  assign n37670 = ~n58215 & ~n58216;
  assign n37671 = ~n37222 & ~n37665;
  assign n37672 = ~n37664 & ~n58217;
  assign n37673 = n37205 & n58116;
  assign n37674 = ~n37213 & ~n37673;
  assign n37675 = n77 & ~n56686;
  assign n37676 = n24302 & n26283;
  assign n37677 = n21969 & n26289;
  assign n37678 = n23459 & n26286;
  assign n37679 = ~n37677 & ~n37678;
  assign n37680 = ~n37676 & n37679;
  assign n37681 = ~n77 & n37680;
  assign n37682 = n56686 & n37680;
  assign n37683 = ~n37681 & ~n37682;
  assign n37684 = ~n37675 & n37680;
  assign n37685 = pi5  & ~n58218;
  assign n37686 = ~pi5  & n58218;
  assign n37687 = ~n37685 & ~n37686;
  assign n37688 = n37674 & ~n37687;
  assign n37689 = n37198 & n58113;
  assign n37690 = ~n37204 & ~n37689;
  assign n37691 = n77 & ~n56721;
  assign n37692 = n24302 & n26286;
  assign n37693 = n21969 & n26292;
  assign n37694 = n23459 & n26289;
  assign n37695 = ~n37693 & ~n37694;
  assign n37696 = ~n37692 & n37695;
  assign n37697 = ~n77 & n37696;
  assign n37698 = n56721 & n37696;
  assign n37699 = ~n37697 & ~n37698;
  assign n37700 = ~n37691 & n37696;
  assign n37701 = pi5  & ~n58219;
  assign n37702 = ~pi5  & n58219;
  assign n37703 = ~n37701 & ~n37702;
  assign n37704 = n37690 & ~n37703;
  assign n37705 = n37189 & n58112;
  assign n37706 = ~n37197 & ~n37705;
  assign n37707 = n77 & n28107;
  assign n37708 = n24302 & n26289;
  assign n37709 = n21969 & n26295;
  assign n37710 = n23459 & n26292;
  assign n37711 = ~n37709 & ~n37710;
  assign n37712 = ~n37708 & n37711;
  assign n37713 = ~n77 & n37712;
  assign n37714 = ~n28107 & n37712;
  assign n37715 = ~n37713 & ~n37714;
  assign n37716 = ~n37707 & n37712;
  assign n37717 = pi5  & ~n58220;
  assign n37718 = ~pi5  & n58220;
  assign n37719 = ~n37717 & ~n37718;
  assign n37720 = n37706 & ~n37719;
  assign n37721 = n77 & n28808;
  assign n37722 = n24302 & n26292;
  assign n37723 = n21969 & n26298;
  assign n37724 = n23459 & n26295;
  assign n37725 = ~n37723 & ~n37724;
  assign n37726 = ~n37722 & n37725;
  assign n37727 = ~n37721 & n37726;
  assign n37728 = pi5  & ~n37727;
  assign n37729 = ~n37727 & ~n37728;
  assign n37730 = ~pi5  & ~n37727;
  assign n37731 = pi5  & ~n37728;
  assign n37732 = pi5  & n37727;
  assign n37733 = ~n58221 & ~n58222;
  assign n37734 = n37185 & ~n37187;
  assign n37735 = ~n37188 & ~n37734;
  assign n37736 = ~n37733 & n37735;
  assign n37737 = n77 & n28493;
  assign n37738 = n24302 & n26295;
  assign n37739 = n21969 & n26301;
  assign n37740 = n23459 & n26298;
  assign n37741 = ~n37739 & ~n37740;
  assign n37742 = ~n37738 & n37741;
  assign n37743 = ~n37737 & n37742;
  assign n37744 = pi5  & ~n37743;
  assign n37745 = ~n37743 & ~n37744;
  assign n37746 = ~pi5  & ~n37743;
  assign n37747 = pi5  & ~n37744;
  assign n37748 = pi5  & n37743;
  assign n37749 = ~n58223 & ~n58224;
  assign n37750 = n37176 & n58109;
  assign n37751 = ~n37176 & ~n37184;
  assign n37752 = ~n37176 & n58109;
  assign n37753 = ~n58109 & ~n37184;
  assign n37754 = n37176 & ~n58109;
  assign n37755 = ~n58225 & ~n58226;
  assign n37756 = ~n37184 & ~n37750;
  assign n37757 = ~n37749 & ~n58227;
  assign n37758 = n77 & ~n56870;
  assign n37759 = n24302 & n26298;
  assign n37760 = n21969 & n26304;
  assign n37761 = n23459 & n26301;
  assign n37762 = ~n37760 & ~n37761;
  assign n37763 = ~n37759 & n37762;
  assign n37764 = ~n37758 & n37763;
  assign n37765 = pi5  & ~n37764;
  assign n37766 = ~n37764 & ~n37765;
  assign n37767 = ~pi5  & ~n37764;
  assign n37768 = pi5  & ~n37765;
  assign n37769 = pi5  & n37764;
  assign n37770 = ~n58228 & ~n58229;
  assign n37771 = n37167 & n58106;
  assign n37772 = ~n37167 & ~n37175;
  assign n37773 = ~n58106 & ~n37175;
  assign n37774 = ~n37772 & ~n37773;
  assign n37775 = ~n37175 & ~n37771;
  assign n37776 = ~n37770 & ~n58230;
  assign n37777 = n37158 & n58103;
  assign n37778 = ~n37166 & ~n37777;
  assign n37779 = n77 & n29446;
  assign n37780 = n24302 & n26301;
  assign n37781 = n21969 & n26307;
  assign n37782 = n23459 & n26304;
  assign n37783 = ~n37781 & ~n37782;
  assign n37784 = ~n37780 & n37783;
  assign n37785 = ~n77 & n37784;
  assign n37786 = ~n29446 & n37784;
  assign n37787 = ~n37785 & ~n37786;
  assign n37788 = ~n37779 & n37784;
  assign n37789 = pi5  & ~n58231;
  assign n37790 = ~pi5  & n58231;
  assign n37791 = ~n37789 & ~n37790;
  assign n37792 = n37778 & ~n37791;
  assign n37793 = n37149 & n58100;
  assign n37794 = ~n37157 & ~n37793;
  assign n37795 = n77 & ~n56867;
  assign n37796 = n24302 & n26304;
  assign n37797 = n21969 & n26310;
  assign n37798 = n23459 & n26307;
  assign n37799 = ~n37797 & ~n37798;
  assign n37800 = ~n37796 & n37799;
  assign n37801 = ~n77 & n37800;
  assign n37802 = n56867 & n37800;
  assign n37803 = ~n37801 & ~n37802;
  assign n37804 = ~n37795 & n37800;
  assign n37805 = pi5  & ~n58232;
  assign n37806 = ~pi5  & n58232;
  assign n37807 = ~n37805 & ~n37806;
  assign n37808 = n37794 & ~n37807;
  assign n37809 = n37142 & n58097;
  assign n37810 = ~n37148 & ~n37809;
  assign n37811 = n77 & ~n56928;
  assign n37812 = n24302 & n26307;
  assign n37813 = n21969 & n26313;
  assign n37814 = n23459 & n26310;
  assign n37815 = ~n37813 & ~n37814;
  assign n37816 = ~n37812 & n37815;
  assign n37817 = ~n77 & n37816;
  assign n37818 = n56928 & n37816;
  assign n37819 = ~n37817 & ~n37818;
  assign n37820 = ~n37811 & n37816;
  assign n37821 = pi5  & ~n58233;
  assign n37822 = ~pi5  & n58233;
  assign n37823 = ~n37821 & ~n37822;
  assign n37824 = n37810 & ~n37823;
  assign n37825 = n77 & ~n57002;
  assign n37826 = n24302 & n26310;
  assign n37827 = n21969 & n26316;
  assign n37828 = n23459 & n26313;
  assign n37829 = ~n37827 & ~n37828;
  assign n37830 = ~n37826 & n37829;
  assign n37831 = ~n37825 & n37830;
  assign n37832 = pi5  & ~n37831;
  assign n37833 = ~n37831 & ~n37832;
  assign n37834 = ~pi5  & ~n37831;
  assign n37835 = pi5  & ~n37832;
  assign n37836 = pi5  & n37831;
  assign n37837 = ~n58234 & ~n58235;
  assign n37838 = n37138 & ~n37140;
  assign n37839 = ~n37141 & ~n37838;
  assign n37840 = ~n37837 & n37839;
  assign n37841 = n77 & n30192;
  assign n37842 = n24302 & n26313;
  assign n37843 = n21969 & n26319;
  assign n37844 = n23459 & n26316;
  assign n37845 = ~n37843 & ~n37844;
  assign n37846 = ~n37842 & n37845;
  assign n37847 = ~n37841 & n37846;
  assign n37848 = pi5  & ~n37847;
  assign n37849 = ~n37847 & ~n37848;
  assign n37850 = ~pi5  & ~n37847;
  assign n37851 = pi5  & ~n37848;
  assign n37852 = pi5  & n37847;
  assign n37853 = ~n58236 & ~n58237;
  assign n37854 = n37129 & n58096;
  assign n37855 = ~n37129 & ~n37137;
  assign n37856 = ~n58096 & ~n37137;
  assign n37857 = ~n37855 & ~n37856;
  assign n37858 = ~n37137 & ~n37854;
  assign n37859 = ~n37853 & ~n58238;
  assign n37860 = n77 & ~n56920;
  assign n37861 = n24302 & n26316;
  assign n37862 = n21969 & n26322;
  assign n37863 = n23459 & n26319;
  assign n37864 = ~n37862 & ~n37863;
  assign n37865 = ~n37861 & n37864;
  assign n37866 = ~n37860 & n37865;
  assign n37867 = pi5  & ~n37866;
  assign n37868 = ~n37866 & ~n37867;
  assign n37869 = ~pi5  & ~n37866;
  assign n37870 = pi5  & ~n37867;
  assign n37871 = pi5  & n37866;
  assign n37872 = ~n58239 & ~n58240;
  assign n37873 = n37120 & n58093;
  assign n37874 = ~n37120 & ~n37128;
  assign n37875 = ~n37120 & n58093;
  assign n37876 = ~n58093 & ~n37128;
  assign n37877 = n37120 & ~n58093;
  assign n37878 = ~n58241 & ~n58242;
  assign n37879 = ~n37128 & ~n37873;
  assign n37880 = ~n37872 & ~n58243;
  assign n37881 = n37111 & n58090;
  assign n37882 = ~n37119 & ~n37881;
  assign n37883 = n77 & n30264;
  assign n37884 = n24302 & n26319;
  assign n37885 = n21969 & n26325;
  assign n37886 = n23459 & n26322;
  assign n37887 = ~n37885 & ~n37886;
  assign n37888 = ~n37884 & n37887;
  assign n37889 = ~n77 & n37888;
  assign n37890 = ~n30264 & n37888;
  assign n37891 = ~n37889 & ~n37890;
  assign n37892 = ~n37883 & n37888;
  assign n37893 = pi5  & ~n58244;
  assign n37894 = ~pi5  & n58244;
  assign n37895 = ~n37893 & ~n37894;
  assign n37896 = n37882 & ~n37895;
  assign n37897 = n37107 & ~n37109;
  assign n37898 = ~n37110 & ~n37897;
  assign n37899 = n77 & ~n57012;
  assign n37900 = n24302 & n26322;
  assign n37901 = n21969 & n26328;
  assign n37902 = n23459 & n26325;
  assign n37903 = ~n37901 & ~n37902;
  assign n37904 = ~n37900 & n37903;
  assign n37905 = ~n77 & n37904;
  assign n37906 = n57012 & n37904;
  assign n37907 = ~n37905 & ~n37906;
  assign n37908 = ~n37899 & n37904;
  assign n37909 = pi5  & ~n58245;
  assign n37910 = ~pi5  & n58245;
  assign n37911 = ~n37909 & ~n37910;
  assign n37912 = n37898 & ~n37911;
  assign n37913 = n37098 & n58087;
  assign n37914 = ~n37106 & ~n37913;
  assign n37915 = n77 & ~n57017;
  assign n37916 = n24302 & n26325;
  assign n37917 = n21969 & n26331;
  assign n37918 = n23459 & n26328;
  assign n37919 = ~n37917 & ~n37918;
  assign n37920 = ~n37916 & n37919;
  assign n37921 = ~n77 & n37920;
  assign n37922 = n57017 & n37920;
  assign n37923 = ~n37921 & ~n37922;
  assign n37924 = ~n37915 & n37920;
  assign n37925 = pi5  & ~n58246;
  assign n37926 = ~pi5  & n58246;
  assign n37927 = ~n37925 & ~n37926;
  assign n37928 = n37914 & ~n37927;
  assign n37929 = n77 & n30470;
  assign n37930 = n24302 & n26328;
  assign n37931 = n21969 & n26334;
  assign n37932 = n23459 & n26331;
  assign n37933 = ~n37931 & ~n37932;
  assign n37934 = ~n37930 & n37933;
  assign n37935 = ~n37929 & n37934;
  assign n37936 = pi5  & ~n37935;
  assign n37937 = ~n37935 & ~n37936;
  assign n37938 = ~pi5  & ~n37935;
  assign n37939 = pi5  & ~n37936;
  assign n37940 = pi5  & n37935;
  assign n37941 = ~n58247 & ~n58248;
  assign n37942 = n37094 & ~n37096;
  assign n37943 = ~n37097 & ~n37942;
  assign n37944 = ~n37941 & n37943;
  assign n37945 = n77 & ~n57033;
  assign n37946 = n24302 & n26331;
  assign n37947 = n21969 & n26337;
  assign n37948 = n23459 & n26334;
  assign n37949 = ~n37947 & ~n37948;
  assign n37950 = ~n37946 & n37949;
  assign n37951 = ~n77 & n37950;
  assign n37952 = n57033 & n37950;
  assign n37953 = ~n37951 & ~n37952;
  assign n37954 = ~n37945 & n37950;
  assign n37955 = pi5  & ~n58249;
  assign n37956 = ~pi5  & n58249;
  assign n37957 = ~n37955 & ~n37956;
  assign n37958 = n37085 & n58084;
  assign n37959 = ~n58084 & ~n37093;
  assign n37960 = ~n37085 & ~n37093;
  assign n37961 = ~n37959 & ~n37960;
  assign n37962 = ~n37093 & ~n37958;
  assign n37963 = ~n37957 & ~n58250;
  assign n37964 = n77 & ~n57042;
  assign n37965 = n24302 & n26334;
  assign n37966 = n21969 & n26340;
  assign n37967 = n23459 & n26337;
  assign n37968 = ~n37966 & ~n37967;
  assign n37969 = ~n37965 & n37968;
  assign n37970 = ~n37964 & n37969;
  assign n37971 = pi5  & ~n37970;
  assign n37972 = ~n37970 & ~n37971;
  assign n37973 = ~pi5  & ~n37970;
  assign n37974 = pi5  & ~n37971;
  assign n37975 = pi5  & n37970;
  assign n37976 = ~n58251 & ~n58252;
  assign n37977 = pi8  & ~n58077;
  assign n37978 = ~n58078 & ~n37977;
  assign n37979 = n58078 & n37977;
  assign n37980 = ~n58077 & n37069;
  assign n37981 = ~n58079 & ~n37980;
  assign n37982 = ~n37978 & ~n37979;
  assign n37983 = ~n37976 & n58253;
  assign n37984 = n77 & n30866;
  assign n37985 = n24302 & n26337;
  assign n37986 = n21969 & n26343;
  assign n37987 = n23459 & n26340;
  assign n37988 = ~n37986 & ~n37987;
  assign n37989 = ~n37985 & n37988;
  assign n37990 = ~n77 & n37989;
  assign n37991 = ~n30866 & n37989;
  assign n37992 = ~n37990 & ~n37991;
  assign n37993 = ~n37984 & n37989;
  assign n37994 = pi5  & ~n58254;
  assign n37995 = ~pi5  & n58254;
  assign n37996 = ~n37994 & ~n37995;
  assign n37997 = pi8  & n37049;
  assign n37998 = ~n37048 & n37997;
  assign n37999 = n37048 & ~n37997;
  assign n38000 = ~n37050 & n37054;
  assign n38001 = ~n58077 & ~n38000;
  assign n38002 = ~n37998 & ~n37999;
  assign n38003 = ~n37996 & n58255;
  assign n38004 = n77 & ~n31019;
  assign n38005 = n23459 & ~n56543;
  assign n38006 = n24302 & n26348;
  assign n38007 = ~n38005 & ~n38006;
  assign n38008 = ~n38004 & n38007;
  assign n38009 = n53439 & ~n56543;
  assign n38010 = pi5  & ~n38009;
  assign n38011 = pi5  & ~n38008;
  assign n38012 = pi5  & ~n38011;
  assign n38013 = ~n38008 & ~n38011;
  assign n38014 = ~n38012 & ~n38013;
  assign n38015 = n38010 & ~n38014;
  assign n38016 = n38008 & n38010;
  assign n38017 = n77 & ~n31140;
  assign n38018 = n24302 & n26343;
  assign n38019 = n21969 & ~n56543;
  assign n38020 = n23459 & n26348;
  assign n38021 = ~n38019 & ~n38020;
  assign n38022 = ~n38018 & n38021;
  assign n38023 = ~n77 & n38022;
  assign n38024 = n31140 & n38022;
  assign n38025 = ~n38023 & ~n38024;
  assign n38026 = ~n38017 & n38022;
  assign n38027 = pi5  & ~n58257;
  assign n38028 = ~pi5  & n58257;
  assign n38029 = ~n38027 & ~n38028;
  assign n38030 = n58256 & ~n38029;
  assign n38031 = n58256 & ~n58257;
  assign n38032 = n37049 & n58258;
  assign n38033 = n77 & n30915;
  assign n38034 = n24302 & n26340;
  assign n38035 = n21969 & n26348;
  assign n38036 = n23459 & n26343;
  assign n38037 = ~n38035 & ~n38036;
  assign n38038 = ~n38034 & n38037;
  assign n38039 = ~n38033 & n38038;
  assign n38040 = pi5  & ~n38039;
  assign n38041 = pi5  & ~n38040;
  assign n38042 = pi5  & n38039;
  assign n38043 = ~n38039 & ~n38040;
  assign n38044 = ~pi5  & ~n38039;
  assign n38045 = ~n58259 & ~n58260;
  assign n38046 = ~n37049 & ~n58258;
  assign n38047 = n58258 & ~n38032;
  assign n38048 = ~n37049 & n58258;
  assign n38049 = n37049 & ~n38032;
  assign n38050 = n37049 & ~n58258;
  assign n38051 = ~n58261 & ~n58262;
  assign n38052 = ~n38032 & ~n38046;
  assign n38053 = ~n38045 & ~n58263;
  assign n38054 = ~n38032 & ~n38053;
  assign n38055 = n37996 & ~n58255;
  assign n38056 = ~n38003 & ~n38055;
  assign n38057 = ~n38054 & n38056;
  assign n38058 = ~n38003 & ~n38057;
  assign n38059 = n37976 & ~n58253;
  assign n38060 = ~n37976 & ~n37983;
  assign n38061 = ~n37976 & ~n58253;
  assign n38062 = n58253 & ~n37983;
  assign n38063 = n37976 & n58253;
  assign n38064 = ~n58264 & ~n58265;
  assign n38065 = ~n37983 & ~n38059;
  assign n38066 = ~n38058 & ~n58266;
  assign n38067 = ~n37983 & ~n38066;
  assign n38068 = n37957 & n58250;
  assign n38069 = ~n37963 & ~n38068;
  assign n38070 = ~n38067 & n38069;
  assign n38071 = ~n37963 & ~n38070;
  assign n38072 = n37941 & ~n37943;
  assign n38073 = ~n37941 & ~n37944;
  assign n38074 = ~n37941 & ~n37943;
  assign n38075 = n37943 & ~n37944;
  assign n38076 = n37941 & n37943;
  assign n38077 = ~n58267 & ~n58268;
  assign n38078 = ~n37944 & ~n38072;
  assign n38079 = ~n38071 & ~n58269;
  assign n38080 = ~n37944 & ~n38079;
  assign n38081 = ~n37914 & n37927;
  assign n38082 = n37914 & ~n37928;
  assign n38083 = n37914 & n37927;
  assign n38084 = ~n37927 & ~n37928;
  assign n38085 = ~n37914 & ~n37927;
  assign n38086 = ~n58270 & ~n58271;
  assign n38087 = ~n37928 & ~n38081;
  assign n38088 = ~n38080 & ~n58272;
  assign n38089 = ~n37928 & ~n38088;
  assign n38090 = ~n37898 & n37911;
  assign n38091 = n37898 & ~n37912;
  assign n38092 = n37898 & n37911;
  assign n38093 = ~n37911 & ~n37912;
  assign n38094 = ~n37898 & ~n37911;
  assign n38095 = ~n58273 & ~n58274;
  assign n38096 = ~n37912 & ~n38090;
  assign n38097 = ~n38089 & ~n58275;
  assign n38098 = ~n37912 & ~n38097;
  assign n38099 = ~n37882 & n37895;
  assign n38100 = ~n37896 & ~n38099;
  assign n38101 = ~n38098 & n38100;
  assign n38102 = ~n37896 & ~n38101;
  assign n38103 = n37872 & n58243;
  assign n38104 = ~n37872 & ~n37880;
  assign n38105 = ~n58243 & ~n37880;
  assign n38106 = ~n38104 & ~n38105;
  assign n38107 = ~n37880 & ~n38103;
  assign n38108 = ~n38102 & ~n58276;
  assign n38109 = ~n37880 & ~n38108;
  assign n38110 = n37853 & n58238;
  assign n38111 = ~n37853 & ~n37859;
  assign n38112 = ~n37853 & n58238;
  assign n38113 = ~n58238 & ~n37859;
  assign n38114 = n37853 & ~n58238;
  assign n38115 = ~n58277 & ~n58278;
  assign n38116 = ~n37859 & ~n38110;
  assign n38117 = ~n38109 & ~n58279;
  assign n38118 = ~n37859 & ~n38117;
  assign n38119 = n37837 & ~n37839;
  assign n38120 = ~n37837 & ~n37840;
  assign n38121 = ~n37837 & ~n37839;
  assign n38122 = n37839 & ~n37840;
  assign n38123 = n37837 & n37839;
  assign n38124 = ~n58280 & ~n58281;
  assign n38125 = ~n37840 & ~n38119;
  assign n38126 = ~n38118 & ~n58282;
  assign n38127 = ~n37840 & ~n38126;
  assign n38128 = ~n37810 & n37823;
  assign n38129 = n37810 & ~n37824;
  assign n38130 = n37810 & n37823;
  assign n38131 = ~n37823 & ~n37824;
  assign n38132 = ~n37810 & ~n37823;
  assign n38133 = ~n58283 & ~n58284;
  assign n38134 = ~n37824 & ~n38128;
  assign n38135 = ~n38127 & ~n58285;
  assign n38136 = ~n37824 & ~n38135;
  assign n38137 = ~n37794 & n37807;
  assign n38138 = n37794 & ~n37808;
  assign n38139 = n37794 & n37807;
  assign n38140 = ~n37807 & ~n37808;
  assign n38141 = ~n37794 & ~n37807;
  assign n38142 = ~n58286 & ~n58287;
  assign n38143 = ~n37808 & ~n38137;
  assign n38144 = ~n38136 & ~n58288;
  assign n38145 = ~n37808 & ~n38144;
  assign n38146 = ~n37778 & n37791;
  assign n38147 = ~n37792 & ~n38146;
  assign n38148 = ~n38145 & n38147;
  assign n38149 = ~n37792 & ~n38148;
  assign n38150 = n37770 & n58230;
  assign n38151 = ~n37770 & ~n37776;
  assign n38152 = ~n37770 & n58230;
  assign n38153 = ~n58230 & ~n37776;
  assign n38154 = n37770 & ~n58230;
  assign n38155 = ~n58289 & ~n58290;
  assign n38156 = ~n37776 & ~n38150;
  assign n38157 = ~n38149 & ~n58291;
  assign n38158 = ~n37776 & ~n38157;
  assign n38159 = n37749 & n58227;
  assign n38160 = ~n37749 & ~n37757;
  assign n38161 = ~n58227 & ~n37757;
  assign n38162 = ~n38160 & ~n38161;
  assign n38163 = ~n37757 & ~n38159;
  assign n38164 = ~n38158 & ~n58292;
  assign n38165 = ~n37757 & ~n38164;
  assign n38166 = n37733 & ~n37735;
  assign n38167 = ~n37733 & ~n37736;
  assign n38168 = ~n37733 & ~n37735;
  assign n38169 = n37735 & ~n37736;
  assign n38170 = n37733 & n37735;
  assign n38171 = ~n58293 & ~n58294;
  assign n38172 = ~n37736 & ~n38166;
  assign n38173 = ~n38165 & ~n58295;
  assign n38174 = ~n37736 & ~n38173;
  assign n38175 = ~n37706 & n37719;
  assign n38176 = n37706 & ~n37720;
  assign n38177 = n37706 & n37719;
  assign n38178 = ~n37719 & ~n37720;
  assign n38179 = ~n37706 & ~n37719;
  assign n38180 = ~n58296 & ~n58297;
  assign n38181 = ~n37720 & ~n38175;
  assign n38182 = ~n38174 & ~n58298;
  assign n38183 = ~n37720 & ~n38182;
  assign n38184 = ~n37690 & n37703;
  assign n38185 = n37690 & ~n37704;
  assign n38186 = n37690 & n37703;
  assign n38187 = ~n37703 & ~n37704;
  assign n38188 = ~n37690 & ~n37703;
  assign n38189 = ~n58299 & ~n58300;
  assign n38190 = ~n37704 & ~n38184;
  assign n38191 = ~n38183 & ~n58301;
  assign n38192 = ~n37704 & ~n38191;
  assign n38193 = ~n37674 & n37687;
  assign n38194 = ~n37688 & ~n38193;
  assign n38195 = ~n38192 & n38194;
  assign n38196 = ~n37688 & ~n38195;
  assign n38197 = n37664 & n58217;
  assign n38198 = ~n37664 & ~n37672;
  assign n38199 = ~n58217 & ~n37672;
  assign n38200 = ~n38198 & ~n38199;
  assign n38201 = ~n37672 & ~n38197;
  assign n38202 = ~n38196 & ~n58302;
  assign n38203 = ~n37672 & ~n38202;
  assign n38204 = n37645 & n58212;
  assign n38205 = ~n37645 & ~n37651;
  assign n38206 = ~n37645 & n58212;
  assign n38207 = ~n58212 & ~n37651;
  assign n38208 = n37645 & ~n58212;
  assign n38209 = ~n58303 & ~n58304;
  assign n38210 = ~n37651 & ~n38204;
  assign n38211 = ~n38203 & ~n58305;
  assign n38212 = ~n37651 & ~n38211;
  assign n38213 = n37629 & ~n37631;
  assign n38214 = ~n37629 & ~n37632;
  assign n38215 = ~n37629 & ~n37631;
  assign n38216 = n37631 & ~n37632;
  assign n38217 = n37629 & n37631;
  assign n38218 = ~n58306 & ~n58307;
  assign n38219 = ~n37632 & ~n38213;
  assign n38220 = ~n38212 & ~n58308;
  assign n38221 = ~n37632 & ~n38220;
  assign n38222 = ~n37602 & n37615;
  assign n38223 = n37602 & ~n37616;
  assign n38224 = n37602 & n37615;
  assign n38225 = ~n37615 & ~n37616;
  assign n38226 = ~n37602 & ~n37615;
  assign n38227 = ~n58309 & ~n58310;
  assign n38228 = ~n37616 & ~n38222;
  assign n38229 = ~n38221 & ~n58311;
  assign n38230 = ~n37616 & ~n38229;
  assign n38231 = ~n37586 & n37599;
  assign n38232 = ~n37600 & ~n38231;
  assign n38233 = ~n38230 & n38232;
  assign n38234 = ~n37600 & ~n38233;
  assign n38235 = n37576 & n58205;
  assign n38236 = ~n37576 & ~n37584;
  assign n38237 = ~n58205 & ~n37584;
  assign n38238 = ~n38236 & ~n38237;
  assign n38239 = ~n37584 & ~n38235;
  assign n38240 = ~n38234 & ~n58312;
  assign n38241 = ~n37584 & ~n38240;
  assign n38242 = n37555 & n58200;
  assign n38243 = ~n37555 & ~n37563;
  assign n38244 = ~n58200 & ~n37563;
  assign n38245 = ~n38243 & ~n38244;
  assign n38246 = ~n37563 & ~n38242;
  assign n38247 = ~n38241 & ~n58313;
  assign n38248 = ~n37563 & ~n38247;
  assign n38249 = n37536 & n58195;
  assign n38250 = ~n37536 & ~n37542;
  assign n38251 = ~n37536 & n58195;
  assign n38252 = ~n58195 & ~n37542;
  assign n38253 = n37536 & ~n58195;
  assign n38254 = ~n58314 & ~n58315;
  assign n38255 = ~n37542 & ~n38249;
  assign n38256 = ~n38248 & ~n58316;
  assign n38257 = ~n37542 & ~n38256;
  assign n38258 = n37517 & n58192;
  assign n38259 = ~n37517 & ~n37523;
  assign n38260 = ~n37517 & n58192;
  assign n38261 = ~n58192 & ~n37523;
  assign n38262 = n37517 & ~n58192;
  assign n38263 = ~n58317 & ~n58318;
  assign n38264 = ~n37523 & ~n38258;
  assign n38265 = ~n38257 & ~n58319;
  assign n38266 = ~n37523 & ~n38265;
  assign n38267 = n37498 & n58189;
  assign n38268 = ~n37498 & ~n37504;
  assign n38269 = ~n37498 & n58189;
  assign n38270 = ~n58189 & ~n37504;
  assign n38271 = n37498 & ~n58189;
  assign n38272 = ~n58320 & ~n58321;
  assign n38273 = ~n37504 & ~n38267;
  assign n38274 = ~n38266 & ~n58322;
  assign n38275 = ~n37504 & ~n38274;
  assign n38276 = n37477 & n58186;
  assign n38277 = ~n37477 & ~n37485;
  assign n38278 = ~n58186 & ~n37485;
  assign n38279 = ~n38277 & ~n38278;
  assign n38280 = ~n37485 & ~n38276;
  assign n38281 = ~n38275 & ~n58323;
  assign n38282 = ~n37485 & ~n38281;
  assign n38283 = n37456 & n58181;
  assign n38284 = ~n37456 & ~n37464;
  assign n38285 = ~n58181 & ~n37464;
  assign n38286 = ~n38284 & ~n38285;
  assign n38287 = ~n37464 & ~n38283;
  assign n38288 = ~n38282 & ~n58324;
  assign n38289 = ~n37464 & ~n38288;
  assign n38290 = n37435 & n58176;
  assign n38291 = ~n37435 & ~n37443;
  assign n38292 = ~n58176 & ~n37443;
  assign n38293 = ~n38291 & ~n38292;
  assign n38294 = ~n37443 & ~n38290;
  assign n38295 = ~n38289 & ~n58325;
  assign n38296 = ~n37443 & ~n38295;
  assign n38297 = n37414 & n58171;
  assign n38298 = ~n37414 & ~n37422;
  assign n38299 = ~n58171 & ~n37422;
  assign n38300 = ~n38298 & ~n38299;
  assign n38301 = ~n37422 & ~n38297;
  assign n38302 = ~n38296 & ~n58326;
  assign n38303 = ~n37422 & ~n38302;
  assign n38304 = ~n56855 & n58163;
  assign n38305 = ~n58163 & ~n37390;
  assign n38306 = n56855 & ~n37390;
  assign n38307 = ~n38305 & ~n38306;
  assign n38308 = ~n37390 & ~n38304;
  assign n38309 = ~n38303 & ~n58327;
  assign n38310 = n38303 & n58327;
  assign n38311 = ~n38309 & ~n38310;
  assign n38312 = n38296 & n58326;
  assign n38313 = ~n38302 & ~n38312;
  assign n38314 = pi2  & n29078;
  assign n38315 = ~n56855 & ~n38314;
  assign n38316 = n38313 & ~n38315;
  assign n38317 = n38289 & n58325;
  assign n38318 = ~n38295 & ~n38317;
  assign n38319 = n24338 & n28624;
  assign n38320 = n25272 & ~n26537;
  assign n38321 = n24337 & n26242;
  assign n38322 = ~n25287 & ~n38321;
  assign n38323 = ~n38320 & ~n38321;
  assign n38324 = ~n25287 & n38323;
  assign n38325 = ~n38320 & n38322;
  assign n38326 = ~n24338 & n58328;
  assign n38327 = ~n28624 & n58328;
  assign n38328 = ~n38326 & ~n38327;
  assign n38329 = ~n38319 & n58328;
  assign n38330 = pi2  & ~n58329;
  assign n38331 = ~pi2  & n58329;
  assign n38332 = ~n38330 & ~n38331;
  assign n38333 = n38318 & ~n38332;
  assign n38334 = n38282 & n58324;
  assign n38335 = ~n38288 & ~n38334;
  assign n38336 = n24338 & ~n56564;
  assign n38337 = n25287 & ~n26537;
  assign n38338 = n24337 & n26244;
  assign n38339 = n25272 & n26242;
  assign n38340 = ~n38338 & ~n38339;
  assign n38341 = ~n38337 & n38340;
  assign n38342 = ~n24338 & n38341;
  assign n38343 = n56564 & n38341;
  assign n38344 = ~n38342 & ~n38343;
  assign n38345 = ~n38336 & n38341;
  assign n38346 = pi2  & ~n58330;
  assign n38347 = ~pi2  & n58330;
  assign n38348 = ~n38346 & ~n38347;
  assign n38349 = n38335 & ~n38348;
  assign n38350 = n38275 & n58323;
  assign n38351 = ~n38281 & ~n38350;
  assign n38352 = n24338 & n27808;
  assign n38353 = n25287 & n26242;
  assign n38354 = n24337 & n26247;
  assign n38355 = n25272 & n26244;
  assign n38356 = ~n38354 & ~n38355;
  assign n38357 = ~n38353 & n38356;
  assign n38358 = ~n24338 & n38357;
  assign n38359 = ~n27808 & n38357;
  assign n38360 = ~n38358 & ~n38359;
  assign n38361 = ~n38352 & n38357;
  assign n38362 = pi2  & ~n58331;
  assign n38363 = ~pi2  & n58331;
  assign n38364 = ~n38362 & ~n38363;
  assign n38365 = n38351 & ~n38364;
  assign n38366 = n38266 & n58322;
  assign n38367 = ~n38274 & ~n38366;
  assign n38368 = n24338 & n27839;
  assign n38369 = n25287 & n26244;
  assign n38370 = n24337 & n26250;
  assign n38371 = n25272 & n26247;
  assign n38372 = ~n38370 & ~n38371;
  assign n38373 = ~n38369 & n38372;
  assign n38374 = ~n24338 & n38373;
  assign n38375 = ~n27839 & n38373;
  assign n38376 = ~n38374 & ~n38375;
  assign n38377 = ~n38368 & n38373;
  assign n38378 = pi2  & ~n58332;
  assign n38379 = ~pi2  & n58332;
  assign n38380 = ~n38378 & ~n38379;
  assign n38381 = n38367 & ~n38380;
  assign n38382 = n38257 & n58319;
  assign n38383 = ~n38265 & ~n38382;
  assign n38384 = n24338 & ~n56567;
  assign n38385 = n25287 & n26247;
  assign n38386 = n24337 & n26253;
  assign n38387 = n25272 & n26250;
  assign n38388 = ~n38386 & ~n38387;
  assign n38389 = ~n38385 & n38388;
  assign n38390 = ~n24338 & n38389;
  assign n38391 = n56567 & n38389;
  assign n38392 = ~n38390 & ~n38391;
  assign n38393 = ~n38384 & n38389;
  assign n38394 = pi2  & ~n58333;
  assign n38395 = ~pi2  & n58333;
  assign n38396 = ~n38394 & ~n38395;
  assign n38397 = n38383 & ~n38396;
  assign n38398 = n38248 & n58316;
  assign n38399 = ~n38256 & ~n38398;
  assign n38400 = n24338 & n27491;
  assign n38401 = n25287 & n26250;
  assign n38402 = n24337 & n26256;
  assign n38403 = n25272 & n26253;
  assign n38404 = ~n38402 & ~n38403;
  assign n38405 = ~n38401 & n38404;
  assign n38406 = ~n24338 & n38405;
  assign n38407 = ~n27491 & n38405;
  assign n38408 = ~n38406 & ~n38407;
  assign n38409 = ~n38400 & n38405;
  assign n38410 = pi2  & ~n58334;
  assign n38411 = ~pi2  & n58334;
  assign n38412 = ~n38410 & ~n38411;
  assign n38413 = n38399 & ~n38412;
  assign n38414 = n38241 & n58313;
  assign n38415 = ~n38247 & ~n38414;
  assign n38416 = n24338 & ~n56668;
  assign n38417 = n25287 & n26253;
  assign n38418 = n24337 & n26259;
  assign n38419 = n25272 & n26256;
  assign n38420 = ~n38418 & ~n38419;
  assign n38421 = ~n38417 & n38420;
  assign n38422 = ~n24338 & n38421;
  assign n38423 = n56668 & n38421;
  assign n38424 = ~n38422 & ~n38423;
  assign n38425 = ~n38416 & n38421;
  assign n38426 = pi2  & ~n58335;
  assign n38427 = ~pi2  & n58335;
  assign n38428 = ~n38426 & ~n38427;
  assign n38429 = n38415 & ~n38428;
  assign n38430 = n38234 & n58312;
  assign n38431 = ~n38240 & ~n38430;
  assign n38432 = n24338 & n27387;
  assign n38433 = n25287 & n26256;
  assign n38434 = n24337 & n26262;
  assign n38435 = n25272 & n26259;
  assign n38436 = ~n38434 & ~n38435;
  assign n38437 = ~n38433 & n38436;
  assign n38438 = ~n24338 & n38437;
  assign n38439 = ~n27387 & n38437;
  assign n38440 = ~n38438 & ~n38439;
  assign n38441 = ~n38432 & n38437;
  assign n38442 = pi2  & ~n58336;
  assign n38443 = ~pi2  & n58336;
  assign n38444 = ~n38442 & ~n38443;
  assign n38445 = n38431 & ~n38444;
  assign n38446 = ~n38431 & n38444;
  assign n38447 = n38431 & ~n38445;
  assign n38448 = n38431 & n38444;
  assign n38449 = ~n38444 & ~n38445;
  assign n38450 = ~n38431 & ~n38444;
  assign n38451 = ~n58337 & ~n58338;
  assign n38452 = ~n38445 & ~n38446;
  assign n38453 = n38230 & ~n38232;
  assign n38454 = ~n38233 & ~n38453;
  assign n38455 = n38221 & ~n58310;
  assign n38456 = ~n58309 & n38455;
  assign n38457 = n38221 & n58311;
  assign n38458 = ~n38229 & ~n58340;
  assign n38459 = n38212 & n58308;
  assign n38460 = ~n38220 & ~n38459;
  assign n38461 = n38203 & n58305;
  assign n38462 = ~n38211 & ~n38461;
  assign n38463 = n24338 & ~n56612;
  assign n38464 = n25287 & n26271;
  assign n38465 = n24337 & n26277;
  assign n38466 = n25272 & n26274;
  assign n38467 = ~n38465 & ~n38466;
  assign n38468 = ~n38464 & n38467;
  assign n38469 = ~n24338 & n38468;
  assign n38470 = n56612 & n38468;
  assign n38471 = ~n38469 & ~n38470;
  assign n38472 = ~n38463 & n38468;
  assign n38473 = pi2  & ~n58341;
  assign n38474 = ~pi2  & n58341;
  assign n38475 = ~n38473 & ~n38474;
  assign n38476 = n38196 & n58302;
  assign n38477 = ~n38202 & ~n38476;
  assign n38478 = n38475 & ~n38477;
  assign n38479 = ~n38475 & n38477;
  assign n38480 = n38183 & ~n58300;
  assign n38481 = ~n58299 & n38480;
  assign n38482 = n38183 & n58301;
  assign n38483 = ~n38191 & ~n58342;
  assign n38484 = n38174 & ~n58297;
  assign n38485 = ~n58296 & n38484;
  assign n38486 = n38174 & n58298;
  assign n38487 = ~n38182 & ~n58343;
  assign n38488 = n38165 & n58295;
  assign n38489 = ~n38173 & ~n38488;
  assign n38490 = n38158 & n58292;
  assign n38491 = ~n38164 & ~n38490;
  assign n38492 = n24338 & n28107;
  assign n38493 = n25287 & n26289;
  assign n38494 = n24337 & n26295;
  assign n38495 = n25272 & n26292;
  assign n38496 = ~n38494 & ~n38495;
  assign n38497 = ~n38493 & n38496;
  assign n38498 = ~n24338 & n38497;
  assign n38499 = ~n28107 & n38497;
  assign n38500 = ~n38498 & ~n38499;
  assign n38501 = ~n38492 & n38497;
  assign n38502 = pi2  & ~n58344;
  assign n38503 = ~pi2  & n58344;
  assign n38504 = ~n38502 & ~n38503;
  assign n38505 = n38149 & n58291;
  assign n38506 = ~n38157 & ~n38505;
  assign n38507 = n38504 & ~n38506;
  assign n38508 = ~n38504 & n38506;
  assign n38509 = n38136 & ~n58287;
  assign n38510 = ~n58286 & n38509;
  assign n38511 = n38136 & n58288;
  assign n38512 = ~n38144 & ~n58345;
  assign n38513 = n38127 & ~n58284;
  assign n38514 = ~n58283 & n38513;
  assign n38515 = n38127 & n58285;
  assign n38516 = ~n38135 & ~n58346;
  assign n38517 = n38118 & n58282;
  assign n38518 = ~n38126 & ~n38517;
  assign n38519 = n38109 & n58279;
  assign n38520 = ~n38117 & ~n38519;
  assign n38521 = n24338 & ~n56928;
  assign n38522 = n25287 & n26307;
  assign n38523 = n24337 & n26313;
  assign n38524 = n25272 & n26310;
  assign n38525 = ~n38523 & ~n38524;
  assign n38526 = ~n38522 & n38525;
  assign n38527 = ~n24338 & n38526;
  assign n38528 = n56928 & n38526;
  assign n38529 = ~n38527 & ~n38528;
  assign n38530 = ~n38521 & n38526;
  assign n38531 = pi2  & ~n58347;
  assign n38532 = ~pi2  & n58347;
  assign n38533 = ~n38531 & ~n38532;
  assign n38534 = n38102 & n58276;
  assign n38535 = ~n38108 & ~n38534;
  assign n38536 = n38533 & ~n38535;
  assign n38537 = ~n38533 & n38535;
  assign n38538 = n38089 & ~n58274;
  assign n38539 = ~n58273 & n38538;
  assign n38540 = n38089 & n58275;
  assign n38541 = ~n38097 & ~n58348;
  assign n38542 = n38080 & ~n58271;
  assign n38543 = ~n58270 & n38542;
  assign n38544 = n38080 & n58272;
  assign n38545 = ~n38088 & ~n58349;
  assign n38546 = n38071 & n58269;
  assign n38547 = ~n38079 & ~n38546;
  assign n38548 = n38067 & ~n38069;
  assign n38549 = ~n38070 & ~n38548;
  assign n38550 = n24338 & ~n57017;
  assign n38551 = n25287 & n26325;
  assign n38552 = n24337 & n26331;
  assign n38553 = n25272 & n26328;
  assign n38554 = ~n38552 & ~n38553;
  assign n38555 = ~n38551 & n38554;
  assign n38556 = ~n24338 & n38555;
  assign n38557 = n57017 & n38555;
  assign n38558 = ~n38556 & ~n38557;
  assign n38559 = ~n38550 & n38555;
  assign n38560 = pi2  & ~n58350;
  assign n38561 = ~pi2  & n58350;
  assign n38562 = ~n38560 & ~n38561;
  assign n38563 = n38058 & n58266;
  assign n38564 = ~n38066 & ~n38563;
  assign n38565 = n38562 & ~n38564;
  assign n38566 = ~n38562 & n38564;
  assign n38567 = n24338 & ~n57033;
  assign n38568 = n25287 & n26331;
  assign n38569 = n24337 & n26337;
  assign n38570 = n25272 & n26334;
  assign n38571 = ~n38569 & ~n38570;
  assign n38572 = ~n38568 & n38571;
  assign n38573 = ~n24338 & n38572;
  assign n38574 = n57033 & n38572;
  assign n38575 = ~n38573 & ~n38574;
  assign n38576 = ~n38567 & n38572;
  assign n38577 = pi2  & ~n58351;
  assign n38578 = ~pi2  & n58351;
  assign n38579 = ~n38577 & ~n38578;
  assign n38580 = n38045 & n58263;
  assign n38581 = ~n38053 & ~n38580;
  assign n38582 = n38579 & ~n38581;
  assign n38583 = ~n38579 & n38581;
  assign n38584 = pi5  & ~n58256;
  assign n38585 = ~n58257 & ~n38584;
  assign n38586 = n58257 & n38584;
  assign n38587 = ~n58256 & n38029;
  assign n38588 = ~n58258 & ~n38587;
  assign n38589 = ~n38585 & ~n38586;
  assign n38590 = n24338 & ~n57042;
  assign n38591 = n25287 & n26334;
  assign n38592 = n24337 & n26340;
  assign n38593 = n25272 & n26337;
  assign n38594 = ~n38592 & ~n38593;
  assign n38595 = ~n38591 & n38594;
  assign n38596 = ~n38590 & n38595;
  assign n38597 = pi2  & ~n38596;
  assign n38598 = ~pi2  & n38596;
  assign n38599 = ~pi2  & ~n38596;
  assign n38600 = pi2  & n38596;
  assign n38601 = ~n38599 & ~n38600;
  assign n38602 = ~n38597 & ~n38598;
  assign n38603 = n58352 & ~n58353;
  assign n38604 = n24338 & n30866;
  assign n38605 = n25287 & n26337;
  assign n38606 = n25272 & n26340;
  assign n38607 = n24337 & n26343;
  assign n38608 = ~n38606 & ~n38607;
  assign n38609 = ~n38605 & n38608;
  assign n38610 = ~n24338 & n38609;
  assign n38611 = ~n30866 & n38609;
  assign n38612 = ~n38610 & ~n38611;
  assign n38613 = ~n38604 & n38609;
  assign n38614 = pi2  & ~n58354;
  assign n38615 = ~pi2  & n58354;
  assign n38616 = ~n38614 & ~n38615;
  assign n38617 = ~n26343 & n31019;
  assign n38618 = n24338 & ~n38617;
  assign n38619 = n25287 & n26343;
  assign n38620 = n26348 & ~n56852;
  assign n38621 = pi2  & n56543;
  assign n38622 = ~n38620 & n38621;
  assign n38623 = ~n38619 & n38622;
  assign n38624 = pi0  & ~n56543;
  assign n38625 = n25558 & ~n31140;
  assign n38626 = n24337 & ~n56543;
  assign n38627 = n25272 & n26348;
  assign n38628 = ~n38626 & ~n38627;
  assign n38629 = ~n38619 & n38628;
  assign n38630 = pi2  & ~n38629;
  assign n38631 = n25558 & ~n31019;
  assign n38632 = n25569 & ~n56543;
  assign n38633 = n25571 & n26348;
  assign n38634 = pi2  & ~n38633;
  assign n38635 = ~n38632 & n38634;
  assign n38636 = ~n38631 & n38635;
  assign n38637 = ~n38630 & n38636;
  assign n38638 = ~n38625 & n38637;
  assign n38639 = ~n38624 & n38638;
  assign n38640 = ~n24330 & ~n56543;
  assign n38641 = pi2  & ~n38624;
  assign n38642 = ~n38632 & n38641;
  assign n38643 = pi2  & ~n38640;
  assign n38644 = ~n38633 & n58356;
  assign n38645 = ~n38631 & n38644;
  assign n38646 = ~n38630 & n38645;
  assign n38647 = ~n38625 & n38646;
  assign n38648 = ~n38625 & n38645;
  assign n38649 = ~n38630 & n38648;
  assign n38650 = ~n38618 & n38623;
  assign n38651 = ~n38009 & ~n58355;
  assign n38652 = n24338 & n30915;
  assign n38653 = n25287 & n26340;
  assign n38654 = n24337 & n26348;
  assign n38655 = n25272 & n26343;
  assign n38656 = ~n38654 & ~n38655;
  assign n38657 = ~n38653 & n38656;
  assign n38658 = ~n38652 & n38657;
  assign n38659 = ~pi2  & ~n38658;
  assign n38660 = pi2  & n38658;
  assign n38661 = pi2  & ~n38658;
  assign n38662 = ~pi2  & n38658;
  assign n38663 = ~n38661 & ~n38662;
  assign n38664 = ~n38659 & ~n38660;
  assign n38665 = ~n38651 & n58357;
  assign n38666 = ~n38616 & n38665;
  assign n38667 = n38616 & ~n38665;
  assign n38668 = pi5  & n38009;
  assign n38669 = n38008 & ~n38668;
  assign n38670 = ~n38008 & n38668;
  assign n38671 = ~n38010 & n38014;
  assign n38672 = ~n58256 & ~n38671;
  assign n38673 = ~n38669 & ~n38670;
  assign n38674 = ~n38667 & n58358;
  assign n38675 = ~n38666 & ~n38674;
  assign n38676 = ~n38603 & n38675;
  assign n38677 = ~n58352 & n58353;
  assign n38678 = n58352 & ~n38675;
  assign n38679 = ~n58352 & n38675;
  assign n38680 = ~n58353 & ~n38679;
  assign n38681 = ~n38678 & ~n38680;
  assign n38682 = ~n38676 & ~n38677;
  assign n38683 = ~n38583 & n58359;
  assign n38684 = ~n38579 & ~n58359;
  assign n38685 = n38579 & n58359;
  assign n38686 = n38581 & ~n38685;
  assign n38687 = ~n38684 & ~n38686;
  assign n38688 = ~n38582 & ~n38683;
  assign n38689 = n38054 & ~n38056;
  assign n38690 = ~n38057 & ~n38689;
  assign n38691 = n24338 & n30470;
  assign n38692 = n25287 & n26328;
  assign n38693 = n24337 & n26334;
  assign n38694 = n25272 & n26331;
  assign n38695 = ~n38693 & ~n38694;
  assign n38696 = ~n38692 & n38695;
  assign n38697 = ~n38691 & n38696;
  assign n38698 = pi2  & ~n38697;
  assign n38699 = ~pi2  & n38697;
  assign n38700 = ~pi2  & ~n38697;
  assign n38701 = pi2  & n38697;
  assign n38702 = ~n38700 & ~n38701;
  assign n38703 = ~n38698 & ~n38699;
  assign n38704 = n38690 & ~n58361;
  assign n38705 = n58360 & ~n38704;
  assign n38706 = ~n38690 & n58361;
  assign n38707 = ~n58360 & n38690;
  assign n38708 = n58360 & ~n38690;
  assign n38709 = ~n58361 & ~n38708;
  assign n38710 = ~n38707 & ~n38709;
  assign n38711 = ~n38705 & ~n38706;
  assign n38712 = ~n38566 & ~n38707;
  assign n38713 = ~n38709 & n38712;
  assign n38714 = ~n38566 & n58362;
  assign n38715 = n38562 & n58362;
  assign n38716 = n38564 & ~n38715;
  assign n38717 = ~n38562 & ~n58362;
  assign n38718 = ~n38716 & ~n38717;
  assign n38719 = ~n38565 & ~n58363;
  assign n38720 = ~n38549 & n58364;
  assign n38721 = n38549 & ~n58364;
  assign n38722 = n24338 & ~n57012;
  assign n38723 = n25287 & n26322;
  assign n38724 = n24337 & n26328;
  assign n38725 = n25272 & n26325;
  assign n38726 = ~n38724 & ~n38725;
  assign n38727 = ~n38723 & n38726;
  assign n38728 = ~n24338 & n38727;
  assign n38729 = n57012 & n38727;
  assign n38730 = ~n38728 & ~n38729;
  assign n38731 = ~n38722 & n38727;
  assign n38732 = pi2  & ~n58365;
  assign n38733 = ~pi2  & n58365;
  assign n38734 = ~n38732 & ~n38733;
  assign n38735 = ~n38721 & n38734;
  assign n38736 = n58364 & n38734;
  assign n38737 = n38549 & ~n38736;
  assign n38738 = ~n58364 & ~n38734;
  assign n38739 = ~n38737 & ~n38738;
  assign n38740 = ~n38720 & ~n38735;
  assign n38741 = ~n38547 & n58366;
  assign n38742 = n38547 & ~n58366;
  assign n38743 = n24338 & n30264;
  assign n38744 = n25287 & n26319;
  assign n38745 = n24337 & n26325;
  assign n38746 = n25272 & n26322;
  assign n38747 = ~n38745 & ~n38746;
  assign n38748 = ~n38744 & n38747;
  assign n38749 = ~n24338 & n38748;
  assign n38750 = ~n30264 & n38748;
  assign n38751 = ~n38749 & ~n38750;
  assign n38752 = ~n38743 & n38748;
  assign n38753 = pi2  & ~n58367;
  assign n38754 = ~pi2  & n58367;
  assign n38755 = ~n38753 & ~n38754;
  assign n38756 = ~n38742 & n38755;
  assign n38757 = n58366 & n38755;
  assign n38758 = n38547 & ~n38757;
  assign n38759 = ~n58366 & ~n38755;
  assign n38760 = ~n38758 & ~n38759;
  assign n38761 = ~n38741 & ~n38756;
  assign n38762 = n38545 & ~n58368;
  assign n38763 = ~n38545 & n58368;
  assign n38764 = n24338 & ~n56920;
  assign n38765 = n25287 & n26316;
  assign n38766 = n24337 & n26322;
  assign n38767 = n25272 & n26319;
  assign n38768 = ~n38766 & ~n38767;
  assign n38769 = ~n38765 & n38768;
  assign n38770 = ~n38764 & n38769;
  assign n38771 = pi2  & ~n38770;
  assign n38772 = ~pi2  & n38770;
  assign n38773 = ~pi2  & ~n38770;
  assign n38774 = pi2  & n38770;
  assign n38775 = ~n38773 & ~n38774;
  assign n38776 = ~n38771 & ~n38772;
  assign n38777 = ~n38763 & ~n58369;
  assign n38778 = ~n38762 & ~n38777;
  assign n38779 = ~n38541 & n38778;
  assign n38780 = n24338 & n30192;
  assign n38781 = n25287 & n26313;
  assign n38782 = n24337 & n26319;
  assign n38783 = n25272 & n26316;
  assign n38784 = ~n38782 & ~n38783;
  assign n38785 = ~n38781 & n38784;
  assign n38786 = ~n38780 & n38785;
  assign n38787 = pi2  & ~n38786;
  assign n38788 = ~pi2  & n38786;
  assign n38789 = ~pi2  & ~n38786;
  assign n38790 = pi2  & n38786;
  assign n38791 = ~n38789 & ~n38790;
  assign n38792 = ~n38787 & ~n38788;
  assign n38793 = ~n38779 & ~n58370;
  assign n38794 = n38541 & ~n38778;
  assign n38795 = n38098 & ~n38100;
  assign n38796 = ~n38101 & ~n38795;
  assign n38797 = n24338 & ~n57002;
  assign n38798 = n25287 & n26310;
  assign n38799 = n24337 & n26316;
  assign n38800 = n25272 & n26313;
  assign n38801 = ~n38799 & ~n38800;
  assign n38802 = ~n38798 & n38801;
  assign n38803 = ~n38797 & n38802;
  assign n38804 = pi2  & ~n38803;
  assign n38805 = ~pi2  & n38803;
  assign n38806 = ~pi2  & ~n38803;
  assign n38807 = pi2  & n38803;
  assign n38808 = ~n38806 & ~n38807;
  assign n38809 = ~n38804 & ~n38805;
  assign n38810 = n38796 & ~n58371;
  assign n38811 = ~n38794 & ~n38810;
  assign n38812 = ~n38793 & n38811;
  assign n38813 = ~n38796 & n58371;
  assign n38814 = ~n38793 & ~n38794;
  assign n38815 = n38796 & ~n38814;
  assign n38816 = ~n38796 & n38814;
  assign n38817 = ~n58371 & ~n38816;
  assign n38818 = ~n38815 & ~n38817;
  assign n38819 = ~n38812 & ~n38813;
  assign n38820 = ~n38537 & ~n38815;
  assign n38821 = ~n38817 & n38820;
  assign n38822 = ~n38537 & n58372;
  assign n38823 = n38533 & n58372;
  assign n38824 = n38535 & ~n38823;
  assign n38825 = ~n38533 & ~n58372;
  assign n38826 = ~n38824 & ~n38825;
  assign n38827 = ~n38536 & ~n58373;
  assign n38828 = ~n38520 & n58374;
  assign n38829 = n38520 & ~n58374;
  assign n38830 = n24338 & ~n56867;
  assign n38831 = n25287 & n26304;
  assign n38832 = n24337 & n26310;
  assign n38833 = n25272 & n26307;
  assign n38834 = ~n38832 & ~n38833;
  assign n38835 = ~n38831 & n38834;
  assign n38836 = ~n24338 & n38835;
  assign n38837 = n56867 & n38835;
  assign n38838 = ~n38836 & ~n38837;
  assign n38839 = ~n38830 & n38835;
  assign n38840 = pi2  & ~n58375;
  assign n38841 = ~pi2  & n58375;
  assign n38842 = ~n38840 & ~n38841;
  assign n38843 = ~n38829 & n38842;
  assign n38844 = n58374 & n38842;
  assign n38845 = n38520 & ~n38844;
  assign n38846 = ~n58374 & ~n38842;
  assign n38847 = ~n38845 & ~n38846;
  assign n38848 = ~n38828 & ~n38843;
  assign n38849 = ~n38518 & n58376;
  assign n38850 = n38518 & ~n58376;
  assign n38851 = n24338 & n29446;
  assign n38852 = n25287 & n26301;
  assign n38853 = n24337 & n26307;
  assign n38854 = n25272 & n26304;
  assign n38855 = ~n38853 & ~n38854;
  assign n38856 = ~n38852 & n38855;
  assign n38857 = ~n24338 & n38856;
  assign n38858 = ~n29446 & n38856;
  assign n38859 = ~n38857 & ~n38858;
  assign n38860 = ~n38851 & n38856;
  assign n38861 = pi2  & ~n58377;
  assign n38862 = ~pi2  & n58377;
  assign n38863 = ~n38861 & ~n38862;
  assign n38864 = ~n38850 & n38863;
  assign n38865 = n58376 & n38863;
  assign n38866 = n38518 & ~n38865;
  assign n38867 = ~n58376 & ~n38863;
  assign n38868 = ~n38866 & ~n38867;
  assign n38869 = ~n38849 & ~n38864;
  assign n38870 = n38516 & ~n58378;
  assign n38871 = ~n38516 & n58378;
  assign n38872 = n24338 & ~n56870;
  assign n38873 = n25287 & n26298;
  assign n38874 = n24337 & n26304;
  assign n38875 = n25272 & n26301;
  assign n38876 = ~n38874 & ~n38875;
  assign n38877 = ~n38873 & n38876;
  assign n38878 = ~n38872 & n38877;
  assign n38879 = pi2  & ~n38878;
  assign n38880 = ~pi2  & n38878;
  assign n38881 = ~pi2  & ~n38878;
  assign n38882 = pi2  & n38878;
  assign n38883 = ~n38881 & ~n38882;
  assign n38884 = ~n38879 & ~n38880;
  assign n38885 = ~n38871 & ~n58379;
  assign n38886 = ~n38870 & ~n38885;
  assign n38887 = ~n38512 & n38886;
  assign n38888 = n24338 & n28493;
  assign n38889 = n25287 & n26295;
  assign n38890 = n24337 & n26301;
  assign n38891 = n25272 & n26298;
  assign n38892 = ~n38890 & ~n38891;
  assign n38893 = ~n38889 & n38892;
  assign n38894 = ~n38888 & n38893;
  assign n38895 = pi2  & ~n38894;
  assign n38896 = ~pi2  & n38894;
  assign n38897 = ~pi2  & ~n38894;
  assign n38898 = pi2  & n38894;
  assign n38899 = ~n38897 & ~n38898;
  assign n38900 = ~n38895 & ~n38896;
  assign n38901 = ~n38887 & ~n58380;
  assign n38902 = n38512 & ~n38886;
  assign n38903 = n38145 & ~n38147;
  assign n38904 = ~n38148 & ~n38903;
  assign n38905 = n24338 & n28808;
  assign n38906 = n25287 & n26292;
  assign n38907 = n24337 & n26298;
  assign n38908 = n25272 & n26295;
  assign n38909 = ~n38907 & ~n38908;
  assign n38910 = ~n38906 & n38909;
  assign n38911 = ~n38905 & n38910;
  assign n38912 = pi2  & ~n38911;
  assign n38913 = ~pi2  & n38911;
  assign n38914 = ~pi2  & ~n38911;
  assign n38915 = pi2  & n38911;
  assign n38916 = ~n38914 & ~n38915;
  assign n38917 = ~n38912 & ~n38913;
  assign n38918 = n38904 & ~n58381;
  assign n38919 = ~n38902 & ~n38918;
  assign n38920 = ~n38901 & n38919;
  assign n38921 = ~n38904 & n58381;
  assign n38922 = ~n38901 & ~n38902;
  assign n38923 = n38904 & ~n38922;
  assign n38924 = ~n38904 & n38922;
  assign n38925 = ~n58381 & ~n38924;
  assign n38926 = ~n38923 & ~n38925;
  assign n38927 = ~n38920 & ~n38921;
  assign n38928 = ~n38508 & ~n38923;
  assign n38929 = ~n38925 & n38928;
  assign n38930 = ~n38508 & n58382;
  assign n38931 = n38504 & n58382;
  assign n38932 = n38506 & ~n38931;
  assign n38933 = ~n38504 & ~n58382;
  assign n38934 = ~n38932 & ~n38933;
  assign n38935 = ~n38507 & ~n58383;
  assign n38936 = ~n38491 & n58384;
  assign n38937 = n38491 & ~n58384;
  assign n38938 = n24338 & ~n56721;
  assign n38939 = n25287 & n26286;
  assign n38940 = n24337 & n26292;
  assign n38941 = n25272 & n26289;
  assign n38942 = ~n38940 & ~n38941;
  assign n38943 = ~n38939 & n38942;
  assign n38944 = ~n24338 & n38943;
  assign n38945 = n56721 & n38943;
  assign n38946 = ~n38944 & ~n38945;
  assign n38947 = ~n38938 & n38943;
  assign n38948 = pi2  & ~n58385;
  assign n38949 = ~pi2  & n58385;
  assign n38950 = ~n38948 & ~n38949;
  assign n38951 = ~n38937 & n38950;
  assign n38952 = n58384 & n38950;
  assign n38953 = n38491 & ~n38952;
  assign n38954 = ~n58384 & ~n38950;
  assign n38955 = ~n38953 & ~n38954;
  assign n38956 = ~n38936 & ~n38951;
  assign n38957 = ~n38489 & n58386;
  assign n38958 = n38489 & ~n58386;
  assign n38959 = n24338 & ~n56686;
  assign n38960 = n25287 & n26283;
  assign n38961 = n24337 & n26289;
  assign n38962 = n25272 & n26286;
  assign n38963 = ~n38961 & ~n38962;
  assign n38964 = ~n38960 & n38963;
  assign n38965 = ~n24338 & n38964;
  assign n38966 = n56686 & n38964;
  assign n38967 = ~n38965 & ~n38966;
  assign n38968 = ~n38959 & n38964;
  assign n38969 = pi2  & ~n58387;
  assign n38970 = ~pi2  & n58387;
  assign n38971 = ~n38969 & ~n38970;
  assign n38972 = ~n38958 & n38971;
  assign n38973 = n58386 & n38971;
  assign n38974 = n38489 & ~n38973;
  assign n38975 = ~n58386 & ~n38971;
  assign n38976 = ~n38974 & ~n38975;
  assign n38977 = ~n38957 & ~n38972;
  assign n38978 = n38487 & ~n58388;
  assign n38979 = ~n38487 & n58388;
  assign n38980 = n24338 & n27743;
  assign n38981 = n25287 & n26280;
  assign n38982 = n24337 & n26286;
  assign n38983 = n25272 & n26283;
  assign n38984 = ~n38982 & ~n38983;
  assign n38985 = ~n38981 & n38984;
  assign n38986 = ~n38980 & n38985;
  assign n38987 = pi2  & ~n38986;
  assign n38988 = ~pi2  & n38986;
  assign n38989 = ~pi2  & ~n38986;
  assign n38990 = pi2  & n38986;
  assign n38991 = ~n38989 & ~n38990;
  assign n38992 = ~n38987 & ~n38988;
  assign n38993 = ~n38979 & ~n58389;
  assign n38994 = ~n38978 & ~n38993;
  assign n38995 = ~n38483 & n38994;
  assign n38996 = n24338 & n27330;
  assign n38997 = n25287 & n26277;
  assign n38998 = n24337 & n26283;
  assign n38999 = n25272 & n26280;
  assign n39000 = ~n38998 & ~n38999;
  assign n39001 = ~n38997 & n39000;
  assign n39002 = ~n38996 & n39001;
  assign n39003 = pi2  & ~n39002;
  assign n39004 = ~pi2  & n39002;
  assign n39005 = ~pi2  & ~n39002;
  assign n39006 = pi2  & n39002;
  assign n39007 = ~n39005 & ~n39006;
  assign n39008 = ~n39003 & ~n39004;
  assign n39009 = ~n38995 & ~n58390;
  assign n39010 = n38483 & ~n38994;
  assign n39011 = n38192 & ~n38194;
  assign n39012 = ~n38195 & ~n39011;
  assign n39013 = n24338 & ~n56648;
  assign n39014 = n25287 & n26274;
  assign n39015 = n24337 & n26280;
  assign n39016 = n25272 & n26277;
  assign n39017 = ~n39015 & ~n39016;
  assign n39018 = ~n39014 & n39017;
  assign n39019 = ~n39013 & n39018;
  assign n39020 = pi2  & ~n39019;
  assign n39021 = ~pi2  & n39019;
  assign n39022 = ~pi2  & ~n39019;
  assign n39023 = pi2  & n39019;
  assign n39024 = ~n39022 & ~n39023;
  assign n39025 = ~n39020 & ~n39021;
  assign n39026 = n39012 & ~n58391;
  assign n39027 = ~n39010 & ~n39026;
  assign n39028 = ~n39009 & n39027;
  assign n39029 = ~n39012 & n58391;
  assign n39030 = ~n39009 & ~n39010;
  assign n39031 = n39012 & ~n39030;
  assign n39032 = ~n39012 & n39030;
  assign n39033 = ~n58391 & ~n39032;
  assign n39034 = ~n39031 & ~n39033;
  assign n39035 = ~n39028 & ~n39029;
  assign n39036 = ~n38479 & ~n39031;
  assign n39037 = ~n39033 & n39036;
  assign n39038 = ~n38479 & n58392;
  assign n39039 = n38475 & n58392;
  assign n39040 = n38477 & ~n39039;
  assign n39041 = ~n38475 & ~n58392;
  assign n39042 = ~n39040 & ~n39041;
  assign n39043 = ~n38478 & ~n58393;
  assign n39044 = ~n38462 & n58394;
  assign n39045 = n38462 & ~n58394;
  assign n39046 = n24338 & ~n56601;
  assign n39047 = n25287 & n26268;
  assign n39048 = n24337 & n26274;
  assign n39049 = n25272 & n26271;
  assign n39050 = ~n39048 & ~n39049;
  assign n39051 = ~n39047 & n39050;
  assign n39052 = ~n24338 & n39051;
  assign n39053 = n56601 & n39051;
  assign n39054 = ~n39052 & ~n39053;
  assign n39055 = ~n39046 & n39051;
  assign n39056 = pi2  & ~n58395;
  assign n39057 = ~pi2  & n58395;
  assign n39058 = ~n39056 & ~n39057;
  assign n39059 = ~n39045 & n39058;
  assign n39060 = n58394 & n39058;
  assign n39061 = n38462 & ~n39060;
  assign n39062 = ~n58394 & ~n39058;
  assign n39063 = ~n39061 & ~n39062;
  assign n39064 = ~n39044 & ~n39059;
  assign n39065 = ~n38460 & n58396;
  assign n39066 = n38460 & ~n58396;
  assign n39067 = n24338 & n27042;
  assign n39068 = n25287 & n26265;
  assign n39069 = n24337 & n26271;
  assign n39070 = n25272 & n26268;
  assign n39071 = ~n39069 & ~n39070;
  assign n39072 = ~n39068 & n39071;
  assign n39073 = ~n24338 & n39072;
  assign n39074 = ~n27042 & n39072;
  assign n39075 = ~n39073 & ~n39074;
  assign n39076 = ~n39067 & n39072;
  assign n39077 = pi2  & ~n58397;
  assign n39078 = ~pi2  & n58397;
  assign n39079 = ~n39077 & ~n39078;
  assign n39080 = ~n39066 & n39079;
  assign n39081 = n58396 & n39079;
  assign n39082 = n38460 & ~n39081;
  assign n39083 = ~n58396 & ~n39079;
  assign n39084 = ~n39082 & ~n39083;
  assign n39085 = ~n39065 & ~n39080;
  assign n39086 = n38458 & ~n58398;
  assign n39087 = ~n38458 & n58398;
  assign n39088 = n24338 & n27466;
  assign n39089 = n25287 & n26262;
  assign n39090 = n24337 & n26268;
  assign n39091 = n25272 & n26265;
  assign n39092 = ~n39090 & ~n39091;
  assign n39093 = ~n39089 & n39092;
  assign n39094 = ~n39088 & n39093;
  assign n39095 = pi2  & ~n39094;
  assign n39096 = ~pi2  & n39094;
  assign n39097 = ~pi2  & ~n39094;
  assign n39098 = pi2  & n39094;
  assign n39099 = ~n39097 & ~n39098;
  assign n39100 = ~n39095 & ~n39096;
  assign n39101 = ~n39087 & ~n58399;
  assign n39102 = ~n39086 & ~n39101;
  assign n39103 = n38454 & ~n39102;
  assign n39104 = ~n38454 & n39102;
  assign n39105 = n24338 & ~n56639;
  assign n39106 = n25287 & n26259;
  assign n39107 = n24337 & n26265;
  assign n39108 = n25272 & n26262;
  assign n39109 = ~n39107 & ~n39108;
  assign n39110 = ~n39106 & n39109;
  assign n39111 = ~n39105 & n39110;
  assign n39112 = pi2  & ~n39111;
  assign n39113 = ~pi2  & n39111;
  assign n39114 = ~pi2  & ~n39111;
  assign n39115 = pi2  & n39111;
  assign n39116 = ~n39114 & ~n39115;
  assign n39117 = ~n39112 & ~n39113;
  assign n39118 = ~n39104 & ~n58400;
  assign n39119 = ~n39103 & ~n39118;
  assign n39120 = ~n58339 & ~n39119;
  assign n39121 = ~n38445 & ~n39120;
  assign n39122 = ~n38415 & n38428;
  assign n39123 = ~n38429 & ~n39122;
  assign n39124 = ~n39121 & n39123;
  assign n39125 = ~n38429 & ~n39124;
  assign n39126 = ~n38399 & n38412;
  assign n39127 = ~n38413 & ~n39126;
  assign n39128 = ~n39125 & n39127;
  assign n39129 = ~n38413 & ~n39128;
  assign n39130 = ~n38383 & n38396;
  assign n39131 = ~n38397 & ~n39130;
  assign n39132 = ~n39129 & n39131;
  assign n39133 = ~n38397 & ~n39132;
  assign n39134 = ~n38367 & n38380;
  assign n39135 = ~n38381 & ~n39134;
  assign n39136 = ~n39133 & n39135;
  assign n39137 = ~n38381 & ~n39136;
  assign n39138 = ~n38351 & n38364;
  assign n39139 = ~n38365 & ~n39138;
  assign n39140 = ~n39137 & n39139;
  assign n39141 = ~n38365 & ~n39140;
  assign n39142 = ~n38335 & n38348;
  assign n39143 = ~n38349 & ~n39142;
  assign n39144 = ~n39141 & n39143;
  assign n39145 = ~n38349 & ~n39144;
  assign n39146 = ~n38318 & n38332;
  assign n39147 = ~n38333 & ~n39146;
  assign n39148 = ~n39145 & n39147;
  assign n39149 = ~n38333 & ~n39148;
  assign n39150 = ~n38313 & n38315;
  assign n39151 = ~n38316 & ~n39150;
  assign n39152 = ~n39149 & n39151;
  assign n39153 = ~n38316 & ~n39152;
  assign n39154 = n38311 & ~n39153;
  assign n39155 = ~n38309 & ~n39154;
  assign n39156 = n37401 & ~n39155;
  assign n39157 = ~n37399 & ~n39156;
  assign n39158 = n37366 & ~n39157;
  assign n39159 = ~n37364 & ~n39158;
  assign n39160 = n36510 & ~n39159;
  assign n39161 = ~n36508 & ~n39160;
  assign n39162 = ~n34940 & n57869;
  assign n39163 = ~n35674 & ~n39162;
  assign n39164 = ~n39161 & n39163;
  assign n39165 = ~n35674 & ~n39164;
  assign n39166 = n34932 & n57753;
  assign n39167 = ~n57753 & ~n34938;
  assign n39168 = n34932 & ~n57753;
  assign n39169 = ~n34932 & ~n34938;
  assign n39170 = ~n34932 & n57753;
  assign n39171 = ~n58401 & ~n58402;
  assign n39172 = ~n34938 & ~n39166;
  assign n39173 = ~n39165 & ~n58403;
  assign n39174 = ~n34938 & ~n39173;
  assign n39175 = n34204 & ~n39174;
  assign n39176 = ~n34202 & ~n39175;
  assign n39177 = ~n32935 & n57514;
  assign n39178 = ~n33549 & ~n39177;
  assign n39179 = ~n39176 & n39178;
  assign n39180 = ~n33549 & ~n39179;
  assign n39181 = n32925 & ~n57402;
  assign n39182 = n57402 & ~n32933;
  assign n39183 = n32925 & n57402;
  assign n39184 = ~n32925 & ~n32933;
  assign n39185 = ~n32925 & ~n57402;
  assign n39186 = ~n58404 & ~n58405;
  assign n39187 = ~n32933 & ~n39181;
  assign n39188 = ~n39180 & ~n58406;
  assign n39189 = ~n32933 & ~n39188;
  assign n39190 = n32352 & ~n39189;
  assign n39191 = ~n32350 & ~n39190;
  assign n39192 = ~n31633 & n57217;
  assign n39193 = ~n31842 & ~n39192;
  assign n39194 = ~n39191 & n39193;
  assign n39195 = ~n31842 & ~n39194;
  assign n39196 = n31625 & n57175;
  assign n39197 = ~n57175 & ~n31631;
  assign n39198 = n31625 & ~n57175;
  assign n39199 = ~n31625 & ~n31631;
  assign n39200 = ~n31625 & n57175;
  assign n39201 = ~n58407 & ~n58408;
  assign n39202 = ~n31631 & ~n39196;
  assign n39203 = ~n39195 & ~n58409;
  assign n39204 = ~n31631 & ~n39203;
  assign n39205 = n31408 & ~n39204;
  assign n39206 = ~n31406 & ~n39205;
  assign n39207 = ~n29926 & n56985;
  assign n39208 = ~n30102 & ~n39207;
  assign n39209 = ~n39206 & n39208;
  assign n39210 = ~n30102 & ~n39209;
  assign n39211 = n29916 & ~n56954;
  assign n39212 = n56954 & ~n29924;
  assign n39213 = n29916 & n56954;
  assign n39214 = ~n29916 & ~n29924;
  assign n39215 = ~n29916 & ~n56954;
  assign n39216 = ~n58410 & ~n58411;
  assign n39217 = ~n29924 & ~n39211;
  assign n39218 = ~n39210 & ~n58412;
  assign n39219 = ~n29924 & ~n39218;
  assign n39220 = n29373 & ~n39219;
  assign n39221 = ~n29371 & ~n39220;
  assign n39222 = ~n28771 & n56835;
  assign n39223 = ~n28950 & ~n39222;
  assign n39224 = ~n39221 & n39223;
  assign n39225 = ~n28950 & ~n39224;
  assign n39226 = n28763 & n56803;
  assign n39227 = ~n56803 & ~n28769;
  assign n39228 = n28763 & ~n56803;
  assign n39229 = ~n28763 & ~n28769;
  assign n39230 = ~n28763 & n56803;
  assign n39231 = ~n58413 & ~n58414;
  assign n39232 = ~n28769 & ~n39226;
  assign n39233 = ~n39225 & ~n58415;
  assign n39234 = ~n28769 & ~n39233;
  assign n39235 = n28623 & ~n39234;
  assign n39236 = ~n28621 & ~n39235;
  assign n39237 = ~n27401 & ~n27409;
  assign n39238 = n123 & n27839;
  assign n39239 = n128 & n26244;
  assign n39240 = n53444 & n26250;
  assign n39241 = n127 & n26247;
  assign n39242 = ~n39240 & ~n39241;
  assign n39243 = ~n39239 & n39242;
  assign n39244 = ~n39238 & n39243;
  assign n39245 = pi26  & ~n39244;
  assign n39246 = pi26  & ~n39245;
  assign n39247 = pi26  & n39244;
  assign n39248 = ~n39244 & ~n39245;
  assign n39249 = ~pi26  & ~n39244;
  assign n39250 = ~n58416 & ~n58417;
  assign n39251 = n11279 & ~n56668;
  assign n39252 = n12584 & n26253;
  assign n39253 = n54410 & n26259;
  assign n39254 = n11267 & n26256;
  assign n39255 = ~n39253 & ~n39254;
  assign n39256 = ~n39252 & n39255;
  assign n39257 = ~n39251 & n39256;
  assign n39258 = pi29  & ~n39257;
  assign n39259 = pi29  & ~n39258;
  assign n39260 = pi29  & n39257;
  assign n39261 = ~n39257 & ~n39258;
  assign n39262 = ~pi29  & ~n39257;
  assign n39263 = ~n58418 & ~n58419;
  assign n39264 = ~n27059 & ~n27383;
  assign n39265 = n1576 & n27466;
  assign n39266 = n11215 & n26262;
  assign n39267 = n54403 & n26268;
  assign n39268 = n10564 & n26265;
  assign n39269 = ~n39267 & ~n39268;
  assign n39270 = ~n39266 & n39269;
  assign n39271 = ~n39265 & n39270;
  assign n39272 = n7755 & n14965;
  assign n39273 = n27169 & n39272;
  assign n39274 = n53702 & n39273;
  assign n39275 = n54278 & n39274;
  assign n39276 = n905 & n4313;
  assign n39277 = ~n983 & ~n1912;
  assign n39278 = ~n1192 & ~n1912;
  assign n39279 = ~n983 & n39278;
  assign n39280 = ~n1192 & n39277;
  assign n39281 = n4224 & n4376;
  assign n39282 = n58420 & n39281;
  assign n39283 = n39276 & n39282;
  assign n39284 = n54002 & n39283;
  assign n39285 = n4224 & n7755;
  assign n39286 = n14965 & n39285;
  assign n39287 = n54278 & n39286;
  assign n39288 = n4224 & n14965;
  assign n39289 = n54278 & n39288;
  assign n39290 = n53702 & n39289;
  assign n39291 = n7755 & n39290;
  assign n39292 = n53702 & n39287;
  assign n39293 = n54002 & n58421;
  assign n39294 = n4313 & n39293;
  assign n39295 = n4376 & n39294;
  assign n39296 = n905 & n39295;
  assign n39297 = ~n416 & n39296;
  assign n39298 = ~n1192 & n39297;
  assign n39299 = ~n983 & n39298;
  assign n39300 = ~n465 & n39299;
  assign n39301 = ~n1912 & n39300;
  assign n39302 = n905 & n27169;
  assign n39303 = n4313 & n4376;
  assign n39304 = n39302 & n39303;
  assign n39305 = n58420 & n39304;
  assign n39306 = n54002 & n39305;
  assign n39307 = n58421 & n39306;
  assign n39308 = n39275 & n39284;
  assign n39309 = n5116 & n5377;
  assign n39310 = n11514 & n39309;
  assign n39311 = ~n346 & ~n623;
  assign n39312 = n1704 & n39311;
  assign n39313 = n4538 & n4914;
  assign n39314 = n39312 & n39313;
  assign n39315 = ~n363 & ~n773;
  assign n39316 = ~n901 & n39315;
  assign n39317 = n12339 & n39316;
  assign n39318 = ~n346 & ~n363;
  assign n39319 = n4538 & n39318;
  assign n39320 = n1704 & n4914;
  assign n39321 = n39319 & n39320;
  assign n39322 = ~n623 & ~n773;
  assign n39323 = ~n901 & n39322;
  assign n39324 = n12339 & n39323;
  assign n39325 = n39321 & n39324;
  assign n39326 = n39314 & n39317;
  assign n39327 = n4914 & n5377;
  assign n39328 = n11514 & n39327;
  assign n39329 = n1704 & n4538;
  assign n39330 = n5116 & n39315;
  assign n39331 = n39329 & n39330;
  assign n39332 = ~n901 & n39311;
  assign n39333 = n12339 & n39332;
  assign n39334 = n39331 & n39333;
  assign n39335 = n39328 & n39334;
  assign n39336 = n4914 & n5116;
  assign n39337 = n5377 & n39336;
  assign n39338 = ~n363 & ~n901;
  assign n39339 = n39322 & n39338;
  assign n39340 = n39329 & n39339;
  assign n39341 = ~n346 & ~n789;
  assign n39342 = ~n2103 & n39341;
  assign n39343 = n12339 & n39342;
  assign n39344 = n39340 & n39343;
  assign n39345 = n39337 & n39344;
  assign n39346 = n39310 & n58423;
  assign n39347 = n53911 & n54320;
  assign n39348 = n58424 & n39347;
  assign n39349 = n58422 & n39348;
  assign n39350 = n4914 & n12339;
  assign n39351 = n54320 & n39350;
  assign n39352 = n53911 & n39351;
  assign n39353 = n5116 & n39352;
  assign n39354 = n58422 & n39353;
  assign n39355 = n54082 & n39354;
  assign n39356 = n1704 & n39355;
  assign n39357 = n4538 & n39356;
  assign n39358 = n5377 & n39357;
  assign n39359 = ~n2103 & n39358;
  assign n39360 = ~n901 & n39359;
  assign n39361 = ~n363 & n39360;
  assign n39362 = ~n773 & n39361;
  assign n39363 = ~n789 & n39362;
  assign n39364 = ~n346 & n39363;
  assign n39365 = ~n623 & n39364;
  assign n39366 = n54082 & n39349;
  assign n39367 = ~n56589 & ~n58425;
  assign n39368 = n56589 & n58425;
  assign n39369 = ~n39367 & ~n39368;
  assign n39370 = n27531 & n39369;
  assign n39371 = ~n27531 & ~n39369;
  assign n39372 = ~n39370 & ~n39371;
  assign n39373 = n27055 & ~n39372;
  assign n39374 = ~n27055 & n39372;
  assign n39375 = ~n39373 & ~n39374;
  assign n39376 = ~n39271 & n39375;
  assign n39377 = n39271 & ~n39375;
  assign n39378 = n39375 & ~n39376;
  assign n39379 = ~n39271 & ~n39376;
  assign n39380 = ~n39378 & ~n39379;
  assign n39381 = ~n39376 & ~n39377;
  assign n39382 = ~n39264 & ~n58426;
  assign n39383 = n39264 & n58426;
  assign n39384 = ~n39382 & ~n39383;
  assign n39385 = ~n39263 & n39384;
  assign n39386 = n39384 & ~n39385;
  assign n39387 = n39263 & n39384;
  assign n39388 = ~n39263 & ~n39385;
  assign n39389 = ~n39263 & ~n39384;
  assign n39390 = n39263 & ~n39384;
  assign n39391 = ~n39385 & ~n39390;
  assign n39392 = ~n58427 & ~n58428;
  assign n39393 = ~n39250 & n58429;
  assign n39394 = n39250 & ~n58429;
  assign n39395 = n58429 & ~n39393;
  assign n39396 = n39250 & n58429;
  assign n39397 = ~n39250 & ~n39393;
  assign n39398 = ~n39250 & ~n58429;
  assign n39399 = ~n58430 & ~n58431;
  assign n39400 = ~n39393 & ~n39394;
  assign n39401 = ~n39237 & ~n58432;
  assign n39402 = n39237 & n58432;
  assign n39403 = ~n39401 & ~n39402;
  assign n39404 = n90 & n28624;
  assign n39405 = n14210 & ~n26537;
  assign n39406 = n54667 & n26242;
  assign n39407 = ~n14236 & ~n39406;
  assign n39408 = ~n39405 & ~n39406;
  assign n39409 = ~n14236 & n39408;
  assign n39410 = ~n39405 & n39407;
  assign n39411 = ~n39404 & n58433;
  assign n39412 = pi23  & ~n39411;
  assign n39413 = pi23  & ~n39412;
  assign n39414 = pi23  & n39411;
  assign n39415 = ~n39411 & ~n39412;
  assign n39416 = ~pi23  & ~n39411;
  assign n39417 = ~n58434 & ~n58435;
  assign n39418 = ~n26557 & ~n27512;
  assign n39419 = ~n27511 & ~n27514;
  assign n39420 = ~n27511 & ~n39418;
  assign n39421 = ~n39417 & ~n58436;
  assign n39422 = n39417 & n58436;
  assign n39423 = ~n58436 & ~n39421;
  assign n39424 = n39417 & ~n58436;
  assign n39425 = ~n39417 & ~n39421;
  assign n39426 = ~n39417 & n58436;
  assign n39427 = ~n58437 & ~n58438;
  assign n39428 = ~n39421 & ~n39422;
  assign n39429 = n39403 & ~n58439;
  assign n39430 = ~n39403 & n58439;
  assign n39431 = ~n39429 & ~n39430;
  assign n39432 = n56665 & ~n27828;
  assign n39433 = ~n27827 & ~n27830;
  assign n39434 = ~n27827 & ~n39432;
  assign n39435 = n39431 & ~n58440;
  assign n39436 = ~n39431 & n58440;
  assign n39437 = ~n39435 & ~n39436;
  assign n39438 = ~n39236 & n39437;
  assign n39439 = n39236 & ~n39437;
  assign n39440 = ~n39438 & ~n39439;
  assign n39441 = ~n39435 & ~n39438;
  assign n39442 = ~n39421 & ~n39429;
  assign n39443 = n54667 & ~n26537;
  assign n39444 = ~n14210 & ~n14236;
  assign n39445 = ~n14210 & ~n39443;
  assign n39446 = ~n14236 & n39445;
  assign n39447 = ~n14236 & ~n39443;
  assign n39448 = ~n14210 & n39447;
  assign n39449 = ~n39443 & n39444;
  assign n39450 = ~n90 & n58441;
  assign n39451 = pi23  & ~n39450;
  assign n39452 = pi23  & ~n39451;
  assign n39453 = pi23  & n39450;
  assign n39454 = ~n39450 & ~n39451;
  assign n39455 = ~pi23  & ~n39450;
  assign n39456 = ~n58442 & ~n58443;
  assign n39457 = ~n39393 & ~n39401;
  assign n39458 = n123 & n27808;
  assign n39459 = n128 & n26242;
  assign n39460 = n53444 & n26247;
  assign n39461 = n127 & n26244;
  assign n39462 = ~n39460 & ~n39461;
  assign n39463 = ~n39459 & n39462;
  assign n39464 = ~n39458 & n39463;
  assign n39465 = pi26  & ~n39464;
  assign n39466 = pi26  & ~n39465;
  assign n39467 = pi26  & n39464;
  assign n39468 = ~n39464 & ~n39465;
  assign n39469 = ~pi26  & ~n39464;
  assign n39470 = ~n58444 & ~n58445;
  assign n39471 = ~n39367 & ~n39370;
  assign n39472 = n53600 & ~n39471;
  assign n39473 = ~n53600 & n39471;
  assign n39474 = ~n39472 & ~n39473;
  assign n39475 = n1576 & ~n56639;
  assign n39476 = n11215 & n26259;
  assign n39477 = n10564 & n26262;
  assign n39478 = n54403 & n26265;
  assign n39479 = ~n39477 & ~n39478;
  assign n39480 = ~n39476 & n39479;
  assign n39481 = ~n39475 & ~n39478;
  assign n39482 = ~n39477 & n39481;
  assign n39483 = ~n39476 & n39482;
  assign n39484 = ~n39475 & n39480;
  assign n39485 = n39474 & ~n58446;
  assign n39486 = ~n39474 & n58446;
  assign n39487 = ~n39485 & ~n39486;
  assign n39488 = n39271 & ~n39374;
  assign n39489 = ~n39374 & ~n39376;
  assign n39490 = ~n39373 & ~n39488;
  assign n39491 = n39487 & ~n58447;
  assign n39492 = ~n39487 & n58447;
  assign n39493 = ~n39491 & ~n39492;
  assign n39494 = n11279 & n27491;
  assign n39495 = n12584 & n26250;
  assign n39496 = n54410 & n26256;
  assign n39497 = n11267 & n26253;
  assign n39498 = ~n39496 & ~n39497;
  assign n39499 = ~n39495 & n39498;
  assign n39500 = ~n11279 & n39499;
  assign n39501 = ~n27491 & n39499;
  assign n39502 = ~n39500 & ~n39501;
  assign n39503 = ~n39494 & n39499;
  assign n39504 = pi29  & ~n58448;
  assign n39505 = ~pi29  & n58448;
  assign n39506 = ~n39504 & ~n39505;
  assign n39507 = n39493 & ~n39506;
  assign n39508 = ~n39493 & n39506;
  assign n39509 = ~n39507 & ~n39508;
  assign n39510 = ~n39263 & ~n39383;
  assign n39511 = ~n39382 & ~n39385;
  assign n39512 = ~n39382 & ~n39510;
  assign n39513 = n39509 & ~n58449;
  assign n39514 = ~n39509 & n58449;
  assign n39515 = ~n39513 & ~n39514;
  assign n39516 = ~n39470 & n39515;
  assign n39517 = n39515 & ~n39516;
  assign n39518 = n39470 & n39515;
  assign n39519 = ~n39470 & ~n39516;
  assign n39520 = ~n39470 & ~n39515;
  assign n39521 = n39470 & ~n39515;
  assign n39522 = ~n39516 & ~n39521;
  assign n39523 = ~n58450 & ~n58451;
  assign n39524 = n39457 & ~n58452;
  assign n39525 = ~n39457 & n58452;
  assign n39526 = ~n39524 & ~n39525;
  assign n39527 = n39456 & ~n39526;
  assign n39528 = ~n39456 & n39526;
  assign n39529 = n39526 & ~n39528;
  assign n39530 = n39456 & n39526;
  assign n39531 = ~n39456 & ~n39528;
  assign n39532 = ~n39456 & ~n39526;
  assign n39533 = ~n58453 & ~n58454;
  assign n39534 = ~n39527 & ~n39528;
  assign n39535 = ~n39442 & ~n58455;
  assign n39536 = n39442 & n58455;
  assign n39537 = ~n58455 & ~n39535;
  assign n39538 = ~n39442 & ~n39535;
  assign n39539 = ~n39537 & ~n39538;
  assign n39540 = ~n39535 & ~n39536;
  assign n39541 = ~n39441 & ~n58456;
  assign n39542 = n39441 & n58456;
  assign n39543 = ~n39541 & ~n39542;
  assign n39544 = n39440 & n39543;
  assign n39545 = ~n28623 & n39234;
  assign n39546 = ~n39235 & ~n39545;
  assign n39547 = n39440 & n39546;
  assign n39548 = n39225 & n58415;
  assign n39549 = ~n39233 & ~n39548;
  assign n39550 = n39546 & n39549;
  assign n39551 = n39221 & ~n39223;
  assign n39552 = ~n39224 & ~n39551;
  assign n39553 = n39549 & n39552;
  assign n39554 = ~n29373 & n39219;
  assign n39555 = ~n39220 & ~n39554;
  assign n39556 = n39552 & n39555;
  assign n39557 = n39210 & n58412;
  assign n39558 = ~n39218 & ~n39557;
  assign n39559 = n39555 & n39558;
  assign n39560 = n39206 & ~n39208;
  assign n39561 = ~n39209 & ~n39560;
  assign n39562 = n39558 & n39561;
  assign n39563 = ~n31408 & n39204;
  assign n39564 = ~n39205 & ~n39563;
  assign n39565 = n39561 & n39564;
  assign n39566 = n39195 & n58409;
  assign n39567 = ~n39203 & ~n39566;
  assign n39568 = n39564 & n39567;
  assign n39569 = n39191 & ~n39193;
  assign n39570 = ~n39194 & ~n39569;
  assign n39571 = n39567 & n39570;
  assign n39572 = ~n32352 & n39189;
  assign n39573 = ~n39190 & ~n39572;
  assign n39574 = n39570 & n39573;
  assign n39575 = n39180 & n58406;
  assign n39576 = ~n39188 & ~n39575;
  assign n39577 = n39573 & n39576;
  assign n39578 = n39176 & ~n39178;
  assign n39579 = ~n39179 & ~n39578;
  assign n39580 = n39576 & n39579;
  assign n39581 = ~n34204 & n39174;
  assign n39582 = ~n39175 & ~n39581;
  assign n39583 = n39579 & n39582;
  assign n39584 = n39165 & n58403;
  assign n39585 = ~n39173 & ~n39584;
  assign n39586 = n39582 & n39585;
  assign n39587 = n39161 & ~n39163;
  assign n39588 = ~n39164 & ~n39587;
  assign n39589 = n39585 & n39588;
  assign n39590 = ~n36510 & n39159;
  assign n39591 = ~n39160 & ~n39590;
  assign n39592 = n39588 & n39591;
  assign n39593 = ~n37366 & n39157;
  assign n39594 = ~n39158 & ~n39593;
  assign n39595 = n39591 & n39594;
  assign n39596 = ~n37401 & n39155;
  assign n39597 = ~n39156 & ~n39596;
  assign n39598 = n39594 & n39597;
  assign n39599 = ~n38311 & n39153;
  assign n39600 = ~n39154 & ~n39599;
  assign n39601 = n39597 & n39600;
  assign n39602 = n39149 & ~n39151;
  assign n39603 = ~n39152 & ~n39602;
  assign n39604 = n39600 & n39603;
  assign n39605 = n39145 & ~n39147;
  assign n39606 = ~n39148 & ~n39605;
  assign n39607 = n39603 & n39606;
  assign n39608 = n39141 & ~n39143;
  assign n39609 = ~n39144 & ~n39608;
  assign n39610 = n39606 & n39609;
  assign n39611 = n39137 & ~n39139;
  assign n39612 = ~n39140 & ~n39611;
  assign n39613 = n39609 & n39612;
  assign n39614 = n39133 & ~n39135;
  assign n39615 = ~n39136 & ~n39614;
  assign n39616 = n39612 & n39615;
  assign n39617 = n39129 & ~n39131;
  assign n39618 = ~n39132 & ~n39617;
  assign n39619 = n39615 & n39618;
  assign n39620 = n39125 & ~n39127;
  assign n39621 = ~n39128 & ~n39620;
  assign n39622 = n39618 & n39621;
  assign n39623 = ~n39618 & ~n39621;
  assign n39624 = ~n39622 & ~n39623;
  assign n39625 = n39121 & ~n39123;
  assign n39626 = ~n39124 & ~n39625;
  assign n39627 = n58339 & n39119;
  assign n39628 = ~n39119 & ~n39120;
  assign n39629 = ~n58339 & ~n39120;
  assign n39630 = ~n39628 & ~n39629;
  assign n39631 = ~n39120 & ~n39627;
  assign n39632 = ~n39621 & n58457;
  assign n39633 = n39621 & n39626;
  assign n39634 = n39626 & ~n58457;
  assign n39635 = ~n39621 & n39634;
  assign n39636 = ~n39633 & ~n39635;
  assign n39637 = n39626 & ~n39632;
  assign n39638 = n39624 & ~n58458;
  assign n39639 = ~n39622 & ~n39638;
  assign n39640 = ~n39615 & ~n39618;
  assign n39641 = ~n39619 & ~n39640;
  assign n39642 = ~n39639 & n39641;
  assign n39643 = ~n39619 & ~n39642;
  assign n39644 = ~n39612 & ~n39615;
  assign n39645 = ~n39616 & ~n39644;
  assign n39646 = ~n39643 & n39645;
  assign n39647 = ~n39616 & ~n39646;
  assign n39648 = ~n39609 & ~n39612;
  assign n39649 = ~n39613 & ~n39648;
  assign n39650 = ~n39647 & n39649;
  assign n39651 = ~n39613 & ~n39650;
  assign n39652 = ~n39606 & ~n39609;
  assign n39653 = ~n39610 & ~n39652;
  assign n39654 = ~n39651 & n39653;
  assign n39655 = ~n39610 & ~n39654;
  assign n39656 = ~n39603 & ~n39606;
  assign n39657 = ~n39607 & ~n39656;
  assign n39658 = ~n39655 & n39657;
  assign n39659 = ~n39607 & ~n39658;
  assign n39660 = ~n39600 & ~n39603;
  assign n39661 = ~n39604 & ~n39660;
  assign n39662 = ~n39604 & ~n39659;
  assign n39663 = ~n39660 & n39662;
  assign n39664 = ~n39659 & n39661;
  assign n39665 = ~n39604 & ~n58459;
  assign n39666 = ~n39597 & ~n39600;
  assign n39667 = ~n39601 & ~n39666;
  assign n39668 = ~n39665 & n39667;
  assign n39669 = ~n39601 & ~n39668;
  assign n39670 = ~n39594 & ~n39597;
  assign n39671 = ~n39598 & ~n39670;
  assign n39672 = ~n39669 & n39671;
  assign n39673 = ~n39598 & ~n39672;
  assign n39674 = ~n39591 & ~n39594;
  assign n39675 = ~n39595 & ~n39674;
  assign n39676 = ~n39673 & n39675;
  assign n39677 = ~n39595 & ~n39676;
  assign n39678 = ~n39588 & ~n39591;
  assign n39679 = ~n39592 & ~n39678;
  assign n39680 = ~n39677 & ~n39678;
  assign n39681 = ~n39592 & n39680;
  assign n39682 = ~n39677 & n39679;
  assign n39683 = ~n39592 & ~n58460;
  assign n39684 = ~n39585 & ~n39588;
  assign n39685 = ~n39589 & ~n39684;
  assign n39686 = ~n39683 & ~n39684;
  assign n39687 = ~n39589 & n39686;
  assign n39688 = ~n39683 & n39685;
  assign n39689 = ~n39589 & ~n58461;
  assign n39690 = ~n39582 & ~n39585;
  assign n39691 = ~n39586 & ~n39690;
  assign n39692 = ~n39689 & n39691;
  assign n39693 = ~n39586 & ~n39692;
  assign n39694 = ~n39579 & ~n39582;
  assign n39695 = ~n39583 & ~n39694;
  assign n39696 = ~n39693 & ~n39694;
  assign n39697 = ~n39583 & n39696;
  assign n39698 = ~n39693 & n39695;
  assign n39699 = ~n39583 & ~n58462;
  assign n39700 = ~n39576 & ~n39579;
  assign n39701 = ~n39580 & ~n39700;
  assign n39702 = ~n39699 & ~n39700;
  assign n39703 = ~n39580 & n39702;
  assign n39704 = ~n39699 & n39701;
  assign n39705 = ~n39580 & ~n58463;
  assign n39706 = ~n39573 & ~n39576;
  assign n39707 = ~n39577 & ~n39706;
  assign n39708 = ~n39705 & n39707;
  assign n39709 = ~n39577 & ~n39708;
  assign n39710 = ~n39570 & ~n39573;
  assign n39711 = ~n39574 & ~n39710;
  assign n39712 = ~n39709 & ~n39710;
  assign n39713 = ~n39574 & n39712;
  assign n39714 = ~n39709 & n39711;
  assign n39715 = ~n39574 & ~n58464;
  assign n39716 = ~n39567 & ~n39570;
  assign n39717 = ~n39571 & ~n39716;
  assign n39718 = ~n39715 & ~n39716;
  assign n39719 = ~n39571 & n39718;
  assign n39720 = ~n39715 & n39717;
  assign n39721 = ~n39571 & ~n58465;
  assign n39722 = ~n39564 & ~n39567;
  assign n39723 = ~n39568 & ~n39722;
  assign n39724 = ~n39721 & n39723;
  assign n39725 = ~n39568 & ~n39724;
  assign n39726 = ~n39561 & ~n39564;
  assign n39727 = ~n39565 & ~n39726;
  assign n39728 = ~n39725 & ~n39726;
  assign n39729 = ~n39565 & n39728;
  assign n39730 = ~n39725 & n39727;
  assign n39731 = ~n39565 & ~n58466;
  assign n39732 = ~n39558 & ~n39561;
  assign n39733 = ~n39562 & ~n39732;
  assign n39734 = ~n39731 & ~n39732;
  assign n39735 = ~n39562 & n39734;
  assign n39736 = ~n39731 & n39733;
  assign n39737 = ~n39562 & ~n58467;
  assign n39738 = ~n39555 & ~n39558;
  assign n39739 = ~n39559 & ~n39738;
  assign n39740 = ~n39737 & n39739;
  assign n39741 = ~n39559 & ~n39740;
  assign n39742 = ~n39552 & ~n39555;
  assign n39743 = ~n39556 & ~n39742;
  assign n39744 = ~n39741 & ~n39742;
  assign n39745 = ~n39556 & n39744;
  assign n39746 = ~n39741 & n39743;
  assign n39747 = ~n39556 & ~n58468;
  assign n39748 = ~n39549 & ~n39552;
  assign n39749 = ~n39553 & ~n39748;
  assign n39750 = ~n39747 & ~n39748;
  assign n39751 = ~n39553 & n39750;
  assign n39752 = ~n39747 & n39749;
  assign n39753 = ~n39553 & ~n58469;
  assign n39754 = ~n39546 & ~n39549;
  assign n39755 = ~n39550 & ~n39754;
  assign n39756 = ~n39753 & n39755;
  assign n39757 = ~n39550 & ~n39756;
  assign n39758 = ~n39440 & ~n39546;
  assign n39759 = ~n39547 & ~n39758;
  assign n39760 = ~n39757 & ~n39758;
  assign n39761 = ~n39547 & n39760;
  assign n39762 = ~n39757 & n39759;
  assign n39763 = ~n39547 & ~n58470;
  assign n39764 = ~n39440 & ~n39543;
  assign n39765 = ~n39544 & ~n39764;
  assign n39766 = ~n39763 & ~n39764;
  assign n39767 = ~n39544 & n39766;
  assign n39768 = ~n39763 & n39765;
  assign n39769 = ~n39544 & ~n58471;
  assign n39770 = ~n54667 & n39444;
  assign n39771 = ~n90 & n39770;
  assign n39772 = ~n53442 & n39444;
  assign n39773 = ~n90 & ~n54667;
  assign n39774 = n39444 & n39773;
  assign n39775 = ~n53442 & n14110;
  assign n39776 = pi23  & n58472;
  assign n39777 = ~pi23  & ~n58472;
  assign n39778 = ~n39776 & ~n39777;
  assign n39779 = ~n39470 & ~n39514;
  assign n39780 = ~n39513 & ~n39516;
  assign n39781 = ~n39513 & ~n39779;
  assign n39782 = ~n39778 & ~n58473;
  assign n39783 = n39778 & n58473;
  assign n39784 = ~n39782 & ~n39783;
  assign n39785 = ~n39491 & ~n39507;
  assign n39786 = n11279 & ~n56567;
  assign n39787 = n12584 & n26247;
  assign n39788 = n54410 & n26253;
  assign n39789 = n11267 & n26250;
  assign n39790 = ~n39788 & ~n39789;
  assign n39791 = ~n39787 & n39790;
  assign n39792 = ~n11279 & n39791;
  assign n39793 = n56567 & n39791;
  assign n39794 = ~n39792 & ~n39793;
  assign n39795 = ~n39786 & n39791;
  assign n39796 = pi29  & ~n58474;
  assign n39797 = ~pi29  & n58474;
  assign n39798 = ~n39796 & ~n39797;
  assign n39799 = ~n39472 & ~n39485;
  assign n39800 = n2140 & n8929;
  assign n39801 = n11793 & n39800;
  assign n39802 = ~n659 & ~n896;
  assign n39803 = n5485 & n39802;
  assign n39804 = n53679 & n39803;
  assign n39805 = n53612 & n11038;
  assign n39806 = n53612 & n53679;
  assign n39807 = n3476 & n39802;
  assign n39808 = n4378 & n5485;
  assign n39809 = n39807 & n39808;
  assign n39810 = n39806 & n39809;
  assign n39811 = n39804 & n39805;
  assign n39812 = n5485 & n39806;
  assign n39813 = n8929 & n39812;
  assign n39814 = n3476 & n39813;
  assign n39815 = n4378 & n39814;
  assign n39816 = ~n896 & n39815;
  assign n39817 = ~n184 & n39816;
  assign n39818 = ~n659 & n39817;
  assign n39819 = ~n357 & n39818;
  assign n39820 = ~n740 & n39819;
  assign n39821 = ~n770 & n39820;
  assign n39822 = n5485 & n8929;
  assign n39823 = n3476 & n39822;
  assign n39824 = n2140 & n11793;
  assign n39825 = n4378 & n39802;
  assign n39826 = n39824 & n39825;
  assign n39827 = n39806 & n39826;
  assign n39828 = n39823 & n39827;
  assign n39829 = n39801 & n58475;
  assign n39830 = n5277 & n9740;
  assign n39831 = n12005 & n39830;
  assign n39832 = ~n275 & n1278;
  assign n39833 = n3474 & n3535;
  assign n39834 = n39832 & n39833;
  assign n39835 = n3535 & n5277;
  assign n39836 = n9740 & n39835;
  assign n39837 = ~n275 & ~n956;
  assign n39838 = ~n275 & ~n618;
  assign n39839 = ~n956 & n39838;
  assign n39840 = ~n618 & n39837;
  assign n39841 = n1278 & n3474;
  assign n39842 = n58477 & n39841;
  assign n39843 = n39836 & n39842;
  assign n39844 = n1278 & n39833;
  assign n39845 = n39830 & n58477;
  assign n39846 = n39844 & n39845;
  assign n39847 = n39831 & n39834;
  assign n39848 = n53692 & n54454;
  assign n39849 = n53692 & n54932;
  assign n39850 = n54454 & n39849;
  assign n39851 = n54932 & n39848;
  assign n39852 = n58478 & n58479;
  assign n39853 = n58476 & n39852;
  assign n39854 = n56575 & n39853;
  assign n39855 = n3474 & n54932;
  assign n39856 = n54454 & n39855;
  assign n39857 = n53692 & n39856;
  assign n39858 = n56575 & n39857;
  assign n39859 = n58476 & n39858;
  assign n39860 = n54623 & n39859;
  assign n39861 = n3535 & n39860;
  assign n39862 = n5277 & n39861;
  assign n39863 = n1278 & n39862;
  assign n39864 = ~n894 & n39863;
  assign n39865 = ~n559 & n39864;
  assign n39866 = ~n956 & n39865;
  assign n39867 = ~n618 & n39866;
  assign n39868 = ~n275 & n39867;
  assign n39869 = n54623 & n39854;
  assign n39870 = ~n53600 & n58480;
  assign n39871 = n53600 & ~n58480;
  assign n39872 = ~n39870 & ~n39871;
  assign n39873 = ~n39799 & ~n39871;
  assign n39874 = ~n39870 & n39873;
  assign n39875 = ~n39799 & n39872;
  assign n39876 = n39799 & ~n39872;
  assign n39877 = ~n39799 & ~n58481;
  assign n39878 = ~n39870 & ~n58481;
  assign n39879 = ~n39871 & n39878;
  assign n39880 = ~n39877 & ~n39879;
  assign n39881 = ~n58481 & ~n39876;
  assign n39882 = n1576 & n27387;
  assign n39883 = n11215 & n26256;
  assign n39884 = n54403 & n26262;
  assign n39885 = n10564 & n26259;
  assign n39886 = ~n39884 & ~n39885;
  assign n39887 = ~n39883 & n39886;
  assign n39888 = ~n39882 & n39887;
  assign n39889 = ~n58482 & ~n39888;
  assign n39890 = n58482 & n39888;
  assign n39891 = ~n58482 & ~n39889;
  assign n39892 = ~n58482 & n39888;
  assign n39893 = ~n39888 & ~n39889;
  assign n39894 = n58482 & ~n39888;
  assign n39895 = ~n58483 & ~n58484;
  assign n39896 = ~n39889 & ~n39890;
  assign n39897 = ~n39798 & ~n58485;
  assign n39898 = n39798 & n58485;
  assign n39899 = ~n39897 & ~n39898;
  assign n39900 = ~n39785 & n39899;
  assign n39901 = n39785 & ~n39899;
  assign n39902 = ~n39900 & ~n39901;
  assign n39903 = n123 & ~n56564;
  assign n39904 = n128 & ~n26537;
  assign n39905 = n53444 & n26244;
  assign n39906 = n127 & n26242;
  assign n39907 = ~n39905 & ~n39906;
  assign n39908 = ~n39904 & n39907;
  assign n39909 = ~n39903 & n39908;
  assign n39910 = pi26  & ~n39909;
  assign n39911 = pi26  & ~n39910;
  assign n39912 = pi26  & n39909;
  assign n39913 = ~n39909 & ~n39910;
  assign n39914 = ~pi26  & ~n39909;
  assign n39915 = ~n58486 & ~n58487;
  assign n39916 = n39902 & ~n39915;
  assign n39917 = ~n39902 & n39915;
  assign n39918 = n39902 & ~n39916;
  assign n39919 = ~n39915 & ~n39916;
  assign n39920 = ~n39918 & ~n39919;
  assign n39921 = ~n39916 & ~n39917;
  assign n39922 = n39784 & ~n58488;
  assign n39923 = ~n39784 & n58488;
  assign n39924 = ~n58488 & ~n39922;
  assign n39925 = n39784 & ~n39922;
  assign n39926 = ~n39924 & ~n39925;
  assign n39927 = ~n39922 & ~n39923;
  assign n39928 = n39456 & ~n39525;
  assign n39929 = ~n39525 & ~n39528;
  assign n39930 = ~n39524 & ~n39928;
  assign n39931 = ~n58489 & ~n58490;
  assign n39932 = n58489 & n58490;
  assign n39933 = ~n39931 & ~n39932;
  assign n39934 = ~n39535 & ~n39541;
  assign n39935 = n39933 & ~n39934;
  assign n39936 = ~n39933 & n39934;
  assign n39937 = ~n39935 & ~n39936;
  assign n39938 = n39543 & n39937;
  assign n39939 = ~n39543 & ~n39937;
  assign n39940 = ~n39938 & ~n39939;
  assign n39941 = ~n39769 & n39940;
  assign n39942 = n39769 & ~n39940;
  assign n39943 = ~n39941 & ~n39942;
  assign n39944 = n77 & n39943;
  assign n39945 = n24302 & n39937;
  assign n39946 = n21969 & n39440;
  assign n39947 = n23459 & n39543;
  assign n39948 = ~n39946 & ~n39947;
  assign n39949 = ~n39945 & n39948;
  assign n39950 = ~n39944 & n39949;
  assign n39951 = pi5  & ~n39950;
  assign n39952 = ~n39950 & ~n39951;
  assign n39953 = ~pi5  & ~n39950;
  assign n39954 = pi5  & ~n39951;
  assign n39955 = pi5  & n39950;
  assign n39956 = ~n58491 & ~n58492;
  assign n39957 = n39725 & ~n39727;
  assign n39958 = ~n39725 & ~n58466;
  assign n39959 = ~n39726 & n39731;
  assign n39960 = ~n39958 & ~n39959;
  assign n39961 = ~n58466 & ~n39957;
  assign n39962 = n18846 & ~n58493;
  assign n39963 = n19541 & n39561;
  assign n39964 = n55247 & n39567;
  assign n39965 = n19509 & n39564;
  assign n39966 = ~n39964 & ~n39965;
  assign n39967 = ~n39963 & n39966;
  assign n39968 = ~n39962 & n39967;
  assign n39969 = pi11  & ~n39968;
  assign n39970 = ~n39968 & ~n39969;
  assign n39971 = ~pi11  & ~n39968;
  assign n39972 = pi11  & ~n39969;
  assign n39973 = pi11  & n39968;
  assign n39974 = ~n58494 & ~n58495;
  assign n39975 = n39705 & ~n39707;
  assign n39976 = ~n39708 & ~n39975;
  assign n39977 = n17265 & n39976;
  assign n39978 = n18588 & n39573;
  assign n39979 = n55041 & n39579;
  assign n39980 = n18556 & n39576;
  assign n39981 = ~n39979 & ~n39980;
  assign n39982 = ~n39978 & n39981;
  assign n39983 = ~n39977 & n39982;
  assign n39984 = pi14  & ~n39983;
  assign n39985 = ~n39983 & ~n39984;
  assign n39986 = ~pi14  & ~n39983;
  assign n39987 = pi14  & ~n39984;
  assign n39988 = pi14  & n39983;
  assign n39989 = ~n58496 & ~n58497;
  assign n39990 = n39647 & ~n39649;
  assign n39991 = ~n39650 & ~n39990;
  assign n39992 = n90 & n39991;
  assign n39993 = n14236 & n39609;
  assign n39994 = n54667 & n39615;
  assign n39995 = n14210 & n39612;
  assign n39996 = ~n39994 & ~n39995;
  assign n39997 = ~n39993 & n39996;
  assign n39998 = ~n90 & n39997;
  assign n39999 = ~n39991 & n39997;
  assign n40000 = ~n39998 & ~n39999;
  assign n40001 = ~n39992 & n39997;
  assign n40002 = pi23  & ~n58498;
  assign n40003 = ~pi23  & n58498;
  assign n40004 = ~n40002 & ~n40003;
  assign n40005 = ~n39624 & n58458;
  assign n40006 = ~n39638 & ~n40005;
  assign n40007 = n123 & n40006;
  assign n40008 = n128 & n39618;
  assign n40009 = n53444 & n39626;
  assign n40010 = n127 & n39621;
  assign n40011 = ~n40009 & ~n40010;
  assign n40012 = ~n40008 & n40011;
  assign n40013 = ~n40007 & n40012;
  assign n40014 = pi26  & ~n40013;
  assign n40015 = pi26  & ~n40014;
  assign n40016 = pi26  & n40013;
  assign n40017 = ~n40013 & ~n40014;
  assign n40018 = ~pi26  & ~n40013;
  assign n40019 = ~n58499 & ~n58500;
  assign n40020 = n54407 & ~n58457;
  assign n40021 = n39626 & n58457;
  assign n40022 = ~n39626 & ~n58457;
  assign n40023 = ~n40021 & ~n40022;
  assign n40024 = n123 & ~n40023;
  assign n40025 = n127 & ~n58457;
  assign n40026 = n128 & n39626;
  assign n40027 = ~n40025 & ~n40026;
  assign n40028 = ~n40024 & n40027;
  assign n40029 = ~n120 & ~n58457;
  assign n40030 = pi26  & ~n40029;
  assign n40031 = pi26  & ~n40028;
  assign n40032 = pi26  & ~n40031;
  assign n40033 = ~n40028 & ~n40031;
  assign n40034 = ~n40032 & ~n40033;
  assign n40035 = n40030 & ~n40034;
  assign n40036 = n40028 & n40030;
  assign n40037 = n39621 & ~n40021;
  assign n40038 = ~n39621 & n40021;
  assign n40039 = ~n40037 & ~n40038;
  assign n40040 = n123 & ~n40039;
  assign n40041 = n128 & n39621;
  assign n40042 = n53444 & ~n58457;
  assign n40043 = n127 & n39626;
  assign n40044 = ~n40042 & ~n40043;
  assign n40045 = ~n40041 & n40044;
  assign n40046 = ~n123 & n40045;
  assign n40047 = n40039 & n40045;
  assign n40048 = ~n40046 & ~n40047;
  assign n40049 = ~n40040 & n40045;
  assign n40050 = pi26  & ~n58502;
  assign n40051 = ~pi26  & n58502;
  assign n40052 = ~n40050 & ~n40051;
  assign n40053 = n58501 & ~n40052;
  assign n40054 = n58501 & ~n58502;
  assign n40055 = n40020 & n58503;
  assign n40056 = ~n40020 & ~n58503;
  assign n40057 = n58503 & ~n40055;
  assign n40058 = ~n40020 & n58503;
  assign n40059 = n40020 & ~n40055;
  assign n40060 = n40020 & ~n58503;
  assign n40061 = ~n58504 & ~n58505;
  assign n40062 = ~n40055 & ~n40056;
  assign n40063 = ~n40019 & ~n58506;
  assign n40064 = n40019 & n58506;
  assign n40065 = ~n58506 & ~n40063;
  assign n40066 = ~n40019 & ~n40063;
  assign n40067 = ~n40065 & ~n40066;
  assign n40068 = ~n40063 & ~n40064;
  assign n40069 = ~n40004 & ~n58507;
  assign n40070 = n39643 & ~n39645;
  assign n40071 = ~n39646 & ~n40070;
  assign n40072 = n90 & n40071;
  assign n40073 = n14236 & n39612;
  assign n40074 = n54667 & n39618;
  assign n40075 = n14210 & n39615;
  assign n40076 = ~n40074 & ~n40075;
  assign n40077 = ~n40073 & n40076;
  assign n40078 = ~n40072 & n40077;
  assign n40079 = pi23  & ~n40078;
  assign n40080 = ~n40078 & ~n40079;
  assign n40081 = ~pi23  & ~n40078;
  assign n40082 = pi23  & ~n40079;
  assign n40083 = pi23  & n40078;
  assign n40084 = ~n58508 & ~n58509;
  assign n40085 = pi26  & ~n58501;
  assign n40086 = ~n58502 & ~n40085;
  assign n40087 = n58502 & n40085;
  assign n40088 = ~n58501 & n40052;
  assign n40089 = ~n58503 & ~n40088;
  assign n40090 = ~n40086 & ~n40087;
  assign n40091 = ~n40084 & n58510;
  assign n40092 = n39639 & ~n39641;
  assign n40093 = ~n39642 & ~n40092;
  assign n40094 = n90 & n40093;
  assign n40095 = n14236 & n39615;
  assign n40096 = n54667 & n39621;
  assign n40097 = n14210 & n39618;
  assign n40098 = ~n40096 & ~n40097;
  assign n40099 = ~n40095 & n40098;
  assign n40100 = ~n90 & n40099;
  assign n40101 = ~n40093 & n40099;
  assign n40102 = ~n40100 & ~n40101;
  assign n40103 = ~n40094 & n40099;
  assign n40104 = pi23  & ~n58511;
  assign n40105 = ~pi23  & n58511;
  assign n40106 = ~n40104 & ~n40105;
  assign n40107 = pi26  & n40029;
  assign n40108 = ~n40028 & n40107;
  assign n40109 = n40028 & ~n40107;
  assign n40110 = ~n40030 & n40034;
  assign n40111 = ~n58501 & ~n40110;
  assign n40112 = ~n40108 & ~n40109;
  assign n40113 = ~n40106 & n58512;
  assign n40114 = n90 & ~n40023;
  assign n40115 = n14210 & ~n58457;
  assign n40116 = n14236 & n39626;
  assign n40117 = ~n40115 & ~n40116;
  assign n40118 = ~n40114 & n40117;
  assign n40119 = n53441 & ~n58457;
  assign n40120 = pi23  & ~n40119;
  assign n40121 = pi23  & ~n40118;
  assign n40122 = pi23  & ~n40121;
  assign n40123 = ~n40118 & ~n40121;
  assign n40124 = ~n40122 & ~n40123;
  assign n40125 = n40120 & ~n40124;
  assign n40126 = n40118 & n40120;
  assign n40127 = n90 & ~n40039;
  assign n40128 = n14236 & n39621;
  assign n40129 = n54667 & ~n58457;
  assign n40130 = n14210 & n39626;
  assign n40131 = ~n40129 & ~n40130;
  assign n40132 = ~n40128 & n40131;
  assign n40133 = ~n90 & n40132;
  assign n40134 = n40039 & n40132;
  assign n40135 = ~n40133 & ~n40134;
  assign n40136 = ~n40127 & n40132;
  assign n40137 = pi23  & ~n58514;
  assign n40138 = ~pi23  & n58514;
  assign n40139 = ~n40137 & ~n40138;
  assign n40140 = n58513 & ~n40139;
  assign n40141 = n58513 & ~n58514;
  assign n40142 = n40029 & n58515;
  assign n40143 = n90 & n40006;
  assign n40144 = n14236 & n39618;
  assign n40145 = n54667 & n39626;
  assign n40146 = n14210 & n39621;
  assign n40147 = ~n40145 & ~n40146;
  assign n40148 = ~n40144 & n40147;
  assign n40149 = ~n40143 & n40148;
  assign n40150 = pi23  & ~n40149;
  assign n40151 = pi23  & ~n40150;
  assign n40152 = pi23  & n40149;
  assign n40153 = ~n40149 & ~n40150;
  assign n40154 = ~pi23  & ~n40149;
  assign n40155 = ~n58516 & ~n58517;
  assign n40156 = ~n40029 & ~n58515;
  assign n40157 = n58515 & ~n40142;
  assign n40158 = ~n40029 & n58515;
  assign n40159 = n40029 & ~n40142;
  assign n40160 = n40029 & ~n58515;
  assign n40161 = ~n58518 & ~n58519;
  assign n40162 = ~n40142 & ~n40156;
  assign n40163 = ~n40155 & ~n58520;
  assign n40164 = ~n40142 & ~n40163;
  assign n40165 = n40106 & ~n58512;
  assign n40166 = ~n40113 & ~n40165;
  assign n40167 = ~n40164 & n40166;
  assign n40168 = ~n40113 & ~n40167;
  assign n40169 = n40084 & ~n58510;
  assign n40170 = ~n40084 & ~n40091;
  assign n40171 = ~n40084 & ~n58510;
  assign n40172 = n58510 & ~n40091;
  assign n40173 = n40084 & n58510;
  assign n40174 = ~n58521 & ~n58522;
  assign n40175 = ~n40091 & ~n40169;
  assign n40176 = ~n40168 & ~n58523;
  assign n40177 = ~n40091 & ~n40176;
  assign n40178 = n40004 & n58507;
  assign n40179 = ~n40069 & ~n40178;
  assign n40180 = ~n40177 & n40179;
  assign n40181 = ~n40069 & ~n40180;
  assign n40182 = n39651 & ~n39653;
  assign n40183 = ~n39654 & ~n40182;
  assign n40184 = n90 & n40183;
  assign n40185 = n14236 & n39606;
  assign n40186 = n54667 & n39612;
  assign n40187 = n14210 & n39609;
  assign n40188 = ~n40186 & ~n40187;
  assign n40189 = ~n40185 & n40188;
  assign n40190 = ~n40184 & n40189;
  assign n40191 = pi23  & ~n40190;
  assign n40192 = ~n40190 & ~n40191;
  assign n40193 = ~pi23  & ~n40190;
  assign n40194 = pi23  & ~n40191;
  assign n40195 = pi23  & n40190;
  assign n40196 = ~n58524 & ~n58525;
  assign n40197 = ~n40055 & ~n40063;
  assign n40198 = n123 & n40093;
  assign n40199 = n128 & n39615;
  assign n40200 = n53444 & n39621;
  assign n40201 = n127 & n39618;
  assign n40202 = ~n40200 & ~n40201;
  assign n40203 = ~n40199 & n40202;
  assign n40204 = ~n123 & n40203;
  assign n40205 = ~n40093 & n40203;
  assign n40206 = ~n40204 & ~n40205;
  assign n40207 = ~n40198 & n40203;
  assign n40208 = pi26  & ~n58526;
  assign n40209 = ~pi26  & n58526;
  assign n40210 = ~n40208 & ~n40209;
  assign n40211 = pi29  & n40020;
  assign n40212 = n11279 & ~n40023;
  assign n40213 = n11267 & ~n58457;
  assign n40214 = n12584 & n39626;
  assign n40215 = ~n40213 & ~n40214;
  assign n40216 = ~n40212 & n40215;
  assign n40217 = n40211 & ~n40216;
  assign n40218 = ~n40211 & n40216;
  assign n40219 = pi29  & ~n40020;
  assign n40220 = pi29  & ~n40216;
  assign n40221 = pi29  & ~n40220;
  assign n40222 = ~n40216 & ~n40220;
  assign n40223 = ~n40221 & ~n40222;
  assign n40224 = n40219 & ~n40223;
  assign n40225 = n40216 & n40219;
  assign n40226 = ~n40219 & n40223;
  assign n40227 = ~n58527 & ~n40226;
  assign n40228 = ~n40217 & ~n40218;
  assign n40229 = ~n40210 & n58528;
  assign n40230 = n40210 & ~n58528;
  assign n40231 = ~n40229 & ~n40230;
  assign n40232 = ~n40197 & n40231;
  assign n40233 = n40197 & ~n40231;
  assign n40234 = ~n40232 & ~n40233;
  assign n40235 = ~n40196 & n40234;
  assign n40236 = n40196 & ~n40234;
  assign n40237 = ~n40196 & ~n40235;
  assign n40238 = ~n40196 & ~n40234;
  assign n40239 = n40234 & ~n40235;
  assign n40240 = n40196 & n40234;
  assign n40241 = ~n58529 & ~n58530;
  assign n40242 = ~n40235 & ~n40236;
  assign n40243 = ~n40181 & ~n58531;
  assign n40244 = n40181 & n58531;
  assign n40245 = ~n40243 & ~n40244;
  assign n40246 = n39665 & ~n39667;
  assign n40247 = ~n39668 & ~n40246;
  assign n40248 = n14413 & n40247;
  assign n40249 = n15921 & n39597;
  assign n40250 = n54719 & n39603;
  assign n40251 = n15901 & n39600;
  assign n40252 = ~n40250 & ~n40251;
  assign n40253 = ~n40249 & n40252;
  assign n40254 = ~n14413 & n40253;
  assign n40255 = ~n40247 & n40253;
  assign n40256 = ~n40254 & ~n40255;
  assign n40257 = ~n40248 & n40253;
  assign n40258 = pi20  & ~n58532;
  assign n40259 = ~pi20  & n58532;
  assign n40260 = ~n40258 & ~n40259;
  assign n40261 = n40245 & ~n40260;
  assign n40262 = n40177 & ~n40179;
  assign n40263 = ~n40180 & ~n40262;
  assign n40264 = n39659 & ~n39661;
  assign n40265 = ~n39659 & ~n58459;
  assign n40266 = ~n39660 & n39665;
  assign n40267 = ~n40265 & ~n40266;
  assign n40268 = ~n58459 & ~n40264;
  assign n40269 = n14413 & ~n58533;
  assign n40270 = n15921 & n39600;
  assign n40271 = n54719 & n39606;
  assign n40272 = n15901 & n39603;
  assign n40273 = ~n40271 & ~n40272;
  assign n40274 = ~n40270 & n40273;
  assign n40275 = ~n14413 & n40274;
  assign n40276 = n58533 & n40274;
  assign n40277 = ~n40275 & ~n40276;
  assign n40278 = ~n40269 & n40274;
  assign n40279 = pi20  & ~n58534;
  assign n40280 = ~pi20  & n58534;
  assign n40281 = ~n40279 & ~n40280;
  assign n40282 = n40263 & ~n40281;
  assign n40283 = n40168 & n58523;
  assign n40284 = ~n40176 & ~n40283;
  assign n40285 = n39655 & ~n39657;
  assign n40286 = ~n39658 & ~n40285;
  assign n40287 = n14413 & n40286;
  assign n40288 = n15921 & n39603;
  assign n40289 = n54719 & n39609;
  assign n40290 = n15901 & n39606;
  assign n40291 = ~n40289 & ~n40290;
  assign n40292 = ~n40288 & n40291;
  assign n40293 = ~n14413 & n40292;
  assign n40294 = ~n40286 & n40292;
  assign n40295 = ~n40293 & ~n40294;
  assign n40296 = ~n40287 & n40292;
  assign n40297 = pi20  & ~n58535;
  assign n40298 = ~pi20  & n58535;
  assign n40299 = ~n40297 & ~n40298;
  assign n40300 = n40284 & ~n40299;
  assign n40301 = n14413 & n40183;
  assign n40302 = n15921 & n39606;
  assign n40303 = n54719 & n39612;
  assign n40304 = n15901 & n39609;
  assign n40305 = ~n40303 & ~n40304;
  assign n40306 = ~n40302 & n40305;
  assign n40307 = ~n40301 & n40306;
  assign n40308 = pi20  & ~n40307;
  assign n40309 = ~n40307 & ~n40308;
  assign n40310 = ~pi20  & ~n40307;
  assign n40311 = pi20  & ~n40308;
  assign n40312 = pi20  & n40307;
  assign n40313 = ~n58536 & ~n58537;
  assign n40314 = n40164 & ~n40166;
  assign n40315 = ~n40167 & ~n40314;
  assign n40316 = ~n40313 & n40315;
  assign n40317 = n14413 & n39991;
  assign n40318 = n15921 & n39609;
  assign n40319 = n54719 & n39615;
  assign n40320 = n15901 & n39612;
  assign n40321 = ~n40319 & ~n40320;
  assign n40322 = ~n40318 & n40321;
  assign n40323 = ~n14413 & n40322;
  assign n40324 = ~n39991 & n40322;
  assign n40325 = ~n40323 & ~n40324;
  assign n40326 = ~n40317 & n40322;
  assign n40327 = pi20  & ~n58538;
  assign n40328 = ~pi20  & n58538;
  assign n40329 = ~n40327 & ~n40328;
  assign n40330 = n40155 & n58520;
  assign n40331 = ~n58520 & ~n40163;
  assign n40332 = ~n40155 & ~n40163;
  assign n40333 = ~n40331 & ~n40332;
  assign n40334 = ~n40163 & ~n40330;
  assign n40335 = ~n40329 & ~n58539;
  assign n40336 = n14413 & n40071;
  assign n40337 = n15921 & n39612;
  assign n40338 = n54719 & n39618;
  assign n40339 = n15901 & n39615;
  assign n40340 = ~n40338 & ~n40339;
  assign n40341 = ~n40337 & n40340;
  assign n40342 = ~n40336 & n40341;
  assign n40343 = pi20  & ~n40342;
  assign n40344 = ~n40342 & ~n40343;
  assign n40345 = ~pi20  & ~n40342;
  assign n40346 = pi20  & ~n40343;
  assign n40347 = pi20  & n40342;
  assign n40348 = ~n58540 & ~n58541;
  assign n40349 = pi23  & ~n58513;
  assign n40350 = ~n58514 & ~n40349;
  assign n40351 = n58514 & n40349;
  assign n40352 = ~n58513 & n40139;
  assign n40353 = ~n58515 & ~n40352;
  assign n40354 = ~n40350 & ~n40351;
  assign n40355 = ~n40348 & n58542;
  assign n40356 = n14413 & n40093;
  assign n40357 = n15921 & n39615;
  assign n40358 = n54719 & n39621;
  assign n40359 = n15901 & n39618;
  assign n40360 = ~n40358 & ~n40359;
  assign n40361 = ~n40357 & n40360;
  assign n40362 = ~n14413 & n40361;
  assign n40363 = ~n40093 & n40361;
  assign n40364 = ~n40362 & ~n40363;
  assign n40365 = ~n40356 & n40361;
  assign n40366 = pi20  & ~n58543;
  assign n40367 = ~pi20  & n58543;
  assign n40368 = ~n40366 & ~n40367;
  assign n40369 = pi23  & n40119;
  assign n40370 = ~n40118 & n40369;
  assign n40371 = n40118 & ~n40369;
  assign n40372 = ~n40120 & n40124;
  assign n40373 = ~n58513 & ~n40372;
  assign n40374 = ~n40370 & ~n40371;
  assign n40375 = ~n40368 & n58544;
  assign n40376 = n14413 & ~n40023;
  assign n40377 = n15901 & ~n58457;
  assign n40378 = n15921 & n39626;
  assign n40379 = ~n40377 & ~n40378;
  assign n40380 = ~n40376 & n40379;
  assign n40381 = n54717 & ~n58457;
  assign n40382 = pi20  & ~n40381;
  assign n40383 = pi20  & ~n40380;
  assign n40384 = pi20  & ~n40383;
  assign n40385 = ~n40380 & ~n40383;
  assign n40386 = ~n40384 & ~n40385;
  assign n40387 = n40382 & ~n40386;
  assign n40388 = n40380 & n40382;
  assign n40389 = n14413 & ~n40039;
  assign n40390 = n15921 & n39621;
  assign n40391 = n54719 & ~n58457;
  assign n40392 = n15901 & n39626;
  assign n40393 = ~n40391 & ~n40392;
  assign n40394 = ~n40390 & n40393;
  assign n40395 = ~n14413 & n40394;
  assign n40396 = n40039 & n40394;
  assign n40397 = ~n40395 & ~n40396;
  assign n40398 = ~n40389 & n40394;
  assign n40399 = pi20  & ~n58546;
  assign n40400 = ~pi20  & n58546;
  assign n40401 = ~n40399 & ~n40400;
  assign n40402 = n58545 & ~n40401;
  assign n40403 = n58545 & ~n58546;
  assign n40404 = n40119 & n58547;
  assign n40405 = n14413 & n40006;
  assign n40406 = n15921 & n39618;
  assign n40407 = n54719 & n39626;
  assign n40408 = n15901 & n39621;
  assign n40409 = ~n40407 & ~n40408;
  assign n40410 = ~n40406 & n40409;
  assign n40411 = ~n40405 & n40410;
  assign n40412 = pi20  & ~n40411;
  assign n40413 = pi20  & ~n40412;
  assign n40414 = pi20  & n40411;
  assign n40415 = ~n40411 & ~n40412;
  assign n40416 = ~pi20  & ~n40411;
  assign n40417 = ~n58548 & ~n58549;
  assign n40418 = ~n40119 & ~n58547;
  assign n40419 = n58547 & ~n40404;
  assign n40420 = ~n40119 & n58547;
  assign n40421 = n40119 & ~n40404;
  assign n40422 = n40119 & ~n58547;
  assign n40423 = ~n58550 & ~n58551;
  assign n40424 = ~n40404 & ~n40418;
  assign n40425 = ~n40417 & ~n58552;
  assign n40426 = ~n40404 & ~n40425;
  assign n40427 = n40368 & ~n58544;
  assign n40428 = ~n40375 & ~n40427;
  assign n40429 = ~n40426 & n40428;
  assign n40430 = ~n40375 & ~n40429;
  assign n40431 = n40348 & ~n58542;
  assign n40432 = ~n40348 & ~n40355;
  assign n40433 = ~n40348 & ~n58542;
  assign n40434 = n58542 & ~n40355;
  assign n40435 = n40348 & n58542;
  assign n40436 = ~n58553 & ~n58554;
  assign n40437 = ~n40355 & ~n40431;
  assign n40438 = ~n40430 & ~n58555;
  assign n40439 = ~n40355 & ~n40438;
  assign n40440 = n40329 & n58539;
  assign n40441 = ~n40335 & ~n40440;
  assign n40442 = ~n40439 & n40441;
  assign n40443 = ~n40335 & ~n40442;
  assign n40444 = n40313 & ~n40315;
  assign n40445 = ~n40313 & ~n40316;
  assign n40446 = ~n40313 & ~n40315;
  assign n40447 = n40315 & ~n40316;
  assign n40448 = n40313 & n40315;
  assign n40449 = ~n58556 & ~n58557;
  assign n40450 = ~n40316 & ~n40444;
  assign n40451 = ~n40443 & ~n58558;
  assign n40452 = ~n40316 & ~n40451;
  assign n40453 = ~n40284 & n40299;
  assign n40454 = n40284 & ~n40300;
  assign n40455 = n40284 & n40299;
  assign n40456 = ~n40299 & ~n40300;
  assign n40457 = ~n40284 & ~n40299;
  assign n40458 = ~n58559 & ~n58560;
  assign n40459 = ~n40300 & ~n40453;
  assign n40460 = ~n40452 & ~n58561;
  assign n40461 = ~n40300 & ~n40460;
  assign n40462 = ~n40263 & n40281;
  assign n40463 = n40263 & ~n40282;
  assign n40464 = n40263 & n40281;
  assign n40465 = ~n40281 & ~n40282;
  assign n40466 = ~n40263 & ~n40281;
  assign n40467 = ~n58562 & ~n58563;
  assign n40468 = ~n40282 & ~n40462;
  assign n40469 = ~n40461 & ~n58564;
  assign n40470 = ~n40282 & ~n40469;
  assign n40471 = ~n40245 & n40260;
  assign n40472 = ~n40261 & ~n40471;
  assign n40473 = ~n40470 & n40472;
  assign n40474 = ~n40261 & ~n40473;
  assign n40475 = n39669 & ~n39671;
  assign n40476 = ~n39672 & ~n40475;
  assign n40477 = n14413 & n40476;
  assign n40478 = n15921 & n39594;
  assign n40479 = n54719 & n39600;
  assign n40480 = n15901 & n39597;
  assign n40481 = ~n40479 & ~n40480;
  assign n40482 = ~n40478 & n40481;
  assign n40483 = ~n40477 & n40482;
  assign n40484 = pi20  & ~n40483;
  assign n40485 = ~n40483 & ~n40484;
  assign n40486 = ~pi20  & ~n40483;
  assign n40487 = pi20  & ~n40484;
  assign n40488 = pi20  & n40483;
  assign n40489 = ~n58565 & ~n58566;
  assign n40490 = ~n40235 & ~n40243;
  assign n40491 = ~n40229 & ~n40232;
  assign n40492 = n123 & n40071;
  assign n40493 = n128 & n39612;
  assign n40494 = n53444 & n39618;
  assign n40495 = n127 & n39615;
  assign n40496 = ~n40494 & ~n40495;
  assign n40497 = ~n40493 & n40496;
  assign n40498 = ~n40492 & n40497;
  assign n40499 = pi26  & ~n40498;
  assign n40500 = ~n40498 & ~n40499;
  assign n40501 = ~pi26  & ~n40498;
  assign n40502 = pi26  & ~n40499;
  assign n40503 = pi26  & n40498;
  assign n40504 = ~n58567 & ~n58568;
  assign n40505 = pi29  & ~n58527;
  assign n40506 = n11279 & ~n40039;
  assign n40507 = n12584 & n39621;
  assign n40508 = n54410 & ~n58457;
  assign n40509 = n11267 & n39626;
  assign n40510 = ~n40508 & ~n40509;
  assign n40511 = ~n40507 & n40510;
  assign n40512 = ~n11279 & n40511;
  assign n40513 = n40039 & n40511;
  assign n40514 = ~n40512 & ~n40513;
  assign n40515 = ~n40506 & n40511;
  assign n40516 = ~n40505 & ~n58569;
  assign n40517 = n40505 & n58569;
  assign n40518 = pi29  & ~n58569;
  assign n40519 = ~pi29  & n58569;
  assign n40520 = ~n40518 & ~n40519;
  assign n40521 = n58527 & ~n40520;
  assign n40522 = n58527 & ~n58569;
  assign n40523 = ~n58527 & n40520;
  assign n40524 = ~n58570 & ~n40523;
  assign n40525 = ~n40516 & ~n40517;
  assign n40526 = ~n40504 & n58571;
  assign n40527 = n40504 & ~n58571;
  assign n40528 = ~n40504 & ~n40526;
  assign n40529 = ~n40504 & ~n58571;
  assign n40530 = n58571 & ~n40526;
  assign n40531 = n40504 & n58571;
  assign n40532 = ~n58572 & ~n58573;
  assign n40533 = ~n40526 & ~n40527;
  assign n40534 = ~n40491 & ~n58574;
  assign n40535 = n40491 & n58574;
  assign n40536 = ~n40534 & ~n40535;
  assign n40537 = n90 & n40286;
  assign n40538 = n14236 & n39603;
  assign n40539 = n54667 & n39609;
  assign n40540 = n14210 & n39606;
  assign n40541 = ~n40539 & ~n40540;
  assign n40542 = ~n40538 & n40541;
  assign n40543 = ~n90 & n40542;
  assign n40544 = ~n40286 & n40542;
  assign n40545 = ~n40543 & ~n40544;
  assign n40546 = ~n40537 & n40542;
  assign n40547 = pi23  & ~n58575;
  assign n40548 = ~pi23  & n58575;
  assign n40549 = ~n40547 & ~n40548;
  assign n40550 = n40536 & ~n40549;
  assign n40551 = ~n40536 & n40549;
  assign n40552 = n40536 & ~n40550;
  assign n40553 = n40536 & n40549;
  assign n40554 = ~n40549 & ~n40550;
  assign n40555 = ~n40536 & ~n40549;
  assign n40556 = ~n58576 & ~n58577;
  assign n40557 = ~n40550 & ~n40551;
  assign n40558 = ~n40490 & ~n58578;
  assign n40559 = n40490 & n58578;
  assign n40560 = ~n40490 & ~n40558;
  assign n40561 = ~n40490 & n58578;
  assign n40562 = ~n58578 & ~n40558;
  assign n40563 = n40490 & ~n58578;
  assign n40564 = ~n58579 & ~n58580;
  assign n40565 = ~n40558 & ~n40559;
  assign n40566 = ~n40489 & ~n58581;
  assign n40567 = n40489 & n58581;
  assign n40568 = ~n40489 & ~n40566;
  assign n40569 = ~n58581 & ~n40566;
  assign n40570 = ~n40568 & ~n40569;
  assign n40571 = ~n40566 & ~n40567;
  assign n40572 = ~n40474 & ~n58582;
  assign n40573 = n40474 & n58582;
  assign n40574 = ~n40572 & ~n40573;
  assign n40575 = n39683 & ~n39685;
  assign n40576 = ~n39683 & ~n58461;
  assign n40577 = ~n39684 & n39689;
  assign n40578 = ~n40576 & ~n40577;
  assign n40579 = ~n58461 & ~n40575;
  assign n40580 = n16079 & ~n58583;
  assign n40581 = n16696 & n39585;
  assign n40582 = n54886 & n39591;
  assign n40583 = n16676 & n39588;
  assign n40584 = ~n40582 & ~n40583;
  assign n40585 = ~n40581 & n40584;
  assign n40586 = ~n16079 & n40585;
  assign n40587 = n58583 & n40585;
  assign n40588 = ~n40586 & ~n40587;
  assign n40589 = ~n40580 & n40585;
  assign n40590 = pi17  & ~n58584;
  assign n40591 = ~pi17  & n58584;
  assign n40592 = ~n40590 & ~n40591;
  assign n40593 = n40574 & ~n40592;
  assign n40594 = n39677 & ~n39679;
  assign n40595 = ~n39677 & ~n58460;
  assign n40596 = ~n39678 & n39683;
  assign n40597 = ~n40595 & ~n40596;
  assign n40598 = ~n58460 & ~n40594;
  assign n40599 = n16079 & ~n58585;
  assign n40600 = n16696 & n39588;
  assign n40601 = n54886 & n39594;
  assign n40602 = n16676 & n39591;
  assign n40603 = ~n40601 & ~n40602;
  assign n40604 = ~n40600 & n40603;
  assign n40605 = ~n40599 & n40604;
  assign n40606 = pi17  & ~n40605;
  assign n40607 = ~n40605 & ~n40606;
  assign n40608 = ~pi17  & ~n40605;
  assign n40609 = pi17  & ~n40606;
  assign n40610 = pi17  & n40605;
  assign n40611 = ~n58586 & ~n58587;
  assign n40612 = n40470 & ~n40472;
  assign n40613 = ~n40473 & ~n40612;
  assign n40614 = ~n40611 & n40613;
  assign n40615 = n39673 & ~n39675;
  assign n40616 = ~n39676 & ~n40615;
  assign n40617 = n16079 & n40616;
  assign n40618 = n16696 & n39591;
  assign n40619 = n54886 & n39597;
  assign n40620 = n16676 & n39594;
  assign n40621 = ~n40619 & ~n40620;
  assign n40622 = ~n40618 & n40621;
  assign n40623 = ~n40617 & n40622;
  assign n40624 = pi17  & ~n40623;
  assign n40625 = ~n40623 & ~n40624;
  assign n40626 = ~pi17  & ~n40623;
  assign n40627 = pi17  & ~n40624;
  assign n40628 = pi17  & n40623;
  assign n40629 = ~n58588 & ~n58589;
  assign n40630 = n40461 & n58564;
  assign n40631 = ~n40461 & ~n40469;
  assign n40632 = ~n58564 & ~n40469;
  assign n40633 = ~n40631 & ~n40632;
  assign n40634 = ~n40469 & ~n40630;
  assign n40635 = ~n40629 & ~n58590;
  assign n40636 = n16079 & n40476;
  assign n40637 = n16696 & n39594;
  assign n40638 = n54886 & n39600;
  assign n40639 = n16676 & n39597;
  assign n40640 = ~n40638 & ~n40639;
  assign n40641 = ~n40637 & n40640;
  assign n40642 = ~n40636 & n40641;
  assign n40643 = pi17  & ~n40642;
  assign n40644 = ~n40642 & ~n40643;
  assign n40645 = ~pi17  & ~n40642;
  assign n40646 = pi17  & ~n40643;
  assign n40647 = pi17  & n40642;
  assign n40648 = ~n58591 & ~n58592;
  assign n40649 = n40452 & n58561;
  assign n40650 = ~n40452 & ~n40460;
  assign n40651 = ~n40452 & n58561;
  assign n40652 = ~n58561 & ~n40460;
  assign n40653 = n40452 & ~n58561;
  assign n40654 = ~n58593 & ~n58594;
  assign n40655 = ~n40460 & ~n40649;
  assign n40656 = ~n40648 & ~n58595;
  assign n40657 = n40443 & n58558;
  assign n40658 = ~n40451 & ~n40657;
  assign n40659 = n16079 & n40247;
  assign n40660 = n16696 & n39597;
  assign n40661 = n54886 & n39603;
  assign n40662 = n16676 & n39600;
  assign n40663 = ~n40661 & ~n40662;
  assign n40664 = ~n40660 & n40663;
  assign n40665 = ~n16079 & n40664;
  assign n40666 = ~n40247 & n40664;
  assign n40667 = ~n40665 & ~n40666;
  assign n40668 = ~n40659 & n40664;
  assign n40669 = pi17  & ~n58596;
  assign n40670 = ~pi17  & n58596;
  assign n40671 = ~n40669 & ~n40670;
  assign n40672 = n40658 & ~n40671;
  assign n40673 = n40439 & ~n40441;
  assign n40674 = ~n40442 & ~n40673;
  assign n40675 = n16079 & ~n58533;
  assign n40676 = n16696 & n39600;
  assign n40677 = n54886 & n39606;
  assign n40678 = n16676 & n39603;
  assign n40679 = ~n40677 & ~n40678;
  assign n40680 = ~n40676 & n40679;
  assign n40681 = ~n16079 & n40680;
  assign n40682 = n58533 & n40680;
  assign n40683 = ~n40681 & ~n40682;
  assign n40684 = ~n40675 & n40680;
  assign n40685 = pi17  & ~n58597;
  assign n40686 = ~pi17  & n58597;
  assign n40687 = ~n40685 & ~n40686;
  assign n40688 = n40674 & ~n40687;
  assign n40689 = n40430 & n58555;
  assign n40690 = ~n40438 & ~n40689;
  assign n40691 = n16079 & n40286;
  assign n40692 = n16696 & n39603;
  assign n40693 = n54886 & n39609;
  assign n40694 = n16676 & n39606;
  assign n40695 = ~n40693 & ~n40694;
  assign n40696 = ~n40692 & n40695;
  assign n40697 = ~n16079 & n40696;
  assign n40698 = ~n40286 & n40696;
  assign n40699 = ~n40697 & ~n40698;
  assign n40700 = ~n40691 & n40696;
  assign n40701 = pi17  & ~n58598;
  assign n40702 = ~pi17  & n58598;
  assign n40703 = ~n40701 & ~n40702;
  assign n40704 = n40690 & ~n40703;
  assign n40705 = n16079 & n40183;
  assign n40706 = n16696 & n39606;
  assign n40707 = n54886 & n39612;
  assign n40708 = n16676 & n39609;
  assign n40709 = ~n40707 & ~n40708;
  assign n40710 = ~n40706 & n40709;
  assign n40711 = ~n40705 & n40710;
  assign n40712 = pi17  & ~n40711;
  assign n40713 = ~n40711 & ~n40712;
  assign n40714 = ~pi17  & ~n40711;
  assign n40715 = pi17  & ~n40712;
  assign n40716 = pi17  & n40711;
  assign n40717 = ~n58599 & ~n58600;
  assign n40718 = n40426 & ~n40428;
  assign n40719 = ~n40429 & ~n40718;
  assign n40720 = ~n40717 & n40719;
  assign n40721 = n16079 & n39991;
  assign n40722 = n16696 & n39609;
  assign n40723 = n54886 & n39615;
  assign n40724 = n16676 & n39612;
  assign n40725 = ~n40723 & ~n40724;
  assign n40726 = ~n40722 & n40725;
  assign n40727 = ~n16079 & n40726;
  assign n40728 = ~n39991 & n40726;
  assign n40729 = ~n40727 & ~n40728;
  assign n40730 = ~n40721 & n40726;
  assign n40731 = pi17  & ~n58601;
  assign n40732 = ~pi17  & n58601;
  assign n40733 = ~n40731 & ~n40732;
  assign n40734 = n40417 & n58552;
  assign n40735 = ~n58552 & ~n40425;
  assign n40736 = ~n40417 & ~n40425;
  assign n40737 = ~n40735 & ~n40736;
  assign n40738 = ~n40425 & ~n40734;
  assign n40739 = ~n40733 & ~n58602;
  assign n40740 = n16079 & n40071;
  assign n40741 = n16696 & n39612;
  assign n40742 = n54886 & n39618;
  assign n40743 = n16676 & n39615;
  assign n40744 = ~n40742 & ~n40743;
  assign n40745 = ~n40741 & n40744;
  assign n40746 = ~n40740 & n40745;
  assign n40747 = pi17  & ~n40746;
  assign n40748 = ~n40746 & ~n40747;
  assign n40749 = ~pi17  & ~n40746;
  assign n40750 = pi17  & ~n40747;
  assign n40751 = pi17  & n40746;
  assign n40752 = ~n58603 & ~n58604;
  assign n40753 = pi20  & ~n58545;
  assign n40754 = ~n58546 & ~n40753;
  assign n40755 = n58546 & n40753;
  assign n40756 = ~n58545 & n40401;
  assign n40757 = ~n58547 & ~n40756;
  assign n40758 = ~n40754 & ~n40755;
  assign n40759 = ~n40752 & n58605;
  assign n40760 = n16079 & n40093;
  assign n40761 = n16696 & n39615;
  assign n40762 = n54886 & n39621;
  assign n40763 = n16676 & n39618;
  assign n40764 = ~n40762 & ~n40763;
  assign n40765 = ~n40761 & n40764;
  assign n40766 = ~n16079 & n40765;
  assign n40767 = ~n40093 & n40765;
  assign n40768 = ~n40766 & ~n40767;
  assign n40769 = ~n40760 & n40765;
  assign n40770 = pi17  & ~n58606;
  assign n40771 = ~pi17  & n58606;
  assign n40772 = ~n40770 & ~n40771;
  assign n40773 = pi20  & n40381;
  assign n40774 = ~n40380 & n40773;
  assign n40775 = n40380 & ~n40773;
  assign n40776 = ~n40382 & n40386;
  assign n40777 = ~n58545 & ~n40776;
  assign n40778 = ~n40774 & ~n40775;
  assign n40779 = ~n40772 & n58607;
  assign n40780 = n16079 & ~n40023;
  assign n40781 = n16676 & ~n58457;
  assign n40782 = n16696 & n39626;
  assign n40783 = ~n40781 & ~n40782;
  assign n40784 = ~n40780 & n40783;
  assign n40785 = n54883 & ~n58457;
  assign n40786 = pi17  & ~n40785;
  assign n40787 = pi17  & ~n40784;
  assign n40788 = pi17  & ~n40787;
  assign n40789 = ~n40784 & ~n40787;
  assign n40790 = ~n40788 & ~n40789;
  assign n40791 = n40786 & ~n40790;
  assign n40792 = n40784 & n40786;
  assign n40793 = n16079 & ~n40039;
  assign n40794 = n16696 & n39621;
  assign n40795 = n54886 & ~n58457;
  assign n40796 = n16676 & n39626;
  assign n40797 = ~n40795 & ~n40796;
  assign n40798 = ~n40794 & n40797;
  assign n40799 = ~n16079 & n40798;
  assign n40800 = n40039 & n40798;
  assign n40801 = ~n40799 & ~n40800;
  assign n40802 = ~n40793 & n40798;
  assign n40803 = pi17  & ~n58609;
  assign n40804 = ~pi17  & n58609;
  assign n40805 = ~n40803 & ~n40804;
  assign n40806 = n58608 & ~n40805;
  assign n40807 = n58608 & ~n58609;
  assign n40808 = n40381 & n58610;
  assign n40809 = n16079 & n40006;
  assign n40810 = n16696 & n39618;
  assign n40811 = n54886 & n39626;
  assign n40812 = n16676 & n39621;
  assign n40813 = ~n40811 & ~n40812;
  assign n40814 = ~n40810 & n40813;
  assign n40815 = ~n40809 & n40814;
  assign n40816 = pi17  & ~n40815;
  assign n40817 = pi17  & ~n40816;
  assign n40818 = pi17  & n40815;
  assign n40819 = ~n40815 & ~n40816;
  assign n40820 = ~pi17  & ~n40815;
  assign n40821 = ~n58611 & ~n58612;
  assign n40822 = ~n40381 & ~n58610;
  assign n40823 = n58610 & ~n40808;
  assign n40824 = ~n40381 & n58610;
  assign n40825 = n40381 & ~n40808;
  assign n40826 = n40381 & ~n58610;
  assign n40827 = ~n58613 & ~n58614;
  assign n40828 = ~n40808 & ~n40822;
  assign n40829 = ~n40821 & ~n58615;
  assign n40830 = ~n40808 & ~n40829;
  assign n40831 = n40772 & ~n58607;
  assign n40832 = ~n40779 & ~n40831;
  assign n40833 = ~n40830 & n40832;
  assign n40834 = ~n40779 & ~n40833;
  assign n40835 = n40752 & ~n58605;
  assign n40836 = ~n40752 & ~n40759;
  assign n40837 = ~n40752 & ~n58605;
  assign n40838 = n58605 & ~n40759;
  assign n40839 = n40752 & n58605;
  assign n40840 = ~n58616 & ~n58617;
  assign n40841 = ~n40759 & ~n40835;
  assign n40842 = ~n40834 & ~n58618;
  assign n40843 = ~n40759 & ~n40842;
  assign n40844 = n40733 & n58602;
  assign n40845 = ~n40739 & ~n40844;
  assign n40846 = ~n40843 & n40845;
  assign n40847 = ~n40739 & ~n40846;
  assign n40848 = n40717 & ~n40719;
  assign n40849 = ~n40717 & ~n40720;
  assign n40850 = ~n40717 & ~n40719;
  assign n40851 = n40719 & ~n40720;
  assign n40852 = n40717 & n40719;
  assign n40853 = ~n58619 & ~n58620;
  assign n40854 = ~n40720 & ~n40848;
  assign n40855 = ~n40847 & ~n58621;
  assign n40856 = ~n40720 & ~n40855;
  assign n40857 = ~n40690 & n40703;
  assign n40858 = n40690 & ~n40704;
  assign n40859 = n40690 & n40703;
  assign n40860 = ~n40703 & ~n40704;
  assign n40861 = ~n40690 & ~n40703;
  assign n40862 = ~n58622 & ~n58623;
  assign n40863 = ~n40704 & ~n40857;
  assign n40864 = ~n40856 & ~n58624;
  assign n40865 = ~n40704 & ~n40864;
  assign n40866 = ~n40674 & n40687;
  assign n40867 = n40674 & ~n40688;
  assign n40868 = n40674 & n40687;
  assign n40869 = ~n40687 & ~n40688;
  assign n40870 = ~n40674 & ~n40687;
  assign n40871 = ~n58625 & ~n58626;
  assign n40872 = ~n40688 & ~n40866;
  assign n40873 = ~n40865 & ~n58627;
  assign n40874 = ~n40688 & ~n40873;
  assign n40875 = ~n40658 & n40671;
  assign n40876 = ~n40672 & ~n40875;
  assign n40877 = ~n40874 & n40876;
  assign n40878 = ~n40672 & ~n40877;
  assign n40879 = n40648 & n58595;
  assign n40880 = ~n40648 & ~n40656;
  assign n40881 = ~n58595 & ~n40656;
  assign n40882 = ~n40880 & ~n40881;
  assign n40883 = ~n40656 & ~n40879;
  assign n40884 = ~n40878 & ~n58628;
  assign n40885 = ~n40656 & ~n40884;
  assign n40886 = n40629 & n58590;
  assign n40887 = ~n40629 & ~n40635;
  assign n40888 = ~n40629 & n58590;
  assign n40889 = ~n58590 & ~n40635;
  assign n40890 = n40629 & ~n58590;
  assign n40891 = ~n58629 & ~n58630;
  assign n40892 = ~n40635 & ~n40886;
  assign n40893 = ~n40885 & ~n58631;
  assign n40894 = ~n40635 & ~n40893;
  assign n40895 = n40611 & ~n40613;
  assign n40896 = ~n40611 & ~n40614;
  assign n40897 = ~n40611 & ~n40613;
  assign n40898 = n40613 & ~n40614;
  assign n40899 = n40611 & n40613;
  assign n40900 = ~n58632 & ~n58633;
  assign n40901 = ~n40614 & ~n40895;
  assign n40902 = ~n40894 & ~n58634;
  assign n40903 = ~n40614 & ~n40902;
  assign n40904 = ~n40574 & n40592;
  assign n40905 = n40574 & ~n40593;
  assign n40906 = n40574 & n40592;
  assign n40907 = ~n40592 & ~n40593;
  assign n40908 = ~n40574 & ~n40592;
  assign n40909 = ~n58635 & ~n58636;
  assign n40910 = ~n40593 & ~n40904;
  assign n40911 = ~n40903 & ~n58637;
  assign n40912 = ~n40593 & ~n40911;
  assign n40913 = ~n40566 & ~n40572;
  assign n40914 = n14413 & n40616;
  assign n40915 = n15921 & n39591;
  assign n40916 = n54719 & n39597;
  assign n40917 = n15901 & n39594;
  assign n40918 = ~n40916 & ~n40917;
  assign n40919 = ~n40915 & n40918;
  assign n40920 = ~n40914 & n40919;
  assign n40921 = pi20  & ~n40920;
  assign n40922 = ~n40920 & ~n40921;
  assign n40923 = ~pi20  & ~n40920;
  assign n40924 = pi20  & ~n40921;
  assign n40925 = pi20  & n40920;
  assign n40926 = ~n58638 & ~n58639;
  assign n40927 = ~n40550 & ~n40558;
  assign n40928 = ~n40526 & ~n40534;
  assign n40929 = n123 & n39991;
  assign n40930 = n128 & n39609;
  assign n40931 = n53444 & n39615;
  assign n40932 = n127 & n39612;
  assign n40933 = ~n40931 & ~n40932;
  assign n40934 = ~n40930 & n40933;
  assign n40935 = ~n40929 & n40934;
  assign n40936 = pi26  & ~n40935;
  assign n40937 = ~n40935 & ~n40936;
  assign n40938 = ~pi26  & ~n40935;
  assign n40939 = pi26  & ~n40936;
  assign n40940 = pi26  & n40935;
  assign n40941 = ~n58640 & ~n58641;
  assign n40942 = n11279 & n40006;
  assign n40943 = n12584 & n39618;
  assign n40944 = n54410 & n39626;
  assign n40945 = n11267 & n39621;
  assign n40946 = ~n40944 & ~n40945;
  assign n40947 = ~n40943 & n40946;
  assign n40948 = ~n40942 & n40947;
  assign n40949 = pi29  & ~n40948;
  assign n40950 = ~n40948 & ~n40949;
  assign n40951 = ~pi29  & ~n40948;
  assign n40952 = pi29  & ~n40949;
  assign n40953 = pi29  & n40948;
  assign n40954 = ~n58642 & ~n58643;
  assign n40955 = ~n94 & ~n58457;
  assign n40956 = n58570 & n40955;
  assign n40957 = ~n58570 & ~n40955;
  assign n40958 = n58570 & ~n40955;
  assign n40959 = ~n58570 & n40955;
  assign n40960 = ~n40958 & ~n40959;
  assign n40961 = ~n40956 & ~n40957;
  assign n40962 = ~n40954 & ~n58644;
  assign n40963 = n40954 & n58644;
  assign n40964 = ~n40962 & ~n40963;
  assign n40965 = ~n40941 & n40964;
  assign n40966 = n40941 & ~n40964;
  assign n40967 = ~n40941 & ~n40965;
  assign n40968 = ~n40941 & ~n40964;
  assign n40969 = n40964 & ~n40965;
  assign n40970 = n40941 & n40964;
  assign n40971 = ~n58645 & ~n58646;
  assign n40972 = ~n40965 & ~n40966;
  assign n40973 = ~n40928 & ~n58647;
  assign n40974 = n40928 & n58647;
  assign n40975 = ~n40973 & ~n40974;
  assign n40976 = n90 & ~n58533;
  assign n40977 = n14236 & n39600;
  assign n40978 = n54667 & n39606;
  assign n40979 = n14210 & n39603;
  assign n40980 = ~n40978 & ~n40979;
  assign n40981 = ~n40977 & n40980;
  assign n40982 = ~n90 & n40981;
  assign n40983 = n58533 & n40981;
  assign n40984 = ~n40982 & ~n40983;
  assign n40985 = ~n40976 & n40981;
  assign n40986 = pi23  & ~n58648;
  assign n40987 = ~pi23  & n58648;
  assign n40988 = ~n40986 & ~n40987;
  assign n40989 = n40975 & ~n40988;
  assign n40990 = ~n40975 & n40988;
  assign n40991 = ~n40989 & ~n40990;
  assign n40992 = ~n40927 & n40991;
  assign n40993 = n40927 & ~n40991;
  assign n40994 = ~n40992 & ~n40993;
  assign n40995 = ~n40926 & n40994;
  assign n40996 = n40926 & ~n40994;
  assign n40997 = ~n40926 & ~n40995;
  assign n40998 = ~n40926 & ~n40994;
  assign n40999 = n40994 & ~n40995;
  assign n41000 = n40926 & n40994;
  assign n41001 = ~n58649 & ~n58650;
  assign n41002 = ~n40995 & ~n40996;
  assign n41003 = ~n40913 & ~n58651;
  assign n41004 = n40913 & n58651;
  assign n41005 = ~n41003 & ~n41004;
  assign n41006 = n39689 & ~n39691;
  assign n41007 = ~n39692 & ~n41006;
  assign n41008 = n16079 & n41007;
  assign n41009 = n16696 & n39582;
  assign n41010 = n54886 & n39588;
  assign n41011 = n16676 & n39585;
  assign n41012 = ~n41010 & ~n41011;
  assign n41013 = ~n41009 & n41012;
  assign n41014 = ~n16079 & n41013;
  assign n41015 = ~n41007 & n41013;
  assign n41016 = ~n41014 & ~n41015;
  assign n41017 = ~n41008 & n41013;
  assign n41018 = pi17  & ~n58652;
  assign n41019 = ~pi17  & n58652;
  assign n41020 = ~n41018 & ~n41019;
  assign n41021 = n41005 & ~n41020;
  assign n41022 = ~n41005 & n41020;
  assign n41023 = ~n41021 & ~n41022;
  assign n41024 = ~n40912 & n41023;
  assign n41025 = n40912 & ~n41023;
  assign n41026 = ~n41024 & ~n41025;
  assign n41027 = ~n39989 & n41026;
  assign n41028 = n39699 & ~n39701;
  assign n41029 = ~n39699 & ~n58463;
  assign n41030 = ~n39700 & n39705;
  assign n41031 = ~n41029 & ~n41030;
  assign n41032 = ~n58463 & ~n41028;
  assign n41033 = n17265 & ~n58653;
  assign n41034 = n18588 & n39576;
  assign n41035 = n55041 & n39582;
  assign n41036 = n18556 & n39579;
  assign n41037 = ~n41035 & ~n41036;
  assign n41038 = ~n41034 & n41037;
  assign n41039 = ~n41033 & n41038;
  assign n41040 = pi14  & ~n41039;
  assign n41041 = ~n41039 & ~n41040;
  assign n41042 = ~pi14  & ~n41039;
  assign n41043 = pi14  & ~n41040;
  assign n41044 = pi14  & n41039;
  assign n41045 = ~n58654 & ~n58655;
  assign n41046 = n40903 & n58637;
  assign n41047 = ~n40903 & ~n40911;
  assign n41048 = ~n58637 & ~n40911;
  assign n41049 = ~n41047 & ~n41048;
  assign n41050 = ~n40911 & ~n41046;
  assign n41051 = ~n41045 & ~n58656;
  assign n41052 = n40894 & n58634;
  assign n41053 = ~n40902 & ~n41052;
  assign n41054 = n39693 & ~n39695;
  assign n41055 = ~n39693 & ~n58462;
  assign n41056 = ~n39694 & n39699;
  assign n41057 = ~n41055 & ~n41056;
  assign n41058 = ~n58462 & ~n41054;
  assign n41059 = n17265 & ~n58657;
  assign n41060 = n18588 & n39579;
  assign n41061 = n55041 & n39585;
  assign n41062 = n18556 & n39582;
  assign n41063 = ~n41061 & ~n41062;
  assign n41064 = ~n41060 & n41063;
  assign n41065 = ~n17265 & n41064;
  assign n41066 = n58657 & n41064;
  assign n41067 = ~n41065 & ~n41066;
  assign n41068 = ~n41059 & n41064;
  assign n41069 = pi14  & ~n58658;
  assign n41070 = ~pi14  & n58658;
  assign n41071 = ~n41069 & ~n41070;
  assign n41072 = n41053 & ~n41071;
  assign n41073 = n40885 & n58631;
  assign n41074 = ~n40893 & ~n41073;
  assign n41075 = n17265 & n41007;
  assign n41076 = n18588 & n39582;
  assign n41077 = n55041 & n39588;
  assign n41078 = n18556 & n39585;
  assign n41079 = ~n41077 & ~n41078;
  assign n41080 = ~n41076 & n41079;
  assign n41081 = ~n17265 & n41080;
  assign n41082 = ~n41007 & n41080;
  assign n41083 = ~n41081 & ~n41082;
  assign n41084 = ~n41075 & n41080;
  assign n41085 = pi14  & ~n58659;
  assign n41086 = ~pi14  & n58659;
  assign n41087 = ~n41085 & ~n41086;
  assign n41088 = n41074 & ~n41087;
  assign n41089 = n40878 & n58628;
  assign n41090 = ~n40884 & ~n41089;
  assign n41091 = n17265 & ~n58583;
  assign n41092 = n18588 & n39585;
  assign n41093 = n55041 & n39591;
  assign n41094 = n18556 & n39588;
  assign n41095 = ~n41093 & ~n41094;
  assign n41096 = ~n41092 & n41095;
  assign n41097 = ~n17265 & n41096;
  assign n41098 = n58583 & n41096;
  assign n41099 = ~n41097 & ~n41098;
  assign n41100 = ~n41091 & n41096;
  assign n41101 = pi14  & ~n58660;
  assign n41102 = ~pi14  & n58660;
  assign n41103 = ~n41101 & ~n41102;
  assign n41104 = n41090 & ~n41103;
  assign n41105 = n17265 & ~n58585;
  assign n41106 = n18588 & n39588;
  assign n41107 = n55041 & n39594;
  assign n41108 = n18556 & n39591;
  assign n41109 = ~n41107 & ~n41108;
  assign n41110 = ~n41106 & n41109;
  assign n41111 = ~n41105 & n41110;
  assign n41112 = pi14  & ~n41111;
  assign n41113 = ~n41111 & ~n41112;
  assign n41114 = ~pi14  & ~n41111;
  assign n41115 = pi14  & ~n41112;
  assign n41116 = pi14  & n41111;
  assign n41117 = ~n58661 & ~n58662;
  assign n41118 = n40874 & ~n40876;
  assign n41119 = ~n40877 & ~n41118;
  assign n41120 = ~n41117 & n41119;
  assign n41121 = n17265 & n40616;
  assign n41122 = n18588 & n39591;
  assign n41123 = n55041 & n39597;
  assign n41124 = n18556 & n39594;
  assign n41125 = ~n41123 & ~n41124;
  assign n41126 = ~n41122 & n41125;
  assign n41127 = ~n41121 & n41126;
  assign n41128 = pi14  & ~n41127;
  assign n41129 = ~n41127 & ~n41128;
  assign n41130 = ~pi14  & ~n41127;
  assign n41131 = pi14  & ~n41128;
  assign n41132 = pi14  & n41127;
  assign n41133 = ~n58663 & ~n58664;
  assign n41134 = n40865 & n58627;
  assign n41135 = ~n40865 & ~n40873;
  assign n41136 = ~n58627 & ~n40873;
  assign n41137 = ~n41135 & ~n41136;
  assign n41138 = ~n40873 & ~n41134;
  assign n41139 = ~n41133 & ~n58665;
  assign n41140 = n17265 & n40476;
  assign n41141 = n18588 & n39594;
  assign n41142 = n55041 & n39600;
  assign n41143 = n18556 & n39597;
  assign n41144 = ~n41142 & ~n41143;
  assign n41145 = ~n41141 & n41144;
  assign n41146 = ~n41140 & n41145;
  assign n41147 = pi14  & ~n41146;
  assign n41148 = ~n41146 & ~n41147;
  assign n41149 = ~pi14  & ~n41146;
  assign n41150 = pi14  & ~n41147;
  assign n41151 = pi14  & n41146;
  assign n41152 = ~n58666 & ~n58667;
  assign n41153 = n40856 & n58624;
  assign n41154 = ~n40856 & ~n40864;
  assign n41155 = ~n40856 & n58624;
  assign n41156 = ~n58624 & ~n40864;
  assign n41157 = n40856 & ~n58624;
  assign n41158 = ~n58668 & ~n58669;
  assign n41159 = ~n40864 & ~n41153;
  assign n41160 = ~n41152 & ~n58670;
  assign n41161 = n40847 & n58621;
  assign n41162 = ~n40855 & ~n41161;
  assign n41163 = n17265 & n40247;
  assign n41164 = n18588 & n39597;
  assign n41165 = n55041 & n39603;
  assign n41166 = n18556 & n39600;
  assign n41167 = ~n41165 & ~n41166;
  assign n41168 = ~n41164 & n41167;
  assign n41169 = ~n17265 & n41168;
  assign n41170 = ~n40247 & n41168;
  assign n41171 = ~n41169 & ~n41170;
  assign n41172 = ~n41163 & n41168;
  assign n41173 = pi14  & ~n58671;
  assign n41174 = ~pi14  & n58671;
  assign n41175 = ~n41173 & ~n41174;
  assign n41176 = n41162 & ~n41175;
  assign n41177 = n40843 & ~n40845;
  assign n41178 = ~n40846 & ~n41177;
  assign n41179 = n17265 & ~n58533;
  assign n41180 = n18588 & n39600;
  assign n41181 = n55041 & n39606;
  assign n41182 = n18556 & n39603;
  assign n41183 = ~n41181 & ~n41182;
  assign n41184 = ~n41180 & n41183;
  assign n41185 = ~n17265 & n41184;
  assign n41186 = n58533 & n41184;
  assign n41187 = ~n41185 & ~n41186;
  assign n41188 = ~n41179 & n41184;
  assign n41189 = pi14  & ~n58672;
  assign n41190 = ~pi14  & n58672;
  assign n41191 = ~n41189 & ~n41190;
  assign n41192 = n41178 & ~n41191;
  assign n41193 = n40834 & n58618;
  assign n41194 = ~n40842 & ~n41193;
  assign n41195 = n17265 & n40286;
  assign n41196 = n18588 & n39603;
  assign n41197 = n55041 & n39609;
  assign n41198 = n18556 & n39606;
  assign n41199 = ~n41197 & ~n41198;
  assign n41200 = ~n41196 & n41199;
  assign n41201 = ~n17265 & n41200;
  assign n41202 = ~n40286 & n41200;
  assign n41203 = ~n41201 & ~n41202;
  assign n41204 = ~n41195 & n41200;
  assign n41205 = pi14  & ~n58673;
  assign n41206 = ~pi14  & n58673;
  assign n41207 = ~n41205 & ~n41206;
  assign n41208 = n41194 & ~n41207;
  assign n41209 = n17265 & n40183;
  assign n41210 = n18588 & n39606;
  assign n41211 = n55041 & n39612;
  assign n41212 = n18556 & n39609;
  assign n41213 = ~n41211 & ~n41212;
  assign n41214 = ~n41210 & n41213;
  assign n41215 = ~n41209 & n41214;
  assign n41216 = pi14  & ~n41215;
  assign n41217 = ~n41215 & ~n41216;
  assign n41218 = ~pi14  & ~n41215;
  assign n41219 = pi14  & ~n41216;
  assign n41220 = pi14  & n41215;
  assign n41221 = ~n58674 & ~n58675;
  assign n41222 = n40830 & ~n40832;
  assign n41223 = ~n40833 & ~n41222;
  assign n41224 = ~n41221 & n41223;
  assign n41225 = n17265 & n39991;
  assign n41226 = n18588 & n39609;
  assign n41227 = n55041 & n39615;
  assign n41228 = n18556 & n39612;
  assign n41229 = ~n41227 & ~n41228;
  assign n41230 = ~n41226 & n41229;
  assign n41231 = ~n17265 & n41230;
  assign n41232 = ~n39991 & n41230;
  assign n41233 = ~n41231 & ~n41232;
  assign n41234 = ~n41225 & n41230;
  assign n41235 = pi14  & ~n58676;
  assign n41236 = ~pi14  & n58676;
  assign n41237 = ~n41235 & ~n41236;
  assign n41238 = n40821 & n58615;
  assign n41239 = ~n58615 & ~n40829;
  assign n41240 = ~n40821 & ~n40829;
  assign n41241 = ~n41239 & ~n41240;
  assign n41242 = ~n40829 & ~n41238;
  assign n41243 = ~n41237 & ~n58677;
  assign n41244 = n17265 & n40071;
  assign n41245 = n18588 & n39612;
  assign n41246 = n55041 & n39618;
  assign n41247 = n18556 & n39615;
  assign n41248 = ~n41246 & ~n41247;
  assign n41249 = ~n41245 & n41248;
  assign n41250 = ~n41244 & n41249;
  assign n41251 = pi14  & ~n41250;
  assign n41252 = ~n41250 & ~n41251;
  assign n41253 = ~pi14  & ~n41250;
  assign n41254 = pi14  & ~n41251;
  assign n41255 = pi14  & n41250;
  assign n41256 = ~n58678 & ~n58679;
  assign n41257 = pi17  & ~n58608;
  assign n41258 = ~n58609 & ~n41257;
  assign n41259 = n58609 & n41257;
  assign n41260 = ~n58608 & n40805;
  assign n41261 = ~n58610 & ~n41260;
  assign n41262 = ~n41258 & ~n41259;
  assign n41263 = ~n41256 & n58680;
  assign n41264 = n17265 & n40093;
  assign n41265 = n18588 & n39615;
  assign n41266 = n55041 & n39621;
  assign n41267 = n18556 & n39618;
  assign n41268 = ~n41266 & ~n41267;
  assign n41269 = ~n41265 & n41268;
  assign n41270 = ~n17265 & n41269;
  assign n41271 = ~n40093 & n41269;
  assign n41272 = ~n41270 & ~n41271;
  assign n41273 = ~n41264 & n41269;
  assign n41274 = pi14  & ~n58681;
  assign n41275 = ~pi14  & n58681;
  assign n41276 = ~n41274 & ~n41275;
  assign n41277 = pi17  & n40785;
  assign n41278 = ~n40784 & n41277;
  assign n41279 = n40784 & ~n41277;
  assign n41280 = ~n40786 & n40790;
  assign n41281 = ~n58608 & ~n41280;
  assign n41282 = ~n41278 & ~n41279;
  assign n41283 = ~n41276 & n58682;
  assign n41284 = n17265 & ~n40023;
  assign n41285 = n18556 & ~n58457;
  assign n41286 = n18588 & n39626;
  assign n41287 = ~n41285 & ~n41286;
  assign n41288 = ~n41284 & n41287;
  assign n41289 = n55039 & ~n58457;
  assign n41290 = pi14  & ~n41289;
  assign n41291 = pi14  & ~n41288;
  assign n41292 = pi14  & ~n41291;
  assign n41293 = ~n41288 & ~n41291;
  assign n41294 = ~n41292 & ~n41293;
  assign n41295 = n41290 & ~n41294;
  assign n41296 = n41288 & n41290;
  assign n41297 = n17265 & ~n40039;
  assign n41298 = n18588 & n39621;
  assign n41299 = n55041 & ~n58457;
  assign n41300 = n18556 & n39626;
  assign n41301 = ~n41299 & ~n41300;
  assign n41302 = ~n41298 & n41301;
  assign n41303 = ~n17265 & n41302;
  assign n41304 = n40039 & n41302;
  assign n41305 = ~n41303 & ~n41304;
  assign n41306 = ~n41297 & n41302;
  assign n41307 = pi14  & ~n58684;
  assign n41308 = ~pi14  & n58684;
  assign n41309 = ~n41307 & ~n41308;
  assign n41310 = n58683 & ~n41309;
  assign n41311 = n58683 & ~n58684;
  assign n41312 = n40785 & n58685;
  assign n41313 = n17265 & n40006;
  assign n41314 = n18588 & n39618;
  assign n41315 = n55041 & n39626;
  assign n41316 = n18556 & n39621;
  assign n41317 = ~n41315 & ~n41316;
  assign n41318 = ~n41314 & n41317;
  assign n41319 = ~n41313 & n41318;
  assign n41320 = pi14  & ~n41319;
  assign n41321 = pi14  & ~n41320;
  assign n41322 = pi14  & n41319;
  assign n41323 = ~n41319 & ~n41320;
  assign n41324 = ~pi14  & ~n41319;
  assign n41325 = ~n58686 & ~n58687;
  assign n41326 = ~n40785 & ~n58685;
  assign n41327 = n58685 & ~n41312;
  assign n41328 = ~n40785 & n58685;
  assign n41329 = n40785 & ~n41312;
  assign n41330 = n40785 & ~n58685;
  assign n41331 = ~n58688 & ~n58689;
  assign n41332 = ~n41312 & ~n41326;
  assign n41333 = ~n41325 & ~n58690;
  assign n41334 = ~n41312 & ~n41333;
  assign n41335 = n41276 & ~n58682;
  assign n41336 = ~n41283 & ~n41335;
  assign n41337 = ~n41334 & n41336;
  assign n41338 = ~n41283 & ~n41337;
  assign n41339 = n41256 & ~n58680;
  assign n41340 = ~n41256 & ~n41263;
  assign n41341 = ~n41256 & ~n58680;
  assign n41342 = n58680 & ~n41263;
  assign n41343 = n41256 & n58680;
  assign n41344 = ~n58691 & ~n58692;
  assign n41345 = ~n41263 & ~n41339;
  assign n41346 = ~n41338 & ~n58693;
  assign n41347 = ~n41263 & ~n41346;
  assign n41348 = n41237 & n58677;
  assign n41349 = ~n41243 & ~n41348;
  assign n41350 = ~n41347 & n41349;
  assign n41351 = ~n41243 & ~n41350;
  assign n41352 = n41221 & ~n41223;
  assign n41353 = ~n41221 & ~n41224;
  assign n41354 = ~n41221 & ~n41223;
  assign n41355 = n41223 & ~n41224;
  assign n41356 = n41221 & n41223;
  assign n41357 = ~n58694 & ~n58695;
  assign n41358 = ~n41224 & ~n41352;
  assign n41359 = ~n41351 & ~n58696;
  assign n41360 = ~n41224 & ~n41359;
  assign n41361 = ~n41194 & n41207;
  assign n41362 = n41194 & ~n41208;
  assign n41363 = n41194 & n41207;
  assign n41364 = ~n41207 & ~n41208;
  assign n41365 = ~n41194 & ~n41207;
  assign n41366 = ~n58697 & ~n58698;
  assign n41367 = ~n41208 & ~n41361;
  assign n41368 = ~n41360 & ~n58699;
  assign n41369 = ~n41208 & ~n41368;
  assign n41370 = ~n41178 & n41191;
  assign n41371 = n41178 & ~n41192;
  assign n41372 = n41178 & n41191;
  assign n41373 = ~n41191 & ~n41192;
  assign n41374 = ~n41178 & ~n41191;
  assign n41375 = ~n58700 & ~n58701;
  assign n41376 = ~n41192 & ~n41370;
  assign n41377 = ~n41369 & ~n58702;
  assign n41378 = ~n41192 & ~n41377;
  assign n41379 = ~n41162 & n41175;
  assign n41380 = ~n41176 & ~n41379;
  assign n41381 = ~n41378 & n41380;
  assign n41382 = ~n41176 & ~n41381;
  assign n41383 = n41152 & n58670;
  assign n41384 = ~n41152 & ~n41160;
  assign n41385 = ~n58670 & ~n41160;
  assign n41386 = ~n41384 & ~n41385;
  assign n41387 = ~n41160 & ~n41383;
  assign n41388 = ~n41382 & ~n58703;
  assign n41389 = ~n41160 & ~n41388;
  assign n41390 = n41133 & n58665;
  assign n41391 = ~n41133 & ~n41139;
  assign n41392 = ~n41133 & n58665;
  assign n41393 = ~n58665 & ~n41139;
  assign n41394 = n41133 & ~n58665;
  assign n41395 = ~n58704 & ~n58705;
  assign n41396 = ~n41139 & ~n41390;
  assign n41397 = ~n41389 & ~n58706;
  assign n41398 = ~n41139 & ~n41397;
  assign n41399 = n41117 & ~n41119;
  assign n41400 = ~n41117 & ~n41120;
  assign n41401 = ~n41117 & ~n41119;
  assign n41402 = n41119 & ~n41120;
  assign n41403 = n41117 & n41119;
  assign n41404 = ~n58707 & ~n58708;
  assign n41405 = ~n41120 & ~n41399;
  assign n41406 = ~n41398 & ~n58709;
  assign n41407 = ~n41120 & ~n41406;
  assign n41408 = ~n41090 & n41103;
  assign n41409 = n41090 & ~n41104;
  assign n41410 = n41090 & n41103;
  assign n41411 = ~n41103 & ~n41104;
  assign n41412 = ~n41090 & ~n41103;
  assign n41413 = ~n58710 & ~n58711;
  assign n41414 = ~n41104 & ~n41408;
  assign n41415 = ~n41407 & ~n58712;
  assign n41416 = ~n41104 & ~n41415;
  assign n41417 = ~n41074 & n41087;
  assign n41418 = n41074 & ~n41088;
  assign n41419 = n41074 & n41087;
  assign n41420 = ~n41087 & ~n41088;
  assign n41421 = ~n41074 & ~n41087;
  assign n41422 = ~n58713 & ~n58714;
  assign n41423 = ~n41088 & ~n41417;
  assign n41424 = ~n41416 & ~n58715;
  assign n41425 = ~n41088 & ~n41424;
  assign n41426 = ~n41053 & n41071;
  assign n41427 = ~n41072 & ~n41426;
  assign n41428 = ~n41425 & n41427;
  assign n41429 = ~n41072 & ~n41428;
  assign n41430 = n41045 & n58656;
  assign n41431 = ~n41045 & ~n41051;
  assign n41432 = ~n41045 & n58656;
  assign n41433 = ~n58656 & ~n41051;
  assign n41434 = n41045 & ~n58656;
  assign n41435 = ~n58716 & ~n58717;
  assign n41436 = ~n41051 & ~n41430;
  assign n41437 = ~n41429 & ~n58718;
  assign n41438 = ~n41051 & ~n41437;
  assign n41439 = n39989 & ~n41026;
  assign n41440 = ~n39989 & ~n41027;
  assign n41441 = ~n39989 & ~n41026;
  assign n41442 = n41026 & ~n41027;
  assign n41443 = n39989 & n41026;
  assign n41444 = ~n58719 & ~n58720;
  assign n41445 = ~n41027 & ~n41439;
  assign n41446 = ~n41438 & ~n58721;
  assign n41447 = ~n41027 & ~n41446;
  assign n41448 = ~n41021 & ~n41024;
  assign n41449 = n16079 & ~n58657;
  assign n41450 = n16696 & n39579;
  assign n41451 = n54886 & n39585;
  assign n41452 = n16676 & n39582;
  assign n41453 = ~n41451 & ~n41452;
  assign n41454 = ~n41450 & n41453;
  assign n41455 = ~n41449 & n41454;
  assign n41456 = pi17  & ~n41455;
  assign n41457 = ~n41455 & ~n41456;
  assign n41458 = ~pi17  & ~n41455;
  assign n41459 = pi17  & ~n41456;
  assign n41460 = pi17  & n41455;
  assign n41461 = ~n58722 & ~n58723;
  assign n41462 = ~n40995 & ~n41003;
  assign n41463 = ~n40989 & ~n40992;
  assign n41464 = n90 & n40247;
  assign n41465 = n14236 & n39597;
  assign n41466 = n54667 & n39603;
  assign n41467 = n14210 & n39600;
  assign n41468 = ~n41466 & ~n41467;
  assign n41469 = ~n41465 & n41468;
  assign n41470 = ~n41464 & n41469;
  assign n41471 = pi23  & ~n41470;
  assign n41472 = ~n41470 & ~n41471;
  assign n41473 = ~pi23  & ~n41470;
  assign n41474 = pi23  & ~n41471;
  assign n41475 = pi23  & n41470;
  assign n41476 = ~n58724 & ~n58725;
  assign n41477 = ~n40965 & ~n40973;
  assign n41478 = n123 & n40183;
  assign n41479 = n128 & n39606;
  assign n41480 = n53444 & n39612;
  assign n41481 = n127 & n39609;
  assign n41482 = ~n41480 & ~n41481;
  assign n41483 = ~n41479 & n41482;
  assign n41484 = ~n123 & n41483;
  assign n41485 = ~n40183 & n41483;
  assign n41486 = ~n41484 & ~n41485;
  assign n41487 = ~n41478 & n41483;
  assign n41488 = pi26  & ~n58726;
  assign n41489 = ~pi26  & n58726;
  assign n41490 = ~n41488 & ~n41489;
  assign n41491 = ~n40956 & ~n40962;
  assign n41492 = n11279 & n40093;
  assign n41493 = n12584 & n39615;
  assign n41494 = n54410 & n39621;
  assign n41495 = n11267 & n39618;
  assign n41496 = ~n41494 & ~n41495;
  assign n41497 = ~n41493 & n41496;
  assign n41498 = ~n41492 & n41497;
  assign n41499 = pi29  & ~n41498;
  assign n41500 = ~n41498 & ~n41499;
  assign n41501 = ~pi29  & ~n41498;
  assign n41502 = pi29  & ~n41499;
  assign n41503 = pi29  & n41498;
  assign n41504 = ~n58727 & ~n58728;
  assign n41505 = n1458 & n1760;
  assign n41506 = n14606 & n41505;
  assign n41507 = ~n219 & ~n560;
  assign n41508 = ~n219 & ~n460;
  assign n41509 = ~n560 & n41508;
  assign n41510 = ~n460 & n41507;
  assign n41511 = n3678 & n3715;
  assign n41512 = n4012 & n4258;
  assign n41513 = n41511 & n41512;
  assign n41514 = n58729 & n41513;
  assign n41515 = n1458 & n41511;
  assign n41516 = n4258 & n41515;
  assign n41517 = n462 & n41516;
  assign n41518 = ~n631 & n41517;
  assign n41519 = ~n219 & n41518;
  assign n41520 = ~n560 & n41519;
  assign n41521 = ~n554 & n41520;
  assign n41522 = ~n493 & n41521;
  assign n41523 = ~n1644 & n41522;
  assign n41524 = ~n465 & n41523;
  assign n41525 = n1760 & n41512;
  assign n41526 = ~n560 & ~n1644;
  assign n41527 = ~n460 & n41526;
  assign n41528 = ~n219 & ~n554;
  assign n41529 = n1458 & n41528;
  assign n41530 = n41511 & n41529;
  assign n41531 = n41527 & n41530;
  assign n41532 = n41525 & n41531;
  assign n41533 = n462 & n1458;
  assign n41534 = n3715 & n41533;
  assign n41535 = ~n554 & n4012;
  assign n41536 = ~n219 & ~n465;
  assign n41537 = n41526 & n41536;
  assign n41538 = n3678 & n4258;
  assign n41539 = n41537 & n41538;
  assign n41540 = n41535 & n41539;
  assign n41541 = n41534 & n41540;
  assign n41542 = n41506 & n41514;
  assign n41543 = ~n356 & ~n495;
  assign n41544 = ~n356 & ~n504;
  assign n41545 = ~n495 & n41544;
  assign n41546 = ~n504 & n41543;
  assign n41547 = n3536 & n3950;
  assign n41548 = n58731 & n41547;
  assign n41549 = n54181 & n18103;
  assign n41550 = n41548 & n41549;
  assign n41551 = n976 & n1670;
  assign n41552 = n2174 & n5873;
  assign n41553 = n41551 & n41552;
  assign n41554 = n53924 & n41553;
  assign n41555 = n57044 & n41554;
  assign n41556 = n58731 & n41552;
  assign n41557 = n41549 & n41556;
  assign n41558 = n41547 & n41551;
  assign n41559 = n53924 & n41558;
  assign n41560 = n57044 & n41559;
  assign n41561 = n41557 & n41560;
  assign n41562 = ~n504 & ~n1476;
  assign n41563 = n3950 & n41562;
  assign n41564 = n41551 & n41563;
  assign n41565 = ~n356 & ~n883;
  assign n41566 = ~n495 & n41565;
  assign n41567 = n54181 & n41566;
  assign n41568 = n41564 & n41567;
  assign n41569 = n3536 & n5873;
  assign n41570 = n18103 & n41569;
  assign n41571 = n53924 & n41570;
  assign n41572 = n57044 & n41571;
  assign n41573 = n41568 & n41572;
  assign n41574 = n41550 & n41555;
  assign n41575 = n58730 & n58732;
  assign n41576 = ~n591 & ~n663;
  assign n41577 = ~n344 & ~n511;
  assign n41578 = ~n344 & ~n591;
  assign n41579 = ~n511 & ~n663;
  assign n41580 = n41578 & n41579;
  assign n41581 = n41576 & n41577;
  assign n41582 = n53629 & n58733;
  assign n41583 = n54594 & n41582;
  assign n41584 = n5113 & n8793;
  assign n41585 = n10182 & n11829;
  assign n41586 = n41584 & n41585;
  assign n41587 = n276 & n2328;
  assign n41588 = n1716 & n3742;
  assign n41589 = n41587 & n41588;
  assign n41590 = n8793 & n10182;
  assign n41591 = n2328 & n11829;
  assign n41592 = n41590 & n41591;
  assign n41593 = n276 & n3742;
  assign n41594 = n1716 & n5113;
  assign n41595 = n3742 & n5113;
  assign n41596 = n276 & n1716;
  assign n41597 = n41595 & n41596;
  assign n41598 = n41593 & n41594;
  assign n41599 = n41592 & n58734;
  assign n41600 = n41586 & n41589;
  assign n41601 = n56678 & n58735;
  assign n41602 = n2328 & n53629;
  assign n41603 = n10182 & n41602;
  assign n41604 = n54594 & n41603;
  assign n41605 = n56678 & n41604;
  assign n41606 = n5113 & n41605;
  assign n41607 = n11829 & n41606;
  assign n41608 = n8793 & n41607;
  assign n41609 = n1716 & n41608;
  assign n41610 = n3742 & n41609;
  assign n41611 = n276 & n41610;
  assign n41612 = ~n663 & n41611;
  assign n41613 = ~n591 & n41612;
  assign n41614 = ~n511 & n41613;
  assign n41615 = ~n344 & n41614;
  assign n41616 = n41583 & n41601;
  assign n41617 = n57028 & n58736;
  assign n41618 = n4974 & n54181;
  assign n41619 = n53924 & n41618;
  assign n41620 = n57044 & n41619;
  assign n41621 = n58736 & n41620;
  assign n41622 = n58730 & n41621;
  assign n41623 = n57028 & n41622;
  assign n41624 = n976 & n41623;
  assign n41625 = n3536 & n41624;
  assign n41626 = n3950 & n41625;
  assign n41627 = n3062 & n41626;
  assign n41628 = n5873 & n41627;
  assign n41629 = n1670 & n41628;
  assign n41630 = ~n883 & n41629;
  assign n41631 = ~n1476 & n41630;
  assign n41632 = ~n495 & n41631;
  assign n41633 = ~n504 & n41632;
  assign n41634 = ~n356 & n41633;
  assign n41635 = n41575 & n41617;
  assign n41636 = n1576 & ~n40023;
  assign n41637 = n11215 & n39626;
  assign n41638 = n10564 & ~n58457;
  assign n41639 = ~n41637 & ~n41638;
  assign n41640 = ~n41636 & ~n41638;
  assign n41641 = ~n41637 & n41640;
  assign n41642 = ~n41636 & n41639;
  assign n41643 = ~n58737 & ~n58738;
  assign n41644 = n58737 & n58738;
  assign n41645 = ~n58737 & ~n41643;
  assign n41646 = ~n58737 & n58738;
  assign n41647 = ~n58738 & ~n41643;
  assign n41648 = n58737 & ~n58738;
  assign n41649 = ~n58739 & ~n58740;
  assign n41650 = ~n41643 & ~n41644;
  assign n41651 = ~n41504 & ~n58741;
  assign n41652 = n41504 & n58741;
  assign n41653 = ~n41504 & ~n41651;
  assign n41654 = ~n58741 & ~n41651;
  assign n41655 = ~n41653 & ~n41654;
  assign n41656 = ~n41651 & ~n41652;
  assign n41657 = ~n41491 & ~n58742;
  assign n41658 = n41491 & n58742;
  assign n41659 = ~n58742 & ~n41657;
  assign n41660 = ~n41491 & ~n41657;
  assign n41661 = ~n41659 & ~n41660;
  assign n41662 = ~n41657 & ~n41658;
  assign n41663 = ~n41490 & ~n58743;
  assign n41664 = n41490 & n58743;
  assign n41665 = ~n58743 & ~n41663;
  assign n41666 = n41490 & ~n58743;
  assign n41667 = ~n41490 & ~n41663;
  assign n41668 = ~n41490 & n58743;
  assign n41669 = ~n58744 & ~n58745;
  assign n41670 = ~n41663 & ~n41664;
  assign n41671 = ~n41477 & ~n58746;
  assign n41672 = n41477 & n58746;
  assign n41673 = ~n41477 & ~n41671;
  assign n41674 = ~n58746 & ~n41671;
  assign n41675 = ~n41673 & ~n41674;
  assign n41676 = ~n41671 & ~n41672;
  assign n41677 = ~n41476 & ~n58747;
  assign n41678 = n41476 & n58747;
  assign n41679 = ~n41476 & ~n41677;
  assign n41680 = ~n41476 & n58747;
  assign n41681 = ~n58747 & ~n41677;
  assign n41682 = n41476 & ~n58747;
  assign n41683 = ~n58748 & ~n58749;
  assign n41684 = ~n41677 & ~n41678;
  assign n41685 = n41463 & n58750;
  assign n41686 = ~n41463 & ~n58750;
  assign n41687 = ~n41685 & ~n41686;
  assign n41688 = n14413 & ~n58585;
  assign n41689 = n15921 & n39588;
  assign n41690 = n54719 & n39594;
  assign n41691 = n15901 & n39591;
  assign n41692 = ~n41690 & ~n41691;
  assign n41693 = ~n41689 & n41692;
  assign n41694 = ~n14413 & n41693;
  assign n41695 = n58585 & n41693;
  assign n41696 = ~n41694 & ~n41695;
  assign n41697 = ~n41688 & n41693;
  assign n41698 = pi20  & ~n58751;
  assign n41699 = ~pi20  & n58751;
  assign n41700 = ~n41698 & ~n41699;
  assign n41701 = n41687 & ~n41700;
  assign n41702 = ~n41687 & n41700;
  assign n41703 = n41687 & ~n41701;
  assign n41704 = n41687 & n41700;
  assign n41705 = ~n41700 & ~n41701;
  assign n41706 = ~n41687 & ~n41700;
  assign n41707 = ~n58752 & ~n58753;
  assign n41708 = ~n41701 & ~n41702;
  assign n41709 = ~n41462 & ~n58754;
  assign n41710 = n41462 & n58754;
  assign n41711 = ~n41462 & ~n41709;
  assign n41712 = ~n41462 & n58754;
  assign n41713 = ~n58754 & ~n41709;
  assign n41714 = n41462 & ~n58754;
  assign n41715 = ~n58755 & ~n58756;
  assign n41716 = ~n41709 & ~n41710;
  assign n41717 = ~n41461 & ~n58757;
  assign n41718 = n41461 & n58757;
  assign n41719 = ~n41461 & ~n41717;
  assign n41720 = ~n58757 & ~n41717;
  assign n41721 = ~n41719 & ~n41720;
  assign n41722 = ~n41717 & ~n41718;
  assign n41723 = ~n41448 & ~n58758;
  assign n41724 = n41448 & n58758;
  assign n41725 = ~n41723 & ~n41724;
  assign n41726 = n39709 & ~n39711;
  assign n41727 = ~n39709 & ~n58464;
  assign n41728 = ~n39710 & n39715;
  assign n41729 = ~n41727 & ~n41728;
  assign n41730 = ~n58464 & ~n41726;
  assign n41731 = n17265 & ~n58759;
  assign n41732 = n18588 & n39570;
  assign n41733 = n55041 & n39576;
  assign n41734 = n18556 & n39573;
  assign n41735 = ~n41733 & ~n41734;
  assign n41736 = ~n41732 & n41735;
  assign n41737 = ~n17265 & n41736;
  assign n41738 = n58759 & n41736;
  assign n41739 = ~n41737 & ~n41738;
  assign n41740 = ~n41731 & n41736;
  assign n41741 = pi14  & ~n58760;
  assign n41742 = ~pi14  & n58760;
  assign n41743 = ~n41741 & ~n41742;
  assign n41744 = n41725 & ~n41743;
  assign n41745 = ~n41725 & n41743;
  assign n41746 = n41725 & ~n41744;
  assign n41747 = n41725 & n41743;
  assign n41748 = ~n41743 & ~n41744;
  assign n41749 = ~n41725 & ~n41743;
  assign n41750 = ~n58761 & ~n58762;
  assign n41751 = ~n41744 & ~n41745;
  assign n41752 = ~n41447 & ~n58763;
  assign n41753 = n41447 & n58763;
  assign n41754 = ~n41447 & ~n41752;
  assign n41755 = ~n58763 & ~n41752;
  assign n41756 = ~n41754 & ~n41755;
  assign n41757 = ~n41752 & ~n41753;
  assign n41758 = ~n39974 & ~n58764;
  assign n41759 = n41438 & n58721;
  assign n41760 = ~n41446 & ~n41759;
  assign n41761 = n39721 & ~n39723;
  assign n41762 = ~n39724 & ~n41761;
  assign n41763 = n18846 & n41762;
  assign n41764 = n19541 & n39564;
  assign n41765 = n55247 & n39570;
  assign n41766 = n19509 & n39567;
  assign n41767 = ~n41765 & ~n41766;
  assign n41768 = ~n41764 & n41767;
  assign n41769 = ~n18846 & n41768;
  assign n41770 = ~n41762 & n41768;
  assign n41771 = ~n41769 & ~n41770;
  assign n41772 = ~n41763 & n41768;
  assign n41773 = pi11  & ~n58765;
  assign n41774 = ~pi11  & n58765;
  assign n41775 = ~n41773 & ~n41774;
  assign n41776 = n41760 & ~n41775;
  assign n41777 = n41429 & n58718;
  assign n41778 = ~n41437 & ~n41777;
  assign n41779 = n39715 & ~n39717;
  assign n41780 = ~n39715 & ~n58465;
  assign n41781 = ~n39716 & n39721;
  assign n41782 = ~n41780 & ~n41781;
  assign n41783 = ~n58465 & ~n41779;
  assign n41784 = n18846 & ~n58766;
  assign n41785 = n19541 & n39567;
  assign n41786 = n55247 & n39573;
  assign n41787 = n19509 & n39570;
  assign n41788 = ~n41786 & ~n41787;
  assign n41789 = ~n41785 & n41788;
  assign n41790 = ~n18846 & n41789;
  assign n41791 = n58766 & n41789;
  assign n41792 = ~n41790 & ~n41791;
  assign n41793 = ~n41784 & n41789;
  assign n41794 = pi11  & ~n58767;
  assign n41795 = ~pi11  & n58767;
  assign n41796 = ~n41794 & ~n41795;
  assign n41797 = n41778 & ~n41796;
  assign n41798 = n18846 & ~n58759;
  assign n41799 = n19541 & n39570;
  assign n41800 = n55247 & n39576;
  assign n41801 = n19509 & n39573;
  assign n41802 = ~n41800 & ~n41801;
  assign n41803 = ~n41799 & n41802;
  assign n41804 = ~n41798 & n41803;
  assign n41805 = pi11  & ~n41804;
  assign n41806 = ~n41804 & ~n41805;
  assign n41807 = ~pi11  & ~n41804;
  assign n41808 = pi11  & ~n41805;
  assign n41809 = pi11  & n41804;
  assign n41810 = ~n58768 & ~n58769;
  assign n41811 = n41425 & ~n41427;
  assign n41812 = ~n41428 & ~n41811;
  assign n41813 = ~n41810 & n41812;
  assign n41814 = n18846 & n39976;
  assign n41815 = n19541 & n39573;
  assign n41816 = n55247 & n39579;
  assign n41817 = n19509 & n39576;
  assign n41818 = ~n41816 & ~n41817;
  assign n41819 = ~n41815 & n41818;
  assign n41820 = ~n41814 & n41819;
  assign n41821 = pi11  & ~n41820;
  assign n41822 = ~n41820 & ~n41821;
  assign n41823 = ~pi11  & ~n41820;
  assign n41824 = pi11  & ~n41821;
  assign n41825 = pi11  & n41820;
  assign n41826 = ~n58770 & ~n58771;
  assign n41827 = n41416 & n58715;
  assign n41828 = ~n41416 & ~n41424;
  assign n41829 = ~n41416 & n58715;
  assign n41830 = ~n58715 & ~n41424;
  assign n41831 = n41416 & ~n58715;
  assign n41832 = ~n58772 & ~n58773;
  assign n41833 = ~n41424 & ~n41827;
  assign n41834 = ~n41826 & ~n58774;
  assign n41835 = n18846 & ~n58653;
  assign n41836 = n19541 & n39576;
  assign n41837 = n55247 & n39582;
  assign n41838 = n19509 & n39579;
  assign n41839 = ~n41837 & ~n41838;
  assign n41840 = ~n41836 & n41839;
  assign n41841 = ~n41835 & n41840;
  assign n41842 = pi11  & ~n41841;
  assign n41843 = ~n41841 & ~n41842;
  assign n41844 = ~pi11  & ~n41841;
  assign n41845 = pi11  & ~n41842;
  assign n41846 = pi11  & n41841;
  assign n41847 = ~n58775 & ~n58776;
  assign n41848 = n41407 & n58712;
  assign n41849 = ~n41407 & ~n41415;
  assign n41850 = ~n58712 & ~n41415;
  assign n41851 = ~n41849 & ~n41850;
  assign n41852 = ~n41415 & ~n41848;
  assign n41853 = ~n41847 & ~n58777;
  assign n41854 = n41398 & n58709;
  assign n41855 = ~n41406 & ~n41854;
  assign n41856 = n18846 & ~n58657;
  assign n41857 = n19541 & n39579;
  assign n41858 = n55247 & n39585;
  assign n41859 = n19509 & n39582;
  assign n41860 = ~n41858 & ~n41859;
  assign n41861 = ~n41857 & n41860;
  assign n41862 = ~n18846 & n41861;
  assign n41863 = n58657 & n41861;
  assign n41864 = ~n41862 & ~n41863;
  assign n41865 = ~n41856 & n41861;
  assign n41866 = pi11  & ~n58778;
  assign n41867 = ~pi11  & n58778;
  assign n41868 = ~n41866 & ~n41867;
  assign n41869 = n41855 & ~n41868;
  assign n41870 = n41389 & n58706;
  assign n41871 = ~n41397 & ~n41870;
  assign n41872 = n18846 & n41007;
  assign n41873 = n19541 & n39582;
  assign n41874 = n55247 & n39588;
  assign n41875 = n19509 & n39585;
  assign n41876 = ~n41874 & ~n41875;
  assign n41877 = ~n41873 & n41876;
  assign n41878 = ~n18846 & n41877;
  assign n41879 = ~n41007 & n41877;
  assign n41880 = ~n41878 & ~n41879;
  assign n41881 = ~n41872 & n41877;
  assign n41882 = pi11  & ~n58779;
  assign n41883 = ~pi11  & n58779;
  assign n41884 = ~n41882 & ~n41883;
  assign n41885 = n41871 & ~n41884;
  assign n41886 = n41382 & n58703;
  assign n41887 = ~n41388 & ~n41886;
  assign n41888 = n18846 & ~n58583;
  assign n41889 = n19541 & n39585;
  assign n41890 = n55247 & n39591;
  assign n41891 = n19509 & n39588;
  assign n41892 = ~n41890 & ~n41891;
  assign n41893 = ~n41889 & n41892;
  assign n41894 = ~n18846 & n41893;
  assign n41895 = n58583 & n41893;
  assign n41896 = ~n41894 & ~n41895;
  assign n41897 = ~n41888 & n41893;
  assign n41898 = pi11  & ~n58780;
  assign n41899 = ~pi11  & n58780;
  assign n41900 = ~n41898 & ~n41899;
  assign n41901 = n41887 & ~n41900;
  assign n41902 = n18846 & ~n58585;
  assign n41903 = n19541 & n39588;
  assign n41904 = n55247 & n39594;
  assign n41905 = n19509 & n39591;
  assign n41906 = ~n41904 & ~n41905;
  assign n41907 = ~n41903 & n41906;
  assign n41908 = ~n41902 & n41907;
  assign n41909 = pi11  & ~n41908;
  assign n41910 = ~n41908 & ~n41909;
  assign n41911 = ~pi11  & ~n41908;
  assign n41912 = pi11  & ~n41909;
  assign n41913 = pi11  & n41908;
  assign n41914 = ~n58781 & ~n58782;
  assign n41915 = n41378 & ~n41380;
  assign n41916 = ~n41381 & ~n41915;
  assign n41917 = ~n41914 & n41916;
  assign n41918 = n18846 & n40616;
  assign n41919 = n19541 & n39591;
  assign n41920 = n55247 & n39597;
  assign n41921 = n19509 & n39594;
  assign n41922 = ~n41920 & ~n41921;
  assign n41923 = ~n41919 & n41922;
  assign n41924 = ~n41918 & n41923;
  assign n41925 = pi11  & ~n41924;
  assign n41926 = ~n41924 & ~n41925;
  assign n41927 = ~pi11  & ~n41924;
  assign n41928 = pi11  & ~n41925;
  assign n41929 = pi11  & n41924;
  assign n41930 = ~n58783 & ~n58784;
  assign n41931 = n41369 & n58702;
  assign n41932 = ~n41369 & ~n41377;
  assign n41933 = ~n58702 & ~n41377;
  assign n41934 = ~n41932 & ~n41933;
  assign n41935 = ~n41377 & ~n41931;
  assign n41936 = ~n41930 & ~n58785;
  assign n41937 = n18846 & n40476;
  assign n41938 = n19541 & n39594;
  assign n41939 = n55247 & n39600;
  assign n41940 = n19509 & n39597;
  assign n41941 = ~n41939 & ~n41940;
  assign n41942 = ~n41938 & n41941;
  assign n41943 = ~n41937 & n41942;
  assign n41944 = pi11  & ~n41943;
  assign n41945 = ~n41943 & ~n41944;
  assign n41946 = ~pi11  & ~n41943;
  assign n41947 = pi11  & ~n41944;
  assign n41948 = pi11  & n41943;
  assign n41949 = ~n58786 & ~n58787;
  assign n41950 = n41360 & n58699;
  assign n41951 = ~n41360 & ~n41368;
  assign n41952 = ~n41360 & n58699;
  assign n41953 = ~n58699 & ~n41368;
  assign n41954 = n41360 & ~n58699;
  assign n41955 = ~n58788 & ~n58789;
  assign n41956 = ~n41368 & ~n41950;
  assign n41957 = ~n41949 & ~n58790;
  assign n41958 = n41351 & n58696;
  assign n41959 = ~n41359 & ~n41958;
  assign n41960 = n18846 & n40247;
  assign n41961 = n19541 & n39597;
  assign n41962 = n55247 & n39603;
  assign n41963 = n19509 & n39600;
  assign n41964 = ~n41962 & ~n41963;
  assign n41965 = ~n41961 & n41964;
  assign n41966 = ~n18846 & n41965;
  assign n41967 = ~n40247 & n41965;
  assign n41968 = ~n41966 & ~n41967;
  assign n41969 = ~n41960 & n41965;
  assign n41970 = pi11  & ~n58791;
  assign n41971 = ~pi11  & n58791;
  assign n41972 = ~n41970 & ~n41971;
  assign n41973 = n41959 & ~n41972;
  assign n41974 = n41347 & ~n41349;
  assign n41975 = ~n41350 & ~n41974;
  assign n41976 = n18846 & ~n58533;
  assign n41977 = n19541 & n39600;
  assign n41978 = n55247 & n39606;
  assign n41979 = n19509 & n39603;
  assign n41980 = ~n41978 & ~n41979;
  assign n41981 = ~n41977 & n41980;
  assign n41982 = ~n18846 & n41981;
  assign n41983 = n58533 & n41981;
  assign n41984 = ~n41982 & ~n41983;
  assign n41985 = ~n41976 & n41981;
  assign n41986 = pi11  & ~n58792;
  assign n41987 = ~pi11  & n58792;
  assign n41988 = ~n41986 & ~n41987;
  assign n41989 = n41975 & ~n41988;
  assign n41990 = n41338 & n58693;
  assign n41991 = ~n41346 & ~n41990;
  assign n41992 = n18846 & n40286;
  assign n41993 = n19541 & n39603;
  assign n41994 = n55247 & n39609;
  assign n41995 = n19509 & n39606;
  assign n41996 = ~n41994 & ~n41995;
  assign n41997 = ~n41993 & n41996;
  assign n41998 = ~n18846 & n41997;
  assign n41999 = ~n40286 & n41997;
  assign n42000 = ~n41998 & ~n41999;
  assign n42001 = ~n41992 & n41997;
  assign n42002 = pi11  & ~n58793;
  assign n42003 = ~pi11  & n58793;
  assign n42004 = ~n42002 & ~n42003;
  assign n42005 = n41991 & ~n42004;
  assign n42006 = n18846 & n40183;
  assign n42007 = n19541 & n39606;
  assign n42008 = n55247 & n39612;
  assign n42009 = n19509 & n39609;
  assign n42010 = ~n42008 & ~n42009;
  assign n42011 = ~n42007 & n42010;
  assign n42012 = ~n42006 & n42011;
  assign n42013 = pi11  & ~n42012;
  assign n42014 = ~n42012 & ~n42013;
  assign n42015 = ~pi11  & ~n42012;
  assign n42016 = pi11  & ~n42013;
  assign n42017 = pi11  & n42012;
  assign n42018 = ~n58794 & ~n58795;
  assign n42019 = n41334 & ~n41336;
  assign n42020 = ~n41337 & ~n42019;
  assign n42021 = ~n42018 & n42020;
  assign n42022 = n18846 & n39991;
  assign n42023 = n19541 & n39609;
  assign n42024 = n55247 & n39615;
  assign n42025 = n19509 & n39612;
  assign n42026 = ~n42024 & ~n42025;
  assign n42027 = ~n42023 & n42026;
  assign n42028 = ~n18846 & n42027;
  assign n42029 = ~n39991 & n42027;
  assign n42030 = ~n42028 & ~n42029;
  assign n42031 = ~n42022 & n42027;
  assign n42032 = pi11  & ~n58796;
  assign n42033 = ~pi11  & n58796;
  assign n42034 = ~n42032 & ~n42033;
  assign n42035 = n41325 & n58690;
  assign n42036 = ~n58690 & ~n41333;
  assign n42037 = ~n41325 & ~n41333;
  assign n42038 = ~n42036 & ~n42037;
  assign n42039 = ~n41333 & ~n42035;
  assign n42040 = ~n42034 & ~n58797;
  assign n42041 = n18846 & n40071;
  assign n42042 = n19541 & n39612;
  assign n42043 = n55247 & n39618;
  assign n42044 = n19509 & n39615;
  assign n42045 = ~n42043 & ~n42044;
  assign n42046 = ~n42042 & n42045;
  assign n42047 = ~n42041 & n42046;
  assign n42048 = pi11  & ~n42047;
  assign n42049 = ~n42047 & ~n42048;
  assign n42050 = ~pi11  & ~n42047;
  assign n42051 = pi11  & ~n42048;
  assign n42052 = pi11  & n42047;
  assign n42053 = ~n58798 & ~n58799;
  assign n42054 = pi14  & ~n58683;
  assign n42055 = ~n58684 & ~n42054;
  assign n42056 = n58684 & n42054;
  assign n42057 = ~n58683 & n41309;
  assign n42058 = ~n58685 & ~n42057;
  assign n42059 = ~n42055 & ~n42056;
  assign n42060 = ~n42053 & n58800;
  assign n42061 = n18846 & n40093;
  assign n42062 = n19541 & n39615;
  assign n42063 = n55247 & n39621;
  assign n42064 = n19509 & n39618;
  assign n42065 = ~n42063 & ~n42064;
  assign n42066 = ~n42062 & n42065;
  assign n42067 = ~n18846 & n42066;
  assign n42068 = ~n40093 & n42066;
  assign n42069 = ~n42067 & ~n42068;
  assign n42070 = ~n42061 & n42066;
  assign n42071 = pi11  & ~n58801;
  assign n42072 = ~pi11  & n58801;
  assign n42073 = ~n42071 & ~n42072;
  assign n42074 = pi14  & n41289;
  assign n42075 = ~n41288 & n42074;
  assign n42076 = n41288 & ~n42074;
  assign n42077 = ~n41290 & n41294;
  assign n42078 = ~n58683 & ~n42077;
  assign n42079 = ~n42075 & ~n42076;
  assign n42080 = ~n42073 & n58802;
  assign n42081 = n18846 & ~n40023;
  assign n42082 = n19509 & ~n58457;
  assign n42083 = n19541 & n39626;
  assign n42084 = ~n42082 & ~n42083;
  assign n42085 = ~n42081 & n42084;
  assign n42086 = n55244 & ~n58457;
  assign n42087 = pi11  & ~n42086;
  assign n42088 = pi11  & ~n42085;
  assign n42089 = pi11  & ~n42088;
  assign n42090 = ~n42085 & ~n42088;
  assign n42091 = ~n42089 & ~n42090;
  assign n42092 = n42087 & ~n42091;
  assign n42093 = n42085 & n42087;
  assign n42094 = n18846 & ~n40039;
  assign n42095 = n19541 & n39621;
  assign n42096 = n55247 & ~n58457;
  assign n42097 = n19509 & n39626;
  assign n42098 = ~n42096 & ~n42097;
  assign n42099 = ~n42095 & n42098;
  assign n42100 = ~n18846 & n42099;
  assign n42101 = n40039 & n42099;
  assign n42102 = ~n42100 & ~n42101;
  assign n42103 = ~n42094 & n42099;
  assign n42104 = pi11  & ~n58804;
  assign n42105 = ~pi11  & n58804;
  assign n42106 = ~n42104 & ~n42105;
  assign n42107 = n58803 & ~n42106;
  assign n42108 = n58803 & ~n58804;
  assign n42109 = n41289 & n58805;
  assign n42110 = n18846 & n40006;
  assign n42111 = n19541 & n39618;
  assign n42112 = n55247 & n39626;
  assign n42113 = n19509 & n39621;
  assign n42114 = ~n42112 & ~n42113;
  assign n42115 = ~n42111 & n42114;
  assign n42116 = ~n42110 & n42115;
  assign n42117 = pi11  & ~n42116;
  assign n42118 = pi11  & ~n42117;
  assign n42119 = pi11  & n42116;
  assign n42120 = ~n42116 & ~n42117;
  assign n42121 = ~pi11  & ~n42116;
  assign n42122 = ~n58806 & ~n58807;
  assign n42123 = ~n41289 & ~n58805;
  assign n42124 = n58805 & ~n42109;
  assign n42125 = ~n41289 & n58805;
  assign n42126 = n41289 & ~n42109;
  assign n42127 = n41289 & ~n58805;
  assign n42128 = ~n58808 & ~n58809;
  assign n42129 = ~n42109 & ~n42123;
  assign n42130 = ~n42122 & ~n58810;
  assign n42131 = ~n42109 & ~n42130;
  assign n42132 = n42073 & ~n58802;
  assign n42133 = ~n42080 & ~n42132;
  assign n42134 = ~n42131 & n42133;
  assign n42135 = ~n42080 & ~n42134;
  assign n42136 = n42053 & ~n58800;
  assign n42137 = ~n42053 & ~n42060;
  assign n42138 = ~n42053 & ~n58800;
  assign n42139 = n58800 & ~n42060;
  assign n42140 = n42053 & n58800;
  assign n42141 = ~n58811 & ~n58812;
  assign n42142 = ~n42060 & ~n42136;
  assign n42143 = ~n42135 & ~n58813;
  assign n42144 = ~n42060 & ~n42143;
  assign n42145 = n42034 & n58797;
  assign n42146 = ~n42040 & ~n42145;
  assign n42147 = ~n42144 & n42146;
  assign n42148 = ~n42040 & ~n42147;
  assign n42149 = n42018 & ~n42020;
  assign n42150 = ~n42018 & ~n42021;
  assign n42151 = ~n42018 & ~n42020;
  assign n42152 = n42020 & ~n42021;
  assign n42153 = n42018 & n42020;
  assign n42154 = ~n58814 & ~n58815;
  assign n42155 = ~n42021 & ~n42149;
  assign n42156 = ~n42148 & ~n58816;
  assign n42157 = ~n42021 & ~n42156;
  assign n42158 = ~n41991 & n42004;
  assign n42159 = n41991 & ~n42005;
  assign n42160 = n41991 & n42004;
  assign n42161 = ~n42004 & ~n42005;
  assign n42162 = ~n41991 & ~n42004;
  assign n42163 = ~n58817 & ~n58818;
  assign n42164 = ~n42005 & ~n42158;
  assign n42165 = ~n42157 & ~n58819;
  assign n42166 = ~n42005 & ~n42165;
  assign n42167 = ~n41975 & n41988;
  assign n42168 = n41975 & ~n41989;
  assign n42169 = n41975 & n41988;
  assign n42170 = ~n41988 & ~n41989;
  assign n42171 = ~n41975 & ~n41988;
  assign n42172 = ~n58820 & ~n58821;
  assign n42173 = ~n41989 & ~n42167;
  assign n42174 = ~n42166 & ~n58822;
  assign n42175 = ~n41989 & ~n42174;
  assign n42176 = ~n41959 & n41972;
  assign n42177 = ~n41973 & ~n42176;
  assign n42178 = ~n42175 & n42177;
  assign n42179 = ~n41973 & ~n42178;
  assign n42180 = n41949 & n58790;
  assign n42181 = ~n41949 & ~n41957;
  assign n42182 = ~n58790 & ~n41957;
  assign n42183 = ~n42181 & ~n42182;
  assign n42184 = ~n41957 & ~n42180;
  assign n42185 = ~n42179 & ~n58823;
  assign n42186 = ~n41957 & ~n42185;
  assign n42187 = n41930 & n58785;
  assign n42188 = ~n41930 & ~n41936;
  assign n42189 = ~n41930 & n58785;
  assign n42190 = ~n58785 & ~n41936;
  assign n42191 = n41930 & ~n58785;
  assign n42192 = ~n58824 & ~n58825;
  assign n42193 = ~n41936 & ~n42187;
  assign n42194 = ~n42186 & ~n58826;
  assign n42195 = ~n41936 & ~n42194;
  assign n42196 = n41914 & ~n41916;
  assign n42197 = ~n41914 & ~n41917;
  assign n42198 = ~n41914 & ~n41916;
  assign n42199 = n41916 & ~n41917;
  assign n42200 = n41914 & n41916;
  assign n42201 = ~n58827 & ~n58828;
  assign n42202 = ~n41917 & ~n42196;
  assign n42203 = ~n42195 & ~n58829;
  assign n42204 = ~n41917 & ~n42203;
  assign n42205 = ~n41887 & n41900;
  assign n42206 = n41887 & ~n41901;
  assign n42207 = n41887 & n41900;
  assign n42208 = ~n41900 & ~n41901;
  assign n42209 = ~n41887 & ~n41900;
  assign n42210 = ~n58830 & ~n58831;
  assign n42211 = ~n41901 & ~n42205;
  assign n42212 = ~n42204 & ~n58832;
  assign n42213 = ~n41901 & ~n42212;
  assign n42214 = ~n41871 & n41884;
  assign n42215 = n41871 & ~n41885;
  assign n42216 = n41871 & n41884;
  assign n42217 = ~n41884 & ~n41885;
  assign n42218 = ~n41871 & ~n41884;
  assign n42219 = ~n58833 & ~n58834;
  assign n42220 = ~n41885 & ~n42214;
  assign n42221 = ~n42213 & ~n58835;
  assign n42222 = ~n41885 & ~n42221;
  assign n42223 = ~n41855 & n41868;
  assign n42224 = ~n41869 & ~n42223;
  assign n42225 = ~n42222 & n42224;
  assign n42226 = ~n41869 & ~n42225;
  assign n42227 = n41847 & n58777;
  assign n42228 = ~n41847 & ~n41853;
  assign n42229 = ~n41847 & n58777;
  assign n42230 = ~n58777 & ~n41853;
  assign n42231 = n41847 & ~n58777;
  assign n42232 = ~n58836 & ~n58837;
  assign n42233 = ~n41853 & ~n42227;
  assign n42234 = ~n42226 & ~n58838;
  assign n42235 = ~n41853 & ~n42234;
  assign n42236 = n41826 & n58774;
  assign n42237 = ~n41826 & ~n41834;
  assign n42238 = ~n58774 & ~n41834;
  assign n42239 = ~n42237 & ~n42238;
  assign n42240 = ~n41834 & ~n42236;
  assign n42241 = ~n42235 & ~n58839;
  assign n42242 = ~n41834 & ~n42241;
  assign n42243 = n41810 & ~n41812;
  assign n42244 = ~n41810 & ~n41813;
  assign n42245 = ~n41810 & ~n41812;
  assign n42246 = n41812 & ~n41813;
  assign n42247 = n41810 & n41812;
  assign n42248 = ~n58840 & ~n58841;
  assign n42249 = ~n41813 & ~n42243;
  assign n42250 = ~n42242 & ~n58842;
  assign n42251 = ~n41813 & ~n42250;
  assign n42252 = ~n41778 & n41796;
  assign n42253 = n41778 & ~n41797;
  assign n42254 = n41778 & n41796;
  assign n42255 = ~n41796 & ~n41797;
  assign n42256 = ~n41778 & ~n41796;
  assign n42257 = ~n58843 & ~n58844;
  assign n42258 = ~n41797 & ~n42252;
  assign n42259 = ~n42251 & ~n58845;
  assign n42260 = ~n41797 & ~n42259;
  assign n42261 = ~n41760 & n41775;
  assign n42262 = ~n41776 & ~n42261;
  assign n42263 = ~n42260 & n42262;
  assign n42264 = ~n41776 & ~n42263;
  assign n42265 = n39974 & n58764;
  assign n42266 = ~n39974 & ~n41758;
  assign n42267 = ~n39974 & n58764;
  assign n42268 = ~n58764 & ~n41758;
  assign n42269 = n39974 & ~n58764;
  assign n42270 = ~n58846 & ~n58847;
  assign n42271 = ~n41758 & ~n42265;
  assign n42272 = ~n42264 & ~n58848;
  assign n42273 = ~n41758 & ~n42272;
  assign n42274 = n39731 & ~n39733;
  assign n42275 = ~n39731 & ~n58467;
  assign n42276 = ~n39732 & n39737;
  assign n42277 = ~n42275 & ~n42276;
  assign n42278 = ~n58467 & ~n42274;
  assign n42279 = n18846 & ~n58849;
  assign n42280 = n19541 & n39558;
  assign n42281 = n55247 & n39564;
  assign n42282 = n19509 & n39561;
  assign n42283 = ~n42281 & ~n42282;
  assign n42284 = ~n42280 & n42283;
  assign n42285 = ~n42279 & n42284;
  assign n42286 = pi11  & ~n42285;
  assign n42287 = ~n42285 & ~n42286;
  assign n42288 = ~pi11  & ~n42285;
  assign n42289 = pi11  & ~n42286;
  assign n42290 = pi11  & n42285;
  assign n42291 = ~n58850 & ~n58851;
  assign n42292 = ~n41744 & ~n41752;
  assign n42293 = ~n41717 & ~n41723;
  assign n42294 = n16079 & ~n58653;
  assign n42295 = n16696 & n39576;
  assign n42296 = n54886 & n39582;
  assign n42297 = n16676 & n39579;
  assign n42298 = ~n42296 & ~n42297;
  assign n42299 = ~n42295 & n42298;
  assign n42300 = ~n42294 & n42299;
  assign n42301 = pi17  & ~n42300;
  assign n42302 = ~n42300 & ~n42301;
  assign n42303 = ~pi17  & ~n42300;
  assign n42304 = pi17  & ~n42301;
  assign n42305 = pi17  & n42300;
  assign n42306 = ~n58852 & ~n58853;
  assign n42307 = ~n41701 & ~n41709;
  assign n42308 = ~n41677 & ~n41686;
  assign n42309 = n90 & n40476;
  assign n42310 = n14236 & n39594;
  assign n42311 = n54667 & n39600;
  assign n42312 = n14210 & n39597;
  assign n42313 = ~n42311 & ~n42312;
  assign n42314 = ~n42310 & n42313;
  assign n42315 = ~n42309 & n42314;
  assign n42316 = pi23  & ~n42315;
  assign n42317 = ~n42315 & ~n42316;
  assign n42318 = ~pi23  & ~n42315;
  assign n42319 = pi23  & ~n42316;
  assign n42320 = pi23  & n42315;
  assign n42321 = ~n58854 & ~n58855;
  assign n42322 = ~n41663 & ~n41671;
  assign n42323 = ~n41651 & ~n41657;
  assign n42324 = n11279 & n40071;
  assign n42325 = n12584 & n39612;
  assign n42326 = n54410 & n39618;
  assign n42327 = n11267 & n39615;
  assign n42328 = ~n42326 & ~n42327;
  assign n42329 = ~n42325 & n42328;
  assign n42330 = ~n42324 & n42329;
  assign n42331 = pi29  & ~n42330;
  assign n42332 = ~n42330 & ~n42331;
  assign n42333 = ~pi29  & ~n42330;
  assign n42334 = pi29  & ~n42331;
  assign n42335 = pi29  & n42330;
  assign n42336 = ~n58856 & ~n58857;
  assign n42337 = ~n443 & ~n493;
  assign n42338 = ~n316 & ~n1478;
  assign n42339 = n42337 & n42338;
  assign n42340 = n8970 & n13807;
  assign n42341 = n27077 & n58858;
  assign n42342 = n53923 & n42341;
  assign n42343 = n54452 & n54539;
  assign n42344 = n42342 & n42343;
  assign n42345 = n1266 & n4376;
  assign n42346 = n5021 & n5874;
  assign n42347 = n42345 & n42346;
  assign n42348 = ~n144 & ~n349;
  assign n42349 = ~n144 & ~n788;
  assign n42350 = ~n349 & n42349;
  assign n42351 = ~n349 & ~n788;
  assign n42352 = ~n144 & n42351;
  assign n42353 = ~n788 & n42348;
  assign n42354 = ~n560 & ~n851;
  assign n42355 = n652 & n42354;
  assign n42356 = n58859 & n42355;
  assign n42357 = n652 & n1266;
  assign n42358 = n4376 & n5021;
  assign n42359 = n42357 & n42358;
  assign n42360 = n5874 & n42354;
  assign n42361 = n58859 & n42360;
  assign n42362 = n42359 & n42361;
  assign n42363 = n42347 & n42356;
  assign n42364 = n54814 & n58860;
  assign n42365 = n27077 & n42357;
  assign n42366 = n53923 & n42365;
  assign n42367 = n42343 & n42366;
  assign n42368 = n42358 & n42360;
  assign n42369 = n58858 & n58859;
  assign n42370 = n42368 & n42369;
  assign n42371 = n54814 & n42370;
  assign n42372 = n42367 & n42371;
  assign n42373 = n42344 & n42364;
  assign n42374 = n55118 & n58861;
  assign n42375 = n27077 & n58859;
  assign n42376 = n1266 & n42375;
  assign n42377 = n54452 & n42376;
  assign n42378 = n652 & n42377;
  assign n42379 = n54539 & n42378;
  assign n42380 = n55118 & n42379;
  assign n42381 = n54814 & n42380;
  assign n42382 = n53923 & n42381;
  assign n42383 = n4376 & n42382;
  assign n42384 = n5874 & n42383;
  assign n42385 = n5021 & n42384;
  assign n42386 = n57028 & n42385;
  assign n42387 = ~n316 & n42386;
  assign n42388 = ~n1478 & n42387;
  assign n42389 = ~n560 & n42388;
  assign n42390 = ~n493 & n42389;
  assign n42391 = ~n851 & n42390;
  assign n42392 = ~n443 & n42391;
  assign n42393 = n57028 & n42374;
  assign n42394 = n41643 & ~n58862;
  assign n42395 = ~n41643 & n58862;
  assign n42396 = ~n42394 & ~n42395;
  assign n42397 = n1576 & ~n40039;
  assign n42398 = n11215 & n39621;
  assign n42399 = n54403 & ~n58457;
  assign n42400 = n10564 & n39626;
  assign n42401 = ~n42399 & ~n42400;
  assign n42402 = ~n42398 & n42401;
  assign n42403 = ~n42397 & n42402;
  assign n42404 = ~n42396 & n42403;
  assign n42405 = n42396 & ~n42403;
  assign n42406 = ~n42403 & ~n42405;
  assign n42407 = n42396 & ~n42405;
  assign n42408 = ~n42406 & ~n42407;
  assign n42409 = ~n42404 & ~n42405;
  assign n42410 = ~n42336 & ~n58863;
  assign n42411 = n42336 & n58863;
  assign n42412 = ~n42336 & ~n42410;
  assign n42413 = ~n58863 & ~n42410;
  assign n42414 = ~n42412 & ~n42413;
  assign n42415 = ~n42410 & ~n42411;
  assign n42416 = n42323 & n58864;
  assign n42417 = ~n42323 & ~n58864;
  assign n42418 = ~n42416 & ~n42417;
  assign n42419 = n123 & n40286;
  assign n42420 = n128 & n39603;
  assign n42421 = n53444 & n39609;
  assign n42422 = n127 & n39606;
  assign n42423 = ~n42421 & ~n42422;
  assign n42424 = ~n42420 & n42423;
  assign n42425 = ~n123 & n42424;
  assign n42426 = ~n40286 & n42424;
  assign n42427 = ~n42425 & ~n42426;
  assign n42428 = ~n42419 & n42424;
  assign n42429 = pi26  & ~n58865;
  assign n42430 = ~pi26  & n58865;
  assign n42431 = ~n42429 & ~n42430;
  assign n42432 = n42418 & ~n42431;
  assign n42433 = ~n42418 & n42431;
  assign n42434 = n42418 & ~n42432;
  assign n42435 = n42418 & n42431;
  assign n42436 = ~n42431 & ~n42432;
  assign n42437 = ~n42418 & ~n42431;
  assign n42438 = ~n58866 & ~n58867;
  assign n42439 = ~n42432 & ~n42433;
  assign n42440 = ~n42322 & ~n58868;
  assign n42441 = n42322 & n58868;
  assign n42442 = ~n42322 & ~n42440;
  assign n42443 = ~n58868 & ~n42440;
  assign n42444 = ~n42442 & ~n42443;
  assign n42445 = ~n42440 & ~n42441;
  assign n42446 = ~n42321 & ~n58869;
  assign n42447 = n42321 & n58869;
  assign n42448 = ~n42321 & ~n42446;
  assign n42449 = ~n42321 & n58869;
  assign n42450 = ~n58869 & ~n42446;
  assign n42451 = n42321 & ~n58869;
  assign n42452 = ~n58870 & ~n58871;
  assign n42453 = ~n42446 & ~n42447;
  assign n42454 = n42308 & n58872;
  assign n42455 = ~n42308 & ~n58872;
  assign n42456 = ~n42454 & ~n42455;
  assign n42457 = n14413 & ~n58583;
  assign n42458 = n15921 & n39585;
  assign n42459 = n54719 & n39591;
  assign n42460 = n15901 & n39588;
  assign n42461 = ~n42459 & ~n42460;
  assign n42462 = ~n42458 & n42461;
  assign n42463 = ~n14413 & n42462;
  assign n42464 = n58583 & n42462;
  assign n42465 = ~n42463 & ~n42464;
  assign n42466 = ~n42457 & n42462;
  assign n42467 = pi20  & ~n58873;
  assign n42468 = ~pi20  & n58873;
  assign n42469 = ~n42467 & ~n42468;
  assign n42470 = n42456 & ~n42469;
  assign n42471 = ~n42456 & n42469;
  assign n42472 = n42456 & ~n42470;
  assign n42473 = n42456 & n42469;
  assign n42474 = ~n42469 & ~n42470;
  assign n42475 = ~n42456 & ~n42469;
  assign n42476 = ~n58874 & ~n58875;
  assign n42477 = ~n42470 & ~n42471;
  assign n42478 = ~n42307 & ~n58876;
  assign n42479 = n42307 & n58876;
  assign n42480 = ~n42307 & ~n42478;
  assign n42481 = ~n42307 & n58876;
  assign n42482 = ~n58876 & ~n42478;
  assign n42483 = n42307 & ~n58876;
  assign n42484 = ~n58877 & ~n58878;
  assign n42485 = ~n42478 & ~n42479;
  assign n42486 = ~n42306 & ~n58879;
  assign n42487 = n42306 & n58879;
  assign n42488 = ~n42306 & ~n42486;
  assign n42489 = ~n58879 & ~n42486;
  assign n42490 = ~n42488 & ~n42489;
  assign n42491 = ~n42486 & ~n42487;
  assign n42492 = n42293 & n58880;
  assign n42493 = ~n42293 & ~n58880;
  assign n42494 = ~n42492 & ~n42493;
  assign n42495 = n17265 & ~n58766;
  assign n42496 = n18588 & n39567;
  assign n42497 = n55041 & n39573;
  assign n42498 = n18556 & n39570;
  assign n42499 = ~n42497 & ~n42498;
  assign n42500 = ~n42496 & n42499;
  assign n42501 = ~n17265 & n42500;
  assign n42502 = n58766 & n42500;
  assign n42503 = ~n42501 & ~n42502;
  assign n42504 = ~n42495 & n42500;
  assign n42505 = pi14  & ~n58881;
  assign n42506 = ~pi14  & n58881;
  assign n42507 = ~n42505 & ~n42506;
  assign n42508 = n42494 & ~n42507;
  assign n42509 = ~n42494 & n42507;
  assign n42510 = n42494 & ~n42508;
  assign n42511 = n42494 & n42507;
  assign n42512 = ~n42507 & ~n42508;
  assign n42513 = ~n42494 & ~n42507;
  assign n42514 = ~n58882 & ~n58883;
  assign n42515 = ~n42508 & ~n42509;
  assign n42516 = ~n42292 & ~n58884;
  assign n42517 = n42292 & n58884;
  assign n42518 = ~n42292 & ~n42516;
  assign n42519 = ~n58884 & ~n42516;
  assign n42520 = ~n42518 & ~n42519;
  assign n42521 = ~n42516 & ~n42517;
  assign n42522 = ~n42291 & ~n58885;
  assign n42523 = n42291 & n58885;
  assign n42524 = ~n42291 & ~n42522;
  assign n42525 = ~n42291 & n58885;
  assign n42526 = ~n58885 & ~n42522;
  assign n42527 = n42291 & ~n58885;
  assign n42528 = ~n58886 & ~n58887;
  assign n42529 = ~n42522 & ~n42523;
  assign n42530 = ~n42273 & ~n58888;
  assign n42531 = n42273 & n58888;
  assign n42532 = ~n42530 & ~n42531;
  assign n42533 = n39747 & ~n39749;
  assign n42534 = ~n39747 & ~n58469;
  assign n42535 = ~n39748 & n39753;
  assign n42536 = ~n42534 & ~n42535;
  assign n42537 = ~n58469 & ~n42533;
  assign n42538 = n20085 & ~n58889;
  assign n42539 = n21269 & n39549;
  assign n42540 = n55472 & n39555;
  assign n42541 = n21237 & n39552;
  assign n42542 = ~n42540 & ~n42541;
  assign n42543 = ~n42539 & n42542;
  assign n42544 = ~n20085 & n42543;
  assign n42545 = n58889 & n42543;
  assign n42546 = ~n42544 & ~n42545;
  assign n42547 = ~n42538 & n42543;
  assign n42548 = pi8  & ~n58890;
  assign n42549 = ~pi8  & n58890;
  assign n42550 = ~n42548 & ~n42549;
  assign n42551 = n42532 & ~n42550;
  assign n42552 = n42264 & n58848;
  assign n42553 = ~n42272 & ~n42552;
  assign n42554 = n39741 & ~n39743;
  assign n42555 = ~n39741 & ~n58468;
  assign n42556 = ~n39742 & n39747;
  assign n42557 = ~n42555 & ~n42556;
  assign n42558 = ~n58468 & ~n42554;
  assign n42559 = n20085 & ~n58891;
  assign n42560 = n21269 & n39552;
  assign n42561 = n55472 & n39558;
  assign n42562 = n21237 & n39555;
  assign n42563 = ~n42561 & ~n42562;
  assign n42564 = ~n42560 & n42563;
  assign n42565 = ~n20085 & n42564;
  assign n42566 = n58891 & n42564;
  assign n42567 = ~n42565 & ~n42566;
  assign n42568 = ~n42559 & n42564;
  assign n42569 = pi8  & ~n58892;
  assign n42570 = ~pi8  & n58892;
  assign n42571 = ~n42569 & ~n42570;
  assign n42572 = n42553 & ~n42571;
  assign n42573 = n39737 & ~n39739;
  assign n42574 = ~n39740 & ~n42573;
  assign n42575 = n20085 & n42574;
  assign n42576 = n21269 & n39555;
  assign n42577 = n55472 & n39561;
  assign n42578 = n21237 & n39558;
  assign n42579 = ~n42577 & ~n42578;
  assign n42580 = ~n42576 & n42579;
  assign n42581 = ~n42575 & n42580;
  assign n42582 = pi8  & ~n42581;
  assign n42583 = ~n42581 & ~n42582;
  assign n42584 = ~pi8  & ~n42581;
  assign n42585 = pi8  & ~n42582;
  assign n42586 = pi8  & n42581;
  assign n42587 = ~n58893 & ~n58894;
  assign n42588 = n42260 & ~n42262;
  assign n42589 = ~n42263 & ~n42588;
  assign n42590 = ~n42587 & n42589;
  assign n42591 = n20085 & ~n58849;
  assign n42592 = n21269 & n39558;
  assign n42593 = n55472 & n39564;
  assign n42594 = n21237 & n39561;
  assign n42595 = ~n42593 & ~n42594;
  assign n42596 = ~n42592 & n42595;
  assign n42597 = ~n42591 & n42596;
  assign n42598 = pi8  & ~n42597;
  assign n42599 = ~n42597 & ~n42598;
  assign n42600 = ~pi8  & ~n42597;
  assign n42601 = pi8  & ~n42598;
  assign n42602 = pi8  & n42597;
  assign n42603 = ~n58895 & ~n58896;
  assign n42604 = n42251 & n58845;
  assign n42605 = ~n42251 & ~n42259;
  assign n42606 = ~n42251 & n58845;
  assign n42607 = ~n58845 & ~n42259;
  assign n42608 = n42251 & ~n58845;
  assign n42609 = ~n58897 & ~n58898;
  assign n42610 = ~n42259 & ~n42604;
  assign n42611 = ~n42603 & ~n58899;
  assign n42612 = n42242 & n58842;
  assign n42613 = ~n42250 & ~n42612;
  assign n42614 = n20085 & ~n58493;
  assign n42615 = n21269 & n39561;
  assign n42616 = n55472 & n39567;
  assign n42617 = n21237 & n39564;
  assign n42618 = ~n42616 & ~n42617;
  assign n42619 = ~n42615 & n42618;
  assign n42620 = ~n20085 & n42619;
  assign n42621 = n58493 & n42619;
  assign n42622 = ~n42620 & ~n42621;
  assign n42623 = ~n42614 & n42619;
  assign n42624 = pi8  & ~n58900;
  assign n42625 = ~pi8  & n58900;
  assign n42626 = ~n42624 & ~n42625;
  assign n42627 = n42613 & ~n42626;
  assign n42628 = n42235 & n58839;
  assign n42629 = ~n42241 & ~n42628;
  assign n42630 = n20085 & n41762;
  assign n42631 = n21269 & n39564;
  assign n42632 = n55472 & n39570;
  assign n42633 = n21237 & n39567;
  assign n42634 = ~n42632 & ~n42633;
  assign n42635 = ~n42631 & n42634;
  assign n42636 = ~n20085 & n42635;
  assign n42637 = ~n41762 & n42635;
  assign n42638 = ~n42636 & ~n42637;
  assign n42639 = ~n42630 & n42635;
  assign n42640 = pi8  & ~n58901;
  assign n42641 = ~pi8  & n58901;
  assign n42642 = ~n42640 & ~n42641;
  assign n42643 = n42629 & ~n42642;
  assign n42644 = n42226 & n58838;
  assign n42645 = ~n42234 & ~n42644;
  assign n42646 = n20085 & ~n58766;
  assign n42647 = n21269 & n39567;
  assign n42648 = n55472 & n39573;
  assign n42649 = n21237 & n39570;
  assign n42650 = ~n42648 & ~n42649;
  assign n42651 = ~n42647 & n42650;
  assign n42652 = ~n20085 & n42651;
  assign n42653 = n58766 & n42651;
  assign n42654 = ~n42652 & ~n42653;
  assign n42655 = ~n42646 & n42651;
  assign n42656 = pi8  & ~n58902;
  assign n42657 = ~pi8  & n58902;
  assign n42658 = ~n42656 & ~n42657;
  assign n42659 = n42645 & ~n42658;
  assign n42660 = n20085 & ~n58759;
  assign n42661 = n21269 & n39570;
  assign n42662 = n55472 & n39576;
  assign n42663 = n21237 & n39573;
  assign n42664 = ~n42662 & ~n42663;
  assign n42665 = ~n42661 & n42664;
  assign n42666 = ~n42660 & n42665;
  assign n42667 = pi8  & ~n42666;
  assign n42668 = ~n42666 & ~n42667;
  assign n42669 = ~pi8  & ~n42666;
  assign n42670 = pi8  & ~n42667;
  assign n42671 = pi8  & n42666;
  assign n42672 = ~n58903 & ~n58904;
  assign n42673 = n42222 & ~n42224;
  assign n42674 = ~n42225 & ~n42673;
  assign n42675 = ~n42672 & n42674;
  assign n42676 = n20085 & n39976;
  assign n42677 = n21269 & n39573;
  assign n42678 = n55472 & n39579;
  assign n42679 = n21237 & n39576;
  assign n42680 = ~n42678 & ~n42679;
  assign n42681 = ~n42677 & n42680;
  assign n42682 = ~n42676 & n42681;
  assign n42683 = pi8  & ~n42682;
  assign n42684 = ~n42682 & ~n42683;
  assign n42685 = ~pi8  & ~n42682;
  assign n42686 = pi8  & ~n42683;
  assign n42687 = pi8  & n42682;
  assign n42688 = ~n58905 & ~n58906;
  assign n42689 = n42213 & n58835;
  assign n42690 = ~n42213 & ~n42221;
  assign n42691 = ~n42213 & n58835;
  assign n42692 = ~n58835 & ~n42221;
  assign n42693 = n42213 & ~n58835;
  assign n42694 = ~n58907 & ~n58908;
  assign n42695 = ~n42221 & ~n42689;
  assign n42696 = ~n42688 & ~n58909;
  assign n42697 = n20085 & ~n58653;
  assign n42698 = n21269 & n39576;
  assign n42699 = n55472 & n39582;
  assign n42700 = n21237 & n39579;
  assign n42701 = ~n42699 & ~n42700;
  assign n42702 = ~n42698 & n42701;
  assign n42703 = ~n42697 & n42702;
  assign n42704 = pi8  & ~n42703;
  assign n42705 = ~n42703 & ~n42704;
  assign n42706 = ~pi8  & ~n42703;
  assign n42707 = pi8  & ~n42704;
  assign n42708 = pi8  & n42703;
  assign n42709 = ~n58910 & ~n58911;
  assign n42710 = n42204 & n58832;
  assign n42711 = ~n42204 & ~n42212;
  assign n42712 = ~n58832 & ~n42212;
  assign n42713 = ~n42711 & ~n42712;
  assign n42714 = ~n42212 & ~n42710;
  assign n42715 = ~n42709 & ~n58912;
  assign n42716 = n42195 & n58829;
  assign n42717 = ~n42203 & ~n42716;
  assign n42718 = n20085 & ~n58657;
  assign n42719 = n21269 & n39579;
  assign n42720 = n55472 & n39585;
  assign n42721 = n21237 & n39582;
  assign n42722 = ~n42720 & ~n42721;
  assign n42723 = ~n42719 & n42722;
  assign n42724 = ~n20085 & n42723;
  assign n42725 = n58657 & n42723;
  assign n42726 = ~n42724 & ~n42725;
  assign n42727 = ~n42718 & n42723;
  assign n42728 = pi8  & ~n58913;
  assign n42729 = ~pi8  & n58913;
  assign n42730 = ~n42728 & ~n42729;
  assign n42731 = n42717 & ~n42730;
  assign n42732 = n42186 & n58826;
  assign n42733 = ~n42194 & ~n42732;
  assign n42734 = n20085 & n41007;
  assign n42735 = n21269 & n39582;
  assign n42736 = n55472 & n39588;
  assign n42737 = n21237 & n39585;
  assign n42738 = ~n42736 & ~n42737;
  assign n42739 = ~n42735 & n42738;
  assign n42740 = ~n20085 & n42739;
  assign n42741 = ~n41007 & n42739;
  assign n42742 = ~n42740 & ~n42741;
  assign n42743 = ~n42734 & n42739;
  assign n42744 = pi8  & ~n58914;
  assign n42745 = ~pi8  & n58914;
  assign n42746 = ~n42744 & ~n42745;
  assign n42747 = n42733 & ~n42746;
  assign n42748 = n42179 & n58823;
  assign n42749 = ~n42185 & ~n42748;
  assign n42750 = n20085 & ~n58583;
  assign n42751 = n21269 & n39585;
  assign n42752 = n55472 & n39591;
  assign n42753 = n21237 & n39588;
  assign n42754 = ~n42752 & ~n42753;
  assign n42755 = ~n42751 & n42754;
  assign n42756 = ~n20085 & n42755;
  assign n42757 = n58583 & n42755;
  assign n42758 = ~n42756 & ~n42757;
  assign n42759 = ~n42750 & n42755;
  assign n42760 = pi8  & ~n58915;
  assign n42761 = ~pi8  & n58915;
  assign n42762 = ~n42760 & ~n42761;
  assign n42763 = n42749 & ~n42762;
  assign n42764 = n20085 & ~n58585;
  assign n42765 = n21269 & n39588;
  assign n42766 = n55472 & n39594;
  assign n42767 = n21237 & n39591;
  assign n42768 = ~n42766 & ~n42767;
  assign n42769 = ~n42765 & n42768;
  assign n42770 = ~n42764 & n42769;
  assign n42771 = pi8  & ~n42770;
  assign n42772 = ~n42770 & ~n42771;
  assign n42773 = ~pi8  & ~n42770;
  assign n42774 = pi8  & ~n42771;
  assign n42775 = pi8  & n42770;
  assign n42776 = ~n58916 & ~n58917;
  assign n42777 = n42175 & ~n42177;
  assign n42778 = ~n42178 & ~n42777;
  assign n42779 = ~n42776 & n42778;
  assign n42780 = n20085 & n40616;
  assign n42781 = n21269 & n39591;
  assign n42782 = n55472 & n39597;
  assign n42783 = n21237 & n39594;
  assign n42784 = ~n42782 & ~n42783;
  assign n42785 = ~n42781 & n42784;
  assign n42786 = ~n42780 & n42785;
  assign n42787 = pi8  & ~n42786;
  assign n42788 = ~n42786 & ~n42787;
  assign n42789 = ~pi8  & ~n42786;
  assign n42790 = pi8  & ~n42787;
  assign n42791 = pi8  & n42786;
  assign n42792 = ~n58918 & ~n58919;
  assign n42793 = n42166 & n58822;
  assign n42794 = ~n42166 & ~n42174;
  assign n42795 = ~n58822 & ~n42174;
  assign n42796 = ~n42794 & ~n42795;
  assign n42797 = ~n42174 & ~n42793;
  assign n42798 = ~n42792 & ~n58920;
  assign n42799 = n20085 & n40476;
  assign n42800 = n21269 & n39594;
  assign n42801 = n55472 & n39600;
  assign n42802 = n21237 & n39597;
  assign n42803 = ~n42801 & ~n42802;
  assign n42804 = ~n42800 & n42803;
  assign n42805 = ~n42799 & n42804;
  assign n42806 = pi8  & ~n42805;
  assign n42807 = ~n42805 & ~n42806;
  assign n42808 = ~pi8  & ~n42805;
  assign n42809 = pi8  & ~n42806;
  assign n42810 = pi8  & n42805;
  assign n42811 = ~n58921 & ~n58922;
  assign n42812 = n42157 & n58819;
  assign n42813 = ~n42157 & ~n42165;
  assign n42814 = ~n42157 & n58819;
  assign n42815 = ~n58819 & ~n42165;
  assign n42816 = n42157 & ~n58819;
  assign n42817 = ~n58923 & ~n58924;
  assign n42818 = ~n42165 & ~n42812;
  assign n42819 = ~n42811 & ~n58925;
  assign n42820 = n42148 & n58816;
  assign n42821 = ~n42156 & ~n42820;
  assign n42822 = n20085 & n40247;
  assign n42823 = n21269 & n39597;
  assign n42824 = n55472 & n39603;
  assign n42825 = n21237 & n39600;
  assign n42826 = ~n42824 & ~n42825;
  assign n42827 = ~n42823 & n42826;
  assign n42828 = ~n20085 & n42827;
  assign n42829 = ~n40247 & n42827;
  assign n42830 = ~n42828 & ~n42829;
  assign n42831 = ~n42822 & n42827;
  assign n42832 = pi8  & ~n58926;
  assign n42833 = ~pi8  & n58926;
  assign n42834 = ~n42832 & ~n42833;
  assign n42835 = n42821 & ~n42834;
  assign n42836 = n42144 & ~n42146;
  assign n42837 = ~n42147 & ~n42836;
  assign n42838 = n20085 & ~n58533;
  assign n42839 = n21269 & n39600;
  assign n42840 = n55472 & n39606;
  assign n42841 = n21237 & n39603;
  assign n42842 = ~n42840 & ~n42841;
  assign n42843 = ~n42839 & n42842;
  assign n42844 = ~n20085 & n42843;
  assign n42845 = n58533 & n42843;
  assign n42846 = ~n42844 & ~n42845;
  assign n42847 = ~n42838 & n42843;
  assign n42848 = pi8  & ~n58927;
  assign n42849 = ~pi8  & n58927;
  assign n42850 = ~n42848 & ~n42849;
  assign n42851 = n42837 & ~n42850;
  assign n42852 = n42135 & n58813;
  assign n42853 = ~n42143 & ~n42852;
  assign n42854 = n20085 & n40286;
  assign n42855 = n21269 & n39603;
  assign n42856 = n55472 & n39609;
  assign n42857 = n21237 & n39606;
  assign n42858 = ~n42856 & ~n42857;
  assign n42859 = ~n42855 & n42858;
  assign n42860 = ~n20085 & n42859;
  assign n42861 = ~n40286 & n42859;
  assign n42862 = ~n42860 & ~n42861;
  assign n42863 = ~n42854 & n42859;
  assign n42864 = pi8  & ~n58928;
  assign n42865 = ~pi8  & n58928;
  assign n42866 = ~n42864 & ~n42865;
  assign n42867 = n42853 & ~n42866;
  assign n42868 = n20085 & n40183;
  assign n42869 = n21269 & n39606;
  assign n42870 = n55472 & n39612;
  assign n42871 = n21237 & n39609;
  assign n42872 = ~n42870 & ~n42871;
  assign n42873 = ~n42869 & n42872;
  assign n42874 = ~n42868 & n42873;
  assign n42875 = pi8  & ~n42874;
  assign n42876 = ~n42874 & ~n42875;
  assign n42877 = ~pi8  & ~n42874;
  assign n42878 = pi8  & ~n42875;
  assign n42879 = pi8  & n42874;
  assign n42880 = ~n58929 & ~n58930;
  assign n42881 = n42131 & ~n42133;
  assign n42882 = ~n42134 & ~n42881;
  assign n42883 = ~n42880 & n42882;
  assign n42884 = n20085 & n39991;
  assign n42885 = n21269 & n39609;
  assign n42886 = n55472 & n39615;
  assign n42887 = n21237 & n39612;
  assign n42888 = ~n42886 & ~n42887;
  assign n42889 = ~n42885 & n42888;
  assign n42890 = ~n20085 & n42889;
  assign n42891 = ~n39991 & n42889;
  assign n42892 = ~n42890 & ~n42891;
  assign n42893 = ~n42884 & n42889;
  assign n42894 = pi8  & ~n58931;
  assign n42895 = ~pi8  & n58931;
  assign n42896 = ~n42894 & ~n42895;
  assign n42897 = n42122 & n58810;
  assign n42898 = ~n58810 & ~n42130;
  assign n42899 = ~n42122 & ~n42130;
  assign n42900 = ~n42898 & ~n42899;
  assign n42901 = ~n42130 & ~n42897;
  assign n42902 = ~n42896 & ~n58932;
  assign n42903 = n20085 & n40071;
  assign n42904 = n21269 & n39612;
  assign n42905 = n55472 & n39618;
  assign n42906 = n21237 & n39615;
  assign n42907 = ~n42905 & ~n42906;
  assign n42908 = ~n42904 & n42907;
  assign n42909 = ~n42903 & n42908;
  assign n42910 = pi8  & ~n42909;
  assign n42911 = ~n42909 & ~n42910;
  assign n42912 = ~pi8  & ~n42909;
  assign n42913 = pi8  & ~n42910;
  assign n42914 = pi8  & n42909;
  assign n42915 = ~n58933 & ~n58934;
  assign n42916 = pi11  & ~n58803;
  assign n42917 = ~n58804 & ~n42916;
  assign n42918 = n58804 & n42916;
  assign n42919 = ~n58803 & n42106;
  assign n42920 = ~n58805 & ~n42919;
  assign n42921 = ~n42917 & ~n42918;
  assign n42922 = ~n42915 & n58935;
  assign n42923 = n20085 & n40093;
  assign n42924 = n21269 & n39615;
  assign n42925 = n55472 & n39621;
  assign n42926 = n21237 & n39618;
  assign n42927 = ~n42925 & ~n42926;
  assign n42928 = ~n42924 & n42927;
  assign n42929 = ~n20085 & n42928;
  assign n42930 = ~n40093 & n42928;
  assign n42931 = ~n42929 & ~n42930;
  assign n42932 = ~n42923 & n42928;
  assign n42933 = pi8  & ~n58936;
  assign n42934 = ~pi8  & n58936;
  assign n42935 = ~n42933 & ~n42934;
  assign n42936 = pi11  & n42086;
  assign n42937 = ~n42085 & n42936;
  assign n42938 = n42085 & ~n42936;
  assign n42939 = ~n42087 & n42091;
  assign n42940 = ~n58803 & ~n42939;
  assign n42941 = ~n42937 & ~n42938;
  assign n42942 = ~n42935 & n58937;
  assign n42943 = n20085 & ~n40023;
  assign n42944 = n21237 & ~n58457;
  assign n42945 = n21269 & n39626;
  assign n42946 = ~n42944 & ~n42945;
  assign n42947 = ~n42943 & n42946;
  assign n42948 = n55469 & ~n58457;
  assign n42949 = pi8  & ~n42948;
  assign n42950 = pi8  & ~n42947;
  assign n42951 = pi8  & ~n42950;
  assign n42952 = ~n42947 & ~n42950;
  assign n42953 = ~n42951 & ~n42952;
  assign n42954 = n42949 & ~n42953;
  assign n42955 = n42947 & n42949;
  assign n42956 = n20085 & ~n40039;
  assign n42957 = n21269 & n39621;
  assign n42958 = n55472 & ~n58457;
  assign n42959 = n21237 & n39626;
  assign n42960 = ~n42958 & ~n42959;
  assign n42961 = ~n42957 & n42960;
  assign n42962 = ~n20085 & n42961;
  assign n42963 = n40039 & n42961;
  assign n42964 = ~n42962 & ~n42963;
  assign n42965 = ~n42956 & n42961;
  assign n42966 = pi8  & ~n58939;
  assign n42967 = ~pi8  & n58939;
  assign n42968 = ~n42966 & ~n42967;
  assign n42969 = n58938 & ~n42968;
  assign n42970 = n58938 & ~n58939;
  assign n42971 = n42086 & n58940;
  assign n42972 = n20085 & n40006;
  assign n42973 = n21269 & n39618;
  assign n42974 = n55472 & n39626;
  assign n42975 = n21237 & n39621;
  assign n42976 = ~n42974 & ~n42975;
  assign n42977 = ~n42973 & n42976;
  assign n42978 = ~n42972 & n42977;
  assign n42979 = pi8  & ~n42978;
  assign n42980 = pi8  & ~n42979;
  assign n42981 = pi8  & n42978;
  assign n42982 = ~n42978 & ~n42979;
  assign n42983 = ~pi8  & ~n42978;
  assign n42984 = ~n58941 & ~n58942;
  assign n42985 = ~n42086 & ~n58940;
  assign n42986 = n58940 & ~n42971;
  assign n42987 = ~n42086 & n58940;
  assign n42988 = n42086 & ~n42971;
  assign n42989 = n42086 & ~n58940;
  assign n42990 = ~n58943 & ~n58944;
  assign n42991 = ~n42971 & ~n42985;
  assign n42992 = ~n42984 & ~n58945;
  assign n42993 = ~n42971 & ~n42992;
  assign n42994 = n42935 & ~n58937;
  assign n42995 = ~n42942 & ~n42994;
  assign n42996 = ~n42993 & n42995;
  assign n42997 = ~n42942 & ~n42996;
  assign n42998 = n42915 & ~n58935;
  assign n42999 = ~n42915 & ~n42922;
  assign n43000 = ~n42915 & ~n58935;
  assign n43001 = n58935 & ~n42922;
  assign n43002 = n42915 & n58935;
  assign n43003 = ~n58946 & ~n58947;
  assign n43004 = ~n42922 & ~n42998;
  assign n43005 = ~n42997 & ~n58948;
  assign n43006 = ~n42922 & ~n43005;
  assign n43007 = n42896 & n58932;
  assign n43008 = ~n42902 & ~n43007;
  assign n43009 = ~n43006 & n43008;
  assign n43010 = ~n42902 & ~n43009;
  assign n43011 = n42880 & ~n42882;
  assign n43012 = ~n42880 & ~n42883;
  assign n43013 = ~n42880 & ~n42882;
  assign n43014 = n42882 & ~n42883;
  assign n43015 = n42880 & n42882;
  assign n43016 = ~n58949 & ~n58950;
  assign n43017 = ~n42883 & ~n43011;
  assign n43018 = ~n43010 & ~n58951;
  assign n43019 = ~n42883 & ~n43018;
  assign n43020 = ~n42853 & n42866;
  assign n43021 = n42853 & ~n42867;
  assign n43022 = n42853 & n42866;
  assign n43023 = ~n42866 & ~n42867;
  assign n43024 = ~n42853 & ~n42866;
  assign n43025 = ~n58952 & ~n58953;
  assign n43026 = ~n42867 & ~n43020;
  assign n43027 = ~n43019 & ~n58954;
  assign n43028 = ~n42867 & ~n43027;
  assign n43029 = ~n42837 & n42850;
  assign n43030 = n42837 & ~n42851;
  assign n43031 = n42837 & n42850;
  assign n43032 = ~n42850 & ~n42851;
  assign n43033 = ~n42837 & ~n42850;
  assign n43034 = ~n58955 & ~n58956;
  assign n43035 = ~n42851 & ~n43029;
  assign n43036 = ~n43028 & ~n58957;
  assign n43037 = ~n42851 & ~n43036;
  assign n43038 = ~n42821 & n42834;
  assign n43039 = ~n42835 & ~n43038;
  assign n43040 = ~n43037 & n43039;
  assign n43041 = ~n42835 & ~n43040;
  assign n43042 = n42811 & n58925;
  assign n43043 = ~n42811 & ~n42819;
  assign n43044 = ~n58925 & ~n42819;
  assign n43045 = ~n43043 & ~n43044;
  assign n43046 = ~n42819 & ~n43042;
  assign n43047 = ~n43041 & ~n58958;
  assign n43048 = ~n42819 & ~n43047;
  assign n43049 = n42792 & n58920;
  assign n43050 = ~n42792 & ~n42798;
  assign n43051 = ~n42792 & n58920;
  assign n43052 = ~n58920 & ~n42798;
  assign n43053 = n42792 & ~n58920;
  assign n43054 = ~n58959 & ~n58960;
  assign n43055 = ~n42798 & ~n43049;
  assign n43056 = ~n43048 & ~n58961;
  assign n43057 = ~n42798 & ~n43056;
  assign n43058 = n42776 & ~n42778;
  assign n43059 = ~n42776 & ~n42779;
  assign n43060 = ~n42776 & ~n42778;
  assign n43061 = n42778 & ~n42779;
  assign n43062 = n42776 & n42778;
  assign n43063 = ~n58962 & ~n58963;
  assign n43064 = ~n42779 & ~n43058;
  assign n43065 = ~n43057 & ~n58964;
  assign n43066 = ~n42779 & ~n43065;
  assign n43067 = ~n42749 & n42762;
  assign n43068 = n42749 & ~n42763;
  assign n43069 = n42749 & n42762;
  assign n43070 = ~n42762 & ~n42763;
  assign n43071 = ~n42749 & ~n42762;
  assign n43072 = ~n58965 & ~n58966;
  assign n43073 = ~n42763 & ~n43067;
  assign n43074 = ~n43066 & ~n58967;
  assign n43075 = ~n42763 & ~n43074;
  assign n43076 = ~n42733 & n42746;
  assign n43077 = n42733 & ~n42747;
  assign n43078 = n42733 & n42746;
  assign n43079 = ~n42746 & ~n42747;
  assign n43080 = ~n42733 & ~n42746;
  assign n43081 = ~n58968 & ~n58969;
  assign n43082 = ~n42747 & ~n43076;
  assign n43083 = ~n43075 & ~n58970;
  assign n43084 = ~n42747 & ~n43083;
  assign n43085 = ~n42717 & n42730;
  assign n43086 = ~n42731 & ~n43085;
  assign n43087 = ~n43084 & n43086;
  assign n43088 = ~n42731 & ~n43087;
  assign n43089 = n42709 & n58912;
  assign n43090 = ~n42709 & ~n42715;
  assign n43091 = ~n42709 & n58912;
  assign n43092 = ~n58912 & ~n42715;
  assign n43093 = n42709 & ~n58912;
  assign n43094 = ~n58971 & ~n58972;
  assign n43095 = ~n42715 & ~n43089;
  assign n43096 = ~n43088 & ~n58973;
  assign n43097 = ~n42715 & ~n43096;
  assign n43098 = n42688 & n58909;
  assign n43099 = ~n42688 & ~n42696;
  assign n43100 = ~n58909 & ~n42696;
  assign n43101 = ~n43099 & ~n43100;
  assign n43102 = ~n42696 & ~n43098;
  assign n43103 = ~n43097 & ~n58974;
  assign n43104 = ~n42696 & ~n43103;
  assign n43105 = n42672 & ~n42674;
  assign n43106 = ~n42672 & ~n42675;
  assign n43107 = ~n42672 & ~n42674;
  assign n43108 = n42674 & ~n42675;
  assign n43109 = n42672 & n42674;
  assign n43110 = ~n58975 & ~n58976;
  assign n43111 = ~n42675 & ~n43105;
  assign n43112 = ~n43104 & ~n58977;
  assign n43113 = ~n42675 & ~n43112;
  assign n43114 = ~n42645 & n42658;
  assign n43115 = n42645 & ~n42659;
  assign n43116 = n42645 & n42658;
  assign n43117 = ~n42658 & ~n42659;
  assign n43118 = ~n42645 & ~n42658;
  assign n43119 = ~n58978 & ~n58979;
  assign n43120 = ~n42659 & ~n43114;
  assign n43121 = ~n43113 & ~n58980;
  assign n43122 = ~n42659 & ~n43121;
  assign n43123 = ~n42629 & n42642;
  assign n43124 = n42629 & ~n42643;
  assign n43125 = n42629 & n42642;
  assign n43126 = ~n42642 & ~n42643;
  assign n43127 = ~n42629 & ~n42642;
  assign n43128 = ~n58981 & ~n58982;
  assign n43129 = ~n42643 & ~n43123;
  assign n43130 = ~n43122 & ~n58983;
  assign n43131 = ~n42643 & ~n43130;
  assign n43132 = ~n42613 & n42626;
  assign n43133 = ~n42627 & ~n43132;
  assign n43134 = ~n43131 & n43133;
  assign n43135 = ~n42627 & ~n43134;
  assign n43136 = n42603 & n58899;
  assign n43137 = ~n42603 & ~n42611;
  assign n43138 = ~n58899 & ~n42611;
  assign n43139 = ~n43137 & ~n43138;
  assign n43140 = ~n42611 & ~n43136;
  assign n43141 = ~n43135 & ~n58984;
  assign n43142 = ~n42611 & ~n43141;
  assign n43143 = n42587 & ~n42589;
  assign n43144 = ~n42587 & ~n42590;
  assign n43145 = ~n42587 & ~n42589;
  assign n43146 = n42589 & ~n42590;
  assign n43147 = n42587 & n42589;
  assign n43148 = ~n58985 & ~n58986;
  assign n43149 = ~n42590 & ~n43143;
  assign n43150 = ~n43142 & ~n58987;
  assign n43151 = ~n42590 & ~n43150;
  assign n43152 = ~n42553 & n42571;
  assign n43153 = n42553 & ~n42572;
  assign n43154 = n42553 & n42571;
  assign n43155 = ~n42571 & ~n42572;
  assign n43156 = ~n42553 & ~n42571;
  assign n43157 = ~n58988 & ~n58989;
  assign n43158 = ~n42572 & ~n43152;
  assign n43159 = ~n43151 & ~n58990;
  assign n43160 = ~n42572 & ~n43159;
  assign n43161 = ~n42532 & n42550;
  assign n43162 = n42532 & ~n42551;
  assign n43163 = n42532 & n42550;
  assign n43164 = ~n42550 & ~n42551;
  assign n43165 = ~n42532 & ~n42550;
  assign n43166 = ~n58991 & ~n58992;
  assign n43167 = ~n42551 & ~n43161;
  assign n43168 = ~n43160 & ~n58993;
  assign n43169 = ~n42551 & ~n43168;
  assign n43170 = ~n42522 & ~n42530;
  assign n43171 = n18846 & n42574;
  assign n43172 = n19541 & n39555;
  assign n43173 = n55247 & n39561;
  assign n43174 = n19509 & n39558;
  assign n43175 = ~n43173 & ~n43174;
  assign n43176 = ~n43172 & n43175;
  assign n43177 = ~n43171 & n43176;
  assign n43178 = pi11  & ~n43177;
  assign n43179 = ~n43177 & ~n43178;
  assign n43180 = ~pi11  & ~n43177;
  assign n43181 = pi11  & ~n43178;
  assign n43182 = pi11  & n43177;
  assign n43183 = ~n58994 & ~n58995;
  assign n43184 = ~n42508 & ~n42516;
  assign n43185 = ~n42486 & ~n42493;
  assign n43186 = n16079 & n39976;
  assign n43187 = n16696 & n39573;
  assign n43188 = n54886 & n39579;
  assign n43189 = n16676 & n39576;
  assign n43190 = ~n43188 & ~n43189;
  assign n43191 = ~n43187 & n43190;
  assign n43192 = ~n43186 & n43191;
  assign n43193 = pi17  & ~n43192;
  assign n43194 = ~n43192 & ~n43193;
  assign n43195 = ~pi17  & ~n43192;
  assign n43196 = pi17  & ~n43193;
  assign n43197 = pi17  & n43192;
  assign n43198 = ~n58996 & ~n58997;
  assign n43199 = ~n42470 & ~n42478;
  assign n43200 = ~n42446 & ~n42455;
  assign n43201 = n90 & n40616;
  assign n43202 = n14236 & n39591;
  assign n43203 = n54667 & n39597;
  assign n43204 = n14210 & n39594;
  assign n43205 = ~n43203 & ~n43204;
  assign n43206 = ~n43202 & n43205;
  assign n43207 = ~n43201 & n43206;
  assign n43208 = pi23  & ~n43207;
  assign n43209 = ~n43207 & ~n43208;
  assign n43210 = ~pi23  & ~n43207;
  assign n43211 = pi23  & ~n43208;
  assign n43212 = pi23  & n43207;
  assign n43213 = ~n58998 & ~n58999;
  assign n43214 = ~n42432 & ~n42440;
  assign n43215 = ~n42410 & ~n42417;
  assign n43216 = n11279 & n39991;
  assign n43217 = n12584 & n39609;
  assign n43218 = n54410 & n39615;
  assign n43219 = n11267 & n39612;
  assign n43220 = ~n43218 & ~n43219;
  assign n43221 = ~n43217 & n43220;
  assign n43222 = ~n43216 & n43221;
  assign n43223 = pi29  & ~n43222;
  assign n43224 = ~n43222 & ~n43223;
  assign n43225 = ~pi29  & ~n43222;
  assign n43226 = pi29  & ~n43223;
  assign n43227 = pi29  & n43222;
  assign n43228 = ~n59000 & ~n59001;
  assign n43229 = ~n42395 & ~n42403;
  assign n43230 = ~n42394 & ~n42405;
  assign n43231 = ~n42394 & ~n43229;
  assign n43232 = ~n564 & ~n733;
  assign n43233 = n755 & n43232;
  assign n43234 = n1673 & n2577;
  assign n43235 = n43233 & n43234;
  assign n43236 = n358 & n1578;
  assign n43237 = ~n101 & ~n1468;
  assign n43238 = ~n1468 & n3014;
  assign n43239 = ~n101 & n43238;
  assign n43240 = n3014 & n43237;
  assign n43241 = n43236 & n59003;
  assign n43242 = n43235 & n43241;
  assign n43243 = n915 & n7904;
  assign n43244 = n14965 & n43243;
  assign n43245 = n54066 & n43244;
  assign n43246 = ~n294 & ~n733;
  assign n43247 = ~n564 & ~n1644;
  assign n43248 = n7904 & n43232;
  assign n43249 = n43246 & n43247;
  assign n43250 = n59003 & n59004;
  assign n43251 = n755 & n2577;
  assign n43252 = n43236 & n43251;
  assign n43253 = n43250 & n43252;
  assign n43254 = n915 & n1673;
  assign n43255 = n14965 & n43254;
  assign n43256 = n54066 & n43255;
  assign n43257 = n43253 & n43256;
  assign n43258 = n358 & n1673;
  assign n43259 = n43251 & n43258;
  assign n43260 = n43250 & n43259;
  assign n43261 = n915 & n1578;
  assign n43262 = n14965 & n43261;
  assign n43263 = n54066 & n43262;
  assign n43264 = n43260 & n43263;
  assign n43265 = n43242 & n43245;
  assign n43266 = n54548 & n54835;
  assign n43267 = n59005 & n43266;
  assign n43268 = n53892 & n43267;
  assign n43269 = n54133 & n14965;
  assign n43270 = n59003 & n43269;
  assign n43271 = n915 & n43270;
  assign n43272 = n54066 & n43271;
  assign n43273 = n54835 & n43272;
  assign n43274 = n53892 & n43273;
  assign n43275 = n54548 & n43274;
  assign n43276 = n1578 & n43275;
  assign n43277 = n1673 & n43276;
  assign n43278 = n358 & n43277;
  assign n43279 = n755 & n43278;
  assign n43280 = n2577 & n43279;
  assign n43281 = ~n294 & n43280;
  assign n43282 = ~n564 & n43281;
  assign n43283 = ~n1644 & n43282;
  assign n43284 = ~n733 & n43283;
  assign n43285 = n54133 & n43268;
  assign n43286 = n1576 & n40006;
  assign n43287 = n11215 & n39618;
  assign n43288 = n10564 & n39621;
  assign n43289 = n54403 & n39626;
  assign n43290 = ~n43288 & ~n43289;
  assign n43291 = ~n43287 & n43290;
  assign n43292 = ~n43286 & ~n43289;
  assign n43293 = ~n43288 & n43292;
  assign n43294 = ~n43287 & n43293;
  assign n43295 = ~n43286 & n43291;
  assign n43296 = ~n59006 & ~n59007;
  assign n43297 = n59006 & n59007;
  assign n43298 = ~n59006 & ~n43296;
  assign n43299 = ~n59006 & n59007;
  assign n43300 = ~n59007 & ~n43296;
  assign n43301 = n59006 & ~n59007;
  assign n43302 = ~n59008 & ~n59009;
  assign n43303 = ~n43296 & ~n43297;
  assign n43304 = ~n59002 & ~n59010;
  assign n43305 = n59002 & n59010;
  assign n43306 = ~n59002 & ~n43304;
  assign n43307 = ~n59010 & ~n43304;
  assign n43308 = ~n43306 & ~n43307;
  assign n43309 = ~n43304 & ~n43305;
  assign n43310 = ~n43228 & ~n59011;
  assign n43311 = n43228 & n59011;
  assign n43312 = ~n43228 & ~n43310;
  assign n43313 = ~n43228 & n59011;
  assign n43314 = ~n59011 & ~n43310;
  assign n43315 = n43228 & ~n59011;
  assign n43316 = ~n59012 & ~n59013;
  assign n43317 = ~n43310 & ~n43311;
  assign n43318 = n43215 & n59014;
  assign n43319 = ~n43215 & ~n59014;
  assign n43320 = ~n43318 & ~n43319;
  assign n43321 = n123 & ~n58533;
  assign n43322 = n128 & n39600;
  assign n43323 = n53444 & n39606;
  assign n43324 = n127 & n39603;
  assign n43325 = ~n43323 & ~n43324;
  assign n43326 = ~n43322 & n43325;
  assign n43327 = ~n123 & n43326;
  assign n43328 = n58533 & n43326;
  assign n43329 = ~n43327 & ~n43328;
  assign n43330 = ~n43321 & n43326;
  assign n43331 = pi26  & ~n59015;
  assign n43332 = ~pi26  & n59015;
  assign n43333 = ~n43331 & ~n43332;
  assign n43334 = n43320 & ~n43333;
  assign n43335 = ~n43320 & n43333;
  assign n43336 = n43320 & ~n43334;
  assign n43337 = n43320 & n43333;
  assign n43338 = ~n43333 & ~n43334;
  assign n43339 = ~n43320 & ~n43333;
  assign n43340 = ~n59016 & ~n59017;
  assign n43341 = ~n43334 & ~n43335;
  assign n43342 = ~n43214 & ~n59018;
  assign n43343 = n43214 & n59018;
  assign n43344 = ~n43214 & ~n43342;
  assign n43345 = ~n43214 & n59018;
  assign n43346 = ~n59018 & ~n43342;
  assign n43347 = n43214 & ~n59018;
  assign n43348 = ~n59019 & ~n59020;
  assign n43349 = ~n43342 & ~n43343;
  assign n43350 = ~n43213 & ~n59021;
  assign n43351 = n43213 & n59021;
  assign n43352 = ~n43213 & ~n43350;
  assign n43353 = ~n59021 & ~n43350;
  assign n43354 = ~n43352 & ~n43353;
  assign n43355 = ~n43350 & ~n43351;
  assign n43356 = n43200 & n59022;
  assign n43357 = ~n43200 & ~n59022;
  assign n43358 = ~n43356 & ~n43357;
  assign n43359 = n14413 & n41007;
  assign n43360 = n15921 & n39582;
  assign n43361 = n54719 & n39588;
  assign n43362 = n15901 & n39585;
  assign n43363 = ~n43361 & ~n43362;
  assign n43364 = ~n43360 & n43363;
  assign n43365 = ~n14413 & n43364;
  assign n43366 = ~n41007 & n43364;
  assign n43367 = ~n43365 & ~n43366;
  assign n43368 = ~n43359 & n43364;
  assign n43369 = pi20  & ~n59023;
  assign n43370 = ~pi20  & n59023;
  assign n43371 = ~n43369 & ~n43370;
  assign n43372 = n43358 & ~n43371;
  assign n43373 = ~n43358 & n43371;
  assign n43374 = n43358 & ~n43372;
  assign n43375 = n43358 & n43371;
  assign n43376 = ~n43371 & ~n43372;
  assign n43377 = ~n43358 & ~n43371;
  assign n43378 = ~n59024 & ~n59025;
  assign n43379 = ~n43372 & ~n43373;
  assign n43380 = ~n43199 & ~n59026;
  assign n43381 = n43199 & n59026;
  assign n43382 = ~n43199 & ~n43380;
  assign n43383 = ~n59026 & ~n43380;
  assign n43384 = ~n43382 & ~n43383;
  assign n43385 = ~n43380 & ~n43381;
  assign n43386 = ~n43198 & ~n59027;
  assign n43387 = n43198 & n59027;
  assign n43388 = ~n43198 & ~n43386;
  assign n43389 = ~n43198 & n59027;
  assign n43390 = ~n59027 & ~n43386;
  assign n43391 = n43198 & ~n59027;
  assign n43392 = ~n59028 & ~n59029;
  assign n43393 = ~n43386 & ~n43387;
  assign n43394 = n43185 & n59030;
  assign n43395 = ~n43185 & ~n59030;
  assign n43396 = ~n43394 & ~n43395;
  assign n43397 = n17265 & n41762;
  assign n43398 = n18588 & n39564;
  assign n43399 = n55041 & n39570;
  assign n43400 = n18556 & n39567;
  assign n43401 = ~n43399 & ~n43400;
  assign n43402 = ~n43398 & n43401;
  assign n43403 = ~n17265 & n43402;
  assign n43404 = ~n41762 & n43402;
  assign n43405 = ~n43403 & ~n43404;
  assign n43406 = ~n43397 & n43402;
  assign n43407 = pi14  & ~n59031;
  assign n43408 = ~pi14  & n59031;
  assign n43409 = ~n43407 & ~n43408;
  assign n43410 = n43396 & ~n43409;
  assign n43411 = ~n43396 & n43409;
  assign n43412 = n43396 & ~n43410;
  assign n43413 = n43396 & n43409;
  assign n43414 = ~n43409 & ~n43410;
  assign n43415 = ~n43396 & ~n43409;
  assign n43416 = ~n59032 & ~n59033;
  assign n43417 = ~n43410 & ~n43411;
  assign n43418 = ~n43184 & ~n59034;
  assign n43419 = n43184 & n59034;
  assign n43420 = ~n43184 & ~n43418;
  assign n43421 = ~n43184 & n59034;
  assign n43422 = ~n59034 & ~n43418;
  assign n43423 = n43184 & ~n59034;
  assign n43424 = ~n59035 & ~n59036;
  assign n43425 = ~n43418 & ~n43419;
  assign n43426 = ~n43183 & ~n59037;
  assign n43427 = n43183 & n59037;
  assign n43428 = ~n43183 & ~n43426;
  assign n43429 = ~n59037 & ~n43426;
  assign n43430 = ~n43428 & ~n43429;
  assign n43431 = ~n43426 & ~n43427;
  assign n43432 = n43170 & n59038;
  assign n43433 = ~n43170 & ~n59038;
  assign n43434 = ~n43432 & ~n43433;
  assign n43435 = n39753 & ~n39755;
  assign n43436 = ~n39756 & ~n43435;
  assign n43437 = n20085 & n43436;
  assign n43438 = n21269 & n39546;
  assign n43439 = n55472 & n39552;
  assign n43440 = n21237 & n39549;
  assign n43441 = ~n43439 & ~n43440;
  assign n43442 = ~n43438 & n43441;
  assign n43443 = ~n20085 & n43442;
  assign n43444 = ~n43436 & n43442;
  assign n43445 = ~n43443 & ~n43444;
  assign n43446 = ~n43437 & n43442;
  assign n43447 = pi8  & ~n59039;
  assign n43448 = ~pi8  & n59039;
  assign n43449 = ~n43447 & ~n43448;
  assign n43450 = n43434 & ~n43449;
  assign n43451 = ~n43434 & n43449;
  assign n43452 = n43434 & ~n43450;
  assign n43453 = n43434 & n43449;
  assign n43454 = ~n43449 & ~n43450;
  assign n43455 = ~n43434 & ~n43449;
  assign n43456 = ~n59040 & ~n59041;
  assign n43457 = ~n43450 & ~n43451;
  assign n43458 = ~n43169 & ~n59042;
  assign n43459 = n43169 & n59042;
  assign n43460 = ~n43169 & ~n43458;
  assign n43461 = ~n59042 & ~n43458;
  assign n43462 = ~n43460 & ~n43461;
  assign n43463 = ~n43458 & ~n43459;
  assign n43464 = ~n39956 & ~n59043;
  assign n43465 = n39763 & ~n39765;
  assign n43466 = ~n39763 & ~n58471;
  assign n43467 = ~n39764 & n39769;
  assign n43468 = ~n43466 & ~n43467;
  assign n43469 = ~n58471 & ~n43465;
  assign n43470 = n77 & ~n59044;
  assign n43471 = n24302 & n39543;
  assign n43472 = n21969 & n39546;
  assign n43473 = n23459 & n39440;
  assign n43474 = ~n43472 & ~n43473;
  assign n43475 = ~n43471 & n43474;
  assign n43476 = ~n43470 & n43475;
  assign n43477 = pi5  & ~n43476;
  assign n43478 = ~n43476 & ~n43477;
  assign n43479 = ~pi5  & ~n43476;
  assign n43480 = pi5  & ~n43477;
  assign n43481 = pi5  & n43476;
  assign n43482 = ~n59045 & ~n59046;
  assign n43483 = n43160 & n58993;
  assign n43484 = ~n43160 & ~n43168;
  assign n43485 = ~n43160 & n58993;
  assign n43486 = ~n58993 & ~n43168;
  assign n43487 = n43160 & ~n58993;
  assign n43488 = ~n59047 & ~n59048;
  assign n43489 = ~n43168 & ~n43483;
  assign n43490 = ~n43482 & ~n59049;
  assign n43491 = n39757 & ~n39759;
  assign n43492 = ~n39757 & ~n58470;
  assign n43493 = ~n39758 & n39763;
  assign n43494 = ~n43492 & ~n43493;
  assign n43495 = ~n58470 & ~n43491;
  assign n43496 = n77 & ~n59050;
  assign n43497 = n24302 & n39440;
  assign n43498 = n21969 & n39549;
  assign n43499 = n23459 & n39546;
  assign n43500 = ~n43498 & ~n43499;
  assign n43501 = ~n43497 & n43500;
  assign n43502 = ~n43496 & n43501;
  assign n43503 = pi5  & ~n43502;
  assign n43504 = ~n43502 & ~n43503;
  assign n43505 = ~pi5  & ~n43502;
  assign n43506 = pi5  & ~n43503;
  assign n43507 = pi5  & n43502;
  assign n43508 = ~n59051 & ~n59052;
  assign n43509 = n43151 & n58990;
  assign n43510 = ~n43151 & ~n43159;
  assign n43511 = ~n43151 & n58990;
  assign n43512 = ~n58990 & ~n43159;
  assign n43513 = n43151 & ~n58990;
  assign n43514 = ~n59053 & ~n59054;
  assign n43515 = ~n43159 & ~n43509;
  assign n43516 = ~n43508 & ~n59055;
  assign n43517 = n43142 & n58987;
  assign n43518 = ~n43150 & ~n43517;
  assign n43519 = n77 & n43436;
  assign n43520 = n24302 & n39546;
  assign n43521 = n21969 & n39552;
  assign n43522 = n23459 & n39549;
  assign n43523 = ~n43521 & ~n43522;
  assign n43524 = ~n43520 & n43523;
  assign n43525 = ~n77 & n43524;
  assign n43526 = ~n43436 & n43524;
  assign n43527 = ~n43525 & ~n43526;
  assign n43528 = ~n43519 & n43524;
  assign n43529 = pi5  & ~n59056;
  assign n43530 = ~pi5  & n59056;
  assign n43531 = ~n43529 & ~n43530;
  assign n43532 = n43518 & ~n43531;
  assign n43533 = n43135 & n58984;
  assign n43534 = ~n43141 & ~n43533;
  assign n43535 = n77 & ~n58889;
  assign n43536 = n24302 & n39549;
  assign n43537 = n21969 & n39555;
  assign n43538 = n23459 & n39552;
  assign n43539 = ~n43537 & ~n43538;
  assign n43540 = ~n43536 & n43539;
  assign n43541 = ~n77 & n43540;
  assign n43542 = n58889 & n43540;
  assign n43543 = ~n43541 & ~n43542;
  assign n43544 = ~n43535 & n43540;
  assign n43545 = pi5  & ~n59057;
  assign n43546 = ~pi5  & n59057;
  assign n43547 = ~n43545 & ~n43546;
  assign n43548 = n43534 & ~n43547;
  assign n43549 = n77 & ~n58891;
  assign n43550 = n24302 & n39552;
  assign n43551 = n21969 & n39558;
  assign n43552 = n23459 & n39555;
  assign n43553 = ~n43551 & ~n43552;
  assign n43554 = ~n43550 & n43553;
  assign n43555 = ~n43549 & n43554;
  assign n43556 = pi5  & ~n43555;
  assign n43557 = ~n43555 & ~n43556;
  assign n43558 = ~pi5  & ~n43555;
  assign n43559 = pi5  & ~n43556;
  assign n43560 = pi5  & n43555;
  assign n43561 = ~n59058 & ~n59059;
  assign n43562 = n43131 & ~n43133;
  assign n43563 = ~n43134 & ~n43562;
  assign n43564 = ~n43561 & n43563;
  assign n43565 = n77 & n42574;
  assign n43566 = n24302 & n39555;
  assign n43567 = n21969 & n39561;
  assign n43568 = n23459 & n39558;
  assign n43569 = ~n43567 & ~n43568;
  assign n43570 = ~n43566 & n43569;
  assign n43571 = ~n43565 & n43570;
  assign n43572 = pi5  & ~n43571;
  assign n43573 = ~n43571 & ~n43572;
  assign n43574 = ~pi5  & ~n43571;
  assign n43575 = pi5  & ~n43572;
  assign n43576 = pi5  & n43571;
  assign n43577 = ~n59060 & ~n59061;
  assign n43578 = n43122 & n58983;
  assign n43579 = ~n43122 & ~n43130;
  assign n43580 = ~n58983 & ~n43130;
  assign n43581 = ~n43579 & ~n43580;
  assign n43582 = ~n43130 & ~n43578;
  assign n43583 = ~n43577 & ~n59062;
  assign n43584 = n77 & ~n58849;
  assign n43585 = n24302 & n39558;
  assign n43586 = n21969 & n39564;
  assign n43587 = n23459 & n39561;
  assign n43588 = ~n43586 & ~n43587;
  assign n43589 = ~n43585 & n43588;
  assign n43590 = ~n43584 & n43589;
  assign n43591 = pi5  & ~n43590;
  assign n43592 = ~n43590 & ~n43591;
  assign n43593 = ~pi5  & ~n43590;
  assign n43594 = pi5  & ~n43591;
  assign n43595 = pi5  & n43590;
  assign n43596 = ~n59063 & ~n59064;
  assign n43597 = n43113 & n58980;
  assign n43598 = ~n43113 & ~n43121;
  assign n43599 = ~n43113 & n58980;
  assign n43600 = ~n58980 & ~n43121;
  assign n43601 = n43113 & ~n58980;
  assign n43602 = ~n59065 & ~n59066;
  assign n43603 = ~n43121 & ~n43597;
  assign n43604 = ~n43596 & ~n59067;
  assign n43605 = n43104 & n58977;
  assign n43606 = ~n43112 & ~n43605;
  assign n43607 = n77 & ~n58493;
  assign n43608 = n24302 & n39561;
  assign n43609 = n21969 & n39567;
  assign n43610 = n23459 & n39564;
  assign n43611 = ~n43609 & ~n43610;
  assign n43612 = ~n43608 & n43611;
  assign n43613 = ~n77 & n43612;
  assign n43614 = n58493 & n43612;
  assign n43615 = ~n43613 & ~n43614;
  assign n43616 = ~n43607 & n43612;
  assign n43617 = pi5  & ~n59068;
  assign n43618 = ~pi5  & n59068;
  assign n43619 = ~n43617 & ~n43618;
  assign n43620 = n43606 & ~n43619;
  assign n43621 = n43097 & n58974;
  assign n43622 = ~n43103 & ~n43621;
  assign n43623 = n77 & n41762;
  assign n43624 = n24302 & n39564;
  assign n43625 = n21969 & n39570;
  assign n43626 = n23459 & n39567;
  assign n43627 = ~n43625 & ~n43626;
  assign n43628 = ~n43624 & n43627;
  assign n43629 = ~n77 & n43628;
  assign n43630 = ~n41762 & n43628;
  assign n43631 = ~n43629 & ~n43630;
  assign n43632 = ~n43623 & n43628;
  assign n43633 = pi5  & ~n59069;
  assign n43634 = ~pi5  & n59069;
  assign n43635 = ~n43633 & ~n43634;
  assign n43636 = n43622 & ~n43635;
  assign n43637 = n43088 & n58973;
  assign n43638 = ~n43096 & ~n43637;
  assign n43639 = n77 & ~n58766;
  assign n43640 = n24302 & n39567;
  assign n43641 = n21969 & n39573;
  assign n43642 = n23459 & n39570;
  assign n43643 = ~n43641 & ~n43642;
  assign n43644 = ~n43640 & n43643;
  assign n43645 = ~n77 & n43644;
  assign n43646 = n58766 & n43644;
  assign n43647 = ~n43645 & ~n43646;
  assign n43648 = ~n43639 & n43644;
  assign n43649 = pi5  & ~n59070;
  assign n43650 = ~pi5  & n59070;
  assign n43651 = ~n43649 & ~n43650;
  assign n43652 = n43638 & ~n43651;
  assign n43653 = n77 & ~n58759;
  assign n43654 = n24302 & n39570;
  assign n43655 = n21969 & n39576;
  assign n43656 = n23459 & n39573;
  assign n43657 = ~n43655 & ~n43656;
  assign n43658 = ~n43654 & n43657;
  assign n43659 = ~n43653 & n43658;
  assign n43660 = pi5  & ~n43659;
  assign n43661 = ~n43659 & ~n43660;
  assign n43662 = ~pi5  & ~n43659;
  assign n43663 = pi5  & ~n43660;
  assign n43664 = pi5  & n43659;
  assign n43665 = ~n59071 & ~n59072;
  assign n43666 = n43084 & ~n43086;
  assign n43667 = ~n43087 & ~n43666;
  assign n43668 = ~n43665 & n43667;
  assign n43669 = n77 & n39976;
  assign n43670 = n24302 & n39573;
  assign n43671 = n21969 & n39579;
  assign n43672 = n23459 & n39576;
  assign n43673 = ~n43671 & ~n43672;
  assign n43674 = ~n43670 & n43673;
  assign n43675 = ~n43669 & n43674;
  assign n43676 = pi5  & ~n43675;
  assign n43677 = ~n43675 & ~n43676;
  assign n43678 = ~pi5  & ~n43675;
  assign n43679 = pi5  & ~n43676;
  assign n43680 = pi5  & n43675;
  assign n43681 = ~n59073 & ~n59074;
  assign n43682 = n43075 & n58970;
  assign n43683 = ~n43075 & ~n43083;
  assign n43684 = ~n43075 & n58970;
  assign n43685 = ~n58970 & ~n43083;
  assign n43686 = n43075 & ~n58970;
  assign n43687 = ~n59075 & ~n59076;
  assign n43688 = ~n43083 & ~n43682;
  assign n43689 = ~n43681 & ~n59077;
  assign n43690 = n77 & ~n58653;
  assign n43691 = n24302 & n39576;
  assign n43692 = n21969 & n39582;
  assign n43693 = n23459 & n39579;
  assign n43694 = ~n43692 & ~n43693;
  assign n43695 = ~n43691 & n43694;
  assign n43696 = ~n43690 & n43695;
  assign n43697 = pi5  & ~n43696;
  assign n43698 = ~n43696 & ~n43697;
  assign n43699 = ~pi5  & ~n43696;
  assign n43700 = pi5  & ~n43697;
  assign n43701 = pi5  & n43696;
  assign n43702 = ~n59078 & ~n59079;
  assign n43703 = n43066 & n58967;
  assign n43704 = ~n43066 & ~n43074;
  assign n43705 = ~n58967 & ~n43074;
  assign n43706 = ~n43704 & ~n43705;
  assign n43707 = ~n43074 & ~n43703;
  assign n43708 = ~n43702 & ~n59080;
  assign n43709 = n43057 & n58964;
  assign n43710 = ~n43065 & ~n43709;
  assign n43711 = n77 & ~n58657;
  assign n43712 = n24302 & n39579;
  assign n43713 = n21969 & n39585;
  assign n43714 = n23459 & n39582;
  assign n43715 = ~n43713 & ~n43714;
  assign n43716 = ~n43712 & n43715;
  assign n43717 = ~n77 & n43716;
  assign n43718 = n58657 & n43716;
  assign n43719 = ~n43717 & ~n43718;
  assign n43720 = ~n43711 & n43716;
  assign n43721 = pi5  & ~n59081;
  assign n43722 = ~pi5  & n59081;
  assign n43723 = ~n43721 & ~n43722;
  assign n43724 = n43710 & ~n43723;
  assign n43725 = n43048 & n58961;
  assign n43726 = ~n43056 & ~n43725;
  assign n43727 = n77 & n41007;
  assign n43728 = n24302 & n39582;
  assign n43729 = n21969 & n39588;
  assign n43730 = n23459 & n39585;
  assign n43731 = ~n43729 & ~n43730;
  assign n43732 = ~n43728 & n43731;
  assign n43733 = ~n77 & n43732;
  assign n43734 = ~n41007 & n43732;
  assign n43735 = ~n43733 & ~n43734;
  assign n43736 = ~n43727 & n43732;
  assign n43737 = pi5  & ~n59082;
  assign n43738 = ~pi5  & n59082;
  assign n43739 = ~n43737 & ~n43738;
  assign n43740 = n43726 & ~n43739;
  assign n43741 = n43041 & n58958;
  assign n43742 = ~n43047 & ~n43741;
  assign n43743 = n77 & ~n58583;
  assign n43744 = n24302 & n39585;
  assign n43745 = n21969 & n39591;
  assign n43746 = n23459 & n39588;
  assign n43747 = ~n43745 & ~n43746;
  assign n43748 = ~n43744 & n43747;
  assign n43749 = ~n77 & n43748;
  assign n43750 = n58583 & n43748;
  assign n43751 = ~n43749 & ~n43750;
  assign n43752 = ~n43743 & n43748;
  assign n43753 = pi5  & ~n59083;
  assign n43754 = ~pi5  & n59083;
  assign n43755 = ~n43753 & ~n43754;
  assign n43756 = n43742 & ~n43755;
  assign n43757 = n77 & ~n58585;
  assign n43758 = n24302 & n39588;
  assign n43759 = n21969 & n39594;
  assign n43760 = n23459 & n39591;
  assign n43761 = ~n43759 & ~n43760;
  assign n43762 = ~n43758 & n43761;
  assign n43763 = ~n43757 & n43762;
  assign n43764 = pi5  & ~n43763;
  assign n43765 = ~n43763 & ~n43764;
  assign n43766 = ~pi5  & ~n43763;
  assign n43767 = pi5  & ~n43764;
  assign n43768 = pi5  & n43763;
  assign n43769 = ~n59084 & ~n59085;
  assign n43770 = n43037 & ~n43039;
  assign n43771 = ~n43040 & ~n43770;
  assign n43772 = ~n43769 & n43771;
  assign n43773 = n77 & n40616;
  assign n43774 = n24302 & n39591;
  assign n43775 = n21969 & n39597;
  assign n43776 = n23459 & n39594;
  assign n43777 = ~n43775 & ~n43776;
  assign n43778 = ~n43774 & n43777;
  assign n43779 = ~n43773 & n43778;
  assign n43780 = pi5  & ~n43779;
  assign n43781 = ~n43779 & ~n43780;
  assign n43782 = ~pi5  & ~n43779;
  assign n43783 = pi5  & ~n43780;
  assign n43784 = pi5  & n43779;
  assign n43785 = ~n59086 & ~n59087;
  assign n43786 = n43028 & n58957;
  assign n43787 = ~n43028 & ~n43036;
  assign n43788 = ~n58957 & ~n43036;
  assign n43789 = ~n43787 & ~n43788;
  assign n43790 = ~n43036 & ~n43786;
  assign n43791 = ~n43785 & ~n59088;
  assign n43792 = n77 & n40476;
  assign n43793 = n24302 & n39594;
  assign n43794 = n21969 & n39600;
  assign n43795 = n23459 & n39597;
  assign n43796 = ~n43794 & ~n43795;
  assign n43797 = ~n43793 & n43796;
  assign n43798 = ~n43792 & n43797;
  assign n43799 = pi5  & ~n43798;
  assign n43800 = ~n43798 & ~n43799;
  assign n43801 = ~pi5  & ~n43798;
  assign n43802 = pi5  & ~n43799;
  assign n43803 = pi5  & n43798;
  assign n43804 = ~n59089 & ~n59090;
  assign n43805 = n43019 & n58954;
  assign n43806 = ~n43019 & ~n43027;
  assign n43807 = ~n43019 & n58954;
  assign n43808 = ~n58954 & ~n43027;
  assign n43809 = n43019 & ~n58954;
  assign n43810 = ~n59091 & ~n59092;
  assign n43811 = ~n43027 & ~n43805;
  assign n43812 = ~n43804 & ~n59093;
  assign n43813 = n43010 & n58951;
  assign n43814 = ~n43018 & ~n43813;
  assign n43815 = n77 & n40247;
  assign n43816 = n24302 & n39597;
  assign n43817 = n21969 & n39603;
  assign n43818 = n23459 & n39600;
  assign n43819 = ~n43817 & ~n43818;
  assign n43820 = ~n43816 & n43819;
  assign n43821 = ~n77 & n43820;
  assign n43822 = ~n40247 & n43820;
  assign n43823 = ~n43821 & ~n43822;
  assign n43824 = ~n43815 & n43820;
  assign n43825 = pi5  & ~n59094;
  assign n43826 = ~pi5  & n59094;
  assign n43827 = ~n43825 & ~n43826;
  assign n43828 = n43814 & ~n43827;
  assign n43829 = n43006 & ~n43008;
  assign n43830 = ~n43009 & ~n43829;
  assign n43831 = n77 & ~n58533;
  assign n43832 = n24302 & n39600;
  assign n43833 = n21969 & n39606;
  assign n43834 = n23459 & n39603;
  assign n43835 = ~n43833 & ~n43834;
  assign n43836 = ~n43832 & n43835;
  assign n43837 = ~n77 & n43836;
  assign n43838 = n58533 & n43836;
  assign n43839 = ~n43837 & ~n43838;
  assign n43840 = ~n43831 & n43836;
  assign n43841 = pi5  & ~n59095;
  assign n43842 = ~pi5  & n59095;
  assign n43843 = ~n43841 & ~n43842;
  assign n43844 = n43830 & ~n43843;
  assign n43845 = n42997 & n58948;
  assign n43846 = ~n43005 & ~n43845;
  assign n43847 = n77 & n40286;
  assign n43848 = n24302 & n39603;
  assign n43849 = n21969 & n39609;
  assign n43850 = n23459 & n39606;
  assign n43851 = ~n43849 & ~n43850;
  assign n43852 = ~n43848 & n43851;
  assign n43853 = ~n77 & n43852;
  assign n43854 = ~n40286 & n43852;
  assign n43855 = ~n43853 & ~n43854;
  assign n43856 = ~n43847 & n43852;
  assign n43857 = pi5  & ~n59096;
  assign n43858 = ~pi5  & n59096;
  assign n43859 = ~n43857 & ~n43858;
  assign n43860 = n43846 & ~n43859;
  assign n43861 = n77 & n40183;
  assign n43862 = n24302 & n39606;
  assign n43863 = n21969 & n39612;
  assign n43864 = n23459 & n39609;
  assign n43865 = ~n43863 & ~n43864;
  assign n43866 = ~n43862 & n43865;
  assign n43867 = ~n43861 & n43866;
  assign n43868 = pi5  & ~n43867;
  assign n43869 = ~n43867 & ~n43868;
  assign n43870 = ~pi5  & ~n43867;
  assign n43871 = pi5  & ~n43868;
  assign n43872 = pi5  & n43867;
  assign n43873 = ~n59097 & ~n59098;
  assign n43874 = n42993 & ~n42995;
  assign n43875 = ~n42996 & ~n43874;
  assign n43876 = ~n43873 & n43875;
  assign n43877 = n77 & n39991;
  assign n43878 = n24302 & n39609;
  assign n43879 = n21969 & n39615;
  assign n43880 = n23459 & n39612;
  assign n43881 = ~n43879 & ~n43880;
  assign n43882 = ~n43878 & n43881;
  assign n43883 = ~n77 & n43882;
  assign n43884 = ~n39991 & n43882;
  assign n43885 = ~n43883 & ~n43884;
  assign n43886 = ~n43877 & n43882;
  assign n43887 = pi5  & ~n59099;
  assign n43888 = ~pi5  & n59099;
  assign n43889 = ~n43887 & ~n43888;
  assign n43890 = n42984 & n58945;
  assign n43891 = ~n58945 & ~n42992;
  assign n43892 = ~n42984 & ~n42992;
  assign n43893 = ~n43891 & ~n43892;
  assign n43894 = ~n42992 & ~n43890;
  assign n43895 = ~n43889 & ~n59100;
  assign n43896 = n77 & n40071;
  assign n43897 = n24302 & n39612;
  assign n43898 = n21969 & n39618;
  assign n43899 = n23459 & n39615;
  assign n43900 = ~n43898 & ~n43899;
  assign n43901 = ~n43897 & n43900;
  assign n43902 = ~n43896 & n43901;
  assign n43903 = pi5  & ~n43902;
  assign n43904 = ~n43902 & ~n43903;
  assign n43905 = ~pi5  & ~n43902;
  assign n43906 = pi5  & ~n43903;
  assign n43907 = pi5  & n43902;
  assign n43908 = ~n59101 & ~n59102;
  assign n43909 = pi8  & ~n58938;
  assign n43910 = ~n58939 & ~n43909;
  assign n43911 = n58939 & n43909;
  assign n43912 = ~n58938 & n42968;
  assign n43913 = ~n58940 & ~n43912;
  assign n43914 = ~n43910 & ~n43911;
  assign n43915 = ~n43908 & n59103;
  assign n43916 = n77 & n40093;
  assign n43917 = n24302 & n39615;
  assign n43918 = n21969 & n39621;
  assign n43919 = n23459 & n39618;
  assign n43920 = ~n43918 & ~n43919;
  assign n43921 = ~n43917 & n43920;
  assign n43922 = ~n77 & n43921;
  assign n43923 = ~n40093 & n43921;
  assign n43924 = ~n43922 & ~n43923;
  assign n43925 = ~n43916 & n43921;
  assign n43926 = pi5  & ~n59104;
  assign n43927 = ~pi5  & n59104;
  assign n43928 = ~n43926 & ~n43927;
  assign n43929 = pi8  & n42948;
  assign n43930 = ~n42947 & n43929;
  assign n43931 = n42947 & ~n43929;
  assign n43932 = ~n42949 & n42953;
  assign n43933 = ~n58938 & ~n43932;
  assign n43934 = ~n43930 & ~n43931;
  assign n43935 = ~n43928 & n59105;
  assign n43936 = n77 & ~n40023;
  assign n43937 = n23459 & ~n58457;
  assign n43938 = n24302 & n39626;
  assign n43939 = ~n43937 & ~n43938;
  assign n43940 = ~n43936 & n43939;
  assign n43941 = n53439 & ~n58457;
  assign n43942 = pi5  & ~n43941;
  assign n43943 = pi5  & ~n43940;
  assign n43944 = pi5  & ~n43943;
  assign n43945 = ~n43940 & ~n43943;
  assign n43946 = ~n43944 & ~n43945;
  assign n43947 = n43942 & ~n43946;
  assign n43948 = n43940 & n43942;
  assign n43949 = n77 & ~n40039;
  assign n43950 = n24302 & n39621;
  assign n43951 = n21969 & ~n58457;
  assign n43952 = n23459 & n39626;
  assign n43953 = ~n43951 & ~n43952;
  assign n43954 = ~n43950 & n43953;
  assign n43955 = ~n77 & n43954;
  assign n43956 = n40039 & n43954;
  assign n43957 = ~n43955 & ~n43956;
  assign n43958 = ~n43949 & n43954;
  assign n43959 = pi5  & ~n59107;
  assign n43960 = ~pi5  & n59107;
  assign n43961 = ~n43959 & ~n43960;
  assign n43962 = n59106 & ~n43961;
  assign n43963 = n59106 & ~n59107;
  assign n43964 = n42948 & n59108;
  assign n43965 = n77 & n40006;
  assign n43966 = n24302 & n39618;
  assign n43967 = n21969 & n39626;
  assign n43968 = n23459 & n39621;
  assign n43969 = ~n43967 & ~n43968;
  assign n43970 = ~n43966 & n43969;
  assign n43971 = ~n43965 & n43970;
  assign n43972 = pi5  & ~n43971;
  assign n43973 = pi5  & ~n43972;
  assign n43974 = pi5  & n43971;
  assign n43975 = ~n43971 & ~n43972;
  assign n43976 = ~pi5  & ~n43971;
  assign n43977 = ~n59109 & ~n59110;
  assign n43978 = ~n42948 & ~n59108;
  assign n43979 = n59108 & ~n43964;
  assign n43980 = ~n42948 & n59108;
  assign n43981 = n42948 & ~n43964;
  assign n43982 = n42948 & ~n59108;
  assign n43983 = ~n59111 & ~n59112;
  assign n43984 = ~n43964 & ~n43978;
  assign n43985 = ~n43977 & ~n59113;
  assign n43986 = ~n43964 & ~n43985;
  assign n43987 = n43928 & ~n59105;
  assign n43988 = ~n43935 & ~n43987;
  assign n43989 = ~n43986 & n43988;
  assign n43990 = ~n43935 & ~n43989;
  assign n43991 = n43908 & ~n59103;
  assign n43992 = ~n43908 & ~n43915;
  assign n43993 = ~n43908 & ~n59103;
  assign n43994 = n59103 & ~n43915;
  assign n43995 = n43908 & n59103;
  assign n43996 = ~n59114 & ~n59115;
  assign n43997 = ~n43915 & ~n43991;
  assign n43998 = ~n43990 & ~n59116;
  assign n43999 = ~n43915 & ~n43998;
  assign n44000 = n43889 & n59100;
  assign n44001 = ~n43895 & ~n44000;
  assign n44002 = ~n43999 & n44001;
  assign n44003 = ~n43895 & ~n44002;
  assign n44004 = n43873 & ~n43875;
  assign n44005 = ~n43873 & ~n43876;
  assign n44006 = ~n43873 & ~n43875;
  assign n44007 = n43875 & ~n43876;
  assign n44008 = n43873 & n43875;
  assign n44009 = ~n59117 & ~n59118;
  assign n44010 = ~n43876 & ~n44004;
  assign n44011 = ~n44003 & ~n59119;
  assign n44012 = ~n43876 & ~n44011;
  assign n44013 = ~n43846 & n43859;
  assign n44014 = n43846 & ~n43860;
  assign n44015 = n43846 & n43859;
  assign n44016 = ~n43859 & ~n43860;
  assign n44017 = ~n43846 & ~n43859;
  assign n44018 = ~n59120 & ~n59121;
  assign n44019 = ~n43860 & ~n44013;
  assign n44020 = ~n44012 & ~n59122;
  assign n44021 = ~n43860 & ~n44020;
  assign n44022 = ~n43830 & n43843;
  assign n44023 = n43830 & ~n43844;
  assign n44024 = n43830 & n43843;
  assign n44025 = ~n43843 & ~n43844;
  assign n44026 = ~n43830 & ~n43843;
  assign n44027 = ~n59123 & ~n59124;
  assign n44028 = ~n43844 & ~n44022;
  assign n44029 = ~n44021 & ~n59125;
  assign n44030 = ~n43844 & ~n44029;
  assign n44031 = ~n43814 & n43827;
  assign n44032 = ~n43828 & ~n44031;
  assign n44033 = ~n44030 & n44032;
  assign n44034 = ~n43828 & ~n44033;
  assign n44035 = n43804 & n59093;
  assign n44036 = ~n43804 & ~n43812;
  assign n44037 = ~n59093 & ~n43812;
  assign n44038 = ~n44036 & ~n44037;
  assign n44039 = ~n43812 & ~n44035;
  assign n44040 = ~n44034 & ~n59126;
  assign n44041 = ~n43812 & ~n44040;
  assign n44042 = n43785 & n59088;
  assign n44043 = ~n43785 & ~n43791;
  assign n44044 = ~n43785 & n59088;
  assign n44045 = ~n59088 & ~n43791;
  assign n44046 = n43785 & ~n59088;
  assign n44047 = ~n59127 & ~n59128;
  assign n44048 = ~n43791 & ~n44042;
  assign n44049 = ~n44041 & ~n59129;
  assign n44050 = ~n43791 & ~n44049;
  assign n44051 = n43769 & ~n43771;
  assign n44052 = ~n43769 & ~n43772;
  assign n44053 = ~n43769 & ~n43771;
  assign n44054 = n43771 & ~n43772;
  assign n44055 = n43769 & n43771;
  assign n44056 = ~n59130 & ~n59131;
  assign n44057 = ~n43772 & ~n44051;
  assign n44058 = ~n44050 & ~n59132;
  assign n44059 = ~n43772 & ~n44058;
  assign n44060 = ~n43742 & n43755;
  assign n44061 = n43742 & ~n43756;
  assign n44062 = n43742 & n43755;
  assign n44063 = ~n43755 & ~n43756;
  assign n44064 = ~n43742 & ~n43755;
  assign n44065 = ~n59133 & ~n59134;
  assign n44066 = ~n43756 & ~n44060;
  assign n44067 = ~n44059 & ~n59135;
  assign n44068 = ~n43756 & ~n44067;
  assign n44069 = ~n43726 & n43739;
  assign n44070 = n43726 & ~n43740;
  assign n44071 = n43726 & n43739;
  assign n44072 = ~n43739 & ~n43740;
  assign n44073 = ~n43726 & ~n43739;
  assign n44074 = ~n59136 & ~n59137;
  assign n44075 = ~n43740 & ~n44069;
  assign n44076 = ~n44068 & ~n59138;
  assign n44077 = ~n43740 & ~n44076;
  assign n44078 = ~n43710 & n43723;
  assign n44079 = ~n43724 & ~n44078;
  assign n44080 = ~n44077 & n44079;
  assign n44081 = ~n43724 & ~n44080;
  assign n44082 = n43702 & n59080;
  assign n44083 = ~n43702 & ~n43708;
  assign n44084 = ~n43702 & n59080;
  assign n44085 = ~n59080 & ~n43708;
  assign n44086 = n43702 & ~n59080;
  assign n44087 = ~n59139 & ~n59140;
  assign n44088 = ~n43708 & ~n44082;
  assign n44089 = ~n44081 & ~n59141;
  assign n44090 = ~n43708 & ~n44089;
  assign n44091 = n43681 & n59077;
  assign n44092 = ~n43681 & ~n43689;
  assign n44093 = ~n59077 & ~n43689;
  assign n44094 = ~n44092 & ~n44093;
  assign n44095 = ~n43689 & ~n44091;
  assign n44096 = ~n44090 & ~n59142;
  assign n44097 = ~n43689 & ~n44096;
  assign n44098 = n43665 & ~n43667;
  assign n44099 = ~n43665 & ~n43668;
  assign n44100 = ~n43665 & ~n43667;
  assign n44101 = n43667 & ~n43668;
  assign n44102 = n43665 & n43667;
  assign n44103 = ~n59143 & ~n59144;
  assign n44104 = ~n43668 & ~n44098;
  assign n44105 = ~n44097 & ~n59145;
  assign n44106 = ~n43668 & ~n44105;
  assign n44107 = ~n43638 & n43651;
  assign n44108 = n43638 & ~n43652;
  assign n44109 = n43638 & n43651;
  assign n44110 = ~n43651 & ~n43652;
  assign n44111 = ~n43638 & ~n43651;
  assign n44112 = ~n59146 & ~n59147;
  assign n44113 = ~n43652 & ~n44107;
  assign n44114 = ~n44106 & ~n59148;
  assign n44115 = ~n43652 & ~n44114;
  assign n44116 = ~n43622 & n43635;
  assign n44117 = n43622 & ~n43636;
  assign n44118 = n43622 & n43635;
  assign n44119 = ~n43635 & ~n43636;
  assign n44120 = ~n43622 & ~n43635;
  assign n44121 = ~n59149 & ~n59150;
  assign n44122 = ~n43636 & ~n44116;
  assign n44123 = ~n44115 & ~n59151;
  assign n44124 = ~n43636 & ~n44123;
  assign n44125 = ~n43606 & n43619;
  assign n44126 = ~n43620 & ~n44125;
  assign n44127 = ~n44124 & n44126;
  assign n44128 = ~n43620 & ~n44127;
  assign n44129 = n43596 & n59067;
  assign n44130 = ~n43596 & ~n43604;
  assign n44131 = ~n59067 & ~n43604;
  assign n44132 = ~n44130 & ~n44131;
  assign n44133 = ~n43604 & ~n44129;
  assign n44134 = ~n44128 & ~n59152;
  assign n44135 = ~n43604 & ~n44134;
  assign n44136 = n43577 & n59062;
  assign n44137 = ~n43577 & ~n43583;
  assign n44138 = ~n43577 & n59062;
  assign n44139 = ~n59062 & ~n43583;
  assign n44140 = n43577 & ~n59062;
  assign n44141 = ~n59153 & ~n59154;
  assign n44142 = ~n43583 & ~n44136;
  assign n44143 = ~n44135 & ~n59155;
  assign n44144 = ~n43583 & ~n44143;
  assign n44145 = n43561 & ~n43563;
  assign n44146 = ~n43561 & ~n43564;
  assign n44147 = ~n43561 & ~n43563;
  assign n44148 = n43563 & ~n43564;
  assign n44149 = n43561 & n43563;
  assign n44150 = ~n59156 & ~n59157;
  assign n44151 = ~n43564 & ~n44145;
  assign n44152 = ~n44144 & ~n59158;
  assign n44153 = ~n43564 & ~n44152;
  assign n44154 = ~n43534 & n43547;
  assign n44155 = n43534 & ~n43548;
  assign n44156 = n43534 & n43547;
  assign n44157 = ~n43547 & ~n43548;
  assign n44158 = ~n43534 & ~n43547;
  assign n44159 = ~n59159 & ~n59160;
  assign n44160 = ~n43548 & ~n44154;
  assign n44161 = ~n44153 & ~n59161;
  assign n44162 = ~n43548 & ~n44161;
  assign n44163 = ~n43518 & n43531;
  assign n44164 = ~n43532 & ~n44163;
  assign n44165 = ~n44162 & n44164;
  assign n44166 = ~n43532 & ~n44165;
  assign n44167 = n43508 & n59055;
  assign n44168 = ~n43508 & ~n43516;
  assign n44169 = ~n59055 & ~n43516;
  assign n44170 = ~n44168 & ~n44169;
  assign n44171 = ~n43516 & ~n44167;
  assign n44172 = ~n44166 & ~n59162;
  assign n44173 = ~n43516 & ~n44172;
  assign n44174 = n43482 & n59049;
  assign n44175 = ~n43482 & ~n43490;
  assign n44176 = ~n59049 & ~n43490;
  assign n44177 = ~n44175 & ~n44176;
  assign n44178 = ~n43490 & ~n44174;
  assign n44179 = ~n44173 & ~n59163;
  assign n44180 = ~n43490 & ~n44179;
  assign n44181 = n39956 & n59043;
  assign n44182 = ~n39956 & ~n43464;
  assign n44183 = ~n39956 & n59043;
  assign n44184 = ~n59043 & ~n43464;
  assign n44185 = n39956 & ~n59043;
  assign n44186 = ~n59164 & ~n59165;
  assign n44187 = ~n43464 & ~n44181;
  assign n44188 = ~n44180 & ~n59166;
  assign n44189 = ~n43464 & ~n44188;
  assign n44190 = ~n39938 & ~n39941;
  assign n44191 = ~n39931 & ~n39935;
  assign n44192 = n123 & n28624;
  assign n44193 = n127 & ~n26537;
  assign n44194 = n53444 & n26242;
  assign n44195 = ~n128 & ~n44194;
  assign n44196 = ~n44193 & ~n44194;
  assign n44197 = ~n128 & n44196;
  assign n44198 = ~n44193 & n44195;
  assign n44199 = ~n44192 & n59167;
  assign n44200 = pi26  & ~n44199;
  assign n44201 = pi26  & ~n44200;
  assign n44202 = pi26  & n44199;
  assign n44203 = ~n44199 & ~n44200;
  assign n44204 = ~pi26  & ~n44199;
  assign n44205 = ~n59168 & ~n59169;
  assign n44206 = ~n39900 & n39915;
  assign n44207 = ~n39900 & ~n39916;
  assign n44208 = ~n39901 & ~n44206;
  assign n44209 = ~n44205 & ~n59170;
  assign n44210 = n44205 & n59170;
  assign n44211 = ~n59170 & ~n44209;
  assign n44212 = n44205 & ~n59170;
  assign n44213 = ~n44205 & ~n44209;
  assign n44214 = ~n44205 & n59170;
  assign n44215 = ~n59171 & ~n59172;
  assign n44216 = ~n44209 & ~n44210;
  assign n44217 = ~n39889 & ~n39897;
  assign n44218 = ~n221 & ~n1881;
  assign n44219 = n358 & n44218;
  assign n44220 = n3272 & n3536;
  assign n44221 = n44219 & n44220;
  assign n44222 = n55106 & n44221;
  assign n44223 = n895 & n1078;
  assign n44224 = n12008 & n17997;
  assign n44225 = n44223 & n44224;
  assign n44226 = n53664 & n44225;
  assign n44227 = ~n255 & ~n1881;
  assign n44228 = ~n221 & ~n894;
  assign n44229 = ~n894 & ~n1881;
  assign n44230 = ~n221 & ~n255;
  assign n44231 = n44229 & n44230;
  assign n44232 = n44227 & n44228;
  assign n44233 = n358 & n3272;
  assign n44234 = n59174 & n44233;
  assign n44235 = n55106 & n44234;
  assign n44236 = n1078 & n3536;
  assign n44237 = n44224 & n44236;
  assign n44238 = n53664 & n44237;
  assign n44239 = n44235 & n44238;
  assign n44240 = n3272 & n17997;
  assign n44241 = n59174 & n44240;
  assign n44242 = n55106 & n44241;
  assign n44243 = n358 & n1078;
  assign n44244 = n3536 & n12008;
  assign n44245 = n44243 & n44244;
  assign n44246 = n53664 & n44245;
  assign n44247 = n44242 & n44246;
  assign n44248 = n44222 & n44226;
  assign n44249 = n54727 & n59175;
  assign n44250 = n56746 & n57073;
  assign n44251 = n44249 & n44250;
  assign n44252 = n3272 & n12008;
  assign n44253 = n55106 & n44252;
  assign n44254 = n54727 & n44253;
  assign n44255 = n57073 & n44254;
  assign n44256 = n56616 & n44255;
  assign n44257 = n56746 & n44256;
  assign n44258 = n1078 & n44257;
  assign n44259 = n358 & n44258;
  assign n44260 = n53664 & n44259;
  assign n44261 = n3536 & n44260;
  assign n44262 = ~n894 & n44261;
  assign n44263 = ~n255 & n44262;
  assign n44264 = ~n221 & n44263;
  assign n44265 = ~n513 & n44264;
  assign n44266 = ~n735 & n44265;
  assign n44267 = ~n1881 & n44266;
  assign n44268 = n56616 & n44251;
  assign n44269 = n58480 & n59176;
  assign n44270 = ~n58480 & ~n59176;
  assign n44271 = ~n44269 & ~n44270;
  assign n44272 = n39778 & n44271;
  assign n44273 = ~n39778 & ~n44271;
  assign n44274 = ~n44272 & ~n44273;
  assign n44275 = ~n39878 & n44274;
  assign n44276 = n39878 & ~n44274;
  assign n44277 = ~n44275 & ~n44276;
  assign n44278 = n1576 & ~n56668;
  assign n44279 = n11215 & n26253;
  assign n44280 = n54403 & n26259;
  assign n44281 = n10564 & n26256;
  assign n44282 = ~n44280 & ~n44281;
  assign n44283 = ~n44279 & n44282;
  assign n44284 = ~n44278 & n44283;
  assign n44285 = n44277 & ~n44284;
  assign n44286 = ~n44277 & n44284;
  assign n44287 = n44277 & ~n44285;
  assign n44288 = ~n44284 & ~n44285;
  assign n44289 = ~n44287 & ~n44288;
  assign n44290 = ~n44285 & ~n44286;
  assign n44291 = n44217 & n59177;
  assign n44292 = ~n44217 & ~n59177;
  assign n44293 = ~n44291 & ~n44292;
  assign n44294 = n11279 & n27839;
  assign n44295 = n12584 & n26244;
  assign n44296 = n54410 & n26250;
  assign n44297 = n11267 & n26247;
  assign n44298 = ~n44296 & ~n44297;
  assign n44299 = ~n44295 & n44298;
  assign n44300 = ~n44294 & n44299;
  assign n44301 = pi29  & ~n44300;
  assign n44302 = pi29  & ~n44301;
  assign n44303 = pi29  & n44300;
  assign n44304 = ~n44300 & ~n44301;
  assign n44305 = ~pi29  & ~n44300;
  assign n44306 = ~n59178 & ~n59179;
  assign n44307 = ~n44293 & n44306;
  assign n44308 = n44293 & ~n44306;
  assign n44309 = n44293 & ~n44308;
  assign n44310 = ~n44306 & ~n44308;
  assign n44311 = ~n44309 & ~n44310;
  assign n44312 = ~n44307 & ~n44308;
  assign n44313 = ~n59173 & ~n59180;
  assign n44314 = n59173 & n59180;
  assign n44315 = ~n59173 & n59180;
  assign n44316 = n59173 & ~n59180;
  assign n44317 = ~n44315 & ~n44316;
  assign n44318 = ~n44313 & ~n44314;
  assign n44319 = ~n39782 & n58488;
  assign n44320 = ~n39782 & ~n39922;
  assign n44321 = ~n39783 & ~n44319;
  assign n44322 = ~n59181 & ~n59182;
  assign n44323 = n59181 & n59182;
  assign n44324 = ~n44322 & ~n44323;
  assign n44325 = ~n44191 & n44324;
  assign n44326 = n44191 & ~n44324;
  assign n44327 = ~n44325 & ~n44326;
  assign n44328 = n39937 & n44327;
  assign n44329 = ~n39937 & ~n44327;
  assign n44330 = ~n44328 & ~n44329;
  assign n44331 = ~n44190 & ~n44329;
  assign n44332 = ~n44328 & n44331;
  assign n44333 = ~n44190 & n44330;
  assign n44334 = n44190 & ~n44330;
  assign n44335 = ~n44190 & ~n59183;
  assign n44336 = ~n44328 & ~n59183;
  assign n44337 = ~n44329 & n44336;
  assign n44338 = ~n44335 & ~n44337;
  assign n44339 = ~n59183 & ~n44334;
  assign n44340 = n77 & ~n59184;
  assign n44341 = n24302 & n44327;
  assign n44342 = n21969 & n39543;
  assign n44343 = n23459 & n39937;
  assign n44344 = ~n44342 & ~n44343;
  assign n44345 = ~n44341 & n44344;
  assign n44346 = ~n44340 & n44345;
  assign n44347 = pi5  & ~n44346;
  assign n44348 = ~n44346 & ~n44347;
  assign n44349 = ~pi5  & ~n44346;
  assign n44350 = pi5  & ~n44347;
  assign n44351 = pi5  & n44346;
  assign n44352 = ~n59185 & ~n59186;
  assign n44353 = ~n43450 & ~n43458;
  assign n44354 = ~n43426 & ~n43433;
  assign n44355 = n18846 & ~n58891;
  assign n44356 = n19541 & n39552;
  assign n44357 = n55247 & n39558;
  assign n44358 = n19509 & n39555;
  assign n44359 = ~n44357 & ~n44358;
  assign n44360 = ~n44356 & n44359;
  assign n44361 = ~n44355 & n44360;
  assign n44362 = pi11  & ~n44361;
  assign n44363 = ~n44361 & ~n44362;
  assign n44364 = ~pi11  & ~n44361;
  assign n44365 = pi11  & ~n44362;
  assign n44366 = pi11  & n44361;
  assign n44367 = ~n59187 & ~n59188;
  assign n44368 = ~n43410 & ~n43418;
  assign n44369 = ~n43386 & ~n43395;
  assign n44370 = n16079 & ~n58759;
  assign n44371 = n16696 & n39570;
  assign n44372 = n54886 & n39576;
  assign n44373 = n16676 & n39573;
  assign n44374 = ~n44372 & ~n44373;
  assign n44375 = ~n44371 & n44374;
  assign n44376 = ~n44370 & n44375;
  assign n44377 = pi17  & ~n44376;
  assign n44378 = ~n44376 & ~n44377;
  assign n44379 = ~pi17  & ~n44376;
  assign n44380 = pi17  & ~n44377;
  assign n44381 = pi17  & n44376;
  assign n44382 = ~n59189 & ~n59190;
  assign n44383 = ~n43372 & ~n43380;
  assign n44384 = ~n43350 & ~n43357;
  assign n44385 = n90 & ~n58585;
  assign n44386 = n14236 & n39588;
  assign n44387 = n54667 & n39594;
  assign n44388 = n14210 & n39591;
  assign n44389 = ~n44387 & ~n44388;
  assign n44390 = ~n44386 & n44389;
  assign n44391 = ~n44385 & n44390;
  assign n44392 = pi23  & ~n44391;
  assign n44393 = ~n44391 & ~n44392;
  assign n44394 = ~pi23  & ~n44391;
  assign n44395 = pi23  & ~n44392;
  assign n44396 = pi23  & n44391;
  assign n44397 = ~n59191 & ~n59192;
  assign n44398 = ~n43334 & ~n43342;
  assign n44399 = ~n43310 & ~n43319;
  assign n44400 = n11279 & n40183;
  assign n44401 = n12584 & n39606;
  assign n44402 = n54410 & n39612;
  assign n44403 = n11267 & n39609;
  assign n44404 = ~n44402 & ~n44403;
  assign n44405 = ~n44401 & n44404;
  assign n44406 = ~n44400 & n44405;
  assign n44407 = pi29  & ~n44406;
  assign n44408 = ~n44406 & ~n44407;
  assign n44409 = ~pi29  & ~n44406;
  assign n44410 = pi29  & ~n44407;
  assign n44411 = pi29  & n44406;
  assign n44412 = ~n59193 & ~n59194;
  assign n44413 = ~n43296 & ~n43304;
  assign n44414 = n3371 & n5445;
  assign n44415 = n54930 & n26696;
  assign n44416 = n44414 & n44415;
  assign n44417 = ~n1127 & ~n1680;
  assign n44418 = ~n1492 & n44417;
  assign n44419 = ~n495 & ~n1059;
  assign n44420 = n27887 & n44419;
  assign n44421 = n44418 & n44420;
  assign n44422 = n56578 & n44421;
  assign n44423 = ~n1059 & ~n1127;
  assign n44424 = ~n495 & ~n1079;
  assign n44425 = n44423 & n44424;
  assign n44426 = n3371 & n44425;
  assign n44427 = n5445 & n54930;
  assign n44428 = n44426 & n44427;
  assign n44429 = ~n733 & ~n1680;
  assign n44430 = n7045 & n44429;
  assign n44431 = n13530 & n44430;
  assign n44432 = n56578 & n44431;
  assign n44433 = n44428 & n44432;
  assign n44434 = ~n495 & ~n1680;
  assign n44435 = ~n1079 & n44434;
  assign n44436 = ~n733 & ~n1059;
  assign n44437 = n7045 & n44436;
  assign n44438 = n44435 & n44437;
  assign n44439 = n3371 & n54930;
  assign n44440 = n44438 & n44439;
  assign n44441 = n1391 & n4893;
  assign n44442 = n13530 & n44441;
  assign n44443 = n56578 & n44442;
  assign n44444 = n44440 & n44443;
  assign n44445 = n44416 & n44422;
  assign n44446 = n56572 & n59195;
  assign n44447 = n58476 & n44446;
  assign n44448 = n7045 & n54930;
  assign n44449 = n13530 & n44448;
  assign n44450 = n4893 & n44449;
  assign n44451 = n3371 & n44450;
  assign n44452 = n58476 & n44451;
  assign n44453 = n56572 & n44452;
  assign n44454 = n56578 & n44453;
  assign n44455 = n57038 & n44454;
  assign n44456 = n1391 & n44455;
  assign n44457 = ~n1079 & n44456;
  assign n44458 = ~n1680 & n44457;
  assign n44459 = ~n1059 & n44458;
  assign n44460 = ~n495 & n44459;
  assign n44461 = ~n733 & n44460;
  assign n44462 = n57038 & n44447;
  assign n44463 = n1576 & n40093;
  assign n44464 = n11215 & n39615;
  assign n44465 = n10564 & n39618;
  assign n44466 = n54403 & n39621;
  assign n44467 = ~n44465 & ~n44466;
  assign n44468 = ~n44464 & n44467;
  assign n44469 = ~n44463 & ~n44466;
  assign n44470 = ~n44465 & n44469;
  assign n44471 = ~n44464 & n44470;
  assign n44472 = ~n44463 & n44468;
  assign n44473 = ~n59196 & ~n59197;
  assign n44474 = n59196 & n59197;
  assign n44475 = ~n59196 & ~n44473;
  assign n44476 = ~n59196 & n59197;
  assign n44477 = ~n59197 & ~n44473;
  assign n44478 = n59196 & ~n59197;
  assign n44479 = ~n59198 & ~n59199;
  assign n44480 = ~n44473 & ~n44474;
  assign n44481 = ~n44413 & ~n59200;
  assign n44482 = n44413 & n59200;
  assign n44483 = ~n44413 & ~n44481;
  assign n44484 = ~n59200 & ~n44481;
  assign n44485 = ~n44483 & ~n44484;
  assign n44486 = ~n44481 & ~n44482;
  assign n44487 = ~n44412 & ~n59201;
  assign n44488 = n44412 & n59201;
  assign n44489 = ~n44412 & ~n44487;
  assign n44490 = ~n44412 & n59201;
  assign n44491 = ~n59201 & ~n44487;
  assign n44492 = n44412 & ~n59201;
  assign n44493 = ~n59202 & ~n59203;
  assign n44494 = ~n44487 & ~n44488;
  assign n44495 = n44399 & n59204;
  assign n44496 = ~n44399 & ~n59204;
  assign n44497 = ~n44495 & ~n44496;
  assign n44498 = n123 & n40247;
  assign n44499 = n128 & n39597;
  assign n44500 = n53444 & n39603;
  assign n44501 = n127 & n39600;
  assign n44502 = ~n44500 & ~n44501;
  assign n44503 = ~n44499 & n44502;
  assign n44504 = ~n123 & n44503;
  assign n44505 = ~n40247 & n44503;
  assign n44506 = ~n44504 & ~n44505;
  assign n44507 = ~n44498 & n44503;
  assign n44508 = pi26  & ~n59205;
  assign n44509 = ~pi26  & n59205;
  assign n44510 = ~n44508 & ~n44509;
  assign n44511 = n44497 & ~n44510;
  assign n44512 = ~n44497 & n44510;
  assign n44513 = n44497 & ~n44511;
  assign n44514 = n44497 & n44510;
  assign n44515 = ~n44510 & ~n44511;
  assign n44516 = ~n44497 & ~n44510;
  assign n44517 = ~n59206 & ~n59207;
  assign n44518 = ~n44511 & ~n44512;
  assign n44519 = ~n44398 & ~n59208;
  assign n44520 = n44398 & n59208;
  assign n44521 = ~n44398 & ~n44519;
  assign n44522 = ~n44398 & n59208;
  assign n44523 = ~n59208 & ~n44519;
  assign n44524 = n44398 & ~n59208;
  assign n44525 = ~n59209 & ~n59210;
  assign n44526 = ~n44519 & ~n44520;
  assign n44527 = ~n44397 & ~n59211;
  assign n44528 = n44397 & n59211;
  assign n44529 = ~n44397 & ~n44527;
  assign n44530 = ~n59211 & ~n44527;
  assign n44531 = ~n44529 & ~n44530;
  assign n44532 = ~n44527 & ~n44528;
  assign n44533 = n44384 & n59212;
  assign n44534 = ~n44384 & ~n59212;
  assign n44535 = ~n44533 & ~n44534;
  assign n44536 = n14413 & ~n58657;
  assign n44537 = n15921 & n39579;
  assign n44538 = n54719 & n39585;
  assign n44539 = n15901 & n39582;
  assign n44540 = ~n44538 & ~n44539;
  assign n44541 = ~n44537 & n44540;
  assign n44542 = ~n14413 & n44541;
  assign n44543 = n58657 & n44541;
  assign n44544 = ~n44542 & ~n44543;
  assign n44545 = ~n44536 & n44541;
  assign n44546 = pi20  & ~n59213;
  assign n44547 = ~pi20  & n59213;
  assign n44548 = ~n44546 & ~n44547;
  assign n44549 = n44535 & ~n44548;
  assign n44550 = ~n44535 & n44548;
  assign n44551 = n44535 & ~n44549;
  assign n44552 = n44535 & n44548;
  assign n44553 = ~n44548 & ~n44549;
  assign n44554 = ~n44535 & ~n44548;
  assign n44555 = ~n59214 & ~n59215;
  assign n44556 = ~n44549 & ~n44550;
  assign n44557 = ~n44383 & ~n59216;
  assign n44558 = n44383 & n59216;
  assign n44559 = ~n44383 & ~n44557;
  assign n44560 = ~n59216 & ~n44557;
  assign n44561 = ~n44559 & ~n44560;
  assign n44562 = ~n44557 & ~n44558;
  assign n44563 = ~n44382 & ~n59217;
  assign n44564 = n44382 & n59217;
  assign n44565 = ~n44382 & ~n44563;
  assign n44566 = ~n44382 & n59217;
  assign n44567 = ~n59217 & ~n44563;
  assign n44568 = n44382 & ~n59217;
  assign n44569 = ~n59218 & ~n59219;
  assign n44570 = ~n44563 & ~n44564;
  assign n44571 = n44369 & n59220;
  assign n44572 = ~n44369 & ~n59220;
  assign n44573 = ~n44571 & ~n44572;
  assign n44574 = n17265 & ~n58493;
  assign n44575 = n18588 & n39561;
  assign n44576 = n55041 & n39567;
  assign n44577 = n18556 & n39564;
  assign n44578 = ~n44576 & ~n44577;
  assign n44579 = ~n44575 & n44578;
  assign n44580 = ~n17265 & n44579;
  assign n44581 = n58493 & n44579;
  assign n44582 = ~n44580 & ~n44581;
  assign n44583 = ~n44574 & n44579;
  assign n44584 = pi14  & ~n59221;
  assign n44585 = ~pi14  & n59221;
  assign n44586 = ~n44584 & ~n44585;
  assign n44587 = n44573 & ~n44586;
  assign n44588 = ~n44573 & n44586;
  assign n44589 = n44573 & ~n44587;
  assign n44590 = n44573 & n44586;
  assign n44591 = ~n44586 & ~n44587;
  assign n44592 = ~n44573 & ~n44586;
  assign n44593 = ~n59222 & ~n59223;
  assign n44594 = ~n44587 & ~n44588;
  assign n44595 = ~n44368 & ~n59224;
  assign n44596 = n44368 & n59224;
  assign n44597 = ~n44368 & ~n44595;
  assign n44598 = ~n44368 & n59224;
  assign n44599 = ~n59224 & ~n44595;
  assign n44600 = n44368 & ~n59224;
  assign n44601 = ~n59225 & ~n59226;
  assign n44602 = ~n44595 & ~n44596;
  assign n44603 = ~n44367 & ~n59227;
  assign n44604 = n44367 & n59227;
  assign n44605 = ~n44367 & ~n44603;
  assign n44606 = ~n59227 & ~n44603;
  assign n44607 = ~n44605 & ~n44606;
  assign n44608 = ~n44603 & ~n44604;
  assign n44609 = n44354 & n59228;
  assign n44610 = ~n44354 & ~n59228;
  assign n44611 = ~n44609 & ~n44610;
  assign n44612 = n20085 & ~n59050;
  assign n44613 = n21269 & n39440;
  assign n44614 = n55472 & n39549;
  assign n44615 = n21237 & n39546;
  assign n44616 = ~n44614 & ~n44615;
  assign n44617 = ~n44613 & n44616;
  assign n44618 = ~n20085 & n44617;
  assign n44619 = n59050 & n44617;
  assign n44620 = ~n44618 & ~n44619;
  assign n44621 = ~n44612 & n44617;
  assign n44622 = pi8  & ~n59229;
  assign n44623 = ~pi8  & n59229;
  assign n44624 = ~n44622 & ~n44623;
  assign n44625 = n44611 & ~n44624;
  assign n44626 = ~n44611 & n44624;
  assign n44627 = n44611 & ~n44625;
  assign n44628 = n44611 & n44624;
  assign n44629 = ~n44624 & ~n44625;
  assign n44630 = ~n44611 & ~n44624;
  assign n44631 = ~n59230 & ~n59231;
  assign n44632 = ~n44625 & ~n44626;
  assign n44633 = ~n44353 & ~n59232;
  assign n44634 = n44353 & n59232;
  assign n44635 = ~n44353 & ~n44633;
  assign n44636 = ~n59232 & ~n44633;
  assign n44637 = ~n44635 & ~n44636;
  assign n44638 = ~n44633 & ~n44634;
  assign n44639 = ~n44352 & ~n59233;
  assign n44640 = n44352 & n59233;
  assign n44641 = ~n44352 & ~n44639;
  assign n44642 = ~n44352 & n59233;
  assign n44643 = ~n59233 & ~n44639;
  assign n44644 = n44352 & ~n59233;
  assign n44645 = ~n59234 & ~n59235;
  assign n44646 = ~n44639 & ~n44640;
  assign n44647 = n44189 & n59236;
  assign n44648 = ~n44189 & ~n59236;
  assign n44649 = ~n44647 & ~n44648;
  assign n44650 = ~n44322 & ~n44325;
  assign n44651 = ~n44209 & ~n44313;
  assign n44652 = n53444 & ~n26537;
  assign n44653 = ~n127 & ~n44652;
  assign n44654 = ~n128 & n44653;
  assign n44655 = ~n128 & ~n44652;
  assign n44656 = ~n127 & n44655;
  assign n44657 = n129 & ~n44652;
  assign n44658 = ~n123 & n59237;
  assign n44659 = pi26  & ~n44658;
  assign n44660 = pi26  & ~n44659;
  assign n44661 = pi26  & n44658;
  assign n44662 = ~n44658 & ~n44659;
  assign n44663 = ~pi26  & ~n44658;
  assign n44664 = ~n59238 & ~n59239;
  assign n44665 = ~n44270 & ~n44272;
  assign n44666 = ~n510 & ~n1658;
  assign n44667 = ~n510 & ~n649;
  assign n44668 = ~n659 & ~n1658;
  assign n44669 = n44667 & n44668;
  assign n44670 = ~n510 & ~n659;
  assign n44671 = ~n649 & ~n1658;
  assign n44672 = n44670 & n44671;
  assign n44673 = n2503 & n44666;
  assign n44674 = n1078 & n59240;
  assign n44675 = n1279 & n55148;
  assign n44676 = n1078 & n55148;
  assign n44677 = n1277 & n44676;
  assign n44678 = n1278 & n44677;
  assign n44679 = ~n659 & n44678;
  assign n44680 = ~n1658 & n44679;
  assign n44681 = ~n510 & n44680;
  assign n44682 = ~n649 & n44681;
  assign n44683 = n1078 & n1277;
  assign n44684 = n1278 & n44683;
  assign n44685 = n55148 & n59240;
  assign n44686 = n44684 & n44685;
  assign n44687 = n44674 & n44675;
  assign n44688 = n462 & ~n1085;
  assign n44689 = n3671 & n3716;
  assign n44690 = n6152 & n8793;
  assign n44691 = n44689 & n44690;
  assign n44692 = ~n662 & ~n1085;
  assign n44693 = ~n1085 & n6152;
  assign n44694 = ~n1457 & n44692;
  assign n44695 = n462 & n3716;
  assign n44696 = n3671 & n8793;
  assign n44697 = n44695 & n44696;
  assign n44698 = n59242 & n44697;
  assign n44699 = n44688 & n44691;
  assign n44700 = n53684 & n59243;
  assign n44701 = n59241 & n44700;
  assign n44702 = n53479 & n44701;
  assign n44703 = n53479 & n3716;
  assign n44704 = n53700 & n44703;
  assign n44705 = n53684 & n44704;
  assign n44706 = n53693 & n44705;
  assign n44707 = n3671 & n44706;
  assign n44708 = n59241 & n44707;
  assign n44709 = n8793 & n44708;
  assign n44710 = n462 & n44709;
  assign n44711 = ~n1085 & n44710;
  assign n44712 = ~n662 & n44711;
  assign n44713 = ~n1457 & n44712;
  assign n44714 = n3060 & n44702;
  assign n44715 = ~n44665 & n59244;
  assign n44716 = n44665 & ~n59244;
  assign n44717 = ~n44715 & ~n44716;
  assign n44718 = n1576 & n27491;
  assign n44719 = n11215 & n26250;
  assign n44720 = n10564 & n26253;
  assign n44721 = n54403 & n26256;
  assign n44722 = ~n44720 & ~n44721;
  assign n44723 = ~n44719 & n44722;
  assign n44724 = ~n44718 & ~n44721;
  assign n44725 = ~n44720 & n44724;
  assign n44726 = ~n44719 & n44725;
  assign n44727 = ~n44718 & n44723;
  assign n44728 = n44717 & ~n59245;
  assign n44729 = ~n44717 & n59245;
  assign n44730 = ~n44728 & ~n44729;
  assign n44731 = ~n44275 & n44284;
  assign n44732 = ~n44275 & ~n44285;
  assign n44733 = ~n44276 & ~n44731;
  assign n44734 = n44730 & ~n59246;
  assign n44735 = ~n44730 & n59246;
  assign n44736 = ~n44734 & ~n44735;
  assign n44737 = n11279 & n27808;
  assign n44738 = n12584 & n26242;
  assign n44739 = n54410 & n26247;
  assign n44740 = n11267 & n26244;
  assign n44741 = ~n44739 & ~n44740;
  assign n44742 = ~n44738 & n44741;
  assign n44743 = ~n11279 & n44742;
  assign n44744 = ~n27808 & n44742;
  assign n44745 = ~n44743 & ~n44744;
  assign n44746 = ~n44737 & n44742;
  assign n44747 = pi29  & ~n59247;
  assign n44748 = ~pi29  & n59247;
  assign n44749 = ~n44747 & ~n44748;
  assign n44750 = n44736 & ~n44749;
  assign n44751 = ~n44736 & n44749;
  assign n44752 = ~n44750 & ~n44751;
  assign n44753 = ~n44292 & n44306;
  assign n44754 = ~n44292 & ~n44308;
  assign n44755 = ~n44291 & ~n44753;
  assign n44756 = ~n44752 & n59248;
  assign n44757 = n44752 & ~n59248;
  assign n44758 = ~n44756 & ~n44757;
  assign n44759 = n44664 & ~n44758;
  assign n44760 = ~n44664 & n44758;
  assign n44761 = n44758 & ~n44760;
  assign n44762 = n44664 & n44758;
  assign n44763 = ~n44664 & ~n44760;
  assign n44764 = ~n44664 & ~n44758;
  assign n44765 = ~n59249 & ~n59250;
  assign n44766 = ~n44759 & ~n44760;
  assign n44767 = ~n44651 & ~n59251;
  assign n44768 = n44651 & n59251;
  assign n44769 = ~n59251 & ~n44767;
  assign n44770 = ~n44651 & ~n44767;
  assign n44771 = ~n44769 & ~n44770;
  assign n44772 = ~n44767 & ~n44768;
  assign n44773 = ~n44650 & ~n59252;
  assign n44774 = n44650 & n59252;
  assign n44775 = ~n44773 & ~n44774;
  assign n44776 = ~n44767 & ~n44773;
  assign n44777 = ~n44715 & ~n44728;
  assign n44778 = ~n1044 & ~n1457;
  assign n44779 = n494 & n44778;
  assign n44780 = n2538 & n16350;
  assign n44781 = n2538 & n44778;
  assign n44782 = n494 & n16350;
  assign n44783 = n44781 & n44782;
  assign n44784 = n16350 & n44778;
  assign n44785 = n494 & n2538;
  assign n44786 = n44784 & n44785;
  assign n44787 = n44779 & n44780;
  assign n44788 = n53825 & n5690;
  assign n44789 = n59253 & n44788;
  assign n44790 = n53542 & n44789;
  assign n44791 = n53649 & n44790;
  assign n44792 = n53479 & n44791;
  assign n44793 = n53649 & n44788;
  assign n44794 = n53677 & n44793;
  assign n44795 = n53479 & n44794;
  assign n44796 = n53542 & n44795;
  assign n44797 = n494 & n44796;
  assign n44798 = n53668 & n44797;
  assign n44799 = ~n1044 & n44798;
  assign n44800 = ~n1457 & n44799;
  assign n44801 = ~n514 & n44800;
  assign n44802 = ~n852 & n44801;
  assign n44803 = ~n1646 & n44802;
  assign n44804 = ~n1634 & n44803;
  assign n44805 = n53677 & n44792;
  assign n44806 = n53668 & n44805;
  assign n44807 = n2875 & n44792;
  assign n44808 = ~n59244 & n59254;
  assign n44809 = n59244 & ~n59254;
  assign n44810 = ~n44808 & ~n44809;
  assign n44811 = n1576 & ~n56567;
  assign n44812 = n11215 & n26247;
  assign n44813 = n54403 & n26253;
  assign n44814 = n10564 & n26250;
  assign n44815 = ~n44813 & ~n44814;
  assign n44816 = ~n44812 & n44815;
  assign n44817 = ~n44811 & n44816;
  assign n44818 = ~n44809 & ~n44817;
  assign n44819 = ~n44808 & n44818;
  assign n44820 = n44810 & ~n44817;
  assign n44821 = ~n44810 & n44817;
  assign n44822 = ~n44817 & ~n59255;
  assign n44823 = ~n44809 & ~n59255;
  assign n44824 = ~n44808 & n44823;
  assign n44825 = ~n44822 & ~n44824;
  assign n44826 = ~n59255 & ~n44821;
  assign n44827 = n44777 & n59256;
  assign n44828 = ~n44777 & ~n59256;
  assign n44829 = ~n44827 & ~n44828;
  assign n44830 = ~n44734 & ~n44750;
  assign n44831 = ~n44829 & n44830;
  assign n44832 = n44829 & ~n44830;
  assign n44833 = ~n44831 & ~n44832;
  assign n44834 = ~n53445 & ~n135;
  assign n44835 = ~pi26  & ~n53445;
  assign n44836 = ~n53446 & ~n59257;
  assign n44837 = n11279 & ~n56564;
  assign n44838 = n12584 & ~n26537;
  assign n44839 = n54410 & n26244;
  assign n44840 = n11267 & n26242;
  assign n44841 = ~n44839 & ~n44840;
  assign n44842 = ~n44838 & n44841;
  assign n44843 = ~n44837 & n44842;
  assign n44844 = pi29  & ~n44843;
  assign n44845 = pi29  & ~n44844;
  assign n44846 = pi29  & n44843;
  assign n44847 = ~n44843 & ~n44844;
  assign n44848 = ~pi29  & ~n44843;
  assign n44849 = ~n59258 & ~n59259;
  assign n44850 = ~n44836 & ~n44849;
  assign n44851 = n44836 & n44849;
  assign n44852 = ~n44836 & ~n44850;
  assign n44853 = ~n44836 & n44849;
  assign n44854 = ~n44849 & ~n44850;
  assign n44855 = n44836 & ~n44849;
  assign n44856 = ~n59260 & ~n59261;
  assign n44857 = ~n44850 & ~n44851;
  assign n44858 = ~n44833 & n59262;
  assign n44859 = n44833 & ~n59262;
  assign n44860 = ~n44858 & ~n44859;
  assign n44861 = n44664 & ~n44757;
  assign n44862 = ~n44664 & ~n44756;
  assign n44863 = ~n44757 & ~n44862;
  assign n44864 = ~n44757 & ~n44760;
  assign n44865 = ~n44756 & ~n44861;
  assign n44866 = n44860 & ~n59263;
  assign n44867 = ~n44860 & n59263;
  assign n44868 = ~n44866 & ~n44867;
  assign n44869 = ~n44776 & n44868;
  assign n44870 = n44776 & ~n44868;
  assign n44871 = ~n44869 & ~n44870;
  assign n44872 = n44775 & n44871;
  assign n44873 = n44327 & n44775;
  assign n44874 = ~n44327 & ~n44775;
  assign n44875 = ~n44873 & ~n44874;
  assign n44876 = ~n44336 & ~n44874;
  assign n44877 = ~n44873 & n44876;
  assign n44878 = ~n44336 & n44875;
  assign n44879 = ~n44873 & ~n59264;
  assign n44880 = ~n44775 & ~n44871;
  assign n44881 = ~n44872 & ~n44880;
  assign n44882 = ~n44879 & ~n44880;
  assign n44883 = ~n44872 & n44882;
  assign n44884 = ~n44879 & n44881;
  assign n44885 = ~n44872 & ~n59265;
  assign n44886 = ~n44866 & ~n44869;
  assign n44887 = ~n44828 & ~n44832;
  assign n44888 = n11279 & n28624;
  assign n44889 = n54410 & n26242;
  assign n44890 = ~n11267 & ~n44889;
  assign n44891 = ~n12584 & ~n44889;
  assign n44892 = ~n11267 & n44891;
  assign n44893 = ~n12584 & n44890;
  assign n44894 = ~n44888 & n59266;
  assign n44895 = pi29  & ~n44894;
  assign n44896 = pi29  & ~n44895;
  assign n44897 = pi29  & n44894;
  assign n44898 = ~n44894 & ~n44895;
  assign n44899 = ~pi29  & ~n44894;
  assign n44900 = ~n59267 & ~n59268;
  assign n44901 = n53564 & n53633;
  assign n44902 = ~n1457 & n44901;
  assign n44903 = n1627 & n53633;
  assign n44904 = ~n852 & ~n1081;
  assign n44905 = n1197 & n44904;
  assign n44906 = n53646 & n44905;
  assign n44907 = n53463 & n44906;
  assign n44908 = n53463 & n53646;
  assign n44909 = n1197 & n44908;
  assign n44910 = n59269 & n44909;
  assign n44911 = ~n1081 & n44910;
  assign n44912 = ~n852 & n44911;
  assign n44913 = n59269 & n44907;
  assign n44914 = n59244 & n59270;
  assign n44915 = ~n59244 & ~n59270;
  assign n44916 = ~n44914 & ~n44915;
  assign n44917 = n44836 & n44916;
  assign n44918 = ~n44836 & ~n44916;
  assign n44919 = ~n44917 & ~n44918;
  assign n44920 = ~n44823 & n44919;
  assign n44921 = n44823 & ~n44919;
  assign n44922 = ~n44920 & ~n44921;
  assign n44923 = n1576 & n27839;
  assign n44924 = n11215 & n26244;
  assign n44925 = n54403 & n26247;
  assign n44926 = n54403 & n26250;
  assign n44927 = n10564 & n26247;
  assign n44928 = ~n59271 & ~n44927;
  assign n44929 = ~n44924 & n44928;
  assign n44930 = ~n44923 & n44929;
  assign n44931 = n44922 & ~n44930;
  assign n44932 = ~n44922 & n44930;
  assign n44933 = n44922 & ~n44931;
  assign n44934 = ~n44930 & ~n44931;
  assign n44935 = ~n44933 & ~n44934;
  assign n44936 = ~n44931 & ~n44932;
  assign n44937 = ~n44900 & ~n59272;
  assign n44938 = n44900 & n59272;
  assign n44939 = ~n59272 & ~n44937;
  assign n44940 = ~n44900 & ~n44937;
  assign n44941 = ~n44939 & ~n44940;
  assign n44942 = ~n44937 & ~n44938;
  assign n44943 = n44887 & n59273;
  assign n44944 = ~n44887 & ~n59273;
  assign n44945 = ~n44943 & ~n44944;
  assign n44946 = ~n44850 & ~n44859;
  assign n44947 = n44945 & ~n44946;
  assign n44948 = ~n44945 & n44946;
  assign n44949 = ~n44947 & ~n44948;
  assign n44950 = n44886 & ~n44949;
  assign n44951 = ~n44886 & n44949;
  assign n44952 = ~n44950 & ~n44951;
  assign n44953 = n44871 & n44952;
  assign n44954 = ~n44871 & ~n44952;
  assign n44955 = ~n44953 & ~n44954;
  assign n44956 = ~n44885 & ~n44954;
  assign n44957 = ~n44953 & n44956;
  assign n44958 = ~n44885 & n44955;
  assign n44959 = n44885 & ~n44955;
  assign n44960 = ~n44885 & ~n59274;
  assign n44961 = ~n44953 & ~n59274;
  assign n44962 = ~n44954 & n44961;
  assign n44963 = ~n44960 & ~n44962;
  assign n44964 = ~n59274 & ~n44959;
  assign n44965 = n24338 & ~n59275;
  assign n44966 = n25287 & n44952;
  assign n44967 = n24337 & n44775;
  assign n44968 = n25272 & n44871;
  assign n44969 = ~n44967 & ~n44968;
  assign n44970 = ~n44966 & n44969;
  assign n44971 = ~n24338 & n44970;
  assign n44972 = n59275 & n44970;
  assign n44973 = ~n44971 & ~n44972;
  assign n44974 = ~n44965 & n44970;
  assign n44975 = pi2  & ~n59276;
  assign n44976 = ~pi2  & n59276;
  assign n44977 = ~n44975 & ~n44976;
  assign n44978 = n44649 & ~n44977;
  assign n44979 = ~n44649 & n44977;
  assign n44980 = n44649 & ~n44978;
  assign n44981 = n44649 & n44977;
  assign n44982 = ~n44977 & ~n44978;
  assign n44983 = ~n44649 & ~n44977;
  assign n44984 = ~n59277 & ~n59278;
  assign n44985 = ~n44978 & ~n44979;
  assign n44986 = n44879 & ~n44881;
  assign n44987 = ~n44879 & ~n59265;
  assign n44988 = ~n44880 & n44885;
  assign n44989 = ~n44987 & ~n44988;
  assign n44990 = ~n59265 & ~n44986;
  assign n44991 = n24338 & ~n59280;
  assign n44992 = n25287 & n44871;
  assign n44993 = n24337 & n44327;
  assign n44994 = n25272 & n44775;
  assign n44995 = ~n44993 & ~n44994;
  assign n44996 = ~n44992 & n44995;
  assign n44997 = ~n24338 & n44996;
  assign n44998 = n59280 & n44996;
  assign n44999 = ~n44997 & ~n44998;
  assign n45000 = ~n44991 & n44996;
  assign n45001 = pi2  & ~n59281;
  assign n45002 = ~pi2  & n59281;
  assign n45003 = ~n45001 & ~n45002;
  assign n45004 = n44336 & ~n44875;
  assign n45005 = ~n44336 & ~n59264;
  assign n45006 = ~n44874 & n44879;
  assign n45007 = ~n45005 & ~n45006;
  assign n45008 = ~n59264 & ~n45004;
  assign n45009 = n24338 & ~n59282;
  assign n45010 = n25287 & n44775;
  assign n45011 = n24337 & n39937;
  assign n45012 = n25272 & n44327;
  assign n45013 = ~n45011 & ~n45012;
  assign n45014 = ~n45010 & n45013;
  assign n45015 = ~n24338 & n45014;
  assign n45016 = n59282 & n45014;
  assign n45017 = ~n45015 & ~n45016;
  assign n45018 = ~n45009 & n45014;
  assign n45019 = pi2  & ~n59283;
  assign n45020 = ~pi2  & n59283;
  assign n45021 = ~n45019 & ~n45020;
  assign n45022 = n24338 & ~n59184;
  assign n45023 = n25287 & n44327;
  assign n45024 = n24337 & n39543;
  assign n45025 = n25272 & n39937;
  assign n45026 = ~n45024 & ~n45025;
  assign n45027 = ~n45023 & n45026;
  assign n45028 = ~n24338 & n45027;
  assign n45029 = n59184 & n45027;
  assign n45030 = ~n45028 & ~n45029;
  assign n45031 = ~n45022 & n45027;
  assign n45032 = pi2  & ~n59284;
  assign n45033 = ~pi2  & n59284;
  assign n45034 = ~n45032 & ~n45033;
  assign n45035 = n44162 & ~n44164;
  assign n45036 = ~n44165 & ~n45035;
  assign n45037 = n44153 & ~n59160;
  assign n45038 = ~n59159 & n45037;
  assign n45039 = n44153 & n59161;
  assign n45040 = ~n44161 & ~n59285;
  assign n45041 = n24338 & ~n59050;
  assign n45042 = n25287 & n39440;
  assign n45043 = n24337 & n39549;
  assign n45044 = n25272 & n39546;
  assign n45045 = ~n45043 & ~n45044;
  assign n45046 = ~n45042 & n45045;
  assign n45047 = ~n24338 & n45046;
  assign n45048 = n59050 & n45046;
  assign n45049 = ~n45047 & ~n45048;
  assign n45050 = ~n45041 & n45046;
  assign n45051 = pi2  & ~n59286;
  assign n45052 = ~pi2  & n59286;
  assign n45053 = ~n45051 & ~n45052;
  assign n45054 = n24338 & n43436;
  assign n45055 = n25287 & n39546;
  assign n45056 = n24337 & n39552;
  assign n45057 = n25272 & n39549;
  assign n45058 = ~n45056 & ~n45057;
  assign n45059 = ~n45055 & n45058;
  assign n45060 = ~n24338 & n45059;
  assign n45061 = ~n43436 & n45059;
  assign n45062 = ~n45060 & ~n45061;
  assign n45063 = ~n45054 & n45059;
  assign n45064 = pi2  & ~n59287;
  assign n45065 = ~pi2  & n59287;
  assign n45066 = ~n45064 & ~n45065;
  assign n45067 = n24338 & ~n58889;
  assign n45068 = n25287 & n39549;
  assign n45069 = n24337 & n39555;
  assign n45070 = n25272 & n39552;
  assign n45071 = ~n45069 & ~n45070;
  assign n45072 = ~n45068 & n45071;
  assign n45073 = ~n24338 & n45072;
  assign n45074 = n58889 & n45072;
  assign n45075 = ~n45073 & ~n45074;
  assign n45076 = ~n45067 & n45072;
  assign n45077 = pi2  & ~n59288;
  assign n45078 = ~pi2  & n59288;
  assign n45079 = ~n45077 & ~n45078;
  assign n45080 = n44124 & ~n44126;
  assign n45081 = ~n44127 & ~n45080;
  assign n45082 = n44115 & ~n59150;
  assign n45083 = ~n59149 & n45082;
  assign n45084 = n44115 & n59151;
  assign n45085 = ~n44123 & ~n59289;
  assign n45086 = n44106 & ~n59147;
  assign n45087 = ~n59146 & n45086;
  assign n45088 = n44106 & n59148;
  assign n45089 = ~n44114 & ~n59290;
  assign n45090 = n24338 & ~n58493;
  assign n45091 = n25287 & n39561;
  assign n45092 = n24337 & n39567;
  assign n45093 = n25272 & n39564;
  assign n45094 = ~n45092 & ~n45093;
  assign n45095 = ~n45091 & n45094;
  assign n45096 = ~n24338 & n45095;
  assign n45097 = n58493 & n45095;
  assign n45098 = ~n45096 & ~n45097;
  assign n45099 = ~n45090 & n45095;
  assign n45100 = pi2  & ~n59291;
  assign n45101 = ~pi2  & n59291;
  assign n45102 = ~n45100 & ~n45101;
  assign n45103 = n24338 & n41762;
  assign n45104 = n25287 & n39564;
  assign n45105 = n24337 & n39570;
  assign n45106 = n25272 & n39567;
  assign n45107 = ~n45105 & ~n45106;
  assign n45108 = ~n45104 & n45107;
  assign n45109 = ~n24338 & n45108;
  assign n45110 = ~n41762 & n45108;
  assign n45111 = ~n45109 & ~n45110;
  assign n45112 = ~n45103 & n45108;
  assign n45113 = pi2  & ~n59292;
  assign n45114 = ~pi2  & n59292;
  assign n45115 = ~n45113 & ~n45114;
  assign n45116 = n24338 & ~n58766;
  assign n45117 = n25287 & n39567;
  assign n45118 = n24337 & n39573;
  assign n45119 = n25272 & n39570;
  assign n45120 = ~n45118 & ~n45119;
  assign n45121 = ~n45117 & n45120;
  assign n45122 = ~n24338 & n45121;
  assign n45123 = n58766 & n45121;
  assign n45124 = ~n45122 & ~n45123;
  assign n45125 = ~n45116 & n45121;
  assign n45126 = pi2  & ~n59293;
  assign n45127 = ~pi2  & n59293;
  assign n45128 = ~n45126 & ~n45127;
  assign n45129 = n44077 & ~n44079;
  assign n45130 = ~n44080 & ~n45129;
  assign n45131 = n44068 & ~n59137;
  assign n45132 = ~n59136 & n45131;
  assign n45133 = n44068 & n59138;
  assign n45134 = ~n44076 & ~n59294;
  assign n45135 = n44059 & ~n59134;
  assign n45136 = ~n59133 & n45135;
  assign n45137 = n44059 & n59135;
  assign n45138 = ~n44067 & ~n59295;
  assign n45139 = n24338 & ~n58657;
  assign n45140 = n25287 & n39579;
  assign n45141 = n24337 & n39585;
  assign n45142 = n25272 & n39582;
  assign n45143 = ~n45141 & ~n45142;
  assign n45144 = ~n45140 & n45143;
  assign n45145 = ~n24338 & n45144;
  assign n45146 = n58657 & n45144;
  assign n45147 = ~n45145 & ~n45146;
  assign n45148 = ~n45139 & n45144;
  assign n45149 = pi2  & ~n59296;
  assign n45150 = ~pi2  & n59296;
  assign n45151 = ~n45149 & ~n45150;
  assign n45152 = n24338 & n41007;
  assign n45153 = n25287 & n39582;
  assign n45154 = n24337 & n39588;
  assign n45155 = n25272 & n39585;
  assign n45156 = ~n45154 & ~n45155;
  assign n45157 = ~n45153 & n45156;
  assign n45158 = ~n24338 & n45157;
  assign n45159 = ~n41007 & n45157;
  assign n45160 = ~n45158 & ~n45159;
  assign n45161 = ~n45152 & n45157;
  assign n45162 = pi2  & ~n59297;
  assign n45163 = ~pi2  & n59297;
  assign n45164 = ~n45162 & ~n45163;
  assign n45165 = n24338 & ~n58583;
  assign n45166 = n25287 & n39585;
  assign n45167 = n24337 & n39591;
  assign n45168 = n25272 & n39588;
  assign n45169 = ~n45167 & ~n45168;
  assign n45170 = ~n45166 & n45169;
  assign n45171 = ~n24338 & n45170;
  assign n45172 = n58583 & n45170;
  assign n45173 = ~n45171 & ~n45172;
  assign n45174 = ~n45165 & n45170;
  assign n45175 = pi2  & ~n59298;
  assign n45176 = ~pi2  & n59298;
  assign n45177 = ~n45175 & ~n45176;
  assign n45178 = n44030 & ~n44032;
  assign n45179 = ~n44033 & ~n45178;
  assign n45180 = n44021 & ~n59124;
  assign n45181 = ~n59123 & n45180;
  assign n45182 = n44021 & ~n59123;
  assign n45183 = ~n59124 & n45182;
  assign n45184 = n44021 & n59125;
  assign n45185 = ~n44029 & ~n59299;
  assign n45186 = n44012 & ~n59121;
  assign n45187 = ~n59120 & n45186;
  assign n45188 = n44012 & n59122;
  assign n45189 = ~n44020 & ~n59300;
  assign n45190 = n24338 & n40247;
  assign n45191 = n25287 & n39597;
  assign n45192 = n24337 & n39603;
  assign n45193 = n25272 & n39600;
  assign n45194 = ~n45192 & ~n45193;
  assign n45195 = ~n45191 & n45194;
  assign n45196 = ~n24338 & n45195;
  assign n45197 = ~n40247 & n45195;
  assign n45198 = ~n45196 & ~n45197;
  assign n45199 = ~n45190 & n45195;
  assign n45200 = pi2  & ~n59301;
  assign n45201 = ~pi2  & n59301;
  assign n45202 = ~n45200 & ~n45201;
  assign n45203 = n24338 & ~n58533;
  assign n45204 = n25287 & n39600;
  assign n45205 = n24337 & n39606;
  assign n45206 = n25272 & n39603;
  assign n45207 = ~n45205 & ~n45206;
  assign n45208 = ~n45204 & n45207;
  assign n45209 = ~n24338 & n45208;
  assign n45210 = n58533 & n45208;
  assign n45211 = ~n45209 & ~n45210;
  assign n45212 = ~n45203 & n45208;
  assign n45213 = pi2  & ~n59302;
  assign n45214 = ~pi2  & n59302;
  assign n45215 = ~n45213 & ~n45214;
  assign n45216 = n24338 & n40286;
  assign n45217 = n25287 & n39603;
  assign n45218 = n24337 & n39609;
  assign n45219 = n25272 & n39606;
  assign n45220 = ~n45218 & ~n45219;
  assign n45221 = ~n45217 & n45220;
  assign n45222 = ~n24338 & n45221;
  assign n45223 = ~n40286 & n45221;
  assign n45224 = ~n45222 & ~n45223;
  assign n45225 = ~n45216 & n45221;
  assign n45226 = pi2  & ~n59303;
  assign n45227 = ~pi2  & n59303;
  assign n45228 = ~n45226 & ~n45227;
  assign n45229 = n43986 & ~n43988;
  assign n45230 = ~n43989 & ~n45229;
  assign n45231 = n24338 & n39991;
  assign n45232 = n25287 & n39609;
  assign n45233 = n24337 & n39615;
  assign n45234 = n25272 & n39612;
  assign n45235 = ~n45233 & ~n45234;
  assign n45236 = ~n45232 & n45235;
  assign n45237 = ~n24338 & n45236;
  assign n45238 = ~n39991 & n45236;
  assign n45239 = ~n45237 & ~n45238;
  assign n45240 = ~n45231 & n45236;
  assign n45241 = pi2  & ~n59304;
  assign n45242 = ~pi2  & n59304;
  assign n45243 = ~n45241 & ~n45242;
  assign n45244 = pi5  & ~n59106;
  assign n45245 = ~n59107 & ~n45244;
  assign n45246 = n59107 & n45244;
  assign n45247 = ~n59106 & n43961;
  assign n45248 = ~n59108 & ~n45247;
  assign n45249 = ~n45245 & ~n45246;
  assign n45250 = n24338 & n40093;
  assign n45251 = n25287 & n39615;
  assign n45252 = n24337 & n39621;
  assign n45253 = n25272 & n39618;
  assign n45254 = ~n45252 & ~n45253;
  assign n45255 = ~n45251 & n45254;
  assign n45256 = ~n24338 & n45255;
  assign n45257 = ~n40093 & n45255;
  assign n45258 = ~n45256 & ~n45257;
  assign n45259 = ~n45250 & n45255;
  assign n45260 = pi2  & ~n59306;
  assign n45261 = ~pi2  & n59306;
  assign n45262 = ~n45260 & ~n45261;
  assign n45263 = ~n39621 & n40023;
  assign n45264 = n24338 & ~n45263;
  assign n45265 = n25287 & n39621;
  assign n45266 = ~n56852 & n39626;
  assign n45267 = pi2  & n58457;
  assign n45268 = ~n45266 & n45267;
  assign n45269 = ~n45265 & n45268;
  assign n45270 = pi0  & ~n58457;
  assign n45271 = n25558 & ~n40039;
  assign n45272 = n24337 & ~n58457;
  assign n45273 = n25272 & n39626;
  assign n45274 = ~n45272 & ~n45273;
  assign n45275 = ~n45265 & n45274;
  assign n45276 = pi2  & ~n45275;
  assign n45277 = n25558 & ~n40023;
  assign n45278 = n25569 & ~n58457;
  assign n45279 = n25571 & n39626;
  assign n45280 = pi2  & ~n45279;
  assign n45281 = ~n45278 & n45280;
  assign n45282 = ~n45277 & n45281;
  assign n45283 = ~n45276 & n45282;
  assign n45284 = ~n45271 & n45283;
  assign n45285 = ~n45270 & n45284;
  assign n45286 = ~n24330 & ~n58457;
  assign n45287 = pi2  & ~n45270;
  assign n45288 = ~n45278 & n45287;
  assign n45289 = pi2  & ~n45286;
  assign n45290 = ~n45279 & n59308;
  assign n45291 = ~n45277 & n45290;
  assign n45292 = ~n45276 & n45291;
  assign n45293 = ~n45271 & n45292;
  assign n45294 = ~n45271 & n45291;
  assign n45295 = ~n45276 & n45294;
  assign n45296 = ~n45264 & n45269;
  assign n45297 = ~n43941 & ~n59307;
  assign n45298 = n24338 & n40006;
  assign n45299 = n25287 & n39618;
  assign n45300 = n24337 & n39626;
  assign n45301 = n25272 & n39621;
  assign n45302 = ~n45300 & ~n45301;
  assign n45303 = ~n45299 & n45302;
  assign n45304 = ~n45298 & n45303;
  assign n45305 = ~pi2  & ~n45304;
  assign n45306 = pi2  & n45304;
  assign n45307 = pi2  & ~n45304;
  assign n45308 = ~pi2  & n45304;
  assign n45309 = ~n45307 & ~n45308;
  assign n45310 = ~n45305 & ~n45306;
  assign n45311 = ~n45297 & n59309;
  assign n45312 = ~n45262 & n45311;
  assign n45313 = n45262 & ~n45311;
  assign n45314 = pi5  & n43941;
  assign n45315 = ~n43940 & n45314;
  assign n45316 = n43940 & ~n45314;
  assign n45317 = ~n43942 & n43946;
  assign n45318 = ~n59106 & ~n45317;
  assign n45319 = ~n45315 & ~n45316;
  assign n45320 = ~n45313 & n59310;
  assign n45321 = ~n45312 & ~n45320;
  assign n45322 = n59305 & ~n45321;
  assign n45323 = ~n59305 & n45321;
  assign n45324 = n24338 & n40071;
  assign n45325 = n25287 & n39612;
  assign n45326 = n24337 & n39618;
  assign n45327 = n25272 & n39615;
  assign n45328 = ~n45326 & ~n45327;
  assign n45329 = ~n45325 & n45328;
  assign n45330 = ~n45324 & n45329;
  assign n45331 = pi2  & ~n45330;
  assign n45332 = ~pi2  & n45330;
  assign n45333 = ~pi2  & ~n45330;
  assign n45334 = pi2  & n45330;
  assign n45335 = ~n45333 & ~n45334;
  assign n45336 = ~n45331 & ~n45332;
  assign n45337 = ~n45323 & ~n59311;
  assign n45338 = ~n45322 & ~n45337;
  assign n45339 = ~n45243 & ~n45338;
  assign n45340 = n45243 & n45338;
  assign n45341 = n43977 & n59113;
  assign n45342 = ~n43985 & ~n45341;
  assign n45343 = ~n45340 & n45342;
  assign n45344 = ~n45339 & ~n45343;
  assign n45345 = n45230 & ~n45344;
  assign n45346 = ~n45230 & n45344;
  assign n45347 = n24338 & n40183;
  assign n45348 = n25287 & n39606;
  assign n45349 = n24337 & n39612;
  assign n45350 = n25272 & n39609;
  assign n45351 = ~n45349 & ~n45350;
  assign n45352 = ~n45348 & n45351;
  assign n45353 = ~n45347 & n45352;
  assign n45354 = pi2  & ~n45353;
  assign n45355 = ~pi2  & n45353;
  assign n45356 = ~pi2  & ~n45353;
  assign n45357 = pi2  & n45353;
  assign n45358 = ~n45356 & ~n45357;
  assign n45359 = ~n45354 & ~n45355;
  assign n45360 = ~n45346 & ~n59312;
  assign n45361 = ~n45345 & ~n45360;
  assign n45362 = ~n45228 & ~n45361;
  assign n45363 = n45228 & n45361;
  assign n45364 = n43990 & n59116;
  assign n45365 = ~n43998 & ~n45364;
  assign n45366 = ~n45363 & n45365;
  assign n45367 = ~n45362 & ~n45366;
  assign n45368 = ~n45215 & ~n45367;
  assign n45369 = n45215 & n45367;
  assign n45370 = n43999 & ~n44001;
  assign n45371 = ~n44002 & ~n45370;
  assign n45372 = ~n45369 & n45371;
  assign n45373 = ~n45368 & ~n45372;
  assign n45374 = ~n45202 & ~n45373;
  assign n45375 = n45202 & n45373;
  assign n45376 = n44003 & n59119;
  assign n45377 = ~n44011 & ~n45376;
  assign n45378 = ~n45375 & n45377;
  assign n45379 = ~n45374 & ~n45378;
  assign n45380 = n45189 & ~n45379;
  assign n45381 = ~n45189 & n45379;
  assign n45382 = n24338 & n40476;
  assign n45383 = n25287 & n39594;
  assign n45384 = n24337 & n39600;
  assign n45385 = n25272 & n39597;
  assign n45386 = ~n45384 & ~n45385;
  assign n45387 = ~n45383 & n45386;
  assign n45388 = ~n45382 & n45387;
  assign n45389 = pi2  & ~n45388;
  assign n45390 = ~pi2  & n45388;
  assign n45391 = ~pi2  & ~n45388;
  assign n45392 = pi2  & n45388;
  assign n45393 = ~n45391 & ~n45392;
  assign n45394 = ~n45389 & ~n45390;
  assign n45395 = ~n45381 & ~n59313;
  assign n45396 = ~n45380 & ~n45395;
  assign n45397 = n45185 & ~n45396;
  assign n45398 = ~n45185 & n45396;
  assign n45399 = n24338 & n40616;
  assign n45400 = n25287 & n39591;
  assign n45401 = n24337 & n39597;
  assign n45402 = n25272 & n39594;
  assign n45403 = ~n45401 & ~n45402;
  assign n45404 = ~n45400 & n45403;
  assign n45405 = ~n45399 & n45404;
  assign n45406 = pi2  & ~n45405;
  assign n45407 = ~pi2  & n45405;
  assign n45408 = ~pi2  & ~n45405;
  assign n45409 = pi2  & n45405;
  assign n45410 = ~n45408 & ~n45409;
  assign n45411 = ~n45406 & ~n45407;
  assign n45412 = ~n45398 & ~n59314;
  assign n45413 = ~n45397 & ~n45412;
  assign n45414 = n45179 & ~n45413;
  assign n45415 = ~n45179 & n45413;
  assign n45416 = n24338 & ~n58585;
  assign n45417 = n25287 & n39588;
  assign n45418 = n24337 & n39594;
  assign n45419 = n25272 & n39591;
  assign n45420 = ~n45418 & ~n45419;
  assign n45421 = ~n45417 & n45420;
  assign n45422 = ~n45416 & n45421;
  assign n45423 = pi2  & ~n45422;
  assign n45424 = ~pi2  & n45422;
  assign n45425 = ~pi2  & ~n45422;
  assign n45426 = pi2  & n45422;
  assign n45427 = ~n45425 & ~n45426;
  assign n45428 = ~n45423 & ~n45424;
  assign n45429 = ~n45415 & ~n59315;
  assign n45430 = ~n45414 & ~n45429;
  assign n45431 = ~n45177 & ~n45430;
  assign n45432 = n45177 & n45430;
  assign n45433 = n44034 & n59126;
  assign n45434 = ~n44040 & ~n45433;
  assign n45435 = ~n45432 & n45434;
  assign n45436 = ~n45431 & ~n45435;
  assign n45437 = ~n45164 & ~n45436;
  assign n45438 = n45164 & n45436;
  assign n45439 = n44041 & n59129;
  assign n45440 = ~n44049 & ~n45439;
  assign n45441 = ~n45438 & n45440;
  assign n45442 = ~n45437 & ~n45441;
  assign n45443 = ~n45151 & ~n45442;
  assign n45444 = n45151 & n45442;
  assign n45445 = n44050 & n59132;
  assign n45446 = ~n44058 & ~n45445;
  assign n45447 = ~n45444 & n45446;
  assign n45448 = ~n45443 & ~n45447;
  assign n45449 = n45138 & ~n45448;
  assign n45450 = ~n45138 & n45448;
  assign n45451 = n24338 & ~n58653;
  assign n45452 = n25287 & n39576;
  assign n45453 = n24337 & n39582;
  assign n45454 = n25272 & n39579;
  assign n45455 = ~n45453 & ~n45454;
  assign n45456 = ~n45452 & n45455;
  assign n45457 = ~n45451 & n45456;
  assign n45458 = pi2  & ~n45457;
  assign n45459 = ~pi2  & n45457;
  assign n45460 = ~pi2  & ~n45457;
  assign n45461 = pi2  & n45457;
  assign n45462 = ~n45460 & ~n45461;
  assign n45463 = ~n45458 & ~n45459;
  assign n45464 = ~n45450 & ~n59316;
  assign n45465 = ~n45449 & ~n45464;
  assign n45466 = n45134 & ~n45465;
  assign n45467 = ~n45134 & n45465;
  assign n45468 = n24338 & n39976;
  assign n45469 = n25287 & n39573;
  assign n45470 = n24337 & n39579;
  assign n45471 = n25272 & n39576;
  assign n45472 = ~n45470 & ~n45471;
  assign n45473 = ~n45469 & n45472;
  assign n45474 = ~n45468 & n45473;
  assign n45475 = pi2  & ~n45474;
  assign n45476 = ~pi2  & n45474;
  assign n45477 = ~pi2  & ~n45474;
  assign n45478 = pi2  & n45474;
  assign n45479 = ~n45477 & ~n45478;
  assign n45480 = ~n45475 & ~n45476;
  assign n45481 = ~n45467 & ~n59317;
  assign n45482 = ~n45466 & ~n45481;
  assign n45483 = n45130 & ~n45482;
  assign n45484 = ~n45130 & n45482;
  assign n45485 = n24338 & ~n58759;
  assign n45486 = n25287 & n39570;
  assign n45487 = n24337 & n39576;
  assign n45488 = n25272 & n39573;
  assign n45489 = ~n45487 & ~n45488;
  assign n45490 = ~n45486 & n45489;
  assign n45491 = ~n45485 & n45490;
  assign n45492 = pi2  & ~n45491;
  assign n45493 = ~pi2  & n45491;
  assign n45494 = ~pi2  & ~n45491;
  assign n45495 = pi2  & n45491;
  assign n45496 = ~n45494 & ~n45495;
  assign n45497 = ~n45492 & ~n45493;
  assign n45498 = ~n45484 & ~n59318;
  assign n45499 = ~n45483 & ~n45498;
  assign n45500 = ~n45128 & ~n45499;
  assign n45501 = n45128 & n45499;
  assign n45502 = n44081 & n59141;
  assign n45503 = ~n44089 & ~n45502;
  assign n45504 = ~n45501 & n45503;
  assign n45505 = ~n45500 & ~n45504;
  assign n45506 = ~n45115 & ~n45505;
  assign n45507 = n45115 & n45505;
  assign n45508 = n44090 & n59142;
  assign n45509 = ~n44096 & ~n45508;
  assign n45510 = ~n45507 & n45509;
  assign n45511 = ~n45506 & ~n45510;
  assign n45512 = ~n45102 & ~n45511;
  assign n45513 = n45102 & n45511;
  assign n45514 = n44097 & n59145;
  assign n45515 = ~n44105 & ~n45514;
  assign n45516 = ~n45513 & n45515;
  assign n45517 = ~n45512 & ~n45516;
  assign n45518 = n45089 & ~n45517;
  assign n45519 = ~n45089 & n45517;
  assign n45520 = n24338 & ~n58849;
  assign n45521 = n25287 & n39558;
  assign n45522 = n24337 & n39564;
  assign n45523 = n25272 & n39561;
  assign n45524 = ~n45522 & ~n45523;
  assign n45525 = ~n45521 & n45524;
  assign n45526 = ~n45520 & n45525;
  assign n45527 = pi2  & ~n45526;
  assign n45528 = ~pi2  & n45526;
  assign n45529 = ~pi2  & ~n45526;
  assign n45530 = pi2  & n45526;
  assign n45531 = ~n45529 & ~n45530;
  assign n45532 = ~n45527 & ~n45528;
  assign n45533 = ~n45519 & ~n59319;
  assign n45534 = ~n45518 & ~n45533;
  assign n45535 = n45085 & ~n45534;
  assign n45536 = ~n45085 & n45534;
  assign n45537 = n24338 & n42574;
  assign n45538 = n25287 & n39555;
  assign n45539 = n24337 & n39561;
  assign n45540 = n25272 & n39558;
  assign n45541 = ~n45539 & ~n45540;
  assign n45542 = ~n45538 & n45541;
  assign n45543 = ~n45537 & n45542;
  assign n45544 = pi2  & ~n45543;
  assign n45545 = ~pi2  & n45543;
  assign n45546 = ~pi2  & ~n45543;
  assign n45547 = pi2  & n45543;
  assign n45548 = ~n45546 & ~n45547;
  assign n45549 = ~n45544 & ~n45545;
  assign n45550 = ~n45536 & ~n59320;
  assign n45551 = ~n45535 & ~n45550;
  assign n45552 = n45081 & ~n45551;
  assign n45553 = ~n45081 & n45551;
  assign n45554 = n24338 & ~n58891;
  assign n45555 = n25287 & n39552;
  assign n45556 = n24337 & n39558;
  assign n45557 = n25272 & n39555;
  assign n45558 = ~n45556 & ~n45557;
  assign n45559 = ~n45555 & n45558;
  assign n45560 = ~n45554 & n45559;
  assign n45561 = pi2  & ~n45560;
  assign n45562 = ~pi2  & n45560;
  assign n45563 = ~pi2  & ~n45560;
  assign n45564 = pi2  & n45560;
  assign n45565 = ~n45563 & ~n45564;
  assign n45566 = ~n45561 & ~n45562;
  assign n45567 = ~n45553 & ~n59321;
  assign n45568 = ~n45552 & ~n45567;
  assign n45569 = ~n45079 & ~n45568;
  assign n45570 = n45079 & n45568;
  assign n45571 = n44128 & n59152;
  assign n45572 = ~n44134 & ~n45571;
  assign n45573 = ~n45570 & n45572;
  assign n45574 = ~n45569 & ~n45573;
  assign n45575 = ~n45066 & ~n45574;
  assign n45576 = n45066 & n45574;
  assign n45577 = n44135 & n59155;
  assign n45578 = ~n44143 & ~n45577;
  assign n45579 = ~n45576 & n45578;
  assign n45580 = ~n45575 & ~n45579;
  assign n45581 = ~n45053 & ~n45580;
  assign n45582 = n45053 & n45580;
  assign n45583 = n44144 & n59158;
  assign n45584 = ~n44152 & ~n45583;
  assign n45585 = ~n45582 & n45584;
  assign n45586 = ~n45581 & ~n45585;
  assign n45587 = n45040 & ~n45586;
  assign n45588 = ~n45040 & n45586;
  assign n45589 = n24338 & ~n59044;
  assign n45590 = n25287 & n39543;
  assign n45591 = n24337 & n39546;
  assign n45592 = n25272 & n39440;
  assign n45593 = ~n45591 & ~n45592;
  assign n45594 = ~n45590 & n45593;
  assign n45595 = ~n45589 & n45594;
  assign n45596 = pi2  & ~n45595;
  assign n45597 = ~pi2  & n45595;
  assign n45598 = ~pi2  & ~n45595;
  assign n45599 = pi2  & n45595;
  assign n45600 = ~n45598 & ~n45599;
  assign n45601 = ~n45596 & ~n45597;
  assign n45602 = ~n45588 & ~n59322;
  assign n45603 = ~n45587 & ~n45602;
  assign n45604 = n45036 & ~n45603;
  assign n45605 = ~n45036 & n45603;
  assign n45606 = n24338 & n39943;
  assign n45607 = n25287 & n39937;
  assign n45608 = n24337 & n39440;
  assign n45609 = n25272 & n39543;
  assign n45610 = ~n45608 & ~n45609;
  assign n45611 = ~n45607 & n45610;
  assign n45612 = ~n45606 & n45611;
  assign n45613 = pi2  & ~n45612;
  assign n45614 = ~pi2  & n45612;
  assign n45615 = ~pi2  & ~n45612;
  assign n45616 = pi2  & n45612;
  assign n45617 = ~n45615 & ~n45616;
  assign n45618 = ~n45613 & ~n45614;
  assign n45619 = ~n45605 & ~n59323;
  assign n45620 = ~n45604 & ~n45619;
  assign n45621 = ~n45034 & ~n45620;
  assign n45622 = n45034 & n45620;
  assign n45623 = n44166 & n59162;
  assign n45624 = ~n44172 & ~n45623;
  assign n45625 = ~n45622 & n45624;
  assign n45626 = ~n45621 & ~n45625;
  assign n45627 = ~n45021 & ~n45626;
  assign n45628 = n45021 & n45626;
  assign n45629 = n44173 & n59163;
  assign n45630 = ~n44179 & ~n45629;
  assign n45631 = ~n45628 & n45630;
  assign n45632 = ~n45627 & ~n45631;
  assign n45633 = ~n45003 & ~n45632;
  assign n45634 = n45003 & n45632;
  assign n45635 = n44180 & n59166;
  assign n45636 = ~n44188 & ~n45635;
  assign n45637 = ~n45634 & n45636;
  assign n45638 = ~n45633 & ~n45637;
  assign n45639 = ~n59279 & ~n45638;
  assign n45640 = ~n44978 & ~n45639;
  assign n45641 = ~n44639 & ~n44648;
  assign n45642 = n77 & ~n59282;
  assign n45643 = n24302 & n44775;
  assign n45644 = n21969 & n39937;
  assign n45645 = n23459 & n44327;
  assign n45646 = ~n45644 & ~n45645;
  assign n45647 = ~n45643 & n45646;
  assign n45648 = ~n45642 & n45647;
  assign n45649 = pi5  & ~n45648;
  assign n45650 = ~n45648 & ~n45649;
  assign n45651 = ~pi5  & ~n45648;
  assign n45652 = pi5  & ~n45649;
  assign n45653 = pi5  & n45648;
  assign n45654 = ~n59324 & ~n59325;
  assign n45655 = ~n44625 & ~n44633;
  assign n45656 = ~n44603 & ~n44610;
  assign n45657 = n18846 & ~n58889;
  assign n45658 = n19541 & n39549;
  assign n45659 = n55247 & n39555;
  assign n45660 = n19509 & n39552;
  assign n45661 = ~n45659 & ~n45660;
  assign n45662 = ~n45658 & n45661;
  assign n45663 = ~n45657 & n45662;
  assign n45664 = pi11  & ~n45663;
  assign n45665 = ~n45663 & ~n45664;
  assign n45666 = ~pi11  & ~n45663;
  assign n45667 = pi11  & ~n45664;
  assign n45668 = pi11  & n45663;
  assign n45669 = ~n59326 & ~n59327;
  assign n45670 = ~n44587 & ~n44595;
  assign n45671 = ~n44563 & ~n44572;
  assign n45672 = n16079 & ~n58766;
  assign n45673 = n16696 & n39567;
  assign n45674 = n54886 & n39573;
  assign n45675 = n16676 & n39570;
  assign n45676 = ~n45674 & ~n45675;
  assign n45677 = ~n45673 & n45676;
  assign n45678 = ~n45672 & n45677;
  assign n45679 = pi17  & ~n45678;
  assign n45680 = ~n45678 & ~n45679;
  assign n45681 = ~pi17  & ~n45678;
  assign n45682 = pi17  & ~n45679;
  assign n45683 = pi17  & n45678;
  assign n45684 = ~n59328 & ~n59329;
  assign n45685 = ~n44549 & ~n44557;
  assign n45686 = ~n44527 & ~n44534;
  assign n45687 = n90 & ~n58583;
  assign n45688 = n14236 & n39585;
  assign n45689 = n54667 & n39591;
  assign n45690 = n14210 & n39588;
  assign n45691 = ~n45689 & ~n45690;
  assign n45692 = ~n45688 & n45691;
  assign n45693 = ~n45687 & n45692;
  assign n45694 = pi23  & ~n45693;
  assign n45695 = ~n45693 & ~n45694;
  assign n45696 = ~pi23  & ~n45693;
  assign n45697 = pi23  & ~n45694;
  assign n45698 = pi23  & n45693;
  assign n45699 = ~n59330 & ~n59331;
  assign n45700 = ~n44511 & ~n44519;
  assign n45701 = ~n44487 & ~n44496;
  assign n45702 = n11279 & n40286;
  assign n45703 = n12584 & n39603;
  assign n45704 = n54410 & n39609;
  assign n45705 = n11267 & n39606;
  assign n45706 = ~n45704 & ~n45705;
  assign n45707 = ~n45703 & n45706;
  assign n45708 = ~n45702 & n45707;
  assign n45709 = pi29  & ~n45708;
  assign n45710 = ~n45708 & ~n45709;
  assign n45711 = ~pi29  & ~n45708;
  assign n45712 = pi29  & ~n45709;
  assign n45713 = pi29  & n45708;
  assign n45714 = ~n59332 & ~n59333;
  assign n45715 = ~n44473 & ~n44481;
  assign n45716 = n916 & n7209;
  assign n45717 = n26637 & n45716;
  assign n45718 = n54732 & n45717;
  assign n45719 = n56590 & n45718;
  assign n45720 = ~n1477 & n3273;
  assign n45721 = n4094 & n6482;
  assign n45722 = n45720 & n45721;
  assign n45723 = n7212 & n54121;
  assign n45724 = n45722 & n45723;
  assign n45725 = n54512 & n45724;
  assign n45726 = n916 & n5390;
  assign n45727 = n3273 & n4094;
  assign n45728 = n45726 & n45727;
  assign n45729 = n54732 & n45728;
  assign n45730 = n56590 & n45729;
  assign n45731 = ~n625 & ~n1641;
  assign n45732 = ~n174 & ~n499;
  assign n45733 = n7209 & n26637;
  assign n45734 = n45731 & n45732;
  assign n45735 = n3014 & n6482;
  assign n45736 = n59334 & n45735;
  assign n45737 = n54121 & n45736;
  assign n45738 = n54512 & n45737;
  assign n45739 = n45730 & n45738;
  assign n45740 = n3014 & n4094;
  assign n45741 = n45726 & n45740;
  assign n45742 = n54732 & n45741;
  assign n45743 = n56590 & n45742;
  assign n45744 = n3273 & n6482;
  assign n45745 = n59334 & n45744;
  assign n45746 = n54121 & n45745;
  assign n45747 = n54512 & n45746;
  assign n45748 = n45743 & n45747;
  assign n45749 = n45719 & n45725;
  assign n45750 = n54626 & n59335;
  assign n45751 = n916 & n56618;
  assign n45752 = n54732 & n45751;
  assign n45753 = n54121 & n45752;
  assign n45754 = n3273 & n45753;
  assign n45755 = n56590 & n45754;
  assign n45756 = n54626 & n45755;
  assign n45757 = n54512 & n45756;
  assign n45758 = n4094 & n45757;
  assign n45759 = n5390 & n45758;
  assign n45760 = n6482 & n45759;
  assign n45761 = n3014 & n45760;
  assign n45762 = ~n174 & n45761;
  assign n45763 = ~n1641 & n45762;
  assign n45764 = ~n499 & n45763;
  assign n45765 = ~n625 & n45764;
  assign n45766 = n56618 & n45750;
  assign n45767 = n1576 & n40071;
  assign n45768 = n11215 & n39612;
  assign n45769 = n10564 & n39615;
  assign n45770 = n54403 & n39618;
  assign n45771 = ~n45769 & ~n45770;
  assign n45772 = ~n45768 & n45771;
  assign n45773 = ~n45767 & ~n45770;
  assign n45774 = ~n45769 & n45773;
  assign n45775 = ~n45768 & n45774;
  assign n45776 = ~n45767 & n45772;
  assign n45777 = ~n59336 & ~n59337;
  assign n45778 = n59336 & n59337;
  assign n45779 = ~n59336 & ~n45777;
  assign n45780 = ~n59336 & n59337;
  assign n45781 = ~n59337 & ~n45777;
  assign n45782 = n59336 & ~n59337;
  assign n45783 = ~n59338 & ~n59339;
  assign n45784 = ~n45777 & ~n45778;
  assign n45785 = ~n45715 & ~n59340;
  assign n45786 = n45715 & n59340;
  assign n45787 = ~n45715 & ~n45785;
  assign n45788 = ~n59340 & ~n45785;
  assign n45789 = ~n45787 & ~n45788;
  assign n45790 = ~n45785 & ~n45786;
  assign n45791 = ~n45714 & ~n59341;
  assign n45792 = n45714 & n59341;
  assign n45793 = ~n45714 & ~n45791;
  assign n45794 = ~n45714 & n59341;
  assign n45795 = ~n59341 & ~n45791;
  assign n45796 = n45714 & ~n59341;
  assign n45797 = ~n59342 & ~n59343;
  assign n45798 = ~n45791 & ~n45792;
  assign n45799 = n45701 & n59344;
  assign n45800 = ~n45701 & ~n59344;
  assign n45801 = ~n45799 & ~n45800;
  assign n45802 = n123 & n40476;
  assign n45803 = n128 & n39594;
  assign n45804 = n53444 & n39600;
  assign n45805 = n127 & n39597;
  assign n45806 = ~n45804 & ~n45805;
  assign n45807 = ~n45803 & n45806;
  assign n45808 = ~n123 & n45807;
  assign n45809 = ~n40476 & n45807;
  assign n45810 = ~n45808 & ~n45809;
  assign n45811 = ~n45802 & n45807;
  assign n45812 = pi26  & ~n59345;
  assign n45813 = ~pi26  & n59345;
  assign n45814 = ~n45812 & ~n45813;
  assign n45815 = n45801 & ~n45814;
  assign n45816 = ~n45801 & n45814;
  assign n45817 = n45801 & ~n45815;
  assign n45818 = n45801 & n45814;
  assign n45819 = ~n45814 & ~n45815;
  assign n45820 = ~n45801 & ~n45814;
  assign n45821 = ~n59346 & ~n59347;
  assign n45822 = ~n45815 & ~n45816;
  assign n45823 = ~n45700 & ~n59348;
  assign n45824 = n45700 & n59348;
  assign n45825 = ~n45700 & ~n45823;
  assign n45826 = ~n45700 & n59348;
  assign n45827 = ~n59348 & ~n45823;
  assign n45828 = n45700 & ~n59348;
  assign n45829 = ~n59349 & ~n59350;
  assign n45830 = ~n45823 & ~n45824;
  assign n45831 = ~n45699 & ~n59351;
  assign n45832 = n45699 & n59351;
  assign n45833 = ~n45699 & ~n45831;
  assign n45834 = ~n59351 & ~n45831;
  assign n45835 = ~n45833 & ~n45834;
  assign n45836 = ~n45831 & ~n45832;
  assign n45837 = n45686 & n59352;
  assign n45838 = ~n45686 & ~n59352;
  assign n45839 = ~n45837 & ~n45838;
  assign n45840 = n14413 & ~n58653;
  assign n45841 = n15921 & n39576;
  assign n45842 = n54719 & n39582;
  assign n45843 = n15901 & n39579;
  assign n45844 = ~n45842 & ~n45843;
  assign n45845 = ~n45841 & n45844;
  assign n45846 = ~n14413 & n45845;
  assign n45847 = n58653 & n45845;
  assign n45848 = ~n45846 & ~n45847;
  assign n45849 = ~n45840 & n45845;
  assign n45850 = pi20  & ~n59353;
  assign n45851 = ~pi20  & n59353;
  assign n45852 = ~n45850 & ~n45851;
  assign n45853 = n45839 & ~n45852;
  assign n45854 = ~n45839 & n45852;
  assign n45855 = n45839 & ~n45853;
  assign n45856 = n45839 & n45852;
  assign n45857 = ~n45852 & ~n45853;
  assign n45858 = ~n45839 & ~n45852;
  assign n45859 = ~n59354 & ~n59355;
  assign n45860 = ~n45853 & ~n45854;
  assign n45861 = ~n45685 & ~n59356;
  assign n45862 = n45685 & n59356;
  assign n45863 = ~n45685 & ~n45861;
  assign n45864 = ~n59356 & ~n45861;
  assign n45865 = ~n45863 & ~n45864;
  assign n45866 = ~n45861 & ~n45862;
  assign n45867 = ~n45684 & ~n59357;
  assign n45868 = n45684 & n59357;
  assign n45869 = ~n45684 & ~n45867;
  assign n45870 = ~n45684 & n59357;
  assign n45871 = ~n59357 & ~n45867;
  assign n45872 = n45684 & ~n59357;
  assign n45873 = ~n59358 & ~n59359;
  assign n45874 = ~n45867 & ~n45868;
  assign n45875 = n45671 & n59360;
  assign n45876 = ~n45671 & ~n59360;
  assign n45877 = ~n45875 & ~n45876;
  assign n45878 = n17265 & ~n58849;
  assign n45879 = n18588 & n39558;
  assign n45880 = n55041 & n39564;
  assign n45881 = n18556 & n39561;
  assign n45882 = ~n45880 & ~n45881;
  assign n45883 = ~n45879 & n45882;
  assign n45884 = ~n17265 & n45883;
  assign n45885 = n58849 & n45883;
  assign n45886 = ~n45884 & ~n45885;
  assign n45887 = ~n45878 & n45883;
  assign n45888 = pi14  & ~n59361;
  assign n45889 = ~pi14  & n59361;
  assign n45890 = ~n45888 & ~n45889;
  assign n45891 = n45877 & ~n45890;
  assign n45892 = ~n45877 & n45890;
  assign n45893 = n45877 & ~n45891;
  assign n45894 = n45877 & n45890;
  assign n45895 = ~n45890 & ~n45891;
  assign n45896 = ~n45877 & ~n45890;
  assign n45897 = ~n59362 & ~n59363;
  assign n45898 = ~n45891 & ~n45892;
  assign n45899 = ~n45670 & ~n59364;
  assign n45900 = n45670 & n59364;
  assign n45901 = ~n45670 & ~n45899;
  assign n45902 = ~n45670 & n59364;
  assign n45903 = ~n59364 & ~n45899;
  assign n45904 = n45670 & ~n59364;
  assign n45905 = ~n59365 & ~n59366;
  assign n45906 = ~n45899 & ~n45900;
  assign n45907 = ~n45669 & ~n59367;
  assign n45908 = n45669 & n59367;
  assign n45909 = ~n45669 & ~n45907;
  assign n45910 = ~n59367 & ~n45907;
  assign n45911 = ~n45909 & ~n45910;
  assign n45912 = ~n45907 & ~n45908;
  assign n45913 = n45656 & n59368;
  assign n45914 = ~n45656 & ~n59368;
  assign n45915 = ~n45913 & ~n45914;
  assign n45916 = n20085 & ~n59044;
  assign n45917 = n21269 & n39543;
  assign n45918 = n55472 & n39546;
  assign n45919 = n21237 & n39440;
  assign n45920 = ~n45918 & ~n45919;
  assign n45921 = ~n45917 & n45920;
  assign n45922 = ~n20085 & n45921;
  assign n45923 = n59044 & n45921;
  assign n45924 = ~n45922 & ~n45923;
  assign n45925 = ~n45916 & n45921;
  assign n45926 = pi8  & ~n59369;
  assign n45927 = ~pi8  & n59369;
  assign n45928 = ~n45926 & ~n45927;
  assign n45929 = n45915 & ~n45928;
  assign n45930 = ~n45915 & n45928;
  assign n45931 = n45915 & ~n45929;
  assign n45932 = n45915 & n45928;
  assign n45933 = ~n45928 & ~n45929;
  assign n45934 = ~n45915 & ~n45928;
  assign n45935 = ~n59370 & ~n59371;
  assign n45936 = ~n45929 & ~n45930;
  assign n45937 = ~n45655 & ~n59372;
  assign n45938 = n45655 & n59372;
  assign n45939 = ~n45655 & ~n45937;
  assign n45940 = ~n59372 & ~n45937;
  assign n45941 = ~n45939 & ~n45940;
  assign n45942 = ~n45937 & ~n45938;
  assign n45943 = ~n45654 & ~n59373;
  assign n45944 = n45654 & n59373;
  assign n45945 = ~n45654 & ~n45943;
  assign n45946 = ~n45654 & n59373;
  assign n45947 = ~n59373 & ~n45943;
  assign n45948 = n45654 & ~n59373;
  assign n45949 = ~n59374 & ~n59375;
  assign n45950 = ~n45943 & ~n45944;
  assign n45951 = n45641 & n59376;
  assign n45952 = ~n45641 & ~n59376;
  assign n45953 = ~n45951 & ~n45952;
  assign n45954 = ~n44947 & ~n44951;
  assign n45955 = ~n44937 & ~n44944;
  assign n45956 = ~n44915 & ~n44917;
  assign n45957 = ~n1081 & n53563;
  assign n45958 = n53640 & n45957;
  assign n45959 = n53563 & n53640;
  assign n45960 = n59269 & n45959;
  assign n45961 = ~n1081 & n45960;
  assign n45962 = n59269 & n45958;
  assign n45963 = ~n45956 & n59377;
  assign n45964 = n45956 & ~n59377;
  assign n45965 = ~n45963 & ~n45964;
  assign n45966 = n1576 & n27808;
  assign n45967 = n11215 & n26242;
  assign n45968 = n10564 & n26244;
  assign n45969 = ~n59271 & ~n45968;
  assign n45970 = ~n45967 & n45969;
  assign n45971 = ~n45966 & n45970;
  assign n45972 = n45965 & ~n45971;
  assign n45973 = ~n45965 & n45971;
  assign n45974 = ~n45971 & ~n45972;
  assign n45975 = n45965 & ~n45972;
  assign n45976 = ~n45974 & ~n45975;
  assign n45977 = ~n45972 & ~n45973;
  assign n45978 = ~n44920 & n44930;
  assign n45979 = ~n44920 & ~n44931;
  assign n45980 = ~n44921 & ~n45978;
  assign n45981 = n59378 & n59379;
  assign n45982 = ~n59378 & ~n59379;
  assign n45983 = ~n45981 & ~n45982;
  assign n45984 = ~n54408 & ~n11279;
  assign n45985 = ~n11267 & ~n12584;
  assign n45986 = ~n11267 & ~n54410;
  assign n45987 = ~n12584 & n45986;
  assign n45988 = ~n54410 & ~n12584;
  assign n45989 = ~n11267 & n45988;
  assign n45990 = ~n54410 & ~n59380;
  assign n45991 = ~n11279 & n59381;
  assign n45992 = ~n54407 & n45986;
  assign n45993 = n54408 & ~n54410;
  assign n45994 = n54408 & ~n54409;
  assign n45995 = pi29  & ~n59382;
  assign n45996 = pi29  & ~n45995;
  assign n45997 = pi29  & n59382;
  assign n45998 = ~n59382 & ~n45995;
  assign n45999 = ~pi29  & ~n59382;
  assign n46000 = ~n59383 & ~n59384;
  assign n46001 = n45983 & ~n46000;
  assign n46002 = ~n45983 & n46000;
  assign n46003 = ~n46001 & ~n46002;
  assign n46004 = ~n45955 & n46003;
  assign n46005 = n45955 & ~n46003;
  assign n46006 = ~n46004 & ~n46005;
  assign n46007 = ~n45954 & n46006;
  assign n46008 = n45954 & ~n46006;
  assign n46009 = ~n46007 & ~n46008;
  assign n46010 = n44952 & n46009;
  assign n46011 = ~n44952 & ~n46009;
  assign n46012 = ~n46010 & ~n46011;
  assign n46013 = ~n44961 & ~n46011;
  assign n46014 = ~n46010 & n46013;
  assign n46015 = ~n44961 & n46012;
  assign n46016 = n44961 & ~n46012;
  assign n46017 = ~n44961 & ~n59385;
  assign n46018 = ~n46010 & ~n59385;
  assign n46019 = ~n46011 & n46018;
  assign n46020 = ~n46017 & ~n46019;
  assign n46021 = ~n59385 & ~n46016;
  assign n46022 = n24338 & ~n59386;
  assign n46023 = n25287 & n46009;
  assign n46024 = n24337 & n44871;
  assign n46025 = n25272 & n44952;
  assign n46026 = ~n46024 & ~n46025;
  assign n46027 = ~n46023 & n46026;
  assign n46028 = ~n24338 & n46027;
  assign n46029 = n59386 & n46027;
  assign n46030 = ~n46028 & ~n46029;
  assign n46031 = ~n46022 & n46027;
  assign n46032 = pi2  & ~n59387;
  assign n46033 = ~pi2  & n59387;
  assign n46034 = ~n46032 & ~n46033;
  assign n46035 = n45953 & ~n46034;
  assign n46036 = ~n45953 & n46034;
  assign n46037 = ~n46035 & ~n46036;
  assign n46038 = ~n45640 & n46037;
  assign n46039 = n45640 & ~n46037;
  assign n46040 = ~n46038 & ~n46039;
  assign n46041 = n59279 & n45638;
  assign n46042 = ~n45638 & ~n45639;
  assign n46043 = n59279 & ~n45638;
  assign n46044 = ~n59279 & ~n45639;
  assign n46045 = ~n59279 & n45638;
  assign n46046 = ~n59388 & ~n59389;
  assign n46047 = ~n45639 & ~n46041;
  assign n46048 = n46040 & ~n59390;
  assign n46049 = ~n46040 & n59390;
  assign n46050 = n46040 & n59390;
  assign n46051 = ~n46040 & ~n59390;
  assign n46052 = ~n46050 & ~n46051;
  assign n46053 = ~n46048 & ~n46049;
  assign n46054 = ~n46035 & ~n46038;
  assign n46055 = ~n45943 & ~n45952;
  assign n46056 = n77 & ~n59280;
  assign n46057 = n24302 & n44871;
  assign n46058 = n21969 & n44327;
  assign n46059 = n23459 & n44775;
  assign n46060 = ~n46058 & ~n46059;
  assign n46061 = ~n46057 & n46060;
  assign n46062 = ~n46056 & n46061;
  assign n46063 = pi5  & ~n46062;
  assign n46064 = ~n46062 & ~n46063;
  assign n46065 = ~pi5  & ~n46062;
  assign n46066 = pi5  & ~n46063;
  assign n46067 = pi5  & n46062;
  assign n46068 = ~n59392 & ~n59393;
  assign n46069 = ~n45929 & ~n45937;
  assign n46070 = ~n45907 & ~n45914;
  assign n46071 = n18846 & n43436;
  assign n46072 = n19541 & n39546;
  assign n46073 = n55247 & n39552;
  assign n46074 = n19509 & n39549;
  assign n46075 = ~n46073 & ~n46074;
  assign n46076 = ~n46072 & n46075;
  assign n46077 = ~n46071 & n46076;
  assign n46078 = pi11  & ~n46077;
  assign n46079 = ~n46077 & ~n46078;
  assign n46080 = ~pi11  & ~n46077;
  assign n46081 = pi11  & ~n46078;
  assign n46082 = pi11  & n46077;
  assign n46083 = ~n59394 & ~n59395;
  assign n46084 = ~n45891 & ~n45899;
  assign n46085 = ~n45867 & ~n45876;
  assign n46086 = n16079 & n41762;
  assign n46087 = n16696 & n39564;
  assign n46088 = n54886 & n39570;
  assign n46089 = n16676 & n39567;
  assign n46090 = ~n46088 & ~n46089;
  assign n46091 = ~n46087 & n46090;
  assign n46092 = ~n46086 & n46091;
  assign n46093 = pi17  & ~n46092;
  assign n46094 = ~n46092 & ~n46093;
  assign n46095 = ~pi17  & ~n46092;
  assign n46096 = pi17  & ~n46093;
  assign n46097 = pi17  & n46092;
  assign n46098 = ~n59396 & ~n59397;
  assign n46099 = ~n45853 & ~n45861;
  assign n46100 = ~n45831 & ~n45838;
  assign n46101 = n90 & n41007;
  assign n46102 = n14236 & n39582;
  assign n46103 = n54667 & n39588;
  assign n46104 = n14210 & n39585;
  assign n46105 = ~n46103 & ~n46104;
  assign n46106 = ~n46102 & n46105;
  assign n46107 = ~n46101 & n46106;
  assign n46108 = pi23  & ~n46107;
  assign n46109 = ~n46107 & ~n46108;
  assign n46110 = ~pi23  & ~n46107;
  assign n46111 = pi23  & ~n46108;
  assign n46112 = pi23  & n46107;
  assign n46113 = ~n59398 & ~n59399;
  assign n46114 = ~n45815 & ~n45823;
  assign n46115 = ~n45791 & ~n45800;
  assign n46116 = n11279 & ~n58533;
  assign n46117 = n12584 & n39600;
  assign n46118 = n54410 & n39606;
  assign n46119 = n11267 & n39603;
  assign n46120 = ~n46118 & ~n46119;
  assign n46121 = ~n46117 & n46120;
  assign n46122 = ~n11279 & n46121;
  assign n46123 = n58533 & n46121;
  assign n46124 = ~n46122 & ~n46123;
  assign n46125 = ~n46116 & n46121;
  assign n46126 = pi29  & ~n59400;
  assign n46127 = ~pi29  & n59400;
  assign n46128 = ~n46126 & ~n46127;
  assign n46129 = ~n45777 & ~n45785;
  assign n46130 = n6482 & n6626;
  assign n46131 = n7005 & n46130;
  assign n46132 = ~n346 & ~n415;
  assign n46133 = ~n496 & ~n1457;
  assign n46134 = ~n346 & ~n496;
  assign n46135 = ~n415 & ~n1457;
  assign n46136 = n46134 & n46135;
  assign n46137 = n46132 & n46133;
  assign n46138 = n424 & n3776;
  assign n46139 = n59401 & n46138;
  assign n46140 = n46131 & n46139;
  assign n46141 = n55112 & n46140;
  assign n46142 = n3476 & n7144;
  assign n46143 = n53752 & n54161;
  assign n46144 = n46142 & n46143;
  assign n46145 = n55132 & n46144;
  assign n46146 = n7005 & n7144;
  assign n46147 = n424 & n46146;
  assign n46148 = ~n415 & ~n496;
  assign n46149 = n3776 & n46148;
  assign n46150 = n3476 & n6482;
  assign n46151 = n46149 & n46150;
  assign n46152 = n46147 & n46151;
  assign n46153 = n55112 & n46152;
  assign n46154 = ~n346 & ~n1457;
  assign n46155 = n6626 & n46154;
  assign n46156 = n53752 & n46155;
  assign n46157 = n54161 & n46156;
  assign n46158 = n55132 & n46157;
  assign n46159 = n46153 & n46158;
  assign n46160 = n3476 & n46146;
  assign n46161 = ~n415 & ~n464;
  assign n46162 = n424 & n46161;
  assign n46163 = n3776 & n6482;
  assign n46164 = n46162 & n46163;
  assign n46165 = n46160 & n46164;
  assign n46166 = n55112 & n46165;
  assign n46167 = ~n268 & ~n346;
  assign n46168 = n46133 & n46167;
  assign n46169 = n54161 & n46168;
  assign n46170 = n53752 & n46169;
  assign n46171 = n55132 & n46170;
  assign n46172 = n46166 & n46171;
  assign n46173 = n46141 & n46145;
  assign n46174 = n54250 & n56744;
  assign n46175 = n59402 & n46174;
  assign n46176 = n53752 & n7005;
  assign n46177 = n54161 & n46176;
  assign n46178 = n55112 & n46177;
  assign n46179 = n56744 & n46178;
  assign n46180 = n55132 & n46179;
  assign n46181 = n53787 & n46180;
  assign n46182 = n3476 & n46181;
  assign n46183 = n7144 & n46182;
  assign n46184 = n424 & n46183;
  assign n46185 = n6482 & n46184;
  assign n46186 = n54250 & n46185;
  assign n46187 = n3776 & n46186;
  assign n46188 = ~n415 & n46187;
  assign n46189 = ~n464 & n46188;
  assign n46190 = ~n1457 & n46189;
  assign n46191 = ~n268 & n46190;
  assign n46192 = ~n496 & n46191;
  assign n46193 = ~n346 & n46192;
  assign n46194 = n53787 & n46175;
  assign n46195 = n1576 & n39991;
  assign n46196 = n11215 & n39609;
  assign n46197 = n10564 & n39612;
  assign n46198 = n54403 & n39615;
  assign n46199 = ~n46197 & ~n46198;
  assign n46200 = ~n46196 & n46199;
  assign n46201 = ~n46195 & ~n46198;
  assign n46202 = ~n46197 & n46201;
  assign n46203 = ~n46196 & n46202;
  assign n46204 = ~n46195 & n46200;
  assign n46205 = ~n59403 & ~n59404;
  assign n46206 = n59403 & n59404;
  assign n46207 = ~n59403 & ~n46205;
  assign n46208 = ~n59403 & n59404;
  assign n46209 = ~n59404 & ~n46205;
  assign n46210 = n59403 & ~n59404;
  assign n46211 = ~n59405 & ~n59406;
  assign n46212 = ~n46205 & ~n46206;
  assign n46213 = ~n46129 & ~n59407;
  assign n46214 = n46129 & n59407;
  assign n46215 = ~n46129 & ~n46213;
  assign n46216 = ~n59407 & ~n46213;
  assign n46217 = ~n46215 & ~n46216;
  assign n46218 = ~n46213 & ~n46214;
  assign n46219 = ~n46128 & ~n59408;
  assign n46220 = n46128 & n59408;
  assign n46221 = ~n46219 & ~n46220;
  assign n46222 = ~n46115 & n46221;
  assign n46223 = n46115 & ~n46221;
  assign n46224 = ~n46222 & ~n46223;
  assign n46225 = n123 & n40616;
  assign n46226 = n128 & n39591;
  assign n46227 = n53444 & n39597;
  assign n46228 = n127 & n39594;
  assign n46229 = ~n46227 & ~n46228;
  assign n46230 = ~n46226 & n46229;
  assign n46231 = ~n123 & n46230;
  assign n46232 = ~n40616 & n46230;
  assign n46233 = ~n46231 & ~n46232;
  assign n46234 = ~n46225 & n46230;
  assign n46235 = pi26  & ~n59409;
  assign n46236 = ~pi26  & n59409;
  assign n46237 = ~n46235 & ~n46236;
  assign n46238 = n46224 & ~n46237;
  assign n46239 = ~n46224 & n46237;
  assign n46240 = n46224 & ~n46238;
  assign n46241 = n46224 & n46237;
  assign n46242 = ~n46237 & ~n46238;
  assign n46243 = ~n46224 & ~n46237;
  assign n46244 = ~n59410 & ~n59411;
  assign n46245 = ~n46238 & ~n46239;
  assign n46246 = ~n46114 & ~n59412;
  assign n46247 = n46114 & n59412;
  assign n46248 = ~n46114 & ~n46246;
  assign n46249 = ~n59412 & ~n46246;
  assign n46250 = ~n46248 & ~n46249;
  assign n46251 = ~n46246 & ~n46247;
  assign n46252 = ~n46113 & ~n59413;
  assign n46253 = n46113 & n59413;
  assign n46254 = ~n46113 & ~n46252;
  assign n46255 = ~n46113 & n59413;
  assign n46256 = ~n59413 & ~n46252;
  assign n46257 = n46113 & ~n59413;
  assign n46258 = ~n59414 & ~n59415;
  assign n46259 = ~n46252 & ~n46253;
  assign n46260 = n46100 & n59416;
  assign n46261 = ~n46100 & ~n59416;
  assign n46262 = ~n46260 & ~n46261;
  assign n46263 = n14413 & n39976;
  assign n46264 = n15921 & n39573;
  assign n46265 = n54719 & n39579;
  assign n46266 = n15901 & n39576;
  assign n46267 = ~n46265 & ~n46266;
  assign n46268 = ~n46264 & n46267;
  assign n46269 = ~n14413 & n46268;
  assign n46270 = ~n39976 & n46268;
  assign n46271 = ~n46269 & ~n46270;
  assign n46272 = ~n46263 & n46268;
  assign n46273 = pi20  & ~n59417;
  assign n46274 = ~pi20  & n59417;
  assign n46275 = ~n46273 & ~n46274;
  assign n46276 = n46262 & ~n46275;
  assign n46277 = ~n46262 & n46275;
  assign n46278 = n46262 & ~n46276;
  assign n46279 = n46262 & n46275;
  assign n46280 = ~n46275 & ~n46276;
  assign n46281 = ~n46262 & ~n46275;
  assign n46282 = ~n59418 & ~n59419;
  assign n46283 = ~n46276 & ~n46277;
  assign n46284 = ~n46099 & ~n59420;
  assign n46285 = n46099 & n59420;
  assign n46286 = ~n46099 & ~n46284;
  assign n46287 = ~n46099 & n59420;
  assign n46288 = ~n59420 & ~n46284;
  assign n46289 = n46099 & ~n59420;
  assign n46290 = ~n59421 & ~n59422;
  assign n46291 = ~n46284 & ~n46285;
  assign n46292 = ~n46098 & ~n59423;
  assign n46293 = n46098 & n59423;
  assign n46294 = ~n46098 & ~n46292;
  assign n46295 = ~n59423 & ~n46292;
  assign n46296 = ~n46294 & ~n46295;
  assign n46297 = ~n46292 & ~n46293;
  assign n46298 = n46085 & n59424;
  assign n46299 = ~n46085 & ~n59424;
  assign n46300 = ~n46298 & ~n46299;
  assign n46301 = n17265 & n42574;
  assign n46302 = n18588 & n39555;
  assign n46303 = n55041 & n39561;
  assign n46304 = n18556 & n39558;
  assign n46305 = ~n46303 & ~n46304;
  assign n46306 = ~n46302 & n46305;
  assign n46307 = ~n17265 & n46306;
  assign n46308 = ~n42574 & n46306;
  assign n46309 = ~n46307 & ~n46308;
  assign n46310 = ~n46301 & n46306;
  assign n46311 = pi14  & ~n59425;
  assign n46312 = ~pi14  & n59425;
  assign n46313 = ~n46311 & ~n46312;
  assign n46314 = n46300 & ~n46313;
  assign n46315 = ~n46300 & n46313;
  assign n46316 = n46300 & ~n46314;
  assign n46317 = n46300 & n46313;
  assign n46318 = ~n46313 & ~n46314;
  assign n46319 = ~n46300 & ~n46313;
  assign n46320 = ~n59426 & ~n59427;
  assign n46321 = ~n46314 & ~n46315;
  assign n46322 = ~n46084 & ~n59428;
  assign n46323 = n46084 & n59428;
  assign n46324 = ~n46084 & ~n46322;
  assign n46325 = ~n59428 & ~n46322;
  assign n46326 = ~n46324 & ~n46325;
  assign n46327 = ~n46322 & ~n46323;
  assign n46328 = ~n46083 & ~n59429;
  assign n46329 = n46083 & n59429;
  assign n46330 = ~n46083 & ~n46328;
  assign n46331 = ~n46083 & n59429;
  assign n46332 = ~n59429 & ~n46328;
  assign n46333 = n46083 & ~n59429;
  assign n46334 = ~n59430 & ~n59431;
  assign n46335 = ~n46328 & ~n46329;
  assign n46336 = n46070 & n59432;
  assign n46337 = ~n46070 & ~n59432;
  assign n46338 = ~n46336 & ~n46337;
  assign n46339 = n20085 & n39943;
  assign n46340 = n21269 & n39937;
  assign n46341 = n55472 & n39440;
  assign n46342 = n21237 & n39543;
  assign n46343 = ~n46341 & ~n46342;
  assign n46344 = ~n46340 & n46343;
  assign n46345 = ~n20085 & n46344;
  assign n46346 = ~n39943 & n46344;
  assign n46347 = ~n46345 & ~n46346;
  assign n46348 = ~n46339 & n46344;
  assign n46349 = pi8  & ~n59433;
  assign n46350 = ~pi8  & n59433;
  assign n46351 = ~n46349 & ~n46350;
  assign n46352 = n46338 & ~n46351;
  assign n46353 = ~n46338 & n46351;
  assign n46354 = n46338 & ~n46352;
  assign n46355 = n46338 & n46351;
  assign n46356 = ~n46351 & ~n46352;
  assign n46357 = ~n46338 & ~n46351;
  assign n46358 = ~n59434 & ~n59435;
  assign n46359 = ~n46352 & ~n46353;
  assign n46360 = ~n46069 & ~n59436;
  assign n46361 = n46069 & n59436;
  assign n46362 = ~n46069 & ~n46360;
  assign n46363 = ~n46069 & n59436;
  assign n46364 = ~n59436 & ~n46360;
  assign n46365 = n46069 & ~n59436;
  assign n46366 = ~n59437 & ~n59438;
  assign n46367 = ~n46360 & ~n46361;
  assign n46368 = ~n46068 & ~n59439;
  assign n46369 = n46068 & n59439;
  assign n46370 = ~n46068 & ~n46368;
  assign n46371 = ~n59439 & ~n46368;
  assign n46372 = ~n46370 & ~n46371;
  assign n46373 = ~n46368 & ~n46369;
  assign n46374 = n46055 & n59440;
  assign n46375 = ~n46055 & ~n59440;
  assign n46376 = ~n46374 & ~n46375;
  assign n46377 = ~n46004 & ~n46007;
  assign n46378 = ~n45982 & ~n46001;
  assign n46379 = n53499 & n53565;
  assign n46380 = n59377 & ~n46379;
  assign n46381 = ~n59377 & n46379;
  assign n46382 = ~n46380 & ~n46381;
  assign n46383 = ~n45963 & n45971;
  assign n46384 = ~n45963 & ~n45972;
  assign n46385 = ~n45964 & ~n46383;
  assign n46386 = ~n46381 & ~n59441;
  assign n46387 = ~n46380 & n46386;
  assign n46388 = n46382 & ~n59441;
  assign n46389 = ~n46382 & n59441;
  assign n46390 = ~n59441 & ~n59442;
  assign n46391 = ~n46381 & ~n59442;
  assign n46392 = ~n46380 & n46391;
  assign n46393 = ~n46390 & ~n46392;
  assign n46394 = ~n59442 & ~n46389;
  assign n46395 = n1576 & ~n56564;
  assign n46396 = n54403 & n26244;
  assign n46397 = n10564 & n26242;
  assign n46398 = ~n46396 & ~n46397;
  assign n46399 = ~n11215 & n46398;
  assign n46400 = ~n46395 & n46399;
  assign n46401 = ~n46000 & ~n46400;
  assign n46402 = n46000 & n46400;
  assign n46403 = ~n46000 & ~n46401;
  assign n46404 = ~n46000 & n46400;
  assign n46405 = ~n46400 & ~n46401;
  assign n46406 = n46000 & ~n46400;
  assign n46407 = ~n59444 & ~n59445;
  assign n46408 = ~n46401 & ~n46402;
  assign n46409 = ~n59443 & ~n59446;
  assign n46410 = n59443 & n59446;
  assign n46411 = ~n59443 & n59446;
  assign n46412 = n59443 & ~n59446;
  assign n46413 = ~n46411 & ~n46412;
  assign n46414 = ~n46409 & ~n46410;
  assign n46415 = ~n46378 & ~n59447;
  assign n46416 = n46378 & n59447;
  assign n46417 = ~n46415 & ~n46416;
  assign n46418 = ~n46377 & n46417;
  assign n46419 = n46377 & ~n46417;
  assign n46420 = ~n46418 & ~n46419;
  assign n46421 = ~n46009 & ~n46420;
  assign n46422 = n46009 & n46420;
  assign n46423 = ~n46421 & ~n46422;
  assign n46424 = ~n46018 & n46423;
  assign n46425 = n46018 & ~n46423;
  assign n46426 = ~n46424 & ~n46425;
  assign n46427 = n24338 & n46426;
  assign n46428 = n25287 & n46420;
  assign n46429 = n24337 & n44952;
  assign n46430 = n25272 & n46009;
  assign n46431 = ~n46429 & ~n46430;
  assign n46432 = ~n46428 & n46431;
  assign n46433 = ~n24338 & n46432;
  assign n46434 = ~n46426 & n46432;
  assign n46435 = ~n46433 & ~n46434;
  assign n46436 = ~n46427 & n46432;
  assign n46437 = pi2  & ~n59448;
  assign n46438 = ~pi2  & n59448;
  assign n46439 = ~n46437 & ~n46438;
  assign n46440 = n46376 & ~n46439;
  assign n46441 = ~n46376 & n46439;
  assign n46442 = ~n46440 & ~n46441;
  assign n46443 = ~n46054 & n46442;
  assign n46444 = n46054 & ~n46442;
  assign n46445 = ~n46443 & ~n46444;
  assign n46446 = n46048 & n46445;
  assign n46447 = ~n46048 & ~n46445;
  assign po1  = ~n46446 & ~n46447;
  assign n46449 = ~n46440 & ~n46443;
  assign n46450 = ~n46368 & ~n46375;
  assign n46451 = n77 & ~n59275;
  assign n46452 = n24302 & n44952;
  assign n46453 = n21969 & n44775;
  assign n46454 = n23459 & n44871;
  assign n46455 = ~n46453 & ~n46454;
  assign n46456 = ~n46452 & n46455;
  assign n46457 = ~n46451 & n46456;
  assign n46458 = pi5  & ~n46457;
  assign n46459 = ~n46457 & ~n46458;
  assign n46460 = ~pi5  & ~n46457;
  assign n46461 = pi5  & ~n46458;
  assign n46462 = pi5  & n46457;
  assign n46463 = ~n59449 & ~n59450;
  assign n46464 = ~n46352 & ~n46360;
  assign n46465 = ~n46328 & ~n46337;
  assign n46466 = n18846 & ~n59050;
  assign n46467 = n19541 & n39440;
  assign n46468 = n55247 & n39549;
  assign n46469 = n19509 & n39546;
  assign n46470 = ~n46468 & ~n46469;
  assign n46471 = ~n46467 & n46470;
  assign n46472 = ~n46466 & n46471;
  assign n46473 = pi11  & ~n46472;
  assign n46474 = ~n46472 & ~n46473;
  assign n46475 = ~pi11  & ~n46472;
  assign n46476 = pi11  & ~n46473;
  assign n46477 = pi11  & n46472;
  assign n46478 = ~n59451 & ~n59452;
  assign n46479 = ~n46314 & ~n46322;
  assign n46480 = ~n46292 & ~n46299;
  assign n46481 = n16079 & ~n58493;
  assign n46482 = n16696 & n39561;
  assign n46483 = n54886 & n39567;
  assign n46484 = n16676 & n39564;
  assign n46485 = ~n46483 & ~n46484;
  assign n46486 = ~n46482 & n46485;
  assign n46487 = ~n46481 & n46486;
  assign n46488 = pi17  & ~n46487;
  assign n46489 = ~n46487 & ~n46488;
  assign n46490 = ~pi17  & ~n46487;
  assign n46491 = pi17  & ~n46488;
  assign n46492 = pi17  & n46487;
  assign n46493 = ~n59453 & ~n59454;
  assign n46494 = ~n46276 & ~n46284;
  assign n46495 = ~n46252 & ~n46261;
  assign n46496 = n90 & ~n58657;
  assign n46497 = n14236 & n39579;
  assign n46498 = n54667 & n39585;
  assign n46499 = n14210 & n39582;
  assign n46500 = ~n46498 & ~n46499;
  assign n46501 = ~n46497 & n46500;
  assign n46502 = ~n46496 & n46501;
  assign n46503 = pi23  & ~n46502;
  assign n46504 = ~n46502 & ~n46503;
  assign n46505 = ~pi23  & ~n46502;
  assign n46506 = pi23  & ~n46503;
  assign n46507 = pi23  & n46502;
  assign n46508 = ~n59455 & ~n59456;
  assign n46509 = ~n46238 & ~n46246;
  assign n46510 = ~n46219 & ~n46222;
  assign n46511 = n11279 & n40247;
  assign n46512 = n12584 & n39597;
  assign n46513 = n54410 & n39603;
  assign n46514 = n11267 & n39600;
  assign n46515 = ~n46513 & ~n46514;
  assign n46516 = ~n46512 & n46515;
  assign n46517 = ~n11279 & n46516;
  assign n46518 = ~n40247 & n46516;
  assign n46519 = ~n46517 & ~n46518;
  assign n46520 = ~n46511 & n46516;
  assign n46521 = pi29  & ~n59457;
  assign n46522 = ~pi29  & n59457;
  assign n46523 = ~n46521 & ~n46522;
  assign n46524 = ~n46205 & ~n46213;
  assign n46525 = n1273 & n1391;
  assign n46526 = n3536 & n9155;
  assign n46527 = n46525 & n46526;
  assign n46528 = ~n166 & ~n663;
  assign n46529 = ~n357 & n46528;
  assign n46530 = n561 & n1647;
  assign n46531 = ~n166 & ~n1646;
  assign n46532 = ~n956 & n46531;
  assign n46533 = ~n357 & ~n663;
  assign n46534 = n561 & n46533;
  assign n46535 = n46532 & n46534;
  assign n46536 = ~n357 & ~n1646;
  assign n46537 = ~n166 & n46536;
  assign n46538 = ~n663 & ~n956;
  assign n46539 = n561 & n46538;
  assign n46540 = n46537 & n46539;
  assign n46541 = n46529 & n46530;
  assign n46542 = n1273 & n3536;
  assign n46543 = n561 & n9155;
  assign n46544 = n46542 & n46543;
  assign n46545 = ~n956 & n46528;
  assign n46546 = n1391 & n46536;
  assign n46547 = n46545 & n46546;
  assign n46548 = n46544 & n46547;
  assign n46549 = n46527 & n59458;
  assign n46550 = n54102 & n18271;
  assign n46551 = n59459 & n46550;
  assign n46552 = n4916 & n27277;
  assign n46553 = n56750 & n46552;
  assign n46554 = n54506 & n46553;
  assign n46555 = n46551 & n46554;
  assign n46556 = n54058 & n46555;
  assign n46557 = n27277 & n56750;
  assign n46558 = n18271 & n46557;
  assign n46559 = n9155 & n46558;
  assign n46560 = n4916 & n46559;
  assign n46561 = n54500 & n46560;
  assign n46562 = n54506 & n46561;
  assign n46563 = n54058 & n46562;
  assign n46564 = n1273 & n46563;
  assign n46565 = n54102 & n46564;
  assign n46566 = n1391 & n46565;
  assign n46567 = n561 & n46566;
  assign n46568 = n3536 & n46567;
  assign n46569 = ~n166 & n46568;
  assign n46570 = ~n663 & n46569;
  assign n46571 = ~n956 & n46570;
  assign n46572 = ~n1646 & n46571;
  assign n46573 = ~n357 & n46572;
  assign n46574 = n54500 & n46556;
  assign n46575 = n1576 & n40183;
  assign n46576 = n11215 & n39606;
  assign n46577 = n10564 & n39609;
  assign n46578 = n54403 & n39612;
  assign n46579 = ~n46577 & ~n46578;
  assign n46580 = ~n46576 & n46579;
  assign n46581 = ~n46575 & ~n46578;
  assign n46582 = ~n46577 & n46581;
  assign n46583 = ~n46576 & n46582;
  assign n46584 = ~n46575 & n46580;
  assign n46585 = ~n59460 & ~n59461;
  assign n46586 = n59460 & n59461;
  assign n46587 = ~n59460 & ~n46585;
  assign n46588 = ~n59460 & n59461;
  assign n46589 = ~n59461 & ~n46585;
  assign n46590 = n59460 & ~n59461;
  assign n46591 = ~n59462 & ~n59463;
  assign n46592 = ~n46585 & ~n46586;
  assign n46593 = ~n46524 & ~n59464;
  assign n46594 = n46524 & n59464;
  assign n46595 = ~n46524 & ~n46593;
  assign n46596 = ~n59464 & ~n46593;
  assign n46597 = ~n46595 & ~n46596;
  assign n46598 = ~n46593 & ~n46594;
  assign n46599 = ~n46523 & ~n59465;
  assign n46600 = n46523 & n59465;
  assign n46601 = ~n46599 & ~n46600;
  assign n46602 = ~n46510 & n46601;
  assign n46603 = n46510 & ~n46601;
  assign n46604 = ~n46602 & ~n46603;
  assign n46605 = n123 & ~n58585;
  assign n46606 = n128 & n39588;
  assign n46607 = n53444 & n39594;
  assign n46608 = n127 & n39591;
  assign n46609 = ~n46607 & ~n46608;
  assign n46610 = ~n46606 & n46609;
  assign n46611 = ~n123 & n46610;
  assign n46612 = n58585 & n46610;
  assign n46613 = ~n46611 & ~n46612;
  assign n46614 = ~n46605 & n46610;
  assign n46615 = pi26  & ~n59466;
  assign n46616 = ~pi26  & n59466;
  assign n46617 = ~n46615 & ~n46616;
  assign n46618 = n46604 & ~n46617;
  assign n46619 = ~n46604 & n46617;
  assign n46620 = n46604 & ~n46618;
  assign n46621 = n46604 & n46617;
  assign n46622 = ~n46617 & ~n46618;
  assign n46623 = ~n46604 & ~n46617;
  assign n46624 = ~n59467 & ~n59468;
  assign n46625 = ~n46618 & ~n46619;
  assign n46626 = ~n46509 & ~n59469;
  assign n46627 = n46509 & n59469;
  assign n46628 = ~n46509 & ~n46626;
  assign n46629 = ~n59469 & ~n46626;
  assign n46630 = ~n46628 & ~n46629;
  assign n46631 = ~n46626 & ~n46627;
  assign n46632 = ~n46508 & ~n59470;
  assign n46633 = n46508 & n59470;
  assign n46634 = ~n46508 & ~n46632;
  assign n46635 = ~n46508 & n59470;
  assign n46636 = ~n59470 & ~n46632;
  assign n46637 = n46508 & ~n59470;
  assign n46638 = ~n59471 & ~n59472;
  assign n46639 = ~n46632 & ~n46633;
  assign n46640 = n46495 & n59473;
  assign n46641 = ~n46495 & ~n59473;
  assign n46642 = ~n46640 & ~n46641;
  assign n46643 = n14413 & ~n58759;
  assign n46644 = n15921 & n39570;
  assign n46645 = n54719 & n39576;
  assign n46646 = n15901 & n39573;
  assign n46647 = ~n46645 & ~n46646;
  assign n46648 = ~n46644 & n46647;
  assign n46649 = ~n14413 & n46648;
  assign n46650 = n58759 & n46648;
  assign n46651 = ~n46649 & ~n46650;
  assign n46652 = ~n46643 & n46648;
  assign n46653 = pi20  & ~n59474;
  assign n46654 = ~pi20  & n59474;
  assign n46655 = ~n46653 & ~n46654;
  assign n46656 = n46642 & ~n46655;
  assign n46657 = ~n46642 & n46655;
  assign n46658 = n46642 & ~n46656;
  assign n46659 = n46642 & n46655;
  assign n46660 = ~n46655 & ~n46656;
  assign n46661 = ~n46642 & ~n46655;
  assign n46662 = ~n59475 & ~n59476;
  assign n46663 = ~n46656 & ~n46657;
  assign n46664 = ~n46494 & ~n59477;
  assign n46665 = n46494 & n59477;
  assign n46666 = ~n46494 & ~n46664;
  assign n46667 = ~n46494 & n59477;
  assign n46668 = ~n59477 & ~n46664;
  assign n46669 = n46494 & ~n59477;
  assign n46670 = ~n59478 & ~n59479;
  assign n46671 = ~n46664 & ~n46665;
  assign n46672 = ~n46493 & ~n59480;
  assign n46673 = n46493 & n59480;
  assign n46674 = ~n46493 & ~n46672;
  assign n46675 = ~n59480 & ~n46672;
  assign n46676 = ~n46674 & ~n46675;
  assign n46677 = ~n46672 & ~n46673;
  assign n46678 = n46480 & n59481;
  assign n46679 = ~n46480 & ~n59481;
  assign n46680 = ~n46678 & ~n46679;
  assign n46681 = n17265 & ~n58891;
  assign n46682 = n18588 & n39552;
  assign n46683 = n55041 & n39558;
  assign n46684 = n18556 & n39555;
  assign n46685 = ~n46683 & ~n46684;
  assign n46686 = ~n46682 & n46685;
  assign n46687 = ~n17265 & n46686;
  assign n46688 = n58891 & n46686;
  assign n46689 = ~n46687 & ~n46688;
  assign n46690 = ~n46681 & n46686;
  assign n46691 = pi14  & ~n59482;
  assign n46692 = ~pi14  & n59482;
  assign n46693 = ~n46691 & ~n46692;
  assign n46694 = n46680 & ~n46693;
  assign n46695 = ~n46680 & n46693;
  assign n46696 = n46680 & ~n46694;
  assign n46697 = n46680 & n46693;
  assign n46698 = ~n46693 & ~n46694;
  assign n46699 = ~n46680 & ~n46693;
  assign n46700 = ~n59483 & ~n59484;
  assign n46701 = ~n46694 & ~n46695;
  assign n46702 = ~n46479 & ~n59485;
  assign n46703 = n46479 & n59485;
  assign n46704 = ~n46479 & ~n46702;
  assign n46705 = ~n59485 & ~n46702;
  assign n46706 = ~n46704 & ~n46705;
  assign n46707 = ~n46702 & ~n46703;
  assign n46708 = ~n46478 & ~n59486;
  assign n46709 = n46478 & n59486;
  assign n46710 = ~n46478 & ~n46708;
  assign n46711 = ~n46478 & n59486;
  assign n46712 = ~n59486 & ~n46708;
  assign n46713 = n46478 & ~n59486;
  assign n46714 = ~n59487 & ~n59488;
  assign n46715 = ~n46708 & ~n46709;
  assign n46716 = n46465 & n59489;
  assign n46717 = ~n46465 & ~n59489;
  assign n46718 = ~n46716 & ~n46717;
  assign n46719 = n20085 & ~n59184;
  assign n46720 = n21269 & n44327;
  assign n46721 = n55472 & n39543;
  assign n46722 = n21237 & n39937;
  assign n46723 = ~n46721 & ~n46722;
  assign n46724 = ~n46720 & n46723;
  assign n46725 = ~n20085 & n46724;
  assign n46726 = n59184 & n46724;
  assign n46727 = ~n46725 & ~n46726;
  assign n46728 = ~n46719 & n46724;
  assign n46729 = pi8  & ~n59490;
  assign n46730 = ~pi8  & n59490;
  assign n46731 = ~n46729 & ~n46730;
  assign n46732 = n46718 & ~n46731;
  assign n46733 = ~n46718 & n46731;
  assign n46734 = n46718 & ~n46732;
  assign n46735 = n46718 & n46731;
  assign n46736 = ~n46731 & ~n46732;
  assign n46737 = ~n46718 & ~n46731;
  assign n46738 = ~n59491 & ~n59492;
  assign n46739 = ~n46732 & ~n46733;
  assign n46740 = ~n46464 & ~n59493;
  assign n46741 = n46464 & n59493;
  assign n46742 = ~n46464 & ~n46740;
  assign n46743 = ~n46464 & n59493;
  assign n46744 = ~n59493 & ~n46740;
  assign n46745 = n46464 & ~n59493;
  assign n46746 = ~n59494 & ~n59495;
  assign n46747 = ~n46740 & ~n46741;
  assign n46748 = ~n46463 & ~n59496;
  assign n46749 = n46463 & n59496;
  assign n46750 = ~n46463 & ~n46748;
  assign n46751 = ~n59496 & ~n46748;
  assign n46752 = ~n46750 & ~n46751;
  assign n46753 = ~n46748 & ~n46749;
  assign n46754 = n46450 & n59497;
  assign n46755 = ~n46450 & ~n59497;
  assign n46756 = ~n46754 & ~n46755;
  assign n46757 = ~n46422 & ~n46424;
  assign n46758 = ~n46415 & ~n46418;
  assign n46759 = ~n46401 & ~n46409;
  assign n46760 = ~n53622 & n46379;
  assign n46761 = n46000 & n46760;
  assign n46762 = ~n46000 & ~n46760;
  assign n46763 = ~n46761 & ~n46762;
  assign n46764 = ~n10564 & ~n54403;
  assign n46765 = ~n11215 & ~n54403;
  assign n46766 = ~n10564 & n46765;
  assign n46767 = ~n10564 & ~n11215;
  assign n46768 = ~n54403 & n46767;
  assign n46769 = ~n11215 & n46764;
  assign n46770 = ~n1576 & n59498;
  assign n46771 = ~pi31  & n266;
  assign n46772 = n46763 & ~n59499;
  assign n46773 = ~n46763 & n59499;
  assign n46774 = n46763 & ~n46772;
  assign n46775 = n46763 & n59499;
  assign n46776 = ~n59499 & ~n46772;
  assign n46777 = ~n46763 & ~n59499;
  assign n46778 = ~n59500 & ~n59501;
  assign n46779 = ~n46772 & ~n46773;
  assign n46780 = ~n46391 & ~n59502;
  assign n46781 = n46391 & n59502;
  assign n46782 = ~n46780 & ~n46781;
  assign n46783 = ~n46759 & n46782;
  assign n46784 = n46759 & ~n46782;
  assign n46785 = ~n46783 & ~n46784;
  assign n46786 = ~n46758 & n46785;
  assign n46787 = n46758 & ~n46785;
  assign n46788 = ~n46786 & ~n46787;
  assign n46789 = ~n46772 & ~n46780;
  assign n46790 = n46379 & ~n46761;
  assign n46791 = ~n53622 & n46790;
  assign n46792 = ~n59499 & ~n46791;
  assign n46793 = n46789 & ~n46792;
  assign n46794 = ~n46789 & n46792;
  assign n46795 = ~n46793 & ~n46794;
  assign n46796 = ~n46783 & ~n46786;
  assign n46797 = ~n46795 & n46796;
  assign n46798 = n46795 & ~n46796;
  assign n46799 = ~n46797 & ~n46798;
  assign n46800 = ~n46420 & ~n46788;
  assign n46801 = n46420 & n46788;
  assign n46802 = ~n59503 & ~n46801;
  assign n46803 = ~n46757 & n46802;
  assign n46804 = n46757 & ~n46802;
  assign n46805 = ~n46803 & ~n46804;
  assign n46806 = n24338 & n46805;
  assign n46807 = n25287 & n46788;
  assign n46808 = n24337 & n46009;
  assign n46809 = n25272 & n46420;
  assign n46810 = ~n46808 & ~n46809;
  assign n46811 = ~n46807 & n46810;
  assign n46812 = ~n24338 & n46811;
  assign n46813 = ~n46805 & n46811;
  assign n46814 = ~n46812 & ~n46813;
  assign n46815 = ~n46806 & n46811;
  assign n46816 = pi2  & ~n59504;
  assign n46817 = ~pi2  & n59504;
  assign n46818 = ~n46816 & ~n46817;
  assign n46819 = n46756 & ~n46818;
  assign n46820 = ~n46756 & n46818;
  assign n46821 = ~n46819 & ~n46820;
  assign n46822 = ~n46449 & n46821;
  assign n46823 = n46449 & ~n46821;
  assign n46824 = ~n46822 & ~n46823;
  assign n46825 = n46446 & n46824;
  assign n46826 = ~n46446 & ~n46824;
  assign po2  = ~n46825 & ~n46826;
  assign n46828 = ~n46819 & ~n46822;
  assign n46829 = ~n46748 & ~n46755;
  assign n46830 = n77 & ~n59386;
  assign n46831 = n24302 & n46009;
  assign n46832 = n21969 & n44871;
  assign n46833 = n23459 & n44952;
  assign n46834 = ~n46832 & ~n46833;
  assign n46835 = ~n46831 & n46834;
  assign n46836 = ~n46830 & n46835;
  assign n46837 = pi5  & ~n46836;
  assign n46838 = ~n46836 & ~n46837;
  assign n46839 = ~pi5  & ~n46836;
  assign n46840 = pi5  & ~n46837;
  assign n46841 = pi5  & n46836;
  assign n46842 = ~n59505 & ~n59506;
  assign n46843 = ~n46732 & ~n46740;
  assign n46844 = ~n46708 & ~n46717;
  assign n46845 = n18846 & ~n59044;
  assign n46846 = n19541 & n39543;
  assign n46847 = n55247 & n39546;
  assign n46848 = n19509 & n39440;
  assign n46849 = ~n46847 & ~n46848;
  assign n46850 = ~n46846 & n46849;
  assign n46851 = ~n46845 & n46850;
  assign n46852 = pi11  & ~n46851;
  assign n46853 = ~n46851 & ~n46852;
  assign n46854 = ~pi11  & ~n46851;
  assign n46855 = pi11  & ~n46852;
  assign n46856 = pi11  & n46851;
  assign n46857 = ~n59507 & ~n59508;
  assign n46858 = ~n46694 & ~n46702;
  assign n46859 = ~n46672 & ~n46679;
  assign n46860 = n16079 & ~n58849;
  assign n46861 = n16696 & n39558;
  assign n46862 = n54886 & n39564;
  assign n46863 = n16676 & n39561;
  assign n46864 = ~n46862 & ~n46863;
  assign n46865 = ~n46861 & n46864;
  assign n46866 = ~n46860 & n46865;
  assign n46867 = pi17  & ~n46866;
  assign n46868 = ~n46866 & ~n46867;
  assign n46869 = ~pi17  & ~n46866;
  assign n46870 = pi17  & ~n46867;
  assign n46871 = pi17  & n46866;
  assign n46872 = ~n59509 & ~n59510;
  assign n46873 = ~n46656 & ~n46664;
  assign n46874 = ~n46632 & ~n46641;
  assign n46875 = n90 & ~n58653;
  assign n46876 = n14236 & n39576;
  assign n46877 = n54667 & n39582;
  assign n46878 = n14210 & n39579;
  assign n46879 = ~n46877 & ~n46878;
  assign n46880 = ~n46876 & n46879;
  assign n46881 = ~n46875 & n46880;
  assign n46882 = pi23  & ~n46881;
  assign n46883 = ~n46881 & ~n46882;
  assign n46884 = ~pi23  & ~n46881;
  assign n46885 = pi23  & ~n46882;
  assign n46886 = pi23  & n46881;
  assign n46887 = ~n59511 & ~n59512;
  assign n46888 = ~n46618 & ~n46626;
  assign n46889 = ~n46599 & ~n46602;
  assign n46890 = n11279 & n40476;
  assign n46891 = n12584 & n39594;
  assign n46892 = n54410 & n39600;
  assign n46893 = n11267 & n39597;
  assign n46894 = ~n46892 & ~n46893;
  assign n46895 = ~n46891 & n46894;
  assign n46896 = ~n11279 & n46895;
  assign n46897 = ~n40476 & n46895;
  assign n46898 = ~n46896 & ~n46897;
  assign n46899 = ~n46890 & n46895;
  assign n46900 = pi29  & ~n59513;
  assign n46901 = ~pi29  & n59513;
  assign n46902 = ~n46900 & ~n46901;
  assign n46903 = ~n46585 & ~n46593;
  assign n46904 = ~n627 & ~n975;
  assign n46905 = n1128 & n46904;
  assign n46906 = n54086 & n46905;
  assign n46907 = n54090 & n54731;
  assign n46908 = n46906 & n46907;
  assign n46909 = n309 & n3389;
  assign n46910 = n903 & n3389;
  assign n46911 = n309 & n46910;
  assign n46912 = n903 & n46909;
  assign n46913 = n3217 & n4584;
  assign n46914 = n9155 & n46913;
  assign n46915 = n59514 & n46914;
  assign n46916 = n3217 & n46904;
  assign n46917 = n54086 & n46916;
  assign n46918 = n46907 & n46917;
  assign n46919 = n1128 & n4584;
  assign n46920 = n9155 & n46919;
  assign n46921 = n59514 & n46920;
  assign n46922 = n46918 & n46921;
  assign n46923 = n4584 & n46904;
  assign n46924 = n54090 & n46923;
  assign n46925 = n54086 & n54731;
  assign n46926 = n46924 & n46925;
  assign n46927 = n1128 & n3217;
  assign n46928 = n9155 & n46927;
  assign n46929 = n59514 & n46928;
  assign n46930 = n46926 & n46929;
  assign n46931 = n46908 & n46915;
  assign n46932 = n57005 & n59515;
  assign n46933 = n54196 & n46932;
  assign n46934 = n54448 & n55151;
  assign n46935 = n54086 & n54090;
  assign n46936 = n59514 & n46935;
  assign n46937 = n9155 & n46936;
  assign n46938 = n54731 & n46937;
  assign n46939 = n57005 & n46938;
  assign n46940 = n55151 & n46939;
  assign n46941 = n54448 & n46940;
  assign n46942 = n54196 & n46941;
  assign n46943 = n4584 & n46942;
  assign n46944 = n3217 & n46943;
  assign n46945 = n1128 & n46944;
  assign n46946 = ~n975 & n46945;
  assign n46947 = ~n627 & n46946;
  assign n46948 = n46933 & n46934;
  assign n46949 = n1576 & n40286;
  assign n46950 = n11215 & n39603;
  assign n46951 = n10564 & n39606;
  assign n46952 = n54403 & n39609;
  assign n46953 = ~n46951 & ~n46952;
  assign n46954 = ~n46950 & n46953;
  assign n46955 = ~n46949 & ~n46952;
  assign n46956 = ~n46951 & n46955;
  assign n46957 = ~n46950 & n46956;
  assign n46958 = ~n46949 & n46954;
  assign n46959 = ~n59516 & ~n59517;
  assign n46960 = n59516 & n59517;
  assign n46961 = ~n59516 & ~n46959;
  assign n46962 = ~n59516 & n59517;
  assign n46963 = ~n59517 & ~n46959;
  assign n46964 = n59516 & ~n59517;
  assign n46965 = ~n59518 & ~n59519;
  assign n46966 = ~n46959 & ~n46960;
  assign n46967 = ~n46903 & ~n59520;
  assign n46968 = n46903 & n59520;
  assign n46969 = ~n46903 & ~n46967;
  assign n46970 = ~n59520 & ~n46967;
  assign n46971 = ~n46969 & ~n46970;
  assign n46972 = ~n46967 & ~n46968;
  assign n46973 = ~n46902 & ~n59521;
  assign n46974 = n46902 & n59521;
  assign n46975 = ~n46973 & ~n46974;
  assign n46976 = ~n46889 & n46975;
  assign n46977 = n46889 & ~n46975;
  assign n46978 = ~n46976 & ~n46977;
  assign n46979 = n123 & ~n58583;
  assign n46980 = n128 & n39585;
  assign n46981 = n53444 & n39591;
  assign n46982 = n127 & n39588;
  assign n46983 = ~n46981 & ~n46982;
  assign n46984 = ~n46980 & n46983;
  assign n46985 = ~n123 & n46984;
  assign n46986 = n58583 & n46984;
  assign n46987 = ~n46985 & ~n46986;
  assign n46988 = ~n46979 & n46984;
  assign n46989 = pi26  & ~n59522;
  assign n46990 = ~pi26  & n59522;
  assign n46991 = ~n46989 & ~n46990;
  assign n46992 = n46978 & ~n46991;
  assign n46993 = ~n46978 & n46991;
  assign n46994 = n46978 & ~n46992;
  assign n46995 = n46978 & n46991;
  assign n46996 = ~n46991 & ~n46992;
  assign n46997 = ~n46978 & ~n46991;
  assign n46998 = ~n59523 & ~n59524;
  assign n46999 = ~n46992 & ~n46993;
  assign n47000 = ~n46888 & ~n59525;
  assign n47001 = n46888 & n59525;
  assign n47002 = ~n46888 & ~n47000;
  assign n47003 = ~n59525 & ~n47000;
  assign n47004 = ~n47002 & ~n47003;
  assign n47005 = ~n47000 & ~n47001;
  assign n47006 = ~n46887 & ~n59526;
  assign n47007 = n46887 & n59526;
  assign n47008 = ~n46887 & ~n47006;
  assign n47009 = ~n46887 & n59526;
  assign n47010 = ~n59526 & ~n47006;
  assign n47011 = n46887 & ~n59526;
  assign n47012 = ~n59527 & ~n59528;
  assign n47013 = ~n47006 & ~n47007;
  assign n47014 = n46874 & n59529;
  assign n47015 = ~n46874 & ~n59529;
  assign n47016 = ~n47014 & ~n47015;
  assign n47017 = n14413 & ~n58766;
  assign n47018 = n15921 & n39567;
  assign n47019 = n54719 & n39573;
  assign n47020 = n15901 & n39570;
  assign n47021 = ~n47019 & ~n47020;
  assign n47022 = ~n47018 & n47021;
  assign n47023 = ~n14413 & n47022;
  assign n47024 = n58766 & n47022;
  assign n47025 = ~n47023 & ~n47024;
  assign n47026 = ~n47017 & n47022;
  assign n47027 = pi20  & ~n59530;
  assign n47028 = ~pi20  & n59530;
  assign n47029 = ~n47027 & ~n47028;
  assign n47030 = n47016 & ~n47029;
  assign n47031 = ~n47016 & n47029;
  assign n47032 = n47016 & ~n47030;
  assign n47033 = n47016 & n47029;
  assign n47034 = ~n47029 & ~n47030;
  assign n47035 = ~n47016 & ~n47029;
  assign n47036 = ~n59531 & ~n59532;
  assign n47037 = ~n47030 & ~n47031;
  assign n47038 = ~n46873 & ~n59533;
  assign n47039 = n46873 & n59533;
  assign n47040 = ~n46873 & ~n47038;
  assign n47041 = ~n46873 & n59533;
  assign n47042 = ~n59533 & ~n47038;
  assign n47043 = n46873 & ~n59533;
  assign n47044 = ~n59534 & ~n59535;
  assign n47045 = ~n47038 & ~n47039;
  assign n47046 = ~n46872 & ~n59536;
  assign n47047 = n46872 & n59536;
  assign n47048 = ~n46872 & ~n47046;
  assign n47049 = ~n59536 & ~n47046;
  assign n47050 = ~n47048 & ~n47049;
  assign n47051 = ~n47046 & ~n47047;
  assign n47052 = n46859 & n59537;
  assign n47053 = ~n46859 & ~n59537;
  assign n47054 = ~n47052 & ~n47053;
  assign n47055 = n17265 & ~n58889;
  assign n47056 = n18588 & n39549;
  assign n47057 = n55041 & n39555;
  assign n47058 = n18556 & n39552;
  assign n47059 = ~n47057 & ~n47058;
  assign n47060 = ~n47056 & n47059;
  assign n47061 = ~n17265 & n47060;
  assign n47062 = n58889 & n47060;
  assign n47063 = ~n47061 & ~n47062;
  assign n47064 = ~n47055 & n47060;
  assign n47065 = pi14  & ~n59538;
  assign n47066 = ~pi14  & n59538;
  assign n47067 = ~n47065 & ~n47066;
  assign n47068 = n47054 & ~n47067;
  assign n47069 = ~n47054 & n47067;
  assign n47070 = n47054 & ~n47068;
  assign n47071 = n47054 & n47067;
  assign n47072 = ~n47067 & ~n47068;
  assign n47073 = ~n47054 & ~n47067;
  assign n47074 = ~n59539 & ~n59540;
  assign n47075 = ~n47068 & ~n47069;
  assign n47076 = ~n46858 & ~n59541;
  assign n47077 = n46858 & n59541;
  assign n47078 = ~n46858 & ~n47076;
  assign n47079 = ~n59541 & ~n47076;
  assign n47080 = ~n47078 & ~n47079;
  assign n47081 = ~n47076 & ~n47077;
  assign n47082 = ~n46857 & ~n59542;
  assign n47083 = n46857 & n59542;
  assign n47084 = ~n46857 & ~n47082;
  assign n47085 = ~n46857 & n59542;
  assign n47086 = ~n59542 & ~n47082;
  assign n47087 = n46857 & ~n59542;
  assign n47088 = ~n59543 & ~n59544;
  assign n47089 = ~n47082 & ~n47083;
  assign n47090 = n46844 & n59545;
  assign n47091 = ~n46844 & ~n59545;
  assign n47092 = ~n47090 & ~n47091;
  assign n47093 = n20085 & ~n59282;
  assign n47094 = n21269 & n44775;
  assign n47095 = n55472 & n39937;
  assign n47096 = n21237 & n44327;
  assign n47097 = ~n47095 & ~n47096;
  assign n47098 = ~n47094 & n47097;
  assign n47099 = ~n20085 & n47098;
  assign n47100 = n59282 & n47098;
  assign n47101 = ~n47099 & ~n47100;
  assign n47102 = ~n47093 & n47098;
  assign n47103 = pi8  & ~n59546;
  assign n47104 = ~pi8  & n59546;
  assign n47105 = ~n47103 & ~n47104;
  assign n47106 = n47092 & ~n47105;
  assign n47107 = ~n47092 & n47105;
  assign n47108 = n47092 & ~n47106;
  assign n47109 = n47092 & n47105;
  assign n47110 = ~n47105 & ~n47106;
  assign n47111 = ~n47092 & ~n47105;
  assign n47112 = ~n59547 & ~n59548;
  assign n47113 = ~n47106 & ~n47107;
  assign n47114 = ~n46843 & ~n59549;
  assign n47115 = n46843 & n59549;
  assign n47116 = ~n46843 & ~n47114;
  assign n47117 = ~n46843 & n59549;
  assign n47118 = ~n59549 & ~n47114;
  assign n47119 = n46843 & ~n59549;
  assign n47120 = ~n59550 & ~n59551;
  assign n47121 = ~n47114 & ~n47115;
  assign n47122 = ~n46842 & ~n59552;
  assign n47123 = n46842 & n59552;
  assign n47124 = ~n46842 & ~n47122;
  assign n47125 = ~n59552 & ~n47122;
  assign n47126 = ~n47124 & ~n47125;
  assign n47127 = ~n47122 & ~n47123;
  assign n47128 = n46829 & n59553;
  assign n47129 = ~n46829 & ~n59553;
  assign n47130 = ~n47128 & ~n47129;
  assign n47131 = ~n46801 & ~n46803;
  assign n47132 = ~n46788 & ~n59503;
  assign n47133 = ~n47131 & ~n47132;
  assign n47134 = n47131 & n47132;
  assign n47135 = ~n47131 & ~n47133;
  assign n47136 = ~n47132 & ~n47133;
  assign n47137 = ~n47135 & ~n47136;
  assign n47138 = ~n47133 & ~n47134;
  assign n47139 = n24338 & ~n59554;
  assign n47140 = n25287 & n59503;
  assign n47141 = n24337 & n46420;
  assign n47142 = n25272 & n46788;
  assign n47143 = ~n47141 & ~n47142;
  assign n47144 = ~n47140 & n47143;
  assign n47145 = ~n24338 & n47144;
  assign n47146 = n59554 & n47144;
  assign n47147 = ~n47145 & ~n47146;
  assign n47148 = ~n47139 & n47144;
  assign n47149 = pi2  & ~n59555;
  assign n47150 = ~pi2  & n59555;
  assign n47151 = ~n47149 & ~n47150;
  assign n47152 = n47130 & ~n47151;
  assign n47153 = ~n47130 & n47151;
  assign n47154 = ~n47152 & ~n47153;
  assign n47155 = ~n46828 & n47154;
  assign n47156 = n46828 & ~n47154;
  assign n47157 = ~n47155 & ~n47156;
  assign n47158 = n46825 & n47157;
  assign n47159 = ~n46825 & ~n47157;
  assign po3  = ~n47158 & ~n47159;
  assign n47161 = ~n47152 & ~n47155;
  assign n47162 = ~n47122 & ~n47129;
  assign n47163 = n77 & n46426;
  assign n47164 = n24302 & n46420;
  assign n47165 = n21969 & n44952;
  assign n47166 = n23459 & n46009;
  assign n47167 = ~n47165 & ~n47166;
  assign n47168 = ~n47164 & n47167;
  assign n47169 = ~n47163 & n47168;
  assign n47170 = pi5  & ~n47169;
  assign n47171 = ~n47169 & ~n47170;
  assign n47172 = ~pi5  & ~n47169;
  assign n47173 = pi5  & ~n47170;
  assign n47174 = pi5  & n47169;
  assign n47175 = ~n59556 & ~n59557;
  assign n47176 = ~n47106 & ~n47114;
  assign n47177 = ~n47082 & ~n47091;
  assign n47178 = n18846 & n39943;
  assign n47179 = n19541 & n39937;
  assign n47180 = n55247 & n39440;
  assign n47181 = n19509 & n39543;
  assign n47182 = ~n47180 & ~n47181;
  assign n47183 = ~n47179 & n47182;
  assign n47184 = ~n47178 & n47183;
  assign n47185 = pi11  & ~n47184;
  assign n47186 = ~n47184 & ~n47185;
  assign n47187 = ~pi11  & ~n47184;
  assign n47188 = pi11  & ~n47185;
  assign n47189 = pi11  & n47184;
  assign n47190 = ~n59558 & ~n59559;
  assign n47191 = ~n47068 & ~n47076;
  assign n47192 = ~n47046 & ~n47053;
  assign n47193 = n16079 & n42574;
  assign n47194 = n16696 & n39555;
  assign n47195 = n54886 & n39561;
  assign n47196 = n16676 & n39558;
  assign n47197 = ~n47195 & ~n47196;
  assign n47198 = ~n47194 & n47197;
  assign n47199 = ~n47193 & n47198;
  assign n47200 = pi17  & ~n47199;
  assign n47201 = ~n47199 & ~n47200;
  assign n47202 = ~pi17  & ~n47199;
  assign n47203 = pi17  & ~n47200;
  assign n47204 = pi17  & n47199;
  assign n47205 = ~n59560 & ~n59561;
  assign n47206 = ~n47030 & ~n47038;
  assign n47207 = ~n47006 & ~n47015;
  assign n47208 = n90 & n39976;
  assign n47209 = n14236 & n39573;
  assign n47210 = n54667 & n39579;
  assign n47211 = n14210 & n39576;
  assign n47212 = ~n47210 & ~n47211;
  assign n47213 = ~n47209 & n47212;
  assign n47214 = ~n47208 & n47213;
  assign n47215 = pi23  & ~n47214;
  assign n47216 = ~n47214 & ~n47215;
  assign n47217 = ~pi23  & ~n47214;
  assign n47218 = pi23  & ~n47215;
  assign n47219 = pi23  & n47214;
  assign n47220 = ~n59562 & ~n59563;
  assign n47221 = ~n46992 & ~n47000;
  assign n47222 = ~n46973 & ~n46976;
  assign n47223 = n11279 & n40616;
  assign n47224 = n12584 & n39591;
  assign n47225 = n54410 & n39597;
  assign n47226 = n11267 & n39594;
  assign n47227 = ~n47225 & ~n47226;
  assign n47228 = ~n47224 & n47227;
  assign n47229 = ~n11279 & n47228;
  assign n47230 = ~n40616 & n47228;
  assign n47231 = ~n47229 & ~n47230;
  assign n47232 = ~n47223 & n47228;
  assign n47233 = pi29  & ~n59564;
  assign n47234 = ~pi29  & n59564;
  assign n47235 = ~n47233 & ~n47234;
  assign n47236 = ~n46959 & ~n46967;
  assign n47237 = n7307 & n8268;
  assign n47238 = n3560 & n3672;
  assign n47239 = n47237 & n47238;
  assign n47240 = n2814 & n4261;
  assign n47241 = n406 & n648;
  assign n47242 = n47240 & n47241;
  assign n47243 = n47239 & n47242;
  assign n47244 = n54158 & n47243;
  assign n47245 = n7144 & n8267;
  assign n47246 = n16874 & n28019;
  assign n47247 = n47245 & n47246;
  assign n47248 = ~n221 & ~n1065;
  assign n47249 = n2037 & n47248;
  assign n47250 = n3476 & n4021;
  assign n47251 = n47249 & n47250;
  assign n47252 = n2037 & n16874;
  assign n47253 = n28019 & n47252;
  assign n47254 = ~n212 & ~n221;
  assign n47255 = ~n1065 & n47254;
  assign n47256 = n12328 & n47255;
  assign n47257 = n46142 & n47256;
  assign n47258 = n47253 & n47257;
  assign n47259 = n4021 & n7144;
  assign n47260 = n3476 & n8267;
  assign n47261 = n4021 & n8267;
  assign n47262 = n3476 & n47261;
  assign n47263 = n7144 & n47262;
  assign n47264 = n47259 & n47260;
  assign n47265 = ~n1065 & n59566;
  assign n47266 = ~n256 & n47265;
  assign n47267 = ~n221 & n47266;
  assign n47268 = ~n402 & n47267;
  assign n47269 = ~n663 & n47268;
  assign n47270 = ~n830 & n47269;
  assign n47271 = ~n1644 & n47270;
  assign n47272 = ~n751 & n47271;
  assign n47273 = ~n212 & ~n663;
  assign n47274 = n16874 & n47273;
  assign n47275 = n28019 & n47274;
  assign n47276 = ~n221 & ~n830;
  assign n47277 = ~n1065 & n47276;
  assign n47278 = n12328 & n47277;
  assign n47279 = n46142 & n47278;
  assign n47280 = n47275 & n47279;
  assign n47281 = n28019 & n47276;
  assign n47282 = ~n663 & ~n1065;
  assign n47283 = n16874 & n47282;
  assign n47284 = n47281 & n47283;
  assign n47285 = n59566 & n47284;
  assign n47286 = n47247 & n47251;
  assign n47287 = ~n464 & ~n1646;
  assign n47288 = ~n1646 & ~n2201;
  assign n47289 = ~n464 & n47288;
  assign n47290 = ~n2201 & n47287;
  assign n47291 = n3262 & n59567;
  assign n47292 = n5848 & n53999;
  assign n47293 = n47291 & n47292;
  assign n47294 = n59565 & n47293;
  assign n47295 = n3262 & n5848;
  assign n47296 = n406 & n2814;
  assign n47297 = n53999 & n47296;
  assign n47298 = n47295 & n47297;
  assign n47299 = n3560 & n4261;
  assign n47300 = n47237 & n47299;
  assign n47301 = n648 & n3672;
  assign n47302 = n59567 & n47301;
  assign n47303 = n47300 & n47302;
  assign n47304 = n54158 & n47303;
  assign n47305 = n47298 & n47304;
  assign n47306 = n59565 & n47305;
  assign n47307 = n406 & n3672;
  assign n47308 = n2814 & n7307;
  assign n47309 = n47307 & n47308;
  assign n47310 = ~n464 & ~n2201;
  assign n47311 = n8268 & n47310;
  assign n47312 = n648 & n4261;
  assign n47313 = n47311 & n47312;
  assign n47314 = n47309 & n47313;
  assign n47315 = n54158 & n47314;
  assign n47316 = ~n1490 & ~n1646;
  assign n47317 = ~n166 & n47316;
  assign n47318 = n5848 & n47317;
  assign n47319 = n3262 & n53999;
  assign n47320 = n47318 & n47319;
  assign n47321 = n59565 & n47320;
  assign n47322 = n47315 & n47321;
  assign n47323 = n47244 & n47294;
  assign n47324 = n54494 & n59568;
  assign n47325 = n5848 & n8268;
  assign n47326 = n3262 & n47325;
  assign n47327 = n53999 & n47326;
  assign n47328 = n648 & n47327;
  assign n47329 = n2814 & n47328;
  assign n47330 = n7307 & n47329;
  assign n47331 = n54494 & n47330;
  assign n47332 = n54641 & n47331;
  assign n47333 = n54158 & n47332;
  assign n47334 = n59565 & n47333;
  assign n47335 = n4261 & n47334;
  assign n47336 = n406 & n47335;
  assign n47337 = n3672 & n47336;
  assign n47338 = ~n464 & n47337;
  assign n47339 = ~n1490 & n47338;
  assign n47340 = ~n166 & n47339;
  assign n47341 = ~n1646 & n47340;
  assign n47342 = ~n2201 & n47341;
  assign n47343 = n54641 & n47324;
  assign n47344 = n1576 & ~n58533;
  assign n47345 = n11215 & n39600;
  assign n47346 = n10564 & n39603;
  assign n47347 = n54403 & n39606;
  assign n47348 = ~n47346 & ~n47347;
  assign n47349 = ~n47345 & n47348;
  assign n47350 = ~n47344 & ~n47347;
  assign n47351 = ~n47346 & n47350;
  assign n47352 = ~n47345 & n47351;
  assign n47353 = ~n47344 & n47349;
  assign n47354 = ~n59569 & ~n59570;
  assign n47355 = n59569 & n59570;
  assign n47356 = ~n59569 & ~n47354;
  assign n47357 = ~n59569 & n59570;
  assign n47358 = ~n59570 & ~n47354;
  assign n47359 = n59569 & ~n59570;
  assign n47360 = ~n59571 & ~n59572;
  assign n47361 = ~n47354 & ~n47355;
  assign n47362 = ~n47236 & ~n59573;
  assign n47363 = n47236 & n59573;
  assign n47364 = ~n47236 & ~n47362;
  assign n47365 = ~n59573 & ~n47362;
  assign n47366 = ~n47364 & ~n47365;
  assign n47367 = ~n47362 & ~n47363;
  assign n47368 = ~n47235 & ~n59574;
  assign n47369 = n47235 & n59574;
  assign n47370 = ~n47368 & ~n47369;
  assign n47371 = ~n47222 & n47370;
  assign n47372 = n47222 & ~n47370;
  assign n47373 = ~n47371 & ~n47372;
  assign n47374 = n123 & n41007;
  assign n47375 = n128 & n39582;
  assign n47376 = n53444 & n39588;
  assign n47377 = n127 & n39585;
  assign n47378 = ~n47376 & ~n47377;
  assign n47379 = ~n47375 & n47378;
  assign n47380 = ~n123 & n47379;
  assign n47381 = ~n41007 & n47379;
  assign n47382 = ~n47380 & ~n47381;
  assign n47383 = ~n47374 & n47379;
  assign n47384 = pi26  & ~n59575;
  assign n47385 = ~pi26  & n59575;
  assign n47386 = ~n47384 & ~n47385;
  assign n47387 = n47373 & ~n47386;
  assign n47388 = ~n47373 & n47386;
  assign n47389 = n47373 & ~n47387;
  assign n47390 = n47373 & n47386;
  assign n47391 = ~n47386 & ~n47387;
  assign n47392 = ~n47373 & ~n47386;
  assign n47393 = ~n59576 & ~n59577;
  assign n47394 = ~n47387 & ~n47388;
  assign n47395 = ~n47221 & ~n59578;
  assign n47396 = n47221 & n59578;
  assign n47397 = ~n47221 & ~n47395;
  assign n47398 = ~n59578 & ~n47395;
  assign n47399 = ~n47397 & ~n47398;
  assign n47400 = ~n47395 & ~n47396;
  assign n47401 = ~n47220 & ~n59579;
  assign n47402 = n47220 & n59579;
  assign n47403 = ~n47220 & ~n47401;
  assign n47404 = ~n47220 & n59579;
  assign n47405 = ~n59579 & ~n47401;
  assign n47406 = n47220 & ~n59579;
  assign n47407 = ~n59580 & ~n59581;
  assign n47408 = ~n47401 & ~n47402;
  assign n47409 = n47207 & n59582;
  assign n47410 = ~n47207 & ~n59582;
  assign n47411 = ~n47409 & ~n47410;
  assign n47412 = n14413 & n41762;
  assign n47413 = n15921 & n39564;
  assign n47414 = n54719 & n39570;
  assign n47415 = n15901 & n39567;
  assign n47416 = ~n47414 & ~n47415;
  assign n47417 = ~n47413 & n47416;
  assign n47418 = ~n14413 & n47417;
  assign n47419 = ~n41762 & n47417;
  assign n47420 = ~n47418 & ~n47419;
  assign n47421 = ~n47412 & n47417;
  assign n47422 = pi20  & ~n59583;
  assign n47423 = ~pi20  & n59583;
  assign n47424 = ~n47422 & ~n47423;
  assign n47425 = n47411 & ~n47424;
  assign n47426 = ~n47411 & n47424;
  assign n47427 = n47411 & ~n47425;
  assign n47428 = n47411 & n47424;
  assign n47429 = ~n47424 & ~n47425;
  assign n47430 = ~n47411 & ~n47424;
  assign n47431 = ~n59584 & ~n59585;
  assign n47432 = ~n47425 & ~n47426;
  assign n47433 = ~n47206 & ~n59586;
  assign n47434 = n47206 & n59586;
  assign n47435 = ~n47206 & ~n47433;
  assign n47436 = ~n47206 & n59586;
  assign n47437 = ~n59586 & ~n47433;
  assign n47438 = n47206 & ~n59586;
  assign n47439 = ~n59587 & ~n59588;
  assign n47440 = ~n47433 & ~n47434;
  assign n47441 = ~n47205 & ~n59589;
  assign n47442 = n47205 & n59589;
  assign n47443 = ~n47205 & ~n47441;
  assign n47444 = ~n59589 & ~n47441;
  assign n47445 = ~n47443 & ~n47444;
  assign n47446 = ~n47441 & ~n47442;
  assign n47447 = n47192 & n59590;
  assign n47448 = ~n47192 & ~n59590;
  assign n47449 = ~n47447 & ~n47448;
  assign n47450 = n17265 & n43436;
  assign n47451 = n18588 & n39546;
  assign n47452 = n55041 & n39552;
  assign n47453 = n18556 & n39549;
  assign n47454 = ~n47452 & ~n47453;
  assign n47455 = ~n47451 & n47454;
  assign n47456 = ~n17265 & n47455;
  assign n47457 = ~n43436 & n47455;
  assign n47458 = ~n47456 & ~n47457;
  assign n47459 = ~n47450 & n47455;
  assign n47460 = pi14  & ~n59591;
  assign n47461 = ~pi14  & n59591;
  assign n47462 = ~n47460 & ~n47461;
  assign n47463 = n47449 & ~n47462;
  assign n47464 = ~n47449 & n47462;
  assign n47465 = n47449 & ~n47463;
  assign n47466 = n47449 & n47462;
  assign n47467 = ~n47462 & ~n47463;
  assign n47468 = ~n47449 & ~n47462;
  assign n47469 = ~n59592 & ~n59593;
  assign n47470 = ~n47463 & ~n47464;
  assign n47471 = ~n47191 & ~n59594;
  assign n47472 = n47191 & n59594;
  assign n47473 = ~n47191 & ~n47471;
  assign n47474 = ~n59594 & ~n47471;
  assign n47475 = ~n47473 & ~n47474;
  assign n47476 = ~n47471 & ~n47472;
  assign n47477 = ~n47190 & ~n59595;
  assign n47478 = n47190 & n59595;
  assign n47479 = ~n47190 & ~n47477;
  assign n47480 = ~n47190 & n59595;
  assign n47481 = ~n59595 & ~n47477;
  assign n47482 = n47190 & ~n59595;
  assign n47483 = ~n59596 & ~n59597;
  assign n47484 = ~n47477 & ~n47478;
  assign n47485 = n47177 & n59598;
  assign n47486 = ~n47177 & ~n59598;
  assign n47487 = ~n47485 & ~n47486;
  assign n47488 = n20085 & ~n59280;
  assign n47489 = n21269 & n44871;
  assign n47490 = n55472 & n44327;
  assign n47491 = n21237 & n44775;
  assign n47492 = ~n47490 & ~n47491;
  assign n47493 = ~n47489 & n47492;
  assign n47494 = ~n20085 & n47493;
  assign n47495 = n59280 & n47493;
  assign n47496 = ~n47494 & ~n47495;
  assign n47497 = ~n47488 & n47493;
  assign n47498 = pi8  & ~n59599;
  assign n47499 = ~pi8  & n59599;
  assign n47500 = ~n47498 & ~n47499;
  assign n47501 = n47487 & ~n47500;
  assign n47502 = ~n47487 & n47500;
  assign n47503 = n47487 & ~n47501;
  assign n47504 = n47487 & n47500;
  assign n47505 = ~n47500 & ~n47501;
  assign n47506 = ~n47487 & ~n47500;
  assign n47507 = ~n59600 & ~n59601;
  assign n47508 = ~n47501 & ~n47502;
  assign n47509 = ~n47176 & ~n59602;
  assign n47510 = n47176 & n59602;
  assign n47511 = ~n47176 & ~n47509;
  assign n47512 = ~n47176 & n59602;
  assign n47513 = ~n59602 & ~n47509;
  assign n47514 = n47176 & ~n59602;
  assign n47515 = ~n59603 & ~n59604;
  assign n47516 = ~n47509 & ~n47510;
  assign n47517 = ~n47175 & ~n59605;
  assign n47518 = n47175 & n59605;
  assign n47519 = ~n47175 & ~n47517;
  assign n47520 = ~n59605 & ~n47517;
  assign n47521 = ~n47519 & ~n47520;
  assign n47522 = ~n47517 & ~n47518;
  assign n47523 = n47162 & n59606;
  assign n47524 = ~n47162 & ~n59606;
  assign n47525 = ~n47523 & ~n47524;
  assign n47526 = ~n59503 & ~n47133;
  assign n47527 = n24338 & ~n47526;
  assign n47528 = n24337 & n46788;
  assign n47529 = n25272 & n59503;
  assign n47530 = ~n47528 & ~n47529;
  assign n47531 = ~n24338 & n47530;
  assign n47532 = n47526 & n47530;
  assign n47533 = ~n47531 & ~n47532;
  assign n47534 = ~n47527 & n47530;
  assign n47535 = pi2  & ~n59607;
  assign n47536 = ~pi2  & n59607;
  assign n47537 = ~n47535 & ~n47536;
  assign n47538 = n47525 & ~n47537;
  assign n47539 = ~n47525 & n47537;
  assign n47540 = ~n47538 & ~n47539;
  assign n47541 = ~n47161 & n47540;
  assign n47542 = n47161 & ~n47540;
  assign n47543 = ~n47541 & ~n47542;
  assign n47544 = n47158 & n47543;
  assign n47545 = ~n47158 & ~n47543;
  assign po4  = ~n47544 & ~n47545;
  assign n47547 = ~n47538 & ~n47541;
  assign n47548 = ~n47517 & ~n47524;
  assign n47549 = n77 & n46805;
  assign n47550 = n24302 & n46788;
  assign n47551 = n21969 & n46009;
  assign n47552 = n23459 & n46420;
  assign n47553 = ~n47551 & ~n47552;
  assign n47554 = ~n47550 & n47553;
  assign n47555 = ~n47549 & n47554;
  assign n47556 = pi5  & ~n47555;
  assign n47557 = ~n47555 & ~n47556;
  assign n47558 = ~pi5  & ~n47555;
  assign n47559 = pi5  & ~n47556;
  assign n47560 = pi5  & n47555;
  assign n47561 = ~n59608 & ~n59609;
  assign n47562 = ~n47501 & ~n47509;
  assign n47563 = ~n47477 & ~n47486;
  assign n47564 = n18846 & ~n59184;
  assign n47565 = n19541 & n44327;
  assign n47566 = n55247 & n39543;
  assign n47567 = n19509 & n39937;
  assign n47568 = ~n47566 & ~n47567;
  assign n47569 = ~n47565 & n47568;
  assign n47570 = ~n47564 & n47569;
  assign n47571 = pi11  & ~n47570;
  assign n47572 = ~n47570 & ~n47571;
  assign n47573 = ~pi11  & ~n47570;
  assign n47574 = pi11  & ~n47571;
  assign n47575 = pi11  & n47570;
  assign n47576 = ~n59610 & ~n59611;
  assign n47577 = ~n47463 & ~n47471;
  assign n47578 = ~n47441 & ~n47448;
  assign n47579 = n16079 & ~n58891;
  assign n47580 = n16696 & n39552;
  assign n47581 = n54886 & n39558;
  assign n47582 = n16676 & n39555;
  assign n47583 = ~n47581 & ~n47582;
  assign n47584 = ~n47580 & n47583;
  assign n47585 = ~n47579 & n47584;
  assign n47586 = pi17  & ~n47585;
  assign n47587 = ~n47585 & ~n47586;
  assign n47588 = ~pi17  & ~n47585;
  assign n47589 = pi17  & ~n47586;
  assign n47590 = pi17  & n47585;
  assign n47591 = ~n59612 & ~n59613;
  assign n47592 = ~n47425 & ~n47433;
  assign n47593 = ~n47401 & ~n47410;
  assign n47594 = n90 & ~n58759;
  assign n47595 = n14236 & n39570;
  assign n47596 = n54667 & n39576;
  assign n47597 = n14210 & n39573;
  assign n47598 = ~n47596 & ~n47597;
  assign n47599 = ~n47595 & n47598;
  assign n47600 = ~n47594 & n47599;
  assign n47601 = pi23  & ~n47600;
  assign n47602 = ~n47600 & ~n47601;
  assign n47603 = ~pi23  & ~n47600;
  assign n47604 = pi23  & ~n47601;
  assign n47605 = pi23  & n47600;
  assign n47606 = ~n59614 & ~n59615;
  assign n47607 = ~n47387 & ~n47395;
  assign n47608 = ~n47368 & ~n47371;
  assign n47609 = n11279 & ~n58585;
  assign n47610 = n12584 & n39588;
  assign n47611 = n54410 & n39594;
  assign n47612 = n11267 & n39591;
  assign n47613 = ~n47611 & ~n47612;
  assign n47614 = ~n47610 & n47613;
  assign n47615 = ~n11279 & n47614;
  assign n47616 = n58585 & n47614;
  assign n47617 = ~n47615 & ~n47616;
  assign n47618 = ~n47609 & n47614;
  assign n47619 = pi29  & ~n59616;
  assign n47620 = ~pi29  & n59616;
  assign n47621 = ~n47619 & ~n47620;
  assign n47622 = ~n47354 & ~n47362;
  assign n47623 = n7024 & n11628;
  assign n47624 = n15060 & n47623;
  assign n47625 = n53714 & n47624;
  assign n47626 = n54449 & n47625;
  assign n47627 = ~n747 & ~n948;
  assign n47628 = ~n1196 & n47627;
  assign n47629 = ~n414 & ~n499;
  assign n47630 = n1541 & n47629;
  assign n47631 = n3369 & n4892;
  assign n47632 = n47630 & n47631;
  assign n47633 = n47628 & n47632;
  assign n47634 = n54432 & n47633;
  assign n47635 = n4892 & n7024;
  assign n47636 = n15060 & n47635;
  assign n47637 = n53714 & n47636;
  assign n47638 = n54449 & n47637;
  assign n47639 = n11628 & n47629;
  assign n47640 = n1541 & n3369;
  assign n47641 = n47639 & n47640;
  assign n47642 = n47628 & n47641;
  assign n47643 = n54432 & n47642;
  assign n47644 = n47638 & n47643;
  assign n47645 = n7024 & n47631;
  assign n47646 = n53714 & n47645;
  assign n47647 = n54449 & n47646;
  assign n47648 = ~n409 & ~n1196;
  assign n47649 = ~n747 & n47648;
  assign n47650 = ~n414 & ~n948;
  assign n47651 = ~n499 & ~n2109;
  assign n47652 = n47650 & n47651;
  assign n47653 = n1541 & n15060;
  assign n47654 = n47652 & n47653;
  assign n47655 = n47649 & n47654;
  assign n47656 = n54432 & n47655;
  assign n47657 = n47647 & n47656;
  assign n47658 = n1541 & n47631;
  assign n47659 = n53714 & n47658;
  assign n47660 = n54449 & n47659;
  assign n47661 = ~n735 & ~n2109;
  assign n47662 = ~n499 & n47661;
  assign n47663 = ~n414 & ~n1196;
  assign n47664 = ~n507 & ~n747;
  assign n47665 = n47663 & n47664;
  assign n47666 = ~n409 & ~n948;
  assign n47667 = n7024 & n47666;
  assign n47668 = n47665 & n47667;
  assign n47669 = n47662 & n47668;
  assign n47670 = n54432 & n47669;
  assign n47671 = n47660 & n47670;
  assign n47672 = n47626 & n47634;
  assign n47673 = n54827 & n59617;
  assign n47674 = n53714 & n3369;
  assign n47675 = n4892 & n47674;
  assign n47676 = n54449 & n47675;
  assign n47677 = n57048 & n47676;
  assign n47678 = n54432 & n47677;
  assign n47679 = n54827 & n47678;
  assign n47680 = n1541 & n47679;
  assign n47681 = ~n948 & n47680;
  assign n47682 = ~n1065 & n47681;
  assign n47683 = ~n414 & n47682;
  assign n47684 = ~n1196 & n47683;
  assign n47685 = ~n852 & n47684;
  assign n47686 = ~n507 & n47685;
  assign n47687 = ~n499 & n47686;
  assign n47688 = ~n409 & n47687;
  assign n47689 = ~n747 & n47688;
  assign n47690 = ~n735 & n47689;
  assign n47691 = ~n2109 & n47690;
  assign n47692 = n57048 & n47673;
  assign n47693 = n1576 & n40247;
  assign n47694 = n11215 & n39597;
  assign n47695 = n10564 & n39600;
  assign n47696 = n54403 & n39603;
  assign n47697 = ~n47695 & ~n47696;
  assign n47698 = ~n47694 & n47697;
  assign n47699 = ~n47693 & ~n47696;
  assign n47700 = ~n47695 & n47699;
  assign n47701 = ~n47694 & n47700;
  assign n47702 = ~n47693 & n47698;
  assign n47703 = ~n59618 & ~n59619;
  assign n47704 = n59618 & n59619;
  assign n47705 = ~n59618 & ~n47703;
  assign n47706 = ~n59618 & n59619;
  assign n47707 = ~n59619 & ~n47703;
  assign n47708 = n59618 & ~n59619;
  assign n47709 = ~n59620 & ~n59621;
  assign n47710 = ~n47703 & ~n47704;
  assign n47711 = ~n47622 & ~n59622;
  assign n47712 = n47622 & n59622;
  assign n47713 = ~n47622 & ~n47711;
  assign n47714 = ~n59622 & ~n47711;
  assign n47715 = ~n47713 & ~n47714;
  assign n47716 = ~n47711 & ~n47712;
  assign n47717 = ~n47621 & ~n59623;
  assign n47718 = n47621 & n59623;
  assign n47719 = ~n47717 & ~n47718;
  assign n47720 = ~n47608 & n47719;
  assign n47721 = n47608 & ~n47719;
  assign n47722 = ~n47720 & ~n47721;
  assign n47723 = n123 & ~n58657;
  assign n47724 = n128 & n39579;
  assign n47725 = n53444 & n39585;
  assign n47726 = n127 & n39582;
  assign n47727 = ~n47725 & ~n47726;
  assign n47728 = ~n47724 & n47727;
  assign n47729 = ~n123 & n47728;
  assign n47730 = n58657 & n47728;
  assign n47731 = ~n47729 & ~n47730;
  assign n47732 = ~n47723 & n47728;
  assign n47733 = pi26  & ~n59624;
  assign n47734 = ~pi26  & n59624;
  assign n47735 = ~n47733 & ~n47734;
  assign n47736 = n47722 & ~n47735;
  assign n47737 = ~n47722 & n47735;
  assign n47738 = n47722 & ~n47736;
  assign n47739 = n47722 & n47735;
  assign n47740 = ~n47735 & ~n47736;
  assign n47741 = ~n47722 & ~n47735;
  assign n47742 = ~n59625 & ~n59626;
  assign n47743 = ~n47736 & ~n47737;
  assign n47744 = ~n47607 & ~n59627;
  assign n47745 = n47607 & n59627;
  assign n47746 = ~n47607 & ~n47744;
  assign n47747 = ~n59627 & ~n47744;
  assign n47748 = ~n47746 & ~n47747;
  assign n47749 = ~n47744 & ~n47745;
  assign n47750 = ~n47606 & ~n59628;
  assign n47751 = n47606 & n59628;
  assign n47752 = ~n47606 & ~n47750;
  assign n47753 = ~n47606 & n59628;
  assign n47754 = ~n59628 & ~n47750;
  assign n47755 = n47606 & ~n59628;
  assign n47756 = ~n59629 & ~n59630;
  assign n47757 = ~n47750 & ~n47751;
  assign n47758 = n47593 & n59631;
  assign n47759 = ~n47593 & ~n59631;
  assign n47760 = ~n47758 & ~n47759;
  assign n47761 = n14413 & ~n58493;
  assign n47762 = n15921 & n39561;
  assign n47763 = n54719 & n39567;
  assign n47764 = n15901 & n39564;
  assign n47765 = ~n47763 & ~n47764;
  assign n47766 = ~n47762 & n47765;
  assign n47767 = ~n14413 & n47766;
  assign n47768 = n58493 & n47766;
  assign n47769 = ~n47767 & ~n47768;
  assign n47770 = ~n47761 & n47766;
  assign n47771 = pi20  & ~n59632;
  assign n47772 = ~pi20  & n59632;
  assign n47773 = ~n47771 & ~n47772;
  assign n47774 = n47760 & ~n47773;
  assign n47775 = ~n47760 & n47773;
  assign n47776 = n47760 & ~n47774;
  assign n47777 = n47760 & n47773;
  assign n47778 = ~n47773 & ~n47774;
  assign n47779 = ~n47760 & ~n47773;
  assign n47780 = ~n59633 & ~n59634;
  assign n47781 = ~n47774 & ~n47775;
  assign n47782 = ~n47592 & ~n59635;
  assign n47783 = n47592 & n59635;
  assign n47784 = ~n47592 & ~n47782;
  assign n47785 = ~n47592 & n59635;
  assign n47786 = ~n59635 & ~n47782;
  assign n47787 = n47592 & ~n59635;
  assign n47788 = ~n59636 & ~n59637;
  assign n47789 = ~n47782 & ~n47783;
  assign n47790 = ~n47591 & ~n59638;
  assign n47791 = n47591 & n59638;
  assign n47792 = ~n47591 & ~n47790;
  assign n47793 = ~n59638 & ~n47790;
  assign n47794 = ~n47792 & ~n47793;
  assign n47795 = ~n47790 & ~n47791;
  assign n47796 = n47578 & n59639;
  assign n47797 = ~n47578 & ~n59639;
  assign n47798 = ~n47796 & ~n47797;
  assign n47799 = n17265 & ~n59050;
  assign n47800 = n18588 & n39440;
  assign n47801 = n55041 & n39549;
  assign n47802 = n18556 & n39546;
  assign n47803 = ~n47801 & ~n47802;
  assign n47804 = ~n47800 & n47803;
  assign n47805 = ~n17265 & n47804;
  assign n47806 = n59050 & n47804;
  assign n47807 = ~n47805 & ~n47806;
  assign n47808 = ~n47799 & n47804;
  assign n47809 = pi14  & ~n59640;
  assign n47810 = ~pi14  & n59640;
  assign n47811 = ~n47809 & ~n47810;
  assign n47812 = n47798 & ~n47811;
  assign n47813 = ~n47798 & n47811;
  assign n47814 = n47798 & ~n47812;
  assign n47815 = n47798 & n47811;
  assign n47816 = ~n47811 & ~n47812;
  assign n47817 = ~n47798 & ~n47811;
  assign n47818 = ~n59641 & ~n59642;
  assign n47819 = ~n47812 & ~n47813;
  assign n47820 = ~n47577 & ~n59643;
  assign n47821 = n47577 & n59643;
  assign n47822 = ~n47577 & ~n47820;
  assign n47823 = ~n59643 & ~n47820;
  assign n47824 = ~n47822 & ~n47823;
  assign n47825 = ~n47820 & ~n47821;
  assign n47826 = ~n47576 & ~n59644;
  assign n47827 = n47576 & n59644;
  assign n47828 = ~n47576 & ~n47826;
  assign n47829 = ~n47576 & n59644;
  assign n47830 = ~n59644 & ~n47826;
  assign n47831 = n47576 & ~n59644;
  assign n47832 = ~n59645 & ~n59646;
  assign n47833 = ~n47826 & ~n47827;
  assign n47834 = n47563 & n59647;
  assign n47835 = ~n47563 & ~n59647;
  assign n47836 = ~n47834 & ~n47835;
  assign n47837 = n20085 & ~n59275;
  assign n47838 = n21269 & n44952;
  assign n47839 = n55472 & n44775;
  assign n47840 = n21237 & n44871;
  assign n47841 = ~n47839 & ~n47840;
  assign n47842 = ~n47838 & n47841;
  assign n47843 = ~n20085 & n47842;
  assign n47844 = n59275 & n47842;
  assign n47845 = ~n47843 & ~n47844;
  assign n47846 = ~n47837 & n47842;
  assign n47847 = pi8  & ~n59648;
  assign n47848 = ~pi8  & n59648;
  assign n47849 = ~n47847 & ~n47848;
  assign n47850 = n47836 & ~n47849;
  assign n47851 = ~n47836 & n47849;
  assign n47852 = n47836 & ~n47850;
  assign n47853 = n47836 & n47849;
  assign n47854 = ~n47849 & ~n47850;
  assign n47855 = ~n47836 & ~n47849;
  assign n47856 = ~n59649 & ~n59650;
  assign n47857 = ~n47850 & ~n47851;
  assign n47858 = ~n47562 & ~n59651;
  assign n47859 = n47562 & n59651;
  assign n47860 = ~n47562 & ~n47858;
  assign n47861 = ~n47562 & n59651;
  assign n47862 = ~n59651 & ~n47858;
  assign n47863 = n47562 & ~n59651;
  assign n47864 = ~n59652 & ~n59653;
  assign n47865 = ~n47858 & ~n47859;
  assign n47866 = ~n47561 & ~n59654;
  assign n47867 = n47561 & n59654;
  assign n47868 = ~n47561 & ~n47866;
  assign n47869 = ~n59654 & ~n47866;
  assign n47870 = ~n47868 & ~n47869;
  assign n47871 = ~n47866 & ~n47867;
  assign n47872 = n47548 & n59655;
  assign n47873 = ~n47548 & ~n59655;
  assign n47874 = ~n47872 & ~n47873;
  assign n47875 = n24337 & n59503;
  assign n47876 = pi2  & ~n47875;
  assign n47877 = n47874 & n47876;
  assign n47878 = ~n47874 & ~n47876;
  assign n47879 = ~n47877 & ~n47878;
  assign n47880 = ~n47547 & n47879;
  assign n47881 = n47547 & ~n47879;
  assign n47882 = ~n47880 & ~n47881;
  assign n47883 = n47544 & n47882;
  assign n47884 = ~n47544 & ~n47882;
  assign po5  = ~n47883 & ~n47884;
  assign n47886 = ~n47866 & ~n47873;
  assign n47887 = n77 & ~n59554;
  assign n47888 = n24302 & n59503;
  assign n47889 = n21969 & n46420;
  assign n47890 = n23459 & n46788;
  assign n47891 = ~n47889 & ~n47890;
  assign n47892 = ~n47888 & n47891;
  assign n47893 = ~n47887 & n47892;
  assign n47894 = pi5  & ~n47893;
  assign n47895 = ~n47893 & ~n47894;
  assign n47896 = ~pi5  & ~n47893;
  assign n47897 = pi5  & ~n47894;
  assign n47898 = pi5  & n47893;
  assign n47899 = ~n59656 & ~n59657;
  assign n47900 = ~n47850 & ~n47858;
  assign n47901 = ~n47826 & ~n47835;
  assign n47902 = n18846 & ~n59282;
  assign n47903 = n19541 & n44775;
  assign n47904 = n55247 & n39937;
  assign n47905 = n19509 & n44327;
  assign n47906 = ~n47904 & ~n47905;
  assign n47907 = ~n47903 & n47906;
  assign n47908 = ~n47902 & n47907;
  assign n47909 = pi11  & ~n47908;
  assign n47910 = ~n47908 & ~n47909;
  assign n47911 = ~pi11  & ~n47908;
  assign n47912 = pi11  & ~n47909;
  assign n47913 = pi11  & n47908;
  assign n47914 = ~n59658 & ~n59659;
  assign n47915 = ~n47812 & ~n47820;
  assign n47916 = ~n47790 & ~n47797;
  assign n47917 = n16079 & ~n58889;
  assign n47918 = n16696 & n39549;
  assign n47919 = n54886 & n39555;
  assign n47920 = n16676 & n39552;
  assign n47921 = ~n47919 & ~n47920;
  assign n47922 = ~n47918 & n47921;
  assign n47923 = ~n47917 & n47922;
  assign n47924 = pi17  & ~n47923;
  assign n47925 = ~n47923 & ~n47924;
  assign n47926 = ~pi17  & ~n47923;
  assign n47927 = pi17  & ~n47924;
  assign n47928 = pi17  & n47923;
  assign n47929 = ~n59660 & ~n59661;
  assign n47930 = ~n47774 & ~n47782;
  assign n47931 = ~n47750 & ~n47759;
  assign n47932 = n90 & ~n58766;
  assign n47933 = n14236 & n39567;
  assign n47934 = n54667 & n39573;
  assign n47935 = n14210 & n39570;
  assign n47936 = ~n47934 & ~n47935;
  assign n47937 = ~n47933 & n47936;
  assign n47938 = ~n47932 & n47937;
  assign n47939 = pi23  & ~n47938;
  assign n47940 = ~n47938 & ~n47939;
  assign n47941 = ~pi23  & ~n47938;
  assign n47942 = pi23  & ~n47939;
  assign n47943 = pi23  & n47938;
  assign n47944 = ~n59662 & ~n59663;
  assign n47945 = ~n47736 & ~n47744;
  assign n47946 = ~n47717 & ~n47720;
  assign n47947 = n11279 & ~n58583;
  assign n47948 = n12584 & n39585;
  assign n47949 = n54410 & n39591;
  assign n47950 = n11267 & n39588;
  assign n47951 = ~n47949 & ~n47950;
  assign n47952 = ~n47948 & n47951;
  assign n47953 = ~n11279 & n47952;
  assign n47954 = n58583 & n47952;
  assign n47955 = ~n47953 & ~n47954;
  assign n47956 = ~n47947 & n47952;
  assign n47957 = pi29  & ~n59664;
  assign n47958 = ~pi29  & n59664;
  assign n47959 = ~n47957 & ~n47958;
  assign n47960 = ~n47703 & ~n47711;
  assign n47961 = n4383 & n4587;
  assign n47962 = n6301 & n47961;
  assign n47963 = n56752 & n47962;
  assign n47964 = n59514 & n47963;
  assign n47965 = ~n560 & ~n975;
  assign n47966 = n2666 & n47965;
  assign n47967 = n1956 & n6897;
  assign n47968 = n14924 & n47967;
  assign n47969 = ~n291 & ~n560;
  assign n47970 = n6897 & n47969;
  assign n47971 = ~n291 & n47967;
  assign n47972 = ~n560 & n47971;
  assign n47973 = n1956 & n47970;
  assign n47974 = ~n975 & n59665;
  assign n47975 = ~n443 & n47974;
  assign n47976 = ~n774 & n47975;
  assign n47977 = ~n735 & n47976;
  assign n47978 = n6897 & n47965;
  assign n47979 = n1956 & n2666;
  assign n47980 = n14924 & n47979;
  assign n47981 = n47978 & n47980;
  assign n47982 = ~n443 & ~n975;
  assign n47983 = n14924 & n47982;
  assign n47984 = n59665 & n47983;
  assign n47985 = n47966 & n47968;
  assign n47986 = ~n177 & ~n268;
  assign n47987 = n3014 & n47986;
  assign n47988 = n3678 & n4319;
  assign n47989 = n47987 & n47988;
  assign n47990 = ~n465 & ~n751;
  assign n47991 = ~n741 & ~n911;
  assign n47992 = n47990 & n47991;
  assign n47993 = n47296 & n47992;
  assign n47994 = ~n268 & ~n465;
  assign n47995 = n3014 & n47994;
  assign n47996 = n47988 & n47995;
  assign n47997 = ~n177 & ~n741;
  assign n47998 = ~n751 & ~n911;
  assign n47999 = n47997 & n47998;
  assign n48000 = n47296 & n47999;
  assign n48001 = n47996 & n48000;
  assign n48002 = n47989 & n47993;
  assign n48003 = n59666 & n59667;
  assign n48004 = n3678 & n4383;
  assign n48005 = n6301 & n48004;
  assign n48006 = n56752 & n48005;
  assign n48007 = n59514 & n48006;
  assign n48008 = n3014 & n4587;
  assign n48009 = n47296 & n48008;
  assign n48010 = ~n465 & ~n741;
  assign n48011 = ~n268 & ~n911;
  assign n48012 = n48010 & n48011;
  assign n48013 = ~n177 & ~n751;
  assign n48014 = n4319 & n48013;
  assign n48015 = n48012 & n48014;
  assign n48016 = n48009 & n48015;
  assign n48017 = n59666 & n48016;
  assign n48018 = n48007 & n48017;
  assign n48019 = n406 & n4587;
  assign n48020 = n2814 & n48019;
  assign n48021 = n56752 & n48020;
  assign n48022 = n59514 & n48021;
  assign n48023 = n3014 & n4319;
  assign n48024 = n48004 & n48023;
  assign n48025 = ~n177 & ~n911;
  assign n48026 = n47994 & n48025;
  assign n48027 = ~n741 & ~n751;
  assign n48028 = n6301 & n48027;
  assign n48029 = n48026 & n48028;
  assign n48030 = n48024 & n48029;
  assign n48031 = n59666 & n48030;
  assign n48032 = n48022 & n48031;
  assign n48033 = n47964 & n48003;
  assign n48034 = n54250 & n54779;
  assign n48035 = n56857 & n48034;
  assign n48036 = n4383 & n59514;
  assign n48037 = n3678 & n48036;
  assign n48038 = n2814 & n48037;
  assign n48039 = n59666 & n48038;
  assign n48040 = n56752 & n48039;
  assign n48041 = n54779 & n48040;
  assign n48042 = n56857 & n48041;
  assign n48043 = n4587 & n48042;
  assign n48044 = n406 & n48043;
  assign n48045 = n4319 & n48044;
  assign n48046 = n54250 & n48045;
  assign n48047 = n3014 & n48046;
  assign n48048 = ~n177 & n48047;
  assign n48049 = ~n911 & n48048;
  assign n48050 = ~n268 & n48049;
  assign n48051 = ~n364 & n48050;
  assign n48052 = ~n465 & n48051;
  assign n48053 = ~n741 & n48052;
  assign n48054 = ~n751 & n48053;
  assign n48055 = ~n625 & n48054;
  assign n48056 = n59668 & n48035;
  assign n48057 = n1576 & n40476;
  assign n48058 = n11215 & n39594;
  assign n48059 = n10564 & n39597;
  assign n48060 = n54403 & n39600;
  assign n48061 = ~n48059 & ~n48060;
  assign n48062 = ~n48058 & n48061;
  assign n48063 = ~n48057 & ~n48060;
  assign n48064 = ~n48059 & n48063;
  assign n48065 = ~n48058 & n48064;
  assign n48066 = ~n48057 & n48062;
  assign n48067 = ~n59669 & ~n59670;
  assign n48068 = n59669 & n59670;
  assign n48069 = ~n59669 & ~n48067;
  assign n48070 = ~n59669 & n59670;
  assign n48071 = ~n59670 & ~n48067;
  assign n48072 = n59669 & ~n59670;
  assign n48073 = ~n59671 & ~n59672;
  assign n48074 = ~n48067 & ~n48068;
  assign n48075 = ~n47960 & ~n59673;
  assign n48076 = n47960 & n59673;
  assign n48077 = ~n47960 & ~n48075;
  assign n48078 = ~n59673 & ~n48075;
  assign n48079 = ~n48077 & ~n48078;
  assign n48080 = ~n48075 & ~n48076;
  assign n48081 = ~n47959 & ~n59674;
  assign n48082 = n47959 & n59674;
  assign n48083 = ~n48081 & ~n48082;
  assign n48084 = ~n47946 & n48083;
  assign n48085 = n47946 & ~n48083;
  assign n48086 = ~n48084 & ~n48085;
  assign n48087 = n123 & ~n58653;
  assign n48088 = n128 & n39576;
  assign n48089 = n53444 & n39582;
  assign n48090 = n127 & n39579;
  assign n48091 = ~n48089 & ~n48090;
  assign n48092 = ~n48088 & n48091;
  assign n48093 = ~n123 & n48092;
  assign n48094 = n58653 & n48092;
  assign n48095 = ~n48093 & ~n48094;
  assign n48096 = ~n48087 & n48092;
  assign n48097 = pi26  & ~n59675;
  assign n48098 = ~pi26  & n59675;
  assign n48099 = ~n48097 & ~n48098;
  assign n48100 = n48086 & ~n48099;
  assign n48101 = ~n48086 & n48099;
  assign n48102 = ~n48100 & ~n48101;
  assign n48103 = ~n47945 & n48102;
  assign n48104 = n47945 & ~n48102;
  assign n48105 = ~n48103 & ~n48104;
  assign n48106 = ~n47944 & n48105;
  assign n48107 = n47944 & ~n48105;
  assign n48108 = ~n47944 & ~n48106;
  assign n48109 = ~n47944 & ~n48105;
  assign n48110 = n48105 & ~n48106;
  assign n48111 = n47944 & n48105;
  assign n48112 = ~n59676 & ~n59677;
  assign n48113 = ~n48106 & ~n48107;
  assign n48114 = n47931 & n59678;
  assign n48115 = ~n47931 & ~n59678;
  assign n48116 = ~n48114 & ~n48115;
  assign n48117 = n14413 & ~n58849;
  assign n48118 = n15921 & n39558;
  assign n48119 = n54719 & n39564;
  assign n48120 = n15901 & n39561;
  assign n48121 = ~n48119 & ~n48120;
  assign n48122 = ~n48118 & n48121;
  assign n48123 = ~n14413 & n48122;
  assign n48124 = n58849 & n48122;
  assign n48125 = ~n48123 & ~n48124;
  assign n48126 = ~n48117 & n48122;
  assign n48127 = pi20  & ~n59679;
  assign n48128 = ~pi20  & n59679;
  assign n48129 = ~n48127 & ~n48128;
  assign n48130 = n48116 & ~n48129;
  assign n48131 = ~n48116 & n48129;
  assign n48132 = ~n48130 & ~n48131;
  assign n48133 = ~n47930 & n48132;
  assign n48134 = n47930 & ~n48132;
  assign n48135 = ~n48133 & ~n48134;
  assign n48136 = ~n47929 & n48135;
  assign n48137 = n47929 & ~n48135;
  assign n48138 = ~n47929 & ~n48136;
  assign n48139 = ~n47929 & ~n48135;
  assign n48140 = n48135 & ~n48136;
  assign n48141 = n47929 & n48135;
  assign n48142 = ~n59680 & ~n59681;
  assign n48143 = ~n48136 & ~n48137;
  assign n48144 = n47916 & n59682;
  assign n48145 = ~n47916 & ~n59682;
  assign n48146 = ~n48144 & ~n48145;
  assign n48147 = n17265 & ~n59044;
  assign n48148 = n18588 & n39543;
  assign n48149 = n55041 & n39546;
  assign n48150 = n18556 & n39440;
  assign n48151 = ~n48149 & ~n48150;
  assign n48152 = ~n48148 & n48151;
  assign n48153 = ~n17265 & n48152;
  assign n48154 = n59044 & n48152;
  assign n48155 = ~n48153 & ~n48154;
  assign n48156 = ~n48147 & n48152;
  assign n48157 = pi14  & ~n59683;
  assign n48158 = ~pi14  & n59683;
  assign n48159 = ~n48157 & ~n48158;
  assign n48160 = n48146 & ~n48159;
  assign n48161 = ~n48146 & n48159;
  assign n48162 = ~n48160 & ~n48161;
  assign n48163 = ~n47915 & n48162;
  assign n48164 = n47915 & ~n48162;
  assign n48165 = ~n48163 & ~n48164;
  assign n48166 = ~n47914 & n48165;
  assign n48167 = n47914 & ~n48165;
  assign n48168 = ~n47914 & ~n48166;
  assign n48169 = ~n47914 & ~n48165;
  assign n48170 = n48165 & ~n48166;
  assign n48171 = n47914 & n48165;
  assign n48172 = ~n59684 & ~n59685;
  assign n48173 = ~n48166 & ~n48167;
  assign n48174 = n47901 & n59686;
  assign n48175 = ~n47901 & ~n59686;
  assign n48176 = ~n48174 & ~n48175;
  assign n48177 = n20085 & ~n59386;
  assign n48178 = n21269 & n46009;
  assign n48179 = n55472 & n44871;
  assign n48180 = n21237 & n44952;
  assign n48181 = ~n48179 & ~n48180;
  assign n48182 = ~n48178 & n48181;
  assign n48183 = ~n20085 & n48182;
  assign n48184 = n59386 & n48182;
  assign n48185 = ~n48183 & ~n48184;
  assign n48186 = ~n48177 & n48182;
  assign n48187 = pi8  & ~n59687;
  assign n48188 = ~pi8  & n59687;
  assign n48189 = ~n48187 & ~n48188;
  assign n48190 = n48176 & ~n48189;
  assign n48191 = ~n48176 & n48189;
  assign n48192 = ~n48190 & ~n48191;
  assign n48193 = ~n47900 & n48192;
  assign n48194 = n47900 & ~n48192;
  assign n48195 = ~n48193 & ~n48194;
  assign n48196 = ~n47899 & n48195;
  assign n48197 = n47899 & ~n48195;
  assign n48198 = ~n47899 & ~n48196;
  assign n48199 = ~n47899 & ~n48195;
  assign n48200 = n48195 & ~n48196;
  assign n48201 = n47899 & n48195;
  assign n48202 = ~n59688 & ~n59689;
  assign n48203 = ~n48196 & ~n48197;
  assign n48204 = pi2  & ~n59690;
  assign n48205 = ~pi2  & n59690;
  assign n48206 = ~n59690 & ~n48204;
  assign n48207 = pi2  & ~n48204;
  assign n48208 = ~n48206 & ~n48207;
  assign n48209 = ~n48204 & ~n48205;
  assign n48210 = n47886 & n59691;
  assign n48211 = ~n47886 & ~n59691;
  assign n48212 = ~n48210 & ~n48211;
  assign n48213 = ~n47877 & ~n47880;
  assign n48214 = ~n48212 & n48213;
  assign n48215 = n48212 & ~n48213;
  assign n48216 = ~n48214 & ~n48215;
  assign n48217 = n47883 & n48216;
  assign n48218 = ~n47883 & ~n48216;
  assign po6  = ~n48217 & ~n48218;
  assign n48220 = ~n48196 & ~n48204;
  assign n48221 = ~n48190 & ~n48193;
  assign n48222 = ~n48166 & ~n48175;
  assign n48223 = ~n48160 & ~n48163;
  assign n48224 = ~n48136 & ~n48145;
  assign n48225 = ~n48130 & ~n48133;
  assign n48226 = ~n48106 & ~n48115;
  assign n48227 = ~n48100 & ~n48103;
  assign n48228 = ~n48081 & ~n48084;
  assign n48229 = ~n48067 & ~n48075;
  assign n48230 = ~n274 & ~n466;
  assign n48231 = ~n852 & ~n894;
  assign n48232 = n48230 & n48231;
  assign n48233 = n54170 & n48232;
  assign n48234 = n56594 & n27949;
  assign n48235 = n48233 & n48234;
  assign n48236 = n2454 & n3475;
  assign n48237 = n9210 & n28007;
  assign n48238 = n48236 & n48237;
  assign n48239 = n55142 & n48238;
  assign n48240 = n48232 & n48236;
  assign n48241 = n54170 & n56594;
  assign n48242 = n48240 & n48241;
  assign n48243 = n27949 & n48237;
  assign n48244 = n55142 & n48243;
  assign n48245 = n48242 & n48244;
  assign n48246 = n54170 & n55142;
  assign n48247 = n56594 & n48246;
  assign n48248 = n3639 & n9210;
  assign n48249 = n48236 & n48248;
  assign n48250 = ~n466 & ~n852;
  assign n48251 = n28007 & n48250;
  assign n48252 = ~n274 & ~n894;
  assign n48253 = n164 & n48252;
  assign n48254 = n48251 & n48253;
  assign n48255 = n48249 & n48254;
  assign n48256 = n48247 & n48255;
  assign n48257 = n48235 & n48239;
  assign n48258 = n53477 & n54128;
  assign n48259 = n54128 & n56587;
  assign n48260 = n53477 & n48259;
  assign n48261 = n56587 & n48258;
  assign n48262 = n59692 & n59693;
  assign n48263 = n54268 & n48262;
  assign n48264 = n54170 & n9210;
  assign n48265 = n55142 & n48264;
  assign n48266 = n56594 & n48265;
  assign n48267 = n3639 & n48266;
  assign n48268 = n56587 & n48267;
  assign n48269 = n2454 & n48268;
  assign n48270 = n53668 & n48269;
  assign n48271 = n54128 & n48270;
  assign n48272 = n3475 & n48271;
  assign n48273 = n53477 & n48272;
  assign n48274 = n54268 & n48273;
  assign n48275 = n164 & n48274;
  assign n48276 = ~n894 & n48275;
  assign n48277 = ~n659 & n48276;
  assign n48278 = ~n852 & n48277;
  assign n48279 = ~n274 & n48278;
  assign n48280 = ~n506 & n48279;
  assign n48281 = ~n466 & n48280;
  assign n48282 = n53668 & n48263;
  assign n48283 = pi2  & ~n59694;
  assign n48284 = ~pi2  & n59694;
  assign n48285 = ~n48283 & ~n48284;
  assign n48286 = n1576 & n40616;
  assign n48287 = n11215 & n39591;
  assign n48288 = n54403 & n39597;
  assign n48289 = n10564 & n39594;
  assign n48290 = ~n48288 & ~n48289;
  assign n48291 = ~n48287 & n48290;
  assign n48292 = ~n48286 & n48291;
  assign n48293 = ~n48285 & n48292;
  assign n48294 = ~n48284 & ~n48292;
  assign n48295 = ~n48283 & n48294;
  assign n48296 = ~n48283 & ~n48292;
  assign n48297 = ~n48284 & n48296;
  assign n48298 = n48285 & ~n48292;
  assign n48299 = ~n48292 & ~n59695;
  assign n48300 = ~n48283 & ~n59695;
  assign n48301 = ~n48283 & ~n48294;
  assign n48302 = ~n48284 & n59696;
  assign n48303 = ~n48299 & ~n48302;
  assign n48304 = ~n48293 & ~n59695;
  assign n48305 = n48229 & n59697;
  assign n48306 = ~n48229 & ~n59697;
  assign n48307 = ~n48305 & ~n48306;
  assign n48308 = n11279 & n41007;
  assign n48309 = n12584 & n39582;
  assign n48310 = n54410 & n39588;
  assign n48311 = n11267 & n39585;
  assign n48312 = ~n48310 & ~n48311;
  assign n48313 = ~n48309 & n48312;
  assign n48314 = ~n11279 & n48313;
  assign n48315 = ~n41007 & n48313;
  assign n48316 = ~n48314 & ~n48315;
  assign n48317 = ~n48308 & n48313;
  assign n48318 = pi29  & ~n59698;
  assign n48319 = ~pi29  & n59698;
  assign n48320 = ~n48318 & ~n48319;
  assign n48321 = n48307 & ~n48320;
  assign n48322 = ~n48307 & n48320;
  assign n48323 = ~n48321 & ~n48322;
  assign n48324 = ~n48228 & n48323;
  assign n48325 = n48228 & ~n48323;
  assign n48326 = ~n48324 & ~n48325;
  assign n48327 = n123 & n39976;
  assign n48328 = n128 & n39573;
  assign n48329 = n53444 & n39579;
  assign n48330 = n127 & n39576;
  assign n48331 = ~n48329 & ~n48330;
  assign n48332 = ~n48328 & n48331;
  assign n48333 = ~n48327 & n48332;
  assign n48334 = pi26  & ~n48333;
  assign n48335 = pi26  & ~n48334;
  assign n48336 = pi26  & n48333;
  assign n48337 = ~n48333 & ~n48334;
  assign n48338 = ~pi26  & ~n48333;
  assign n48339 = ~n59699 & ~n59700;
  assign n48340 = n48326 & ~n48339;
  assign n48341 = ~n48326 & n48339;
  assign n48342 = n48326 & ~n48340;
  assign n48343 = ~n48339 & ~n48340;
  assign n48344 = ~n48342 & ~n48343;
  assign n48345 = ~n48340 & ~n48341;
  assign n48346 = n48227 & n59701;
  assign n48347 = ~n48227 & ~n59701;
  assign n48348 = ~n48346 & ~n48347;
  assign n48349 = n90 & n41762;
  assign n48350 = n14236 & n39564;
  assign n48351 = n54667 & n39570;
  assign n48352 = n14210 & n39567;
  assign n48353 = ~n48351 & ~n48352;
  assign n48354 = ~n48350 & n48353;
  assign n48355 = ~n48349 & n48354;
  assign n48356 = pi23  & ~n48355;
  assign n48357 = pi23  & ~n48356;
  assign n48358 = pi23  & n48355;
  assign n48359 = ~n48355 & ~n48356;
  assign n48360 = ~pi23  & ~n48355;
  assign n48361 = ~n59702 & ~n59703;
  assign n48362 = ~n48348 & n48361;
  assign n48363 = n48348 & ~n48361;
  assign n48364 = n48348 & ~n48363;
  assign n48365 = ~n48361 & ~n48363;
  assign n48366 = ~n48364 & ~n48365;
  assign n48367 = ~n48362 & ~n48363;
  assign n48368 = n48226 & n59704;
  assign n48369 = ~n48226 & ~n59704;
  assign n48370 = ~n48368 & ~n48369;
  assign n48371 = n14413 & n42574;
  assign n48372 = n15921 & n39555;
  assign n48373 = n54719 & n39561;
  assign n48374 = n15901 & n39558;
  assign n48375 = ~n48373 & ~n48374;
  assign n48376 = ~n48372 & n48375;
  assign n48377 = ~n48371 & n48376;
  assign n48378 = pi20  & ~n48377;
  assign n48379 = pi20  & ~n48378;
  assign n48380 = pi20  & n48377;
  assign n48381 = ~n48377 & ~n48378;
  assign n48382 = ~pi20  & ~n48377;
  assign n48383 = ~n59705 & ~n59706;
  assign n48384 = n48370 & ~n48383;
  assign n48385 = ~n48370 & n48383;
  assign n48386 = n48370 & ~n48384;
  assign n48387 = ~n48383 & ~n48384;
  assign n48388 = ~n48386 & ~n48387;
  assign n48389 = ~n48384 & ~n48385;
  assign n48390 = n48225 & n59707;
  assign n48391 = ~n48225 & ~n59707;
  assign n48392 = ~n48390 & ~n48391;
  assign n48393 = n16079 & n43436;
  assign n48394 = n16696 & n39546;
  assign n48395 = n54886 & n39552;
  assign n48396 = n16676 & n39549;
  assign n48397 = ~n48395 & ~n48396;
  assign n48398 = ~n48394 & n48397;
  assign n48399 = ~n48393 & n48398;
  assign n48400 = pi17  & ~n48399;
  assign n48401 = pi17  & ~n48400;
  assign n48402 = pi17  & n48399;
  assign n48403 = ~n48399 & ~n48400;
  assign n48404 = ~pi17  & ~n48399;
  assign n48405 = ~n59708 & ~n59709;
  assign n48406 = ~n48392 & n48405;
  assign n48407 = n48392 & ~n48405;
  assign n48408 = n48392 & ~n48407;
  assign n48409 = ~n48405 & ~n48407;
  assign n48410 = ~n48408 & ~n48409;
  assign n48411 = ~n48406 & ~n48407;
  assign n48412 = n48224 & n59710;
  assign n48413 = ~n48224 & ~n59710;
  assign n48414 = ~n48412 & ~n48413;
  assign n48415 = n17265 & n39943;
  assign n48416 = n18588 & n39937;
  assign n48417 = n55041 & n39440;
  assign n48418 = n18556 & n39543;
  assign n48419 = ~n48417 & ~n48418;
  assign n48420 = ~n48416 & n48419;
  assign n48421 = ~n48415 & n48420;
  assign n48422 = pi14  & ~n48421;
  assign n48423 = pi14  & ~n48422;
  assign n48424 = pi14  & n48421;
  assign n48425 = ~n48421 & ~n48422;
  assign n48426 = ~pi14  & ~n48421;
  assign n48427 = ~n59711 & ~n59712;
  assign n48428 = n48414 & ~n48427;
  assign n48429 = ~n48414 & n48427;
  assign n48430 = n48414 & ~n48428;
  assign n48431 = ~n48427 & ~n48428;
  assign n48432 = ~n48430 & ~n48431;
  assign n48433 = ~n48428 & ~n48429;
  assign n48434 = n48223 & n59713;
  assign n48435 = ~n48223 & ~n59713;
  assign n48436 = ~n48434 & ~n48435;
  assign n48437 = n18846 & ~n59280;
  assign n48438 = n19541 & n44871;
  assign n48439 = n55247 & n44327;
  assign n48440 = n19509 & n44775;
  assign n48441 = ~n48439 & ~n48440;
  assign n48442 = ~n48438 & n48441;
  assign n48443 = ~n48437 & n48442;
  assign n48444 = pi11  & ~n48443;
  assign n48445 = pi11  & ~n48444;
  assign n48446 = pi11  & n48443;
  assign n48447 = ~n48443 & ~n48444;
  assign n48448 = ~pi11  & ~n48443;
  assign n48449 = ~n59714 & ~n59715;
  assign n48450 = ~n48436 & n48449;
  assign n48451 = n48436 & ~n48449;
  assign n48452 = n48436 & ~n48451;
  assign n48453 = ~n48449 & ~n48451;
  assign n48454 = ~n48452 & ~n48453;
  assign n48455 = ~n48450 & ~n48451;
  assign n48456 = n48222 & n59716;
  assign n48457 = ~n48222 & ~n59716;
  assign n48458 = ~n48456 & ~n48457;
  assign n48459 = n20085 & n46426;
  assign n48460 = n21269 & n46420;
  assign n48461 = n55472 & n44952;
  assign n48462 = n21237 & n46009;
  assign n48463 = ~n48461 & ~n48462;
  assign n48464 = ~n48460 & n48463;
  assign n48465 = ~n48459 & n48464;
  assign n48466 = pi8  & ~n48465;
  assign n48467 = pi8  & ~n48466;
  assign n48468 = pi8  & n48465;
  assign n48469 = ~n48465 & ~n48466;
  assign n48470 = ~pi8  & ~n48465;
  assign n48471 = ~n59717 & ~n59718;
  assign n48472 = n48458 & ~n48471;
  assign n48473 = ~n48458 & n48471;
  assign n48474 = n48458 & ~n48472;
  assign n48475 = ~n48471 & ~n48472;
  assign n48476 = ~n48474 & ~n48475;
  assign n48477 = ~n48472 & ~n48473;
  assign n48478 = n48221 & n59719;
  assign n48479 = ~n48221 & ~n59719;
  assign n48480 = ~n48478 & ~n48479;
  assign n48481 = n77 & ~n47526;
  assign n48482 = n21969 & n46788;
  assign n48483 = n23459 & n59503;
  assign n48484 = ~n48482 & ~n48483;
  assign n48485 = ~n48481 & n48484;
  assign n48486 = pi5  & ~n48485;
  assign n48487 = pi5  & ~n48486;
  assign n48488 = pi5  & n48485;
  assign n48489 = ~n48485 & ~n48486;
  assign n48490 = ~pi5  & ~n48485;
  assign n48491 = ~n59720 & ~n59721;
  assign n48492 = ~n48480 & n48491;
  assign n48493 = n48480 & ~n48491;
  assign n48494 = n48480 & ~n48493;
  assign n48495 = ~n48491 & ~n48493;
  assign n48496 = ~n48494 & ~n48495;
  assign n48497 = ~n48492 & ~n48493;
  assign n48498 = n48220 & n59722;
  assign n48499 = ~n48220 & ~n59722;
  assign n48500 = ~n48498 & ~n48499;
  assign n48501 = ~n48211 & ~n48215;
  assign n48502 = ~n48500 & n48501;
  assign n48503 = n48500 & ~n48501;
  assign n48504 = ~n48502 & ~n48503;
  assign n48505 = n48217 & n48504;
  assign n48506 = ~n48217 & ~n48504;
  assign po7  = ~n48505 & ~n48506;
  assign n48508 = n123 & ~n58759;
  assign n48509 = n128 & n39570;
  assign n48510 = n53444 & n39576;
  assign n48511 = n127 & n39573;
  assign n48512 = ~n48510 & ~n48511;
  assign n48513 = ~n48509 & n48512;
  assign n48514 = ~n48508 & n48513;
  assign n48515 = pi26  & ~n48514;
  assign n48516 = pi26  & ~n48515;
  assign n48517 = pi26  & n48514;
  assign n48518 = ~n48514 & ~n48515;
  assign n48519 = ~pi26  & ~n48514;
  assign n48520 = ~n59723 & ~n59724;
  assign n48521 = ~n48306 & ~n48321;
  assign n48522 = ~n269 & ~n622;
  assign n48523 = n257 & n48522;
  assign n48524 = n10240 & n48523;
  assign n48525 = n58859 & n48524;
  assign n48526 = n6530 & n7646;
  assign n48527 = n9155 & n11829;
  assign n48528 = n48526 & n48527;
  assign n48529 = n4381 & n4710;
  assign n48530 = n5377 & n5849;
  assign n48531 = n48529 & n48530;
  assign n48532 = n48528 & n48531;
  assign n48533 = ~n307 & ~n622;
  assign n48534 = ~n269 & ~n754;
  assign n48535 = ~n622 & ~n754;
  assign n48536 = ~n269 & ~n307;
  assign n48537 = n48535 & n48536;
  assign n48538 = n48533 & n48534;
  assign n48539 = n10240 & n59725;
  assign n48540 = n58859 & n48539;
  assign n48541 = n257 & n5377;
  assign n48542 = n48529 & n48541;
  assign n48543 = n48528 & n48542;
  assign n48544 = n48540 & n48543;
  assign n48545 = n424 & n7646;
  assign n48546 = n59725 & n48545;
  assign n48547 = n58859 & n48546;
  assign n48548 = n257 & n6530;
  assign n48549 = n48527 & n48548;
  assign n48550 = n2326 & n4381;
  assign n48551 = n4710 & n5377;
  assign n48552 = n48550 & n48551;
  assign n48553 = n48549 & n48552;
  assign n48554 = n48547 & n48553;
  assign n48555 = n48525 & n48532;
  assign n48556 = ~n108 & ~n751;
  assign n48557 = ~n751 & ~n1124;
  assign n48558 = ~n108 & n48557;
  assign n48559 = ~n1124 & n48556;
  assign n48560 = n749 & n59727;
  assign n48561 = n749 & n57071;
  assign n48562 = ~n1124 & n48561;
  assign n48563 = ~n108 & n48562;
  assign n48564 = ~n751 & n48563;
  assign n48565 = n57071 & n48560;
  assign n48566 = n53994 & n59728;
  assign n48567 = n59726 & n48566;
  assign n48568 = n54182 & n48567;
  assign n48569 = n257 & n58859;
  assign n48570 = n6530 & n48569;
  assign n48571 = n9155 & n48570;
  assign n48572 = n59728 & n48571;
  assign n48573 = n57065 & n48572;
  assign n48574 = n53994 & n48573;
  assign n48575 = n7646 & n48574;
  assign n48576 = n5377 & n48575;
  assign n48577 = n2326 & n48576;
  assign n48578 = n4710 & n48577;
  assign n48579 = n424 & n48578;
  assign n48580 = n54182 & n48579;
  assign n48581 = n11829 & n48580;
  assign n48582 = n4381 & n48581;
  assign n48583 = ~n307 & n48582;
  assign n48584 = ~n269 & n48583;
  assign n48585 = ~n754 & n48584;
  assign n48586 = ~n622 & n48585;
  assign n48587 = n57065 & n48568;
  assign n48588 = pi2  & ~n59729;
  assign n48589 = ~pi2  & n59729;
  assign n48590 = ~n48588 & ~n48589;
  assign n48591 = ~n59696 & ~n48589;
  assign n48592 = ~n48588 & n48591;
  assign n48593 = ~n59696 & n48590;
  assign n48594 = n59696 & ~n48590;
  assign n48595 = ~n59696 & ~n59730;
  assign n48596 = ~n48588 & ~n59730;
  assign n48597 = ~n48589 & n48596;
  assign n48598 = ~n48595 & ~n48597;
  assign n48599 = ~n59730 & ~n48594;
  assign n48600 = n1576 & ~n58585;
  assign n48601 = n11215 & n39588;
  assign n48602 = n54403 & n39594;
  assign n48603 = n10564 & n39591;
  assign n48604 = ~n48602 & ~n48603;
  assign n48605 = ~n48601 & n48604;
  assign n48606 = ~n48600 & n48605;
  assign n48607 = ~n59731 & ~n48606;
  assign n48608 = n59731 & n48606;
  assign n48609 = ~n59731 & ~n48607;
  assign n48610 = ~n59731 & n48606;
  assign n48611 = ~n48606 & ~n48607;
  assign n48612 = n59731 & ~n48606;
  assign n48613 = ~n59732 & ~n59733;
  assign n48614 = ~n48607 & ~n48608;
  assign n48615 = n48521 & n59734;
  assign n48616 = ~n48521 & ~n59734;
  assign n48617 = ~n48615 & ~n48616;
  assign n48618 = n11279 & ~n58657;
  assign n48619 = n12584 & n39579;
  assign n48620 = n54410 & n39585;
  assign n48621 = n11267 & n39582;
  assign n48622 = ~n48620 & ~n48621;
  assign n48623 = ~n48619 & n48622;
  assign n48624 = ~n48618 & n48623;
  assign n48625 = pi29  & ~n48624;
  assign n48626 = pi29  & ~n48625;
  assign n48627 = pi29  & n48624;
  assign n48628 = ~n48624 & ~n48625;
  assign n48629 = ~pi29  & ~n48624;
  assign n48630 = ~n59735 & ~n59736;
  assign n48631 = n48617 & ~n48630;
  assign n48632 = ~n48617 & n48630;
  assign n48633 = n48617 & ~n48631;
  assign n48634 = n48617 & n48630;
  assign n48635 = ~n48630 & ~n48631;
  assign n48636 = ~n48617 & ~n48630;
  assign n48637 = ~n59737 & ~n59738;
  assign n48638 = ~n48631 & ~n48632;
  assign n48639 = ~n48520 & ~n59739;
  assign n48640 = n48520 & n59739;
  assign n48641 = ~n59739 & ~n48639;
  assign n48642 = n48520 & ~n59739;
  assign n48643 = ~n48520 & ~n48639;
  assign n48644 = ~n48520 & n59739;
  assign n48645 = ~n59740 & ~n59741;
  assign n48646 = ~n48639 & ~n48640;
  assign n48647 = ~n48324 & n48339;
  assign n48648 = ~n48324 & ~n48340;
  assign n48649 = ~n48325 & ~n48647;
  assign n48650 = n59742 & n59743;
  assign n48651 = ~n59742 & ~n59743;
  assign n48652 = ~n48650 & ~n48651;
  assign n48653 = n90 & ~n58493;
  assign n48654 = n14236 & n39561;
  assign n48655 = n54667 & n39567;
  assign n48656 = n14210 & n39564;
  assign n48657 = ~n48655 & ~n48656;
  assign n48658 = ~n48654 & n48657;
  assign n48659 = ~n48653 & n48658;
  assign n48660 = pi23  & ~n48659;
  assign n48661 = pi23  & ~n48660;
  assign n48662 = pi23  & n48659;
  assign n48663 = ~n48659 & ~n48660;
  assign n48664 = ~pi23  & ~n48659;
  assign n48665 = ~n59744 & ~n59745;
  assign n48666 = n48652 & ~n48665;
  assign n48667 = ~n48652 & n48665;
  assign n48668 = n48652 & ~n48666;
  assign n48669 = ~n48665 & ~n48666;
  assign n48670 = ~n48668 & ~n48669;
  assign n48671 = ~n48666 & ~n48667;
  assign n48672 = ~n48347 & n48361;
  assign n48673 = ~n48347 & ~n48363;
  assign n48674 = ~n48346 & ~n48672;
  assign n48675 = n59746 & n59747;
  assign n48676 = ~n59746 & ~n59747;
  assign n48677 = ~n48675 & ~n48676;
  assign n48678 = n14413 & ~n58891;
  assign n48679 = n15921 & n39552;
  assign n48680 = n54719 & n39558;
  assign n48681 = n15901 & n39555;
  assign n48682 = ~n48680 & ~n48681;
  assign n48683 = ~n48679 & n48682;
  assign n48684 = ~n48678 & n48683;
  assign n48685 = pi20  & ~n48684;
  assign n48686 = pi20  & ~n48685;
  assign n48687 = pi20  & n48684;
  assign n48688 = ~n48684 & ~n48685;
  assign n48689 = ~pi20  & ~n48684;
  assign n48690 = ~n59748 & ~n59749;
  assign n48691 = ~n48677 & n48690;
  assign n48692 = n48677 & ~n48690;
  assign n48693 = n48677 & ~n48692;
  assign n48694 = ~n48690 & ~n48692;
  assign n48695 = ~n48693 & ~n48694;
  assign n48696 = ~n48691 & ~n48692;
  assign n48697 = ~n48369 & n48383;
  assign n48698 = ~n48369 & ~n48384;
  assign n48699 = ~n48368 & ~n48697;
  assign n48700 = n59750 & n59751;
  assign n48701 = ~n59750 & ~n59751;
  assign n48702 = ~n48700 & ~n48701;
  assign n48703 = n16079 & ~n59050;
  assign n48704 = n16696 & n39440;
  assign n48705 = n54886 & n39549;
  assign n48706 = n16676 & n39546;
  assign n48707 = ~n48705 & ~n48706;
  assign n48708 = ~n48704 & n48707;
  assign n48709 = ~n48703 & n48708;
  assign n48710 = pi17  & ~n48709;
  assign n48711 = pi17  & ~n48710;
  assign n48712 = pi17  & n48709;
  assign n48713 = ~n48709 & ~n48710;
  assign n48714 = ~pi17  & ~n48709;
  assign n48715 = ~n59752 & ~n59753;
  assign n48716 = n48702 & ~n48715;
  assign n48717 = ~n48702 & n48715;
  assign n48718 = n48702 & ~n48716;
  assign n48719 = ~n48715 & ~n48716;
  assign n48720 = ~n48718 & ~n48719;
  assign n48721 = ~n48716 & ~n48717;
  assign n48722 = ~n48391 & n48405;
  assign n48723 = ~n48391 & ~n48407;
  assign n48724 = ~n48390 & ~n48722;
  assign n48725 = n59754 & n59755;
  assign n48726 = ~n59754 & ~n59755;
  assign n48727 = ~n48725 & ~n48726;
  assign n48728 = n17265 & ~n59184;
  assign n48729 = n18588 & n44327;
  assign n48730 = n55041 & n39543;
  assign n48731 = n18556 & n39937;
  assign n48732 = ~n48730 & ~n48731;
  assign n48733 = ~n48729 & n48732;
  assign n48734 = ~n48728 & n48733;
  assign n48735 = pi14  & ~n48734;
  assign n48736 = pi14  & ~n48735;
  assign n48737 = pi14  & n48734;
  assign n48738 = ~n48734 & ~n48735;
  assign n48739 = ~pi14  & ~n48734;
  assign n48740 = ~n59756 & ~n59757;
  assign n48741 = ~n48727 & n48740;
  assign n48742 = n48727 & ~n48740;
  assign n48743 = n48727 & ~n48742;
  assign n48744 = ~n48740 & ~n48742;
  assign n48745 = ~n48743 & ~n48744;
  assign n48746 = ~n48741 & ~n48742;
  assign n48747 = ~n48413 & n48427;
  assign n48748 = ~n48413 & ~n48428;
  assign n48749 = ~n48412 & ~n48747;
  assign n48750 = n59758 & n59759;
  assign n48751 = ~n59758 & ~n59759;
  assign n48752 = ~n48750 & ~n48751;
  assign n48753 = n18846 & ~n59275;
  assign n48754 = n19541 & n44952;
  assign n48755 = n55247 & n44775;
  assign n48756 = n19509 & n44871;
  assign n48757 = ~n48755 & ~n48756;
  assign n48758 = ~n48754 & n48757;
  assign n48759 = ~n48753 & n48758;
  assign n48760 = pi11  & ~n48759;
  assign n48761 = pi11  & ~n48760;
  assign n48762 = pi11  & n48759;
  assign n48763 = ~n48759 & ~n48760;
  assign n48764 = ~pi11  & ~n48759;
  assign n48765 = ~n59760 & ~n59761;
  assign n48766 = n48752 & ~n48765;
  assign n48767 = ~n48752 & n48765;
  assign n48768 = n48752 & ~n48766;
  assign n48769 = ~n48765 & ~n48766;
  assign n48770 = ~n48768 & ~n48769;
  assign n48771 = ~n48766 & ~n48767;
  assign n48772 = ~n48435 & n48449;
  assign n48773 = ~n48435 & ~n48451;
  assign n48774 = ~n48434 & ~n48772;
  assign n48775 = n59762 & n59763;
  assign n48776 = ~n59762 & ~n59763;
  assign n48777 = ~n48775 & ~n48776;
  assign n48778 = n20085 & n46805;
  assign n48779 = n21269 & n46788;
  assign n48780 = n55472 & n46009;
  assign n48781 = n21237 & n46420;
  assign n48782 = ~n48780 & ~n48781;
  assign n48783 = ~n48779 & n48782;
  assign n48784 = ~n48778 & n48783;
  assign n48785 = pi8  & ~n48784;
  assign n48786 = pi8  & ~n48785;
  assign n48787 = pi8  & n48784;
  assign n48788 = ~n48784 & ~n48785;
  assign n48789 = ~pi8  & ~n48784;
  assign n48790 = ~n59764 & ~n59765;
  assign n48791 = ~n48777 & n48790;
  assign n48792 = n48777 & ~n48790;
  assign n48793 = n48777 & ~n48792;
  assign n48794 = ~n48790 & ~n48792;
  assign n48795 = ~n48793 & ~n48794;
  assign n48796 = ~n48791 & ~n48792;
  assign n48797 = ~n48457 & n48471;
  assign n48798 = ~n48457 & ~n48472;
  assign n48799 = ~n48456 & ~n48797;
  assign n48800 = n59766 & n59767;
  assign n48801 = ~n59766 & ~n59767;
  assign n48802 = ~n48800 & ~n48801;
  assign n48803 = n21969 & n59503;
  assign n48804 = pi5  & n48803;
  assign n48805 = pi5  & ~n48804;
  assign n48806 = pi5  & ~n48803;
  assign n48807 = n48803 & ~n48804;
  assign n48808 = ~pi5  & n48803;
  assign n48809 = ~n59768 & ~n59769;
  assign n48810 = n48802 & ~n48809;
  assign n48811 = ~n48802 & n48809;
  assign n48812 = n48802 & ~n48810;
  assign n48813 = ~n48809 & ~n48810;
  assign n48814 = ~n48812 & ~n48813;
  assign n48815 = ~n48810 & ~n48811;
  assign n48816 = ~n48479 & n48491;
  assign n48817 = ~n48479 & ~n48493;
  assign n48818 = ~n48478 & ~n48816;
  assign n48819 = n59770 & n59771;
  assign n48820 = ~n59770 & ~n59771;
  assign n48821 = ~n48819 & ~n48820;
  assign n48822 = ~n48499 & ~n48503;
  assign n48823 = ~n48821 & n48822;
  assign n48824 = n48821 & ~n48822;
  assign n48825 = ~n48823 & ~n48824;
  assign n48826 = n48505 & n48825;
  assign n48827 = ~n48505 & ~n48825;
  assign po8  = ~n48826 & ~n48827;
  assign n48829 = ~n48776 & n48790;
  assign n48830 = ~n48776 & ~n48792;
  assign n48831 = ~n48775 & ~n48829;
  assign n48832 = pi5  & ~n59772;
  assign n48833 = ~pi5  & n59772;
  assign n48834 = ~n48832 & ~n48833;
  assign n48835 = ~n48631 & ~n48639;
  assign n48836 = n123 & ~n58766;
  assign n48837 = n128 & n39567;
  assign n48838 = n53444 & n39573;
  assign n48839 = n127 & n39570;
  assign n48840 = ~n48838 & ~n48839;
  assign n48841 = ~n48837 & n48840;
  assign n48842 = ~n48836 & n48841;
  assign n48843 = pi26  & ~n48842;
  assign n48844 = pi26  & ~n48843;
  assign n48845 = pi26  & n48842;
  assign n48846 = ~n48842 & ~n48843;
  assign n48847 = ~pi26  & ~n48842;
  assign n48848 = ~n59773 & ~n59774;
  assign n48849 = ~n48607 & ~n48616;
  assign n48850 = n1128 & n5733;
  assign n48851 = n9211 & n10301;
  assign n48852 = n48850 & n48851;
  assign n48853 = n54438 & n48852;
  assign n48854 = n56904 & n48853;
  assign n48855 = ~n901 & ~n1492;
  assign n48856 = ~n901 & ~n1471;
  assign n48857 = ~n1492 & n48856;
  assign n48858 = ~n1471 & n48855;
  assign n48859 = ~n354 & ~n628;
  assign n48860 = n1035 & n48859;
  assign n48861 = ~n628 & n48855;
  assign n48862 = ~n354 & ~n1471;
  assign n48863 = n1035 & n48862;
  assign n48864 = n48861 & n48863;
  assign n48865 = ~n354 & n48855;
  assign n48866 = ~n628 & ~n1471;
  assign n48867 = n1035 & n48866;
  assign n48868 = n48865 & n48867;
  assign n48869 = n59775 & n48860;
  assign n48870 = n9331 & n59776;
  assign n48871 = n53842 & n48870;
  assign n48872 = n54817 & n48870;
  assign n48873 = n53842 & n48872;
  assign n48874 = n54817 & n48871;
  assign n48875 = n48854 & n59777;
  assign n48876 = n54187 & n48875;
  assign n48877 = n9211 & n56904;
  assign n48878 = n10301 & n48877;
  assign n48879 = n5733 & n48878;
  assign n48880 = n54438 & n48879;
  assign n48881 = n54817 & n48880;
  assign n48882 = n53872 & n48881;
  assign n48883 = n53842 & n48882;
  assign n48884 = n1128 & n48883;
  assign n48885 = n9331 & n48884;
  assign n48886 = n1035 & n48885;
  assign n48887 = n54187 & n48886;
  assign n48888 = ~n1471 & n48887;
  assign n48889 = ~n628 & n48888;
  assign n48890 = ~n901 & n48889;
  assign n48891 = ~n1492 & n48890;
  assign n48892 = ~n354 & n48891;
  assign n48893 = n53872 & n48876;
  assign n48894 = pi2  & ~n59778;
  assign n48895 = ~pi2  & n59778;
  assign n48896 = ~n48894 & ~n48895;
  assign n48897 = ~n48596 & ~n48895;
  assign n48898 = ~n48894 & n48897;
  assign n48899 = ~n48596 & n48896;
  assign n48900 = n48596 & ~n48896;
  assign n48901 = ~n48596 & ~n59779;
  assign n48902 = ~n48894 & ~n59779;
  assign n48903 = ~n48895 & n48902;
  assign n48904 = ~n48901 & ~n48903;
  assign n48905 = ~n59779 & ~n48900;
  assign n48906 = n1576 & ~n58583;
  assign n48907 = n11215 & n39585;
  assign n48908 = n54403 & n39591;
  assign n48909 = n10564 & n39588;
  assign n48910 = ~n48908 & ~n48909;
  assign n48911 = ~n48907 & n48910;
  assign n48912 = ~n48906 & n48911;
  assign n48913 = ~n59780 & ~n48912;
  assign n48914 = n59780 & n48912;
  assign n48915 = ~n59780 & ~n48913;
  assign n48916 = ~n59780 & n48912;
  assign n48917 = ~n48912 & ~n48913;
  assign n48918 = n59780 & ~n48912;
  assign n48919 = ~n59781 & ~n59782;
  assign n48920 = ~n48913 & ~n48914;
  assign n48921 = n48849 & n59783;
  assign n48922 = ~n48849 & ~n59783;
  assign n48923 = ~n48921 & ~n48922;
  assign n48924 = n11279 & ~n58653;
  assign n48925 = n12584 & n39576;
  assign n48926 = n54410 & n39582;
  assign n48927 = n11267 & n39579;
  assign n48928 = ~n48926 & ~n48927;
  assign n48929 = ~n48925 & n48928;
  assign n48930 = ~n48924 & n48929;
  assign n48931 = pi29  & ~n48930;
  assign n48932 = pi29  & ~n48931;
  assign n48933 = pi29  & n48930;
  assign n48934 = ~n48930 & ~n48931;
  assign n48935 = ~pi29  & ~n48930;
  assign n48936 = ~n59784 & ~n59785;
  assign n48937 = n48923 & ~n48936;
  assign n48938 = ~n48923 & n48936;
  assign n48939 = n48923 & ~n48937;
  assign n48940 = n48923 & n48936;
  assign n48941 = ~n48936 & ~n48937;
  assign n48942 = ~n48923 & ~n48936;
  assign n48943 = ~n59786 & ~n59787;
  assign n48944 = ~n48937 & ~n48938;
  assign n48945 = ~n48848 & ~n59788;
  assign n48946 = n48848 & n59788;
  assign n48947 = ~n59788 & ~n48945;
  assign n48948 = n48848 & ~n59788;
  assign n48949 = ~n48848 & ~n48945;
  assign n48950 = ~n48848 & n59788;
  assign n48951 = ~n59789 & ~n59790;
  assign n48952 = ~n48945 & ~n48946;
  assign n48953 = n48835 & n59791;
  assign n48954 = ~n48835 & ~n59791;
  assign n48955 = ~n48953 & ~n48954;
  assign n48956 = n90 & ~n58849;
  assign n48957 = n14236 & n39558;
  assign n48958 = n54667 & n39564;
  assign n48959 = n14210 & n39561;
  assign n48960 = ~n48958 & ~n48959;
  assign n48961 = ~n48957 & n48960;
  assign n48962 = ~n48956 & n48961;
  assign n48963 = pi23  & ~n48962;
  assign n48964 = pi23  & ~n48963;
  assign n48965 = pi23  & n48962;
  assign n48966 = ~n48962 & ~n48963;
  assign n48967 = ~pi23  & ~n48962;
  assign n48968 = ~n59792 & ~n59793;
  assign n48969 = n48955 & ~n48968;
  assign n48970 = ~n48955 & n48968;
  assign n48971 = n48955 & ~n48969;
  assign n48972 = ~n48968 & ~n48969;
  assign n48973 = ~n48971 & ~n48972;
  assign n48974 = ~n48969 & ~n48970;
  assign n48975 = ~n48651 & n48665;
  assign n48976 = ~n48651 & ~n48666;
  assign n48977 = ~n48650 & ~n48975;
  assign n48978 = n59794 & n59795;
  assign n48979 = ~n59794 & ~n59795;
  assign n48980 = ~n48978 & ~n48979;
  assign n48981 = n14413 & ~n58889;
  assign n48982 = n15921 & n39549;
  assign n48983 = n54719 & n39555;
  assign n48984 = n15901 & n39552;
  assign n48985 = ~n48983 & ~n48984;
  assign n48986 = ~n48982 & n48985;
  assign n48987 = ~n48981 & n48986;
  assign n48988 = pi20  & ~n48987;
  assign n48989 = pi20  & ~n48988;
  assign n48990 = pi20  & n48987;
  assign n48991 = ~n48987 & ~n48988;
  assign n48992 = ~pi20  & ~n48987;
  assign n48993 = ~n59796 & ~n59797;
  assign n48994 = ~n48980 & n48993;
  assign n48995 = n48980 & ~n48993;
  assign n48996 = n48980 & ~n48995;
  assign n48997 = ~n48993 & ~n48995;
  assign n48998 = ~n48996 & ~n48997;
  assign n48999 = ~n48994 & ~n48995;
  assign n49000 = ~n48676 & n48690;
  assign n49001 = ~n48676 & ~n48692;
  assign n49002 = ~n48675 & ~n49000;
  assign n49003 = n59798 & n59799;
  assign n49004 = ~n59798 & ~n59799;
  assign n49005 = ~n49003 & ~n49004;
  assign n49006 = n16079 & ~n59044;
  assign n49007 = n16696 & n39543;
  assign n49008 = n54886 & n39546;
  assign n49009 = n16676 & n39440;
  assign n49010 = ~n49008 & ~n49009;
  assign n49011 = ~n49007 & n49010;
  assign n49012 = ~n49006 & n49011;
  assign n49013 = pi17  & ~n49012;
  assign n49014 = pi17  & ~n49013;
  assign n49015 = pi17  & n49012;
  assign n49016 = ~n49012 & ~n49013;
  assign n49017 = ~pi17  & ~n49012;
  assign n49018 = ~n59800 & ~n59801;
  assign n49019 = n49005 & ~n49018;
  assign n49020 = ~n49005 & n49018;
  assign n49021 = n49005 & ~n49019;
  assign n49022 = ~n49018 & ~n49019;
  assign n49023 = ~n49021 & ~n49022;
  assign n49024 = ~n49019 & ~n49020;
  assign n49025 = ~n48701 & n48715;
  assign n49026 = ~n48701 & ~n48716;
  assign n49027 = ~n48700 & ~n49025;
  assign n49028 = n59802 & n59803;
  assign n49029 = ~n59802 & ~n59803;
  assign n49030 = ~n49028 & ~n49029;
  assign n49031 = n17265 & ~n59282;
  assign n49032 = n18588 & n44775;
  assign n49033 = n55041 & n39937;
  assign n49034 = n18556 & n44327;
  assign n49035 = ~n49033 & ~n49034;
  assign n49036 = ~n49032 & n49035;
  assign n49037 = ~n49031 & n49036;
  assign n49038 = pi14  & ~n49037;
  assign n49039 = pi14  & ~n49038;
  assign n49040 = pi14  & n49037;
  assign n49041 = ~n49037 & ~n49038;
  assign n49042 = ~pi14  & ~n49037;
  assign n49043 = ~n59804 & ~n59805;
  assign n49044 = ~n49030 & n49043;
  assign n49045 = n49030 & ~n49043;
  assign n49046 = n49030 & ~n49045;
  assign n49047 = ~n49043 & ~n49045;
  assign n49048 = ~n49046 & ~n49047;
  assign n49049 = ~n49044 & ~n49045;
  assign n49050 = ~n48726 & n48740;
  assign n49051 = ~n48726 & ~n48742;
  assign n49052 = ~n48725 & ~n49050;
  assign n49053 = n59806 & n59807;
  assign n49054 = ~n59806 & ~n59807;
  assign n49055 = ~n49053 & ~n49054;
  assign n49056 = n18846 & ~n59386;
  assign n49057 = n19541 & n46009;
  assign n49058 = n55247 & n44871;
  assign n49059 = n19509 & n44952;
  assign n49060 = ~n49058 & ~n49059;
  assign n49061 = ~n49057 & n49060;
  assign n49062 = ~n49056 & n49061;
  assign n49063 = pi11  & ~n49062;
  assign n49064 = pi11  & ~n49063;
  assign n49065 = pi11  & n49062;
  assign n49066 = ~n49062 & ~n49063;
  assign n49067 = ~pi11  & ~n49062;
  assign n49068 = ~n59808 & ~n59809;
  assign n49069 = n49055 & ~n49068;
  assign n49070 = ~n49055 & n49068;
  assign n49071 = n49055 & ~n49069;
  assign n49072 = ~n49068 & ~n49069;
  assign n49073 = ~n49071 & ~n49072;
  assign n49074 = ~n49069 & ~n49070;
  assign n49075 = ~n48751 & n48765;
  assign n49076 = ~n48751 & ~n48766;
  assign n49077 = ~n48750 & ~n49075;
  assign n49078 = n59810 & n59811;
  assign n49079 = ~n59810 & ~n59811;
  assign n49080 = ~n49078 & ~n49079;
  assign n49081 = n20085 & ~n59554;
  assign n49082 = n21269 & n59503;
  assign n49083 = n55472 & n46420;
  assign n49084 = n21237 & n46788;
  assign n49085 = ~n49083 & ~n49084;
  assign n49086 = ~n49082 & n49085;
  assign n49087 = ~n49081 & n49086;
  assign n49088 = pi8  & ~n49087;
  assign n49089 = pi8  & ~n49088;
  assign n49090 = pi8  & n49087;
  assign n49091 = ~n49087 & ~n49088;
  assign n49092 = ~pi8  & ~n49087;
  assign n49093 = ~n59812 & ~n59813;
  assign n49094 = ~n49080 & n49093;
  assign n49095 = n49080 & ~n49093;
  assign n49096 = n49080 & ~n49095;
  assign n49097 = ~n49093 & ~n49095;
  assign n49098 = ~n49096 & ~n49097;
  assign n49099 = ~n49094 & ~n49095;
  assign n49100 = n48834 & ~n59814;
  assign n49101 = ~n48834 & n59814;
  assign n49102 = ~n59814 & ~n49100;
  assign n49103 = n48834 & ~n49100;
  assign n49104 = ~n49102 & ~n49103;
  assign n49105 = ~n49100 & ~n49101;
  assign n49106 = ~n48801 & n48809;
  assign n49107 = ~n48801 & ~n48810;
  assign n49108 = ~n48800 & ~n49106;
  assign n49109 = n59815 & n59816;
  assign n49110 = ~n59815 & ~n59816;
  assign n49111 = ~n49109 & ~n49110;
  assign n49112 = ~n48820 & ~n48824;
  assign n49113 = ~n49111 & n49112;
  assign n49114 = n49111 & ~n49112;
  assign n49115 = ~n49113 & ~n49114;
  assign n49116 = n48826 & n49115;
  assign n49117 = ~n48826 & ~n49115;
  assign po9  = ~n49116 & ~n49117;
  assign n49119 = ~n49110 & ~n49114;
  assign n49120 = ~n48937 & ~n48945;
  assign n49121 = n123 & n41762;
  assign n49122 = n128 & n39564;
  assign n49123 = n53444 & n39570;
  assign n49124 = n127 & n39567;
  assign n49125 = ~n49123 & ~n49124;
  assign n49126 = ~n49122 & n49125;
  assign n49127 = ~n49121 & n49126;
  assign n49128 = pi26  & ~n49127;
  assign n49129 = pi26  & ~n49128;
  assign n49130 = pi26  & n49127;
  assign n49131 = ~n49127 & ~n49128;
  assign n49132 = ~pi26  & ~n49127;
  assign n49133 = ~n59817 & ~n59818;
  assign n49134 = ~n48913 & ~n48922;
  assign n49135 = ~n750 & ~n777;
  assign n49136 = ~n1044 & ~n1478;
  assign n49137 = n49135 & n49136;
  assign n49138 = n648 & n850;
  assign n49139 = n49137 & n49138;
  assign n49140 = n14974 & n49139;
  assign n49141 = n2004 & n5952;
  assign n49142 = n9511 & n13737;
  assign n49143 = n49141 & n49142;
  assign n49144 = n56630 & n49143;
  assign n49145 = n648 & n2004;
  assign n49146 = n850 & n5952;
  assign n49147 = n49145 & n49146;
  assign n49148 = n49137 & n49147;
  assign n49149 = n1278 & n9511;
  assign n49150 = n13737 & n13912;
  assign n49151 = n49149 & n49150;
  assign n49152 = n56630 & n49151;
  assign n49153 = n49148 & n49152;
  assign n49154 = n49140 & n49144;
  assign n49155 = n58730 & n59819;
  assign n49156 = n54480 & n49155;
  assign n49157 = n54105 & n13737;
  assign n49158 = n5952 & n49157;
  assign n49159 = n13912 & n49158;
  assign n49160 = n2004 & n49159;
  assign n49161 = n648 & n49160;
  assign n49162 = n56630 & n49161;
  assign n49163 = n54480 & n49162;
  assign n49164 = n9511 & n49163;
  assign n49165 = n1278 & n49164;
  assign n49166 = n850 & n49165;
  assign n49167 = n58730 & n49166;
  assign n49168 = ~n1044 & n49167;
  assign n49169 = ~n1478 & n49168;
  assign n49170 = ~n777 & n49169;
  assign n49171 = ~n750 & n49170;
  assign n49172 = n54105 & n49156;
  assign n49173 = ~pi2  & ~n59820;
  assign n49174 = pi2  & n59820;
  assign n49175 = ~pi2  & n59820;
  assign n49176 = pi2  & ~n59820;
  assign n49177 = ~n49175 & ~n49176;
  assign n49178 = ~n49173 & ~n49174;
  assign n49179 = ~pi5  & ~n59821;
  assign n49180 = pi5  & n59821;
  assign n49181 = ~n59821 & ~n49179;
  assign n49182 = ~pi5  & ~n49179;
  assign n49183 = ~n49181 & ~n49182;
  assign n49184 = ~n49179 & ~n49180;
  assign n49185 = ~n48902 & ~n59822;
  assign n49186 = n48902 & n59822;
  assign n49187 = ~n48902 & n59822;
  assign n49188 = n48902 & ~n59822;
  assign n49189 = ~n49187 & ~n49188;
  assign n49190 = ~n49185 & ~n49186;
  assign n49191 = n1576 & n41007;
  assign n49192 = n11215 & n39582;
  assign n49193 = n54403 & n39588;
  assign n49194 = n10564 & n39585;
  assign n49195 = ~n49193 & ~n49194;
  assign n49196 = ~n49192 & n49195;
  assign n49197 = ~n49191 & n49196;
  assign n49198 = ~n59823 & ~n49197;
  assign n49199 = n59823 & n49197;
  assign n49200 = ~n49198 & ~n49199;
  assign n49201 = n49134 & ~n49200;
  assign n49202 = ~n49134 & n49200;
  assign n49203 = ~n49201 & ~n49202;
  assign n49204 = n11279 & n39976;
  assign n49205 = n12584 & n39573;
  assign n49206 = n54410 & n39579;
  assign n49207 = n11267 & n39576;
  assign n49208 = ~n49206 & ~n49207;
  assign n49209 = ~n49205 & n49208;
  assign n49210 = ~n49204 & n49209;
  assign n49211 = pi29  & ~n49210;
  assign n49212 = pi29  & ~n49211;
  assign n49213 = pi29  & n49210;
  assign n49214 = ~n49210 & ~n49211;
  assign n49215 = ~pi29  & ~n49210;
  assign n49216 = ~n59824 & ~n59825;
  assign n49217 = n49203 & ~n49216;
  assign n49218 = ~n49203 & n49216;
  assign n49219 = n49203 & ~n49217;
  assign n49220 = ~n49216 & ~n49217;
  assign n49221 = ~n49219 & ~n49220;
  assign n49222 = ~n49217 & ~n49218;
  assign n49223 = ~n49133 & ~n59826;
  assign n49224 = n49133 & n59826;
  assign n49225 = ~n59826 & ~n49223;
  assign n49226 = ~n49133 & ~n49223;
  assign n49227 = ~n49225 & ~n49226;
  assign n49228 = ~n49223 & ~n49224;
  assign n49229 = n49120 & n59827;
  assign n49230 = ~n49120 & ~n59827;
  assign n49231 = ~n49229 & ~n49230;
  assign n49232 = n90 & n42574;
  assign n49233 = n14236 & n39555;
  assign n49234 = n54667 & n39561;
  assign n49235 = n14210 & n39558;
  assign n49236 = ~n49234 & ~n49235;
  assign n49237 = ~n49233 & n49236;
  assign n49238 = ~n49232 & n49237;
  assign n49239 = pi23  & ~n49238;
  assign n49240 = pi23  & ~n49239;
  assign n49241 = pi23  & n49238;
  assign n49242 = ~n49238 & ~n49239;
  assign n49243 = ~pi23  & ~n49238;
  assign n49244 = ~n59828 & ~n59829;
  assign n49245 = n49231 & ~n49244;
  assign n49246 = ~n49231 & n49244;
  assign n49247 = n49231 & ~n49245;
  assign n49248 = n49231 & n49244;
  assign n49249 = ~n49244 & ~n49245;
  assign n49250 = ~n49231 & ~n49244;
  assign n49251 = ~n59830 & ~n59831;
  assign n49252 = ~n49245 & ~n49246;
  assign n49253 = ~n48954 & n48968;
  assign n49254 = ~n48954 & ~n48969;
  assign n49255 = ~n48953 & ~n49253;
  assign n49256 = n59832 & n59833;
  assign n49257 = ~n59832 & ~n59833;
  assign n49258 = ~n49256 & ~n49257;
  assign n49259 = n14413 & n43436;
  assign n49260 = n15921 & n39546;
  assign n49261 = n54719 & n39552;
  assign n49262 = n15901 & n39549;
  assign n49263 = ~n49261 & ~n49262;
  assign n49264 = ~n49260 & n49263;
  assign n49265 = ~n49259 & n49264;
  assign n49266 = pi20  & ~n49265;
  assign n49267 = pi20  & ~n49266;
  assign n49268 = pi20  & n49265;
  assign n49269 = ~n49265 & ~n49266;
  assign n49270 = ~pi20  & ~n49265;
  assign n49271 = ~n59834 & ~n59835;
  assign n49272 = n49258 & ~n49271;
  assign n49273 = ~n49258 & n49271;
  assign n49274 = n49258 & ~n49272;
  assign n49275 = n49258 & n49271;
  assign n49276 = ~n49271 & ~n49272;
  assign n49277 = ~n49258 & ~n49271;
  assign n49278 = ~n59836 & ~n59837;
  assign n49279 = ~n49272 & ~n49273;
  assign n49280 = ~n48979 & n48993;
  assign n49281 = ~n48979 & ~n48995;
  assign n49282 = ~n48978 & ~n49280;
  assign n49283 = n59838 & n59839;
  assign n49284 = ~n59838 & ~n59839;
  assign n49285 = ~n49283 & ~n49284;
  assign n49286 = n16079 & n39943;
  assign n49287 = n16696 & n39937;
  assign n49288 = n54886 & n39440;
  assign n49289 = n16676 & n39543;
  assign n49290 = ~n49288 & ~n49289;
  assign n49291 = ~n49287 & n49290;
  assign n49292 = ~n49286 & n49291;
  assign n49293 = pi17  & ~n49292;
  assign n49294 = pi17  & ~n49293;
  assign n49295 = pi17  & n49292;
  assign n49296 = ~n49292 & ~n49293;
  assign n49297 = ~pi17  & ~n49292;
  assign n49298 = ~n59840 & ~n59841;
  assign n49299 = n49285 & ~n49298;
  assign n49300 = ~n49285 & n49298;
  assign n49301 = n49285 & ~n49299;
  assign n49302 = n49285 & n49298;
  assign n49303 = ~n49298 & ~n49299;
  assign n49304 = ~n49285 & ~n49298;
  assign n49305 = ~n59842 & ~n59843;
  assign n49306 = ~n49299 & ~n49300;
  assign n49307 = ~n49004 & n49018;
  assign n49308 = ~n49004 & ~n49019;
  assign n49309 = ~n49003 & ~n49307;
  assign n49310 = n59844 & n59845;
  assign n49311 = ~n59844 & ~n59845;
  assign n49312 = ~n49310 & ~n49311;
  assign n49313 = n17265 & ~n59280;
  assign n49314 = n18588 & n44871;
  assign n49315 = n55041 & n44327;
  assign n49316 = n18556 & n44775;
  assign n49317 = ~n49315 & ~n49316;
  assign n49318 = ~n49314 & n49317;
  assign n49319 = ~n49313 & n49318;
  assign n49320 = pi14  & ~n49319;
  assign n49321 = pi14  & ~n49320;
  assign n49322 = pi14  & n49319;
  assign n49323 = ~n49319 & ~n49320;
  assign n49324 = ~pi14  & ~n49319;
  assign n49325 = ~n59846 & ~n59847;
  assign n49326 = ~n49029 & n49043;
  assign n49327 = ~n49029 & ~n49045;
  assign n49328 = ~n49028 & ~n49326;
  assign n49329 = ~n49325 & ~n59848;
  assign n49330 = n49325 & n59848;
  assign n49331 = ~n59848 & ~n49329;
  assign n49332 = n49325 & ~n59848;
  assign n49333 = ~n49325 & ~n49329;
  assign n49334 = ~n49325 & n59848;
  assign n49335 = ~n59849 & ~n59850;
  assign n49336 = ~n49329 & ~n49330;
  assign n49337 = ~n49312 & n59851;
  assign n49338 = n49312 & ~n59851;
  assign n49339 = ~n49337 & ~n49338;
  assign n49340 = n18846 & n46426;
  assign n49341 = n19541 & n46420;
  assign n49342 = n55247 & n44952;
  assign n49343 = n19509 & n46009;
  assign n49344 = ~n49342 & ~n49343;
  assign n49345 = ~n49341 & n49344;
  assign n49346 = ~n49340 & n49345;
  assign n49347 = pi11  & ~n49346;
  assign n49348 = pi11  & ~n49347;
  assign n49349 = pi11  & n49346;
  assign n49350 = ~n49346 & ~n49347;
  assign n49351 = ~pi11  & ~n49346;
  assign n49352 = ~n59852 & ~n59853;
  assign n49353 = n49339 & ~n49352;
  assign n49354 = ~n49339 & n49352;
  assign n49355 = n49339 & ~n49353;
  assign n49356 = n49339 & n49352;
  assign n49357 = ~n49352 & ~n49353;
  assign n49358 = ~n49339 & ~n49352;
  assign n49359 = ~n59854 & ~n59855;
  assign n49360 = ~n49353 & ~n49354;
  assign n49361 = ~n49054 & n49068;
  assign n49362 = ~n49054 & ~n49069;
  assign n49363 = ~n49053 & ~n49361;
  assign n49364 = n59856 & n59857;
  assign n49365 = ~n59856 & ~n59857;
  assign n49366 = ~n49364 & ~n49365;
  assign n49367 = n20085 & ~n47526;
  assign n49368 = n55472 & n46788;
  assign n49369 = n21237 & n59503;
  assign n49370 = ~n49368 & ~n49369;
  assign n49371 = ~n49367 & n49370;
  assign n49372 = pi8  & ~n49371;
  assign n49373 = pi8  & ~n49372;
  assign n49374 = pi8  & n49371;
  assign n49375 = ~n49371 & ~n49372;
  assign n49376 = ~pi8  & ~n49371;
  assign n49377 = ~n59858 & ~n59859;
  assign n49378 = ~n49079 & n49093;
  assign n49379 = ~n49079 & ~n49095;
  assign n49380 = ~n49078 & ~n49378;
  assign n49381 = ~n49377 & ~n59860;
  assign n49382 = n49377 & n59860;
  assign n49383 = ~n59860 & ~n49381;
  assign n49384 = n49377 & ~n59860;
  assign n49385 = ~n49377 & ~n49381;
  assign n49386 = ~n49377 & n59860;
  assign n49387 = ~n59861 & ~n59862;
  assign n49388 = ~n49381 & ~n49382;
  assign n49389 = ~n49366 & n59863;
  assign n49390 = n49366 & ~n59863;
  assign n49391 = ~n49389 & ~n49390;
  assign n49392 = ~n48832 & n59814;
  assign n49393 = ~n48832 & ~n49100;
  assign n49394 = ~n48833 & ~n49392;
  assign n49395 = n49391 & ~n59864;
  assign n49396 = ~n49391 & n59864;
  assign n49397 = ~n49395 & ~n49396;
  assign n49398 = ~n49119 & n49397;
  assign n49399 = n49119 & ~n49397;
  assign n49400 = ~n49398 & ~n49399;
  assign n49401 = ~n49116 & ~n49400;
  assign n49402 = n49116 & n49400;
  assign po10  = ~n49401 & ~n49402;
  assign n49404 = ~n49395 & ~n49398;
  assign n49405 = ~n49381 & ~n49390;
  assign n49406 = ~n49353 & ~n49365;
  assign n49407 = n18846 & n46805;
  assign n49408 = n19541 & n46788;
  assign n49409 = n55247 & n46009;
  assign n49410 = n19509 & n46420;
  assign n49411 = ~n49409 & ~n49410;
  assign n49412 = ~n49408 & n49411;
  assign n49413 = ~n49407 & n49412;
  assign n49414 = pi11  & ~n49413;
  assign n49415 = pi11  & ~n49414;
  assign n49416 = pi11  & n49413;
  assign n49417 = ~n49413 & ~n49414;
  assign n49418 = ~pi11  & ~n49413;
  assign n49419 = ~n59865 & ~n59866;
  assign n49420 = ~n49329 & ~n49338;
  assign n49421 = ~n49299 & ~n49311;
  assign n49422 = ~n49272 & ~n49284;
  assign n49423 = ~n49245 & ~n49257;
  assign n49424 = ~n49223 & ~n49230;
  assign n49425 = ~n49185 & ~n49198;
  assign n49426 = ~n49173 & ~n49179;
  assign n49427 = n5377 & n6300;
  assign n49428 = n6481 & n49427;
  assign n49429 = n54993 & n49428;
  assign n49430 = n55141 & n49429;
  assign n49431 = ~n141 & ~n416;
  assign n49432 = n2693 & n49431;
  assign n49433 = n2976 & n4833;
  assign n49434 = n49432 & n49433;
  assign n49435 = n53967 & n49434;
  assign n49436 = n53759 & n49435;
  assign n49437 = n6300 & n54993;
  assign n49438 = n53967 & n49437;
  assign n49439 = n6481 & n49438;
  assign n49440 = n55141 & n49439;
  assign n49441 = n4833 & n49440;
  assign n49442 = n53759 & n49441;
  assign n49443 = n5377 & n49442;
  assign n49444 = n2693 & n49443;
  assign n49445 = ~n416 & n49444;
  assign n49446 = ~n307 & n49445;
  assign n49447 = ~n141 & n49446;
  assign n49448 = ~n402 & n49447;
  assign n49449 = n2693 & n6300;
  assign n49450 = n6481 & n49449;
  assign n49451 = n54993 & n49450;
  assign n49452 = n55141 & n49451;
  assign n49453 = ~n307 & ~n416;
  assign n49454 = ~n141 & ~n402;
  assign n49455 = n49453 & n49454;
  assign n49456 = n4833 & n5377;
  assign n49457 = n49455 & n49456;
  assign n49458 = n53967 & n49457;
  assign n49459 = n53759 & n49458;
  assign n49460 = n49452 & n49459;
  assign n49461 = n49430 & n49436;
  assign n49462 = n882 & n4013;
  assign n49463 = n11990 & n12286;
  assign n49464 = n49462 & n49463;
  assign n49465 = n53855 & n49464;
  assign n49466 = n55134 & n49465;
  assign n49467 = ~n585 & ~n628;
  assign n49468 = n3776 & n49467;
  assign n49469 = n4026 & n4083;
  assign n49470 = n49468 & n49469;
  assign n49471 = ~n415 & ~n499;
  assign n49472 = ~n830 & n49471;
  assign n49473 = n54339 & n49472;
  assign n49474 = ~n499 & ~n628;
  assign n49475 = n3776 & n49474;
  assign n49476 = n49469 & n49475;
  assign n49477 = ~n415 & ~n585;
  assign n49478 = ~n830 & n49477;
  assign n49479 = n54339 & n49478;
  assign n49480 = n49476 & n49479;
  assign n49481 = n49470 & n49473;
  assign n49482 = n54028 & n59868;
  assign n49483 = n882 & n4083;
  assign n49484 = n49463 & n49483;
  assign n49485 = n53855 & n49484;
  assign n49486 = n55134 & n49485;
  assign n49487 = ~n499 & ~n830;
  assign n49488 = n3776 & n49487;
  assign n49489 = n4013 & n4026;
  assign n49490 = n49488 & n49489;
  assign n49491 = ~n628 & n49477;
  assign n49492 = n54339 & n49491;
  assign n49493 = n49490 & n49492;
  assign n49494 = n54028 & n49493;
  assign n49495 = n49486 & n49494;
  assign n49496 = n882 & n3776;
  assign n49497 = n4013 & n12286;
  assign n49498 = n49496 & n49497;
  assign n49499 = n53855 & n49498;
  assign n49500 = n55134 & n49499;
  assign n49501 = ~n415 & ~n628;
  assign n49502 = ~n585 & ~n830;
  assign n49503 = n49501 & n49502;
  assign n49504 = n49469 & n49503;
  assign n49505 = ~n499 & n11990;
  assign n49506 = n54339 & n49505;
  assign n49507 = n49504 & n49506;
  assign n49508 = n54028 & n49507;
  assign n49509 = n49500 & n49508;
  assign n49510 = n49466 & n49482;
  assign n49511 = n59867 & n59869;
  assign n49512 = n12286 & n49462;
  assign n49513 = n55134 & n49512;
  assign n49514 = n59867 & n49513;
  assign n49515 = n54028 & n49514;
  assign n49516 = n54339 & n49515;
  assign n49517 = n53855 & n49516;
  assign n49518 = n53832 & n49517;
  assign n49519 = n4083 & n49518;
  assign n49520 = n4026 & n49519;
  assign n49521 = n3776 & n49520;
  assign n49522 = ~n628 & n49521;
  assign n49523 = ~n415 & n49522;
  assign n49524 = ~n310 & n49523;
  assign n49525 = ~n660 & n49524;
  assign n49526 = ~n830 & n49525;
  assign n49527 = ~n499 & n49526;
  assign n49528 = ~n585 & n49527;
  assign n49529 = n53832 & n49511;
  assign n49530 = ~n49426 & n59870;
  assign n49531 = n49426 & ~n59870;
  assign n49532 = ~n49530 & ~n49531;
  assign n49533 = n1576 & ~n58657;
  assign n49534 = n11215 & n39579;
  assign n49535 = n54403 & n39585;
  assign n49536 = n10564 & n39582;
  assign n49537 = ~n49535 & ~n49536;
  assign n49538 = ~n49534 & n49537;
  assign n49539 = ~n49533 & n49538;
  assign n49540 = n49532 & ~n49539;
  assign n49541 = ~n49532 & n49539;
  assign n49542 = ~n49539 & ~n49540;
  assign n49543 = n49532 & ~n49540;
  assign n49544 = ~n49542 & ~n49543;
  assign n49545 = ~n49540 & ~n49541;
  assign n49546 = n49425 & n59871;
  assign n49547 = ~n49425 & ~n59871;
  assign n49548 = ~n49546 & ~n49547;
  assign n49549 = n11279 & ~n58759;
  assign n49550 = n12584 & n39570;
  assign n49551 = n54410 & n39576;
  assign n49552 = n11267 & n39573;
  assign n49553 = ~n49551 & ~n49552;
  assign n49554 = ~n49550 & n49553;
  assign n49555 = ~n11279 & n49554;
  assign n49556 = n58759 & n49554;
  assign n49557 = ~n49555 & ~n49556;
  assign n49558 = ~n49549 & n49554;
  assign n49559 = pi29  & ~n59872;
  assign n49560 = ~pi29  & n59872;
  assign n49561 = ~n49559 & ~n49560;
  assign n49562 = n49548 & ~n49561;
  assign n49563 = ~n49548 & n49561;
  assign n49564 = ~n49562 & ~n49563;
  assign n49565 = ~n49202 & n49216;
  assign n49566 = ~n49202 & ~n49217;
  assign n49567 = ~n49201 & ~n49565;
  assign n49568 = n49564 & ~n59873;
  assign n49569 = ~n49564 & n59873;
  assign n49570 = ~n49568 & ~n49569;
  assign n49571 = n123 & ~n58493;
  assign n49572 = n128 & n39561;
  assign n49573 = n53444 & n39567;
  assign n49574 = n127 & n39564;
  assign n49575 = ~n49573 & ~n49574;
  assign n49576 = ~n49572 & n49575;
  assign n49577 = ~n49571 & n49576;
  assign n49578 = pi26  & ~n49577;
  assign n49579 = pi26  & ~n49578;
  assign n49580 = pi26  & n49577;
  assign n49581 = ~n49577 & ~n49578;
  assign n49582 = ~pi26  & ~n49577;
  assign n49583 = ~n59874 & ~n59875;
  assign n49584 = n49570 & ~n49583;
  assign n49585 = ~n49570 & n49583;
  assign n49586 = n49570 & ~n49584;
  assign n49587 = ~n49583 & ~n49584;
  assign n49588 = ~n49586 & ~n49587;
  assign n49589 = ~n49584 & ~n49585;
  assign n49590 = n49424 & n59876;
  assign n49591 = ~n49424 & ~n59876;
  assign n49592 = ~n49590 & ~n49591;
  assign n49593 = n90 & ~n58891;
  assign n49594 = n14236 & n39552;
  assign n49595 = n54667 & n39558;
  assign n49596 = n14210 & n39555;
  assign n49597 = ~n49595 & ~n49596;
  assign n49598 = ~n49594 & n49597;
  assign n49599 = ~n49593 & n49598;
  assign n49600 = pi23  & ~n49599;
  assign n49601 = pi23  & ~n49600;
  assign n49602 = pi23  & n49599;
  assign n49603 = ~n49599 & ~n49600;
  assign n49604 = ~pi23  & ~n49599;
  assign n49605 = ~n59877 & ~n59878;
  assign n49606 = ~n49592 & n49605;
  assign n49607 = n49592 & ~n49605;
  assign n49608 = n49592 & ~n49607;
  assign n49609 = ~n49605 & ~n49607;
  assign n49610 = ~n49608 & ~n49609;
  assign n49611 = ~n49606 & ~n49607;
  assign n49612 = n49423 & n59879;
  assign n49613 = ~n49423 & ~n59879;
  assign n49614 = ~n49612 & ~n49613;
  assign n49615 = n14413 & ~n59050;
  assign n49616 = n15921 & n39440;
  assign n49617 = n54719 & n39549;
  assign n49618 = n15901 & n39546;
  assign n49619 = ~n49617 & ~n49618;
  assign n49620 = ~n49616 & n49619;
  assign n49621 = ~n49615 & n49620;
  assign n49622 = pi20  & ~n49621;
  assign n49623 = pi20  & ~n49622;
  assign n49624 = pi20  & n49621;
  assign n49625 = ~n49621 & ~n49622;
  assign n49626 = ~pi20  & ~n49621;
  assign n49627 = ~n59880 & ~n59881;
  assign n49628 = n49614 & ~n49627;
  assign n49629 = ~n49614 & n49627;
  assign n49630 = n49614 & ~n49628;
  assign n49631 = ~n49627 & ~n49628;
  assign n49632 = ~n49630 & ~n49631;
  assign n49633 = ~n49628 & ~n49629;
  assign n49634 = n49422 & n59882;
  assign n49635 = ~n49422 & ~n59882;
  assign n49636 = ~n49634 & ~n49635;
  assign n49637 = n16079 & ~n59184;
  assign n49638 = n16696 & n44327;
  assign n49639 = n54886 & n39543;
  assign n49640 = n16676 & n39937;
  assign n49641 = ~n49639 & ~n49640;
  assign n49642 = ~n49638 & n49641;
  assign n49643 = ~n49637 & n49642;
  assign n49644 = pi17  & ~n49643;
  assign n49645 = pi17  & ~n49644;
  assign n49646 = pi17  & n49643;
  assign n49647 = ~n49643 & ~n49644;
  assign n49648 = ~pi17  & ~n49643;
  assign n49649 = ~n59883 & ~n59884;
  assign n49650 = ~n49636 & n49649;
  assign n49651 = n49636 & ~n49649;
  assign n49652 = n49636 & ~n49651;
  assign n49653 = ~n49649 & ~n49651;
  assign n49654 = ~n49652 & ~n49653;
  assign n49655 = ~n49650 & ~n49651;
  assign n49656 = n49421 & n59885;
  assign n49657 = ~n49421 & ~n59885;
  assign n49658 = ~n49656 & ~n49657;
  assign n49659 = n17265 & ~n59275;
  assign n49660 = n18588 & n44952;
  assign n49661 = n55041 & n44775;
  assign n49662 = n18556 & n44871;
  assign n49663 = ~n49661 & ~n49662;
  assign n49664 = ~n49660 & n49663;
  assign n49665 = ~n49659 & n49664;
  assign n49666 = pi14  & ~n49665;
  assign n49667 = pi14  & ~n49666;
  assign n49668 = pi14  & n49665;
  assign n49669 = ~n49665 & ~n49666;
  assign n49670 = ~pi14  & ~n49665;
  assign n49671 = ~n59886 & ~n59887;
  assign n49672 = n49658 & ~n49671;
  assign n49673 = ~n49658 & n49671;
  assign n49674 = n49658 & ~n49672;
  assign n49675 = ~n49671 & ~n49672;
  assign n49676 = ~n49674 & ~n49675;
  assign n49677 = ~n49672 & ~n49673;
  assign n49678 = ~n49420 & ~n59888;
  assign n49679 = n49420 & n59888;
  assign n49680 = ~n59888 & ~n49678;
  assign n49681 = n49420 & ~n59888;
  assign n49682 = ~n49420 & ~n49678;
  assign n49683 = ~n49420 & n59888;
  assign n49684 = ~n59889 & ~n59890;
  assign n49685 = ~n49678 & ~n49679;
  assign n49686 = ~n49419 & ~n59891;
  assign n49687 = n49419 & n59891;
  assign n49688 = ~n59891 & ~n49686;
  assign n49689 = ~n49419 & ~n49686;
  assign n49690 = ~n49688 & ~n49689;
  assign n49691 = ~n49686 & ~n49687;
  assign n49692 = n49406 & n59892;
  assign n49693 = ~n49406 & ~n59892;
  assign n49694 = ~n49692 & ~n49693;
  assign n49695 = n55472 & n59503;
  assign n49696 = pi8  & n49695;
  assign n49697 = pi8  & ~n49696;
  assign n49698 = pi8  & ~n49695;
  assign n49699 = n49695 & ~n49696;
  assign n49700 = ~pi8  & n49695;
  assign n49701 = ~n59893 & ~n59894;
  assign n49702 = n49694 & ~n49701;
  assign n49703 = ~n49694 & n49701;
  assign n49704 = n49694 & ~n49702;
  assign n49705 = ~n49701 & ~n49702;
  assign n49706 = ~n49704 & ~n49705;
  assign n49707 = ~n49702 & ~n49703;
  assign n49708 = ~n49405 & ~n59895;
  assign n49709 = n49405 & n59895;
  assign n49710 = ~n59895 & ~n49708;
  assign n49711 = ~n49405 & ~n49708;
  assign n49712 = ~n49710 & ~n49711;
  assign n49713 = ~n49708 & ~n49709;
  assign n49714 = n49404 & n59896;
  assign n49715 = ~n49404 & ~n59896;
  assign n49716 = ~n49714 & ~n49715;
  assign n49717 = n49402 & n49716;
  assign n49718 = ~n49402 & ~n49716;
  assign po11  = ~n49717 & ~n49718;
  assign n49720 = ~n49678 & ~n49686;
  assign n49721 = pi8  & ~n49720;
  assign n49722 = ~pi8  & n49720;
  assign n49723 = ~n49721 & ~n49722;
  assign n49724 = n123 & ~n58849;
  assign n49725 = n128 & n39558;
  assign n49726 = n53444 & n39564;
  assign n49727 = n127 & n39561;
  assign n49728 = ~n49726 & ~n49727;
  assign n49729 = ~n49725 & n49728;
  assign n49730 = ~n49724 & n49729;
  assign n49731 = pi26  & ~n49730;
  assign n49732 = pi26  & ~n49731;
  assign n49733 = pi26  & n49730;
  assign n49734 = ~n49730 & ~n49731;
  assign n49735 = ~pi26  & ~n49730;
  assign n49736 = ~n59897 & ~n59898;
  assign n49737 = ~n49547 & ~n49562;
  assign n49738 = ~n975 & ~n1234;
  assign n49739 = ~n1191 & n49738;
  assign n49740 = ~n258 & ~n748;
  assign n49741 = n3085 & n49740;
  assign n49742 = ~n975 & ~n1646;
  assign n49743 = ~n1191 & n49742;
  assign n49744 = n1541 & n49740;
  assign n49745 = n49743 & n49744;
  assign n49746 = n49739 & n49741;
  assign n49747 = n10952 & n13598;
  assign n49748 = n59899 & n49747;
  assign n49749 = n1458 & n9330;
  assign n49750 = n1458 & n9337;
  assign n49751 = n9330 & n49750;
  assign n49752 = n9337 & n49749;
  assign n49753 = n53901 & n59900;
  assign n49754 = ~n748 & ~n975;
  assign n49755 = ~n1191 & n49754;
  assign n49756 = ~n258 & ~n1646;
  assign n49757 = n9330 & n49756;
  assign n49758 = ~n748 & ~n1646;
  assign n49759 = ~n1191 & n49758;
  assign n49760 = ~n258 & ~n975;
  assign n49761 = n9330 & n49760;
  assign n49762 = n49759 & n49761;
  assign n49763 = n49755 & n49757;
  assign n49764 = n49747 & n59901;
  assign n49765 = n1541 & n49750;
  assign n49766 = n53901 & n49765;
  assign n49767 = n49764 & n49766;
  assign n49768 = n49748 & n49753;
  assign n49769 = n9330 & n10952;
  assign n49770 = n53901 & n49769;
  assign n49771 = n13598 & n49770;
  assign n49772 = n9337 & n49771;
  assign n49773 = n1541 & n49772;
  assign n49774 = n54242 & n49773;
  assign n49775 = n1458 & n49774;
  assign n49776 = ~n1191 & n49775;
  assign n49777 = ~n258 & n49776;
  assign n49778 = ~n748 & n49777;
  assign n49779 = ~n975 & n49778;
  assign n49780 = ~n1646 & n49779;
  assign n49781 = n54242 & n59902;
  assign n49782 = ~n1280 & ~n1881;
  assign n49783 = ~n901 & n49782;
  assign n49784 = ~n361 & ~n559;
  assign n49785 = n5660 & n49784;
  assign n49786 = ~n222 & ~n361;
  assign n49787 = ~n321 & ~n410;
  assign n49788 = ~n559 & ~n830;
  assign n49789 = n49787 & n49788;
  assign n49790 = n49786 & n49789;
  assign n49791 = n9981 & n49785;
  assign n49792 = ~n559 & ~n901;
  assign n49793 = ~n321 & n49792;
  assign n49794 = ~n222 & n49793;
  assign n49795 = ~n1280 & n49794;
  assign n49796 = ~n830 & n49795;
  assign n49797 = ~n361 & n49796;
  assign n49798 = ~n410 & n49797;
  assign n49799 = ~n1881 & n49798;
  assign n49800 = ~n410 & n49792;
  assign n49801 = ~n361 & ~n1881;
  assign n49802 = ~n222 & ~n321;
  assign n49803 = ~n830 & ~n1280;
  assign n49804 = n49802 & n49803;
  assign n49805 = n49801 & n49804;
  assign n49806 = n49800 & n49805;
  assign n49807 = ~n410 & n49802;
  assign n49808 = ~n559 & ~n1280;
  assign n49809 = ~n830 & ~n901;
  assign n49810 = n49801 & n49809;
  assign n49811 = n49808 & n49810;
  assign n49812 = n49807 & n49811;
  assign n49813 = n49783 & n59904;
  assign n49814 = ~n349 & ~n774;
  assign n49815 = ~n1033 & ~n1466;
  assign n49816 = n49814 & n49815;
  assign n49817 = ~n271 & ~n274;
  assign n49818 = n834 & n49817;
  assign n49819 = ~n271 & ~n774;
  assign n49820 = n49815 & n49819;
  assign n49821 = ~n274 & ~n349;
  assign n49822 = n834 & n49821;
  assign n49823 = n49820 & n49822;
  assign n49824 = ~n774 & ~n1033;
  assign n49825 = n834 & n49824;
  assign n49826 = ~n271 & ~n1466;
  assign n49827 = ~n349 & ~n1466;
  assign n49828 = n49817 & n49827;
  assign n49829 = n49821 & n49826;
  assign n49830 = n49825 & n59907;
  assign n49831 = n49816 & n49818;
  assign n49832 = n55108 & n56581;
  assign n49833 = n59906 & n49832;
  assign n49834 = n54471 & n49833;
  assign n49835 = n59905 & n49834;
  assign n49836 = n54456 & n49835;
  assign n49837 = n59903 & n49836;
  assign n49838 = n56581 & n56626;
  assign n49839 = n55108 & n49838;
  assign n49840 = n59903 & n49839;
  assign n49841 = n59905 & n49840;
  assign n49842 = n54471 & n49841;
  assign n49843 = n54456 & n49842;
  assign n49844 = ~n1033 & n49843;
  assign n49845 = ~n1466 & n49844;
  assign n49846 = ~n271 & n49845;
  assign n49847 = ~n833 & n49846;
  assign n49848 = ~n832 & n49847;
  assign n49849 = ~n274 & n49848;
  assign n49850 = ~n349 & n49849;
  assign n49851 = ~n774 & n49850;
  assign n49852 = n56626 & n49837;
  assign n49853 = ~n59870 & n59908;
  assign n49854 = n59870 & ~n59908;
  assign n49855 = ~n49853 & ~n49854;
  assign n49856 = ~n49530 & n49539;
  assign n49857 = ~n49530 & ~n49540;
  assign n49858 = ~n49531 & ~n49856;
  assign n49859 = ~n49854 & ~n59909;
  assign n49860 = ~n49853 & n49859;
  assign n49861 = n49855 & ~n59909;
  assign n49862 = ~n49855 & n59909;
  assign n49863 = ~n59909 & ~n59910;
  assign n49864 = ~n49854 & ~n59910;
  assign n49865 = ~n49853 & n49864;
  assign n49866 = ~n49863 & ~n49865;
  assign n49867 = ~n59910 & ~n49862;
  assign n49868 = n1576 & ~n58653;
  assign n49869 = n11215 & n39576;
  assign n49870 = n54403 & n39582;
  assign n49871 = n10564 & n39579;
  assign n49872 = ~n49870 & ~n49871;
  assign n49873 = ~n49869 & n49872;
  assign n49874 = ~n49868 & n49873;
  assign n49875 = ~n59911 & ~n49874;
  assign n49876 = n59911 & n49874;
  assign n49877 = ~n59911 & ~n49875;
  assign n49878 = ~n59911 & n49874;
  assign n49879 = ~n49874 & ~n49875;
  assign n49880 = n59911 & ~n49874;
  assign n49881 = ~n59912 & ~n59913;
  assign n49882 = ~n49875 & ~n49876;
  assign n49883 = n49737 & n59914;
  assign n49884 = ~n49737 & ~n59914;
  assign n49885 = ~n49883 & ~n49884;
  assign n49886 = n11279 & ~n58766;
  assign n49887 = n12584 & n39567;
  assign n49888 = n54410 & n39573;
  assign n49889 = n11267 & n39570;
  assign n49890 = ~n49888 & ~n49889;
  assign n49891 = ~n49887 & n49890;
  assign n49892 = ~n49886 & n49891;
  assign n49893 = pi29  & ~n49892;
  assign n49894 = pi29  & ~n49893;
  assign n49895 = pi29  & n49892;
  assign n49896 = ~n49892 & ~n49893;
  assign n49897 = ~pi29  & ~n49892;
  assign n49898 = ~n59915 & ~n59916;
  assign n49899 = n49885 & ~n49898;
  assign n49900 = ~n49885 & n49898;
  assign n49901 = n49885 & ~n49899;
  assign n49902 = n49885 & n49898;
  assign n49903 = ~n49898 & ~n49899;
  assign n49904 = ~n49885 & ~n49898;
  assign n49905 = ~n59917 & ~n59918;
  assign n49906 = ~n49899 & ~n49900;
  assign n49907 = ~n49736 & ~n59919;
  assign n49908 = n49736 & n59919;
  assign n49909 = ~n59919 & ~n49907;
  assign n49910 = n49736 & ~n59919;
  assign n49911 = ~n49736 & ~n49907;
  assign n49912 = ~n49736 & n59919;
  assign n49913 = ~n59920 & ~n59921;
  assign n49914 = ~n49907 & ~n49908;
  assign n49915 = ~n49568 & n49583;
  assign n49916 = ~n49568 & ~n49584;
  assign n49917 = ~n49569 & ~n49915;
  assign n49918 = n59922 & n59923;
  assign n49919 = ~n59922 & ~n59923;
  assign n49920 = ~n49918 & ~n49919;
  assign n49921 = n90 & ~n58889;
  assign n49922 = n14236 & n39549;
  assign n49923 = n54667 & n39555;
  assign n49924 = n14210 & n39552;
  assign n49925 = ~n49923 & ~n49924;
  assign n49926 = ~n49922 & n49925;
  assign n49927 = ~n49921 & n49926;
  assign n49928 = pi23  & ~n49927;
  assign n49929 = pi23  & ~n49928;
  assign n49930 = pi23  & n49927;
  assign n49931 = ~n49927 & ~n49928;
  assign n49932 = ~pi23  & ~n49927;
  assign n49933 = ~n59924 & ~n59925;
  assign n49934 = n49920 & ~n49933;
  assign n49935 = ~n49920 & n49933;
  assign n49936 = n49920 & ~n49934;
  assign n49937 = ~n49933 & ~n49934;
  assign n49938 = ~n49936 & ~n49937;
  assign n49939 = ~n49934 & ~n49935;
  assign n49940 = ~n49591 & n49605;
  assign n49941 = ~n49591 & ~n49607;
  assign n49942 = ~n49590 & ~n49940;
  assign n49943 = n59926 & n59927;
  assign n49944 = ~n59926 & ~n59927;
  assign n49945 = ~n49943 & ~n49944;
  assign n49946 = n14413 & ~n59044;
  assign n49947 = n15921 & n39543;
  assign n49948 = n54719 & n39546;
  assign n49949 = n15901 & n39440;
  assign n49950 = ~n49948 & ~n49949;
  assign n49951 = ~n49947 & n49950;
  assign n49952 = ~n49946 & n49951;
  assign n49953 = pi20  & ~n49952;
  assign n49954 = pi20  & ~n49953;
  assign n49955 = pi20  & n49952;
  assign n49956 = ~n49952 & ~n49953;
  assign n49957 = ~pi20  & ~n49952;
  assign n49958 = ~n59928 & ~n59929;
  assign n49959 = ~n49945 & n49958;
  assign n49960 = n49945 & ~n49958;
  assign n49961 = n49945 & ~n49960;
  assign n49962 = ~n49958 & ~n49960;
  assign n49963 = ~n49961 & ~n49962;
  assign n49964 = ~n49959 & ~n49960;
  assign n49965 = ~n49613 & n49627;
  assign n49966 = ~n49613 & ~n49628;
  assign n49967 = ~n49612 & ~n49965;
  assign n49968 = n59930 & n59931;
  assign n49969 = ~n59930 & ~n59931;
  assign n49970 = ~n49968 & ~n49969;
  assign n49971 = n16079 & ~n59282;
  assign n49972 = n16696 & n44775;
  assign n49973 = n54886 & n39937;
  assign n49974 = n16676 & n44327;
  assign n49975 = ~n49973 & ~n49974;
  assign n49976 = ~n49972 & n49975;
  assign n49977 = ~n49971 & n49976;
  assign n49978 = pi17  & ~n49977;
  assign n49979 = pi17  & ~n49978;
  assign n49980 = pi17  & n49977;
  assign n49981 = ~n49977 & ~n49978;
  assign n49982 = ~pi17  & ~n49977;
  assign n49983 = ~n59932 & ~n59933;
  assign n49984 = n49970 & ~n49983;
  assign n49985 = ~n49970 & n49983;
  assign n49986 = n49970 & ~n49984;
  assign n49987 = ~n49983 & ~n49984;
  assign n49988 = ~n49986 & ~n49987;
  assign n49989 = ~n49984 & ~n49985;
  assign n49990 = ~n49635 & n49649;
  assign n49991 = ~n49635 & ~n49651;
  assign n49992 = ~n49634 & ~n49990;
  assign n49993 = n59934 & n59935;
  assign n49994 = ~n59934 & ~n59935;
  assign n49995 = ~n49993 & ~n49994;
  assign n49996 = n17265 & ~n59386;
  assign n49997 = n18588 & n46009;
  assign n49998 = n55041 & n44871;
  assign n49999 = n18556 & n44952;
  assign n50000 = ~n49998 & ~n49999;
  assign n50001 = ~n49997 & n50000;
  assign n50002 = ~n49996 & n50001;
  assign n50003 = pi14  & ~n50002;
  assign n50004 = pi14  & ~n50003;
  assign n50005 = pi14  & n50002;
  assign n50006 = ~n50002 & ~n50003;
  assign n50007 = ~pi14  & ~n50002;
  assign n50008 = ~n59936 & ~n59937;
  assign n50009 = ~n49995 & n50008;
  assign n50010 = n49995 & ~n50008;
  assign n50011 = n49995 & ~n50010;
  assign n50012 = ~n50008 & ~n50010;
  assign n50013 = ~n50011 & ~n50012;
  assign n50014 = ~n50009 & ~n50010;
  assign n50015 = ~n49657 & n49671;
  assign n50016 = ~n49657 & ~n49672;
  assign n50017 = ~n49656 & ~n50015;
  assign n50018 = n59938 & n59939;
  assign n50019 = ~n59938 & ~n59939;
  assign n50020 = ~n50018 & ~n50019;
  assign n50021 = n18846 & ~n59554;
  assign n50022 = n19541 & n59503;
  assign n50023 = n55247 & n46420;
  assign n50024 = n19509 & n46788;
  assign n50025 = ~n50023 & ~n50024;
  assign n50026 = ~n50022 & n50025;
  assign n50027 = ~n50021 & n50026;
  assign n50028 = pi11  & ~n50027;
  assign n50029 = pi11  & ~n50028;
  assign n50030 = pi11  & n50027;
  assign n50031 = ~n50027 & ~n50028;
  assign n50032 = ~pi11  & ~n50027;
  assign n50033 = ~n59940 & ~n59941;
  assign n50034 = n50020 & ~n50033;
  assign n50035 = ~n50020 & n50033;
  assign n50036 = n50020 & ~n50034;
  assign n50037 = ~n50033 & ~n50034;
  assign n50038 = ~n50036 & ~n50037;
  assign n50039 = ~n50034 & ~n50035;
  assign n50040 = n49723 & ~n59942;
  assign n50041 = ~n49723 & n59942;
  assign n50042 = ~n59942 & ~n50040;
  assign n50043 = n49723 & ~n50040;
  assign n50044 = ~n50042 & ~n50043;
  assign n50045 = ~n50040 & ~n50041;
  assign n50046 = ~n49693 & n49701;
  assign n50047 = ~n49693 & ~n49702;
  assign n50048 = ~n49692 & ~n50046;
  assign n50049 = n59943 & n59944;
  assign n50050 = ~n59943 & ~n59944;
  assign n50051 = ~n50049 & ~n50050;
  assign n50052 = ~n49708 & ~n49715;
  assign n50053 = ~n50051 & n50052;
  assign n50054 = n50051 & ~n50052;
  assign n50055 = ~n50053 & ~n50054;
  assign n50056 = n49717 & n50055;
  assign n50057 = ~n49717 & ~n50055;
  assign po12  = ~n50056 & ~n50057;
  assign n50059 = ~n50050 & ~n50054;
  assign n50060 = ~n49899 & ~n49907;
  assign n50061 = ~n49875 & ~n49884;
  assign n50062 = n11279 & n41762;
  assign n50063 = n12584 & n39564;
  assign n50064 = n54410 & n39570;
  assign n50065 = n11267 & n39567;
  assign n50066 = ~n50064 & ~n50065;
  assign n50067 = ~n50063 & n50066;
  assign n50068 = ~n50062 & n50067;
  assign n50069 = pi29  & ~n50068;
  assign n50070 = pi29  & ~n50069;
  assign n50071 = pi29  & n50068;
  assign n50072 = ~n50068 & ~n50069;
  assign n50073 = ~pi29  & ~n50068;
  assign n50074 = ~n59945 & ~n59946;
  assign n50075 = n53809 & n54022;
  assign n50076 = n27165 & n50075;
  assign n50077 = n3001 & n3389;
  assign n50078 = n2004 & n50077;
  assign n50079 = ~n275 & ~n1997;
  assign n50080 = n494 & n50079;
  assign n50081 = n53761 & n50080;
  assign n50082 = n2004 & n3001;
  assign n50083 = n494 & n50082;
  assign n50084 = n3389 & n50079;
  assign n50085 = n53761 & n50084;
  assign n50086 = n50083 & n50085;
  assign n50087 = n50078 & n50081;
  assign n50088 = n56615 & n59947;
  assign n50089 = n53761 & n50075;
  assign n50090 = n494 & n27165;
  assign n50091 = n50082 & n50084;
  assign n50092 = n50090 & n50091;
  assign n50093 = n56615 & n50092;
  assign n50094 = n50089 & n50093;
  assign n50095 = n50076 & n50088;
  assign n50096 = n54157 & n59948;
  assign n50097 = n53782 & n54331;
  assign n50098 = n2004 & n53761;
  assign n50099 = n54022 & n50098;
  assign n50100 = n3001 & n50099;
  assign n50101 = n56615 & n50100;
  assign n50102 = n54157 & n50101;
  assign n50103 = n7144 & n50102;
  assign n50104 = n54331 & n50103;
  assign n50105 = n53809 & n50104;
  assign n50106 = n53782 & n50105;
  assign n50107 = n9477 & n50106;
  assign n50108 = n494 & n50107;
  assign n50109 = n3389 & n50108;
  assign n50110 = ~n1997 & n50109;
  assign n50111 = ~n275 & n50110;
  assign n50112 = n50096 & n50097;
  assign n50113 = n59870 & n59949;
  assign n50114 = ~n59870 & ~n59949;
  assign n50115 = ~n50113 & ~n50114;
  assign n50116 = ~pi8  & n50115;
  assign n50117 = pi8  & ~n50115;
  assign n50118 = ~n50116 & ~n50117;
  assign n50119 = ~n49864 & n50118;
  assign n50120 = n49864 & ~n50118;
  assign n50121 = ~n50119 & ~n50120;
  assign n50122 = n1576 & n39976;
  assign n50123 = n11215 & n39573;
  assign n50124 = n54403 & n39579;
  assign n50125 = n10564 & n39576;
  assign n50126 = ~n50124 & ~n50125;
  assign n50127 = ~n50123 & n50126;
  assign n50128 = ~n50122 & n50127;
  assign n50129 = n50121 & ~n50128;
  assign n50130 = ~n50121 & n50128;
  assign n50131 = n50121 & ~n50129;
  assign n50132 = ~n50128 & ~n50129;
  assign n50133 = ~n50131 & ~n50132;
  assign n50134 = ~n50129 & ~n50130;
  assign n50135 = ~n50074 & ~n59950;
  assign n50136 = n50074 & n59950;
  assign n50137 = ~n59950 & ~n50135;
  assign n50138 = ~n50074 & ~n50135;
  assign n50139 = ~n50137 & ~n50138;
  assign n50140 = ~n50135 & ~n50136;
  assign n50141 = n50061 & n59951;
  assign n50142 = ~n50061 & ~n59951;
  assign n50143 = ~n50141 & ~n50142;
  assign n50144 = n123 & n42574;
  assign n50145 = n128 & n39555;
  assign n50146 = n53444 & n39561;
  assign n50147 = n127 & n39558;
  assign n50148 = ~n50146 & ~n50147;
  assign n50149 = ~n50145 & n50148;
  assign n50150 = ~n50144 & n50149;
  assign n50151 = pi26  & ~n50150;
  assign n50152 = pi26  & ~n50151;
  assign n50153 = pi26  & n50150;
  assign n50154 = ~n50150 & ~n50151;
  assign n50155 = ~pi26  & ~n50150;
  assign n50156 = ~n59952 & ~n59953;
  assign n50157 = n50143 & ~n50156;
  assign n50158 = ~n50143 & n50156;
  assign n50159 = n50143 & ~n50157;
  assign n50160 = n50143 & n50156;
  assign n50161 = ~n50156 & ~n50157;
  assign n50162 = ~n50143 & ~n50156;
  assign n50163 = ~n59954 & ~n59955;
  assign n50164 = ~n50157 & ~n50158;
  assign n50165 = n50060 & n59956;
  assign n50166 = ~n50060 & ~n59956;
  assign n50167 = ~n50165 & ~n50166;
  assign n50168 = n90 & n43436;
  assign n50169 = n14236 & n39546;
  assign n50170 = n54667 & n39552;
  assign n50171 = n14210 & n39549;
  assign n50172 = ~n50170 & ~n50171;
  assign n50173 = ~n50169 & n50172;
  assign n50174 = ~n50168 & n50173;
  assign n50175 = pi23  & ~n50174;
  assign n50176 = pi23  & ~n50175;
  assign n50177 = pi23  & n50174;
  assign n50178 = ~n50174 & ~n50175;
  assign n50179 = ~pi23  & ~n50174;
  assign n50180 = ~n59957 & ~n59958;
  assign n50181 = n50167 & ~n50180;
  assign n50182 = ~n50167 & n50180;
  assign n50183 = n50167 & ~n50181;
  assign n50184 = n50167 & n50180;
  assign n50185 = ~n50180 & ~n50181;
  assign n50186 = ~n50167 & ~n50180;
  assign n50187 = ~n59959 & ~n59960;
  assign n50188 = ~n50181 & ~n50182;
  assign n50189 = ~n49919 & n49933;
  assign n50190 = ~n49919 & ~n49934;
  assign n50191 = ~n49918 & ~n50189;
  assign n50192 = n59961 & n59962;
  assign n50193 = ~n59961 & ~n59962;
  assign n50194 = ~n50192 & ~n50193;
  assign n50195 = n14413 & n39943;
  assign n50196 = n15921 & n39937;
  assign n50197 = n54719 & n39440;
  assign n50198 = n15901 & n39543;
  assign n50199 = ~n50197 & ~n50198;
  assign n50200 = ~n50196 & n50199;
  assign n50201 = ~n50195 & n50200;
  assign n50202 = pi20  & ~n50201;
  assign n50203 = pi20  & ~n50202;
  assign n50204 = pi20  & n50201;
  assign n50205 = ~n50201 & ~n50202;
  assign n50206 = ~pi20  & ~n50201;
  assign n50207 = ~n59963 & ~n59964;
  assign n50208 = n50194 & ~n50207;
  assign n50209 = ~n50194 & n50207;
  assign n50210 = n50194 & ~n50208;
  assign n50211 = n50194 & n50207;
  assign n50212 = ~n50207 & ~n50208;
  assign n50213 = ~n50194 & ~n50207;
  assign n50214 = ~n59965 & ~n59966;
  assign n50215 = ~n50208 & ~n50209;
  assign n50216 = ~n49944 & n49958;
  assign n50217 = ~n49944 & ~n49960;
  assign n50218 = ~n49943 & ~n50216;
  assign n50219 = n59967 & n59968;
  assign n50220 = ~n59967 & ~n59968;
  assign n50221 = ~n50219 & ~n50220;
  assign n50222 = n16079 & ~n59280;
  assign n50223 = n16696 & n44871;
  assign n50224 = n54886 & n44327;
  assign n50225 = n16676 & n44775;
  assign n50226 = ~n50224 & ~n50225;
  assign n50227 = ~n50223 & n50226;
  assign n50228 = ~n50222 & n50227;
  assign n50229 = pi17  & ~n50228;
  assign n50230 = pi17  & ~n50229;
  assign n50231 = pi17  & n50228;
  assign n50232 = ~n50228 & ~n50229;
  assign n50233 = ~pi17  & ~n50228;
  assign n50234 = ~n59969 & ~n59970;
  assign n50235 = ~n49969 & n49983;
  assign n50236 = ~n49969 & ~n49984;
  assign n50237 = ~n49968 & ~n50235;
  assign n50238 = ~n50234 & ~n59971;
  assign n50239 = n50234 & n59971;
  assign n50240 = ~n59971 & ~n50238;
  assign n50241 = n50234 & ~n59971;
  assign n50242 = ~n50234 & ~n50238;
  assign n50243 = ~n50234 & n59971;
  assign n50244 = ~n59972 & ~n59973;
  assign n50245 = ~n50238 & ~n50239;
  assign n50246 = ~n50221 & n59974;
  assign n50247 = n50221 & ~n59974;
  assign n50248 = ~n50246 & ~n50247;
  assign n50249 = n17265 & n46426;
  assign n50250 = n18588 & n46420;
  assign n50251 = n55041 & n44952;
  assign n50252 = n18556 & n46009;
  assign n50253 = ~n50251 & ~n50252;
  assign n50254 = ~n50250 & n50253;
  assign n50255 = ~n50249 & n50254;
  assign n50256 = pi14  & ~n50255;
  assign n50257 = pi14  & ~n50256;
  assign n50258 = pi14  & n50255;
  assign n50259 = ~n50255 & ~n50256;
  assign n50260 = ~pi14  & ~n50255;
  assign n50261 = ~n59975 & ~n59976;
  assign n50262 = n50248 & ~n50261;
  assign n50263 = ~n50248 & n50261;
  assign n50264 = n50248 & ~n50262;
  assign n50265 = n50248 & n50261;
  assign n50266 = ~n50261 & ~n50262;
  assign n50267 = ~n50248 & ~n50261;
  assign n50268 = ~n59977 & ~n59978;
  assign n50269 = ~n50262 & ~n50263;
  assign n50270 = ~n49994 & n50008;
  assign n50271 = ~n49994 & ~n50010;
  assign n50272 = ~n49993 & ~n50270;
  assign n50273 = n59979 & n59980;
  assign n50274 = ~n59979 & ~n59980;
  assign n50275 = ~n50273 & ~n50274;
  assign n50276 = n18846 & ~n47526;
  assign n50277 = n55247 & n46788;
  assign n50278 = n19509 & n59503;
  assign n50279 = ~n50277 & ~n50278;
  assign n50280 = ~n50276 & n50279;
  assign n50281 = pi11  & ~n50280;
  assign n50282 = pi11  & ~n50281;
  assign n50283 = pi11  & n50280;
  assign n50284 = ~n50280 & ~n50281;
  assign n50285 = ~pi11  & ~n50280;
  assign n50286 = ~n59981 & ~n59982;
  assign n50287 = ~n50019 & n50033;
  assign n50288 = ~n50019 & ~n50034;
  assign n50289 = ~n50018 & ~n50287;
  assign n50290 = ~n50286 & ~n59983;
  assign n50291 = n50286 & n59983;
  assign n50292 = ~n59983 & ~n50290;
  assign n50293 = n50286 & ~n59983;
  assign n50294 = ~n50286 & ~n50290;
  assign n50295 = ~n50286 & n59983;
  assign n50296 = ~n59984 & ~n59985;
  assign n50297 = ~n50290 & ~n50291;
  assign n50298 = ~n50275 & n59986;
  assign n50299 = n50275 & ~n59986;
  assign n50300 = ~n50298 & ~n50299;
  assign n50301 = ~n49721 & n59942;
  assign n50302 = ~n49721 & ~n50040;
  assign n50303 = ~n49722 & ~n50301;
  assign n50304 = n50300 & ~n59987;
  assign n50305 = ~n50300 & n59987;
  assign n50306 = ~n50304 & ~n50305;
  assign n50307 = ~n50059 & n50306;
  assign n50308 = n50059 & ~n50306;
  assign n50309 = ~n50307 & ~n50308;
  assign n50310 = ~n50056 & ~n50309;
  assign n50311 = n50056 & n50309;
  assign po13  = ~n50310 & ~n50311;
  assign n50313 = ~n50304 & ~n50307;
  assign n50314 = ~n50290 & ~n50299;
  assign n50315 = ~n50262 & ~n50274;
  assign n50316 = n17265 & n46805;
  assign n50317 = n18588 & n46788;
  assign n50318 = n55041 & n46009;
  assign n50319 = n18556 & n46420;
  assign n50320 = ~n50318 & ~n50319;
  assign n50321 = ~n50317 & n50320;
  assign n50322 = ~n50316 & n50321;
  assign n50323 = pi14  & ~n50322;
  assign n50324 = pi14  & ~n50323;
  assign n50325 = pi14  & n50322;
  assign n50326 = ~n50322 & ~n50323;
  assign n50327 = ~pi14  & ~n50322;
  assign n50328 = ~n59988 & ~n59989;
  assign n50329 = ~n50238 & ~n50247;
  assign n50330 = ~n50208 & ~n50220;
  assign n50331 = ~n50181 & ~n50193;
  assign n50332 = ~n50157 & ~n50166;
  assign n50333 = ~n50135 & ~n50142;
  assign n50334 = ~n50114 & ~n50116;
  assign n50335 = ~n450 & ~n493;
  assign n50336 = ~n450 & ~n1881;
  assign n50337 = ~n493 & n50336;
  assign n50338 = ~n1881 & n50335;
  assign n50339 = n53585 & n59990;
  assign n50340 = n53518 & n57026;
  assign n50341 = n50339 & n50340;
  assign n50342 = n3000 & n9861;
  assign n50343 = n10901 & n29675;
  assign n50344 = n3000 & n10901;
  assign n50345 = n9861 & n29675;
  assign n50346 = n50344 & n50345;
  assign n50347 = n50342 & n50343;
  assign n50348 = n54729 & n59991;
  assign n50349 = ~n660 & n29675;
  assign n50350 = n53585 & n50349;
  assign n50351 = n50340 & n50350;
  assign n50352 = ~n414 & ~n450;
  assign n50353 = ~n493 & ~n1881;
  assign n50354 = n50352 & n50353;
  assign n50355 = n50344 & n50354;
  assign n50356 = n54729 & n50355;
  assign n50357 = n50351 & n50356;
  assign n50358 = n50341 & n50348;
  assign n50359 = n56715 & n59992;
  assign n50360 = n53740 & n50359;
  assign n50361 = n53585 & n3000;
  assign n50362 = n57026 & n50361;
  assign n50363 = n56715 & n50362;
  assign n50364 = n54729 & n50363;
  assign n50365 = n10901 & n50364;
  assign n50366 = n54084 & n50365;
  assign n50367 = n53740 & n50366;
  assign n50368 = n53518 & n50367;
  assign n50369 = ~n414 & n50368;
  assign n50370 = ~n1492 & n50369;
  assign n50371 = ~n660 & n50370;
  assign n50372 = ~n956 & n50371;
  assign n50373 = ~n493 & n50372;
  assign n50374 = ~n450 & n50373;
  assign n50375 = ~n1881 & n50374;
  assign n50376 = n54084 & n50360;
  assign n50377 = ~n50334 & n59993;
  assign n50378 = n50334 & ~n59993;
  assign n50379 = ~n50377 & ~n50378;
  assign n50380 = n1576 & ~n58759;
  assign n50381 = n11215 & n39570;
  assign n50382 = n54403 & n39576;
  assign n50383 = n10564 & n39573;
  assign n50384 = ~n50382 & ~n50383;
  assign n50385 = ~n50381 & n50384;
  assign n50386 = ~n50380 & n50385;
  assign n50387 = n50379 & ~n50386;
  assign n50388 = ~n50379 & n50386;
  assign n50389 = ~n50386 & ~n50387;
  assign n50390 = n50379 & ~n50387;
  assign n50391 = ~n50389 & ~n50390;
  assign n50392 = ~n50387 & ~n50388;
  assign n50393 = ~n50119 & n50128;
  assign n50394 = ~n50119 & ~n50129;
  assign n50395 = ~n50120 & ~n50393;
  assign n50396 = n59994 & n59995;
  assign n50397 = ~n59994 & ~n59995;
  assign n50398 = ~n50396 & ~n50397;
  assign n50399 = n11279 & ~n58493;
  assign n50400 = n12584 & n39561;
  assign n50401 = n54410 & n39567;
  assign n50402 = n11267 & n39564;
  assign n50403 = ~n50401 & ~n50402;
  assign n50404 = ~n50400 & n50403;
  assign n50405 = ~n11279 & n50404;
  assign n50406 = n58493 & n50404;
  assign n50407 = ~n50405 & ~n50406;
  assign n50408 = ~n50399 & n50404;
  assign n50409 = pi29  & ~n59996;
  assign n50410 = ~pi29  & n59996;
  assign n50411 = ~n50409 & ~n50410;
  assign n50412 = n50398 & ~n50411;
  assign n50413 = ~n50398 & n50411;
  assign n50414 = ~n50412 & ~n50413;
  assign n50415 = ~n50333 & n50414;
  assign n50416 = n50333 & ~n50414;
  assign n50417 = ~n50415 & ~n50416;
  assign n50418 = n123 & ~n58891;
  assign n50419 = n128 & n39552;
  assign n50420 = n53444 & n39558;
  assign n50421 = n127 & n39555;
  assign n50422 = ~n50420 & ~n50421;
  assign n50423 = ~n50419 & n50422;
  assign n50424 = ~n50418 & n50423;
  assign n50425 = pi26  & ~n50424;
  assign n50426 = pi26  & ~n50425;
  assign n50427 = pi26  & n50424;
  assign n50428 = ~n50424 & ~n50425;
  assign n50429 = ~pi26  & ~n50424;
  assign n50430 = ~n59997 & ~n59998;
  assign n50431 = n50417 & ~n50430;
  assign n50432 = ~n50417 & n50430;
  assign n50433 = n50417 & ~n50431;
  assign n50434 = ~n50430 & ~n50431;
  assign n50435 = ~n50433 & ~n50434;
  assign n50436 = ~n50431 & ~n50432;
  assign n50437 = n50332 & n59999;
  assign n50438 = ~n50332 & ~n59999;
  assign n50439 = ~n50437 & ~n50438;
  assign n50440 = n90 & ~n59050;
  assign n50441 = n14236 & n39440;
  assign n50442 = n54667 & n39549;
  assign n50443 = n14210 & n39546;
  assign n50444 = ~n50442 & ~n50443;
  assign n50445 = ~n50441 & n50444;
  assign n50446 = ~n50440 & n50445;
  assign n50447 = pi23  & ~n50446;
  assign n50448 = pi23  & ~n50447;
  assign n50449 = pi23  & n50446;
  assign n50450 = ~n50446 & ~n50447;
  assign n50451 = ~pi23  & ~n50446;
  assign n50452 = ~n60000 & ~n60001;
  assign n50453 = ~n50439 & n50452;
  assign n50454 = n50439 & ~n50452;
  assign n50455 = n50439 & ~n50454;
  assign n50456 = ~n50452 & ~n50454;
  assign n50457 = ~n50455 & ~n50456;
  assign n50458 = ~n50453 & ~n50454;
  assign n50459 = n50331 & n60002;
  assign n50460 = ~n50331 & ~n60002;
  assign n50461 = ~n50459 & ~n50460;
  assign n50462 = n14413 & ~n59184;
  assign n50463 = n15921 & n44327;
  assign n50464 = n54719 & n39543;
  assign n50465 = n15901 & n39937;
  assign n50466 = ~n50464 & ~n50465;
  assign n50467 = ~n50463 & n50466;
  assign n50468 = ~n50462 & n50467;
  assign n50469 = pi20  & ~n50468;
  assign n50470 = pi20  & ~n50469;
  assign n50471 = pi20  & n50468;
  assign n50472 = ~n50468 & ~n50469;
  assign n50473 = ~pi20  & ~n50468;
  assign n50474 = ~n60003 & ~n60004;
  assign n50475 = n50461 & ~n50474;
  assign n50476 = ~n50461 & n50474;
  assign n50477 = n50461 & ~n50475;
  assign n50478 = ~n50474 & ~n50475;
  assign n50479 = ~n50477 & ~n50478;
  assign n50480 = ~n50475 & ~n50476;
  assign n50481 = n50330 & n60005;
  assign n50482 = ~n50330 & ~n60005;
  assign n50483 = ~n50481 & ~n50482;
  assign n50484 = n16079 & ~n59275;
  assign n50485 = n16696 & n44952;
  assign n50486 = n54886 & n44775;
  assign n50487 = n16676 & n44871;
  assign n50488 = ~n50486 & ~n50487;
  assign n50489 = ~n50485 & n50488;
  assign n50490 = ~n50484 & n50489;
  assign n50491 = pi17  & ~n50490;
  assign n50492 = pi17  & ~n50491;
  assign n50493 = pi17  & n50490;
  assign n50494 = ~n50490 & ~n50491;
  assign n50495 = ~pi17  & ~n50490;
  assign n50496 = ~n60006 & ~n60007;
  assign n50497 = ~n50483 & n50496;
  assign n50498 = n50483 & ~n50496;
  assign n50499 = n50483 & ~n50498;
  assign n50500 = ~n50496 & ~n50498;
  assign n50501 = ~n50499 & ~n50500;
  assign n50502 = ~n50497 & ~n50498;
  assign n50503 = ~n50329 & ~n60008;
  assign n50504 = n50329 & n60008;
  assign n50505 = ~n60008 & ~n50503;
  assign n50506 = n50329 & ~n60008;
  assign n50507 = ~n50329 & ~n50503;
  assign n50508 = ~n50329 & n60008;
  assign n50509 = ~n60009 & ~n60010;
  assign n50510 = ~n50503 & ~n50504;
  assign n50511 = ~n50328 & ~n60011;
  assign n50512 = n50328 & n60011;
  assign n50513 = ~n60011 & ~n50511;
  assign n50514 = ~n50328 & ~n50511;
  assign n50515 = ~n50513 & ~n50514;
  assign n50516 = ~n50511 & ~n50512;
  assign n50517 = n50315 & n60012;
  assign n50518 = ~n50315 & ~n60012;
  assign n50519 = ~n50517 & ~n50518;
  assign n50520 = n55247 & n59503;
  assign n50521 = pi11  & n50520;
  assign n50522 = pi11  & ~n50521;
  assign n50523 = pi11  & ~n50520;
  assign n50524 = n50520 & ~n50521;
  assign n50525 = ~pi11  & n50520;
  assign n50526 = ~n60013 & ~n60014;
  assign n50527 = n50519 & ~n50526;
  assign n50528 = ~n50519 & n50526;
  assign n50529 = n50519 & ~n50527;
  assign n50530 = ~n50526 & ~n50527;
  assign n50531 = ~n50529 & ~n50530;
  assign n50532 = ~n50527 & ~n50528;
  assign n50533 = ~n50314 & ~n60015;
  assign n50534 = n50314 & n60015;
  assign n50535 = ~n60015 & ~n50533;
  assign n50536 = ~n50314 & ~n50533;
  assign n50537 = ~n50535 & ~n50536;
  assign n50538 = ~n50533 & ~n50534;
  assign n50539 = n50313 & n60016;
  assign n50540 = ~n50313 & ~n60016;
  assign n50541 = ~n50539 & ~n50540;
  assign n50542 = n50311 & n50541;
  assign n50543 = ~n50311 & ~n50541;
  assign po14  = ~n50542 & ~n50543;
  assign n50545 = ~n50503 & ~n50511;
  assign n50546 = pi11  & ~n50545;
  assign n50547 = ~pi11  & n50545;
  assign n50548 = ~n50546 & ~n50547;
  assign n50549 = ~n50397 & ~n50412;
  assign n50550 = n11279 & ~n58849;
  assign n50551 = n12584 & n39558;
  assign n50552 = n54410 & n39564;
  assign n50553 = n11267 & n39561;
  assign n50554 = ~n50552 & ~n50553;
  assign n50555 = ~n50551 & n50554;
  assign n50556 = ~n11279 & n50555;
  assign n50557 = n58849 & n50555;
  assign n50558 = ~n50556 & ~n50557;
  assign n50559 = ~n50550 & n50555;
  assign n50560 = pi29  & ~n60017;
  assign n50561 = ~pi29  & n60017;
  assign n50562 = ~n50560 & ~n50561;
  assign n50563 = ~n466 & ~n564;
  assign n50564 = ~n564 & ~n1641;
  assign n50565 = ~n466 & n50564;
  assign n50566 = ~n1641 & n50563;
  assign n50567 = n3528 & n60018;
  assign n50568 = n54321 & n50567;
  assign n50569 = n3214 & n5538;
  assign n50570 = n2094 & n10300;
  assign n50571 = n50569 & n50570;
  assign n50572 = n3780 & n4795;
  assign n50573 = n5021 & n5362;
  assign n50574 = n50572 & n50573;
  assign n50575 = n50571 & n50574;
  assign n50576 = n3214 & n3780;
  assign n50577 = n60018 & n50576;
  assign n50578 = n54321 & n50577;
  assign n50579 = n5362 & n5538;
  assign n50580 = n50570 & n50579;
  assign n50581 = n4795 & n5021;
  assign n50582 = n3528 & n50581;
  assign n50583 = n50580 & n50582;
  assign n50584 = n50578 & n50583;
  assign n50585 = n1673 & n4795;
  assign n50586 = n60018 & n50585;
  assign n50587 = n54321 & n50586;
  assign n50588 = n3214 & n3463;
  assign n50589 = n3780 & n10300;
  assign n50590 = n50588 & n50589;
  assign n50591 = n2094 & n5538;
  assign n50592 = n50573 & n50591;
  assign n50593 = n50590 & n50592;
  assign n50594 = n50587 & n50593;
  assign n50595 = n50568 & n50575;
  assign n50596 = n56622 & n56910;
  assign n50597 = n60019 & n50596;
  assign n50598 = n54827 & n50597;
  assign n50599 = n54321 & n10300;
  assign n50600 = n3463 & n50599;
  assign n50601 = n5538 & n50600;
  assign n50602 = n5362 & n50601;
  assign n50603 = n56622 & n50602;
  assign n50604 = n56910 & n50603;
  assign n50605 = n54827 & n50604;
  assign n50606 = n3780 & n50605;
  assign n50607 = n1673 & n50606;
  assign n50608 = n3214 & n50607;
  assign n50609 = n59867 & n50608;
  assign n50610 = n5021 & n50609;
  assign n50611 = n2094 & n50610;
  assign n50612 = ~n1469 & n50611;
  assign n50613 = ~n272 & n50612;
  assign n50614 = ~n564 & n50613;
  assign n50615 = ~n1641 & n50614;
  assign n50616 = ~n466 & n50615;
  assign n50617 = n59867 & n50598;
  assign n50618 = ~n59993 & n60020;
  assign n50619 = n59993 & ~n60020;
  assign n50620 = ~n50618 & ~n50619;
  assign n50621 = ~n50377 & n50386;
  assign n50622 = ~n50377 & ~n50387;
  assign n50623 = ~n50378 & ~n50621;
  assign n50624 = ~n50619 & ~n60021;
  assign n50625 = ~n50618 & n50624;
  assign n50626 = n50620 & ~n60021;
  assign n50627 = ~n50620 & n60021;
  assign n50628 = ~n60021 & ~n60022;
  assign n50629 = ~n50619 & ~n60022;
  assign n50630 = ~n50618 & n50629;
  assign n50631 = ~n50628 & ~n50630;
  assign n50632 = ~n60022 & ~n50627;
  assign n50633 = n1576 & ~n58766;
  assign n50634 = n11215 & n39567;
  assign n50635 = n54403 & n39573;
  assign n50636 = n10564 & n39570;
  assign n50637 = ~n50635 & ~n50636;
  assign n50638 = ~n50634 & n50637;
  assign n50639 = ~n50633 & n50638;
  assign n50640 = ~n60023 & ~n50639;
  assign n50641 = n60023 & n50639;
  assign n50642 = ~n60023 & ~n50640;
  assign n50643 = ~n60023 & n50639;
  assign n50644 = ~n50639 & ~n50640;
  assign n50645 = n60023 & ~n50639;
  assign n50646 = ~n60024 & ~n60025;
  assign n50647 = ~n50640 & ~n50641;
  assign n50648 = ~n50562 & ~n60026;
  assign n50649 = n50562 & n60026;
  assign n50650 = ~n50648 & ~n50649;
  assign n50651 = ~n50549 & n50650;
  assign n50652 = n50549 & ~n50650;
  assign n50653 = ~n50651 & ~n50652;
  assign n50654 = n123 & ~n58889;
  assign n50655 = n128 & n39549;
  assign n50656 = n53444 & n39555;
  assign n50657 = n127 & n39552;
  assign n50658 = ~n50656 & ~n50657;
  assign n50659 = ~n50655 & n50658;
  assign n50660 = ~n50654 & n50659;
  assign n50661 = pi26  & ~n50660;
  assign n50662 = pi26  & ~n50661;
  assign n50663 = pi26  & n50660;
  assign n50664 = ~n50660 & ~n50661;
  assign n50665 = ~pi26  & ~n50660;
  assign n50666 = ~n60027 & ~n60028;
  assign n50667 = n50653 & ~n50666;
  assign n50668 = ~n50653 & n50666;
  assign n50669 = n50653 & ~n50667;
  assign n50670 = ~n50666 & ~n50667;
  assign n50671 = ~n50669 & ~n50670;
  assign n50672 = ~n50667 & ~n50668;
  assign n50673 = ~n50415 & n50430;
  assign n50674 = ~n50415 & ~n50431;
  assign n50675 = ~n50416 & ~n50673;
  assign n50676 = n60029 & n60030;
  assign n50677 = ~n60029 & ~n60030;
  assign n50678 = ~n50676 & ~n50677;
  assign n50679 = n90 & ~n59044;
  assign n50680 = n14236 & n39543;
  assign n50681 = n54667 & n39546;
  assign n50682 = n14210 & n39440;
  assign n50683 = ~n50681 & ~n50682;
  assign n50684 = ~n50680 & n50683;
  assign n50685 = ~n50679 & n50684;
  assign n50686 = pi23  & ~n50685;
  assign n50687 = pi23  & ~n50686;
  assign n50688 = pi23  & n50685;
  assign n50689 = ~n50685 & ~n50686;
  assign n50690 = ~pi23  & ~n50685;
  assign n50691 = ~n60031 & ~n60032;
  assign n50692 = ~n50678 & n50691;
  assign n50693 = n50678 & ~n50691;
  assign n50694 = n50678 & ~n50693;
  assign n50695 = ~n50691 & ~n50693;
  assign n50696 = ~n50694 & ~n50695;
  assign n50697 = ~n50692 & ~n50693;
  assign n50698 = ~n50438 & n50452;
  assign n50699 = ~n50438 & ~n50454;
  assign n50700 = ~n50437 & ~n50698;
  assign n50701 = n60033 & n60034;
  assign n50702 = ~n60033 & ~n60034;
  assign n50703 = ~n50701 & ~n50702;
  assign n50704 = n14413 & ~n59282;
  assign n50705 = n15921 & n44775;
  assign n50706 = n54719 & n39937;
  assign n50707 = n15901 & n44327;
  assign n50708 = ~n50706 & ~n50707;
  assign n50709 = ~n50705 & n50708;
  assign n50710 = ~n50704 & n50709;
  assign n50711 = pi20  & ~n50710;
  assign n50712 = pi20  & ~n50711;
  assign n50713 = pi20  & n50710;
  assign n50714 = ~n50710 & ~n50711;
  assign n50715 = ~pi20  & ~n50710;
  assign n50716 = ~n60035 & ~n60036;
  assign n50717 = n50703 & ~n50716;
  assign n50718 = ~n50703 & n50716;
  assign n50719 = n50703 & ~n50717;
  assign n50720 = ~n50716 & ~n50717;
  assign n50721 = ~n50719 & ~n50720;
  assign n50722 = ~n50717 & ~n50718;
  assign n50723 = ~n50460 & n50474;
  assign n50724 = ~n50460 & ~n50475;
  assign n50725 = ~n50459 & ~n50723;
  assign n50726 = n60037 & n60038;
  assign n50727 = ~n60037 & ~n60038;
  assign n50728 = ~n50726 & ~n50727;
  assign n50729 = n16079 & ~n59386;
  assign n50730 = n16696 & n46009;
  assign n50731 = n54886 & n44871;
  assign n50732 = n16676 & n44952;
  assign n50733 = ~n50731 & ~n50732;
  assign n50734 = ~n50730 & n50733;
  assign n50735 = ~n50729 & n50734;
  assign n50736 = pi17  & ~n50735;
  assign n50737 = pi17  & ~n50736;
  assign n50738 = pi17  & n50735;
  assign n50739 = ~n50735 & ~n50736;
  assign n50740 = ~pi17  & ~n50735;
  assign n50741 = ~n60039 & ~n60040;
  assign n50742 = ~n50728 & n50741;
  assign n50743 = n50728 & ~n50741;
  assign n50744 = n50728 & ~n50743;
  assign n50745 = ~n50741 & ~n50743;
  assign n50746 = ~n50744 & ~n50745;
  assign n50747 = ~n50742 & ~n50743;
  assign n50748 = ~n50482 & n50496;
  assign n50749 = ~n50482 & ~n50498;
  assign n50750 = ~n50481 & ~n50748;
  assign n50751 = n60041 & n60042;
  assign n50752 = ~n60041 & ~n60042;
  assign n50753 = ~n50751 & ~n50752;
  assign n50754 = n17265 & ~n59554;
  assign n50755 = n18588 & n59503;
  assign n50756 = n55041 & n46420;
  assign n50757 = n18556 & n46788;
  assign n50758 = ~n50756 & ~n50757;
  assign n50759 = ~n50755 & n50758;
  assign n50760 = ~n50754 & n50759;
  assign n50761 = pi14  & ~n50760;
  assign n50762 = pi14  & ~n50761;
  assign n50763 = pi14  & n50760;
  assign n50764 = ~n50760 & ~n50761;
  assign n50765 = ~pi14  & ~n50760;
  assign n50766 = ~n60043 & ~n60044;
  assign n50767 = n50753 & ~n50766;
  assign n50768 = ~n50753 & n50766;
  assign n50769 = n50753 & ~n50767;
  assign n50770 = ~n50766 & ~n50767;
  assign n50771 = ~n50769 & ~n50770;
  assign n50772 = ~n50767 & ~n50768;
  assign n50773 = n50548 & ~n60045;
  assign n50774 = ~n50548 & n60045;
  assign n50775 = ~n60045 & ~n50773;
  assign n50776 = n50548 & ~n50773;
  assign n50777 = ~n50775 & ~n50776;
  assign n50778 = ~n50773 & ~n50774;
  assign n50779 = ~n50518 & n50526;
  assign n50780 = ~n50518 & ~n50527;
  assign n50781 = ~n50517 & ~n50779;
  assign n50782 = n60046 & n60047;
  assign n50783 = ~n60046 & ~n60047;
  assign n50784 = ~n50782 & ~n50783;
  assign n50785 = ~n50533 & ~n50540;
  assign n50786 = ~n50784 & n50785;
  assign n50787 = n50784 & ~n50785;
  assign n50788 = ~n50786 & ~n50787;
  assign n50789 = n50542 & n50788;
  assign n50790 = ~n50542 & ~n50788;
  assign po15  = ~n50789 & ~n50790;
  assign n50792 = ~n50783 & ~n50787;
  assign n50793 = n123 & n43436;
  assign n50794 = n128 & n39546;
  assign n50795 = n53444 & n39552;
  assign n50796 = n127 & n39549;
  assign n50797 = ~n50795 & ~n50796;
  assign n50798 = ~n50794 & n50797;
  assign n50799 = ~n50793 & n50798;
  assign n50800 = pi26  & ~n50799;
  assign n50801 = pi26  & ~n50800;
  assign n50802 = pi26  & n50799;
  assign n50803 = ~n50799 & ~n50800;
  assign n50804 = ~pi26  & ~n50799;
  assign n50805 = ~n60048 & ~n60049;
  assign n50806 = n11279 & n42574;
  assign n50807 = n12584 & n39555;
  assign n50808 = n54410 & n39561;
  assign n50809 = n11267 & n39558;
  assign n50810 = ~n50808 & ~n50809;
  assign n50811 = ~n50807 & n50810;
  assign n50812 = ~n50806 & n50811;
  assign n50813 = pi29  & ~n50812;
  assign n50814 = pi29  & ~n50813;
  assign n50815 = pi29  & n50812;
  assign n50816 = ~n50812 & ~n50813;
  assign n50817 = ~pi29  & ~n50812;
  assign n50818 = ~n60050 & ~n60051;
  assign n50819 = ~n50640 & ~n50648;
  assign n50820 = ~n271 & ~n622;
  assign n50821 = ~n414 & ~n447;
  assign n50822 = ~n414 & ~n622;
  assign n50823 = ~n271 & ~n447;
  assign n50824 = n50822 & n50823;
  assign n50825 = ~n447 & ~n622;
  assign n50826 = ~n271 & ~n414;
  assign n50827 = n50825 & n50826;
  assign n50828 = n50820 & n50821;
  assign n50829 = n1278 & n2367;
  assign n50830 = n60052 & n50829;
  assign n50831 = n54773 & n39276;
  assign n50832 = n50830 & n50831;
  assign n50833 = n1060 & n3670;
  assign n50834 = n10184 & n50833;
  assign n50835 = n54188 & n50834;
  assign n50836 = n54776 & n50835;
  assign n50837 = n1060 & n2367;
  assign n50838 = n39276 & n50837;
  assign n50839 = n54773 & n60052;
  assign n50840 = n50838 & n50839;
  assign n50841 = n3670 & n10184;
  assign n50842 = n1278 & n50841;
  assign n50843 = n54188 & n50842;
  assign n50844 = n54776 & n50843;
  assign n50845 = n50840 & n50844;
  assign n50846 = n50832 & n50836;
  assign n50847 = n54009 & n60053;
  assign n50848 = n53749 & n54019;
  assign n50849 = n1060 & n54188;
  assign n50850 = n54773 & n50849;
  assign n50851 = n10184 & n50850;
  assign n50852 = n54776 & n50851;
  assign n50853 = n54019 & n50852;
  assign n50854 = n53749 & n50853;
  assign n50855 = n4313 & n50854;
  assign n50856 = n54009 & n50855;
  assign n50857 = n3670 & n50856;
  assign n50858 = n905 & n50857;
  assign n50859 = n1278 & n50858;
  assign n50860 = n2367 & n50859;
  assign n50861 = ~n414 & n50860;
  assign n50862 = ~n271 & n50861;
  assign n50863 = ~n447 & n50862;
  assign n50864 = ~n622 & n50863;
  assign n50865 = n50847 & n50848;
  assign n50866 = n59993 & n60054;
  assign n50867 = ~n59993 & ~n60054;
  assign n50868 = ~n50866 & ~n50867;
  assign n50869 = ~pi11  & n50868;
  assign n50870 = pi11  & ~n50868;
  assign n50871 = ~n50869 & ~n50870;
  assign n50872 = n1576 & n41762;
  assign n50873 = n11215 & n39564;
  assign n50874 = n54403 & n39570;
  assign n50875 = n10564 & n39567;
  assign n50876 = ~n50874 & ~n50875;
  assign n50877 = ~n50873 & n50876;
  assign n50878 = ~n50872 & n50877;
  assign n50879 = n50871 & ~n50878;
  assign n50880 = ~n50871 & n50878;
  assign n50881 = n50871 & ~n50879;
  assign n50882 = n50871 & n50878;
  assign n50883 = ~n50878 & ~n50879;
  assign n50884 = ~n50871 & ~n50878;
  assign n50885 = ~n60055 & ~n60056;
  assign n50886 = ~n50879 & ~n50880;
  assign n50887 = ~n50629 & ~n60057;
  assign n50888 = n50629 & n60057;
  assign n50889 = ~n60057 & ~n50887;
  assign n50890 = n50629 & ~n60057;
  assign n50891 = ~n50629 & ~n50887;
  assign n50892 = ~n50629 & n60057;
  assign n50893 = ~n60058 & ~n60059;
  assign n50894 = ~n50887 & ~n50888;
  assign n50895 = ~n50819 & ~n60060;
  assign n50896 = n50819 & n60060;
  assign n50897 = ~n50819 & ~n50895;
  assign n50898 = ~n60060 & ~n50895;
  assign n50899 = ~n50897 & ~n50898;
  assign n50900 = ~n50895 & ~n50896;
  assign n50901 = n50818 & n60061;
  assign n50902 = ~n50818 & ~n60061;
  assign n50903 = ~n60061 & ~n50902;
  assign n50904 = ~n50818 & ~n50902;
  assign n50905 = ~n50903 & ~n50904;
  assign n50906 = ~n50901 & ~n50902;
  assign n50907 = ~n50805 & ~n60062;
  assign n50908 = n50805 & n60062;
  assign n50909 = ~n60062 & ~n50907;
  assign n50910 = n50805 & ~n60062;
  assign n50911 = ~n50805 & ~n50907;
  assign n50912 = ~n50805 & n60062;
  assign n50913 = ~n60063 & ~n60064;
  assign n50914 = ~n50907 & ~n50908;
  assign n50915 = ~n50651 & n50666;
  assign n50916 = ~n50651 & ~n50667;
  assign n50917 = ~n50652 & ~n50915;
  assign n50918 = n60065 & n60066;
  assign n50919 = ~n60065 & ~n60066;
  assign n50920 = ~n50918 & ~n50919;
  assign n50921 = n90 & n39943;
  assign n50922 = n14236 & n39937;
  assign n50923 = n54667 & n39440;
  assign n50924 = n14210 & n39543;
  assign n50925 = ~n50923 & ~n50924;
  assign n50926 = ~n50922 & n50925;
  assign n50927 = ~n50921 & n50926;
  assign n50928 = pi23  & ~n50927;
  assign n50929 = pi23  & ~n50928;
  assign n50930 = pi23  & n50927;
  assign n50931 = ~n50927 & ~n50928;
  assign n50932 = ~pi23  & ~n50927;
  assign n50933 = ~n60067 & ~n60068;
  assign n50934 = n50920 & ~n50933;
  assign n50935 = ~n50920 & n50933;
  assign n50936 = n50920 & ~n50934;
  assign n50937 = n50920 & n50933;
  assign n50938 = ~n50933 & ~n50934;
  assign n50939 = ~n50920 & ~n50933;
  assign n50940 = ~n60069 & ~n60070;
  assign n50941 = ~n50934 & ~n50935;
  assign n50942 = ~n50677 & n50691;
  assign n50943 = ~n50677 & ~n50693;
  assign n50944 = ~n50676 & ~n50942;
  assign n50945 = n60071 & n60072;
  assign n50946 = ~n60071 & ~n60072;
  assign n50947 = ~n50945 & ~n50946;
  assign n50948 = n14413 & ~n59280;
  assign n50949 = n15921 & n44871;
  assign n50950 = n54719 & n44327;
  assign n50951 = n15901 & n44775;
  assign n50952 = ~n50950 & ~n50951;
  assign n50953 = ~n50949 & n50952;
  assign n50954 = ~n50948 & n50953;
  assign n50955 = pi20  & ~n50954;
  assign n50956 = pi20  & ~n50955;
  assign n50957 = pi20  & n50954;
  assign n50958 = ~n50954 & ~n50955;
  assign n50959 = ~pi20  & ~n50954;
  assign n50960 = ~n60073 & ~n60074;
  assign n50961 = ~n50702 & n50716;
  assign n50962 = ~n50702 & ~n50717;
  assign n50963 = ~n50701 & ~n50961;
  assign n50964 = ~n50960 & ~n60075;
  assign n50965 = n50960 & n60075;
  assign n50966 = ~n60075 & ~n50964;
  assign n50967 = n50960 & ~n60075;
  assign n50968 = ~n50960 & ~n50964;
  assign n50969 = ~n50960 & n60075;
  assign n50970 = ~n60076 & ~n60077;
  assign n50971 = ~n50964 & ~n50965;
  assign n50972 = ~n50947 & n60078;
  assign n50973 = n50947 & ~n60078;
  assign n50974 = ~n50972 & ~n50973;
  assign n50975 = n16079 & n46426;
  assign n50976 = n16696 & n46420;
  assign n50977 = n54886 & n44952;
  assign n50978 = n16676 & n46009;
  assign n50979 = ~n50977 & ~n50978;
  assign n50980 = ~n50976 & n50979;
  assign n50981 = ~n50975 & n50980;
  assign n50982 = pi17  & ~n50981;
  assign n50983 = pi17  & ~n50982;
  assign n50984 = pi17  & n50981;
  assign n50985 = ~n50981 & ~n50982;
  assign n50986 = ~pi17  & ~n50981;
  assign n50987 = ~n60079 & ~n60080;
  assign n50988 = n50974 & ~n50987;
  assign n50989 = ~n50974 & n50987;
  assign n50990 = n50974 & ~n50988;
  assign n50991 = n50974 & n50987;
  assign n50992 = ~n50987 & ~n50988;
  assign n50993 = ~n50974 & ~n50987;
  assign n50994 = ~n60081 & ~n60082;
  assign n50995 = ~n50988 & ~n50989;
  assign n50996 = ~n50727 & n50741;
  assign n50997 = ~n50727 & ~n50743;
  assign n50998 = ~n50726 & ~n50996;
  assign n50999 = n60083 & n60084;
  assign n51000 = ~n60083 & ~n60084;
  assign n51001 = ~n50999 & ~n51000;
  assign n51002 = n17265 & ~n47526;
  assign n51003 = n55041 & n46788;
  assign n51004 = n18556 & n59503;
  assign n51005 = ~n51003 & ~n51004;
  assign n51006 = ~n51002 & n51005;
  assign n51007 = pi14  & ~n51006;
  assign n51008 = pi14  & ~n51007;
  assign n51009 = pi14  & n51006;
  assign n51010 = ~n51006 & ~n51007;
  assign n51011 = ~pi14  & ~n51006;
  assign n51012 = ~n60085 & ~n60086;
  assign n51013 = ~n50752 & n50766;
  assign n51014 = ~n50752 & ~n50767;
  assign n51015 = ~n50751 & ~n51013;
  assign n51016 = ~n51012 & ~n60087;
  assign n51017 = n51012 & n60087;
  assign n51018 = ~n60087 & ~n51016;
  assign n51019 = n51012 & ~n60087;
  assign n51020 = ~n51012 & ~n51016;
  assign n51021 = ~n51012 & n60087;
  assign n51022 = ~n60088 & ~n60089;
  assign n51023 = ~n51016 & ~n51017;
  assign n51024 = ~n51001 & n60090;
  assign n51025 = n51001 & ~n60090;
  assign n51026 = ~n51024 & ~n51025;
  assign n51027 = ~n50546 & n60045;
  assign n51028 = ~n50546 & ~n50773;
  assign n51029 = ~n50547 & ~n51027;
  assign n51030 = n51026 & ~n60091;
  assign n51031 = ~n51026 & n60091;
  assign n51032 = ~n51030 & ~n51031;
  assign n51033 = ~n50792 & n51032;
  assign n51034 = n50792 & ~n51032;
  assign n51035 = ~n51033 & ~n51034;
  assign n51036 = ~n50789 & ~n51035;
  assign n51037 = n50789 & n51035;
  assign po16  = ~n51036 & ~n51037;
  assign n51039 = ~n51030 & ~n51033;
  assign n51040 = ~n51016 & ~n51025;
  assign n51041 = ~n50988 & ~n51000;
  assign n51042 = n16079 & n46805;
  assign n51043 = n16696 & n46788;
  assign n51044 = n54886 & n46009;
  assign n51045 = n16676 & n46420;
  assign n51046 = ~n51044 & ~n51045;
  assign n51047 = ~n51043 & n51046;
  assign n51048 = ~n51042 & n51047;
  assign n51049 = pi17  & ~n51048;
  assign n51050 = pi17  & ~n51049;
  assign n51051 = pi17  & n51048;
  assign n51052 = ~n51048 & ~n51049;
  assign n51053 = ~pi17  & ~n51048;
  assign n51054 = ~n60092 & ~n60093;
  assign n51055 = ~n50964 & ~n50973;
  assign n51056 = ~n50934 & ~n50946;
  assign n51057 = ~n50907 & ~n50919;
  assign n51058 = ~n50879 & ~n50887;
  assign n51059 = ~n50867 & ~n50869;
  assign n51060 = ~n948 & n8865;
  assign n51061 = n3284 & n4013;
  assign n51062 = ~n948 & ~n1485;
  assign n51063 = ~n1044 & n51062;
  assign n51064 = n3062 & n3284;
  assign n51065 = n51063 & n51064;
  assign n51066 = n51060 & n51061;
  assign n51067 = n53589 & n2404;
  assign n51068 = n60094 & n51067;
  assign n51069 = n1076 & n1803;
  assign n51070 = n8453 & n51069;
  assign n51071 = n56604 & n51070;
  assign n51072 = ~n357 & ~n1485;
  assign n51073 = ~n1044 & n51072;
  assign n51074 = ~n259 & ~n948;
  assign n51075 = n1076 & n51074;
  assign n51076 = n51073 & n51075;
  assign n51077 = n51067 & n51076;
  assign n51078 = n1803 & n3062;
  assign n51079 = n8453 & n51078;
  assign n51080 = n56604 & n51079;
  assign n51081 = n51077 & n51080;
  assign n51082 = n51068 & n51071;
  assign n51083 = n59565 & n59666;
  assign n51084 = n59666 & n60095;
  assign n51085 = n59565 & n51084;
  assign n51086 = n60095 & n51083;
  assign n51087 = n56911 & n58422;
  assign n51088 = n53589 & n8453;
  assign n51089 = n1076 & n51088;
  assign n51090 = n2404 & n51089;
  assign n51091 = n56604 & n51090;
  assign n51092 = n59565 & n51091;
  assign n51093 = n58422 & n51092;
  assign n51094 = n56911 & n51093;
  assign n51095 = n59666 & n51094;
  assign n51096 = n1803 & n51095;
  assign n51097 = n3062 & n51096;
  assign n51098 = ~n948 & n51097;
  assign n51099 = ~n1044 & n51098;
  assign n51100 = ~n1485 & n51099;
  assign n51101 = ~n259 & n51100;
  assign n51102 = ~n357 & n51101;
  assign n51103 = n58422 & n60096;
  assign n51104 = n56911 & n51103;
  assign n51105 = n60096 & n51087;
  assign n51106 = ~n51059 & n60097;
  assign n51107 = n51059 & ~n60097;
  assign n51108 = ~n51106 & ~n51107;
  assign n51109 = n1576 & ~n58493;
  assign n51110 = n11215 & n39561;
  assign n51111 = n54403 & n39567;
  assign n51112 = n10564 & n39564;
  assign n51113 = ~n51111 & ~n51112;
  assign n51114 = ~n51110 & n51113;
  assign n51115 = ~n51109 & n51114;
  assign n51116 = n51108 & ~n51115;
  assign n51117 = ~n51108 & n51115;
  assign n51118 = ~n51115 & ~n51116;
  assign n51119 = n51108 & ~n51116;
  assign n51120 = ~n51118 & ~n51119;
  assign n51121 = ~n51116 & ~n51117;
  assign n51122 = n51058 & n60098;
  assign n51123 = ~n51058 & ~n60098;
  assign n51124 = ~n51122 & ~n51123;
  assign n51125 = n11279 & ~n58891;
  assign n51126 = n12584 & n39552;
  assign n51127 = n54410 & n39558;
  assign n51128 = n11267 & n39555;
  assign n51129 = ~n51127 & ~n51128;
  assign n51130 = ~n51126 & n51129;
  assign n51131 = ~n11279 & n51130;
  assign n51132 = n58891 & n51130;
  assign n51133 = ~n51131 & ~n51132;
  assign n51134 = ~n51125 & n51130;
  assign n51135 = pi29  & ~n60099;
  assign n51136 = ~pi29  & n60099;
  assign n51137 = ~n51135 & ~n51136;
  assign n51138 = n51124 & ~n51137;
  assign n51139 = ~n51124 & n51137;
  assign n51140 = ~n51138 & ~n51139;
  assign n51141 = n50818 & ~n50895;
  assign n51142 = ~n50895 & ~n50902;
  assign n51143 = ~n50896 & ~n51141;
  assign n51144 = n51140 & ~n60100;
  assign n51145 = ~n51140 & n60100;
  assign n51146 = ~n51144 & ~n51145;
  assign n51147 = n123 & ~n59050;
  assign n51148 = n128 & n39440;
  assign n51149 = n53444 & n39549;
  assign n51150 = n127 & n39546;
  assign n51151 = ~n51149 & ~n51150;
  assign n51152 = ~n51148 & n51151;
  assign n51153 = ~n51147 & n51152;
  assign n51154 = pi26  & ~n51153;
  assign n51155 = pi26  & ~n51154;
  assign n51156 = pi26  & n51153;
  assign n51157 = ~n51153 & ~n51154;
  assign n51158 = ~pi26  & ~n51153;
  assign n51159 = ~n60101 & ~n60102;
  assign n51160 = n51146 & ~n51159;
  assign n51161 = ~n51146 & n51159;
  assign n51162 = n51146 & ~n51160;
  assign n51163 = ~n51159 & ~n51160;
  assign n51164 = ~n51162 & ~n51163;
  assign n51165 = ~n51160 & ~n51161;
  assign n51166 = n51057 & n60103;
  assign n51167 = ~n51057 & ~n60103;
  assign n51168 = ~n51166 & ~n51167;
  assign n51169 = n90 & ~n59184;
  assign n51170 = n14236 & n44327;
  assign n51171 = n54667 & n39543;
  assign n51172 = n14210 & n39937;
  assign n51173 = ~n51171 & ~n51172;
  assign n51174 = ~n51170 & n51173;
  assign n51175 = ~n51169 & n51174;
  assign n51176 = pi23  & ~n51175;
  assign n51177 = pi23  & ~n51176;
  assign n51178 = pi23  & n51175;
  assign n51179 = ~n51175 & ~n51176;
  assign n51180 = ~pi23  & ~n51175;
  assign n51181 = ~n60104 & ~n60105;
  assign n51182 = ~n51168 & n51181;
  assign n51183 = n51168 & ~n51181;
  assign n51184 = n51168 & ~n51183;
  assign n51185 = ~n51181 & ~n51183;
  assign n51186 = ~n51184 & ~n51185;
  assign n51187 = ~n51182 & ~n51183;
  assign n51188 = n51056 & n60106;
  assign n51189 = ~n51056 & ~n60106;
  assign n51190 = ~n51188 & ~n51189;
  assign n51191 = n14413 & ~n59275;
  assign n51192 = n15921 & n44952;
  assign n51193 = n54719 & n44775;
  assign n51194 = n15901 & n44871;
  assign n51195 = ~n51193 & ~n51194;
  assign n51196 = ~n51192 & n51195;
  assign n51197 = ~n51191 & n51196;
  assign n51198 = pi20  & ~n51197;
  assign n51199 = pi20  & ~n51198;
  assign n51200 = pi20  & n51197;
  assign n51201 = ~n51197 & ~n51198;
  assign n51202 = ~pi20  & ~n51197;
  assign n51203 = ~n60107 & ~n60108;
  assign n51204 = n51190 & ~n51203;
  assign n51205 = ~n51190 & n51203;
  assign n51206 = n51190 & ~n51204;
  assign n51207 = ~n51203 & ~n51204;
  assign n51208 = ~n51206 & ~n51207;
  assign n51209 = ~n51204 & ~n51205;
  assign n51210 = ~n51055 & ~n60109;
  assign n51211 = n51055 & n60109;
  assign n51212 = ~n60109 & ~n51210;
  assign n51213 = n51055 & ~n60109;
  assign n51214 = ~n51055 & ~n51210;
  assign n51215 = ~n51055 & n60109;
  assign n51216 = ~n60110 & ~n60111;
  assign n51217 = ~n51210 & ~n51211;
  assign n51218 = ~n51054 & ~n60112;
  assign n51219 = n51054 & n60112;
  assign n51220 = ~n60112 & ~n51218;
  assign n51221 = ~n51054 & ~n51218;
  assign n51222 = ~n51220 & ~n51221;
  assign n51223 = ~n51218 & ~n51219;
  assign n51224 = n51041 & n60113;
  assign n51225 = ~n51041 & ~n60113;
  assign n51226 = ~n51224 & ~n51225;
  assign n51227 = n55041 & n59503;
  assign n51228 = pi14  & n51227;
  assign n51229 = pi14  & ~n51228;
  assign n51230 = pi14  & ~n51227;
  assign n51231 = n51227 & ~n51228;
  assign n51232 = ~pi14  & n51227;
  assign n51233 = ~n60114 & ~n60115;
  assign n51234 = n51226 & ~n51233;
  assign n51235 = ~n51226 & n51233;
  assign n51236 = n51226 & ~n51234;
  assign n51237 = ~n51233 & ~n51234;
  assign n51238 = ~n51236 & ~n51237;
  assign n51239 = ~n51234 & ~n51235;
  assign n51240 = ~n51040 & ~n60116;
  assign n51241 = n51040 & n60116;
  assign n51242 = ~n60116 & ~n51240;
  assign n51243 = ~n51040 & ~n51240;
  assign n51244 = ~n51242 & ~n51243;
  assign n51245 = ~n51240 & ~n51241;
  assign n51246 = n51039 & n60117;
  assign n51247 = ~n51039 & ~n60117;
  assign n51248 = ~n51246 & ~n51247;
  assign n51249 = n51037 & n51248;
  assign n51250 = ~n51037 & ~n51248;
  assign po17  = ~n51249 & ~n51250;
  assign n51252 = ~n51210 & ~n51218;
  assign n51253 = pi14  & ~n51252;
  assign n51254 = ~pi14  & n51252;
  assign n51255 = ~n51253 & ~n51254;
  assign n51256 = n123 & ~n59044;
  assign n51257 = n128 & n39543;
  assign n51258 = n53444 & n39546;
  assign n51259 = n127 & n39440;
  assign n51260 = ~n51258 & ~n51259;
  assign n51261 = ~n51257 & n51260;
  assign n51262 = ~n51256 & n51261;
  assign n51263 = pi26  & ~n51262;
  assign n51264 = pi26  & ~n51263;
  assign n51265 = pi26  & n51262;
  assign n51266 = ~n51262 & ~n51263;
  assign n51267 = ~pi26  & ~n51262;
  assign n51268 = ~n60118 & ~n60119;
  assign n51269 = n53513 & n53688;
  assign n51270 = n53688 & n54814;
  assign n51271 = n53513 & n51270;
  assign n51272 = n54814 & n51269;
  assign n51273 = n4914 & n9187;
  assign n51274 = n11043 & n51273;
  assign n51275 = ~n141 & ~n444;
  assign n51276 = ~n448 & ~n1486;
  assign n51277 = n51275 & n51276;
  assign n51278 = ~n258 & ~n660;
  assign n51279 = n180 & n51278;
  assign n51280 = n51277 & n51279;
  assign n51281 = n180 & n4914;
  assign n51282 = n180 & n11043;
  assign n51283 = n4914 & n51282;
  assign n51284 = n11043 & n51281;
  assign n51285 = ~n141 & ~n660;
  assign n51286 = ~n444 & ~n1486;
  assign n51287 = n51285 & n51286;
  assign n51288 = ~n258 & ~n448;
  assign n51289 = n9187 & n51288;
  assign n51290 = ~n141 & ~n822;
  assign n51291 = ~n1485 & ~n1486;
  assign n51292 = n51290 & n51291;
  assign n51293 = ~n444 & ~n448;
  assign n51294 = n51278 & n51293;
  assign n51295 = n51292 & n51294;
  assign n51296 = ~n822 & ~n1486;
  assign n51297 = ~n141 & ~n258;
  assign n51298 = n51296 & n51297;
  assign n51299 = ~n444 & ~n660;
  assign n51300 = ~n448 & ~n1485;
  assign n51301 = n51299 & n51300;
  assign n51302 = n51298 & n51301;
  assign n51303 = n51287 & n51289;
  assign n51304 = n60121 & n60122;
  assign n51305 = n51274 & n51280;
  assign n51306 = n54189 & n54380;
  assign n51307 = n60123 & n51306;
  assign n51308 = n54257 & n51307;
  assign n51309 = n60120 & n51308;
  assign n51310 = n4914 & n54189;
  assign n51311 = n11043 & n51310;
  assign n51312 = n54487 & n51311;
  assign n51313 = n54380 & n51312;
  assign n51314 = n53513 & n51313;
  assign n51315 = n53688 & n51314;
  assign n51316 = n54257 & n51315;
  assign n51317 = n54814 & n51316;
  assign n51318 = n180 & n51317;
  assign n51319 = ~n1486 & n51318;
  assign n51320 = ~n1485 & n51319;
  assign n51321 = ~n258 & n51320;
  assign n51322 = ~n141 & n51321;
  assign n51323 = ~n660 & n51322;
  assign n51324 = ~n822 & n51323;
  assign n51325 = ~n444 & n51324;
  assign n51326 = ~n448 & n51325;
  assign n51327 = n54487 & n51309;
  assign n51328 = ~n60097 & n60124;
  assign n51329 = n60097 & ~n60124;
  assign n51330 = ~n51328 & ~n51329;
  assign n51331 = n1576 & ~n58849;
  assign n51332 = n11215 & n39558;
  assign n51333 = n54403 & n39564;
  assign n51334 = n10564 & n39561;
  assign n51335 = ~n51333 & ~n51334;
  assign n51336 = ~n51332 & n51335;
  assign n51337 = ~n51331 & n51336;
  assign n51338 = ~n51329 & ~n51337;
  assign n51339 = ~n51328 & n51338;
  assign n51340 = n51330 & ~n51337;
  assign n51341 = ~n51330 & n51337;
  assign n51342 = ~n51337 & ~n60125;
  assign n51343 = ~n51329 & ~n60125;
  assign n51344 = ~n51328 & n51343;
  assign n51345 = ~n51342 & ~n51344;
  assign n51346 = ~n60125 & ~n51341;
  assign n51347 = ~n51106 & n51115;
  assign n51348 = ~n51106 & ~n51116;
  assign n51349 = ~n51107 & ~n51347;
  assign n51350 = n60126 & n60127;
  assign n51351 = ~n60126 & ~n60127;
  assign n51352 = ~n51350 & ~n51351;
  assign n51353 = ~n51123 & ~n51138;
  assign n51354 = ~n51352 & n51353;
  assign n51355 = n51352 & ~n51353;
  assign n51356 = ~n51354 & ~n51355;
  assign n51357 = n11279 & ~n58889;
  assign n51358 = n12584 & n39549;
  assign n51359 = n54410 & n39555;
  assign n51360 = n11267 & n39552;
  assign n51361 = ~n51359 & ~n51360;
  assign n51362 = ~n51358 & n51361;
  assign n51363 = ~n51357 & n51362;
  assign n51364 = pi29  & ~n51363;
  assign n51365 = pi29  & ~n51364;
  assign n51366 = pi29  & n51363;
  assign n51367 = ~n51363 & ~n51364;
  assign n51368 = ~pi29  & ~n51363;
  assign n51369 = ~n60128 & ~n60129;
  assign n51370 = n51356 & ~n51369;
  assign n51371 = ~n51356 & n51369;
  assign n51372 = n51356 & ~n51370;
  assign n51373 = n51356 & n51369;
  assign n51374 = ~n51369 & ~n51370;
  assign n51375 = ~n51356 & ~n51369;
  assign n51376 = ~n60130 & ~n60131;
  assign n51377 = ~n51370 & ~n51371;
  assign n51378 = ~n51268 & ~n60132;
  assign n51379 = n51268 & n60132;
  assign n51380 = ~n60132 & ~n51378;
  assign n51381 = ~n51268 & ~n51378;
  assign n51382 = ~n51380 & ~n51381;
  assign n51383 = ~n51378 & ~n51379;
  assign n51384 = ~n51144 & n51159;
  assign n51385 = ~n51144 & ~n51160;
  assign n51386 = ~n51145 & ~n51384;
  assign n51387 = n60133 & n60134;
  assign n51388 = ~n60133 & ~n60134;
  assign n51389 = ~n51387 & ~n51388;
  assign n51390 = n90 & ~n59282;
  assign n51391 = n14236 & n44775;
  assign n51392 = n54667 & n39937;
  assign n51393 = n14210 & n44327;
  assign n51394 = ~n51392 & ~n51393;
  assign n51395 = ~n51391 & n51394;
  assign n51396 = ~n51390 & n51395;
  assign n51397 = pi23  & ~n51396;
  assign n51398 = pi23  & ~n51397;
  assign n51399 = pi23  & n51396;
  assign n51400 = ~n51396 & ~n51397;
  assign n51401 = ~pi23  & ~n51396;
  assign n51402 = ~n60135 & ~n60136;
  assign n51403 = n51389 & ~n51402;
  assign n51404 = ~n51389 & n51402;
  assign n51405 = n51389 & ~n51403;
  assign n51406 = ~n51402 & ~n51403;
  assign n51407 = ~n51405 & ~n51406;
  assign n51408 = ~n51403 & ~n51404;
  assign n51409 = ~n51167 & n51181;
  assign n51410 = ~n51167 & ~n51183;
  assign n51411 = ~n51166 & ~n51409;
  assign n51412 = n60137 & n60138;
  assign n51413 = ~n60137 & ~n60138;
  assign n51414 = ~n51412 & ~n51413;
  assign n51415 = n14413 & ~n59386;
  assign n51416 = n15921 & n46009;
  assign n51417 = n54719 & n44871;
  assign n51418 = n15901 & n44952;
  assign n51419 = ~n51417 & ~n51418;
  assign n51420 = ~n51416 & n51419;
  assign n51421 = ~n51415 & n51420;
  assign n51422 = pi20  & ~n51421;
  assign n51423 = pi20  & ~n51422;
  assign n51424 = pi20  & n51421;
  assign n51425 = ~n51421 & ~n51422;
  assign n51426 = ~pi20  & ~n51421;
  assign n51427 = ~n60139 & ~n60140;
  assign n51428 = ~n51414 & n51427;
  assign n51429 = n51414 & ~n51427;
  assign n51430 = n51414 & ~n51429;
  assign n51431 = ~n51427 & ~n51429;
  assign n51432 = ~n51430 & ~n51431;
  assign n51433 = ~n51428 & ~n51429;
  assign n51434 = ~n51189 & n51203;
  assign n51435 = ~n51189 & ~n51204;
  assign n51436 = ~n51188 & ~n51434;
  assign n51437 = n60141 & n60142;
  assign n51438 = ~n60141 & ~n60142;
  assign n51439 = ~n51437 & ~n51438;
  assign n51440 = n16079 & ~n59554;
  assign n51441 = n16696 & n59503;
  assign n51442 = n54886 & n46420;
  assign n51443 = n16676 & n46788;
  assign n51444 = ~n51442 & ~n51443;
  assign n51445 = ~n51441 & n51444;
  assign n51446 = ~n51440 & n51445;
  assign n51447 = pi17  & ~n51446;
  assign n51448 = pi17  & ~n51447;
  assign n51449 = pi17  & n51446;
  assign n51450 = ~n51446 & ~n51447;
  assign n51451 = ~pi17  & ~n51446;
  assign n51452 = ~n60143 & ~n60144;
  assign n51453 = n51439 & ~n51452;
  assign n51454 = ~n51439 & n51452;
  assign n51455 = n51439 & ~n51453;
  assign n51456 = ~n51452 & ~n51453;
  assign n51457 = ~n51455 & ~n51456;
  assign n51458 = ~n51453 & ~n51454;
  assign n51459 = n51255 & ~n60145;
  assign n51460 = ~n51255 & n60145;
  assign n51461 = ~n60145 & ~n51459;
  assign n51462 = n51255 & ~n51459;
  assign n51463 = ~n51461 & ~n51462;
  assign n51464 = ~n51459 & ~n51460;
  assign n51465 = ~n51225 & n51233;
  assign n51466 = ~n51225 & ~n51234;
  assign n51467 = ~n51224 & ~n51465;
  assign n51468 = n60146 & n60147;
  assign n51469 = ~n60146 & ~n60147;
  assign n51470 = ~n51468 & ~n51469;
  assign n51471 = ~n51240 & ~n51247;
  assign n51472 = ~n51470 & n51471;
  assign n51473 = n51470 & ~n51471;
  assign n51474 = ~n51472 & ~n51473;
  assign n51475 = n51249 & n51474;
  assign n51476 = ~n51249 & ~n51474;
  assign po18  = ~n51475 & ~n51476;
  assign n51478 = ~n51469 & ~n51473;
  assign n51479 = ~n51370 & ~n51378;
  assign n51480 = ~n51351 & ~n51355;
  assign n51481 = n11279 & n43436;
  assign n51482 = n12584 & n39546;
  assign n51483 = n54410 & n39552;
  assign n51484 = n11267 & n39549;
  assign n51485 = ~n51483 & ~n51484;
  assign n51486 = ~n51482 & n51485;
  assign n51487 = ~n51481 & n51486;
  assign n51488 = pi29  & ~n51487;
  assign n51489 = pi29  & ~n51488;
  assign n51490 = pi29  & n51487;
  assign n51491 = ~n51487 & ~n51488;
  assign n51492 = ~pi29  & ~n51487;
  assign n51493 = ~n60148 & ~n60149;
  assign n51494 = n53777 & n54272;
  assign n51495 = n54477 & n51494;
  assign n51496 = ~n405 & ~n1658;
  assign n51497 = ~n660 & n51496;
  assign n51498 = ~n1658 & n4095;
  assign n51499 = n1672 & n7755;
  assign n51500 = n60150 & n51499;
  assign n51501 = n56725 & n51500;
  assign n51502 = n51495 & n51501;
  assign n51503 = n53925 & n55147;
  assign n51504 = n51502 & n51503;
  assign n51505 = n56679 & n51504;
  assign n51506 = n54272 & n54477;
  assign n51507 = n56725 & n51506;
  assign n51508 = n7755 & n51507;
  assign n51509 = n56679 & n51508;
  assign n51510 = n55147 & n51509;
  assign n51511 = n53986 & n51510;
  assign n51512 = n53925 & n51511;
  assign n51513 = n1672 & n51512;
  assign n51514 = n53777 & n51513;
  assign n51515 = ~n660 & n51514;
  assign n51516 = ~n405 & n51515;
  assign n51517 = ~n1658 & n51516;
  assign n51518 = n53986 & n51505;
  assign n51519 = n60097 & n60151;
  assign n51520 = ~n60097 & ~n60151;
  assign n51521 = ~n51519 & ~n51520;
  assign n51522 = ~pi14  & n51521;
  assign n51523 = pi14  & ~n51521;
  assign n51524 = ~n51522 & ~n51523;
  assign n51525 = ~n51343 & n51524;
  assign n51526 = n51343 & ~n51524;
  assign n51527 = ~n51525 & ~n51526;
  assign n51528 = n1576 & n42574;
  assign n51529 = n11215 & n39555;
  assign n51530 = n54403 & n39561;
  assign n51531 = n10564 & n39558;
  assign n51532 = ~n51530 & ~n51531;
  assign n51533 = ~n51529 & n51532;
  assign n51534 = ~n51528 & n51533;
  assign n51535 = n51527 & ~n51534;
  assign n51536 = ~n51527 & n51534;
  assign n51537 = n51527 & ~n51535;
  assign n51538 = ~n51534 & ~n51535;
  assign n51539 = ~n51537 & ~n51538;
  assign n51540 = ~n51535 & ~n51536;
  assign n51541 = ~n51493 & ~n60152;
  assign n51542 = n51493 & n60152;
  assign n51543 = ~n60152 & ~n51541;
  assign n51544 = ~n51493 & ~n51541;
  assign n51545 = ~n51543 & ~n51544;
  assign n51546 = ~n51541 & ~n51542;
  assign n51547 = n51480 & n60153;
  assign n51548 = ~n51480 & ~n60153;
  assign n51549 = ~n51547 & ~n51548;
  assign n51550 = n123 & n39943;
  assign n51551 = n128 & n39937;
  assign n51552 = n53444 & n39440;
  assign n51553 = n127 & n39543;
  assign n51554 = ~n51552 & ~n51553;
  assign n51555 = ~n51551 & n51554;
  assign n51556 = ~n51550 & n51555;
  assign n51557 = pi26  & ~n51556;
  assign n51558 = pi26  & ~n51557;
  assign n51559 = pi26  & n51556;
  assign n51560 = ~n51556 & ~n51557;
  assign n51561 = ~pi26  & ~n51556;
  assign n51562 = ~n60154 & ~n60155;
  assign n51563 = n51549 & ~n51562;
  assign n51564 = ~n51549 & n51562;
  assign n51565 = n51549 & ~n51563;
  assign n51566 = n51549 & n51562;
  assign n51567 = ~n51562 & ~n51563;
  assign n51568 = ~n51549 & ~n51562;
  assign n51569 = ~n60156 & ~n60157;
  assign n51570 = ~n51563 & ~n51564;
  assign n51571 = n51479 & n60158;
  assign n51572 = ~n51479 & ~n60158;
  assign n51573 = ~n51571 & ~n51572;
  assign n51574 = n90 & ~n59280;
  assign n51575 = n14236 & n44871;
  assign n51576 = n54667 & n44327;
  assign n51577 = n14210 & n44775;
  assign n51578 = ~n51576 & ~n51577;
  assign n51579 = ~n51575 & n51578;
  assign n51580 = ~n51574 & n51579;
  assign n51581 = pi23  & ~n51580;
  assign n51582 = pi23  & ~n51581;
  assign n51583 = pi23  & n51580;
  assign n51584 = ~n51580 & ~n51581;
  assign n51585 = ~pi23  & ~n51580;
  assign n51586 = ~n60159 & ~n60160;
  assign n51587 = ~n51388 & n51402;
  assign n51588 = ~n51388 & ~n51403;
  assign n51589 = ~n51387 & ~n51587;
  assign n51590 = ~n51586 & ~n60161;
  assign n51591 = n51586 & n60161;
  assign n51592 = ~n60161 & ~n51590;
  assign n51593 = n51586 & ~n60161;
  assign n51594 = ~n51586 & ~n51590;
  assign n51595 = ~n51586 & n60161;
  assign n51596 = ~n60162 & ~n60163;
  assign n51597 = ~n51590 & ~n51591;
  assign n51598 = ~n51573 & n60164;
  assign n51599 = n51573 & ~n60164;
  assign n51600 = ~n51598 & ~n51599;
  assign n51601 = n14413 & n46426;
  assign n51602 = n15921 & n46420;
  assign n51603 = n54719 & n44952;
  assign n51604 = n15901 & n46009;
  assign n51605 = ~n51603 & ~n51604;
  assign n51606 = ~n51602 & n51605;
  assign n51607 = ~n51601 & n51606;
  assign n51608 = pi20  & ~n51607;
  assign n51609 = pi20  & ~n51608;
  assign n51610 = pi20  & n51607;
  assign n51611 = ~n51607 & ~n51608;
  assign n51612 = ~pi20  & ~n51607;
  assign n51613 = ~n60165 & ~n60166;
  assign n51614 = n51600 & ~n51613;
  assign n51615 = ~n51600 & n51613;
  assign n51616 = n51600 & ~n51614;
  assign n51617 = n51600 & n51613;
  assign n51618 = ~n51613 & ~n51614;
  assign n51619 = ~n51600 & ~n51613;
  assign n51620 = ~n60167 & ~n60168;
  assign n51621 = ~n51614 & ~n51615;
  assign n51622 = ~n51413 & n51427;
  assign n51623 = ~n51413 & ~n51429;
  assign n51624 = ~n51412 & ~n51622;
  assign n51625 = n60169 & n60170;
  assign n51626 = ~n60169 & ~n60170;
  assign n51627 = ~n51625 & ~n51626;
  assign n51628 = n16079 & ~n47526;
  assign n51629 = n54886 & n46788;
  assign n51630 = n16676 & n59503;
  assign n51631 = ~n51629 & ~n51630;
  assign n51632 = ~n51628 & n51631;
  assign n51633 = pi17  & ~n51632;
  assign n51634 = pi17  & ~n51633;
  assign n51635 = pi17  & n51632;
  assign n51636 = ~n51632 & ~n51633;
  assign n51637 = ~pi17  & ~n51632;
  assign n51638 = ~n60171 & ~n60172;
  assign n51639 = ~n51438 & n51452;
  assign n51640 = ~n51438 & ~n51453;
  assign n51641 = ~n51437 & ~n51639;
  assign n51642 = ~n51638 & ~n60173;
  assign n51643 = n51638 & n60173;
  assign n51644 = ~n60173 & ~n51642;
  assign n51645 = n51638 & ~n60173;
  assign n51646 = ~n51638 & ~n51642;
  assign n51647 = ~n51638 & n60173;
  assign n51648 = ~n60174 & ~n60175;
  assign n51649 = ~n51642 & ~n51643;
  assign n51650 = ~n51627 & n60176;
  assign n51651 = n51627 & ~n60176;
  assign n51652 = ~n51650 & ~n51651;
  assign n51653 = ~n51253 & n60145;
  assign n51654 = ~n51253 & ~n51459;
  assign n51655 = ~n51254 & ~n51653;
  assign n51656 = n51652 & ~n60177;
  assign n51657 = ~n51652 & n60177;
  assign n51658 = ~n51656 & ~n51657;
  assign n51659 = ~n51478 & n51658;
  assign n51660 = n51478 & ~n51658;
  assign n51661 = ~n51659 & ~n51660;
  assign n51662 = ~n51475 & ~n51661;
  assign n51663 = n51475 & n51661;
  assign po19  = ~n51662 & ~n51663;
  assign n51665 = ~n51656 & ~n51659;
  assign n51666 = ~n51642 & ~n51651;
  assign n51667 = ~n51614 & ~n51626;
  assign n51668 = n14413 & n46805;
  assign n51669 = n15921 & n46788;
  assign n51670 = n54719 & n46009;
  assign n51671 = n15901 & n46420;
  assign n51672 = ~n51670 & ~n51671;
  assign n51673 = ~n51669 & n51672;
  assign n51674 = ~n51668 & n51673;
  assign n51675 = pi20  & ~n51674;
  assign n51676 = pi20  & ~n51675;
  assign n51677 = pi20  & n51674;
  assign n51678 = ~n51674 & ~n51675;
  assign n51679 = ~pi20  & ~n51674;
  assign n51680 = ~n60178 & ~n60179;
  assign n51681 = ~n51590 & ~n51599;
  assign n51682 = ~n51563 & ~n51572;
  assign n51683 = ~n51541 & ~n51548;
  assign n51684 = ~n51520 & ~n51522;
  assign n51685 = ~n750 & ~n1061;
  assign n51686 = n3082 & n51685;
  assign n51687 = n3134 & n5652;
  assign n51688 = n3082 & n5652;
  assign n51689 = n3134 & n51685;
  assign n51690 = n51688 & n51689;
  assign n51691 = n51686 & n51687;
  assign n51692 = n54026 & n43236;
  assign n51693 = n43236 & n51688;
  assign n51694 = n54026 & n51689;
  assign n51695 = n51693 & n51694;
  assign n51696 = n60180 & n51692;
  assign n51697 = n1067 & n7646;
  assign n51698 = n30933 & n51697;
  assign n51699 = n53691 & n51698;
  assign n51700 = n5652 & n7646;
  assign n51701 = n358 & n1067;
  assign n51702 = n51700 & n51701;
  assign n51703 = ~n409 & ~n750;
  assign n51704 = ~n207 & ~n1061;
  assign n51705 = n51703 & n51704;
  assign n51706 = n54026 & n51705;
  assign n51707 = n51702 & n51706;
  assign n51708 = n1578 & n3082;
  assign n51709 = n3134 & n51708;
  assign n51710 = n53691 & n51709;
  assign n51711 = n51707 & n51710;
  assign n51712 = n60181 & n51699;
  assign n51713 = n54939 & n56742;
  assign n51714 = n60182 & n51713;
  assign n51715 = n54777 & n51714;
  assign n51716 = n53691 & n54026;
  assign n51717 = n3134 & n51716;
  assign n51718 = n56742 & n51717;
  assign n51719 = n54777 & n51718;
  assign n51720 = n54939 & n51719;
  assign n51721 = n5652 & n51720;
  assign n51722 = n3082 & n51721;
  assign n51723 = n1067 & n51722;
  assign n51724 = n1578 & n51723;
  assign n51725 = n54331 & n51724;
  assign n51726 = n358 & n51725;
  assign n51727 = n7646 & n51726;
  assign n51728 = ~n1061 & n51727;
  assign n51729 = ~n207 & n51728;
  assign n51730 = ~n409 & n51729;
  assign n51731 = ~n750 & n51730;
  assign n51732 = n54331 & n51715;
  assign n51733 = ~n51684 & n60183;
  assign n51734 = n51684 & ~n60183;
  assign n51735 = ~n51733 & ~n51734;
  assign n51736 = n1576 & ~n58891;
  assign n51737 = n11215 & n39552;
  assign n51738 = n54403 & n39558;
  assign n51739 = n10564 & n39555;
  assign n51740 = ~n51738 & ~n51739;
  assign n51741 = ~n51737 & n51740;
  assign n51742 = ~n51736 & n51741;
  assign n51743 = n51735 & ~n51742;
  assign n51744 = ~n51735 & n51742;
  assign n51745 = ~n51742 & ~n51743;
  assign n51746 = n51735 & ~n51743;
  assign n51747 = ~n51745 & ~n51746;
  assign n51748 = ~n51743 & ~n51744;
  assign n51749 = ~n51525 & n51534;
  assign n51750 = ~n51525 & ~n51535;
  assign n51751 = ~n51526 & ~n51749;
  assign n51752 = n60184 & n60185;
  assign n51753 = ~n60184 & ~n60185;
  assign n51754 = ~n51752 & ~n51753;
  assign n51755 = n11279 & ~n59050;
  assign n51756 = n12584 & n39440;
  assign n51757 = n54410 & n39549;
  assign n51758 = n11267 & n39546;
  assign n51759 = ~n51757 & ~n51758;
  assign n51760 = ~n51756 & n51759;
  assign n51761 = ~n11279 & n51760;
  assign n51762 = n59050 & n51760;
  assign n51763 = ~n51761 & ~n51762;
  assign n51764 = ~n51755 & n51760;
  assign n51765 = pi29  & ~n60186;
  assign n51766 = ~pi29  & n60186;
  assign n51767 = ~n51765 & ~n51766;
  assign n51768 = n51754 & ~n51767;
  assign n51769 = ~n51754 & n51767;
  assign n51770 = ~n51768 & ~n51769;
  assign n51771 = ~n51683 & n51770;
  assign n51772 = n51683 & ~n51770;
  assign n51773 = ~n51771 & ~n51772;
  assign n51774 = n123 & ~n59184;
  assign n51775 = n128 & n44327;
  assign n51776 = n53444 & n39543;
  assign n51777 = n127 & n39937;
  assign n51778 = ~n51776 & ~n51777;
  assign n51779 = ~n51775 & n51778;
  assign n51780 = ~n51774 & n51779;
  assign n51781 = pi26  & ~n51780;
  assign n51782 = pi26  & ~n51781;
  assign n51783 = pi26  & n51780;
  assign n51784 = ~n51780 & ~n51781;
  assign n51785 = ~pi26  & ~n51780;
  assign n51786 = ~n60187 & ~n60188;
  assign n51787 = n51773 & ~n51786;
  assign n51788 = ~n51773 & n51786;
  assign n51789 = n51773 & ~n51787;
  assign n51790 = ~n51786 & ~n51787;
  assign n51791 = ~n51789 & ~n51790;
  assign n51792 = ~n51787 & ~n51788;
  assign n51793 = n51682 & n60189;
  assign n51794 = ~n51682 & ~n60189;
  assign n51795 = ~n51793 & ~n51794;
  assign n51796 = n90 & ~n59275;
  assign n51797 = n14236 & n44952;
  assign n51798 = n54667 & n44775;
  assign n51799 = n14210 & n44871;
  assign n51800 = ~n51798 & ~n51799;
  assign n51801 = ~n51797 & n51800;
  assign n51802 = ~n51796 & n51801;
  assign n51803 = pi23  & ~n51802;
  assign n51804 = pi23  & ~n51803;
  assign n51805 = pi23  & n51802;
  assign n51806 = ~n51802 & ~n51803;
  assign n51807 = ~pi23  & ~n51802;
  assign n51808 = ~n60190 & ~n60191;
  assign n51809 = ~n51795 & n51808;
  assign n51810 = n51795 & ~n51808;
  assign n51811 = n51795 & ~n51810;
  assign n51812 = ~n51808 & ~n51810;
  assign n51813 = ~n51811 & ~n51812;
  assign n51814 = ~n51809 & ~n51810;
  assign n51815 = ~n51681 & ~n60192;
  assign n51816 = n51681 & n60192;
  assign n51817 = ~n60192 & ~n51815;
  assign n51818 = n51681 & ~n60192;
  assign n51819 = ~n51681 & ~n51815;
  assign n51820 = ~n51681 & n60192;
  assign n51821 = ~n60193 & ~n60194;
  assign n51822 = ~n51815 & ~n51816;
  assign n51823 = ~n51680 & ~n60195;
  assign n51824 = n51680 & n60195;
  assign n51825 = ~n60195 & ~n51823;
  assign n51826 = ~n51680 & ~n51823;
  assign n51827 = ~n51825 & ~n51826;
  assign n51828 = ~n51823 & ~n51824;
  assign n51829 = n51667 & n60196;
  assign n51830 = ~n51667 & ~n60196;
  assign n51831 = ~n51829 & ~n51830;
  assign n51832 = n54886 & n59503;
  assign n51833 = pi17  & n51832;
  assign n51834 = pi17  & ~n51833;
  assign n51835 = pi17  & ~n51832;
  assign n51836 = n51832 & ~n51833;
  assign n51837 = ~pi17  & n51832;
  assign n51838 = ~n60197 & ~n60198;
  assign n51839 = n51831 & ~n51838;
  assign n51840 = ~n51831 & n51838;
  assign n51841 = n51831 & ~n51839;
  assign n51842 = ~n51838 & ~n51839;
  assign n51843 = ~n51841 & ~n51842;
  assign n51844 = ~n51839 & ~n51840;
  assign n51845 = ~n51666 & ~n60199;
  assign n51846 = n51666 & n60199;
  assign n51847 = ~n60199 & ~n51845;
  assign n51848 = ~n51666 & ~n51845;
  assign n51849 = ~n51847 & ~n51848;
  assign n51850 = ~n51845 & ~n51846;
  assign n51851 = n51665 & n60200;
  assign n51852 = ~n51665 & ~n60200;
  assign n51853 = ~n51851 & ~n51852;
  assign n51854 = n51663 & n51853;
  assign n51855 = ~n51663 & ~n51853;
  assign po20  = ~n51854 & ~n51855;
  assign n51857 = ~n51815 & ~n51823;
  assign n51858 = pi17  & ~n51857;
  assign n51859 = ~pi17  & n51857;
  assign n51860 = ~n51858 & ~n51859;
  assign n51861 = ~n51753 & ~n51768;
  assign n51862 = n11279 & ~n59044;
  assign n51863 = n12584 & n39543;
  assign n51864 = n54410 & n39546;
  assign n51865 = n11267 & n39440;
  assign n51866 = ~n51864 & ~n51865;
  assign n51867 = ~n51863 & n51866;
  assign n51868 = ~n11279 & n51867;
  assign n51869 = n59044 & n51867;
  assign n51870 = ~n51868 & ~n51869;
  assign n51871 = ~n51862 & n51867;
  assign n51872 = pi29  & ~n60201;
  assign n51873 = ~pi29  & n60201;
  assign n51874 = ~n51872 & ~n51873;
  assign n51875 = ~n414 & ~n1680;
  assign n51876 = ~n414 & n6150;
  assign n51877 = ~n1680 & n51876;
  assign n51878 = n6150 & n51875;
  assign n51879 = ~n646 & ~n829;
  assign n51880 = ~n776 & ~n922;
  assign n51881 = ~n646 & ~n776;
  assign n51882 = ~n829 & ~n922;
  assign n51883 = n51881 & n51882;
  assign n51884 = n51879 & n51880;
  assign n51885 = n4013 & n4212;
  assign n51886 = n60203 & n51885;
  assign n51887 = n60202 & n51886;
  assign n51888 = n1803 & n4512;
  assign n51889 = n586 & n8196;
  assign n51890 = n51888 & n51889;
  assign n51891 = n53665 & n51890;
  assign n51892 = n54259 & n51891;
  assign n51893 = n4212 & n4512;
  assign n51894 = n60203 & n51893;
  assign n51895 = n60202 & n51894;
  assign n51896 = n586 & n1803;
  assign n51897 = n4013 & n8196;
  assign n51898 = n51896 & n51897;
  assign n51899 = n54259 & n51898;
  assign n51900 = n53665 & n51899;
  assign n51901 = n51895 & n51900;
  assign n51902 = n51887 & n51892;
  assign n51903 = n54395 & n60204;
  assign n51904 = n53961 & n54808;
  assign n51905 = n4212 & n8196;
  assign n51906 = n60202 & n51905;
  assign n51907 = n4013 & n51906;
  assign n51908 = n54808 & n51907;
  assign n51909 = n54395 & n51908;
  assign n51910 = n53961 & n51909;
  assign n51911 = n54259 & n51910;
  assign n51912 = n586 & n51911;
  assign n51913 = n53665 & n51912;
  assign n51914 = n1803 & n51913;
  assign n51915 = ~n922 & n51914;
  assign n51916 = ~n272 & n51915;
  assign n51917 = ~n829 & n51916;
  assign n51918 = ~n733 & n51917;
  assign n51919 = ~n646 & n51918;
  assign n51920 = ~n776 & n51919;
  assign n51921 = n51903 & n51904;
  assign n51922 = n60183 & ~n60205;
  assign n51923 = ~n60183 & n60205;
  assign n51924 = ~n51922 & ~n51923;
  assign n51925 = ~n51733 & n51742;
  assign n51926 = ~n51733 & ~n51743;
  assign n51927 = ~n51734 & ~n51925;
  assign n51928 = ~n51923 & ~n60206;
  assign n51929 = ~n51922 & n51928;
  assign n51930 = n51924 & ~n60206;
  assign n51931 = ~n51924 & n60206;
  assign n51932 = ~n60206 & ~n60207;
  assign n51933 = ~n51923 & ~n60207;
  assign n51934 = ~n51922 & n51933;
  assign n51935 = ~n51932 & ~n51934;
  assign n51936 = ~n60207 & ~n51931;
  assign n51937 = n1576 & ~n58889;
  assign n51938 = n11215 & n39549;
  assign n51939 = n54403 & n39555;
  assign n51940 = n10564 & n39552;
  assign n51941 = ~n51939 & ~n51940;
  assign n51942 = ~n51938 & n51941;
  assign n51943 = ~n51937 & n51942;
  assign n51944 = ~n60208 & ~n51943;
  assign n51945 = n60208 & n51943;
  assign n51946 = ~n60208 & ~n51944;
  assign n51947 = ~n60208 & n51943;
  assign n51948 = ~n51943 & ~n51944;
  assign n51949 = n60208 & ~n51943;
  assign n51950 = ~n60209 & ~n60210;
  assign n51951 = ~n51944 & ~n51945;
  assign n51952 = ~n51874 & ~n60211;
  assign n51953 = n51874 & n60211;
  assign n51954 = ~n51952 & ~n51953;
  assign n51955 = ~n51861 & n51954;
  assign n51956 = n51861 & ~n51954;
  assign n51957 = ~n51955 & ~n51956;
  assign n51958 = n123 & ~n59282;
  assign n51959 = n128 & n44775;
  assign n51960 = n53444 & n39937;
  assign n51961 = n127 & n44327;
  assign n51962 = ~n51960 & ~n51961;
  assign n51963 = ~n51959 & n51962;
  assign n51964 = ~n51958 & n51963;
  assign n51965 = pi26  & ~n51964;
  assign n51966 = pi26  & ~n51965;
  assign n51967 = pi26  & n51964;
  assign n51968 = ~n51964 & ~n51965;
  assign n51969 = ~pi26  & ~n51964;
  assign n51970 = ~n60212 & ~n60213;
  assign n51971 = n51957 & ~n51970;
  assign n51972 = ~n51957 & n51970;
  assign n51973 = n51957 & ~n51971;
  assign n51974 = ~n51970 & ~n51971;
  assign n51975 = ~n51973 & ~n51974;
  assign n51976 = ~n51971 & ~n51972;
  assign n51977 = ~n51771 & n51786;
  assign n51978 = ~n51771 & ~n51787;
  assign n51979 = ~n51772 & ~n51977;
  assign n51980 = n60214 & n60215;
  assign n51981 = ~n60214 & ~n60215;
  assign n51982 = ~n51980 & ~n51981;
  assign n51983 = n90 & ~n59386;
  assign n51984 = n14236 & n46009;
  assign n51985 = n54667 & n44871;
  assign n51986 = n14210 & n44952;
  assign n51987 = ~n51985 & ~n51986;
  assign n51988 = ~n51984 & n51987;
  assign n51989 = ~n51983 & n51988;
  assign n51990 = pi23  & ~n51989;
  assign n51991 = pi23  & ~n51990;
  assign n51992 = pi23  & n51989;
  assign n51993 = ~n51989 & ~n51990;
  assign n51994 = ~pi23  & ~n51989;
  assign n51995 = ~n60216 & ~n60217;
  assign n51996 = ~n51982 & n51995;
  assign n51997 = n51982 & ~n51995;
  assign n51998 = n51982 & ~n51997;
  assign n51999 = ~n51995 & ~n51997;
  assign n52000 = ~n51998 & ~n51999;
  assign n52001 = ~n51996 & ~n51997;
  assign n52002 = ~n51794 & n51808;
  assign n52003 = ~n51794 & ~n51810;
  assign n52004 = ~n51793 & ~n52002;
  assign n52005 = n60218 & n60219;
  assign n52006 = ~n60218 & ~n60219;
  assign n52007 = ~n52005 & ~n52006;
  assign n52008 = n14413 & ~n59554;
  assign n52009 = n15921 & n59503;
  assign n52010 = n54719 & n46420;
  assign n52011 = n15901 & n46788;
  assign n52012 = ~n52010 & ~n52011;
  assign n52013 = ~n52009 & n52012;
  assign n52014 = ~n52008 & n52013;
  assign n52015 = pi20  & ~n52014;
  assign n52016 = pi20  & ~n52015;
  assign n52017 = pi20  & n52014;
  assign n52018 = ~n52014 & ~n52015;
  assign n52019 = ~pi20  & ~n52014;
  assign n52020 = ~n60220 & ~n60221;
  assign n52021 = n52007 & ~n52020;
  assign n52022 = ~n52007 & n52020;
  assign n52023 = n52007 & ~n52021;
  assign n52024 = ~n52020 & ~n52021;
  assign n52025 = ~n52023 & ~n52024;
  assign n52026 = ~n52021 & ~n52022;
  assign n52027 = n51860 & ~n60222;
  assign n52028 = ~n51860 & n60222;
  assign n52029 = ~n60222 & ~n52027;
  assign n52030 = n51860 & ~n52027;
  assign n52031 = ~n52029 & ~n52030;
  assign n52032 = ~n52027 & ~n52028;
  assign n52033 = ~n51830 & n51838;
  assign n52034 = ~n51830 & ~n51839;
  assign n52035 = ~n51829 & ~n52033;
  assign n52036 = n60223 & n60224;
  assign n52037 = ~n60223 & ~n60224;
  assign n52038 = ~n52036 & ~n52037;
  assign n52039 = ~n51845 & ~n51852;
  assign n52040 = ~n52038 & n52039;
  assign n52041 = n52038 & ~n52039;
  assign n52042 = ~n52040 & ~n52041;
  assign n52043 = n51854 & n52042;
  assign n52044 = ~n51854 & ~n52042;
  assign po21  = ~n52043 & ~n52044;
  assign n52046 = ~n52037 & ~n52041;
  assign n52047 = n90 & n46426;
  assign n52048 = n14236 & n46420;
  assign n52049 = n54667 & n44952;
  assign n52050 = n14210 & n46009;
  assign n52051 = ~n52049 & ~n52050;
  assign n52052 = ~n52048 & n52051;
  assign n52053 = ~n52047 & n52052;
  assign n52054 = pi23  & ~n52053;
  assign n52055 = pi23  & ~n52054;
  assign n52056 = pi23  & n52053;
  assign n52057 = ~n52053 & ~n52054;
  assign n52058 = ~pi23  & ~n52053;
  assign n52059 = ~n60225 & ~n60226;
  assign n52060 = n123 & ~n59280;
  assign n52061 = n128 & n44871;
  assign n52062 = n53444 & n44327;
  assign n52063 = n127 & n44775;
  assign n52064 = ~n52062 & ~n52063;
  assign n52065 = ~n52061 & n52064;
  assign n52066 = ~n52060 & n52065;
  assign n52067 = pi26  & ~n52066;
  assign n52068 = pi26  & ~n52067;
  assign n52069 = pi26  & n52066;
  assign n52070 = ~n52066 & ~n52067;
  assign n52071 = ~pi26  & ~n52066;
  assign n52072 = ~n60227 & ~n60228;
  assign n52073 = ~n51955 & n51970;
  assign n52074 = ~n51955 & ~n51971;
  assign n52075 = ~n51956 & ~n52073;
  assign n52076 = ~n52072 & ~n60229;
  assign n52077 = n52072 & n60229;
  assign n52078 = ~n60229 & ~n52076;
  assign n52079 = n52072 & ~n60229;
  assign n52080 = ~n52072 & ~n52076;
  assign n52081 = ~n52072 & n60229;
  assign n52082 = ~n60230 & ~n60231;
  assign n52083 = ~n52076 & ~n52077;
  assign n52084 = n11279 & n39943;
  assign n52085 = n12584 & n39937;
  assign n52086 = n54410 & n39440;
  assign n52087 = n11267 & n39543;
  assign n52088 = ~n52086 & ~n52087;
  assign n52089 = ~n52085 & n52088;
  assign n52090 = ~n52084 & n52089;
  assign n52091 = pi29  & ~n52090;
  assign n52092 = pi29  & ~n52091;
  assign n52093 = pi29  & n52090;
  assign n52094 = ~n52090 & ~n52091;
  assign n52095 = ~pi29  & ~n52090;
  assign n52096 = ~n60233 & ~n60234;
  assign n52097 = ~n51944 & ~n51952;
  assign n52098 = ~n321 & ~n646;
  assign n52099 = ~n416 & ~n646;
  assign n52100 = ~n321 & n52099;
  assign n52101 = ~n416 & n52098;
  assign n52102 = n4381 & n5341;
  assign n52103 = ~n321 & n5341;
  assign n52104 = n4381 & n52099;
  assign n52105 = n52103 & n52104;
  assign n52106 = n60235 & n52102;
  assign n52107 = n53943 & n59003;
  assign n52108 = n60236 & n52107;
  assign n52109 = n53899 & n54333;
  assign n52110 = n53899 & n56574;
  assign n52111 = n54333 & n52110;
  assign n52112 = n56574 & n52109;
  assign n52113 = n52108 & n60237;
  assign n52114 = n53824 & n52113;
  assign n52115 = n54546 & n54733;
  assign n52116 = n54333 & n52107;
  assign n52117 = n54733 & n52116;
  assign n52118 = n54546 & n52117;
  assign n52119 = n56574 & n52118;
  assign n52120 = n53899 & n52119;
  assign n52121 = n53824 & n52120;
  assign n52122 = n4381 & n52121;
  assign n52123 = ~n416 & n52122;
  assign n52124 = ~n1465 & n52123;
  assign n52125 = ~n321 & n52124;
  assign n52126 = ~n646 & n52125;
  assign n52127 = ~n346 & n52126;
  assign n52128 = n52114 & n52115;
  assign n52129 = n60205 & n60238;
  assign n52130 = ~n60205 & ~n60238;
  assign n52131 = ~n52129 & ~n52130;
  assign n52132 = ~pi17  & n52131;
  assign n52133 = pi17  & ~n52131;
  assign n52134 = ~n52132 & ~n52133;
  assign n52135 = n1576 & n43436;
  assign n52136 = n11215 & n39546;
  assign n52137 = n54403 & n39552;
  assign n52138 = n10564 & n39549;
  assign n52139 = ~n52137 & ~n52138;
  assign n52140 = ~n52136 & n52139;
  assign n52141 = ~n52135 & n52140;
  assign n52142 = n52134 & ~n52141;
  assign n52143 = ~n52134 & n52141;
  assign n52144 = n52134 & ~n52142;
  assign n52145 = n52134 & n52141;
  assign n52146 = ~n52141 & ~n52142;
  assign n52147 = ~n52134 & ~n52141;
  assign n52148 = ~n60239 & ~n60240;
  assign n52149 = ~n52142 & ~n52143;
  assign n52150 = ~n51933 & ~n60241;
  assign n52151 = n51933 & n60241;
  assign n52152 = ~n60241 & ~n52150;
  assign n52153 = n51933 & ~n60241;
  assign n52154 = ~n51933 & ~n52150;
  assign n52155 = ~n51933 & n60241;
  assign n52156 = ~n60242 & ~n60243;
  assign n52157 = ~n52150 & ~n52151;
  assign n52158 = ~n52097 & ~n60244;
  assign n52159 = n52097 & n60244;
  assign n52160 = ~n52097 & ~n52158;
  assign n52161 = ~n60244 & ~n52158;
  assign n52162 = ~n52160 & ~n52161;
  assign n52163 = ~n52158 & ~n52159;
  assign n52164 = n52096 & n60245;
  assign n52165 = ~n52096 & ~n60245;
  assign n52166 = ~n60245 & ~n52165;
  assign n52167 = ~n52096 & ~n52165;
  assign n52168 = ~n52166 & ~n52167;
  assign n52169 = ~n52164 & ~n52165;
  assign n52170 = ~n60232 & ~n60246;
  assign n52171 = n60232 & n60246;
  assign n52172 = ~n60232 & n60246;
  assign n52173 = n60232 & ~n60246;
  assign n52174 = ~n52172 & ~n52173;
  assign n52175 = ~n52170 & ~n52171;
  assign n52176 = ~n52059 & ~n60247;
  assign n52177 = n52059 & n60247;
  assign n52178 = ~n52176 & ~n52177;
  assign n52179 = ~n51981 & n51995;
  assign n52180 = ~n51981 & ~n51997;
  assign n52181 = ~n51980 & ~n52179;
  assign n52182 = ~n52178 & n60248;
  assign n52183 = n52178 & ~n60248;
  assign n52184 = ~n52182 & ~n52183;
  assign n52185 = n14413 & ~n47526;
  assign n52186 = n54719 & n46788;
  assign n52187 = n15901 & n59503;
  assign n52188 = ~n52186 & ~n52187;
  assign n52189 = ~n52185 & n52188;
  assign n52190 = pi20  & ~n52189;
  assign n52191 = pi20  & ~n52190;
  assign n52192 = pi20  & n52189;
  assign n52193 = ~n52189 & ~n52190;
  assign n52194 = ~pi20  & ~n52189;
  assign n52195 = ~n60249 & ~n60250;
  assign n52196 = ~n52006 & n52020;
  assign n52197 = ~n52006 & ~n52021;
  assign n52198 = ~n52005 & ~n52196;
  assign n52199 = ~n52195 & ~n60251;
  assign n52200 = n52195 & n60251;
  assign n52201 = ~n60251 & ~n52199;
  assign n52202 = n52195 & ~n60251;
  assign n52203 = ~n52195 & ~n52199;
  assign n52204 = ~n52195 & n60251;
  assign n52205 = ~n60252 & ~n60253;
  assign n52206 = ~n52199 & ~n52200;
  assign n52207 = ~n52184 & n60254;
  assign n52208 = n52184 & ~n60254;
  assign n52209 = ~n52207 & ~n52208;
  assign n52210 = ~n51858 & n60222;
  assign n52211 = ~n51858 & ~n52027;
  assign n52212 = ~n51859 & ~n52210;
  assign n52213 = n52209 & ~n60255;
  assign n52214 = ~n52209 & n60255;
  assign n52215 = ~n52213 & ~n52214;
  assign n52216 = ~n52046 & n52215;
  assign n52217 = n52046 & ~n52215;
  assign n52218 = ~n52216 & ~n52217;
  assign n52219 = ~n52043 & ~n52218;
  assign n52220 = n52043 & n52218;
  assign po22  = ~n52219 & ~n52220;
  assign n52222 = ~n52213 & ~n52216;
  assign n52223 = ~n52199 & ~n52208;
  assign n52224 = ~n52176 & ~n52183;
  assign n52225 = n90 & n46805;
  assign n52226 = n14236 & n46788;
  assign n52227 = n54667 & n46009;
  assign n52228 = n14210 & n46420;
  assign n52229 = ~n52227 & ~n52228;
  assign n52230 = ~n52226 & n52229;
  assign n52231 = ~n52225 & n52230;
  assign n52232 = pi23  & ~n52231;
  assign n52233 = pi23  & ~n52232;
  assign n52234 = pi23  & n52231;
  assign n52235 = ~n52231 & ~n52232;
  assign n52236 = ~pi23  & ~n52231;
  assign n52237 = ~n60256 & ~n60257;
  assign n52238 = ~n52076 & ~n52170;
  assign n52239 = ~n52142 & ~n52150;
  assign n52240 = ~n52130 & ~n52132;
  assign n52241 = n1705 & n4530;
  assign n52242 = n13164 & n52241;
  assign n52243 = ~n630 & ~n659;
  assign n52244 = ~n163 & ~n1478;
  assign n52245 = n52243 & n52244;
  assign n52246 = n3742 & n4225;
  assign n52247 = ~n659 & ~n1478;
  assign n52248 = n4225 & n52247;
  assign n52249 = ~n163 & ~n630;
  assign n52250 = n3742 & n52249;
  assign n52251 = n52248 & n52250;
  assign n52252 = ~n659 & ~n1127;
  assign n52253 = n52244 & n52252;
  assign n52254 = ~n464 & ~n630;
  assign n52255 = n3742 & n52254;
  assign n52256 = n52253 & n52255;
  assign n52257 = n52245 & n52246;
  assign n52258 = n1940 & n54301;
  assign n52259 = n60258 & n52258;
  assign n52260 = n52242 & n52259;
  assign n52261 = n53748 & n54275;
  assign n52262 = n52260 & n52261;
  assign n52263 = n55100 & n52262;
  assign n52264 = n1705 & n1940;
  assign n52265 = n54301 & n52264;
  assign n52266 = n55100 & n52265;
  assign n52267 = n54275 & n52266;
  assign n52268 = n53748 & n52267;
  assign n52269 = n59903 & n52268;
  assign n52270 = n4530 & n52269;
  assign n52271 = n3742 & n52270;
  assign n52272 = n13164 & n52271;
  assign n52273 = ~n464 & n52272;
  assign n52274 = ~n1127 & n52273;
  assign n52275 = ~n1478 & n52274;
  assign n52276 = ~n163 & n52275;
  assign n52277 = ~n659 & n52276;
  assign n52278 = ~n630 & n52277;
  assign n52279 = n59903 & n52263;
  assign n52280 = ~n52240 & n60259;
  assign n52281 = n52240 & ~n60259;
  assign n52282 = ~n52280 & ~n52281;
  assign n52283 = n1576 & ~n59050;
  assign n52284 = n11215 & n39440;
  assign n52285 = n54403 & n39549;
  assign n52286 = n10564 & n39546;
  assign n52287 = ~n52285 & ~n52286;
  assign n52288 = ~n52284 & n52287;
  assign n52289 = ~n52283 & n52288;
  assign n52290 = n52282 & ~n52289;
  assign n52291 = ~n52282 & n52289;
  assign n52292 = ~n52289 & ~n52290;
  assign n52293 = n52282 & ~n52290;
  assign n52294 = ~n52292 & ~n52293;
  assign n52295 = ~n52290 & ~n52291;
  assign n52296 = n52239 & n60260;
  assign n52297 = ~n52239 & ~n60260;
  assign n52298 = ~n52296 & ~n52297;
  assign n52299 = n11279 & ~n59184;
  assign n52300 = n12584 & n44327;
  assign n52301 = n54410 & n39543;
  assign n52302 = n11267 & n39937;
  assign n52303 = ~n52301 & ~n52302;
  assign n52304 = ~n52300 & n52303;
  assign n52305 = ~n11279 & n52304;
  assign n52306 = n59184 & n52304;
  assign n52307 = ~n52305 & ~n52306;
  assign n52308 = ~n52299 & n52304;
  assign n52309 = pi29  & ~n60261;
  assign n52310 = ~pi29  & n60261;
  assign n52311 = ~n52309 & ~n52310;
  assign n52312 = n52298 & ~n52311;
  assign n52313 = ~n52298 & n52311;
  assign n52314 = ~n52312 & ~n52313;
  assign n52315 = n52096 & ~n52158;
  assign n52316 = ~n52158 & ~n52165;
  assign n52317 = ~n52159 & ~n52315;
  assign n52318 = n52314 & ~n60262;
  assign n52319 = ~n52314 & n60262;
  assign n52320 = ~n52318 & ~n52319;
  assign n52321 = n123 & ~n59275;
  assign n52322 = n128 & n44952;
  assign n52323 = n53444 & n44775;
  assign n52324 = n127 & n44871;
  assign n52325 = ~n52323 & ~n52324;
  assign n52326 = ~n52322 & n52325;
  assign n52327 = ~n52321 & n52326;
  assign n52328 = pi26  & ~n52327;
  assign n52329 = pi26  & ~n52328;
  assign n52330 = pi26  & n52327;
  assign n52331 = ~n52327 & ~n52328;
  assign n52332 = ~pi26  & ~n52327;
  assign n52333 = ~n60263 & ~n60264;
  assign n52334 = n52320 & ~n52333;
  assign n52335 = ~n52320 & n52333;
  assign n52336 = n52320 & ~n52334;
  assign n52337 = ~n52333 & ~n52334;
  assign n52338 = ~n52336 & ~n52337;
  assign n52339 = ~n52334 & ~n52335;
  assign n52340 = ~n52238 & ~n60265;
  assign n52341 = n52238 & n60265;
  assign n52342 = ~n60265 & ~n52340;
  assign n52343 = ~n52238 & ~n52340;
  assign n52344 = ~n52342 & ~n52343;
  assign n52345 = ~n52340 & ~n52341;
  assign n52346 = ~n52237 & ~n60266;
  assign n52347 = ~n60266 & ~n52346;
  assign n52348 = n52237 & ~n60266;
  assign n52349 = ~n52237 & ~n52346;
  assign n52350 = ~n52237 & n60266;
  assign n52351 = n52237 & n60266;
  assign n52352 = ~n52346 & ~n52351;
  assign n52353 = ~n60267 & ~n60268;
  assign n52354 = n52224 & ~n60269;
  assign n52355 = ~n52224 & n60269;
  assign n52356 = ~n52354 & ~n52355;
  assign n52357 = n54719 & n59503;
  assign n52358 = pi20  & n52357;
  assign n52359 = pi20  & ~n52358;
  assign n52360 = pi20  & ~n52357;
  assign n52361 = n52357 & ~n52358;
  assign n52362 = ~pi20  & n52357;
  assign n52363 = ~n60270 & ~n60271;
  assign n52364 = n52356 & ~n52363;
  assign n52365 = ~n52356 & n52363;
  assign n52366 = n52356 & ~n52364;
  assign n52367 = ~n52363 & ~n52364;
  assign n52368 = ~n52366 & ~n52367;
  assign n52369 = ~n52364 & ~n52365;
  assign n52370 = ~n52223 & ~n60272;
  assign n52371 = n52223 & n60272;
  assign n52372 = ~n60272 & ~n52370;
  assign n52373 = n52223 & ~n60272;
  assign n52374 = ~n52223 & ~n52370;
  assign n52375 = ~n52223 & n60272;
  assign n52376 = ~n60273 & ~n60274;
  assign n52377 = ~n52370 & ~n52371;
  assign n52378 = n52222 & n60275;
  assign n52379 = ~n52222 & ~n60275;
  assign n52380 = ~n52378 & ~n52379;
  assign n52381 = n52220 & n52380;
  assign n52382 = ~n52220 & ~n52380;
  assign po23  = ~n52381 & ~n52382;
  assign n52384 = n52237 & ~n52340;
  assign n52385 = ~n52340 & ~n52346;
  assign n52386 = ~n52341 & ~n52384;
  assign n52387 = pi20  & ~n60276;
  assign n52388 = ~pi20  & n60276;
  assign n52389 = ~n52387 & ~n52388;
  assign n52390 = n123 & ~n59386;
  assign n52391 = n128 & n46009;
  assign n52392 = n53444 & n44871;
  assign n52393 = n127 & n44952;
  assign n52394 = ~n52392 & ~n52393;
  assign n52395 = ~n52391 & n52394;
  assign n52396 = ~n52390 & n52395;
  assign n52397 = pi26  & ~n52396;
  assign n52398 = pi26  & ~n52397;
  assign n52399 = pi26  & n52396;
  assign n52400 = ~n52396 & ~n52397;
  assign n52401 = ~pi26  & ~n52396;
  assign n52402 = ~n60277 & ~n60278;
  assign n52403 = n4317 & n10238;
  assign n52404 = n27212 & n52403;
  assign n52405 = ~n174 & ~n1634;
  assign n52406 = n3780 & n52405;
  assign n52407 = n56585 & n52406;
  assign n52408 = n60202 & n52407;
  assign n52409 = n3780 & n52403;
  assign n52410 = n27212 & n52405;
  assign n52411 = n56585 & n52410;
  assign n52412 = n60202 & n52411;
  assign n52413 = n52409 & n52412;
  assign n52414 = n52404 & n52408;
  assign n52415 = n54544 & n59728;
  assign n52416 = n60279 & n52415;
  assign n52417 = n54646 & n55109;
  assign n52418 = n52416 & n52417;
  assign n52419 = n56585 & n60202;
  assign n52420 = n54646 & n52419;
  assign n52421 = n55109 & n52420;
  assign n52422 = n54544 & n52421;
  assign n52423 = n3780 & n52422;
  assign n52424 = n10238 & n52423;
  assign n52425 = n4317 & n52424;
  assign n52426 = n53832 & n52425;
  assign n52427 = n59728 & n52426;
  assign n52428 = ~n1490 & n52427;
  assign n52429 = ~n174 & n52428;
  assign n52430 = ~n1634 & n52429;
  assign n52431 = ~n770 & n52430;
  assign n52432 = n53832 & n52418;
  assign n52433 = ~n60259 & n60280;
  assign n52434 = n60259 & ~n60280;
  assign n52435 = ~n52433 & ~n52434;
  assign n52436 = n1576 & ~n59044;
  assign n52437 = n11215 & n39543;
  assign n52438 = n54403 & n39546;
  assign n52439 = n10564 & n39440;
  assign n52440 = ~n52438 & ~n52439;
  assign n52441 = ~n52437 & n52440;
  assign n52442 = ~n52436 & n52441;
  assign n52443 = ~n52434 & ~n52442;
  assign n52444 = ~n52433 & n52443;
  assign n52445 = n52435 & ~n52442;
  assign n52446 = ~n52435 & n52442;
  assign n52447 = ~n52442 & ~n60281;
  assign n52448 = ~n52434 & ~n60281;
  assign n52449 = ~n52433 & n52448;
  assign n52450 = ~n52447 & ~n52449;
  assign n52451 = ~n60281 & ~n52446;
  assign n52452 = ~n52280 & n52289;
  assign n52453 = ~n52280 & ~n52290;
  assign n52454 = ~n52281 & ~n52452;
  assign n52455 = n60282 & n60283;
  assign n52456 = ~n60282 & ~n60283;
  assign n52457 = ~n52455 & ~n52456;
  assign n52458 = ~n52297 & ~n52312;
  assign n52459 = ~n52457 & n52458;
  assign n52460 = n52457 & ~n52458;
  assign n52461 = ~n52459 & ~n52460;
  assign n52462 = n11279 & ~n59282;
  assign n52463 = n12584 & n44775;
  assign n52464 = n54410 & n39937;
  assign n52465 = n11267 & n44327;
  assign n52466 = ~n52464 & ~n52465;
  assign n52467 = ~n52463 & n52466;
  assign n52468 = ~n52462 & n52467;
  assign n52469 = pi29  & ~n52468;
  assign n52470 = pi29  & ~n52469;
  assign n52471 = pi29  & n52468;
  assign n52472 = ~n52468 & ~n52469;
  assign n52473 = ~pi29  & ~n52468;
  assign n52474 = ~n60284 & ~n60285;
  assign n52475 = n52461 & ~n52474;
  assign n52476 = ~n52461 & n52474;
  assign n52477 = n52461 & ~n52475;
  assign n52478 = n52461 & n52474;
  assign n52479 = ~n52474 & ~n52475;
  assign n52480 = ~n52461 & ~n52474;
  assign n52481 = ~n60286 & ~n60287;
  assign n52482 = ~n52475 & ~n52476;
  assign n52483 = ~n52402 & ~n60288;
  assign n52484 = n52402 & n60288;
  assign n52485 = ~n60288 & ~n52483;
  assign n52486 = ~n52402 & ~n52483;
  assign n52487 = ~n52485 & ~n52486;
  assign n52488 = ~n52483 & ~n52484;
  assign n52489 = ~n52318 & n52333;
  assign n52490 = ~n52318 & ~n52334;
  assign n52491 = ~n52319 & ~n52489;
  assign n52492 = n60289 & n60290;
  assign n52493 = ~n60289 & ~n60290;
  assign n52494 = ~n52492 & ~n52493;
  assign n52495 = n90 & ~n59554;
  assign n52496 = n14236 & n59503;
  assign n52497 = n54667 & n46420;
  assign n52498 = n14210 & n46788;
  assign n52499 = ~n52497 & ~n52498;
  assign n52500 = ~n52496 & n52499;
  assign n52501 = ~n52495 & n52500;
  assign n52502 = pi23  & ~n52501;
  assign n52503 = pi23  & ~n52502;
  assign n52504 = pi23  & n52501;
  assign n52505 = ~n52501 & ~n52502;
  assign n52506 = ~pi23  & ~n52501;
  assign n52507 = ~n60291 & ~n60292;
  assign n52508 = n52494 & ~n52507;
  assign n52509 = ~n52494 & n52507;
  assign n52510 = n52494 & ~n52508;
  assign n52511 = ~n52507 & ~n52508;
  assign n52512 = ~n52510 & ~n52511;
  assign n52513 = ~n52508 & ~n52509;
  assign n52514 = n52389 & ~n60293;
  assign n52515 = ~n52389 & n60293;
  assign n52516 = ~n60293 & ~n52514;
  assign n52517 = n52389 & ~n52514;
  assign n52518 = ~n52516 & ~n52517;
  assign n52519 = ~n52514 & ~n52515;
  assign n52520 = ~n52355 & n52363;
  assign n52521 = ~n52355 & ~n52364;
  assign n52522 = ~n52354 & ~n52520;
  assign n52523 = n60294 & n60295;
  assign n52524 = ~n60294 & ~n60295;
  assign n52525 = ~n52523 & ~n52524;
  assign n52526 = ~n52370 & ~n52379;
  assign n52527 = ~n52525 & n52526;
  assign n52528 = n52525 & ~n52526;
  assign n52529 = ~n52527 & ~n52528;
  assign n52530 = n52381 & n52529;
  assign n52531 = ~n52381 & ~n52529;
  assign po24  = ~n52530 & ~n52531;
  assign n52533 = ~n52524 & ~n52528;
  assign n52534 = ~n52475 & ~n52483;
  assign n52535 = n123 & n46426;
  assign n52536 = n128 & n46420;
  assign n52537 = n53444 & n44952;
  assign n52538 = n127 & n46009;
  assign n52539 = ~n52537 & ~n52538;
  assign n52540 = ~n52536 & n52539;
  assign n52541 = ~n52535 & n52540;
  assign n52542 = pi26  & ~n52541;
  assign n52543 = pi26  & ~n52542;
  assign n52544 = pi26  & n52541;
  assign n52545 = ~n52541 & ~n52542;
  assign n52546 = ~pi26  & ~n52541;
  assign n52547 = ~n60296 & ~n60297;
  assign n52548 = ~n52456 & ~n52460;
  assign n52549 = n1186 & n5116;
  assign n52550 = n5789 & n52549;
  assign n52551 = ~n316 & ~n1658;
  assign n52552 = ~n1476 & ~n1486;
  assign n52553 = ~n316 & ~n1476;
  assign n52554 = ~n1486 & ~n1658;
  assign n52555 = n52553 & n52554;
  assign n52556 = n52551 & n52552;
  assign n52557 = n3475 & n3675;
  assign n52558 = n60298 & n52557;
  assign n52559 = n1186 & n52557;
  assign n52560 = n5116 & n5789;
  assign n52561 = n60298 & n52560;
  assign n52562 = n52559 & n52561;
  assign n52563 = n3675 & n5116;
  assign n52564 = n3475 & n52563;
  assign n52565 = ~n419 & ~n1486;
  assign n52566 = n52551 & n52565;
  assign n52567 = ~n1455 & ~n1476;
  assign n52568 = n1186 & n52567;
  assign n52569 = n52566 & n52568;
  assign n52570 = n52564 & n52569;
  assign n52571 = n52550 & n52558;
  assign n52572 = n54259 & n56858;
  assign n52573 = n60299 & n52572;
  assign n52574 = n802 & n53706;
  assign n52575 = n53706 & n10078;
  assign n52576 = n802 & n52575;
  assign n52577 = n802 & n10078;
  assign n52578 = n53706 & n52577;
  assign n52579 = n10078 & n52574;
  assign n52580 = n57047 & n60300;
  assign n52581 = n52573 & n52580;
  assign n52582 = n53916 & n52581;
  assign n52583 = n1186 & n52575;
  assign n52584 = n56858 & n52583;
  assign n52585 = n57047 & n52584;
  assign n52586 = n54623 & n52585;
  assign n52587 = n53916 & n52586;
  assign n52588 = n5116 & n52587;
  assign n52589 = n802 & n52588;
  assign n52590 = n54259 & n52589;
  assign n52591 = n3675 & n52590;
  assign n52592 = n3475 & n52591;
  assign n52593 = ~n1486 & n52592;
  assign n52594 = ~n316 & n52593;
  assign n52595 = ~n1476 & n52594;
  assign n52596 = ~n1455 & n52595;
  assign n52597 = ~n1658 & n52596;
  assign n52598 = ~n419 & n52597;
  assign n52599 = n54623 & n52582;
  assign n52600 = n60259 & n60301;
  assign n52601 = ~n60259 & ~n60301;
  assign n52602 = ~n52600 & ~n52601;
  assign n52603 = ~pi20  & n52602;
  assign n52604 = pi20  & ~n52602;
  assign n52605 = ~n52603 & ~n52604;
  assign n52606 = ~n52448 & n52605;
  assign n52607 = n52448 & ~n52605;
  assign n52608 = ~n52606 & ~n52607;
  assign n52609 = n1576 & n39943;
  assign n52610 = n11215 & n39937;
  assign n52611 = n54403 & n39440;
  assign n52612 = n10564 & n39543;
  assign n52613 = ~n52611 & ~n52612;
  assign n52614 = ~n52610 & n52613;
  assign n52615 = ~n52609 & n52614;
  assign n52616 = n52608 & ~n52615;
  assign n52617 = ~n52608 & n52615;
  assign n52618 = n52608 & ~n52616;
  assign n52619 = ~n52615 & ~n52616;
  assign n52620 = ~n52618 & ~n52619;
  assign n52621 = ~n52616 & ~n52617;
  assign n52622 = n52548 & n60302;
  assign n52623 = ~n52548 & ~n60302;
  assign n52624 = ~n52622 & ~n52623;
  assign n52625 = n11279 & ~n59280;
  assign n52626 = n12584 & n44871;
  assign n52627 = n54410 & n44327;
  assign n52628 = n11267 & n44775;
  assign n52629 = ~n52627 & ~n52628;
  assign n52630 = ~n52626 & n52629;
  assign n52631 = ~n52625 & n52630;
  assign n52632 = pi29  & ~n52631;
  assign n52633 = pi29  & ~n52632;
  assign n52634 = pi29  & n52631;
  assign n52635 = ~n52631 & ~n52632;
  assign n52636 = ~pi29  & ~n52631;
  assign n52637 = ~n60303 & ~n60304;
  assign n52638 = ~n52624 & n52637;
  assign n52639 = n52624 & ~n52637;
  assign n52640 = n52624 & ~n52639;
  assign n52641 = ~n52637 & ~n52639;
  assign n52642 = ~n52640 & ~n52641;
  assign n52643 = ~n52638 & ~n52639;
  assign n52644 = ~n52547 & ~n60305;
  assign n52645 = n52547 & n60305;
  assign n52646 = ~n60305 & ~n52644;
  assign n52647 = n52547 & ~n60305;
  assign n52648 = ~n52547 & ~n52644;
  assign n52649 = ~n52547 & n60305;
  assign n52650 = ~n60306 & ~n60307;
  assign n52651 = ~n52644 & ~n52645;
  assign n52652 = n52534 & n60308;
  assign n52653 = ~n52534 & ~n60308;
  assign n52654 = ~n52652 & ~n52653;
  assign n52655 = n90 & ~n47526;
  assign n52656 = n54667 & n46788;
  assign n52657 = n14210 & n59503;
  assign n52658 = ~n52656 & ~n52657;
  assign n52659 = ~n52655 & n52658;
  assign n52660 = pi23  & ~n52659;
  assign n52661 = pi23  & ~n52660;
  assign n52662 = pi23  & n52659;
  assign n52663 = ~n52659 & ~n52660;
  assign n52664 = ~pi23  & ~n52659;
  assign n52665 = ~n60309 & ~n60310;
  assign n52666 = ~n52493 & n52507;
  assign n52667 = ~n52493 & ~n52508;
  assign n52668 = ~n52492 & ~n52666;
  assign n52669 = ~n52665 & ~n60311;
  assign n52670 = n52665 & n60311;
  assign n52671 = ~n60311 & ~n52669;
  assign n52672 = n52665 & ~n60311;
  assign n52673 = ~n52665 & ~n52669;
  assign n52674 = ~n52665 & n60311;
  assign n52675 = ~n60312 & ~n60313;
  assign n52676 = ~n52669 & ~n52670;
  assign n52677 = ~n52654 & n60314;
  assign n52678 = n52654 & ~n60314;
  assign n52679 = ~n52677 & ~n52678;
  assign n52680 = ~n52387 & n60293;
  assign n52681 = ~n52387 & ~n52514;
  assign n52682 = ~n52388 & ~n52680;
  assign n52683 = n52679 & ~n60315;
  assign n52684 = ~n52679 & n60315;
  assign n52685 = ~n52683 & ~n52684;
  assign n52686 = ~n52533 & n52685;
  assign n52687 = n52533 & ~n52685;
  assign n52688 = ~n52686 & ~n52687;
  assign n52689 = ~n52530 & ~n52688;
  assign n52690 = n52530 & n52688;
  assign po25  = ~n52689 & ~n52690;
  assign n52692 = ~n52683 & ~n52686;
  assign n52693 = ~n52669 & ~n52678;
  assign n52694 = ~n52644 & ~n52653;
  assign n52695 = ~n52601 & ~n52603;
  assign n52696 = ~n415 & ~n441;
  assign n52697 = ~n441 & ~n2109;
  assign n52698 = ~n415 & n52697;
  assign n52699 = ~n2109 & n52696;
  assign n52700 = n905 & n7004;
  assign n52701 = n60316 & n52700;
  assign n52702 = n1675 & n52701;
  assign n52703 = n1532 & n14520;
  assign n52704 = n15313 & n52703;
  assign n52705 = n54069 & n52704;
  assign n52706 = ~n441 & ~n1490;
  assign n52707 = ~n2109 & n52706;
  assign n52708 = ~n415 & ~n824;
  assign n52709 = n905 & n52708;
  assign n52710 = n52707 & n52709;
  assign n52711 = n1675 & n52710;
  assign n52712 = n1532 & n7004;
  assign n52713 = n7004 & n52703;
  assign n52714 = n14520 & n52712;
  assign n52715 = n54069 & n60317;
  assign n52716 = n52711 & n52715;
  assign n52717 = n52702 & n52705;
  assign n52718 = n54475 & n57062;
  assign n52719 = n60318 & n52718;
  assign n52720 = n54075 & n56746;
  assign n52721 = n52719 & n52720;
  assign n52722 = n56746 & n52715;
  assign n52723 = n1675 & n52722;
  assign n52724 = n54546 & n52723;
  assign n52725 = n54075 & n52724;
  assign n52726 = n54475 & n52725;
  assign n52727 = n57062 & n52726;
  assign n52728 = n905 & n52727;
  assign n52729 = ~n415 & n52728;
  assign n52730 = ~n1490 & n52729;
  assign n52731 = ~n824 & n52730;
  assign n52732 = ~n441 & n52731;
  assign n52733 = ~n2109 & n52732;
  assign n52734 = n54546 & n52721;
  assign n52735 = ~n52695 & n60319;
  assign n52736 = n52695 & ~n60319;
  assign n52737 = ~n52735 & ~n52736;
  assign n52738 = n1576 & ~n59184;
  assign n52739 = n11215 & n44327;
  assign n52740 = n54403 & n39543;
  assign n52741 = n10564 & n39937;
  assign n52742 = ~n52740 & ~n52741;
  assign n52743 = ~n52739 & n52742;
  assign n52744 = ~n52738 & n52743;
  assign n52745 = n52737 & ~n52744;
  assign n52746 = ~n52737 & n52744;
  assign n52747 = ~n52744 & ~n52745;
  assign n52748 = n52737 & ~n52745;
  assign n52749 = ~n52747 & ~n52748;
  assign n52750 = ~n52745 & ~n52746;
  assign n52751 = ~n52606 & n52615;
  assign n52752 = ~n52606 & ~n52616;
  assign n52753 = ~n52607 & ~n52751;
  assign n52754 = n60320 & n60321;
  assign n52755 = ~n60320 & ~n60321;
  assign n52756 = ~n52754 & ~n52755;
  assign n52757 = n11279 & ~n59275;
  assign n52758 = n12584 & n44952;
  assign n52759 = n54410 & n44775;
  assign n52760 = n11267 & n44871;
  assign n52761 = ~n52759 & ~n52760;
  assign n52762 = ~n52758 & n52761;
  assign n52763 = ~n11279 & n52762;
  assign n52764 = n59275 & n52762;
  assign n52765 = ~n52763 & ~n52764;
  assign n52766 = ~n52757 & n52762;
  assign n52767 = pi29  & ~n60322;
  assign n52768 = ~pi29  & n60322;
  assign n52769 = ~n52767 & ~n52768;
  assign n52770 = n52756 & ~n52769;
  assign n52771 = ~n52756 & n52769;
  assign n52772 = ~n52770 & ~n52771;
  assign n52773 = ~n52623 & n52637;
  assign n52774 = ~n52623 & ~n52639;
  assign n52775 = ~n52622 & ~n52773;
  assign n52776 = n52772 & ~n60323;
  assign n52777 = ~n52772 & n60323;
  assign n52778 = ~n52776 & ~n52777;
  assign n52779 = n123 & n46805;
  assign n52780 = n128 & n46788;
  assign n52781 = n53444 & n46009;
  assign n52782 = n127 & n46420;
  assign n52783 = ~n52781 & ~n52782;
  assign n52784 = ~n52780 & n52783;
  assign n52785 = ~n52779 & n52784;
  assign n52786 = pi26  & ~n52785;
  assign n52787 = pi26  & ~n52786;
  assign n52788 = pi26  & n52785;
  assign n52789 = ~n52785 & ~n52786;
  assign n52790 = ~pi26  & ~n52785;
  assign n52791 = ~n60324 & ~n60325;
  assign n52792 = n52778 & ~n52791;
  assign n52793 = ~n52778 & n52791;
  assign n52794 = n52778 & ~n52792;
  assign n52795 = ~n52791 & ~n52792;
  assign n52796 = ~n52794 & ~n52795;
  assign n52797 = ~n52792 & ~n52793;
  assign n52798 = n52694 & n60326;
  assign n52799 = ~n52694 & ~n60326;
  assign n52800 = ~n52798 & ~n52799;
  assign n52801 = n54667 & n59503;
  assign n52802 = pi23  & n52801;
  assign n52803 = pi23  & ~n52802;
  assign n52804 = pi23  & ~n52801;
  assign n52805 = n52801 & ~n52802;
  assign n52806 = ~pi23  & n52801;
  assign n52807 = ~n60327 & ~n60328;
  assign n52808 = ~n52800 & n52807;
  assign n52809 = n52800 & ~n52807;
  assign n52810 = n52800 & ~n52809;
  assign n52811 = ~n52807 & ~n52809;
  assign n52812 = ~n52810 & ~n52811;
  assign n52813 = ~n52808 & ~n52809;
  assign n52814 = ~n52693 & ~n60329;
  assign n52815 = n52693 & n60329;
  assign n52816 = ~n60329 & ~n52814;
  assign n52817 = n52693 & ~n60329;
  assign n52818 = ~n52693 & ~n52814;
  assign n52819 = ~n52693 & n60329;
  assign n52820 = ~n60330 & ~n60331;
  assign n52821 = ~n52814 & ~n52815;
  assign n52822 = n52692 & n60332;
  assign n52823 = ~n52692 & ~n60332;
  assign n52824 = ~n52822 & ~n52823;
  assign n52825 = n52690 & n52824;
  assign n52826 = ~n52690 & ~n52824;
  assign po26  = ~n52825 & ~n52826;
  assign n52828 = ~n52776 & n52791;
  assign n52829 = ~n52776 & ~n52792;
  assign n52830 = ~n52777 & ~n52828;
  assign n52831 = pi23  & ~n60333;
  assign n52832 = ~pi23  & n60333;
  assign n52833 = ~n52831 & ~n52832;
  assign n52834 = n123 & ~n59554;
  assign n52835 = n128 & n59503;
  assign n52836 = n53444 & n46420;
  assign n52837 = n127 & n46788;
  assign n52838 = ~n52836 & ~n52837;
  assign n52839 = ~n52835 & n52838;
  assign n52840 = ~n52834 & n52839;
  assign n52841 = pi26  & ~n52840;
  assign n52842 = pi26  & ~n52841;
  assign n52843 = pi26  & n52840;
  assign n52844 = ~n52840 & ~n52841;
  assign n52845 = ~pi26  & ~n52840;
  assign n52846 = ~n60334 & ~n60335;
  assign n52847 = ~n52755 & ~n52770;
  assign n52848 = n3780 & n4378;
  assign n52849 = n905 & n5955;
  assign n52850 = n52848 & n52849;
  assign n52851 = ~n144 & ~n179;
  assign n52852 = ~n401 & ~n823;
  assign n52853 = ~n144 & ~n823;
  assign n52854 = ~n179 & ~n401;
  assign n52855 = n52853 & n52854;
  assign n52856 = ~n144 & ~n401;
  assign n52857 = ~n179 & ~n823;
  assign n52858 = n52856 & n52857;
  assign n52859 = n52851 & n52852;
  assign n52860 = n749 & n3801;
  assign n52861 = n60336 & n52860;
  assign n52862 = n53596 & n57031;
  assign n52863 = n52861 & n52862;
  assign n52864 = n52849 & n52860;
  assign n52865 = n52848 & n60336;
  assign n52866 = n52862 & n52865;
  assign n52867 = n52864 & n52866;
  assign n52868 = n749 & n5955;
  assign n52869 = n3780 & n3801;
  assign n52870 = n52868 & n52869;
  assign n52871 = n905 & n4378;
  assign n52872 = n60336 & n52871;
  assign n52873 = n52862 & n52872;
  assign n52874 = n52870 & n52873;
  assign n52875 = n52850 & n52863;
  assign n52876 = n59241 & n59905;
  assign n52877 = n60337 & n52876;
  assign n52878 = n58736 & n52877;
  assign n52879 = n53596 & n3801;
  assign n52880 = n5955 & n52879;
  assign n52881 = n57031 & n52880;
  assign n52882 = n59241 & n52881;
  assign n52883 = n54359 & n52882;
  assign n52884 = n3780 & n52883;
  assign n52885 = n59905 & n52884;
  assign n52886 = n4378 & n52885;
  assign n52887 = n905 & n52886;
  assign n52888 = n749 & n52887;
  assign n52889 = n58736 & n52888;
  assign n52890 = ~n179 & n52889;
  assign n52891 = ~n144 & n52890;
  assign n52892 = ~n401 & n52891;
  assign n52893 = ~n823 & n52892;
  assign n52894 = n54359 & n52878;
  assign n52895 = n60319 & ~n60338;
  assign n52896 = ~n60319 & n60338;
  assign n52897 = ~n52895 & ~n52896;
  assign n52898 = ~n52735 & n52744;
  assign n52899 = ~n52735 & ~n52745;
  assign n52900 = ~n52736 & ~n52898;
  assign n52901 = ~n52896 & ~n60339;
  assign n52902 = ~n52895 & n52901;
  assign n52903 = n52897 & ~n60339;
  assign n52904 = ~n52897 & n60339;
  assign n52905 = ~n60339 & ~n60340;
  assign n52906 = ~n52896 & ~n60340;
  assign n52907 = ~n52895 & n52906;
  assign n52908 = ~n52905 & ~n52907;
  assign n52909 = ~n60340 & ~n52904;
  assign n52910 = n1576 & ~n59282;
  assign n52911 = n11215 & n44775;
  assign n52912 = n54403 & n39937;
  assign n52913 = n10564 & n44327;
  assign n52914 = ~n52912 & ~n52913;
  assign n52915 = ~n52911 & n52914;
  assign n52916 = ~n52910 & n52915;
  assign n52917 = ~n60341 & ~n52916;
  assign n52918 = n60341 & n52916;
  assign n52919 = ~n60341 & ~n52917;
  assign n52920 = ~n60341 & n52916;
  assign n52921 = ~n52916 & ~n52917;
  assign n52922 = n60341 & ~n52916;
  assign n52923 = ~n60342 & ~n60343;
  assign n52924 = ~n52917 & ~n52918;
  assign n52925 = n52847 & n60344;
  assign n52926 = ~n52847 & ~n60344;
  assign n52927 = ~n52925 & ~n52926;
  assign n52928 = n11279 & ~n59386;
  assign n52929 = n12584 & n46009;
  assign n52930 = n54410 & n44871;
  assign n52931 = n11267 & n44952;
  assign n52932 = ~n52930 & ~n52931;
  assign n52933 = ~n52929 & n52932;
  assign n52934 = ~n52928 & n52933;
  assign n52935 = pi29  & ~n52934;
  assign n52936 = pi29  & ~n52935;
  assign n52937 = pi29  & n52934;
  assign n52938 = ~n52934 & ~n52935;
  assign n52939 = ~pi29  & ~n52934;
  assign n52940 = ~n60345 & ~n60346;
  assign n52941 = n52927 & ~n52940;
  assign n52942 = ~n52927 & n52940;
  assign n52943 = n52927 & ~n52941;
  assign n52944 = n52927 & n52940;
  assign n52945 = ~n52940 & ~n52941;
  assign n52946 = ~n52927 & ~n52940;
  assign n52947 = ~n60347 & ~n60348;
  assign n52948 = ~n52941 & ~n52942;
  assign n52949 = ~n52846 & ~n60349;
  assign n52950 = n52846 & n60349;
  assign n52951 = ~n60349 & ~n52949;
  assign n52952 = n52846 & ~n60349;
  assign n52953 = ~n52846 & ~n52949;
  assign n52954 = ~n52846 & n60349;
  assign n52955 = ~n60350 & ~n60351;
  assign n52956 = ~n52949 & ~n52950;
  assign n52957 = n52833 & ~n60352;
  assign n52958 = ~n52833 & n60352;
  assign n52959 = ~n60352 & ~n52957;
  assign n52960 = n52833 & ~n52957;
  assign n52961 = ~n52959 & ~n52960;
  assign n52962 = ~n52957 & ~n52958;
  assign n52963 = ~n52799 & n52807;
  assign n52964 = ~n52799 & ~n52809;
  assign n52965 = ~n52798 & ~n52963;
  assign n52966 = n60353 & n60354;
  assign n52967 = ~n60353 & ~n60354;
  assign n52968 = ~n52966 & ~n52967;
  assign n52969 = ~n52814 & ~n52823;
  assign n52970 = ~n52968 & n52969;
  assign n52971 = n52968 & ~n52969;
  assign n52972 = ~n52970 & ~n52971;
  assign n52973 = n52825 & n52972;
  assign n52974 = ~n52825 & ~n52972;
  assign po27  = ~n52973 & ~n52974;
  assign n52976 = ~n52967 & ~n52971;
  assign n52977 = ~n52941 & ~n52949;
  assign n52978 = n123 & ~n47526;
  assign n52979 = n53444 & n46788;
  assign n52980 = n127 & n59503;
  assign n52981 = ~n52979 & ~n52980;
  assign n52982 = ~n52978 & n52981;
  assign n52983 = pi26  & ~n52982;
  assign n52984 = pi26  & ~n52983;
  assign n52985 = pi26  & n52982;
  assign n52986 = ~n52982 & ~n52983;
  assign n52987 = ~pi26  & ~n52982;
  assign n52988 = ~n60355 & ~n60356;
  assign n52989 = ~n52977 & ~n52988;
  assign n52990 = n52977 & n52988;
  assign n52991 = ~n52977 & ~n52989;
  assign n52992 = ~n52977 & n52988;
  assign n52993 = ~n52988 & ~n52989;
  assign n52994 = n52977 & ~n52988;
  assign n52995 = ~n60357 & ~n60358;
  assign n52996 = ~n52989 & ~n52990;
  assign n52997 = ~n52917 & ~n52926;
  assign n52998 = n452 & n2401;
  assign n52999 = n53474 & n52998;
  assign n53000 = n30483 & n52999;
  assign n53001 = n4002 & n7092;
  assign n53002 = n14916 & n53001;
  assign n53003 = n54734 & n53002;
  assign n53004 = n452 & n7092;
  assign n53005 = n53474 & n53004;
  assign n53006 = n30483 & n53005;
  assign n53007 = n2401 & n4002;
  assign n53008 = n14916 & n53007;
  assign n53009 = n54734 & n53008;
  assign n53010 = n53006 & n53009;
  assign n53011 = ~n422 & ~n560;
  assign n53012 = ~n628 & ~n1059;
  assign n53013 = n53011 & n53012;
  assign n53014 = n53474 & n53013;
  assign n53015 = n30483 & n53014;
  assign n53016 = n452 & n4002;
  assign n53017 = n14916 & n53016;
  assign n53018 = n54734 & n53017;
  assign n53019 = n53015 & n53018;
  assign n53020 = ~n584 & ~n1059;
  assign n53021 = ~n342 & ~n628;
  assign n53022 = n53020 & n53021;
  assign n53023 = n1642 & n53011;
  assign n53024 = n53022 & n53023;
  assign n53025 = n53474 & n53024;
  assign n53026 = n1035 & n4002;
  assign n53027 = n452 & n53026;
  assign n53028 = n54734 & n53027;
  assign n53029 = n53025 & n53028;
  assign n53030 = n53000 & n53003;
  assign n53031 = n53457 & n60360;
  assign n53032 = n53627 & n60360;
  assign n53033 = n53457 & n53032;
  assign n53034 = n53627 & n53031;
  assign n53035 = n53549 & n54734;
  assign n53036 = n452 & n53035;
  assign n53037 = n53457 & n53036;
  assign n53038 = n53627 & n53037;
  assign n53039 = n4002 & n53038;
  assign n53040 = n1035 & n53039;
  assign n53041 = n53474 & n53040;
  assign n53042 = n1642 & n53041;
  assign n53043 = ~n422 & n53042;
  assign n53044 = ~n628 & n53043;
  assign n53045 = ~n560 & n53044;
  assign n53046 = ~n584 & n53045;
  assign n53047 = ~n1059 & n53046;
  assign n53048 = ~n342 & n53047;
  assign n53049 = n53549 & n60361;
  assign n53050 = n60338 & n60362;
  assign n53051 = ~n60338 & ~n60362;
  assign n53052 = ~n53050 & ~n53051;
  assign n53053 = ~pi23  & n53052;
  assign n53054 = pi23  & ~n53052;
  assign n53055 = ~n53053 & ~n53054;
  assign n53056 = ~n52906 & n53055;
  assign n53057 = n52906 & ~n53055;
  assign n53058 = ~n53056 & ~n53057;
  assign n53059 = n1576 & ~n59280;
  assign n53060 = n11215 & n44871;
  assign n53061 = n54403 & n44327;
  assign n53062 = n10564 & n44775;
  assign n53063 = ~n53061 & ~n53062;
  assign n53064 = ~n53060 & n53063;
  assign n53065 = ~n53059 & n53064;
  assign n53066 = n53058 & ~n53065;
  assign n53067 = ~n53058 & n53065;
  assign n53068 = n53058 & ~n53066;
  assign n53069 = ~n53065 & ~n53066;
  assign n53070 = ~n53068 & ~n53069;
  assign n53071 = ~n53066 & ~n53067;
  assign n53072 = n52997 & n60363;
  assign n53073 = ~n52997 & ~n60363;
  assign n53074 = ~n53072 & ~n53073;
  assign n53075 = n11279 & n46426;
  assign n53076 = n12584 & n46420;
  assign n53077 = n54410 & n44952;
  assign n53078 = n11267 & n46009;
  assign n53079 = ~n53077 & ~n53078;
  assign n53080 = ~n53076 & n53079;
  assign n53081 = ~n53075 & n53080;
  assign n53082 = pi29  & ~n53081;
  assign n53083 = pi29  & ~n53082;
  assign n53084 = pi29  & n53081;
  assign n53085 = ~n53081 & ~n53082;
  assign n53086 = ~pi29  & ~n53081;
  assign n53087 = ~n60364 & ~n60365;
  assign n53088 = ~n53074 & n53087;
  assign n53089 = n53074 & ~n53087;
  assign n53090 = n53074 & ~n53089;
  assign n53091 = ~n53087 & ~n53089;
  assign n53092 = ~n53090 & ~n53091;
  assign n53093 = ~n53088 & ~n53089;
  assign n53094 = ~n60359 & ~n60366;
  assign n53095 = n60359 & n60366;
  assign n53096 = ~n60359 & n60366;
  assign n53097 = n60359 & ~n60366;
  assign n53098 = ~n53096 & ~n53097;
  assign n53099 = ~n53094 & ~n53095;
  assign n53100 = ~n52831 & n60352;
  assign n53101 = ~n52831 & ~n52957;
  assign n53102 = ~n52832 & ~n53100;
  assign n53103 = ~n60367 & ~n60368;
  assign n53104 = n60367 & n60368;
  assign n53105 = ~n53103 & ~n53104;
  assign n53106 = ~n52976 & n53105;
  assign n53107 = n52976 & ~n53105;
  assign n53108 = ~n53106 & ~n53107;
  assign n53109 = ~n52973 & ~n53108;
  assign n53110 = n52973 & n53108;
  assign po28  = ~n53109 & ~n53110;
  assign n53112 = ~n53103 & ~n53106;
  assign n53113 = ~n52989 & ~n53094;
  assign n53114 = ~n53051 & ~n53053;
  assign n53115 = n755 & n3083;
  assign n53116 = n1067 & n4214;
  assign n53117 = n53115 & n53116;
  assign n53118 = ~n316 & ~n441;
  assign n53119 = n322 & n53118;
  assign n53120 = n56849 & n53119;
  assign n53121 = n53117 & n53120;
  assign n53122 = n906 & n7350;
  assign n53123 = n12490 & n53122;
  assign n53124 = n55117 & n53123;
  assign n53125 = n906 & n4214;
  assign n53126 = n322 & n3083;
  assign n53127 = n53125 & n53126;
  assign n53128 = n755 & n53118;
  assign n53129 = n56849 & n53128;
  assign n53130 = n53127 & n53129;
  assign n53131 = n1067 & n7350;
  assign n53132 = n12490 & n53131;
  assign n53133 = n55117 & n53132;
  assign n53134 = n53130 & n53133;
  assign n53135 = n1067 & n3083;
  assign n53136 = n53125 & n53135;
  assign n53137 = n12490 & n53118;
  assign n53138 = n56849 & n53137;
  assign n53139 = n53136 & n53138;
  assign n53140 = n755 & n7350;
  assign n53141 = n322 & n53140;
  assign n53142 = n55117 & n53141;
  assign n53143 = n53139 & n53142;
  assign n53144 = n53121 & n53124;
  assign n53145 = n53453 & n53652;
  assign n53146 = n53453 & n60369;
  assign n53147 = n53652 & n53146;
  assign n53148 = n60369 & n53145;
  assign n53149 = n57025 & n60370;
  assign n53150 = n7350 & n56849;
  assign n53151 = n3083 & n53150;
  assign n53152 = n55117 & n53151;
  assign n53153 = n59269 & n53152;
  assign n53154 = n57025 & n53153;
  assign n53155 = n53652 & n53154;
  assign n53156 = n53453 & n53155;
  assign n53157 = n1067 & n53156;
  assign n53158 = n755 & n53157;
  assign n53159 = n906 & n53158;
  assign n53160 = n322 & n53159;
  assign n53161 = n4214 & n53160;
  assign n53162 = ~n316 & n53161;
  assign n53163 = ~n832 & n53162;
  assign n53164 = ~n441 & n53163;
  assign n53165 = ~n747 & n53164;
  assign n53166 = n59269 & n53149;
  assign n53167 = ~n53114 & n60371;
  assign n53168 = n53114 & ~n60371;
  assign n53169 = ~n53167 & ~n53168;
  assign n53170 = n1576 & ~n59275;
  assign n53171 = n11215 & n44952;
  assign n53172 = n54403 & n44775;
  assign n53173 = n10564 & n44871;
  assign n53174 = ~n53172 & ~n53173;
  assign n53175 = ~n53171 & n53174;
  assign n53176 = ~n53170 & n53175;
  assign n53177 = n53169 & ~n53176;
  assign n53178 = ~n53169 & n53176;
  assign n53179 = ~n53176 & ~n53177;
  assign n53180 = n53169 & ~n53177;
  assign n53181 = ~n53179 & ~n53180;
  assign n53182 = ~n53177 & ~n53178;
  assign n53183 = ~n53056 & n53065;
  assign n53184 = ~n53056 & ~n53066;
  assign n53185 = ~n53057 & ~n53183;
  assign n53186 = n60372 & n60373;
  assign n53187 = ~n60372 & ~n60373;
  assign n53188 = ~n53186 & ~n53187;
  assign n53189 = n11279 & n46805;
  assign n53190 = n12584 & n46788;
  assign n53191 = n54410 & n46009;
  assign n53192 = n11267 & n46420;
  assign n53193 = ~n53191 & ~n53192;
  assign n53194 = ~n53190 & n53193;
  assign n53195 = ~n11279 & n53194;
  assign n53196 = ~n46805 & n53194;
  assign n53197 = ~n53195 & ~n53196;
  assign n53198 = ~n53189 & n53194;
  assign n53199 = pi29  & ~n60374;
  assign n53200 = ~pi29  & n60374;
  assign n53201 = ~n53199 & ~n53200;
  assign n53202 = n53188 & ~n53201;
  assign n53203 = ~n53188 & n53201;
  assign n53204 = ~n53202 & ~n53203;
  assign n53205 = ~n53073 & n53087;
  assign n53206 = ~n53073 & ~n53089;
  assign n53207 = ~n53072 & ~n53205;
  assign n53208 = n53204 & ~n60375;
  assign n53209 = ~n53204 & n60375;
  assign n53210 = ~n53208 & ~n53209;
  assign n53211 = n53444 & n59503;
  assign n53212 = pi26  & n53211;
  assign n53213 = pi26  & ~n53212;
  assign n53214 = pi26  & ~n53211;
  assign n53215 = n53211 & ~n53212;
  assign n53216 = ~pi26  & n53211;
  assign n53217 = ~n60376 & ~n60377;
  assign n53218 = n53210 & ~n53217;
  assign n53219 = ~n53210 & n53217;
  assign n53220 = n53210 & ~n53218;
  assign n53221 = ~n53217 & ~n53218;
  assign n53222 = ~n53220 & ~n53221;
  assign n53223 = ~n53218 & ~n53219;
  assign n53224 = ~n53113 & ~n60378;
  assign n53225 = n53113 & n60378;
  assign n53226 = ~n60378 & ~n53224;
  assign n53227 = ~n53113 & ~n53224;
  assign n53228 = ~n53226 & ~n53227;
  assign n53229 = ~n53224 & ~n53225;
  assign n53230 = n53112 & n60379;
  assign n53231 = ~n53112 & ~n60379;
  assign n53232 = ~n53230 & ~n53231;
  assign n53233 = n53110 & n53232;
  assign n53234 = ~n53110 & ~n53232;
  assign po29  = ~n53233 & ~n53234;
  assign n53236 = ~n53224 & ~n53231;
  assign n53237 = ~n53187 & ~n53202;
  assign n53238 = n53464 & n26220;
  assign n53239 = n53464 & ~n584;
  assign n53240 = n53477 & n26220;
  assign n53241 = n53239 & n53240;
  assign n53242 = n596 & n53238;
  assign n53243 = n53451 & n53492;
  assign n53244 = n53492 & ~n53622;
  assign n53245 = n53451 & n53244;
  assign n53246 = ~n53622 & n53243;
  assign n53247 = n53451 & n26220;
  assign n53248 = n53464 & n53247;
  assign n53249 = n53451 & n53238;
  assign n53250 = n596 & n53492;
  assign n53251 = ~n53622 & n53250;
  assign n53252 = n60382 & n53251;
  assign n53253 = n53492 & n53238;
  assign n53254 = n53451 & n596;
  assign n53255 = ~n53622 & n53254;
  assign n53256 = n53253 & n53255;
  assign n53257 = n60380 & n60381;
  assign n53258 = ~n53622 & n60382;
  assign n53259 = n53492 & n53258;
  assign n53260 = n59269 & n53259;
  assign n53261 = n53477 & n53260;
  assign n53262 = ~n584 & n53261;
  assign n53263 = n59269 & n60383;
  assign n53264 = ~n60371 & n60384;
  assign n53265 = n60371 & ~n60384;
  assign n53266 = ~n53264 & ~n53265;
  assign n53267 = ~n53167 & n53176;
  assign n53268 = ~n53167 & ~n53177;
  assign n53269 = ~n53168 & ~n53267;
  assign n53270 = ~n53265 & ~n60385;
  assign n53271 = ~n53264 & n53270;
  assign n53272 = n53266 & ~n60385;
  assign n53273 = ~n53266 & n60385;
  assign n53274 = ~n60385 & ~n60386;
  assign n53275 = ~n53265 & ~n60386;
  assign n53276 = ~n53264 & n53275;
  assign n53277 = ~n53274 & ~n53276;
  assign n53278 = ~n60386 & ~n53273;
  assign n53279 = n1576 & ~n59386;
  assign n53280 = n11215 & n46009;
  assign n53281 = n54403 & n44871;
  assign n53282 = n10564 & n44952;
  assign n53283 = ~n53281 & ~n53282;
  assign n53284 = ~n53280 & n53283;
  assign n53285 = ~n53279 & n53284;
  assign n53286 = ~n60387 & ~n53285;
  assign n53287 = n60387 & n53285;
  assign n53288 = ~n60387 & ~n53286;
  assign n53289 = ~n60387 & n53285;
  assign n53290 = ~n53285 & ~n53286;
  assign n53291 = n60387 & ~n53285;
  assign n53292 = ~n60388 & ~n60389;
  assign n53293 = ~n53286 & ~n53287;
  assign n53294 = n53237 & n60390;
  assign n53295 = ~n53237 & ~n60390;
  assign n53296 = ~n53294 & ~n53295;
  assign n53297 = n11279 & ~n59554;
  assign n53298 = n12584 & n59503;
  assign n53299 = n54410 & n46420;
  assign n53300 = n11267 & n46788;
  assign n53301 = ~n53299 & ~n53300;
  assign n53302 = ~n53298 & n53301;
  assign n53303 = ~n53297 & n53302;
  assign n53304 = pi29  & ~n53303;
  assign n53305 = pi29  & ~n53304;
  assign n53306 = pi29  & n53303;
  assign n53307 = ~n53303 & ~n53304;
  assign n53308 = ~pi29  & ~n53303;
  assign n53309 = ~n60391 & ~n60392;
  assign n53310 = pi26  & ~n53309;
  assign n53311 = ~pi26  & n53309;
  assign n53312 = pi26  & ~n53310;
  assign n53313 = pi26  & n53309;
  assign n53314 = ~n53309 & ~n53310;
  assign n53315 = ~pi26  & ~n53309;
  assign n53316 = ~n60393 & ~n60394;
  assign n53317 = ~n53310 & ~n53311;
  assign n53318 = ~n53296 & n60395;
  assign n53319 = n53296 & ~n60395;
  assign n53320 = ~n53318 & ~n53319;
  assign n53321 = ~n53208 & n53217;
  assign n53322 = ~n53208 & ~n53218;
  assign n53323 = ~n53209 & ~n53321;
  assign n53324 = n53320 & ~n60396;
  assign n53325 = ~n53320 & n60396;
  assign n53326 = ~n53324 & ~n53325;
  assign n53327 = ~n53236 & n53326;
  assign n53328 = n53236 & ~n53326;
  assign n53329 = ~n53327 & ~n53328;
  assign n53330 = ~n53233 & ~n53329;
  assign n53331 = n53233 & n53329;
  assign po30  = ~n53330 & ~n53331;
  assign n53333 = ~n53324 & ~n53327;
  assign n53334 = ~n53310 & ~n53319;
  assign n53335 = ~n60371 & n53334;
  assign n53336 = n60371 & ~n53334;
  assign n53337 = ~n53335 & ~n53336;
  assign n53338 = n53333 & n53337;
  assign n53339 = ~n53333 & ~n53337;
  assign n53340 = n53333 & ~n53334;
  assign n53341 = ~n53333 & n53334;
  assign n53342 = ~n53340 & ~n53341;
  assign n53343 = n60371 & ~n53342;
  assign n53344 = ~n60371 & n53342;
  assign n53345 = ~n53343 & ~n53344;
  assign n53346 = n60371 & n53342;
  assign n53347 = ~n60371 & ~n53342;
  assign n53348 = ~n53346 & ~n53347;
  assign n53349 = ~n53338 & ~n53339;
  assign n53350 = n1576 & n46426;
  assign n53351 = n11215 & n46420;
  assign n53352 = n54403 & n44952;
  assign n53353 = n10564 & n46009;
  assign n53354 = ~n53352 & ~n53353;
  assign n53355 = ~n53351 & n53354;
  assign n53356 = ~n53350 & n53355;
  assign n53357 = n11279 & ~n47526;
  assign n53358 = n54410 & n46788;
  assign n53359 = ~n53357 & ~n53358;
  assign n53360 = n53275 & ~n53359;
  assign n53361 = ~n53275 & n53359;
  assign n53362 = ~n53360 & ~n53361;
  assign n53363 = ~n53286 & ~n53295;
  assign n53364 = n53563 & n2388;
  assign n53365 = ~n852 & n53364;
  assign n53366 = n1628 & n2388;
  assign n53367 = pi26  & ~n60398;
  assign n53368 = ~pi26  & n60398;
  assign n53369 = ~n53367 & ~n53368;
  assign n53370 = pi29  & ~n53369;
  assign n53371 = ~pi29  & n53369;
  assign n53372 = ~n53370 & ~n53371;
  assign n53373 = n53363 & n53372;
  assign n53374 = ~n53363 & ~n53372;
  assign n53375 = ~n53373 & ~n53374;
  assign n53376 = n53362 & ~n53375;
  assign n53377 = ~n53362 & n53375;
  assign n53378 = ~n53275 & n53363;
  assign n53379 = n53275 & ~n53363;
  assign n53380 = ~n53378 & ~n53379;
  assign n53381 = pi29  & ~n53380;
  assign n53382 = ~pi29  & n53380;
  assign n53383 = ~n53381 & ~n53382;
  assign n53384 = n53359 & n53383;
  assign n53385 = ~n53359 & ~n53383;
  assign n53386 = ~n53384 & ~n53385;
  assign n53387 = n53369 & ~n53386;
  assign n53388 = ~n53369 & n53386;
  assign n53389 = ~n53387 & ~n53388;
  assign n53390 = ~n53376 & ~n53377;
  assign n53391 = n53356 & ~n60399;
  assign n53392 = ~n53356 & n60399;
  assign n53393 = n53356 & n60399;
  assign n53394 = ~n53356 & ~n60399;
  assign n53395 = ~n53393 & ~n53394;
  assign n53396 = pi29  & ~n53359;
  assign n53397 = ~pi29  & n53359;
  assign n53398 = ~n53396 & ~n53397;
  assign n53399 = ~n53356 & n53398;
  assign n53400 = n53356 & ~n53398;
  assign n53401 = ~n53399 & ~n53400;
  assign n53402 = n53380 & n53401;
  assign n53403 = ~n53380 & ~n53401;
  assign n53404 = pi29  & ~n53363;
  assign n53405 = ~pi29  & n53363;
  assign n53406 = ~n53404 & ~n53405;
  assign n53407 = n53359 & n53406;
  assign n53408 = ~n53359 & ~n53406;
  assign n53409 = ~n53407 & ~n53408;
  assign n53410 = n53275 & ~n53356;
  assign n53411 = ~n53275 & n53356;
  assign n53412 = ~n53410 & ~n53411;
  assign n53413 = n53409 & ~n53412;
  assign n53414 = ~n53409 & n53412;
  assign n53415 = ~n53413 & ~n53414;
  assign n53416 = ~n53402 & ~n53403;
  assign n53417 = n53369 & ~n60401;
  assign n53418 = ~n53369 & n60401;
  assign n53419 = ~n53417 & ~n53418;
  assign n53420 = ~n53391 & ~n53392;
  assign n53421 = ~n53331 & ~n60400;
  assign n53422 = n53331 & n60400;
  assign n53423 = ~n53421 & ~n53422;
  assign n53424 = n60397 & n53423;
  assign n53425 = ~n60397 & ~n53423;
  assign n53426 = ~n53331 & n60397;
  assign n53427 = n53331 & ~n60397;
  assign n53428 = ~n53426 & ~n53427;
  assign n53429 = ~n60400 & n53428;
  assign n53430 = n60400 & ~n53428;
  assign n53431 = ~n53429 & ~n53430;
  assign n53432 = ~n60397 & n60400;
  assign n53433 = n60397 & ~n60400;
  assign n53434 = ~n53432 & ~n53433;
  assign n53435 = ~n53331 & n53434;
  assign n53436 = n53331 & ~n53434;
  assign n53437 = ~n53435 & ~n53436;
  assign n53438 = ~n53424 & ~n53425;
  assign n53439 = n69 | ~n70;
  assign n53440 = n75 | ~n76;
  assign n53441 = n82 | ~n83;
  assign n53442 = n88 | ~n89;
  assign n53443 = n95 | n96;
  assign n53444 = n125 | n126;
  assign n53445 = n134 | n131 | n133;
  assign n53446 = n138 | n136 | n137;
  assign n53447 = n148 | n149;
  assign n53448 = n159 | n153 | n158;
  assign n53449 = n191 | n192;
  assign n53450 = n198 | n193 | n197;
  assign n53451 = n204 | n205;
  assign n53452 = n226 | n227;
  assign n53453 = n234 | n238 | n244 | n245;
  assign n53454 = n253 | n254;
  assign n53455 = n264 | n265;
  assign n53456 = n279 | n280;
  assign n53457 = n287 | n288;
  assign n53458 = n299 | n300;
  assign n53459 = n306 | n303 | n305;
  assign n53460 = n314 | n315;
  assign n53461 = n325 | n326;
  assign n53462 = n328 | n329;
  assign n53463 = n337 | n338;
  assign n53464 = n391 | n376 | n384 | n398 | n399;
  assign n53465 = n430 | n431;
  assign n53466 = n433 | n434;
  assign n53467 = n436 | n437;
  assign n53468 = n456 | n457;
  assign n53469 = n469 | n470;
  assign n53470 = n490 | n481 | n489;
  assign n53471 = n526 | n534 | n545 | n546;
  assign n53472 = n543 | n544;
  assign n53473 = n550 | n551;
  assign n53474 = n557 | n558;
  assign n53475 = n572 | n573;
  assign n53476 = n575 | n576;
  assign n53477 = n582 | n583;
  assign n53478 = n597 | n598;
  assign n53479 = n602 | n606 | n609 | n610;
  assign n53480 = n637 | n638;
  assign n53481 = n641 | n642;
  assign n53482 = n644 | n645;
  assign n53483 = n658 | n655 | n657;
  assign n53484 = n677 | n670 | n674 | n679 | n680;
  assign n53485 = n691 | n692;
  assign n53486 = n695 | n696;
  assign n53487 = n706 | n707;
  assign n53488 = n710 | n711;
  assign n53489 = n715 | n716;
  assign n53490 = n721 | n722;
  assign n53491 = n724 | n725;
  assign n53492 = n731 | n732;
  assign n53493 = n738 | n739;
  assign n53494 = n745 | n746;
  assign n53495 = n758 | n759;
  assign n53496 = n769 | n764 | n768;
  assign n53497 = n781 | n782;
  assign n53498 = n786 | n787;
  assign n53499 = n796 | n797;
  assign n53500 = n813 | n808 | n812;
  assign n53501 = n816 | n817;
  assign n53502 = n821 | n818 | n820;
  assign n53503 = n827 | n828;
  assign n53504 = n845 | n840 | n844;
  assign n53505 = n856 | n857;
  assign n53506 = n859 | n860;
  assign n53507 = n863 | n864;
  assign n53508 = n873 | n874;
  assign n53509 = n889 | n886 | n888;
  assign n53510 = n892 | n893;
  assign n53511 = n920 | n921;
  assign n53512 = n925 | n926;
  assign n53513 = n947 | n939 | n946;
  assign n53514 = n954 | n951 | n953;
  assign n53515 = n961 | n962;
  assign n53516 = n973 | n974;
  assign n53517 = n980 | n981;
  assign n53518 = n993 | n990 | n992;
  assign n53519 = n1000 | n997 | n999;
  assign n53520 = n1016 | n1017;
  assign n53521 = n1023 | n1024;
  assign n53522 = n1029 | n1030;
  assign n53523 = n1041 | n1038 | n1040;
  assign n53524 = n1058 | n1050 | n1057;
  assign n53525 = n1055 | n1056;
  assign n53526 = n1071 | n1072;
  assign n53527 = n1098 | n1099;
  assign n53528 = n1105 | n1114 | n1118 | n1119;
  assign n53529 = n1110 | n1111;
  assign n53530 = n1134 | n1135;
  assign n53531 = n1153 | n1166 | n1182 | n1183;
  assign n53532 = n1203 | n1204;
  assign n53533 = n1211 | n1207 | n1210;
  assign n53534 = n1233 | n1224 | n1232;
  assign n53535 = n1237 | n1238;
  assign n53536 = n1241 | n1242;
  assign n53537 = n1263 | n1264;
  assign n53538 = n1320 | n1298 | n1308 | n1334 | n1335;
  assign n53539 = n1340 | n1341;
  assign n53540 = n1344 | n1345;
  assign n53541 = n1351 | n1352;
  assign n53542 = n1356 | n1357;
  assign n53543 = n1375 | n1380 | n1385 | n1386;
  assign n53544 = n1377 | n1378;
  assign n53545 = n1389 | n1390;
  assign n53546 = n1394 | n1395;
  assign n53547 = n1411 | n1423 | n1437 | n1438;
  assign n53548 = n1453 | n1454;
  assign n53549 = n1463 | n1464;
  assign n53550 = n1484 | n1481 | n1483;
  assign n53551 = n1495 | n1496;
  assign n53552 = n1506 | n1514 | n1527 | n1528;
  assign n53553 = n1518 | n1519;
  assign n53554 = n1521 | n1522;
  assign n53555 = n1525 | n1526;
  assign n53556 = n1543 | n1544;
  assign n53557 = n1546 | n1547;
  assign n53558 = n1554 | n1555;
  assign n53559 = n1565 | n1566;
  assign n53560 = n1571 | n1572;
  assign n53561 = n1581 | n1582;
  assign n53562 = n1597 | n1590 | n1596;
  assign n53563 = n1607 | n1608;
  assign n53564 = n1615 | n1619 | n1623 | n1624;
  assign n53565 = n1633 | n1629 | n1632;
  assign n53566 = n1640 | n1637 | n1639;
  assign n53567 = n1651 | n1652;
  assign n53568 = n1655 | n1656;
  assign n53569 = n1668 | ~n1669;
  assign n53570 = n1678 | n1679;
  assign n53571 = n1686 | n1687;
  assign n53572 = n1701 | n1694 | n1700;
  assign n53573 = n1719 | n1720;
  assign n53574 = n1723 | n1724;
  assign n53575 = n1732 | n1739 | n1744 | n1745;
  assign n53576 = n1756 | n1757;
  assign n53577 = n1768 | n1765 | n1767;
  assign n53578 = n1790 | n1780 | n1789;
  assign n53579 = n1800 | n1801;
  assign n53580 = n1815 | n1809 | n1814;
  assign n53581 = n1812 | n1813;
  assign n53582 = n1823 | n1824;
  assign n53583 = n1836 | n1829 | n1835;
  assign n53584 = n1844 | n1845;
  assign n53585 = n1848 | n1849;
  assign n53586 = n1857 | n1858;
  assign n53587 = n1864 | n1865;
  assign n53588 = n1872 | n1873;
  assign n53589 = n1880 | n1877 | n1879;
  assign n53590 = n1897 | n1892 | n1896;
  assign n53591 = n1910 | n1911;
  assign n53592 = n1918 | n1915 | n1917;
  assign n53593 = n1923 | n1924;
  assign n53594 = n1928 | n1929;
  assign n53595 = n1934 | n1935;
  assign n53596 = n1943 | n1944;
  assign n53597 = n1949 | n1950;
  assign n53598 = n1953 | n1954;
  assign n53599 = n1979 | n1967 | n1978;
  assign n53600 = n1995 | n1996;
  assign n53601 = n2017 | n2025 | n2035 | n2036;
  assign n53602 = n2050 | n2046 | n2049;
  assign n53603 = n2068 | n2081 | n2090 | n2091;
  assign n53604 = n2078 | n2079;
  assign n53605 = n2107 | n2108;
  assign n53606 = n2115 | n2112 | n2114;
  assign n53607 = n2139 | n2126 | n2138;
  assign n53608 = n2135 | n2136;
  assign n53609 = n2151 | n2148 | n2150;
  assign n53610 = n2155 | n2156;
  assign n53611 = n2159 | n2160;
  assign n53612 = n2170 | n2171;
  assign n53613 = n2185 | n2180 | n2184;
  assign n53614 = n2191 | n2192;
  assign n53615 = n2198 | n2195 | n2197;
  assign n53616 = n2230 | n2217 | n2229;
  assign n53617 = n2246 | n2247;
  assign n53618 = n2250 | n2251;
  assign n53619 = n2254 | n2255;
  assign n53620 = n2261 | n2262;
  assign n53621 = n2268 | n2265 | n2267;
  assign n53622 = n2323 | ~n2324 | ~n2297 | n2283 | ~n2296;
  assign n53623 = n2288 | n2289;
  assign n53624 = n2315 | n2308 | n2314;
  assign n53625 = n2331 | n2332;
  assign n53626 = n2336 | n2337;
  assign n53627 = n2351 | n2359 | n2365 | n2366;
  assign n53628 = n2355 | n2356;
  assign n53629 = n2370 | n2371;
  assign n53630 = n2376 | n2377;
  assign n53631 = n2379 | n2380;
  assign n53632 = n2381 | n2382;
  assign n53633 = n2386 | n2387;
  assign n53634 = n2393 | n2394;
  assign n53635 = n2399 | n2396 | n2398;
  assign n53636 = n2411 | n2412;
  assign n53637 = n2415 | n2416;
  assign n53638 = n2418 | n2419;
  assign n53639 = n2426 | n2427;
  assign n53640 = n2441 | n2442;
  assign n53641 = n2447 | n2448;
  assign n53642 = n2451 | n2452;
  assign n53643 = n2458 | n2459;
  assign n53644 = n2474 | n2466 | n2473;
  assign n53645 = n2488 | n2483 | n2487;
  assign n53646 = n2495 | n2496;
  assign n53647 = n2499 | n2500;
  assign n53648 = n2509 | n2513 | n2517 | n2518;
  assign n53649 = n2524 | n2525;
  assign n53650 = n2534 | n2535;
  assign n53651 = n2554 | n2555;
  assign n53652 = n2565 | n2556 | n2564;
  assign n53653 = n2575 | n2576;
  assign n53654 = n2583 | n2584;
  assign n53655 = n2605 | n2595 | n2604;
  assign n53656 = n2608 | n2609;
  assign n53657 = n2624 | n2625;
  assign n53658 = n2634 | n2631 | n2633;
  assign n53659 = n2644 | n2645;
  assign n53660 = n2648 | n2649;
  assign n53661 = n2651 | n2652;
  assign n53662 = n2656 | n2657;
  assign n53663 = n2660 | n2661;
  assign n53664 = n2671 | n2672;
  assign n53665 = n2689 | n2682 | n2688;
  assign n53666 = n2698 | n2699;
  assign n53667 = n2725 | n2711 | n2724;
  assign n53668 = n2738 | n2739;
  assign n53669 = n2748 | n2749;
  assign n53670 = n2770 | n2759 | n2769;
  assign n53671 = n2762 | n2763;
  assign n53672 = n2767 | n2768;
  assign n53673 = n2779 | n2775 | n2778;
  assign n53674 = n2791 | n2787 | n2790;
  assign n53675 = n2794 | n2795;
  assign n53676 = n2798 | n2799;
  assign n53677 = n2812 | n2813;
  assign n53678 = n2818 | n2819;
  assign n53679 = n2825 | n2822 | n2824;
  assign n53680 = n2837 | n2838;
  assign n53681 = n2848 | n2842 | n2847;
  assign n53682 = n2850 | n2851;
  assign n53683 = n2859 | n2860;
  assign n53684 = n2871 | n2863 | n2870;
  assign n53685 = n2890 | n2876 | n2889;
  assign n53686 = n2894 | n2895;
  assign n53687 = n2904 | n2905;
  assign n53688 = n2911 | n2912;
  assign n53689 = n2924 | n2921 | n2923;
  assign n53690 = n2932 | n2939 | n2947 | n2948;
  assign n53691 = n2952 | n2953;
  assign n53692 = n2958 | n2959;
  assign n53693 = n2972 | n2973;
  assign n53694 = n2985 | n2986;
  assign n53695 = n2991 | n2992;
  assign n53696 = n2998 | n2999;
  assign n53697 = n3004 | n3005;
  assign n53698 = n3009 | n3010;
  assign n53699 = n3018 | n3019;
  assign n53700 = n3038 | n3047 | n3058 | n3059;
  assign n53701 = n3069 | n3070;
  assign n53702 = n3081 | n3077 | n3080;
  assign n53703 = n3097 | n3109 | n3123 | n3124;
  assign n53704 = n3133 | n3129 | n3132;
  assign n53705 = n3138 | n3139;
  assign n53706 = n3145 | n3142 | n3144;
  assign n53707 = n3151 | n3148 | n3150;
  assign n53708 = n3159 | n3160;
  assign n53709 = n3163 | n3164;
  assign n53710 = n3169 | n3170;
  assign n53711 = n3176 | n3182 | n3188 | n3189;
  assign n53712 = n3212 | n3209 | n3211;
  assign n53713 = n3215 | n3216;
  assign n53714 = n3226 | n3223 | n3225;
  assign n53715 = n3231 | n3232;
  assign n53716 = n3240 | n3245 | n3250 | n3251;
  assign n53717 = n3271 | n3267 | n3270;
  assign n53718 = n3281 | n3282;
  assign n53719 = n3286 | n3287;
  assign n53720 = n3295 | n3292 | n3294;
  assign n53721 = n3307 | n3308;
  assign n53722 = n3311 | n3312;
  assign n53723 = n3332 | n3317 | n3331;
  assign n53724 = n3338 | n3339;
  assign n53725 = n3345 | n3342 | n3344;
  assign n53726 = n3368 | n3356 | n3367;
  assign n53727 = n3360 | n3361;
  assign n53728 = n3364 | n3365;
  assign n53729 = n3376 | n3377;
  assign n53730 = n3384 | n3385;
  assign n53731 = n3396 | n3397;
  assign n53732 = n3420 | n3407 | n3419;
  assign n53733 = n3434 | n3435;
  assign n53734 = n3438 | n3439;
  assign n53735 = n3445 | n3442 | n3444;
  assign n53736 = n3455 | n3459 | n3461 | n3462;
  assign n53737 = n3469 | n3466 | n3468;
  assign n53738 = n3472 | n3473;
  assign n53739 = n3479 | n3480;
  assign n53740 = n3500 | n3492 | n3499;
  assign n53741 = n3519 | n3520;
  assign n53742 = n3533 | n3534;
  assign n53743 = n3543 | n3550 | n3558 | n3559;
  assign n53744 = n3573 | n3574;
  assign n53745 = n3584 | n3591 | n3599 | n3600;
  assign n53746 = n3603 | n3604;
  assign n53747 = n3611 | n3612;
  assign n53748 = n3619 | n3620;
  assign n53749 = n3634 | n3635;
  assign n53750 = n3646 | n3643 | n3645;
  assign n53751 = n3648 | n3649;
  assign n53752 = n3652 | n3653;
  assign n53753 = n3659 | n3656 | n3658;
  assign n53754 = n3668 | n3669;
  assign n53755 = n3684 | n3685;
  assign n53756 = n3687 | n3688;
  assign n53757 = n3696 | n3702 | n3709 | n3710;
  assign n53758 = n3713 | n3714;
  assign n53759 = n3725 | n3731 | n3735 | n3736;
  assign n53760 = n3740 | n3741;
  assign n53761 = n3745 | n3746;
  assign n53762 = n3752 | n3749 | n3751;
  assign n53763 = n3758 | n3755 | n3757;
  assign n53764 = n3774 | n3775;
  assign n53765 = n3777 | n3778;
  assign n53766 = n3783 | n3784;
  assign n53767 = n3793 | n3789 | n3792;
  assign n53768 = n3797 | n3798;
  assign n53769 = n3808 | n3812 | n3817 | n3818;
  assign n53770 = n3829 | n3825 | n3828;
  assign n53771 = n3832 | n3833;
  assign n53772 = n3838 | n3839;
  assign n53773 = n3858 | n3849 | n3857;
  assign n53774 = n3874 | n3875;
  assign n53775 = n3886 | n3887;
  assign n53776 = n3915 | n3900 | n3907 | n3923 | n3924;
  assign n53777 = n3927 | n3928;
  assign n53778 = n3946 | n3941 | n3945;
  assign n53779 = n3943 | n3944;
  assign n53780 = n3979 | n3961 | n3978;
  assign n53781 = n3972 | n3973;
  assign n53782 = n3993 | n3994;
  assign n53783 = n3999 | n4000;
  assign n53784 = n4009 | n4006 | n4008;
  assign n53785 = n4019 | n4016 | n4018;
  assign n53786 = n4038 | n4033 | n4037;
  assign n53787 = n4068 | n4055 | n4067;
  assign n53788 = n4076 | n4079 | n4081 | n4082;
  assign n53789 = n4091 | n4088 | n4090;
  assign n53790 = n4099 | n4100;
  assign n53791 = n4110 | n4106 | n4109;
  assign n53792 = n4115 | n4116;
  assign n53793 = n4123 | n4124;
  assign n53794 = n4132 | n4133;
  assign n53795 = n4136 | n4137;
  assign n53796 = n4142 | n4143;
  assign n53797 = n4146 | n4147;
  assign n53798 = n4174 | n4159 | n4173;
  assign n53799 = n4195 | n4192 | n4194;
  assign n53800 = n4203 | n4200 | n4202;
  assign n53801 = n4210 | n4211;
  assign n53802 = n4217 | n4218;
  assign n53803 = n4221 | n4222;
  assign n53804 = n4229 | n4230;
  assign n53805 = n4242 | n4249 | n4256 | n4257;
  assign n53806 = n4266 | n4267;
  assign n53807 = n4273 | n4270 | n4272;
  assign n53808 = n4301 | n4288 | n4300;
  assign n53809 = n4304 | n4305;
  assign n53810 = n4308 | n4309;
  assign n53811 = n4328 | n4329;
  assign n53812 = n4331 | n4332;
  assign n53813 = n4338 | n4339;
  assign n53814 = n4345 | n4355 | n4359 | n4360;
  assign n53815 = n4366 | n4367;
  assign n53816 = n4374 | n4375;
  assign n53817 = n4391 | n4392;
  assign n53818 = n4408 | n4419 | n4435 | n4436;
  assign n53819 = n4454 | n4455;
  assign n53820 = n4467 | n4461 | n4466;
  assign n53821 = n4464 | n4465;
  assign n53822 = n4476 | n4477;
  assign n53823 = n4491 | n4483 | n4490;
  assign n53824 = n4499 | n4500;
  assign n53825 = n4506 | n4507;
  assign n53826 = n4510 | n4511;
  assign n53827 = n4523 | n4518 | n4522;
  assign n53828 = n4536 | n4537;
  assign n53829 = n4546 | n4543 | n4545;
  assign n53830 = n4551 | n4552;
  assign n53831 = n4565 | n4554 | n4564;
  assign n53832 = n4578 | n4579;
  assign n53833 = n4582 | n4583;
  assign n53834 = n4598 | n4599;
  assign n53835 = n4604 | n4605;
  assign n53836 = n4611 | n4608 | n4610;
  assign n53837 = n4631 | n4646 | n4661 | n4662;
  assign n53838 = n4678 | n4679;
  assign n53839 = n4682 | n4683;
  assign n53840 = n4695 | n4687 | n4694;
  assign n53841 = n4705 | n4702 | n4704;
  assign n53842 = n4736 | n4720 | n4727 | n4745 | n4746;
  assign n53843 = n4749 | n4750;
  assign n53844 = n4766 | n4761 | n4765;
  assign n53845 = n4783 | n4784;
  assign n53846 = n4788 | n4789;
  assign n53847 = n4801 | n4802;
  assign n53848 = n4816 | n4806 | n4815;
  assign n53849 = n4813 | n4809 | n4812;
  assign n53850 = n4822 | n4823;
  assign n53851 = n4825 | n4827 | n4830 | n4831;
  assign n53852 = n4843 | n4844;
  assign n53853 = n4869 | n4853 | n4860 | n4876 | n4877;
  assign n53854 = n4882 | n4883;
  assign n53855 = n4889 | n4890;
  assign n53856 = n4898 | n4899;
  assign n53857 = n4907 | n4908;
  assign n53858 = n4912 | n4913;
  assign n53859 = n4931 | n4932;
  assign n53860 = n4949 | n4950;
  assign n53861 = n4954 | n4955;
  assign n53862 = n4958 | n4959;
  assign n53863 = n4967 | n4962 | n4966;
  assign n53864 = n4964 | n4965;
  assign n53865 = n4970 | n4971;
  assign n53866 = n4985 | n4979 | n4984;
  assign n53867 = n4991 | n4988 | n4990;
  assign n53868 = n4996 | n4997;
  assign n53869 = n5017 | n5008 | n5016;
  assign n53870 = n5039 | n5032 | n5038;
  assign n53871 = n5042 | n5043;
  assign n53872 = n5056 | n5057;
  assign n53873 = n5063 | n5064;
  assign n53874 = n5067 | n5068;
  assign n53875 = n5071 | n5072;
  assign n53876 = n5091 | n5084 | n5090;
  assign n53877 = n5100 | n5096 | n5099;
  assign n53878 = n5112 | n5109 | n5111;
  assign n53879 = n5138 | n5127 | n5137;
  assign n53880 = n5150 | n5151;
  assign n53881 = n5161 | n5162;
  assign n53882 = n5179 | n5170 | n5178;
  assign n53883 = n5184 | n5185;
  assign n53884 = n5190 | n5187 | n5189;
  assign n53885 = n5193 | n5194;
  assign n53886 = n5212 | n5213;
  assign n53887 = n5222 | n5229 | n5234 | n5235;
  assign n53888 = n5253 | n5254;
  assign n53889 = n5260 | n5261;
  assign n53890 = n5270 | n5271;
  assign n53891 = n5275 | n5276;
  assign n53892 = n5315 | n5299 | n5314;
  assign n53893 = n5320 | n5321;
  assign n53894 = n5330 | n5331;
  assign n53895 = n5340 | n5336 | n5339;
  assign n53896 = n5343 | n5344;
  assign n53897 = n5347 | n5348;
  assign n53898 = n5356 | n5357;
  assign n53899 = n5367 | n5368;
  assign n53900 = n5371 | n5372;
  assign n53901 = n5375 | n5376;
  assign n53902 = n5381 | n5382;
  assign n53903 = n5385 | n5386;
  assign n53904 = n5397 | n5393 | n5396;
  assign n53905 = n5408 | n5409;
  assign n53906 = n5417 | n5418;
  assign n53907 = n5438 | n5439;
  assign n53908 = n5443 | n5444;
  assign n53909 = n5450 | n5451;
  assign n53910 = n5455 | n5456;
  assign n53911 = n5462 | n5463;
  assign n53912 = n5474 | n5475;
  assign n53913 = n5481 | n5478 | n5480;
  assign n53914 = n5501 | n5495 | n5500;
  assign n53915 = n5516 | n5517;
  assign n53916 = n5533 | n5534;
  assign n53917 = n5562 | n5550 | n5556 | n5569 | n5570;
  assign n53918 = n5581 | n5582;
  assign n53919 = n5585 | n5586;
  assign n53920 = n5611 | n5602 | n5610;
  assign n53921 = n5624 | n5625;
  assign n53922 = n5630 | n5631;
  assign n53923 = n5636 | n5637;
  assign n53924 = n5644 | n5647 | n5649 | n5650;
  assign n53925 = n5683 | n5671 | n5677 | n5688 | n5689;
  assign n53926 = n5698 | n5699;
  assign n53927 = n5702 | n5703;
  assign n53928 = n5708 | n5709;
  assign n53929 = n5713 | n5714;
  assign n53930 = n5731 | n5728 | n5730;
  assign n53931 = n5742 | n5738 | n5741;
  assign n53932 = n5746 | n5747;
  assign n53933 = n5754 | n5755;
  assign n53934 = n5767 | n5771 | n5781 | n5782;
  assign n53935 = n5788 | n5785 | n5787;
  assign n53936 = n5792 | n5793;
  assign n53937 = n5797 | n5798;
  assign n53938 = n5803 | n5804;
  assign n53939 = n5811 | n5812;
  assign n53940 = n5818 | n5820 | n5822 | n5823;
  assign n53941 = n5845 | n5834 | n5844;
  assign n53942 = n5853 | n5856 | n5858 | n5859;
  assign n53943 = n5863 | n5864;
  assign n53944 = n5870 | n5867 | n5869;
  assign n53945 = n5877 | n5878;
  assign n53946 = n5883 | n5884;
  assign n53947 = n5889 | n5890;
  assign n53948 = n5893 | n5894;
  assign n53949 = n5898 | n5899;
  assign n53950 = n5902 | n5903;
  assign n53951 = n5911 | n5912;
  assign n53952 = n5917 | n5914 | n5916;
  assign n53953 = n5922 | n5923;
  assign n53954 = n5927 | n5928;
  assign n53955 = n5934 | n5937 | n5940 | n5941;
  assign n53956 = n5946 | n5947;
  assign n53957 = n5964 | n5965;
  assign n53958 = n5980 | n5968 | n5974 | n5982 | n5983;
  assign n53959 = n5994 | n5995;
  assign n53960 = n6003 | n6004;
  assign n53961 = n6035 | n6020 | n6034;
  assign n53962 = n6050 | n6051;
  assign n53963 = n6063 | n6059 | n6062;
  assign n53964 = n6069 | n6066 | n6068;
  assign n53965 = n6081 | n6078 | n6080;
  assign n53966 = n6092 | n6100 | n6109 | n6110;
  assign n53967 = n6116 | n6113 | n6115;
  assign n53968 = n6123 | n6124;
  assign n53969 = n6129 | n6130;
  assign n53970 = n6147 | n6148;
  assign n53971 = n6188 | n6167 | n6187;
  assign n53972 = n6175 | n6171 | n6174;
  assign n53973 = n6182 | n6178 | n6181;
  assign n53974 = n6185 | n6186;
  assign n53975 = n6191 | n6192;
  assign n53976 = n6196 | n6197;
  assign n53977 = n6200 | n6201;
  assign n53978 = n6208 | n6209;
  assign n53979 = n6216 | n6217;
  assign n53980 = n6221 | n6222;
  assign n53981 = n6228 | n6229;
  assign n53982 = n6240 | n6233 | n6239;
  assign n53983 = n6237 | n6238;
  assign n53984 = n6246 | n6243 | n6245;
  assign n53985 = n6269 | n6258 | n6268;
  assign n53986 = n6286 | n6287;
  assign n53987 = n6291 | n6292;
  assign n53988 = n6298 | n6299;
  assign n53989 = n6307 | n6308;
  assign n53990 = n6320 | n6321;
  assign n53991 = n6338 | n6346 | n6354 | n6355;
  assign n53992 = n6358 | n6359;
  assign n53993 = n6366 | n6370 | n6373 | n6374;
  assign n53994 = n6379 | n6380;
  assign n53995 = n6393 | n6394;
  assign n53996 = n6399 | n6400;
  assign n53997 = n6406 | n6403 | n6405;
  assign n53998 = n6423 | n6431 | n6441 | n6442;
  assign n53999 = n6446 | n6449 | n6452 | n6453;
  assign n54000 = n6458 | n6459;
  assign n54001 = n6460 | n6461;
  assign n54002 = n6466 | n6467;
  assign n54003 = n6476 | n6477;
  assign n54004 = n6507 | n6495 | n6506;
  assign n54005 = n6527 | n6528;
  assign n54006 = n6533 | n6534;
  assign n54007 = n6538 | n6539;
  assign n54008 = n6542 | n6543;
  assign n54009 = n6552 | n6553;
  assign n54010 = n6560 | n6557 | n6559;
  assign n54011 = n6567 | n6568;
  assign n54012 = n6573 | n6574;
  assign n54013 = n6581 | n6582;
  assign n54014 = n6593 | n6594;
  assign n54015 = n6608 | n6609;
  assign n54016 = n6612 | n6613;
  assign n54017 = n6618 | n6619;
  assign n54018 = n6634 | n6630 | n6633;
  assign n54019 = n6653 | n6659 | n6669 | n6670;
  assign n54020 = n6675 | n6676;
  assign n54021 = n6682 | n6679 | n6681;
  assign n54022 = n6690 | n6687 | n6689;
  assign n54023 = n6695 | n6696;
  assign n54024 = n6706 | n6707;
  assign n54025 = n6713 | n6714;
  assign n54026 = n6720 | n6717 | n6719;
  assign n54027 = n6724 | n6725;
  assign n54028 = n6731 | n6732;
  assign n54029 = n6737 | n6738;
  assign n54030 = n6748 | n6749;
  assign n54031 = n6752 | n6753;
  assign n54032 = n6775 | n6761 | n6774;
  assign n54033 = n6772 | n6773;
  assign n54034 = n6792 | n6793;
  assign n54035 = n6797 | n6798;
  assign n54036 = n6803 | n6804;
  assign n54037 = n6817 | n6818;
  assign n54038 = n6824 | n6821 | n6823;
  assign n54039 = n6840 | n6841;
  assign n54040 = n6857 | n6858;
  assign n54041 = n6864 | n6865;
  assign n54042 = n6872 | n6869 | n6871;
  assign n54043 = n6880 | n6881;
  assign n54044 = n6882 | n6883;
  assign n54045 = n6889 | n6890;
  assign n54046 = n6896 | n6893 | n6895;
  assign n54047 = n6900 | n6901;
  assign n54048 = n6904 | n6905;
  assign n54049 = n6908 | n6909;
  assign n54050 = n6928 | n6925 | n6927;
  assign n54051 = n6932 | n6933;
  assign n54052 = n6940 | n6937 | n6939;
  assign n54053 = n6949 | n6950;
  assign n54054 = n6958 | n6959;
  assign n54055 = n6967 | n6964 | n6966;
  assign n54056 = n6985 | n6976 | n6984;
  assign n54057 = n6979 | n6980;
  assign n54058 = n6996 | n6997;
  assign n54059 = n7002 | n7003;
  assign n54060 = n7008 | n7009;
  assign n54061 = n7013 | n7014;
  assign n54062 = n7022 | n7023;
  assign n54063 = n7043 | n7034 | n7042;
  assign n54064 = n7056 | n7051 | n7055;
  assign n54065 = n7060 | n7061;
  assign n54066 = n7070 | n7063 | n7067 | n7073 | n7074;
  assign n54067 = n7090 | n7091;
  assign n54068 = n7106 | n7107;
  assign n54069 = n7111 | n7112;
  assign n54070 = n7114 | n7115;
  assign n54071 = n7124 | n7120 | n7123;
  assign n54072 = n7143 | n7159 | n7175 | n7176;
  assign n54073 = n7199 | n7196 | n7198;
  assign n54074 = n7210 | n7211;
  assign n54075 = n7224 | n7235 | n7242 | n7243;
  assign n54076 = n7249 | n7246 | n7248;
  assign n54077 = n7252 | n7253;
  assign n54078 = n7269 | n7264 | n7268 | n7273 | n7274;
  assign n54079 = n7280 | n7281;
  assign n54080 = n7285 | n7286;
  assign n54081 = n7292 | n7293;
  assign n54082 = n7305 | n7306;
  assign n54083 = n7321 | n7322;
  assign n54084 = n7332 | n7333;
  assign n54085 = n7341 | n7342;
  assign n54086 = n7345 | n7346;
  assign n54087 = n7388 | n7368 | n7387;
  assign n54088 = n7378 | n7379;
  assign n54089 = n7383 | n7384;
  assign n54090 = n7394 | n7391 | n7393;
  assign n54091 = n7397 | n7398;
  assign n54092 = n7403 | n7404;
  assign n54093 = n7407 | n7408;
  assign n54094 = n7414 | n7415;
  assign n54095 = n7423 | n7424;
  assign n54096 = n7428 | n7429;
  assign n54097 = n7450 | n7439 | n7449;
  assign n54098 = n7468 | n7469;
  assign n54099 = n7486 | n7483 | n7485;
  assign n54100 = n7504 | n7493 | n7503;
  assign n54101 = n7501 | n7502;
  assign n54102 = n7524 | n7519 | n7523;
  assign n54103 = n7540 | n7548 | n7560 | n7561;
  assign n54104 = n7574 | n7575;
  assign n54105 = n7578 | n7579;
  assign n54106 = n7585 | n7582 | n7584;
  assign n54107 = n7590 | n7591;
  assign n54108 = n7600 | n7601;
  assign n54109 = n7611 | n7612;
  assign n54110 = n7618 | n7619;
  assign n54111 = n7630 | n7622 | n7629;
  assign n54112 = n7644 | n7645;
  assign n54113 = n7651 | n7652;
  assign n54114 = n7665 | n7671 | n7678 | n7679;
  assign n54115 = n7684 | n7685;
  assign n54116 = n7691 | n7692;
  assign n54117 = n7702 | n7707 | n7712 | n7713;
  assign n54118 = n7734 | n7727 | n7733;
  assign n54119 = n7752 | n7753;
  assign n54120 = n7758 | n7759;
  assign n54121 = n7768 | n7764 | n7767;
  assign n54122 = n7774 | n7771 | n7773;
  assign n54123 = n7777 | n7778;
  assign n54124 = n7781 | n7782;
  assign n54125 = n7785 | n7786;
  assign n54126 = n7792 | n7793;
  assign n54127 = n7795 | n7796;
  assign n54128 = n7799 | n7802 | n7804 | n7805;
  assign n54129 = n7808 | n7809;
  assign n54130 = n7815 | n7816;
  assign n54131 = n7822 | n7819 | n7821;
  assign n54132 = n7843 | n7844;
  assign n54133 = n7848 | n7849;
  assign n54134 = n7857 | n7854 | n7856;
  assign n54135 = n7876 | n7869 | n7875;
  assign n54136 = n7885 | n7886;
  assign n54137 = n7892 | n7889 | n7891;
  assign n54138 = n7898 | n7895 | n7897;
  assign n54139 = n7901 | n7902;
  assign n54140 = n7911 | n7912;
  assign n54141 = n7935 | n7919 | n7934;
  assign n54142 = n7920 | n7921;
  assign n54143 = n7932 | n7933;
  assign n54144 = n7950 | n7951;
  assign n54145 = n7986 | n7968 | n7976 | n7991 | n7992;
  assign n54146 = n7982 | n7983;
  assign n54147 = n7995 | n7996;
  assign n54148 = n8002 | n8003;
  assign n54149 = n8019 | n8010 | n8018;
  assign n54150 = n8040 | n8041;
  assign n54151 = n8044 | n8045;
  assign n54152 = n8051 | n8048 | n8050;
  assign n54153 = n8063 | n8064;
  assign n54154 = n8086 | n8087;
  assign n54155 = n8096 | n8097;
  assign n54156 = n8103 | n8100 | n8102;
  assign n54157 = n8117 | n8123 | n8131 | n8132;
  assign n54158 = n8147 | n8144 | n8146;
  assign n54159 = n8155 | n8152 | n8154;
  assign n54160 = n8183 | n8169 | n8182;
  assign n54161 = n8189 | n8190;
  assign n54162 = n8217 | n8230 | n8243 | n8244;
  assign n54163 = n8262 | n8263;
  assign n54164 = n8272 | n8273;
  assign n54165 = n8277 | n8278;
  assign n54166 = n8285 | n8286;
  assign n54167 = n8300 | n8294 | n8299;
  assign n54168 = n8317 | n8314 | n8316;
  assign n54169 = n8356 | n8339 | n8355;
  assign n54170 = n8360 | n8361;
  assign n54171 = n8377 | n8382 | n8387 | n8388;
  assign n54172 = n8424 | n8408 | n8423;
  assign n54173 = n8410 | n8411;
  assign n54174 = n8420 | n8421;
  assign n54175 = n8434 | n8430 | n8433;
  assign n54176 = n8441 | n8442;
  assign n54177 = n8449 | n8450;
  assign n54178 = n8462 | n8463;
  assign n54179 = n8466 | n8467;
  assign n54180 = n8474 | n8482 | n8487 | n8488;
  assign n54181 = n8491 | n8492;
  assign n54182 = n8508 | n8509;
  assign n54183 = n8528 | n8529;
  assign n54184 = n8531 | n8532;
  assign n54185 = n8535 | n8536;
  assign n54186 = n8542 | n8543;
  assign n54187 = n8558 | n8562 | n8574 | n8575;
  assign n54188 = n8578 | n8579;
  assign n54189 = n8582 | n8583;
  assign n54190 = n8589 | n8586 | n8588;
  assign n54191 = n8595 | n8592 | n8594;
  assign n54192 = n8603 | n8600 | n8602;
  assign n54193 = n8611 | n8612;
  assign n54194 = n8629 | n8630;
  assign n54195 = n8644 | n8645;
  assign n54196 = n8654 | n8655;
  assign n54197 = n8667 | n8672 | n8676 | n8677;
  assign n54198 = n8684 | n8687 | n8690 | n8691;
  assign n54199 = n8718 | n8710 | n8717;
  assign n54200 = n8731 | n8732;
  assign n54201 = n8750 | n8751;
  assign n54202 = n8757 | n8758;
  assign n54203 = n8764 | n8765;
  assign n54204 = n8781 | n8773 | n8779 | n8787 | n8788;
  assign n54205 = n8791 | n8792;
  assign n54206 = n8796 | n8797;
  assign n54207 = n8800 | n8801;
  assign n54208 = n8814 | n8809 | n8813;
  assign n54209 = n8811 | n8812;
  assign n54210 = n8819 | n8820;
  assign n54211 = n8839 | n8832 | n8838;
  assign n54212 = n8856 | n8857;
  assign n54213 = n8868 | n8869;
  assign n54214 = n8894 | n8883 | n8893;
  assign n54215 = n8897 | n8898;
  assign n54216 = n8908 | n8913 | n8918 | n8919;
  assign n54217 = n8926 | n8927;
  assign n54218 = n8955 | n8947 | n8954;
  assign n54219 = n8962 | n8963;
  assign n54220 = n8968 | n8969;
  assign n54221 = n8990 | n8981 | n8989;
  assign n54222 = n8996 | n8993 | n8995;
  assign n54223 = n8999 | n9000;
  assign n54224 = n9009 | n9005 | n9008;
  assign n54225 = n9020 | n9025 | n9029 | n9030;
  assign n54226 = n9035 | n9036;
  assign n54227 = n9049 | n9050;
  assign n54228 = n9063 | n9057 | n9062;
  assign n54229 = n9060 | n9061;
  assign n54230 = n9066 | n9067;
  assign n54231 = n9073 | n9070 | n9072;
  assign n54232 = n9076 | n9077;
  assign n54233 = n9083 | n9080 | n9082;
  assign n54234 = n9090 | n9091;
  assign n54235 = n9094 | n9095;
  assign n54236 = n9104 | n9105;
  assign n54237 = n9109 | n9110;
  assign n54238 = n9112 | n9113;
  assign n54239 = n9127 | n9128;
  assign n54240 = n9146 | n9147;
  assign n54241 = n9153 | n9154;
  assign n54242 = n9164 | n9170 | n9177 | n9178;
  assign n54243 = n9181 | n9182;
  assign n54244 = n9194 | n9195;
  assign n54245 = n9202 | n9197 | n9199 | n9206 | n9207;
  assign n54246 = n9234 | n9223 | n9233;
  assign n54247 = n9245 | n9246;
  assign n54248 = n9248 | n9249;
  assign n54249 = n9270 | n9271;
  assign n54250 = n9304 | n9282 | n9291 | n9314 | n9315;
  assign n54251 = n9328 | n9329;
  assign n54252 = n9334 | n9335;
  assign n54253 = n9370 | n9355 | n9369;
  assign n54254 = n9392 | n9393;
  assign n54255 = n9403 | n9404;
  assign n54256 = n9415 | n9411 | n9414;
  assign n54257 = n9430 | n9435 | n9447 | n9448;
  assign n54258 = n9451 | n9452;
  assign n54259 = n9465 | n9460 | n9464;
  assign n54260 = n9472 | n9469 | n9471;
  assign n54261 = n9475 | n9476;
  assign n54262 = n9488 | n9489;
  assign n54263 = n9506 | n9498 | n9505;
  assign n54264 = n9524 | n9525;
  assign n54265 = n9529 | n9530;
  assign n54266 = n9543 | n9544;
  assign n54267 = n9552 | n9545 | n9551;
  assign n54268 = n9565 | n9566;
  assign n54269 = n9585 | n9586;
  assign n54270 = n9593 | n9594;
  assign n54271 = n9607 | n9613 | n9620 | n9621;
  assign n54272 = n9625 | n9626;
  assign n54273 = n9629 | n9630;
  assign n54274 = n9637 | n9638;
  assign n54275 = n9644 | n9645;
  assign n54276 = n9673 | n9662 | n9672;
  assign n54277 = n9690 | n9691;
  assign n54278 = n9695 | n9696;
  assign n54279 = n9705 | n9701 | n9704;
  assign n54280 = n9710 | n9707 | n9709;
  assign n54281 = n9715 | n9716;
  assign n54282 = n9728 | n9729;
  assign n54283 = n9738 | n9734 | n9737;
  assign n54284 = n9744 | n9745;
  assign n54285 = n9754 | n9749 | n9753;
  assign n54286 = n9760 | n9757 | n9759;
  assign n54287 = n9770 | n9771;
  assign n54288 = n9780 | n9781;
  assign n54289 = n9790 | n9791;
  assign n54290 = n9807 | n9808;
  assign n54291 = n9814 | n9815;
  assign n54292 = n9820 | n9821;
  assign n54293 = n9835 | n9836;
  assign n54294 = n9849 | n9850;
  assign n54295 = n9853 | n9854;
  assign n54296 = n9860 | n9857 | n9859;
  assign n54297 = n9865 | n9866;
  assign n54298 = n9872 | n9873;
  assign n54299 = n9884 | n9889 | n9896 | n9897;
  assign n54300 = n9901 | n9902;
  assign n54301 = n9908 | n9909;
  assign n54302 = n9919 | n9920;
  assign n54303 = n9926 | n9923 | n9925;
  assign n54304 = n9942 | n9943;
  assign n54305 = n9964 | n9965;
  assign n54306 = n9975 | n9976;
  assign n54307 = n9989 | n9994 | n9999 | n10000;
  assign n54308 = n9996 | n9997;
  assign n54309 = n10009 | n10010;
  assign n54310 = n10013 | n10014;
  assign n54311 = n10016 | n10017;
  assign n54312 = n10029 | n10030;
  assign n54313 = n10034 | n10035;
  assign n54314 = n10047 | n10048;
  assign n54315 = n10053 | n10054;
  assign n54316 = n10073 | n10064 | n10072;
  assign n54317 = n10086 | n10087;
  assign n54318 = n10104 | n10116 | n10131 | n10132;
  assign n54319 = n10144 | n10145;
  assign n54320 = n10152 | n10159 | n10165 | n10166;
  assign n54321 = n10172 | n10173;
  assign n54322 = n10178 | n10179;
  assign n54323 = n10187 | n10188;
  assign n54324 = n10201 | n10202;
  assign n54325 = n10225 | n10222 | n10224;
  assign n54326 = n10231 | n10232;
  assign n54327 = n10235 | n10236;
  assign n54328 = n10250 | n10251;
  assign n54329 = n10257 | n10254 | n10256;
  assign n54330 = n10262 | n10263;
  assign n54331 = n10277 | n10278;
  assign n54332 = n10288 | n10285 | n10287;
  assign n54333 = n10291 | n10292;
  assign n54334 = n10296 | n10297;
  assign n54335 = n10305 | n10306;
  assign n54336 = n10311 | n10312;
  assign n54337 = n10318 | n10319;
  assign n54338 = n10327 | n10335 | n10342 | n10343;
  assign n54339 = n10351 | n10347 | n10350;
  assign n54340 = n10357 | n10354 | n10356;
  assign n54341 = n10362 | n10363;
  assign n54342 = n10366 | n10367;
  assign n54343 = n10388 | n10378 | n10387;
  assign n54344 = n10404 | n10405;
  assign n54345 = n10409 | n10410;
  assign n54346 = n10411 | ~n10412;
  assign n54347 = n10542 | n10543;
  assign n54348 = n10544 | ~n10545;
  assign n54349 = n10549 | n10550;
  assign n54350 = n10553 | n10554;
  assign n54351 = n10555 | ~n10556;
  assign n54352 = n10562 | ~n10563;
  assign n54353 = ~n10573 | n10569 | ~n10572;
  assign n54354 = n10582 | n10583;
  assign n54355 = n10589 | n10586 | n10588;
  assign n54356 = n10603 | n10604;
  assign n54357 = n10609 | n10610;
  assign n54358 = n10613 | n10614;
  assign n54359 = n10627 | n10628;
  assign n54360 = n10634 | n10631 | n10633;
  assign n54361 = n10660 | n10670 | n10683 | n10684;
  assign n54362 = n10692 | n10689 | n10691;
  assign n54363 = n10695 | n10696;
  assign n54364 = n10728 | n10711 | n10727;
  assign n54365 = n10714 | n10715;
  assign n54366 = n10725 | n10726;
  assign n54367 = n10735 | n10736;
  assign n54368 = n10748 | n10753 | n10763 | n10764;
  assign n54369 = n10783 | n10784;
  assign n54370 = n10792 | n10793;
  assign n54371 = n10798 | n10799;
  assign n54372 = n10805 | n10802 | n10804;
  assign n54373 = n10811 | n10808 | n10810;
  assign n54374 = n10819 | n10820;
  assign n54375 = n10823 | n10824;
  assign n54376 = n10836 | n10837;
  assign n54377 = n10865 | n10852 | n10864;
  assign n54378 = n10878 | n10879;
  assign n54379 = n10884 | n10885;
  assign n54380 = n10899 | n10893 | n10898;
  assign n54381 = n10938 | n10926 | n10934 | n10948 | n10949;
  assign n54382 = n10955 | n10956;
  assign n54383 = n10986 | n10971 | n10985;
  assign n54384 = n11005 | n11006;
  assign n54385 = n11011 | n11012;
  assign n54386 = n11031 | n11021 | n11030;
  assign n54387 = n11025 | n11026;
  assign n54388 = n11037 | n11034 | n11036;
  assign n54389 = n11064 | n11065;
  assign n54390 = n11080 | n11066 | n11079;
  assign n54391 = n11096 | n11097;
  assign n54392 = n11106 | n11102 | n11105;
  assign n54393 = n11114 | n11115;
  assign n54394 = n11121 | n11122;
  assign n54395 = n11129 | n11130;
  assign n54396 = n11137 | n11138;
  assign n54397 = n11143 | n11144;
  assign n54398 = n11149 | n11150;
  assign n54399 = n11153 | n11154;
  assign n54400 = n11168 | n11177 | n11183 | n11184;
  assign n54401 = n11201 | n11202;
  assign n54402 = n11207 | n11208;
  assign n54403 = n11217 | n11218;
  assign n54404 = ~n11230 | n11226 | ~n11229;
  assign n54405 = n11232 | n11233;
  assign n54406 = n11253 | ~n11254;
  assign n54407 = n11265 | ~n11266;
  assign n54408 = n11268 | n11269;
  assign n54409 = n11274 | ~n11275;
  assign n54410 = n11277 | n11278;
  assign n54411 = n11282 | n11283;
  assign n54412 = n11293 | n11294;
  assign n54413 = n11301 | ~n11302;
  assign n54414 = n11306 | ~n11307;
  assign n54415 = n11309 | ~n11310;
  assign n54416 = n11316 | n11317;
  assign n54417 = n11323 | n11320 | n11322;
  assign n54418 = n11332 | n11328 | n11331;
  assign n54419 = n11340 | n11341;
  assign n54420 = n11354 | n11355;
  assign n54421 = n11367 | n11368;
  assign n54422 = n11371 | n11372;
  assign n54423 = n11387 | n11388;
  assign n54424 = n11393 | n11394;
  assign n54425 = n11398 | ~n11399;
  assign n54426 = n11408 | n11409;
  assign n54427 = n11410 | n11411;
  assign n54428 = n11416 | n11417;
  assign n54429 = n11425 | ~n11426;
  assign n54430 = n11448 | n11457 | n11467 | n11468;
  assign n54431 = n11487 | n11480 | n11486;
  assign n54432 = n11509 | n11502 | n11508;
  assign n54433 = n11512 | n11513;
  assign n54434 = n11528 | n11521 | n11527;
  assign n54435 = n11542 | n11543;
  assign n54436 = n11561 | n11554 | n11560;
  assign n54437 = n11565 | n11566;
  assign n54438 = n11569 | n11570;
  assign n54439 = n11583 | n11584;
  assign n54440 = n11592 | n11593;
  assign n54441 = n11602 | n11603;
  assign n54442 = n11606 | n11607;
  assign n54443 = n11621 | n11622;
  assign n54444 = n11625 | n11626;
  assign n54445 = n11632 | n11634 | n11637 | n11638;
  assign n54446 = n11644 | n11641 | n11643;
  assign n54447 = n11657 | n11658;
  assign n54448 = n11688 | n11673 | n11687;
  assign n54449 = n11703 | n11699 | n11702;
  assign n54450 = n11708 | n11709;
  assign n54451 = n11731 | n11746 | n11759 | n11760;
  assign n54452 = n11765 | n11766;
  assign n54453 = n11769 | n11770;
  assign n54454 = n11773 | n11774;
  assign n54455 = n11777 | n11778;
  assign n54456 = n11790 | n11787 | n11789;
  assign n54457 = n11801 | n11805 | n11811 | n11812;
  assign n54458 = n11826 | n11822 | n11825;
  assign n54459 = n11838 | n11839;
  assign n54460 = n11844 | n11845;
  assign n54461 = n11858 | n11847 | n11857;
  assign n54462 = n11877 | n11878;
  assign n54463 = n11883 | n11884;
  assign n54464 = n11896 | n11897;
  assign n54465 = ~n11905 | n11901 | n11904;
  assign n54466 = n11920 | n11921;
  assign n54467 = n11924 | n11925;
  assign n54468 = n11932 | n11929 | n11931;
  assign n54469 = n11936 | n11937;
  assign n54470 = n11939 | n11940;
  assign n54471 = n11946 | n11947;
  assign n54472 = n11959 | n11967 | n11975 | n11976;
  assign n54473 = n11984 | n11981 | n11983;
  assign n54474 = n11995 | n11996;
  assign n54475 = n12003 | n12004;
  assign n54476 = n12012 | n12013;
  assign n54477 = n12023 | n12020 | n12022;
  assign n54478 = n12029 | n12030;
  assign n54479 = n12043 | n12036 | n12042;
  assign n54480 = n12055 | n12056;
  assign n54481 = n12072 | n12073;
  assign n54482 = n12081 | n12082;
  assign n54483 = n12108 | n12098 | n12107;
  assign n54484 = n12119 | n12120;
  assign n54485 = n12142 | n12132 | n12141;
  assign n54486 = n12158 | n12165 | n12172 | n12173;
  assign n54487 = n12188 | n12189;
  assign n54488 = n12192 | n12193;
  assign n54489 = n12196 | n12197;
  assign n54490 = n12200 | n12201;
  assign n54491 = n12206 | n12207;
  assign n54492 = n12211 | n12212;
  assign n54493 = n12224 | n12218 | n12223;
  assign n54494 = n12237 | n12238;
  assign n54495 = n12257 | n12258;
  assign n54496 = n12265 | n12266;
  assign n54497 = n12269 | n12270;
  assign n54498 = n12285 | n12280 | n12284;
  assign n54499 = n12282 | n12283;
  assign n54500 = n12308 | n12316 | n12326 | n12327;
  assign n54501 = n12337 | n12334 | n12336;
  assign n54502 = n12362 | n12349 | n12361;
  assign n54503 = n12353 | n12354;
  assign n54504 = n12359 | n12360;
  assign n54505 = n12375 | n12376;
  assign n54506 = n12387 | n12398 | n12407 | n12408;
  assign n54507 = n12420 | n12421;
  assign n54508 = n12429 | n12430;
  assign n54509 = n12476 | n12457 | n12464 | n12488 | n12489;
  assign n54510 = n12498 | n12495 | n12497;
  assign n54511 = n12501 | n12502;
  assign n54512 = n12517 | n12510 | n12516;
  assign n54513 = n12521 | n12522;
  assign n54514 = n12539 | n12536 | n12538;
  assign n54515 = n12544 | n12545;
  assign n54516 = n12557 | n12558;
  assign n54517 = ~n12566 | n12562 | n12565;
  assign n54518 = n12568 | n12569;
  assign n54519 = n12578 | ~n12579;
  assign n54520 = n12592 | ~n12593;
  assign n54521 = n12604 | ~n12605;
  assign n54522 = n12613 | n12614;
  assign n54523 = n12617 | n12618;
  assign n54524 = n12619 | n12620;
  assign n54525 = n12625 | ~n12626;
  assign n54526 = n12630 | n12631;
  assign n54527 = n12632 | n12633;
  assign n54528 = n12634 | ~n12635;
  assign n54529 = n12643 | ~n12644;
  assign n54530 = n12646 | n12647;
  assign n54531 = n12648 | n12649;
  assign n54532 = n12657 | n12658;
  assign n54533 = n12661 | n12662;
  assign n54534 = n12663 | n12664;
  assign n54535 = n12672 | ~n12673;
  assign n54536 = n12679 | ~n12680;
  assign n54537 = n12687 | ~n12688;
  assign n54538 = n12699 | n12700;
  assign n54539 = n12704 | n12705;
  assign n54540 = n12715 | n12712 | n12714;
  assign n54541 = n12717 | n12718;
  assign n54542 = n12721 | n12722;
  assign n54543 = n12726 | n12727;
  assign n54544 = n12740 | n12746 | n12753 | n12754;
  assign n54545 = n12763 | n12759 | n12762;
  assign n54546 = n12790 | n12780 | n12789;
  assign n54547 = n12799 | n12800;
  assign n54548 = n12806 | n12810 | n12816 | n12817;
  assign n54549 = n12825 | n12826;
  assign n54550 = n12845 | n12837 | n12840 | n12850 | n12851;
  assign n54551 = n12864 | n12865;
  assign n54552 = n12876 | n12877;
  assign n54553 = n12883 | n12880 | n12882;
  assign n54554 = n12886 | n12887;
  assign n54555 = n12913 | n12910 | n12912;
  assign n54556 = n12925 | n12926;
  assign n54557 = n12929 | n12930;
  assign n54558 = n12945 | n12946;
  assign n54559 = n12951 | n12952;
  assign n54560 = n12956 | ~n12957;
  assign n54561 = n12967 | n12968;
  assign n54562 = n12971 | ~n12972;
  assign n54563 = n12979 | n12980;
  assign n54564 = n12981 | n12982;
  assign n54565 = n12983 | ~n12984;
  assign n54566 = n12997 | n12998;
  assign n54567 = n13001 | n13002;
  assign n54568 = n13003 | n13004;
  assign n54569 = n13009 | ~n13010;
  assign n54570 = n13018 | n13019;
  assign n54571 = n13020 | n13021;
  assign n54572 = n13026 | ~n13027;
  assign n54573 = n13039 | n13040;
  assign n54574 = n13043 | ~n13044;
  assign n54575 = n13054 | n13055;
  assign n54576 = n13058 | ~n13059;
  assign n54577 = n13066 | ~n13067;
  assign n54578 = n13076 | n13077;
  assign n54579 = n13080 | n13081;
  assign n54580 = n13082 | n13083;
  assign n54581 = n13088 | ~n13089;
  assign n54582 = n13092 | n13093;
  assign n54583 = n13094 | n13095;
  assign n54584 = n13096 | ~n13097;
  assign n54585 = n13098 | n13099;
  assign n54586 = n13100 | n13101;
  assign n54587 = n13106 | n13107;
  assign n54588 = n13114 | n13111 | n13113;
  assign n54589 = n13122 | n13123;
  assign n54590 = n13126 | n13127;
  assign n54591 = n13128 | n13129;
  assign n54592 = n13134 | ~n13135;
  assign n54593 = n13140 | ~n13141;
  assign n54594 = n13151 | n13148 | n13150;
  assign n54595 = n13160 | n13156 | n13159;
  assign n54596 = n13184 | n13175 | n13183;
  assign n54597 = n13204 | n13205;
  assign n54598 = n13212 | n13213;
  assign n54599 = n13229 | n13225 | n13228;
  assign n54600 = n13237 | n13238;
  assign n54601 = n13243 | n13244;
  assign n54602 = n13272 | n13261 | n13271;
  assign n54603 = n13279 | n13280;
  assign n54604 = n13292 | n13293;
  assign n54605 = n13305 | n13306;
  assign n54606 = n13324 | n13325;
  assign n54607 = n13330 | n13331;
  assign n54608 = n13343 | n13344;
  assign n54609 = ~n13352 | n13348 | ~n13351;
  assign n54610 = n13367 | n13368;
  assign n54611 = n13371 | n13372;
  assign n54612 = n13416 | n13400 | n13415;
  assign n54613 = n13419 | n13420;
  assign n54614 = n13462 | n13444 | n13452 | n13474 | n13475;
  assign n54615 = n13487 | n13482 | n13486;
  assign n54616 = n13493 | n13494;
  assign n54617 = n13515 | n13516;
  assign n54618 = n13522 | n13523;
  assign n54619 = n13542 | n13536 | n13541;
  assign n54620 = n13539 | n13540;
  assign n54621 = n13549 | n13550;
  assign n54622 = n13575 | n13563 | n13574;
  assign n54623 = n13588 | n13589;
  assign n54624 = n13596 | n13592 | n13595;
  assign n54625 = n13607 | n13608;
  assign n54626 = n13625 | n13637 | n13648 | n13649;
  assign n54627 = n13657 | n13654 | n13656;
  assign n54628 = n13676 | n13692 | n13704 | n13705;
  assign n54629 = n13689 | n13690;
  assign n54630 = n13711 | n13708 | n13710;
  assign n54631 = n13717 | n13714 | n13716;
  assign n54632 = n13724 | n13725;
  assign n54633 = n13733 | n13734;
  assign n54634 = n13741 | n13742;
  assign n54635 = n13761 | n13750 | n13760;
  assign n54636 = n13780 | n13781;
  assign n54637 = n13789 | n13786 | n13788;
  assign n54638 = n13806 | n13800 | n13805;
  assign n54639 = n13819 | n13820;
  assign n54640 = n13827 | n13828;
  assign n54641 = n13842 | n13843;
  assign n54642 = n13856 | n13857;
  assign n54643 = n13876 | n13894 | n13910 | n13911;
  assign n54644 = n13891 | n13892;
  assign n54645 = n13919 | n13920;
  assign n54646 = n13940 | n13931 | n13939;
  assign n54647 = n13948 | n13945 | n13947;
  assign n54648 = n13953 | n13954;
  assign n54649 = n13981 | n13971 | n13980;
  assign n54650 = n13973 | n13974;
  assign n54651 = n13988 | n13989;
  assign n54652 = n14008 | n14009;
  assign n54653 = n14014 | n14015;
  assign n54654 = n14027 | n14028;
  assign n54655 = ~n14036 | n14032 | ~n14035;
  assign n54656 = n14038 | n14039;
  assign n54657 = n14048 | ~n14049;
  assign n54658 = n14059 | n14060;
  assign n54659 = n14063 | ~n14064;
  assign n54660 = n14073 | n14074;
  assign n54661 = n14075 | n14076;
  assign n54662 = n14077 | ~n14078;
  assign n54663 = n14092 | n14093;
  assign n54664 = n14094 | n14095;
  assign n54665 = n14100 | ~n14101;
  assign n54666 = n14108 | ~n14109;
  assign n54667 = n14112 | n14113;
  assign n54668 = n14119 | n14120;
  assign n54669 = n14126 | n14127;
  assign n54670 = n14128 | n14129;
  assign n54671 = n14134 | ~n14135;
  assign n54672 = n14145 | n14146;
  assign n54673 = n14149 | ~n14150;
  assign n54674 = n14163 | n14164;
  assign n54675 = n14167 | ~n14168;
  assign n54676 = n14179 | n14180;
  assign n54677 = n14183 | n14184;
  assign n54678 = n14185 | n14186;
  assign n54679 = n14192 | n14193;
  assign n54680 = n14195 | n14196;
  assign n54681 = n14197 | n14198;
  assign n54682 = n14199 | ~n14200;
  assign n54683 = n14204 | n14205;
  assign n54684 = n14215 | n14216;
  assign n54685 = n14217 | n14218;
  assign n54686 = n14227 | ~n14228;
  assign n54687 = n14241 | n14242;
  assign n54688 = n14245 | ~n14246;
  assign n54689 = n14253 | ~n14254;
  assign n54690 = n14260 | ~n14261;
  assign n54691 = n14270 | n14271;
  assign n54692 = n14274 | n14275;
  assign n54693 = n14283 | n14284;
  assign n54694 = n14287 | n14288;
  assign n54695 = n14289 | n14290;
  assign n54696 = n14293 | n14294;
  assign n54697 = n14295 | n14296;
  assign n54698 = n14297 | ~n14298;
  assign n54699 = n14311 | n14312;
  assign n54700 = n14315 | n14316;
  assign n54701 = n14317 | n14318;
  assign n54702 = n14323 | n14324;
  assign n54703 = n14333 | n14334;
  assign n54704 = n14337 | n14338;
  assign n54705 = n14339 | n14340;
  assign n54706 = n14345 | n14346;
  assign n54707 = n14355 | n14356;
  assign n54708 = n14359 | n14360;
  assign n54709 = n14361 | n14362;
  assign n54710 = n14367 | n14368;
  assign n54711 = n14372 | n14373;
  assign n54712 = n14374 | n14375;
  assign n54713 = n14376 | ~n14377;
  assign n54714 = n14381 | n14382;
  assign n54715 = n14387 | ~n14388;
  assign n54716 = n14393 | ~n14394;
  assign n54717 = n14399 | ~n14400;
  assign n54718 = n14405 | ~n14406;
  assign n54719 = n14412 | n14409 | n14411;
  assign n54720 = n14419 | n14420;
  assign n54721 = n14430 | n14431;
  assign n54722 = n14434 | ~n14435;
  assign n54723 = n14442 | ~n14443;
  assign n54724 = n14453 | n14457 | n14459 | n14460;
  assign n54725 = n14463 | n14464;
  assign n54726 = n14473 | n14469 | n14472;
  assign n54727 = n14483 | n14484;
  assign n54728 = n14487 | n14488;
  assign n54729 = n14512 | n14503 | n14507 | n14516 | n14517;
  assign n54730 = n14533 | n14534;
  assign n54731 = n14541 | n14542;
  assign n54732 = n14552 | n14549 | n14551;
  assign n54733 = n14572 | n14583 | n14597 | n14598;
  assign n54734 = n14604 | n14601 | n14603;
  assign n54735 = n14609 | n14610;
  assign n54736 = n14635 | n14648 | n14664 | n14665;
  assign n54737 = n14682 | n14683;
  assign n54738 = n14695 | n14696;
  assign n54739 = n14699 | n14700;
  assign n54740 = n14715 | n14716;
  assign n54741 = n14721 | n14722;
  assign n54742 = n14726 | ~n14727;
  assign n54743 = n14737 | n14738;
  assign n54744 = n14741 | ~n14742;
  assign n54745 = n14751 | ~n14752;
  assign n54746 = n14761 | n14762;
  assign n54747 = n14765 | n14766;
  assign n54748 = n14767 | n14768;
  assign n54749 = n14773 | n14774;
  assign n54750 = n14780 | ~n14781;
  assign n54751 = n14792 | n14793;
  assign n54752 = n14794 | n14795;
  assign n54753 = n14800 | n14801;
  assign n54754 = n14807 | ~n14808;
  assign n54755 = n14812 | n14813;
  assign n54756 = n14820 | ~n14821;
  assign n54757 = n14828 | n14829;
  assign n54758 = n14832 | n14833;
  assign n54759 = n14834 | n14835;
  assign n54760 = n14841 | n14842;
  assign n54761 = n14843 | n14844;
  assign n54762 = n14845 | ~n14846;
  assign n54763 = n14850 | ~n14851;
  assign n54764 = n14858 | n14859;
  assign n54765 = n14862 | n14863;
  assign n54766 = n14864 | n14865;
  assign n54767 = n14870 | ~n14871;
  assign n54768 = n14876 | ~n14877;
  assign n54769 = n14883 | n14880 | n14882;
  assign n54770 = n14889 | n14890;
  assign n54771 = n14892 | n14893;
  assign n54772 = n14899 | n14896 | n14898;
  assign n54773 = n14902 | n14903;
  assign n54774 = n14913 | n14914;
  assign n54775 = n14918 | n14919;
  assign n54776 = n14935 | n14931 | n14934;
  assign n54777 = n14964 | n14953 | n14963;
  assign n54778 = n14970 | n14971;
  assign n54779 = n14987 | n14991 | n15001 | n15002;
  assign n54780 = n15017 | n15018;
  assign n54781 = n15023 | n15024;
  assign n54782 = n15032 | n15028 | n15031;
  assign n54783 = n15038 | n15035 | n15037;
  assign n54784 = n15045 | n15046;
  assign n54785 = n15055 | n15052 | n15054;
  assign n54786 = n15074 | n15083 | n15098 | n15099;
  assign n54787 = n15115 | n15116;
  assign n54788 = n15159 | n15143 | n15158;
  assign n54789 = n15183 | n15184;
  assign n54790 = n15189 | n15190;
  assign n54791 = n15202 | n15203;
  assign n54792 = ~n15211 | n15207 | ~n15210;
  assign n54793 = n15228 | n15229;
  assign n54794 = n15236 | n15237;
  assign n54795 = n15240 | n15241;
  assign n54796 = n15253 | n15250 | n15252;
  assign n54797 = n15259 | n15260;
  assign n54798 = n15281 | n15270 | n15280;
  assign n54799 = n15299 | n15300;
  assign n54800 = n15305 | n15306;
  assign n54801 = n15311 | n15312;
  assign n54802 = n15333 | n15327 | n15332;
  assign n54803 = n15363 | n15350 | n15362;
  assign n54804 = n15366 | n15367;
  assign n54805 = n15383 | n15384;
  assign n54806 = n15387 | n15388;
  assign n54807 = n15404 | n15395 | n15403;
  assign n54808 = n15419 | n15420;
  assign n54809 = n15427 | n15428;
  assign n54810 = n15433 | n15434;
  assign n54811 = n15451 | n15452;
  assign n54812 = n15460 | n15461;
  assign n54813 = n15474 | n15468 | n15473;
  assign n54814 = n15482 | n15483;
  assign n54815 = n15492 | n15488 | n15491;
  assign n54816 = n15496 | n15497;
  assign n54817 = n15503 | n15504;
  assign n54818 = n15520 | n15521;
  assign n54819 = n15537 | n15538;
  assign n54820 = n15552 | n15553;
  assign n54821 = n15564 | n15561 | n15563;
  assign n54822 = n15572 | n15569 | n15571;
  assign n54823 = n15580 | n15581;
  assign n54824 = n15593 | n15587 | n15592;
  assign n54825 = n15601 | n15602;
  assign n54826 = n15605 | n15606;
  assign n54827 = n15624 | n15639 | n15648 | n15649;
  assign n54828 = n15633 | n15634;
  assign n54829 = n15654 | n15655;
  assign n54830 = n15679 | n15670 | n15678;
  assign n54831 = n15704 | n15693 | n15697 | n15710 | n15711;
  assign n54832 = n15720 | n15721;
  assign n54833 = n15723 | n15724;
  assign n54834 = n15732 | n15728 | n15731;
  assign n54835 = n15748 | n15739 | n15747;
  assign n54836 = n15745 | n15746;
  assign n54837 = n15767 | n15768;
  assign n54838 = n15773 | n15774;
  assign n54839 = n15789 | n15786 | n15788;
  assign n54840 = ~n15797 | n15793 | ~n15796;
  assign n54841 = n15799 | n15800;
  assign n54842 = n15809 | ~n15810;
  assign n54843 = n15820 | n15821;
  assign n54844 = n15824 | ~n15825;
  assign n54845 = n15834 | n15835;
  assign n54846 = n15836 | n15837;
  assign n54847 = n15838 | ~n15839;
  assign n54848 = n15852 | n15853;
  assign n54849 = n15856 | n15857;
  assign n54850 = n15858 | n15859;
  assign n54851 = n15864 | n15865;
  assign n54852 = n15874 | n15875;
  assign n54853 = n15878 | n15879;
  assign n54854 = n15880 | n15881;
  assign n54855 = n15886 | n15887;
  assign n54856 = n15890 | n15891;
  assign n54857 = n15892 | n15893;
  assign n54858 = n15895 | ~n15896;
  assign n54859 = n15906 | n15907;
  assign n54860 = n15908 | n15909;
  assign n54861 = n15914 | n15915;
  assign n54862 = n15926 | n15927;
  assign n54863 = n15930 | ~n15931;
  assign n54864 = n15938 | ~n15939;
  assign n54865 = n15948 | n15949;
  assign n54866 = n15952 | ~n15953;
  assign n54867 = n15968 | n15969;
  assign n54868 = n15972 | ~n15973;
  assign n54869 = n15984 | n15985;
  assign n54870 = n15988 | n15989;
  assign n54871 = n15990 | n15991;
  assign n54872 = n15997 | n15998;
  assign n54873 = n16004 | ~n16005;
  assign n54874 = n16014 | n16015;
  assign n54875 = n16018 | n16019;
  assign n54876 = n16020 | n16021;
  assign n54877 = n16026 | n16027;
  assign n54878 = n16036 | n16037;
  assign n54879 = n16040 | n16041;
  assign n54880 = n16042 | n16043;
  assign n54881 = n16048 | n16049;
  assign n54882 = n16060 | ~n16061;
  assign n54883 = n16071 | ~n16072;
  assign n54884 = n16077 | ~n16078;
  assign n54885 = n16085 | ~n16086;
  assign n54886 = n16089 | n16090;
  assign n54887 = n16095 | n16096;
  assign n54888 = n16106 | n16107;
  assign n54889 = n16110 | n16111;
  assign n54890 = n16112 | n16113;
  assign n54891 = n16119 | n16120;
  assign n54892 = n16121 | n16122;
  assign n54893 = n16123 | ~n16124;
  assign n54894 = n16128 | ~n16129;
  assign n54895 = n16135 | ~n16136;
  assign n54896 = n16147 | n16148;
  assign n54897 = n16156 | n16157;
  assign n54898 = n16160 | n16161;
  assign n54899 = n16162 | n16163;
  assign n54900 = n16166 | n16167;
  assign n54901 = n16168 | n16169;
  assign n54902 = n16170 | ~n16171;
  assign n54903 = n16184 | n16185;
  assign n54904 = n16188 | n16189;
  assign n54905 = n16190 | n16191;
  assign n54906 = n16196 | n16197;
  assign n54907 = n16206 | n16207;
  assign n54908 = n16210 | n16211;
  assign n54909 = n16212 | n16213;
  assign n54910 = n16218 | n16219;
  assign n54911 = n16228 | n16229;
  assign n54912 = n16232 | n16233;
  assign n54913 = n16234 | n16235;
  assign n54914 = n16240 | n16241;
  assign n54915 = n16244 | n16245;
  assign n54916 = n16246 | n16247;
  assign n54917 = n16249 | ~n16250;
  assign n54918 = n16261 | n16262;
  assign n54919 = n16263 | n16264;
  assign n54920 = n16269 | n16270;
  assign n54921 = n16276 | ~n16277;
  assign n54922 = n16281 | n16282;
  assign n54923 = n16287 | ~n16288;
  assign n54924 = n16297 | n16298;
  assign n54925 = n16301 | ~n16302;
  assign n54926 = n16312 | ~n16313;
  assign n54927 = n16320 | n16321;
  assign n54928 = n16324 | ~n16325;
  assign n54929 = n16332 | ~n16333;
  assign n54930 = n16342 | n16339 | n16341;
  assign n54931 = n16362 | n16363;
  assign n54932 = n16375 | n16372 | n16374;
  assign n54933 = n16392 | n16401 | n16415 | n16416;
  assign n54934 = n16408 | n16409;
  assign n54935 = n16435 | n16436;
  assign n54936 = n16442 | n16443;
  assign n54937 = n16470 | n16457 | n16469;
  assign n54938 = n16473 | n16474;
  assign n54939 = n16489 | n16482 | n16488;
  assign n54940 = n16509 | n16510;
  assign n54941 = n16515 | ~n16516;
  assign n54942 = n16529 | n16530;
  assign n54943 = n16535 | n16536;
  assign n54944 = n16538 | n16539;
  assign n54945 = n16554 | n16555;
  assign n54946 = n16560 | n16561;
  assign n54947 = n16565 | ~n16566;
  assign n54948 = n16576 | n16577;
  assign n54949 = n16580 | ~n16581;
  assign n54950 = n16590 | ~n16591;
  assign n54951 = n16600 | n16601;
  assign n54952 = n16604 | n16605;
  assign n54953 = n16606 | n16607;
  assign n54954 = n16612 | n16613;
  assign n54955 = n16619 | ~n16620;
  assign n54956 = n16629 | n16630;
  assign n54957 = n16633 | n16634;
  assign n54958 = n16635 | n16636;
  assign n54959 = n16641 | n16642;
  assign n54960 = n16651 | n16652;
  assign n54961 = n16655 | n16656;
  assign n54962 = n16657 | n16658;
  assign n54963 = n16663 | n16664;
  assign n54964 = n16670 | ~n16671;
  assign n54965 = n16681 | n16682;
  assign n54966 = n16683 | n16684;
  assign n54967 = n16689 | n16690;
  assign n54968 = n16701 | n16702;
  assign n54969 = n16705 | ~n16706;
  assign n54970 = n16713 | ~n16714;
  assign n54971 = n16721 | n16722;
  assign n54972 = n16725 | n16726;
  assign n54973 = n16727 | n16728;
  assign n54974 = n16734 | n16735;
  assign n54975 = n16736 | n16737;
  assign n54976 = n16738 | ~n16739;
  assign n54977 = n16743 | ~n16744;
  assign n54978 = n16751 | n16752;
  assign n54979 = n16755 | n16756;
  assign n54980 = n16757 | n16758;
  assign n54981 = n16763 | ~n16764;
  assign n54982 = n16769 | ~n16770;
  assign n54983 = n16779 | n16780;
  assign n54984 = n16783 | n16784;
  assign n54985 = n16789 | ~n16790;
  assign n54986 = n16793 | n16794;
  assign n54987 = n16806 | n16800 | n16805;
  assign n54988 = n16816 | n16813 | n16815;
  assign n54989 = n16821 | n16822;
  assign n54990 = n16828 | n16829;
  assign n54991 = n16854 | n16844 | n16853;
  assign n54992 = n16871 | n16872;
  assign n54993 = n16880 | n16881;
  assign n54994 = n16892 | n16888 | n16891;
  assign n54995 = n16907 | n16908;
  assign n54996 = n16927 | n16928;
  assign n54997 = n16943 | n16944;
  assign n54998 = n16961 | n16952 | n16960;
  assign n54999 = n16975 | n16976;
  assign n55000 = n16990 | n16995 | n16999 | n17000;
  assign n55001 = n17018 | n17011 | n17017;
  assign n55002 = n17035 | n17036;
  assign n55003 = n17048 | n17049;
  assign n55004 = n17052 | n17053;
  assign n55005 = n17058 | n17059;
  assign n55006 = n17064 | n17065;
  assign n55007 = n17083 | n17084;
  assign n55008 = n17097 | n17094 | n17096;
  assign n55009 = n17100 | ~n17101;
  assign n55010 = n17108 | n17109;
  assign n55011 = n17110 | n17111;
  assign n55012 = n17112 | ~n17113;
  assign n55013 = n17117 | n17118;
  assign n55014 = n17119 | n17120;
  assign n55015 = n17121 | ~n17122;
  assign n55016 = n17135 | n17136;
  assign n55017 = n17139 | n17140;
  assign n55018 = n17141 | n17142;
  assign n55019 = n17147 | n17148;
  assign n55020 = n17157 | n17158;
  assign n55021 = n17161 | n17162;
  assign n55022 = n17163 | n17164;
  assign n55023 = n17169 | n17170;
  assign n55024 = n17173 | n17174;
  assign n55025 = n17175 | n17176;
  assign n55026 = n17178 | ~n17179;
  assign n55027 = n17188 | n17189;
  assign n55028 = n17192 | n17193;
  assign n55029 = n17194 | n17195;
  assign n55030 = n17200 | n17201;
  assign n55031 = n17210 | n17211;
  assign n55032 = n17214 | n17215;
  assign n55033 = n17216 | n17217;
  assign n55034 = n17222 | n17223;
  assign n55035 = n17231 | n17232;
  assign n55036 = n17233 | n17234;
  assign n55037 = n17236 | ~n17237;
  assign n55038 = n17247 | ~n17248;
  assign n55039 = n17253 | ~n17254;
  assign n55040 = n17260 | ~n17261;
  assign n55041 = n17263 | n17264;
  assign n55042 = n17271 | n17272;
  assign n55043 = n17284 | n17285;
  assign n55044 = n17288 | ~n17289;
  assign n55045 = n17299 | ~n17300;
  assign n55046 = n17309 | n17310;
  assign n55047 = n17313 | ~n17314;
  assign n55048 = n17327 | n17328;
  assign n55049 = n17331 | ~n17332;
  assign n55050 = n17339 | ~n17340;
  assign n55051 = n17349 | n17350;
  assign n55052 = n17353 | n17354;
  assign n55053 = n17355 | n17356;
  assign n55054 = n17361 | n17362;
  assign n55055 = n17368 | ~n17369;
  assign n55056 = n17378 | n17379;
  assign n55057 = n17382 | n17383;
  assign n55058 = n17384 | n17385;
  assign n55059 = n17390 | n17391;
  assign n55060 = n17400 | n17401;
  assign n55061 = n17404 | n17405;
  assign n55062 = n17406 | n17407;
  assign n55063 = n17412 | n17413;
  assign n55064 = n17419 | ~n17420;
  assign n55065 = n17431 | n17432;
  assign n55066 = n17433 | n17434;
  assign n55067 = n17439 | n17440;
  assign n55068 = n17446 | ~n17447;
  assign n55069 = n17451 | n17452;
  assign n55070 = n17462 | n17463;
  assign n55071 = n17466 | n17467;
  assign n55072 = n17468 | n17469;
  assign n55073 = n17475 | n17476;
  assign n55074 = n17477 | n17478;
  assign n55075 = n17479 | ~n17480;
  assign n55076 = n17484 | ~n17485;
  assign n55077 = n17492 | n17493;
  assign n55078 = n17496 | n17497;
  assign n55079 = n17498 | n17499;
  assign n55080 = n17505 | n17506;
  assign n55081 = n17507 | n17508;
  assign n55082 = n17509 | ~n17510;
  assign n55083 = n17514 | ~n17515;
  assign n55084 = n17521 | ~n17522;
  assign n55085 = n17531 | n17532;
  assign n55086 = n17535 | n17536;
  assign n55087 = n17541 | ~n17542;
  assign n55088 = n17553 | n17554;
  assign n55089 = n17558 | n17559;
  assign n55090 = n17563 | n17564;
  assign n55091 = n17567 | n17568;
  assign n55092 = n17578 | n17579;
  assign n55093 = n17588 | n17589;
  assign n55094 = n17590 | n17591;
  assign n55095 = n17593 | n17594;
  assign n55096 = n17600 | n17601;
  assign n55097 = n17604 | n17605;
  assign n55098 = n17615 | n17616;
  assign n55099 = n17627 | n17628;
  assign n55100 = n17639 | n17640;
  assign n55101 = n17657 | n17658;
  assign n55102 = n17667 | n17668;
  assign n55103 = n17671 | n17672;
  assign n55104 = n17684 | n17679 | n17683;
  assign n55105 = n17696 | n17697;
  assign n55106 = n17702 | n17703;
  assign n55107 = n17727 | n17716 | n17726;
  assign n55108 = n17733 | n17734;
  assign n55109 = n17770 | n17752 | n17761 | n17780 | n17781;
  assign n55110 = n17801 | n17802;
  assign n55111 = n17813 | n17814;
  assign n55112 = n17820 | n17821;
  assign n55113 = n17833 | n17834;
  assign n55114 = n17842 | n17843;
  assign n55115 = n17861 | n17852 | n17860;
  assign n55116 = n17867 | n17868;
  assign n55117 = n17884 | n17880 | n17883;
  assign n55118 = n17901 | n17910 | n17921 | n17922;
  assign n55119 = n17936 | n17937;
  assign n55120 = n17948 | n17949;
  assign n55121 = n17955 | n17956;
  assign n55122 = n17970 | n17964 | n17969;
  assign n55123 = n17982 | n17983;
  assign n55124 = n17988 | n17989;
  assign n55125 = n17993 | n17994;
  assign n55126 = n18001 | n18002;
  assign n55127 = n18010 | n18011;
  assign n55128 = n18018 | n18019;
  assign n55129 = n18033 | n18034;
  assign n55130 = n18053 | n18054;
  assign n55131 = n18065 | n18066;
  assign n55132 = n18080 | n18086 | n18093 | n18094;
  assign n55133 = n18099 | n18100;
  assign n55134 = n18108 | n18109;
  assign n55135 = n18126 | n18127;
  assign n55136 = n18150 | n18151;
  assign n55137 = n18154 | n18155;
  assign n55138 = n18165 | n18166;
  assign n55139 = n18176 | n18182 | n18187 | n18188;
  assign n55140 = n18196 | n18197;
  assign n55141 = n18209 | n18200 | n18204 | n18212 | n18213;
  assign n55142 = n18218 | n18215 | n18217;
  assign n55143 = n18221 | n18222;
  assign n55144 = n18226 | n18227;
  assign n55145 = n18231 | n18232;
  assign n55146 = n18241 | n18237 | n18240;
  assign n55147 = n18249 | n18250;
  assign n55148 = n18257 | n18258;
  assign n55149 = n18269 | n18270;
  assign n55150 = n18300 | n18287 | n18299;
  assign n55151 = n18315 | n18316;
  assign n55152 = n18331 | n18332;
  assign n55153 = n18343 | n18344;
  assign n55154 = n18349 | n18350;
  assign n55155 = n18352 | n18353;
  assign n55156 = n18354 | n18355;
  assign n55157 = n18356 | ~n18357;
  assign n55158 = n18361 | n18362;
  assign n55159 = n18363 | n18364;
  assign n55160 = n18365 | ~n18366;
  assign n55161 = n18370 | n18371;
  assign n55162 = n18372 | n18373;
  assign n55163 = n18374 | ~n18375;
  assign n55164 = n18379 | n18380;
  assign n55165 = n18381 | n18382;
  assign n55166 = n18383 | ~n18384;
  assign n55167 = n18390 | ~n18391;
  assign n55168 = n18403 | ~n18404;
  assign n55169 = n18411 | n18412;
  assign n55170 = n18413 | n18414;
  assign n55171 = n18415 | ~n18416;
  assign n55172 = n18420 | n18421;
  assign n55173 = n18422 | n18423;
  assign n55174 = n18424 | ~n18425;
  assign n55175 = n18431 | ~n18432;
  assign n55176 = n18441 | n18442;
  assign n55177 = n18445 | n18446;
  assign n55178 = n18447 | n18448;
  assign n55179 = n18453 | n18454;
  assign n55180 = n18463 | n18464;
  assign n55181 = n18467 | n18468;
  assign n55182 = n18469 | n18470;
  assign n55183 = n18475 | n18476;
  assign n55184 = n18485 | n18486;
  assign n55185 = n18489 | n18490;
  assign n55186 = n18491 | n18492;
  assign n55187 = n18497 | n18498;
  assign n55188 = n18501 | n18502;
  assign n55189 = n18503 | n18504;
  assign n55190 = n18506 | ~n18507;
  assign n55191 = n18516 | n18517;
  assign n55192 = n18520 | n18521;
  assign n55193 = n18522 | n18523;
  assign n55194 = n18528 | n18529;
  assign n55195 = n18538 | n18539;
  assign n55196 = n18542 | n18543;
  assign n55197 = n18544 | n18545;
  assign n55198 = n18550 | n18551;
  assign n55199 = n18561 | ~n18562;
  assign n55200 = n18569 | n18570;
  assign n55201 = n18571 | n18572;
  assign n55202 = n18574 | ~n18575;
  assign n55203 = n18581 | ~n18582;
  assign n55204 = n18593 | n18594;
  assign n55205 = n18597 | ~n18598;
  assign n55206 = n18605 | ~n18606;
  assign n55207 = n18615 | n18616;
  assign n55208 = n18619 | ~n18620;
  assign n55209 = n18630 | ~n18631;
  assign n55210 = n18638 | n18639;
  assign n55211 = n18642 | ~n18643;
  assign n55212 = n18647 | n18648;
  assign n55213 = n18649 | n18650;
  assign n55214 = n18652 | ~n18653;
  assign n55215 = n18663 | n18664;
  assign n55216 = n18667 | ~n18668;
  assign n55217 = n18675 | ~n18676;
  assign n55218 = n18685 | n18686;
  assign n55219 = n18689 | n18690;
  assign n55220 = n18691 | n18692;
  assign n55221 = n18697 | n18698;
  assign n55222 = n18704 | ~n18705;
  assign n55223 = n18714 | n18715;
  assign n55224 = n18718 | n18719;
  assign n55225 = n18720 | n18721;
  assign n55226 = n18726 | n18727;
  assign n55227 = n18736 | n18737;
  assign n55228 = n18740 | n18741;
  assign n55229 = n18742 | n18743;
  assign n55230 = n18748 | n18749;
  assign n55231 = n18755 | ~n18756;
  assign n55232 = n18765 | n18766;
  assign n55233 = n18769 | n18770;
  assign n55234 = n18771 | n18772;
  assign n55235 = n18777 | n18778;
  assign n55236 = n18787 | n18788;
  assign n55237 = n18791 | n18792;
  assign n55238 = n18793 | n18794;
  assign n55239 = n18799 | n18800;
  assign n55240 = n18805 | n18806;
  assign n55241 = n18807 | n18808;
  assign n55242 = n18809 | ~n18810;
  assign n55243 = n18820 | n18817 | n18819;
  assign n55244 = n18826 | ~n18827;
  assign n55245 = n18832 | ~n18833;
  assign n55246 = n18839 | ~n18840;
  assign n55247 = n18845 | n18842 | n18844;
  assign n55248 = n18852 | n18853;
  assign n55249 = n18863 | n18864;
  assign n55250 = n18867 | n18868;
  assign n55251 = n18869 | n18870;
  assign n55252 = n18876 | n18877;
  assign n55253 = n18878 | n18879;
  assign n55254 = n18880 | ~n18881;
  assign n55255 = n18885 | ~n18886;
  assign n55256 = n18893 | n18894;
  assign n55257 = n18897 | n18898;
  assign n55258 = n18899 | n18900;
  assign n55259 = n18906 | n18907;
  assign n55260 = n18908 | n18909;
  assign n55261 = n18910 | ~n18911;
  assign n55262 = n18915 | ~n18916;
  assign n55263 = n18923 | n18924;
  assign n55264 = n18927 | ~n18928;
  assign n55265 = n18935 | ~n18936;
  assign n55266 = n18948 | n18945 | n18947;
  assign n55267 = n18951 | n18952;
  assign n55268 = n18953 | n18954;
  assign n55269 = n18959 | n18960;
  assign n55270 = n18969 | n18970;
  assign n55271 = n18973 | n18974;
  assign n55272 = n18975 | n18976;
  assign n55273 = n18981 | n18982;
  assign n55274 = n18985 | n18986;
  assign n55275 = n18987 | n18988;
  assign n55276 = n18990 | ~n18991;
  assign n55277 = n19000 | n19001;
  assign n55278 = n19004 | n19005;
  assign n55279 = n19006 | n19007;
  assign n55280 = n19012 | n19013;
  assign n55281 = n19022 | n19023;
  assign n55282 = n19026 | n19027;
  assign n55283 = n19028 | n19029;
  assign n55284 = n19034 | n19035;
  assign n55285 = n19038 | n19039;
  assign n55286 = n19040 | n19041;
  assign n55287 = n19043 | ~n19044;
  assign n55288 = n19055 | n19056;
  assign n55289 = n19057 | n19058;
  assign n55290 = n19063 | n19064;
  assign n55291 = n19070 | ~n19071;
  assign n55292 = n19075 | n19076;
  assign n55293 = n19086 | n19087;
  assign n55294 = n19090 | ~n19091;
  assign n55295 = n19097 | n19098;
  assign n55296 = n19099 | n19100;
  assign n55297 = n19101 | ~n19102;
  assign n55298 = n19106 | ~n19107;
  assign n55299 = n19116 | n19117;
  assign n55300 = n19120 | ~n19121;
  assign n55301 = n19131 | ~n19132;
  assign n55302 = n19139 | n19140;
  assign n55303 = n19143 | ~n19144;
  assign n55304 = n19151 | ~n19152;
  assign n55305 = n19160 | n19161;
  assign n55306 = n19164 | ~n19165;
  assign n55307 = n19172 | ~n19173;
  assign n55308 = n19181 | n19182;
  assign n55309 = n19185 | n19186;
  assign n55310 = n19187 | n19188;
  assign n55311 = n19193 | ~n19194;
  assign n55312 = n19202 | n19203;
  assign n55313 = n19206 | n19207;
  assign n55314 = n19208 | n19209;
  assign n55315 = n19214 | ~n19215;
  assign n55316 = n19223 | n19224;
  assign n55317 = n19227 | n19228;
  assign n55318 = n19229 | n19230;
  assign n55319 = n19235 | ~n19236;
  assign n55320 = n19246 | n19247;
  assign n55321 = n19248 | n19249;
  assign n55322 = n19252 | n19253;
  assign n55323 = n19254 | n19255;
  assign n55324 = n19256 | ~n19257;
  assign n55325 = n19265 | n19266;
  assign n55326 = n19269 | n19270;
  assign n55327 = n19271 | n19272;
  assign n55328 = n19294 | n19295;
  assign n55329 = n19304 | ~n19305;
  assign n55330 = n19309 | n19310;
  assign n55331 = n19318 | n19319;
  assign n55332 = n19322 | n19323;
  assign n55333 = n19324 | n19325;
  assign n55334 = n19330 | ~n19331;
  assign n55335 = n19335 | n19336;
  assign n55336 = n19337 | n19338;
  assign n55337 = n19339 | ~n19340;
  assign n55338 = n19346 | ~n19347;
  assign n55339 = n19353 | ~n19354;
  assign n55340 = n19358 | n19359;
  assign n55341 = n19360 | n19361;
  assign n55342 = n19362 | ~n19363;
  assign n55343 = n19367 | n19368;
  assign n55344 = n19369 | n19370;
  assign n55345 = n19371 | ~n19372;
  assign n55346 = n19392 | n19393;
  assign n55347 = n19396 | n19397;
  assign n55348 = n19398 | n19399;
  assign n55349 = n19408 | ~n19409;
  assign n55350 = n19418 | n19419;
  assign n55351 = n19422 | n19423;
  assign n55352 = n19424 | n19425;
  assign n55353 = n19430 | n19431;
  assign n55354 = n19440 | n19441;
  assign n55355 = n19444 | n19445;
  assign n55356 = n19446 | n19447;
  assign n55357 = n19452 | n19453;
  assign n55358 = n19459 | ~n19460;
  assign n55359 = n19469 | n19470;
  assign n55360 = n19473 | n19474;
  assign n55361 = n19475 | n19476;
  assign n55362 = n19481 | n19482;
  assign n55363 = n19491 | n19492;
  assign n55364 = n19495 | n19496;
  assign n55365 = n19497 | n19498;
  assign n55366 = n19503 | n19504;
  assign n55367 = n19514 | ~n19515;
  assign n55368 = n19525 | ~n19526;
  assign n55369 = n19532 | ~n19533;
  assign n55370 = n19546 | n19547;
  assign n55371 = n19550 | ~n19551;
  assign n55372 = n19558 | ~n19559;
  assign n55373 = n19566 | n19567;
  assign n55374 = n19570 | n19571;
  assign n55375 = n19572 | n19573;
  assign n55376 = n19579 | n19580;
  assign n55377 = n19581 | n19582;
  assign n55378 = n19583 | ~n19584;
  assign n55379 = n19588 | ~n19589;
  assign n55380 = n19598 | n19599;
  assign n55381 = n19602 | ~n19603;
  assign n55382 = n19616 | n19617;
  assign n55383 = n19620 | ~n19621;
  assign n55384 = n19636 | ~n19637;
  assign n55385 = n19650 | n19651;
  assign n55386 = n19654 | ~n19655;
  assign n55387 = n19668 | n19669;
  assign n55388 = n19672 | ~n19673;
  assign n55389 = n19686 | n19687;
  assign n55390 = n19690 | ~n19691;
  assign n55391 = n19702 | n19703;
  assign n55392 = n19706 | ~n19707;
  assign n55393 = n19714 | ~n19715;
  assign n55394 = n19723 | n19724;
  assign n55395 = n19727 | n19728;
  assign n55396 = n19729 | n19730;
  assign n55397 = n19743 | n19744;
  assign n55398 = n19745 | n19746;
  assign n55399 = n19752 | n19753;
  assign n55400 = n19761 | n19762;
  assign n55401 = n19765 | ~n19766;
  assign n55402 = n19774 | n19775;
  assign n55403 = n19788 | n19789;
  assign n55404 = n19798 | ~n19799;
  assign n55405 = n19803 | n19804;
  assign n55406 = n19812 | n19813;
  assign n55407 = n19816 | n19817;
  assign n55408 = n19818 | n19819;
  assign n55409 = n19822 | n19823;
  assign n55410 = n19824 | n19825;
  assign n55411 = n19826 | ~n19827;
  assign n55412 = n19835 | n19836;
  assign n55413 = n19837 | n19838;
  assign n55414 = n19839 | ~n19840;
  assign n55415 = n19844 | n19845;
  assign n55416 = n19846 | n19847;
  assign n55417 = n19848 | ~n19849;
  assign n55418 = n19853 | n19854;
  assign n55419 = n19855 | n19856;
  assign n55420 = n19857 | ~n19858;
  assign n55421 = n19862 | n19863;
  assign n55422 = n19864 | n19865;
  assign n55423 = n19866 | ~n19867;
  assign n55424 = n19871 | n19872;
  assign n55425 = n19873 | n19874;
  assign n55426 = n19875 | ~n19876;
  assign n55427 = n19880 | n19881;
  assign n55428 = n19882 | n19883;
  assign n55429 = n19884 | ~n19885;
  assign n55430 = n19889 | n19890;
  assign n55431 = n19891 | n19892;
  assign n55432 = n19893 | ~n19894;
  assign n55433 = n19898 | n19899;
  assign n55434 = n19900 | n19901;
  assign n55435 = n19902 | ~n19903;
  assign n55436 = n19907 | n19908;
  assign n55437 = n19909 | n19910;
  assign n55438 = n19911 | ~n19912;
  assign n55439 = n19924 | n19925;
  assign n55440 = n19928 | n19929;
  assign n55441 = n19930 | n19931;
  assign n55442 = n19937 | n19938;
  assign n55443 = n19939 | n19940;
  assign n55444 = n19942 | ~n19943;
  assign n55445 = n19952 | n19953;
  assign n55446 = n19956 | n19957;
  assign n55447 = n19958 | n19959;
  assign n55448 = n19964 | n19965;
  assign n55449 = n19974 | n19975;
  assign n55450 = n19978 | n19979;
  assign n55451 = n19980 | n19981;
  assign n55452 = n19986 | n19987;
  assign n55453 = n19990 | n19991;
  assign n55454 = n19992 | n19993;
  assign n55455 = n19995 | ~n19996;
  assign n55456 = n20005 | n20006;
  assign n55457 = n20009 | n20010;
  assign n55458 = n20011 | n20012;
  assign n55459 = n20017 | n20018;
  assign n55460 = n20027 | n20028;
  assign n55461 = n20031 | n20032;
  assign n55462 = n20033 | n20034;
  assign n55463 = n20039 | n20040;
  assign n55464 = n20044 | n20045;
  assign n55465 = n20046 | n20047;
  assign n55466 = n20048 | ~n20049;
  assign n55467 = n20053 | n20054;
  assign n55468 = n20059 | ~n20060;
  assign n55469 = n20065 | ~n20066;
  assign n55470 = n20071 | ~n20072;
  assign n55471 = n20078 | ~n20079;
  assign n55472 = n20084 | n20081 | n20083;
  assign n55473 = n20091 | n20092;
  assign n55474 = n20104 | n20105;
  assign n55475 = n20108 | ~n20109;
  assign n55476 = n20119 | ~n20120;
  assign n55477 = n20127 | n20128;
  assign n55478 = n20131 | n20132;
  assign n55479 = n20133 | n20134;
  assign n55480 = n20139 | ~n20140;
  assign n55481 = n20151 | n20148 | n20150;
  assign n55482 = n20154 | n20155;
  assign n55483 = n20156 | n20157;
  assign n55484 = n20162 | ~n20163;
  assign n55485 = n20171 | n20172;
  assign n55486 = n20175 | n20176;
  assign n55487 = n20177 | n20178;
  assign n55488 = n20181 | n20182;
  assign n55489 = n20183 | n20184;
  assign n55490 = n20185 | ~n20186;
  assign n55491 = n20194 | n20195;
  assign n55492 = n20198 | n20199;
  assign n55493 = n20200 | n20201;
  assign n55494 = n20204 | n20205;
  assign n55495 = n20206 | n20207;
  assign n55496 = n20208 | ~n20209;
  assign n55497 = n20217 | n20218;
  assign n55498 = n20221 | n20222;
  assign n55499 = n20223 | n20224;
  assign n55500 = n20229 | ~n20230;
  assign n55501 = n20240 | n20241;
  assign n55502 = n20242 | n20243;
  assign n55503 = n20248 | ~n20249;
  assign n55504 = n20257 | n20258;
  assign n55505 = n20261 | n20262;
  assign n55506 = n20263 | n20264;
  assign n55507 = n20267 | n20268;
  assign n55508 = n20269 | n20270;
  assign n55509 = n20271 | ~n20272;
  assign n55510 = n20282 | n20283;
  assign n55511 = n20286 | ~n20287;
  assign n55512 = n20300 | n20301;
  assign n55513 = n20304 | ~n20305;
  assign n55514 = n20316 | n20317;
  assign n55515 = n20320 | n20321;
  assign n55516 = n20322 | n20323;
  assign n55517 = n20334 | n20335;
  assign n55518 = n20338 | ~n20339;
  assign n55519 = n20346 | ~n20347;
  assign n55520 = n20357 | n20358;
  assign n55521 = n20359 | n20360;
  assign n55522 = n20366 | n20367;
  assign n55523 = n20375 | n20376;
  assign n55524 = n20379 | ~n20380;
  assign n55525 = n20388 | n20389;
  assign n55526 = n20402 | n20403;
  assign n55527 = n20412 | ~n20413;
  assign n55528 = n20417 | n20418;
  assign n55529 = n20426 | n20427;
  assign n55530 = n20430 | n20431;
  assign n55531 = n20432 | n20433;
  assign n55532 = n20436 | n20437;
  assign n55533 = n20438 | n20439;
  assign n55534 = n20440 | ~n20441;
  assign n55535 = n20449 | n20450;
  assign n55536 = n20451 | n20452;
  assign n55537 = n20453 | ~n20454;
  assign n55538 = n20462 | n20463;
  assign n55539 = n20464 | n20465;
  assign n55540 = n20466 | ~n20467;
  assign n55541 = n20471 | n20472;
  assign n55542 = n20473 | n20474;
  assign n55543 = n20475 | ~n20476;
  assign n55544 = n20486 | ~n20487;
  assign n55545 = n20491 | n20492;
  assign n55546 = n20493 | n20494;
  assign n55547 = n20495 | ~n20496;
  assign n55548 = n20500 | n20501;
  assign n55549 = n20502 | n20503;
  assign n55550 = n20504 | ~n20505;
  assign n55551 = n20511 | ~n20512;
  assign n55552 = n20518 | ~n20519;
  assign n55553 = n20523 | n20524;
  assign n55554 = n20525 | n20526;
  assign n55555 = n20527 | ~n20528;
  assign n55556 = n20532 | n20533;
  assign n55557 = n20534 | n20535;
  assign n55558 = n20536 | ~n20537;
  assign n55559 = n20549 | n20550;
  assign n55560 = n20553 | n20554;
  assign n55561 = n20555 | n20556;
  assign n55562 = n20565 | ~n20566;
  assign n55563 = n20575 | n20576;
  assign n55564 = n20579 | n20580;
  assign n55565 = n20581 | n20582;
  assign n55566 = n20587 | n20588;
  assign n55567 = n20597 | n20598;
  assign n55568 = n20601 | n20602;
  assign n55569 = n20603 | n20604;
  assign n55570 = n20609 | n20610;
  assign n55571 = n20616 | ~n20617;
  assign n55572 = n20628 | n20629;
  assign n55573 = n20630 | n20631;
  assign n55574 = n20636 | n20637;
  assign n55575 = n20643 | ~n20644;
  assign n55576 = n20648 | n20649;
  assign n55577 = n20659 | n20660;
  assign n55578 = n20663 | ~n20664;
  assign n55579 = n20671 | ~n20672;
  assign n55580 = n20681 | n20682;
  assign n55581 = n20685 | ~n20686;
  assign n55582 = n20699 | n20700;
  assign n55583 = n20703 | ~n20704;
  assign n55584 = n20717 | n20718;
  assign n55585 = n20721 | ~n20722;
  assign n55586 = n20735 | n20736;
  assign n55587 = n20739 | ~n20740;
  assign n55588 = n20756 | n20753 | n20755;
  assign n55589 = n20759 | ~n20760;
  assign n55590 = n20773 | n20774;
  assign n55591 = n20777 | ~n20778;
  assign n55592 = n20791 | n20792;
  assign n55593 = n20795 | ~n20796;
  assign n55594 = n20807 | n20808;
  assign n55595 = n20811 | n20812;
  assign n55596 = n20813 | n20814;
  assign n55597 = n20827 | n20828;
  assign n55598 = n20829 | n20830;
  assign n55599 = n20833 | n20834;
  assign n55600 = n20835 | n20836;
  assign n55601 = n20837 | ~n20838;
  assign n55602 = n20848 | n20849;
  assign n55603 = n20852 | ~n20853;
  assign n55604 = n20866 | n20867;
  assign n55605 = n20870 | ~n20871;
  assign n55606 = n20884 | n20885;
  assign n55607 = n20888 | ~n20889;
  assign n55608 = n20900 | n20901;
  assign n55609 = n20904 | n20905;
  assign n55610 = n20906 | n20907;
  assign n55611 = n20918 | n20919;
  assign n55612 = n20922 | ~n20923;
  assign n55613 = n20930 | ~n20931;
  assign n55614 = n20941 | n20942;
  assign n55615 = n20943 | n20944;
  assign n55616 = n20950 | n20951;
  assign n55617 = n20959 | n20960;
  assign n55618 = n20963 | ~n20964;
  assign n55619 = n20972 | n20973;
  assign n55620 = n20986 | n20987;
  assign n55621 = n20996 | ~n20997;
  assign n55622 = n21001 | n21002;
  assign n55623 = n21010 | n21011;
  assign n55624 = n21014 | n21015;
  assign n55625 = n21016 | n21017;
  assign n55626 = n21020 | n21021;
  assign n55627 = n21022 | n21023;
  assign n55628 = n21024 | ~n21025;
  assign n55629 = n21033 | n21034;
  assign n55630 = n21035 | n21036;
  assign n55631 = n21037 | ~n21038;
  assign n55632 = n21046 | n21047;
  assign n55633 = n21048 | n21049;
  assign n55634 = n21050 | ~n21051;
  assign n55635 = n21055 | n21056;
  assign n55636 = n21057 | n21058;
  assign n55637 = n21059 | ~n21060;
  assign n55638 = n21064 | n21065;
  assign n55639 = n21066 | n21067;
  assign n55640 = n21068 | ~n21069;
  assign n55641 = n21079 | ~n21080;
  assign n55642 = n21084 | n21085;
  assign n55643 = n21086 | n21087;
  assign n55644 = n21088 | ~n21089;
  assign n55645 = n21093 | n21094;
  assign n55646 = n21095 | n21096;
  assign n55647 = n21097 | ~n21098;
  assign n55648 = n21102 | n21103;
  assign n55649 = n21104 | n21105;
  assign n55650 = n21106 | ~n21107;
  assign n55651 = n21111 | n21112;
  assign n55652 = n21113 | n21114;
  assign n55653 = n21115 | ~n21116;
  assign n55654 = n21120 | n21121;
  assign n55655 = n21122 | n21123;
  assign n55656 = n21124 | ~n21125;
  assign n55657 = n21129 | n21130;
  assign n55658 = n21131 | n21132;
  assign n55659 = n21133 | ~n21134;
  assign n55660 = n21138 | n21139;
  assign n55661 = n21140 | n21141;
  assign n55662 = n21142 | ~n21143;
  assign n55663 = n21147 | n21148;
  assign n55664 = n21149 | n21150;
  assign n55665 = n21151 | ~n21152;
  assign n55666 = n21164 | n21165;
  assign n55667 = n21168 | n21169;
  assign n55668 = n21170 | n21171;
  assign n55669 = n21177 | n21178;
  assign n55670 = n21179 | n21180;
  assign n55671 = n21182 | ~n21183;
  assign n55672 = n21192 | n21193;
  assign n55673 = n21196 | n21197;
  assign n55674 = n21198 | n21199;
  assign n55675 = n21204 | n21205;
  assign n55676 = n21214 | n21215;
  assign n55677 = n21218 | n21219;
  assign n55678 = n21220 | n21221;
  assign n55679 = n21226 | n21227;
  assign n55680 = n21242 | ~n21243;
  assign n55681 = n21250 | n21251;
  assign n55682 = n21252 | n21253;
  assign n55683 = n21255 | ~n21256;
  assign n55684 = n21262 | ~n21263;
  assign n55685 = n21274 | n21275;
  assign n55686 = n21278 | ~n21279;
  assign n55687 = n21286 | ~n21287;
  assign n55688 = n21294 | n21295;
  assign n55689 = n21298 | n21299;
  assign n55690 = n21300 | n21301;
  assign n55691 = n21304 | n21305;
  assign n55692 = n21306 | n21307;
  assign n55693 = n21308 | ~n21309;
  assign n55694 = n21317 | n21318;
  assign n55695 = n21321 | n21322;
  assign n55696 = n21323 | n21324;
  assign n55697 = n21327 | n21328;
  assign n55698 = n21329 | n21330;
  assign n55699 = n21331 | ~n21332;
  assign n55700 = n21340 | n21341;
  assign n55701 = n21344 | n21345;
  assign n55702 = n21346 | n21347;
  assign n55703 = n21352 | ~n21353;
  assign n55704 = n21361 | n21362;
  assign n55705 = n21365 | n21366;
  assign n55706 = n21367 | n21368;
  assign n55707 = n21373 | ~n21374;
  assign n55708 = n21382 | n21383;
  assign n55709 = n21386 | n21387;
  assign n55710 = n21388 | n21389;
  assign n55711 = n21392 | n21393;
  assign n55712 = n21394 | n21395;
  assign n55713 = n21396 | ~n21397;
  assign n55714 = n21405 | n21406;
  assign n55715 = n21409 | n21410;
  assign n55716 = n21411 | n21412;
  assign n55717 = n21415 | n21416;
  assign n55718 = n21417 | n21418;
  assign n55719 = n21419 | ~n21420;
  assign n55720 = n21428 | n21429;
  assign n55721 = n21432 | n21433;
  assign n55722 = n21434 | n21435;
  assign n55723 = n21440 | ~n21441;
  assign n55724 = n21454 | n21451 | n21453;
  assign n55725 = n21457 | ~n21458;
  assign n55726 = n21471 | n21472;
  assign n55727 = n21475 | ~n21476;
  assign n55728 = n21487 | n21488;
  assign n55729 = n21491 | n21492;
  assign n55730 = n21493 | n21494;
  assign n55731 = n21505 | n21506;
  assign n55732 = n21509 | n21510;
  assign n55733 = n21511 | n21512;
  assign n55734 = n21517 | ~n21518;
  assign n55735 = n21528 | n21529;
  assign n55736 = n21530 | n21531;
  assign n55737 = n21534 | n21535;
  assign n55738 = n21536 | n21537;
  assign n55739 = n21538 | ~n21539;
  assign n55740 = n21549 | n21550;
  assign n55741 = n21553 | ~n21554;
  assign n55742 = n21567 | n21568;
  assign n55743 = n21571 | ~n21572;
  assign n55744 = n21585 | n21586;
  assign n55745 = n21589 | ~n21590;
  assign n55746 = n21601 | n21602;
  assign n55747 = n21605 | n21606;
  assign n55748 = n21607 | n21608;
  assign n55749 = n21619 | n21620;
  assign n55750 = n21623 | ~n21624;
  assign n55751 = n21631 | ~n21632;
  assign n55752 = n21642 | n21643;
  assign n55753 = n21644 | n21645;
  assign n55754 = n21651 | n21652;
  assign n55755 = n21660 | n21661;
  assign n55756 = n21664 | ~n21665;
  assign n55757 = n21673 | n21674;
  assign n55758 = n21687 | n21688;
  assign n55759 = n21697 | ~n21698;
  assign n55760 = n21702 | n21703;
  assign n55761 = n21711 | n21712;
  assign n55762 = n21715 | n21716;
  assign n55763 = n21717 | n21718;
  assign n55764 = n21721 | n21722;
  assign n55765 = n21723 | n21724;
  assign n55766 = n21725 | ~n21726;
  assign n55767 = n21734 | n21735;
  assign n55768 = n21736 | n21737;
  assign n55769 = n21738 | ~n21739;
  assign n55770 = n21747 | n21748;
  assign n55771 = n21749 | n21750;
  assign n55772 = n21751 | ~n21752;
  assign n55773 = n21756 | n21757;
  assign n55774 = n21758 | n21759;
  assign n55775 = n21760 | ~n21761;
  assign n55776 = n21765 | n21766;
  assign n55777 = n21767 | n21768;
  assign n55778 = n21769 | ~n21770;
  assign n55779 = n21780 | ~n21781;
  assign n55780 = n21785 | n21786;
  assign n55781 = n21787 | n21788;
  assign n55782 = n21789 | ~n21790;
  assign n55783 = n21794 | n21795;
  assign n55784 = n21796 | n21797;
  assign n55785 = n21798 | ~n21799;
  assign n55786 = n21803 | n21804;
  assign n55787 = n21805 | n21806;
  assign n55788 = n21807 | ~n21808;
  assign n55789 = n21816 | n21817;
  assign n55790 = n21818 | n21819;
  assign n55791 = n21820 | ~n21821;
  assign n55792 = n21827 | ~n21828;
  assign n55793 = n21834 | ~n21835;
  assign n55794 = n21839 | n21840;
  assign n55795 = n21841 | n21842;
  assign n55796 = n21843 | ~n21844;
  assign n55797 = n21848 | n21849;
  assign n55798 = n21850 | n21851;
  assign n55799 = n21852 | ~n21853;
  assign n55800 = n21859 | ~n21860;
  assign n55801 = n21866 | ~n21867;
  assign n55802 = n21879 | n21880;
  assign n55803 = n21883 | n21884;
  assign n55804 = n21885 | n21886;
  assign n55805 = n21895 | ~n21896;
  assign n55806 = n21905 | n21906;
  assign n55807 = n21909 | n21910;
  assign n55808 = n21911 | n21912;
  assign n55809 = n21917 | n21918;
  assign n55810 = n21927 | n21928;
  assign n55811 = n21931 | n21932;
  assign n55812 = n21933 | n21934;
  assign n55813 = n21939 | n21940;
  assign n55814 = n21945 | n21946;
  assign n55815 = n21947 | n21948;
  assign n55816 = n21949 | ~n21950;
  assign n55817 = n21960 | n21957 | n21959;
  assign n55818 = n21967 | ~n21968;
  assign n55819 = n21975 | n21976;
  assign n55820 = n21988 | n21989;
  assign n55821 = n21992 | ~n21993;
  assign n55822 = n22006 | n22007;
  assign n55823 = n22010 | ~n22011;
  assign n55824 = n22024 | n22025;
  assign n55825 = n22028 | ~n22029;
  assign n55826 = n22042 | n22043;
  assign n55827 = n22046 | ~n22047;
  assign n55828 = n22060 | n22061;
  assign n55829 = n22064 | ~n22065;
  assign n55830 = n22078 | n22079;
  assign n55831 = n22082 | ~n22083;
  assign n55832 = n22096 | n22097;
  assign n55833 = n22100 | ~n22101;
  assign n55834 = n22112 | n22113;
  assign n55835 = n22116 | n22117;
  assign n55836 = n22118 | n22119;
  assign n55837 = n22130 | n22131;
  assign n55838 = n22134 | n22135;
  assign n55839 = n22136 | n22137;
  assign n55840 = n22142 | ~n22143;
  assign n55841 = n22153 | n22154;
  assign n55842 = n22157 | ~n22158;
  assign n55843 = n22174 | n22171 | n22173;
  assign n55844 = n22177 | ~n22178;
  assign n55845 = n22191 | n22192;
  assign n55846 = n22195 | ~n22196;
  assign n55847 = n22207 | n22208;
  assign n55848 = n22211 | n22212;
  assign n55849 = n22213 | n22214;
  assign n55850 = n22225 | n22226;
  assign n55851 = n22229 | n22230;
  assign n55852 = n22231 | n22232;
  assign n55853 = n22237 | ~n22238;
  assign n55854 = n22248 | n22249;
  assign n55855 = n22250 | n22251;
  assign n55856 = n22254 | n22255;
  assign n55857 = n22256 | n22257;
  assign n55858 = n22258 | ~n22259;
  assign n55859 = n22269 | n22270;
  assign n55860 = n22273 | ~n22274;
  assign n55861 = n22287 | n22288;
  assign n55862 = n22291 | ~n22292;
  assign n55863 = n22305 | n22306;
  assign n55864 = n22309 | ~n22310;
  assign n55865 = n22321 | n22322;
  assign n55866 = n22325 | n22326;
  assign n55867 = n22327 | n22328;
  assign n55868 = n22339 | n22340;
  assign n55869 = n22343 | ~n22344;
  assign n55870 = n22351 | ~n22352;
  assign n55871 = n22362 | n22363;
  assign n55872 = n22364 | n22365;
  assign n55873 = n22371 | n22372;
  assign n55874 = n22380 | n22381;
  assign n55875 = n22384 | ~n22385;
  assign n55876 = n22393 | n22394;
  assign n55877 = n22407 | n22408;
  assign n55878 = n22417 | ~n22418;
  assign n55879 = n22422 | n22423;
  assign n55880 = n22431 | n22432;
  assign n55881 = n22435 | n22436;
  assign n55882 = n22437 | n22438;
  assign n55883 = n22441 | n22442;
  assign n55884 = n22443 | n22444;
  assign n55885 = n22445 | ~n22446;
  assign n55886 = n22454 | n22455;
  assign n55887 = n22456 | n22457;
  assign n55888 = n22458 | ~n22459;
  assign n55889 = n22467 | n22468;
  assign n55890 = n22469 | n22470;
  assign n55891 = n22471 | ~n22472;
  assign n55892 = n22476 | n22477;
  assign n55893 = n22478 | n22479;
  assign n55894 = n22480 | ~n22481;
  assign n55895 = n22485 | n22486;
  assign n55896 = n22487 | n22488;
  assign n55897 = n22489 | ~n22490;
  assign n55898 = n22500 | ~n22501;
  assign n55899 = n22505 | n22506;
  assign n55900 = n22507 | n22508;
  assign n55901 = n22509 | ~n22510;
  assign n55902 = n22514 | n22515;
  assign n55903 = n22516 | n22517;
  assign n55904 = n22518 | ~n22519;
  assign n55905 = n22523 | n22524;
  assign n55906 = n22525 | n22526;
  assign n55907 = n22527 | ~n22528;
  assign n55908 = n22532 | n22533;
  assign n55909 = n22534 | n22535;
  assign n55910 = n22536 | ~n22537;
  assign n55911 = n22545 | n22546;
  assign n55912 = n22547 | n22548;
  assign n55913 = n22549 | ~n22550;
  assign n55914 = n22554 | n22555;
  assign n55915 = n22556 | n22557;
  assign n55916 = n22558 | ~n22559;
  assign n55917 = n22563 | n22564;
  assign n55918 = n22565 | n22566;
  assign n55919 = n22567 | ~n22568;
  assign n55920 = n22572 | n22573;
  assign n55921 = n22574 | n22575;
  assign n55922 = n22576 | ~n22577;
  assign n55923 = n22581 | n22582;
  assign n55924 = n22583 | n22584;
  assign n55925 = n22585 | ~n22586;
  assign n55926 = n22590 | n22591;
  assign n55927 = n22592 | n22593;
  assign n55928 = n22594 | ~n22595;
  assign n55929 = n22599 | n22600;
  assign n55930 = n22601 | n22602;
  assign n55931 = n22603 | ~n22604;
  assign n55932 = n22608 | n22609;
  assign n55933 = n22610 | n22611;
  assign n55934 = n22612 | ~n22613;
  assign n55935 = n22617 | n22618;
  assign n55936 = n22619 | n22620;
  assign n55937 = n22621 | ~n22622;
  assign n55938 = n22634 | n22635;
  assign n55939 = n22638 | n22639;
  assign n55940 = n22640 | n22641;
  assign n55941 = n22647 | n22648;
  assign n55942 = n22649 | n22650;
  assign n55943 = n22652 | ~n22653;
  assign n55944 = n22664 | n22665;
  assign n55945 = n22666 | n22667;
  assign n55946 = n22672 | n22673;
  assign n55947 = n22679 | ~n22680;
  assign n55948 = n22684 | n22685;
  assign n55949 = n22693 | n22694;
  assign n55950 = n22697 | n22698;
  assign n55951 = n22699 | n22700;
  assign n55952 = n22705 | ~n22706;
  assign n55953 = n22714 | n22715;
  assign n55954 = n22718 | n22719;
  assign n55955 = n22720 | n22721;
  assign n55956 = n22726 | ~n22727;
  assign n55957 = n22735 | n22736;
  assign n55958 = n22739 | n22740;
  assign n55959 = n22741 | n22742;
  assign n55960 = n22745 | n22746;
  assign n55961 = n22747 | n22748;
  assign n55962 = n22749 | ~n22750;
  assign n55963 = n22758 | n22759;
  assign n55964 = n22762 | n22763;
  assign n55965 = n22764 | n22765;
  assign n55966 = n22768 | n22769;
  assign n55967 = n22770 | n22771;
  assign n55968 = n22772 | ~n22773;
  assign n55969 = n22781 | n22782;
  assign n55970 = n22785 | n22786;
  assign n55971 = n22787 | n22788;
  assign n55972 = n22793 | ~n22794;
  assign n55973 = n22802 | n22803;
  assign n55974 = n22806 | n22807;
  assign n55975 = n22808 | n22809;
  assign n55976 = n22814 | ~n22815;
  assign n55977 = n22823 | n22824;
  assign n55978 = n22827 | n22828;
  assign n55979 = n22829 | n22830;
  assign n55980 = n22833 | n22834;
  assign n55981 = n22835 | n22836;
  assign n55982 = n22837 | ~n22838;
  assign n55983 = n22848 | n22849;
  assign n55984 = n22852 | ~n22853;
  assign n55985 = n22866 | n22867;
  assign n55986 = n22870 | ~n22871;
  assign n55987 = n22882 | n22883;
  assign n55988 = n22886 | n22887;
  assign n55989 = n22888 | n22889;
  assign n55990 = n22900 | n22901;
  assign n55991 = n22904 | n22905;
  assign n55992 = n22906 | n22907;
  assign n55993 = n22910 | n22911;
  assign n55994 = n22912 | n22913;
  assign n55995 = n22914 | ~n22915;
  assign n55996 = n22923 | n22924;
  assign n55997 = n22927 | n22928;
  assign n55998 = n22929 | n22930;
  assign n55999 = n22935 | ~n22936;
  assign n56000 = n22946 | n22947;
  assign n56001 = n22950 | ~n22951;
  assign n56002 = n22967 | n22964 | n22966;
  assign n56003 = n22970 | ~n22971;
  assign n56004 = n22984 | n22985;
  assign n56005 = n22988 | ~n22989;
  assign n56006 = n23000 | n23001;
  assign n56007 = n23004 | n23005;
  assign n56008 = n23006 | n23007;
  assign n56009 = n23018 | n23019;
  assign n56010 = n23022 | n23023;
  assign n56011 = n23024 | n23025;
  assign n56012 = n23030 | ~n23031;
  assign n56013 = n23041 | n23042;
  assign n56014 = n23043 | n23044;
  assign n56015 = n23047 | n23048;
  assign n56016 = n23049 | n23050;
  assign n56017 = n23051 | ~n23052;
  assign n56018 = n23062 | n23063;
  assign n56019 = n23066 | ~n23067;
  assign n56020 = n23080 | n23081;
  assign n56021 = n23084 | ~n23085;
  assign n56022 = n23098 | n23099;
  assign n56023 = n23102 | ~n23103;
  assign n56024 = n23114 | n23115;
  assign n56025 = n23118 | n23119;
  assign n56026 = n23120 | n23121;
  assign n56027 = n23132 | n23133;
  assign n56028 = n23136 | ~n23137;
  assign n56029 = n23144 | ~n23145;
  assign n56030 = n23155 | n23156;
  assign n56031 = n23157 | n23158;
  assign n56032 = n23164 | n23165;
  assign n56033 = n23173 | n23174;
  assign n56034 = n23177 | ~n23178;
  assign n56035 = n23186 | n23187;
  assign n56036 = n23200 | n23201;
  assign n56037 = n23210 | ~n23211;
  assign n56038 = n23215 | n23216;
  assign n56039 = n23224 | n23225;
  assign n56040 = n23228 | n23229;
  assign n56041 = n23230 | n23231;
  assign n56042 = n23234 | n23235;
  assign n56043 = n23236 | n23237;
  assign n56044 = n23238 | ~n23239;
  assign n56045 = n23247 | n23248;
  assign n56046 = n23249 | n23250;
  assign n56047 = n23251 | ~n23252;
  assign n56048 = n23260 | n23261;
  assign n56049 = n23262 | n23263;
  assign n56050 = n23264 | ~n23265;
  assign n56051 = n23269 | n23270;
  assign n56052 = n23271 | n23272;
  assign n56053 = n23273 | ~n23274;
  assign n56054 = n23278 | n23279;
  assign n56055 = n23280 | n23281;
  assign n56056 = n23282 | ~n23283;
  assign n56057 = n23293 | ~n23294;
  assign n56058 = n23298 | n23299;
  assign n56059 = n23300 | n23301;
  assign n56060 = n23302 | ~n23303;
  assign n56061 = n23307 | n23308;
  assign n56062 = n23309 | n23310;
  assign n56063 = n23311 | ~n23312;
  assign n56064 = n23316 | n23317;
  assign n56065 = n23318 | n23319;
  assign n56066 = n23320 | ~n23321;
  assign n56067 = n23325 | n23326;
  assign n56068 = n23327 | n23328;
  assign n56069 = n23329 | ~n23330;
  assign n56070 = n23338 | n23339;
  assign n56071 = n23340 | n23341;
  assign n56072 = n23342 | ~n23343;
  assign n56073 = n23349 | ~n23350;
  assign n56074 = n23354 | n23355;
  assign n56075 = n23356 | n23357;
  assign n56076 = n23358 | ~n23359;
  assign n56077 = n23363 | n23364;
  assign n56078 = n23365 | n23366;
  assign n56079 = n23367 | ~n23368;
  assign n56080 = n23378 | ~n23379;
  assign n56081 = n23383 | n23384;
  assign n56082 = n23385 | n23386;
  assign n56083 = n23387 | ~n23388;
  assign n56084 = n23392 | n23393;
  assign n56085 = n23394 | n23395;
  assign n56086 = n23396 | ~n23397;
  assign n56087 = n23403 | ~n23404;
  assign n56088 = n23410 | ~n23411;
  assign n56089 = n23415 | n23416;
  assign n56090 = n23417 | n23418;
  assign n56091 = n23419 | ~n23420;
  assign n56092 = n23424 | n23425;
  assign n56093 = n23426 | n23427;
  assign n56094 = n23428 | ~n23429;
  assign n56095 = n23441 | n23442;
  assign n56096 = n23445 | n23446;
  assign n56097 = n23447 | n23448;
  assign n56098 = n23453 | ~n23454;
  assign n56099 = n23464 | ~n23465;
  assign n56100 = n23475 | ~n23476;
  assign n56101 = n23482 | ~n23483;
  assign n56102 = n23495 | n23496;
  assign n56103 = n23499 | ~n23500;
  assign n56104 = n23513 | n23514;
  assign n56105 = n23517 | ~n23518;
  assign n56106 = n23531 | n23532;
  assign n56107 = n23535 | ~n23536;
  assign n56108 = n23549 | n23550;
  assign n56109 = n23553 | ~n23554;
  assign n56110 = n23567 | n23568;
  assign n56111 = n23571 | ~n23572;
  assign n56112 = n23585 | n23586;
  assign n56113 = n23589 | ~n23590;
  assign n56114 = n23603 | n23604;
  assign n56115 = n23607 | ~n23608;
  assign n56116 = n23619 | n23620;
  assign n56117 = n23623 | n23624;
  assign n56118 = n23625 | n23626;
  assign n56119 = n23637 | n23638;
  assign n56120 = n23641 | n23642;
  assign n56121 = n23643 | n23644;
  assign n56122 = n23647 | n23648;
  assign n56123 = n23649 | n23650;
  assign n56124 = n23651 | ~n23652;
  assign n56125 = n23662 | n23663;
  assign n56126 = n23666 | ~n23667;
  assign n56127 = n23680 | n23681;
  assign n56128 = n23684 | ~n23685;
  assign n56129 = n23698 | n23699;
  assign n56130 = n23702 | ~n23703;
  assign n56131 = n23714 | n23715;
  assign n56132 = n23718 | n23719;
  assign n56133 = n23720 | n23721;
  assign n56134 = n23732 | n23733;
  assign n56135 = n23736 | n23737;
  assign n56136 = n23738 | n23739;
  assign n56137 = n23742 | n23743;
  assign n56138 = n23744 | n23745;
  assign n56139 = n23746 | ~n23747;
  assign n56140 = n23755 | n23756;
  assign n56141 = n23759 | n23760;
  assign n56142 = n23761 | n23762;
  assign n56143 = n23767 | ~n23768;
  assign n56144 = n23778 | n23779;
  assign n56145 = n23782 | ~n23783;
  assign n56146 = n23799 | n23796 | n23798;
  assign n56147 = n23802 | ~n23803;
  assign n56148 = n23816 | n23817;
  assign n56149 = n23820 | ~n23821;
  assign n56150 = n23832 | n23833;
  assign n56151 = n23836 | n23837;
  assign n56152 = n23838 | n23839;
  assign n56153 = n23850 | n23851;
  assign n56154 = n23854 | n23855;
  assign n56155 = n23856 | n23857;
  assign n56156 = n23862 | ~n23863;
  assign n56157 = n23873 | n23874;
  assign n56158 = n23875 | n23876;
  assign n56159 = n23879 | n23880;
  assign n56160 = n23881 | n23882;
  assign n56161 = n23883 | ~n23884;
  assign n56162 = n23894 | n23895;
  assign n56163 = n23898 | ~n23899;
  assign n56164 = n23912 | n23913;
  assign n56165 = n23916 | ~n23917;
  assign n56166 = n23930 | n23931;
  assign n56167 = n23934 | ~n23935;
  assign n56168 = n23946 | n23947;
  assign n56169 = n23950 | n23951;
  assign n56170 = n23952 | n23953;
  assign n56171 = n23964 | n23965;
  assign n56172 = n23968 | ~n23969;
  assign n56173 = n23976 | ~n23977;
  assign n56174 = n23987 | n23988;
  assign n56175 = n23989 | n23990;
  assign n56176 = n23996 | n23997;
  assign n56177 = n24005 | n24006;
  assign n56178 = n24009 | ~n24010;
  assign n56179 = n24018 | n24019;
  assign n56180 = n24032 | n24033;
  assign n56181 = n24042 | ~n24043;
  assign n56182 = n24047 | n24048;
  assign n56183 = n24056 | n24057;
  assign n56184 = n24060 | n24061;
  assign n56185 = n24062 | n24063;
  assign n56186 = n24066 | n24067;
  assign n56187 = n24068 | n24069;
  assign n56188 = n24070 | ~n24071;
  assign n56189 = n24079 | n24080;
  assign n56190 = n24081 | n24082;
  assign n56191 = n24083 | ~n24084;
  assign n56192 = n24092 | n24093;
  assign n56193 = n24094 | n24095;
  assign n56194 = n24096 | ~n24097;
  assign n56195 = n24101 | n24102;
  assign n56196 = n24103 | n24104;
  assign n56197 = n24105 | ~n24106;
  assign n56198 = n24110 | n24111;
  assign n56199 = n24112 | n24113;
  assign n56200 = n24114 | ~n24115;
  assign n56201 = n24125 | ~n24126;
  assign n56202 = n24130 | n24131;
  assign n56203 = n24132 | n24133;
  assign n56204 = n24134 | ~n24135;
  assign n56205 = n24139 | n24140;
  assign n56206 = n24141 | n24142;
  assign n56207 = n24143 | ~n24144;
  assign n56208 = n24148 | n24149;
  assign n56209 = n24150 | n24151;
  assign n56210 = n24152 | ~n24153;
  assign n56211 = n24157 | n24158;
  assign n56212 = n24159 | n24160;
  assign n56213 = n24161 | ~n24162;
  assign n56214 = n24170 | n24171;
  assign n56215 = n24172 | n24173;
  assign n56216 = n24174 | ~n24175;
  assign n56217 = n24181 | ~n24182;
  assign n56218 = n24186 | n24187;
  assign n56219 = n24188 | n24189;
  assign n56220 = n24190 | ~n24191;
  assign n56221 = n24195 | n24196;
  assign n56222 = n24197 | n24198;
  assign n56223 = n24199 | ~n24200;
  assign n56224 = n24204 | n24205;
  assign n56225 = n24206 | n24207;
  assign n56226 = n24208 | ~n24209;
  assign n56227 = n24219 | ~n24220;
  assign n56228 = n24224 | n24225;
  assign n56229 = n24226 | n24227;
  assign n56230 = n24228 | ~n24229;
  assign n56231 = n24233 | n24234;
  assign n56232 = n24235 | n24236;
  assign n56233 = n24237 | ~n24238;
  assign n56234 = n24242 | n24243;
  assign n56235 = n24244 | n24245;
  assign n56236 = n24246 | ~n24247;
  assign n56237 = n24251 | n24252;
  assign n56238 = n24253 | n24254;
  assign n56239 = n24255 | ~n24256;
  assign n56240 = n24260 | n24261;
  assign n56241 = n24262 | n24263;
  assign n56242 = n24264 | ~n24265;
  assign n56243 = n24269 | n24270;
  assign n56244 = n24271 | n24272;
  assign n56245 = n24273 | ~n24274;
  assign n56246 = n24278 | n24279;
  assign n56247 = n24280 | n24281;
  assign n56248 = n24282 | ~n24283;
  assign n56249 = n24287 | n24288;
  assign n56250 = n24289 | n24290;
  assign n56251 = n24291 | ~n24292;
  assign n56252 = n24296 | n24297;
  assign n56253 = n24307 | n24308;
  assign n56254 = n24311 | n24312;
  assign n56255 = n24313 | n24314;
  assign n56256 = n24319 | ~n24320;
  assign n56257 = n24327 | n24328;
  assign n56258 = n24335 | ~n24336;
  assign n56259 = n24343 | ~n24344;
  assign n56260 = n24346 | n24347;
  assign n56261 = n24348 | n24349;
  assign n56262 = n24357 | n24358;
  assign n56263 = n24361 | n24362;
  assign n56264 = n24363 | n24364;
  assign n56265 = n24369 | n24370;
  assign n56266 = n24371 | n24372;
  assign n56267 = n24373 | ~n24374;
  assign n56268 = n24378 | ~n24379;
  assign n56269 = n24381 | n24382;
  assign n56270 = n24392 | n24393;
  assign n56271 = n24394 | n24395;
  assign n56272 = n24398 | n24399;
  assign n56273 = n24400 | n24401;
  assign n56274 = n24402 | ~n24403;
  assign n56275 = n24411 | n24412;
  assign n56276 = n24415 | n24416;
  assign n56277 = n24417 | n24418;
  assign n56278 = n24423 | ~n24424;
  assign n56279 = n24432 | n24433;
  assign n56280 = n24436 | n24437;
  assign n56281 = n24438 | n24439;
  assign n56282 = n24444 | ~n24445;
  assign n56283 = n24453 | n24454;
  assign n56284 = n24457 | n24458;
  assign n56285 = n24459 | n24460;
  assign n56286 = n24463 | n24464;
  assign n56287 = n24465 | n24466;
  assign n56288 = n24467 | ~n24468;
  assign n56289 = n24476 | n24477;
  assign n56290 = n24480 | n24481;
  assign n56291 = n24482 | n24483;
  assign n56292 = n24486 | n24487;
  assign n56293 = n24488 | n24489;
  assign n56294 = n24490 | ~n24491;
  assign n56295 = n24499 | n24500;
  assign n56296 = n24503 | n24504;
  assign n56297 = n24505 | n24506;
  assign n56298 = n24511 | ~n24512;
  assign n56299 = n24522 | n24523;
  assign n56300 = n24526 | ~n24527;
  assign n56301 = n24540 | n24541;
  assign n56302 = n24544 | ~n24545;
  assign n56303 = n24556 | n24557;
  assign n56304 = n24560 | n24561;
  assign n56305 = n24562 | n24563;
  assign n56306 = n24574 | n24575;
  assign n56307 = n24578 | n24579;
  assign n56308 = n24580 | n24581;
  assign n56309 = n24586 | ~n24587;
  assign n56310 = n24595 | n24596;
  assign n56311 = n24599 | n24600;
  assign n56312 = n24601 | n24602;
  assign n56313 = n24605 | n24606;
  assign n56314 = n24607 | n24608;
  assign n56315 = n24609 | ~n24610;
  assign n56316 = n24620 | n24621;
  assign n56317 = n24624 | ~n24625;
  assign n56318 = n24638 | n24639;
  assign n56319 = n24642 | ~n24643;
  assign n56320 = n24656 | n24657;
  assign n56321 = n24660 | ~n24661;
  assign n56322 = n24672 | n24673;
  assign n56323 = n24676 | n24677;
  assign n56324 = n24678 | n24679;
  assign n56325 = n24690 | n24691;
  assign n56326 = n24694 | n24695;
  assign n56327 = n24696 | n24697;
  assign n56328 = n24700 | n24701;
  assign n56329 = n24702 | n24703;
  assign n56330 = n24704 | ~n24705;
  assign n56331 = n24713 | n24714;
  assign n56332 = n24717 | n24718;
  assign n56333 = n24719 | n24720;
  assign n56334 = n24725 | ~n24726;
  assign n56335 = n24736 | n24737;
  assign n56336 = n24740 | ~n24741;
  assign n56337 = n24757 | n24754 | n24756;
  assign n56338 = n24760 | ~n24761;
  assign n56339 = n24774 | n24775;
  assign n56340 = n24778 | ~n24779;
  assign n56341 = n24790 | n24791;
  assign n56342 = n24794 | n24795;
  assign n56343 = n24796 | n24797;
  assign n56344 = n24808 | n24809;
  assign n56345 = n24812 | n24813;
  assign n56346 = n24814 | n24815;
  assign n56347 = n24820 | ~n24821;
  assign n56348 = n24831 | n24832;
  assign n56349 = n24833 | n24834;
  assign n56350 = n24837 | n24838;
  assign n56351 = n24839 | n24840;
  assign n56352 = n24841 | ~n24842;
  assign n56353 = n24852 | n24853;
  assign n56354 = n24856 | ~n24857;
  assign n56355 = n24870 | n24871;
  assign n56356 = n24874 | ~n24875;
  assign n56357 = n24888 | n24889;
  assign n56358 = n24892 | ~n24893;
  assign n56359 = n24904 | n24905;
  assign n56360 = n24908 | n24909;
  assign n56361 = n24910 | n24911;
  assign n56362 = n24922 | n24923;
  assign n56363 = n24926 | ~n24927;
  assign n56364 = n24934 | ~n24935;
  assign n56365 = n24945 | n24946;
  assign n56366 = n24947 | n24948;
  assign n56367 = n24954 | n24955;
  assign n56368 = n24963 | n24964;
  assign n56369 = n24967 | ~n24968;
  assign n56370 = n24976 | n24977;
  assign n56371 = n24990 | n24991;
  assign n56372 = n25000 | ~n25001;
  assign n56373 = n25005 | n25006;
  assign n56374 = n25014 | n25015;
  assign n56375 = n25018 | n25019;
  assign n56376 = n25020 | n25021;
  assign n56377 = n25024 | n25025;
  assign n56378 = n25026 | n25027;
  assign n56379 = n25028 | ~n25029;
  assign n56380 = n25037 | n25038;
  assign n56381 = n25039 | n25040;
  assign n56382 = n25041 | ~n25042;
  assign n56383 = n25050 | n25051;
  assign n56384 = n25052 | n25053;
  assign n56385 = n25054 | ~n25055;
  assign n56386 = n25059 | n25060;
  assign n56387 = n25061 | n25062;
  assign n56388 = n25063 | ~n25064;
  assign n56389 = n25068 | n25069;
  assign n56390 = n25070 | n25071;
  assign n56391 = n25072 | ~n25073;
  assign n56392 = n25083 | ~n25084;
  assign n56393 = n25088 | n25089;
  assign n56394 = n25090 | n25091;
  assign n56395 = n25092 | ~n25093;
  assign n56396 = n25097 | n25098;
  assign n56397 = n25099 | n25100;
  assign n56398 = n25101 | ~n25102;
  assign n56399 = n25106 | n25107;
  assign n56400 = n25108 | n25109;
  assign n56401 = n25110 | ~n25111;
  assign n56402 = n25115 | n25116;
  assign n56403 = n25117 | n25118;
  assign n56404 = n25119 | ~n25120;
  assign n56405 = n25128 | n25129;
  assign n56406 = n25130 | n25131;
  assign n56407 = n25132 | ~n25133;
  assign n56408 = n25139 | ~n25140;
  assign n56409 = n25144 | n25145;
  assign n56410 = n25146 | n25147;
  assign n56411 = n25148 | ~n25149;
  assign n56412 = n25153 | n25154;
  assign n56413 = n25155 | n25156;
  assign n56414 = n25157 | ~n25158;
  assign n56415 = n25162 | n25163;
  assign n56416 = n25164 | n25165;
  assign n56417 = n25166 | ~n25167;
  assign n56418 = n25177 | ~n25178;
  assign n56419 = n25182 | n25183;
  assign n56420 = n25184 | n25185;
  assign n56421 = n25186 | ~n25187;
  assign n56422 = n25191 | n25192;
  assign n56423 = n25193 | n25194;
  assign n56424 = n25195 | ~n25196;
  assign n56425 = n25200 | n25201;
  assign n56426 = n25202 | n25203;
  assign n56427 = n25204 | ~n25205;
  assign n56428 = n25213 | n25214;
  assign n56429 = n25215 | n25216;
  assign n56430 = n25217 | ~n25218;
  assign n56431 = n25224 | ~n25225;
  assign n56432 = n25231 | ~n25232;
  assign n56433 = n25236 | n25237;
  assign n56434 = n25238 | n25239;
  assign n56435 = n25240 | ~n25241;
  assign n56436 = n25245 | n25246;
  assign n56437 = n25247 | n25248;
  assign n56438 = n25249 | ~n25250;
  assign n56439 = n25256 | ~n25257;
  assign n56440 = n25263 | ~n25264;
  assign n56441 = n25277 | ~n25278;
  assign n56442 = n25292 | n25293;
  assign n56443 = n25296 | ~n25297;
  assign n56444 = n25310 | n25311;
  assign n56445 = n25314 | ~n25315;
  assign n56446 = n25330 | ~n25331;
  assign n56447 = n25344 | n25345;
  assign n56448 = n25348 | ~n25349;
  assign n56449 = n25360 | n25361;
  assign n56450 = n25364 | ~n25365;
  assign n56451 = n25375 | n25376;
  assign n56452 = n25388 | n25389;
  assign n56453 = n25392 | ~n25393;
  assign n56454 = n25403 | n25404;
  assign n56455 = n25407 | n25408;
  assign n56456 = n25420 | n25421;
  assign n56457 = n25424 | ~n25425;
  assign n56458 = n25435 | n25436;
  assign n56459 = n25439 | n25440;
  assign n56460 = n25452 | n25453;
  assign n56461 = n25456 | ~n25457;
  assign n56462 = n25467 | n25468;
  assign n56463 = n25471 | n25472;
  assign n56464 = n25484 | n25485;
  assign n56465 = n25488 | ~n25489;
  assign n56466 = n25509 | ~n25510;
  assign n56467 = ~n25519 | n25516 | n25518;
  assign n56468 = n25527 | n25528;
  assign n56469 = n25531 | ~n25532;
  assign n56470 = n25542 | n25543;
  assign n56471 = n25556 | ~n25557;
  assign n56472 = n25577 | n25578;
  assign n56473 = n25579 | n25580;
  assign n56474 = n25592 | n25587 | n25591;
  assign n56475 = n25596 | ~n25597;
  assign n56476 = n25598 | n25599;
  assign n56477 = n25606 | n25607;
  assign n56478 = n25618 | n25615 | ~n25617;
  assign n56479 = n25627 | n25628;
  assign n56480 = n25631 | ~n25632;
  assign n56481 = n25647 | n25642 | ~n25646;
  assign n56482 = n25655 | n25656;
  assign n56483 = n25662 | ~n25663;
  assign n56484 = n25673 | ~n25674;
  assign n56485 = n25683 | n25684;
  assign n56486 = n25687 | ~n25688;
  assign n56487 = n25696 | ~n25697;
  assign n56488 = n25706 | n25707;
  assign n56489 = n25710 | ~n25711;
  assign n56490 = n25719 | ~n25720;
  assign n56491 = n25734 | ~n25735;
  assign n56492 = n25746 | n25747;
  assign n56493 = n25753 | ~n25754;
  assign n56494 = n25764 | n25765;
  assign n56495 = n25771 | ~n25772;
  assign n56496 = n25782 | ~n25783;
  assign n56497 = n25795 | n25792 | n25794;
  assign n56498 = n25798 | ~n25799;
  assign n56499 = n25807 | ~n25808;
  assign n56500 = n25817 | n25818;
  assign n56501 = n25821 | ~n25822;
  assign n56502 = n25830 | ~n25831;
  assign n56503 = n25840 | n25841;
  assign n56504 = n25847 | ~n25848;
  assign n56505 = n25859 | n25860;
  assign n56506 = n25866 | ~n25867;
  assign n56507 = n25877 | n25878;
  assign n56508 = n25884 | ~n25885;
  assign n56509 = n25895 | ~n25896;
  assign n56510 = n25905 | n25906;
  assign n56511 = n25909 | ~n25910;
  assign n56512 = n25918 | ~n25919;
  assign n56513 = n25928 | n25929;
  assign n56514 = n25932 | ~n25933;
  assign n56515 = n25941 | ~n25942;
  assign n56516 = n25951 | n25952;
  assign n56517 = n25958 | ~n25959;
  assign n56518 = n25970 | n25971;
  assign n56519 = n25977 | ~n25978;
  assign n56520 = n25988 | n25989;
  assign n56521 = n25995 | ~n25996;
  assign n56522 = n26006 | ~n26007;
  assign n56523 = n26016 | n26017;
  assign n56524 = n26020 | ~n26021;
  assign n56525 = n26029 | ~n26030;
  assign n56526 = n26039 | n26040;
  assign n56527 = n26043 | ~n26044;
  assign n56528 = n26052 | ~n26053;
  assign n56529 = n26062 | n26063;
  assign n56530 = n26069 | ~n26070;
  assign n56531 = n26080 | n26081;
  assign n56532 = n26087 | ~n26088;
  assign n56533 = n26098 | ~n26099;
  assign n56534 = n26101 | n26102;
  assign n56535 = n26103 | n26104;
  assign n56536 = n26105 | ~n26106;
  assign n56537 = n26202 | ~n26203;
  assign n56538 = n26223 | n26224;
  assign n56539 = n26225 | n26226;
  assign n56540 = n26234 | n26235;
  assign n56541 = n26350 | n26351;
  assign n56542 = n26352 | n26353;
  assign n56543 = n26354 | ~n26355;
  assign n56544 = n26360 | ~n26361;
  assign n56545 = n26371 | n26372;
  assign n56546 = n26377 | n26378;
  assign n56547 = n26387 | n26388;
  assign n56548 = n26393 | n26394;
  assign n56549 = n26403 | n26404;
  assign n56550 = n26413 | n26414;
  assign n56551 = n26419 | n26420;
  assign n56552 = n26425 | n26426;
  assign n56553 = n26435 | n26436;
  assign n56554 = n26453 | n26454;
  assign n56555 = n26459 | n26460;
  assign n56556 = n26473 | n26474;
  assign n56557 = n26479 | n26480;
  assign n56558 = n26485 | n26486;
  assign n56559 = n26499 | n26500;
  assign n56560 = n26509 | n26510;
  assign n56561 = n26519 | n26520;
  assign n56562 = n26532 | n26533;
  assign n56563 = n26534 | n26535;
  assign n56564 = n26543 | ~n26544;
  assign n56565 = n26553 | n26554;
  assign n56566 = n26555 | n26556;
  assign n56567 = n26561 | ~n26562;
  assign n56568 = n26571 | n26572;
  assign n56569 = n26573 | n26574;
  assign n56570 = n26578 | n26579;
  assign n56571 = n26584 | n26585;
  assign n56572 = n26594 | n26595;
  assign n56573 = n26598 | n26599;
  assign n56574 = n26613 | n26608 | n26612;
  assign n56575 = n26622 | n26623;
  assign n56576 = n26628 | n26629;
  assign n56577 = n26642 | n26643;
  assign n56578 = n26647 | n26653 | n26656 | n26657;
  assign n56579 = n26675 | n26667 | n26674;
  assign n56580 = n26671 | n26672;
  assign n56581 = n26677 | n26678;
  assign n56582 = n26690 | n26691;
  assign n56583 = n26702 | n26699 | n26701;
  assign n56584 = n26709 | n26703 | n26708;
  assign n56585 = n26712 | n26713;
  assign n56586 = n26716 | n26717;
  assign n56587 = n26720 | n26721;
  assign n56588 = n26724 | n26725;
  assign n56589 = n26738 | n26739;
  assign n56590 = n26755 | n26748 | n26754;
  assign n56591 = n26799 | n26786 | n26798;
  assign n56592 = n26818 | n26819;
  assign n56593 = n26822 | n26823;
  assign n56594 = n26827 | n26828;
  assign n56595 = n26831 | n26832;
  assign n56596 = n26837 | n26838;
  assign n56597 = n26843 | n26844;
  assign n56598 = n26850 | n26851;
  assign n56599 = n26867 | n26868;
  assign n56600 = n26871 | n26873 | n26875 | n26876;
  assign n56601 = n26890 | ~n26891;
  assign n56602 = n26900 | n26901;
  assign n56603 = n26910 | n26911;
  assign n56604 = n26918 | n26919;
  assign n56605 = n26952 | n26937 | n26951;
  assign n56606 = n26986 | n26987;
  assign n56607 = n27001 | n26988 | n27000;
  assign n56608 = n27016 | n27017;
  assign n56609 = n27036 | n27037;
  assign n56610 = n27051 | n27052;
  assign n56611 = n27057 | ~n27058;
  assign n56612 = n27067 | ~n27068;
  assign n56613 = n27084 | n27085;
  assign n56614 = n27093 | n27094;
  assign n56615 = n27108 | n27102 | n27107;
  assign n56616 = n27123 | n27124;
  assign n56617 = n27125 | n27126;
  assign n56618 = n27128 | n27129;
  assign n56619 = n27134 | n27135;
  assign n56620 = n27142 | n27143;
  assign n56621 = n27146 | n27147;
  assign n56622 = n27161 | n27154 | n27160;
  assign n56623 = n27173 | n27174;
  assign n56624 = n27185 | n27186;
  assign n56625 = n27204 | n27205;
  assign n56626 = n27209 | n27210;
  assign n56627 = n27232 | n27223 | n27231;
  assign n56628 = n27248 | n27249;
  assign n56629 = n27252 | n27253;
  assign n56630 = n27266 | n27269 | n27273 | n27274;
  assign n56631 = n27292 | n27293;
  assign n56632 = n27310 | n27311;
  assign n56633 = n27318 | n27315 | n27317;
  assign n56634 = n27339 | n27340;
  assign n56635 = n27346 | n27347;
  assign n56636 = n27350 | n27351;
  assign n56637 = n27352 | n27353;
  assign n56638 = n27354 | ~n27355;
  assign n56639 = n27366 | ~n27367;
  assign n56640 = n27376 | ~n27377;
  assign n56641 = n27396 | n27397;
  assign n56642 = n27398 | n27399;
  assign n56643 = n27403 | n27404;
  assign n56644 = n27405 | n27406;
  assign n56645 = n27407 | ~n27408;
  assign n56646 = n27413 | ~n27414;
  assign n56647 = n27420 | ~n27421;
  assign n56648 = n27425 | ~n27426;
  assign n56649 = n27443 | ~n27444;
  assign n56650 = n27449 | n27450;
  assign n56651 = n27451 | n27452;
  assign n56652 = n27453 | ~n27454;
  assign n56653 = n27458 | n27459;
  assign n56654 = n27460 | n27461;
  assign n56655 = n27462 | ~n27463;
  assign n56656 = n27475 | n27476;
  assign n56657 = n27477 | n27478;
  assign n56658 = n27484 | ~n27485;
  assign n56659 = n27487 | n27488;
  assign n56660 = n27500 | n27501;
  assign n56661 = n27502 | n27503;
  assign n56662 = n27509 | n27510;
  assign n56663 = n27515 | n27516;
  assign n56664 = n27517 | n27518;
  assign n56665 = n27520 | ~n27521;
  assign n56666 = n27522 | ~n27523;
  assign n56667 = n27528 | n27525 | n27527;
  assign n56668 = n27535 | ~n27536;
  assign n56669 = n27545 | n27546;
  assign n56670 = n27547 | n27548;
  assign n56671 = n27550 | n27551;
  assign n56672 = n27552 | n27553;
  assign n56673 = n27555 | ~n27556;
  assign n56674 = n27559 | n27560;
  assign n56675 = n27561 | n27562;
  assign n56676 = n27563 | ~n27564;
  assign n56677 = n27575 | n27576;
  assign n56678 = n27586 | n27581 | n27585;
  assign n56679 = n27605 | n27612 | n27623 | n27624;
  assign n56680 = n27633 | n27634;
  assign n56681 = n27643 | n27639 | n27642;
  assign n56682 = n27652 | n27653;
  assign n56683 = n27661 | n27662;
  assign n56684 = n27698 | n27681 | n27697;
  assign n56685 = n27717 | n27718;
  assign n56686 = n27725 | ~n27726;
  assign n56687 = n27735 | n27736;
  assign n56688 = n27754 | n27755;
  assign n56689 = n27767 | ~n27768;
  assign n56690 = n27786 | n27787;
  assign n56691 = n27788 | n27789;
  assign n56692 = n27794 | n27795;
  assign n56693 = n27798 | n27799;
  assign n56694 = n27800 | n27801;
  assign n56695 = n27803 | ~n27804;
  assign n56696 = n27817 | n27818;
  assign n56697 = n27819 | n27820;
  assign n56698 = n27825 | n27826;
  assign n56699 = n27834 | ~n27835;
  assign n56700 = n27848 | n27849;
  assign n56701 = n27850 | n27851;
  assign n56702 = n27855 | n27856;
  assign n56703 = n27857 | n27858;
  assign n56704 = n27859 | ~n27860;
  assign n56705 = n27864 | ~n27865;
  assign n56706 = n27874 | n27875;
  assign n56707 = n27876 | n27877;
  assign n56708 = n27882 | ~n27883;
  assign n56709 = n27893 | n27896 | n27899 | n27900;
  assign n56710 = n27924 | n27931 | n27940 | n27941;
  assign n56711 = n27946 | n27947;
  assign n56712 = n27963 | n27976 | n27985 | n27986;
  assign n56713 = n28003 | n28004;
  assign n56714 = n28010 | n28011;
  assign n56715 = n28015 | n28016;
  assign n56716 = n28035 | n28029 | n28034;
  assign n56717 = n28042 | n28043;
  assign n56718 = n28059 | n28060;
  assign n56719 = n28062 | ~n28063;
  assign n56720 = n28068 | n28065 | n28067;
  assign n56721 = n28082 | ~n28083;
  assign n56722 = n28092 | n28093;
  assign n56723 = n28099 | ~n28100;
  assign n56724 = n28121 | n28118 | n28120;
  assign n56725 = n28124 | n28125;
  assign n56726 = n28135 | n28132 | n28134;
  assign n56727 = n28138 | n28139;
  assign n56728 = n28146 | n28147;
  assign n56729 = n28170 | n28158 | n28169;
  assign n56730 = n28185 | n28186;
  assign n56731 = n28193 | n28194;
  assign n56732 = n28201 | n28206 | n28210 | n28211;
  assign n56733 = n28216 | n28217;
  assign n56734 = n28224 | n28225;
  assign n56735 = n28235 | n28236;
  assign n56736 = n28254 | n28255;
  assign n56737 = n28261 | n28262;
  assign n56738 = n28267 | n28268;
  assign n56739 = n28272 | n28273;
  assign n56740 = n28276 | n28277;
  assign n56741 = n28280 | n28281;
  assign n56742 = n28289 | n28290;
  assign n56743 = n28296 | n28293 | n28295;
  assign n56744 = n28328 | n28316 | n28322 | n28336 | n28337;
  assign n56745 = n28344 | n28345;
  assign n56746 = n28356 | n28362 | n28371 | n28372;
  assign n56747 = n28389 | n28390;
  assign n56748 = n28398 | n28399;
  assign n56749 = n28407 | n28408;
  assign n56750 = n28418 | n28419;
  assign n56751 = n28423 | n28424;
  assign n56752 = n28428 | n28429;
  assign n56753 = n28454 | n28445 | n28453;
  assign n56754 = n28472 | n28473;
  assign n56755 = n28475 | ~n28476;
  assign n56756 = n28481 | n28478 | n28480;
  assign n56757 = n28502 | n28503;
  assign n56758 = n28509 | n28510;
  assign n56759 = n28513 | n28514;
  assign n56760 = n28515 | n28516;
  assign n56761 = n28517 | ~n28518;
  assign n56762 = n28534 | ~n28535;
  assign n56763 = n28546 | ~n28547;
  assign n56764 = n28562 | n28563;
  assign n56765 = n28564 | n28565;
  assign n56766 = n28570 | n28571;
  assign n56767 = n28582 | n28583;
  assign n56768 = n28584 | n28585;
  assign n56769 = n28590 | n28591;
  assign n56770 = n28595 | n28596;
  assign n56771 = n28597 | n28598;
  assign n56772 = n28599 | ~n28600;
  assign n56773 = n28608 | n28605 | n28607;
  assign n56774 = n28611 | n28612;
  assign n56775 = n28613 | n28614;
  assign n56776 = n28619 | n28620;
  assign n56777 = n28630 | n28631;
  assign n56778 = n28634 | n28635;
  assign n56779 = n28636 | n28637;
  assign n56780 = n28642 | ~n28643;
  assign n56781 = n28654 | n28655;
  assign n56782 = n28656 | n28657;
  assign n56783 = n28670 | n28671;
  assign n56784 = n28672 | n28673;
  assign n56785 = n28684 | n28685;
  assign n56786 = n28686 | n28687;
  assign n56787 = n28690 | n28691;
  assign n56788 = n28692 | n28693;
  assign n56789 = n28694 | ~n28695;
  assign n56790 = n28699 | n28700;
  assign n56791 = n28701 | n28702;
  assign n56792 = n28703 | ~n28704;
  assign n56793 = n28710 | ~n28711;
  assign n56794 = n28722 | n28723;
  assign n56795 = n28724 | n28725;
  assign n56796 = n28730 | n28731;
  assign n56797 = n28742 | n28743;
  assign n56798 = n28744 | n28745;
  assign n56799 = n28750 | n28751;
  assign n56800 = n28756 | n28757;
  assign n56801 = n28758 | n28759;
  assign n56802 = n28760 | ~n28761;
  assign n56803 = n28767 | ~n28768;
  assign n56804 = n28782 | n28783;
  assign n56805 = n28784 | n28785;
  assign n56806 = n28789 | n28790;
  assign n56807 = n28791 | n28792;
  assign n56808 = n28793 | ~n28794;
  assign n56809 = n28798 | ~n28799;
  assign n56810 = n28805 | ~n28806;
  assign n56811 = n28825 | ~n28826;
  assign n56812 = n28831 | n28832;
  assign n56813 = n28833 | n28834;
  assign n56814 = n28835 | ~n28836;
  assign n56815 = n28840 | n28841;
  assign n56816 = n28842 | n28843;
  assign n56817 = n28844 | ~n28845;
  assign n56818 = n28856 | n28857;
  assign n56819 = n28858 | n28859;
  assign n56820 = n28864 | ~n28865;
  assign n56821 = n28867 | n28868;
  assign n56822 = n28879 | n28880;
  assign n56823 = n28881 | n28882;
  assign n56824 = n28887 | n28888;
  assign n56825 = n28899 | n28900;
  assign n56826 = n28901 | n28902;
  assign n56827 = n28907 | n28908;
  assign n56828 = n28911 | n28912;
  assign n56829 = n28913 | n28914;
  assign n56830 = n28916 | ~n28917;
  assign n56831 = n28928 | n28929;
  assign n56832 = n28930 | n28931;
  assign n56833 = n28936 | n28937;
  assign n56834 = n28943 | ~n28944;
  assign n56835 = n28948 | n28949;
  assign n56836 = n28954 | ~n28955;
  assign n56837 = n28966 | n28967;
  assign n56838 = n28968 | n28969;
  assign n56839 = n28973 | n28974;
  assign n56840 = n28975 | n28976;
  assign n56841 = n28977 | ~n28978;
  assign n56842 = n28982 | ~n28983;
  assign n56843 = n28992 | n28993;
  assign n56844 = n28994 | n28995;
  assign n56845 = n29000 | ~n29001;
  assign n56846 = n29004 | n29005;
  assign n56847 = n29006 | n29007;
  assign n56848 = n29008 | ~n29009;
  assign n56849 = n29019 | n29020;
  assign n56850 = n29046 | n29033 | n29045;
  assign n56851 = n29064 | n29065;
  assign n56852 = n29067 | ~n29068;
  assign n56853 = n29070 | n29071;
  assign n56854 = n29077 | n29074 | n29076;
  assign n56855 = n29079 | n29080;
  assign n56856 = n29092 | n29093;
  assign n56857 = n29103 | n29113 | n29121 | n29122;
  assign n56858 = n29127 | n29128;
  assign n56859 = n29142 | n29143;
  assign n56860 = n29153 | n29154;
  assign n56861 = n29171 | n29165 | n29170;
  assign n56862 = n29188 | n29189;
  assign n56863 = n29197 | n29193 | n29196;
  assign n56864 = n29194 | n29195;
  assign n56865 = n29204 | ~n29205;
  assign n56866 = n29207 | n29208;
  assign n56867 = n29216 | ~n29217;
  assign n56868 = n29226 | n29227;
  assign n56869 = n29233 | n29234;
  assign n56870 = n29243 | ~n29244;
  assign n56871 = n29255 | n29256;
  assign n56872 = n29268 | ~n29269;
  assign n56873 = n29287 | n29288;
  assign n56874 = n29289 | n29290;
  assign n56875 = n29295 | n29296;
  assign n56876 = n29302 | ~n29303;
  assign n56877 = n29314 | n29315;
  assign n56878 = n29316 | n29317;
  assign n56879 = n29322 | n29323;
  assign n56880 = n29334 | n29335;
  assign n56881 = n29336 | n29337;
  assign n56882 = n29342 | n29343;
  assign n56883 = n29349 | ~n29350;
  assign n56884 = n29358 | n29355 | n29357;
  assign n56885 = n29361 | n29362;
  assign n56886 = n29363 | n29364;
  assign n56887 = n29369 | n29370;
  assign n56888 = n29379 | n29380;
  assign n56889 = n29383 | n29384;
  assign n56890 = n29385 | n29386;
  assign n56891 = n29391 | ~n29392;
  assign n56892 = n29403 | n29404;
  assign n56893 = n29405 | n29406;
  assign n56894 = n29410 | n29411;
  assign n56895 = n29412 | n29413;
  assign n56896 = n29414 | ~n29415;
  assign n56897 = n29419 | ~n29420;
  assign n56898 = n29429 | n29430;
  assign n56899 = n29431 | n29432;
  assign n56900 = n29437 | ~n29438;
  assign n56901 = n29443 | ~n29444;
  assign n56902 = n29482 | n29472 | n29481;
  assign n56903 = n29503 | n29504;
  assign n56904 = n29508 | n29509;
  assign n56905 = n29550 | n29534 | n29549;
  assign n56906 = n29569 | n29570;
  assign n56907 = n29578 | n29579;
  assign n56908 = n29591 | n29592;
  assign n56909 = n29602 | n29603;
  assign n56910 = n29606 | n29612 | n29615 | n29616;
  assign n56911 = n29628 | n29629;
  assign n56912 = n29632 | n29633;
  assign n56913 = n29638 | n29639;
  assign n56914 = n29645 | n29646;
  assign n56915 = n29655 | n29656;
  assign n56916 = n29663 | n29664;
  assign n56917 = n29671 | n29672;
  assign n56918 = n29700 | n29688 | n29699;
  assign n56919 = n29717 | n29718;
  assign n56920 = n29724 | ~n29725;
  assign n56921 = n29738 | n29735 | n29737;
  assign n56922 = n29739 | n29740;
  assign n56923 = n29742 | n29743;
  assign n56924 = n29748 | n29749;
  assign n56925 = n29754 | n29755;
  assign n56926 = n29756 | ~n29757;
  assign n56927 = n29762 | ~n29763;
  assign n56928 = n29767 | ~n29768;
  assign n56929 = n29791 | ~n29792;
  assign n56930 = n29799 | n29800;
  assign n56931 = n29801 | n29802;
  assign n56932 = n29803 | ~n29804;
  assign n56933 = n29810 | ~n29811;
  assign n56934 = n29826 | n29827;
  assign n56935 = n29828 | n29829;
  assign n56936 = n29834 | n29835;
  assign n56937 = n29846 | n29847;
  assign n56938 = n29848 | n29849;
  assign n56939 = n29854 | n29855;
  assign n56940 = n29858 | n29859;
  assign n56941 = n29860 | n29861;
  assign n56942 = n29863 | ~n29864;
  assign n56943 = n29875 | n29876;
  assign n56944 = n29877 | n29878;
  assign n56945 = n29883 | n29884;
  assign n56946 = n29895 | n29896;
  assign n56947 = n29897 | n29898;
  assign n56948 = n29903 | n29904;
  assign n56949 = n29909 | n29910;
  assign n56950 = n29911 | n29912;
  assign n56951 = n29913 | ~n29914;
  assign n56952 = n29917 | n29918;
  assign n56953 = n29919 | n29920;
  assign n56954 = n29922 | ~n29923;
  assign n56955 = n29937 | n29938;
  assign n56956 = n29939 | n29940;
  assign n56957 = n29944 | n29945;
  assign n56958 = n29946 | n29947;
  assign n56959 = n29948 | ~n29949;
  assign n56960 = n29953 | ~n29954;
  assign n56961 = n29965 | n29966;
  assign n56962 = n29967 | n29968;
  assign n56963 = n29981 | n29982;
  assign n56964 = n29983 | n29984;
  assign n56965 = n29995 | n29996;
  assign n56966 = n29997 | n29998;
  assign n56967 = n30001 | n30002;
  assign n56968 = n30003 | n30004;
  assign n56969 = n30005 | ~n30006;
  assign n56970 = n30010 | n30011;
  assign n56971 = n30012 | n30013;
  assign n56972 = n30014 | ~n30015;
  assign n56973 = n30021 | ~n30022;
  assign n56974 = n30033 | n30034;
  assign n56975 = n30035 | n30036;
  assign n56976 = n30041 | n30042;
  assign n56977 = n30053 | n30054;
  assign n56978 = n30055 | n30056;
  assign n56979 = n30061 | n30062;
  assign n56980 = n30068 | ~n30069;
  assign n56981 = n30080 | n30081;
  assign n56982 = n30082 | n30083;
  assign n56983 = n30088 | n30089;
  assign n56984 = n30095 | ~n30096;
  assign n56985 = n30100 | n30101;
  assign n56986 = n30106 | ~n30107;
  assign n56987 = n30118 | n30119;
  assign n56988 = n30120 | n30121;
  assign n56989 = n30125 | n30126;
  assign n56990 = n30127 | n30128;
  assign n56991 = n30129 | ~n30130;
  assign n56992 = n30134 | ~n30135;
  assign n56993 = n30146 | n30147;
  assign n56994 = n30148 | n30149;
  assign n56995 = n30153 | n30154;
  assign n56996 = n30155 | n30156;
  assign n56997 = n30157 | ~n30158;
  assign n56998 = n30160 | n30161;
  assign n56999 = n30162 | n30163;
  assign n57000 = n30164 | ~n30165;
  assign n57001 = n30171 | ~n30172;
  assign n57002 = n30176 | ~n30177;
  assign n57003 = n30189 | ~n30190;
  assign n57004 = n30216 | n30211 | n30215;
  assign n57005 = n30221 | n30222;
  assign n57006 = n30229 | n30230;
  assign n57007 = n30244 | n30245;
  assign n57008 = n30261 | n30262;
  assign n57009 = n30273 | n30274;
  assign n57010 = n30293 | n30285 | n30292;
  assign n57011 = n30316 | n30317;
  assign n57012 = n30321 | ~n30322;
  assign n57013 = n30331 | n30332;
  assign n57014 = n30349 | n30350;
  assign n57015 = n30370 | n30361 | n30369;
  assign n57016 = n30385 | n30386;
  assign n57017 = n30390 | ~n30391;
  assign n57018 = n30400 | n30401;
  assign n57019 = n30411 | n30407 | n30410;
  assign n57020 = n30424 | n30420 | n30423;
  assign n57021 = n30429 | n30430;
  assign n57022 = n30448 | n30440 | n30447;
  assign n57023 = n30468 | n30465 | n30467;
  assign n57024 = n30479 | n30480;
  assign n57025 = n30505 | n30511 | n30521 | n30522;
  assign n57026 = n30531 | n30528 | n30530;
  assign n57027 = n30546 | n30557 | n30567 | n30568;
  assign n57028 = n30580 | n30581;
  assign n57029 = n30592 | n30588 | n30591;
  assign n57030 = n30606 | n30598 | n30605;
  assign n57031 = n30611 | n30612;
  assign n57032 = n30635 | n30632 | n30634;
  assign n57033 = n30639 | ~n30640;
  assign n57034 = n30649 | n30650;
  assign n57035 = n30660 | n30656 | n30659;
  assign n57036 = n30663 | n30664;
  assign n57037 = n30675 | n30676;
  assign n57038 = n30692 | n30693;
  assign n57039 = n30716 | n30705 | n30715;
  assign n57040 = n30720 | n30721;
  assign n57041 = n30735 | n30736;
  assign n57042 = n30740 | ~n30741;
  assign n57043 = n30750 | n30751;
  assign n57044 = n30761 | n30762;
  assign n57045 = n30775 | n30785 | n30795 | n30796;
  assign n57046 = n30799 | n30800;
  assign n57047 = n30805 | n30806;
  assign n57048 = n30821 | n30822;
  assign n57049 = n30825 | n30826;
  assign n57050 = n30839 | n30840;
  assign n57051 = n30844 | n30845;
  assign n57052 = n30848 | n30849;
  assign n57053 = n30850 | n30851;
  assign n57054 = n30863 | n30864;
  assign n57055 = n30875 | n30876;
  assign n57056 = n30882 | n30883;
  assign n57057 = n30892 | n30888 | n30891;
  assign n57058 = n30912 | n30913;
  assign n57059 = n30924 | n30925;
  assign n57060 = n30931 | n30932;
  assign n57061 = n30939 | n30940;
  assign n57062 = n30946 | n30947;
  assign n57063 = n30952 | n30953;
  assign n57064 = n30962 | n30958 | n30961;
  assign n57065 = n30977 | n30978;
  assign n57066 = n30981 | n30982;
  assign n57067 = n30987 | n30988;
  assign n57068 = n30998 | n30994 | n30997;
  assign n57069 = n31015 | n31016;
  assign n57070 = n31025 | n31026;
  assign n57071 = n31036 | n31037;
  assign n57072 = n31044 | n31045;
  assign n57073 = n31056 | n31064 | n31071 | n31072;
  assign n57074 = n31084 | n31085;
  assign n57075 = n31094 | n31095;
  assign n57076 = n31114 | n31101 | n31113;
  assign n57077 = n31134 | n31135;
  assign n57078 = n31151 | n31152;
  assign n57079 = n31154 | n31155;
  assign n57080 = n31156 | n31157;
  assign n57081 = n31158 | ~n31159;
  assign n57082 = n31163 | n31164;
  assign n57083 = n31165 | n31166;
  assign n57084 = n31167 | ~n31168;
  assign n57085 = n31172 | n31173;
  assign n57086 = n31174 | n31175;
  assign n57087 = n31176 | ~n31177;
  assign n57088 = n31181 | n31182;
  assign n57089 = n31183 | n31184;
  assign n57090 = n31185 | ~n31186;
  assign n57091 = n31190 | n31191;
  assign n57092 = n31192 | n31193;
  assign n57093 = n31194 | ~n31195;
  assign n57094 = n31199 | n31200;
  assign n57095 = n31201 | n31202;
  assign n57096 = n31203 | ~n31204;
  assign n57097 = n31208 | n31209;
  assign n57098 = n31210 | n31211;
  assign n57099 = n31212 | ~n31213;
  assign n57100 = n31217 | n31218;
  assign n57101 = n31219 | n31220;
  assign n57102 = n31221 | ~n31222;
  assign n57103 = n31228 | ~n31229;
  assign n57104 = n31241 | ~n31242;
  assign n57105 = n31249 | n31250;
  assign n57106 = n31251 | n31252;
  assign n57107 = n31253 | ~n31254;
  assign n57108 = n31258 | n31259;
  assign n57109 = n31260 | n31261;
  assign n57110 = n31262 | ~n31263;
  assign n57111 = n31278 | n31279;
  assign n57112 = n31280 | n31281;
  assign n57113 = n31286 | n31287;
  assign n57114 = n31298 | n31299;
  assign n57115 = n31300 | n31301;
  assign n57116 = n31306 | n31307;
  assign n57117 = n31318 | n31319;
  assign n57118 = n31320 | n31321;
  assign n57119 = n31326 | n31327;
  assign n57120 = n31330 | n31331;
  assign n57121 = n31332 | n31333;
  assign n57122 = n31335 | ~n31336;
  assign n57123 = n31347 | n31348;
  assign n57124 = n31349 | n31350;
  assign n57125 = n31355 | n31356;
  assign n57126 = n31367 | n31368;
  assign n57127 = n31369 | n31370;
  assign n57128 = n31375 | n31376;
  assign n57129 = n31379 | n31380;
  assign n57130 = n31381 | n31382;
  assign n57131 = n31384 | ~n31385;
  assign n57132 = n31393 | n31390 | n31392;
  assign n57133 = n31396 | n31397;
  assign n57134 = n31398 | n31399;
  assign n57135 = n31404 | n31405;
  assign n57136 = n31414 | n31415;
  assign n57137 = n31418 | n31419;
  assign n57138 = n31420 | n31421;
  assign n57139 = n31426 | ~n31427;
  assign n57140 = n31438 | n31439;
  assign n57141 = n31440 | n31441;
  assign n57142 = n31445 | n31446;
  assign n57143 = n31447 | n31448;
  assign n57144 = n31449 | ~n31450;
  assign n57145 = n31454 | ~n31455;
  assign n57146 = n31464 | n31465;
  assign n57147 = n31466 | n31467;
  assign n57148 = n31472 | ~n31473;
  assign n57149 = n31485 | n31486;
  assign n57150 = n31487 | n31488;
  assign n57151 = n31497 | n31498;
  assign n57152 = n31501 | n31502;
  assign n57153 = n31503 | n31504;
  assign n57154 = n31507 | n31508;
  assign n57155 = n31509 | n31510;
  assign n57156 = n31511 | ~n31512;
  assign n57157 = n31518 | ~n31519;
  assign n57158 = n31525 | ~n31526;
  assign n57159 = n31537 | n31538;
  assign n57160 = n31539 | n31540;
  assign n57161 = n31545 | n31546;
  assign n57162 = n31557 | n31558;
  assign n57163 = n31559 | n31560;
  assign n57164 = n31565 | n31566;
  assign n57165 = n31572 | ~n31573;
  assign n57166 = n31584 | n31585;
  assign n57167 = n31586 | n31587;
  assign n57168 = n31592 | n31593;
  assign n57169 = n31604 | n31605;
  assign n57170 = n31606 | n31607;
  assign n57171 = n31612 | n31613;
  assign n57172 = n31618 | n31619;
  assign n57173 = n31620 | n31621;
  assign n57174 = n31622 | ~n31623;
  assign n57175 = n31629 | ~n31630;
  assign n57176 = n31644 | n31645;
  assign n57177 = n31646 | n31647;
  assign n57178 = n31651 | n31652;
  assign n57179 = n31653 | n31654;
  assign n57180 = n31655 | ~n31656;
  assign n57181 = n31660 | ~n31661;
  assign n57182 = n31672 | n31673;
  assign n57183 = n31674 | n31675;
  assign n57184 = n31679 | n31680;
  assign n57185 = n31681 | n31682;
  assign n57186 = n31683 | ~n31684;
  assign n57187 = n31695 | n31696;
  assign n57188 = n31697 | n31698;
  assign n57189 = n31707 | n31708;
  assign n57190 = n31711 | n31712;
  assign n57191 = n31713 | n31714;
  assign n57192 = n31717 | n31718;
  assign n57193 = n31719 | n31720;
  assign n57194 = n31721 | ~n31722;
  assign n57195 = n31726 | n31727;
  assign n57196 = n31728 | n31729;
  assign n57197 = n31730 | ~n31731;
  assign n57198 = n31742 | n31743;
  assign n57199 = n31744 | n31745;
  assign n57200 = n31750 | n31751;
  assign n57201 = n31754 | n31755;
  assign n57202 = n31756 | n31757;
  assign n57203 = n31759 | ~n31760;
  assign n57204 = n31771 | n31772;
  assign n57205 = n31773 | n31774;
  assign n57206 = n31779 | n31780;
  assign n57207 = n31791 | n31792;
  assign n57208 = n31793 | n31794;
  assign n57209 = n31799 | n31800;
  assign n57210 = n31803 | n31804;
  assign n57211 = n31805 | n31806;
  assign n57212 = n31808 | ~n31809;
  assign n57213 = n31820 | n31821;
  assign n57214 = n31822 | n31823;
  assign n57215 = n31828 | n31829;
  assign n57216 = n31835 | ~n31836;
  assign n57217 = n31840 | n31841;
  assign n57218 = n31846 | ~n31847;
  assign n57219 = n31858 | n31859;
  assign n57220 = n31860 | n31861;
  assign n57221 = n31865 | n31866;
  assign n57222 = n31867 | n31868;
  assign n57223 = n31869 | ~n31870;
  assign n57224 = n31874 | ~n31875;
  assign n57225 = n31886 | n31887;
  assign n57226 = n31888 | n31889;
  assign n57227 = n31893 | n31894;
  assign n57228 = n31895 | n31896;
  assign n57229 = n31897 | ~n31898;
  assign n57230 = n31902 | ~n31903;
  assign n57231 = n31905 | n31906;
  assign n57232 = n31907 | n31908;
  assign n57233 = n31909 | ~n31910;
  assign n57234 = n31919 | ~n31920;
  assign n57235 = n31927 | ~n31928;
  assign n57236 = n31938 | ~n31939;
  assign n57237 = n31946 | ~n31947;
  assign n57238 = n31957 | ~n31958;
  assign n57239 = n31965 | ~n31966;
  assign n57240 = n31976 | ~n31977;
  assign n57241 = n31984 | ~n31985;
  assign n57242 = n31995 | ~n31996;
  assign n57243 = n32003 | ~n32004;
  assign n57244 = n32014 | n32015;
  assign n57245 = n32016 | n32017;
  assign n57246 = n32022 | ~n32023;
  assign n57247 = n32033 | n32034;
  assign n57248 = n32035 | n32036;
  assign n57249 = n32041 | ~n32042;
  assign n57250 = n32052 | n32053;
  assign n57251 = n32054 | n32055;
  assign n57252 = n32060 | ~n32061;
  assign n57253 = n32071 | n32072;
  assign n57254 = n32073 | n32074;
  assign n57255 = n32079 | ~n32080;
  assign n57256 = n32090 | n32091;
  assign n57257 = n32092 | n32093;
  assign n57258 = n32096 | n32097;
  assign n57259 = n32098 | n32099;
  assign n57260 = n32100 | ~n32101;
  assign n57261 = n32115 | n32116;
  assign n57262 = n32125 | ~n32126;
  assign n57263 = n32130 | n32131;
  assign n57264 = n32141 | n32142;
  assign n57265 = n32143 | n32144;
  assign n57266 = n32149 | ~n32150;
  assign n57267 = n32156 | ~n32157;
  assign n57268 = n32163 | ~n32164;
  assign n57269 = n32168 | n32169;
  assign n57270 = n32170 | n32171;
  assign n57271 = n32172 | ~n32173;
  assign n57272 = n32177 | n32178;
  assign n57273 = n32179 | n32180;
  assign n57274 = n32181 | ~n32182;
  assign n57275 = n32186 | n32187;
  assign n57276 = n32188 | n32189;
  assign n57277 = n32190 | ~n32191;
  assign n57278 = n32226 | n32227;
  assign n57279 = n32228 | n32229;
  assign n57280 = n32234 | n32235;
  assign n57281 = n32246 | n32247;
  assign n57282 = n32248 | n32249;
  assign n57283 = n32254 | n32255;
  assign n57284 = n32266 | n32267;
  assign n57285 = n32268 | n32269;
  assign n57286 = n32274 | n32275;
  assign n57287 = n32281 | ~n32282;
  assign n57288 = n32293 | n32294;
  assign n57289 = n32295 | n32296;
  assign n57290 = n32301 | n32302;
  assign n57291 = n32313 | n32314;
  assign n57292 = n32315 | n32316;
  assign n57293 = n32321 | n32322;
  assign n57294 = n32328 | ~n32329;
  assign n57295 = n32337 | n32334 | n32336;
  assign n57296 = n32340 | n32341;
  assign n57297 = n32342 | n32343;
  assign n57298 = n32348 | n32349;
  assign n57299 = n32358 | n32359;
  assign n57300 = n32362 | n32363;
  assign n57301 = n32364 | n32365;
  assign n57302 = n32370 | ~n32371;
  assign n57303 = n32382 | n32383;
  assign n57304 = n32384 | n32385;
  assign n57305 = n32389 | n32390;
  assign n57306 = n32391 | n32392;
  assign n57307 = n32393 | ~n32394;
  assign n57308 = n32398 | ~n32399;
  assign n57309 = n32403 | ~n32404;
  assign n57310 = n32415 | ~n32416;
  assign n57311 = n32431 | ~n32432;
  assign n57312 = n32447 | ~n32448;
  assign n57313 = n32463 | ~n32464;
  assign n57314 = n32479 | ~n32480;
  assign n57315 = n32495 | ~n32496;
  assign n57316 = n32509 | n32510;
  assign n57317 = n32513 | ~n32514;
  assign n57318 = n32527 | n32528;
  assign n57319 = n32531 | ~n32532;
  assign n57320 = n32545 | n32546;
  assign n57321 = n32549 | ~n32550;
  assign n57322 = n32561 | n32562;
  assign n57323 = n32565 | ~n32566;
  assign n57324 = n32573 | ~n32574;
  assign n57325 = n32582 | n32583;
  assign n57326 = n32586 | n32587;
  assign n57327 = n32588 | n32589;
  assign n57328 = n32600 | n32601;
  assign n57329 = n32604 | n32605;
  assign n57330 = n32606 | n32607;
  assign n57331 = n32613 | n32614;
  assign n57332 = n32622 | n32623;
  assign n57333 = n32626 | ~n32627;
  assign n57334 = n32635 | n32636;
  assign n57335 = n32649 | n32650;
  assign n57336 = n32657 | n32658;
  assign n57337 = n32661 | ~n32662;
  assign n57338 = n32666 | n32667;
  assign n57339 = n32675 | n32676;
  assign n57340 = n32679 | n32680;
  assign n57341 = n32681 | n32682;
  assign n57342 = n32685 | n32686;
  assign n57343 = n32687 | n32688;
  assign n57344 = n32689 | ~n32690;
  assign n57345 = n32698 | n32699;
  assign n57346 = n32700 | n32701;
  assign n57347 = n32702 | ~n32703;
  assign n57348 = n32707 | n32708;
  assign n57349 = n32709 | n32710;
  assign n57350 = n32711 | ~n32712;
  assign n57351 = n32716 | n32717;
  assign n57352 = n32718 | n32719;
  assign n57353 = n32720 | ~n32721;
  assign n57354 = n32725 | n32726;
  assign n57355 = n32727 | n32728;
  assign n57356 = n32729 | ~n32730;
  assign n57357 = n32734 | n32735;
  assign n57358 = n32736 | n32737;
  assign n57359 = n32738 | ~n32739;
  assign n57360 = n32743 | n32744;
  assign n57361 = n32745 | n32746;
  assign n57362 = n32747 | ~n32748;
  assign n57363 = n32752 | n32753;
  assign n57364 = n32754 | n32755;
  assign n57365 = n32756 | ~n32757;
  assign n57366 = n32761 | n32762;
  assign n57367 = n32763 | n32764;
  assign n57368 = n32765 | ~n32766;
  assign n57369 = n32770 | n32771;
  assign n57370 = n32772 | n32773;
  assign n57371 = n32774 | ~n32775;
  assign n57372 = n32779 | n32780;
  assign n57373 = n32781 | n32782;
  assign n57374 = n32783 | ~n32784;
  assign n57375 = n32788 | n32789;
  assign n57376 = n32790 | n32791;
  assign n57377 = n32792 | ~n32793;
  assign n57378 = n32803 | ~n32804;
  assign n57379 = n32815 | n32816;
  assign n57380 = n32817 | n32818;
  assign n57381 = n32823 | n32824;
  assign n57382 = n32835 | n32836;
  assign n57383 = n32837 | n32838;
  assign n57384 = n32843 | n32844;
  assign n57385 = n32855 | n32856;
  assign n57386 = n32857 | n32858;
  assign n57387 = n32863 | n32864;
  assign n57388 = n32867 | n32868;
  assign n57389 = n32869 | n32870;
  assign n57390 = n32872 | ~n32873;
  assign n57391 = n32884 | n32885;
  assign n57392 = n32886 | n32887;
  assign n57393 = n32892 | n32893;
  assign n57394 = n32904 | n32905;
  assign n57395 = n32906 | n32907;
  assign n57396 = n32912 | n32913;
  assign n57397 = n32918 | n32919;
  assign n57398 = n32920 | n32921;
  assign n57399 = n32922 | ~n32923;
  assign n57400 = n32926 | n32927;
  assign n57401 = n32928 | n32929;
  assign n57402 = n32931 | ~n32932;
  assign n57403 = n32946 | n32947;
  assign n57404 = n32948 | n32949;
  assign n57405 = n32953 | n32954;
  assign n57406 = n32955 | n32956;
  assign n57407 = n32957 | ~n32958;
  assign n57408 = n32962 | ~n32963;
  assign n57409 = n32967 | ~n32968;
  assign n57410 = n32977 | n32978;
  assign n57411 = n32979 | n32980;
  assign n57412 = n32993 | n32994;
  assign n57413 = n32995 | n32996;
  assign n57414 = n33001 | ~n33002;
  assign n57415 = n33012 | n33013;
  assign n57416 = n33014 | n33015;
  assign n57417 = n33020 | ~n33021;
  assign n57418 = n33031 | n33032;
  assign n57419 = n33033 | n33034;
  assign n57420 = n33039 | ~n33040;
  assign n57421 = n33050 | n33051;
  assign n57422 = n33052 | n33053;
  assign n57423 = n33058 | ~n33059;
  assign n57424 = n33069 | n33070;
  assign n57425 = n33071 | n33072;
  assign n57426 = n33075 | n33076;
  assign n57427 = n33077 | n33078;
  assign n57428 = n33079 | ~n33080;
  assign n57429 = n33090 | n33091;
  assign n57430 = n33092 | n33093;
  assign n57431 = n33096 | n33097;
  assign n57432 = n33098 | n33099;
  assign n57433 = n33100 | ~n33101;
  assign n57434 = n33111 | n33112;
  assign n57435 = n33113 | n33114;
  assign n57436 = n33117 | n33118;
  assign n57437 = n33119 | n33120;
  assign n57438 = n33121 | ~n33122;
  assign n57439 = n33132 | n33133;
  assign n57440 = n33134 | n33135;
  assign n57441 = n33140 | ~n33141;
  assign n57442 = n33151 | n33152;
  assign n57443 = n33153 | n33154;
  assign n57444 = n33159 | ~n33160;
  assign n57445 = n33172 | ~n33173;
  assign n57446 = n33188 | ~n33189;
  assign n57447 = n33202 | n33203;
  assign n57448 = n33204 | n33205;
  assign n57449 = n33218 | ~n33219;
  assign n57450 = n33226 | ~n33227;
  assign n57451 = n33237 | n33238;
  assign n57452 = n33239 | n33240;
  assign n57453 = n33246 | n33247;
  assign n57454 = n33257 | ~n33258;
  assign n57455 = n33266 | n33267;
  assign n57456 = n33280 | n33281;
  assign n57457 = n33290 | ~n33291;
  assign n57458 = n33295 | n33296;
  assign n57459 = n33306 | n33307;
  assign n57460 = n33308 | n33309;
  assign n57461 = n33312 | n33313;
  assign n57462 = n33314 | n33315;
  assign n57463 = n33316 | ~n33317;
  assign n57464 = n33325 | n33326;
  assign n57465 = n33327 | n33328;
  assign n57466 = n33329 | ~n33330;
  assign n57467 = n33338 | n33339;
  assign n57468 = n33340 | n33341;
  assign n57469 = n33342 | ~n33343;
  assign n57470 = n33347 | n33348;
  assign n57471 = n33349 | n33350;
  assign n57472 = n33351 | ~n33352;
  assign n57473 = n33360 | n33361;
  assign n57474 = n33362 | n33363;
  assign n57475 = n33364 | ~n33365;
  assign n57476 = n33369 | n33370;
  assign n57477 = n33371 | n33372;
  assign n57478 = n33373 | ~n33374;
  assign n57479 = n33380 | ~n33381;
  assign n57480 = n33387 | ~n33388;
  assign n57481 = n33394 | ~n33395;
  assign n57482 = n33399 | n33400;
  assign n57483 = n33401 | n33402;
  assign n57484 = n33403 | ~n33404;
  assign n57485 = n33408 | n33409;
  assign n57486 = n33410 | n33411;
  assign n57487 = n33412 | ~n33413;
  assign n57488 = n33417 | n33418;
  assign n57489 = n33419 | n33420;
  assign n57490 = n33421 | ~n33422;
  assign n57491 = n33426 | n33427;
  assign n57492 = n33428 | n33429;
  assign n57493 = n33430 | ~n33431;
  assign n57494 = n33435 | n33436;
  assign n57495 = n33437 | n33438;
  assign n57496 = n33439 | ~n33440;
  assign n57497 = n33443 | n33444;
  assign n57498 = n33445 | n33446;
  assign n57499 = n33448 | ~n33449;
  assign n57500 = n33460 | n33461;
  assign n57501 = n33462 | n33463;
  assign n57502 = n33468 | n33469;
  assign n57503 = n33480 | n33481;
  assign n57504 = n33482 | n33483;
  assign n57505 = n33488 | n33489;
  assign n57506 = n33500 | n33501;
  assign n57507 = n33502 | n33503;
  assign n57508 = n33508 | n33509;
  assign n57509 = n33515 | ~n33516;
  assign n57510 = n33527 | n33528;
  assign n57511 = n33529 | n33530;
  assign n57512 = n33535 | n33536;
  assign n57513 = n33542 | ~n33543;
  assign n57514 = n33547 | n33548;
  assign n57515 = n33553 | ~n33554;
  assign n57516 = n33565 | n33566;
  assign n57517 = n33567 | n33568;
  assign n57518 = n33572 | n33573;
  assign n57519 = n33574 | n33575;
  assign n57520 = n33576 | ~n33577;
  assign n57521 = n33581 | ~n33582;
  assign n57522 = n33586 | ~n33587;
  assign n57523 = n33598 | ~n33599;
  assign n57524 = n33614 | ~n33615;
  assign n57525 = n33630 | ~n33631;
  assign n57526 = n33646 | ~n33647;
  assign n57527 = n33662 | ~n33663;
  assign n57528 = n33678 | ~n33679;
  assign n57529 = n33694 | ~n33695;
  assign n57530 = n33710 | ~n33711;
  assign n57531 = n33726 | ~n33727;
  assign n57532 = n33742 | ~n33743;
  assign n57533 = n33756 | n33757;
  assign n57534 = n33758 | n33759;
  assign n57535 = n33772 | n33773;
  assign n57536 = n33774 | n33775;
  assign n57537 = n33778 | n33779;
  assign n57538 = n33780 | n33781;
  assign n57539 = n33782 | ~n33783;
  assign n57540 = n33795 | ~n33796;
  assign n57541 = n33811 | ~n33812;
  assign n57542 = n33827 | ~n33828;
  assign n57543 = n33841 | n33842;
  assign n57544 = n33843 | n33844;
  assign n57545 = n33857 | ~n33858;
  assign n57546 = n33865 | ~n33866;
  assign n57547 = n33876 | n33877;
  assign n57548 = n33878 | n33879;
  assign n57549 = n33885 | n33886;
  assign n57550 = n33896 | ~n33897;
  assign n57551 = n33905 | n33906;
  assign n57552 = n33919 | n33920;
  assign n57553 = n33929 | ~n33930;
  assign n57554 = n33934 | n33935;
  assign n57555 = n33945 | n33946;
  assign n57556 = n33947 | n33948;
  assign n57557 = n33951 | n33952;
  assign n57558 = n33953 | n33954;
  assign n57559 = n33955 | ~n33956;
  assign n57560 = n33964 | n33965;
  assign n57561 = n33966 | n33967;
  assign n57562 = n33968 | ~n33969;
  assign n57563 = n33977 | n33978;
  assign n57564 = n33979 | n33980;
  assign n57565 = n33981 | ~n33982;
  assign n57566 = n33986 | n33987;
  assign n57567 = n33988 | n33989;
  assign n57568 = n33990 | ~n33991;
  assign n57569 = n33995 | n33996;
  assign n57570 = n33997 | n33998;
  assign n57571 = n33999 | ~n34000;
  assign n57572 = n34010 | ~n34011;
  assign n57573 = n34015 | n34016;
  assign n57574 = n34017 | n34018;
  assign n57575 = n34019 | ~n34020;
  assign n57576 = n34024 | n34025;
  assign n57577 = n34026 | n34027;
  assign n57578 = n34028 | ~n34029;
  assign n57579 = n34033 | n34034;
  assign n57580 = n34035 | n34036;
  assign n57581 = n34037 | ~n34038;
  assign n57582 = n34042 | n34043;
  assign n57583 = n34044 | n34045;
  assign n57584 = n34046 | ~n34047;
  assign n57585 = n34051 | n34052;
  assign n57586 = n34053 | n34054;
  assign n57587 = n34055 | ~n34056;
  assign n57588 = n34060 | n34061;
  assign n57589 = n34062 | n34063;
  assign n57590 = n34064 | ~n34065;
  assign n57591 = n34069 | n34070;
  assign n57592 = n34071 | n34072;
  assign n57593 = n34073 | ~n34074;
  assign n57594 = n34078 | n34079;
  assign n57595 = n34080 | n34081;
  assign n57596 = n34082 | ~n34083;
  assign n57597 = n34087 | n34088;
  assign n57598 = n34089 | n34090;
  assign n57599 = n34091 | ~n34092;
  assign n57600 = n34096 | n34097;
  assign n57601 = n34098 | n34099;
  assign n57602 = n34100 | ~n34101;
  assign n57603 = n34111 | ~n34112;
  assign n57604 = n34123 | n34124;
  assign n57605 = n34125 | n34126;
  assign n57606 = n34131 | n34132;
  assign n57607 = n34143 | n34144;
  assign n57608 = n34145 | n34146;
  assign n57609 = n34151 | n34152;
  assign n57610 = n34163 | n34164;
  assign n57611 = n34165 | n34166;
  assign n57612 = n34171 | n34172;
  assign n57613 = n34175 | n34176;
  assign n57614 = n34177 | n34178;
  assign n57615 = n34180 | ~n34181;
  assign n57616 = n34189 | n34186 | n34188;
  assign n57617 = n34192 | n34193;
  assign n57618 = n34194 | n34195;
  assign n57619 = n34200 | n34201;
  assign n57620 = n34210 | n34211;
  assign n57621 = n34214 | n34215;
  assign n57622 = n34216 | n34217;
  assign n57623 = n34222 | ~n34223;
  assign n57624 = n34227 | ~n34228;
  assign n57625 = n34237 | n34238;
  assign n57626 = n34239 | n34240;
  assign n57627 = n34253 | n34254;
  assign n57628 = n34255 | n34256;
  assign n57629 = n34259 | n34260;
  assign n57630 = n34261 | n34262;
  assign n57631 = n34263 | ~n34264;
  assign n57632 = n34274 | n34275;
  assign n57633 = n34276 | n34277;
  assign n57634 = n34280 | n34281;
  assign n57635 = n34282 | n34283;
  assign n57636 = n34284 | ~n34285;
  assign n57637 = n34295 | n34296;
  assign n57638 = n34297 | n34298;
  assign n57639 = n34301 | n34302;
  assign n57640 = n34303 | n34304;
  assign n57641 = n34305 | ~n34306;
  assign n57642 = n34316 | n34317;
  assign n57643 = n34318 | n34319;
  assign n57644 = n34322 | n34323;
  assign n57645 = n34324 | n34325;
  assign n57646 = n34326 | ~n34327;
  assign n57647 = n34337 | n34338;
  assign n57648 = n34339 | n34340;
  assign n57649 = n34345 | ~n34346;
  assign n57650 = n34356 | n34357;
  assign n57651 = n34358 | n34359;
  assign n57652 = n34364 | ~n34365;
  assign n57653 = n34375 | n34376;
  assign n57654 = n34377 | n34378;
  assign n57655 = n34383 | ~n34384;
  assign n57656 = n34394 | n34395;
  assign n57657 = n34396 | n34397;
  assign n57658 = n34400 | n34401;
  assign n57659 = n34402 | n34403;
  assign n57660 = n34404 | ~n34405;
  assign n57661 = n34415 | n34416;
  assign n57662 = n34417 | n34418;
  assign n57663 = n34421 | n34422;
  assign n57664 = n34423 | n34424;
  assign n57665 = n34425 | ~n34426;
  assign n57666 = n34438 | ~n34439;
  assign n57667 = n34454 | ~n34455;
  assign n57668 = n34468 | n34469;
  assign n57669 = n34470 | n34471;
  assign n57670 = n34484 | n34485;
  assign n57671 = n34486 | n34487;
  assign n57672 = n34492 | ~n34493;
  assign n57673 = n34503 | n34504;
  assign n57674 = n34505 | n34506;
  assign n57675 = n34509 | n34510;
  assign n57676 = n34511 | n34512;
  assign n57677 = n34513 | ~n34514;
  assign n57678 = n34526 | ~n34527;
  assign n57679 = n34542 | ~n34543;
  assign n57680 = n34558 | ~n34559;
  assign n57681 = n34572 | n34573;
  assign n57682 = n34574 | n34575;
  assign n57683 = n34588 | ~n34589;
  assign n57684 = n34596 | ~n34597;
  assign n57685 = n34607 | n34608;
  assign n57686 = n34609 | n34610;
  assign n57687 = n34616 | n34617;
  assign n57688 = n34627 | ~n34628;
  assign n57689 = n34636 | n34637;
  assign n57690 = n34650 | n34651;
  assign n57691 = n34660 | ~n34661;
  assign n57692 = n34665 | n34666;
  assign n57693 = n34676 | n34677;
  assign n57694 = n34678 | n34679;
  assign n57695 = n34682 | n34683;
  assign n57696 = n34684 | n34685;
  assign n57697 = n34686 | ~n34687;
  assign n57698 = n34695 | n34696;
  assign n57699 = n34697 | n34698;
  assign n57700 = n34699 | ~n34700;
  assign n57701 = n34708 | n34709;
  assign n57702 = n34710 | n34711;
  assign n57703 = n34712 | ~n34713;
  assign n57704 = n34717 | n34718;
  assign n57705 = n34719 | n34720;
  assign n57706 = n34721 | ~n34722;
  assign n57707 = n34726 | n34727;
  assign n57708 = n34728 | n34729;
  assign n57709 = n34730 | ~n34731;
  assign n57710 = n34741 | ~n34742;
  assign n57711 = n34746 | n34747;
  assign n57712 = n34748 | n34749;
  assign n57713 = n34750 | ~n34751;
  assign n57714 = n34755 | n34756;
  assign n57715 = n34757 | n34758;
  assign n57716 = n34759 | ~n34760;
  assign n57717 = n34764 | n34765;
  assign n57718 = n34766 | n34767;
  assign n57719 = n34768 | ~n34769;
  assign n57720 = n34779 | ~n34780;
  assign n57721 = n34786 | ~n34787;
  assign n57722 = n34791 | n34792;
  assign n57723 = n34793 | n34794;
  assign n57724 = n34795 | ~n34796;
  assign n57725 = n34800 | n34801;
  assign n57726 = n34802 | n34803;
  assign n57727 = n34804 | ~n34805;
  assign n57728 = n34809 | n34810;
  assign n57729 = n34811 | n34812;
  assign n57730 = n34813 | ~n34814;
  assign n57731 = n34820 | ~n34821;
  assign n57732 = n34827 | ~n34828;
  assign n57733 = n34834 | ~n34835;
  assign n57734 = n34841 | ~n34842;
  assign n57735 = n34846 | n34847;
  assign n57736 = n34848 | n34849;
  assign n57737 = n34850 | ~n34851;
  assign n57738 = n34854 | n34855;
  assign n57739 = n34856 | n34857;
  assign n57740 = n34859 | ~n34860;
  assign n57741 = n34871 | n34872;
  assign n57742 = n34873 | n34874;
  assign n57743 = n34879 | n34880;
  assign n57744 = n34891 | n34892;
  assign n57745 = n34893 | n34894;
  assign n57746 = n34899 | n34900;
  assign n57747 = n34911 | n34912;
  assign n57748 = n34913 | n34914;
  assign n57749 = n34919 | n34920;
  assign n57750 = n34925 | n34926;
  assign n57751 = n34927 | n34928;
  assign n57752 = n34929 | ~n34930;
  assign n57753 = n34936 | ~n34937;
  assign n57754 = n34944 | ~n34945;
  assign n57755 = n34956 | ~n34957;
  assign n57756 = n34972 | ~n34973;
  assign n57757 = n34988 | ~n34989;
  assign n57758 = n35004 | ~n35005;
  assign n57759 = n35020 | ~n35021;
  assign n57760 = n35036 | ~n35037;
  assign n57761 = n35052 | ~n35053;
  assign n57762 = n35068 | ~n35069;
  assign n57763 = n35084 | ~n35085;
  assign n57764 = n35100 | ~n35101;
  assign n57765 = n35114 | n35115;
  assign n57766 = n35116 | n35117;
  assign n57767 = n35130 | n35131;
  assign n57768 = n35132 | n35133;
  assign n57769 = n35138 | ~n35139;
  assign n57770 = n35151 | ~n35152;
  assign n57771 = n35167 | ~n35168;
  assign n57772 = n35183 | ~n35184;
  assign n57773 = n35197 | n35198;
  assign n57774 = n35199 | n35200;
  assign n57775 = n35213 | n35214;
  assign n57776 = n35215 | n35216;
  assign n57777 = n35221 | ~n35222;
  assign n57778 = n35232 | n35233;
  assign n57779 = n35234 | n35235;
  assign n57780 = n35238 | n35239;
  assign n57781 = n35240 | n35241;
  assign n57782 = n35242 | ~n35243;
  assign n57783 = n35255 | ~n35256;
  assign n57784 = n35271 | ~n35272;
  assign n57785 = n35287 | ~n35288;
  assign n57786 = n35301 | n35302;
  assign n57787 = n35303 | n35304;
  assign n57788 = n35317 | ~n35318;
  assign n57789 = n35325 | ~n35326;
  assign n57790 = n35336 | n35337;
  assign n57791 = n35338 | n35339;
  assign n57792 = n35345 | n35346;
  assign n57793 = n35356 | ~n35357;
  assign n57794 = n35365 | n35366;
  assign n57795 = n35379 | n35380;
  assign n57796 = n35389 | ~n35390;
  assign n57797 = n35394 | n35395;
  assign n57798 = n35405 | n35406;
  assign n57799 = n35407 | n35408;
  assign n57800 = n35411 | n35412;
  assign n57801 = n35413 | n35414;
  assign n57802 = n35415 | ~n35416;
  assign n57803 = n35424 | n35425;
  assign n57804 = n35426 | n35427;
  assign n57805 = n35428 | ~n35429;
  assign n57806 = n35437 | n35438;
  assign n57807 = n35439 | n35440;
  assign n57808 = n35441 | ~n35442;
  assign n57809 = n35446 | n35447;
  assign n57810 = n35448 | n35449;
  assign n57811 = n35450 | ~n35451;
  assign n57812 = n35455 | n35456;
  assign n57813 = n35457 | n35458;
  assign n57814 = n35459 | ~n35460;
  assign n57815 = n35470 | ~n35471;
  assign n57816 = n35475 | n35476;
  assign n57817 = n35477 | n35478;
  assign n57818 = n35479 | ~n35480;
  assign n57819 = n35484 | n35485;
  assign n57820 = n35486 | n35487;
  assign n57821 = n35488 | ~n35489;
  assign n57822 = n35493 | n35494;
  assign n57823 = n35495 | n35496;
  assign n57824 = n35497 | ~n35498;
  assign n57825 = n35502 | n35503;
  assign n57826 = n35504 | n35505;
  assign n57827 = n35506 | ~n35507;
  assign n57828 = n35515 | n35516;
  assign n57829 = n35517 | n35518;
  assign n57830 = n35519 | ~n35520;
  assign n57831 = n35524 | n35525;
  assign n57832 = n35526 | n35527;
  assign n57833 = n35528 | ~n35529;
  assign n57834 = n35533 | n35534;
  assign n57835 = n35535 | n35536;
  assign n57836 = n35537 | ~n35538;
  assign n57837 = n35542 | n35543;
  assign n57838 = n35544 | n35545;
  assign n57839 = n35546 | ~n35547;
  assign n57840 = n35551 | n35552;
  assign n57841 = n35553 | n35554;
  assign n57842 = n35555 | ~n35556;
  assign n57843 = n35560 | n35561;
  assign n57844 = n35562 | n35563;
  assign n57845 = n35564 | ~n35565;
  assign n57846 = n35569 | n35570;
  assign n57847 = n35571 | n35572;
  assign n57848 = n35573 | ~n35574;
  assign n57849 = n35578 | n35579;
  assign n57850 = n35580 | n35581;
  assign n57851 = n35582 | ~n35583;
  assign n57852 = n35587 | n35588;
  assign n57853 = n35589 | n35590;
  assign n57854 = n35591 | ~n35592;
  assign n57855 = n35596 | n35597;
  assign n57856 = n35598 | n35599;
  assign n57857 = n35600 | ~n35601;
  assign n57858 = n35605 | n35606;
  assign n57859 = n35607 | n35608;
  assign n57860 = n35609 | ~n35610;
  assign n57861 = n35620 | ~n35621;
  assign n57862 = n35632 | n35633;
  assign n57863 = n35634 | n35635;
  assign n57864 = n35640 | n35641;
  assign n57865 = n35652 | n35653;
  assign n57866 = n35654 | n35655;
  assign n57867 = n35660 | n35661;
  assign n57868 = n35667 | ~n35668;
  assign n57869 = n35672 | n35673;
  assign n57870 = n35678 | ~n35679;
  assign n57871 = n35683 | ~n35684;
  assign n57872 = n35693 | n35694;
  assign n57873 = n35695 | n35696;
  assign n57874 = n35709 | n35710;
  assign n57875 = n35711 | n35712;
  assign n57876 = n35717 | ~n35718;
  assign n57877 = n35728 | n35729;
  assign n57878 = n35730 | n35731;
  assign n57879 = n35736 | ~n35737;
  assign n57880 = n35747 | n35748;
  assign n57881 = n35749 | n35750;
  assign n57882 = n35755 | ~n35756;
  assign n57883 = n35766 | n35767;
  assign n57884 = n35768 | n35769;
  assign n57885 = n35774 | ~n35775;
  assign n57886 = n35785 | n35786;
  assign n57887 = n35787 | n35788;
  assign n57888 = n35791 | n35792;
  assign n57889 = n35793 | n35794;
  assign n57890 = n35795 | ~n35796;
  assign n57891 = n35806 | n35807;
  assign n57892 = n35808 | n35809;
  assign n57893 = n35812 | n35813;
  assign n57894 = n35814 | n35815;
  assign n57895 = n35816 | ~n35817;
  assign n57896 = n35827 | n35828;
  assign n57897 = n35829 | n35830;
  assign n57898 = n35833 | n35834;
  assign n57899 = n35835 | n35836;
  assign n57900 = n35837 | ~n35838;
  assign n57901 = n35848 | n35849;
  assign n57902 = n35850 | n35851;
  assign n57903 = n35856 | ~n35857;
  assign n57904 = n35867 | n35868;
  assign n57905 = n35869 | n35870;
  assign n57906 = n35875 | ~n35876;
  assign n57907 = n35888 | ~n35889;
  assign n57908 = n35904 | ~n35905;
  assign n57909 = n35918 | n35919;
  assign n57910 = n35920 | n35921;
  assign n57911 = n35934 | n35935;
  assign n57912 = n35936 | n35937;
  assign n57913 = n35940 | n35941;
  assign n57914 = n35942 | n35943;
  assign n57915 = n35944 | ~n35945;
  assign n57916 = n35955 | n35956;
  assign n57917 = n35957 | n35958;
  assign n57918 = n35963 | ~n35964;
  assign n57919 = n35976 | ~n35977;
  assign n57920 = n35992 | ~n35993;
  assign n57921 = n36008 | ~n36009;
  assign n57922 = n36022 | n36023;
  assign n57923 = n36024 | n36025;
  assign n57924 = n36038 | n36039;
  assign n57925 = n36040 | n36041;
  assign n57926 = n36046 | ~n36047;
  assign n57927 = n36057 | n36058;
  assign n57928 = n36059 | n36060;
  assign n57929 = n36063 | n36064;
  assign n57930 = n36065 | n36066;
  assign n57931 = n36067 | ~n36068;
  assign n57932 = n36080 | ~n36081;
  assign n57933 = n36096 | ~n36097;
  assign n57934 = n36112 | ~n36113;
  assign n57935 = n36126 | n36127;
  assign n57936 = n36128 | n36129;
  assign n57937 = n36142 | ~n36143;
  assign n57938 = n36150 | ~n36151;
  assign n57939 = n36161 | n36162;
  assign n57940 = n36163 | n36164;
  assign n57941 = n36170 | n36171;
  assign n57942 = n36181 | ~n36182;
  assign n57943 = n36190 | n36191;
  assign n57944 = n36204 | n36205;
  assign n57945 = n36214 | ~n36215;
  assign n57946 = n36219 | n36220;
  assign n57947 = n36230 | n36231;
  assign n57948 = n36232 | n36233;
  assign n57949 = n36236 | n36237;
  assign n57950 = n36238 | n36239;
  assign n57951 = n36240 | ~n36241;
  assign n57952 = n36249 | n36250;
  assign n57953 = n36251 | n36252;
  assign n57954 = n36253 | ~n36254;
  assign n57955 = n36262 | n36263;
  assign n57956 = n36264 | n36265;
  assign n57957 = n36266 | ~n36267;
  assign n57958 = n36271 | n36272;
  assign n57959 = n36273 | n36274;
  assign n57960 = n36275 | ~n36276;
  assign n57961 = n36280 | n36281;
  assign n57962 = n36282 | n36283;
  assign n57963 = n36284 | ~n36285;
  assign n57964 = n36295 | ~n36296;
  assign n57965 = n36300 | n36301;
  assign n57966 = n36302 | n36303;
  assign n57967 = n36304 | ~n36305;
  assign n57968 = n36309 | n36310;
  assign n57969 = n36311 | n36312;
  assign n57970 = n36313 | ~n36314;
  assign n57971 = n36318 | n36319;
  assign n57972 = n36320 | n36321;
  assign n57973 = n36322 | ~n36323;
  assign n57974 = n36327 | n36328;
  assign n57975 = n36329 | n36330;
  assign n57976 = n36331 | ~n36332;
  assign n57977 = n36340 | n36341;
  assign n57978 = n36342 | n36343;
  assign n57979 = n36344 | ~n36345;
  assign n57980 = n36351 | ~n36352;
  assign n57981 = n36356 | n36357;
  assign n57982 = n36358 | n36359;
  assign n57983 = n36360 | ~n36361;
  assign n57984 = n36365 | n36366;
  assign n57985 = n36367 | n36368;
  assign n57986 = n36369 | ~n36370;
  assign n57987 = n36378 | n36379;
  assign n57988 = n36380 | n36381;
  assign n57989 = n36382 | ~n36383;
  assign n57990 = n36387 | n36388;
  assign n57991 = n36389 | n36390;
  assign n57992 = n36391 | ~n36392;
  assign n57993 = n36398 | ~n36399;
  assign n57994 = n36405 | ~n36406;
  assign n57995 = n36412 | ~n36413;
  assign n57996 = n36417 | n36418;
  assign n57997 = n36419 | n36420;
  assign n57998 = n36421 | ~n36422;
  assign n57999 = n36426 | n36427;
  assign n58000 = n36428 | n36429;
  assign n58001 = n36430 | ~n36431;
  assign n58002 = n36435 | n36436;
  assign n58003 = n36437 | n36438;
  assign n58004 = n36439 | ~n36440;
  assign n58005 = n36444 | n36445;
  assign n58006 = n36446 | n36447;
  assign n58007 = n36448 | ~n36449;
  assign n58008 = n36453 | n36454;
  assign n58009 = n36455 | n36456;
  assign n58010 = n36457 | ~n36458;
  assign n58011 = n36461 | n36462;
  assign n58012 = n36463 | n36464;
  assign n58013 = n36466 | ~n36467;
  assign n58014 = n36478 | n36479;
  assign n58015 = n36480 | n36481;
  assign n58016 = n36486 | n36487;
  assign n58017 = n36495 | n36492 | n36494;
  assign n58018 = n36498 | n36499;
  assign n58019 = n36500 | n36501;
  assign n58020 = n36506 | n36507;
  assign n58021 = n36514 | ~n36515;
  assign n58022 = n36526 | ~n36527;
  assign n58023 = n36542 | ~n36543;
  assign n58024 = n36558 | ~n36559;
  assign n58025 = n36574 | ~n36575;
  assign n58026 = n36590 | ~n36591;
  assign n58027 = n36606 | ~n36607;
  assign n58028 = n36622 | ~n36623;
  assign n58029 = n36638 | ~n36639;
  assign n58030 = n36654 | ~n36655;
  assign n58031 = n36670 | ~n36671;
  assign n58032 = n36684 | n36685;
  assign n58033 = n36686 | n36687;
  assign n58034 = n36700 | n36701;
  assign n58035 = n36702 | n36703;
  assign n58036 = n36706 | n36707;
  assign n58037 = n36708 | n36709;
  assign n58038 = n36710 | ~n36711;
  assign n58039 = n36723 | ~n36724;
  assign n58040 = n36739 | ~n36740;
  assign n58041 = n36755 | ~n36756;
  assign n58042 = n36769 | n36770;
  assign n58043 = n36771 | n36772;
  assign n58044 = n36785 | n36786;
  assign n58045 = n36787 | n36788;
  assign n58046 = n36791 | n36792;
  assign n58047 = n36793 | n36794;
  assign n58048 = n36795 | ~n36796;
  assign n58049 = n36806 | n36807;
  assign n58050 = n36808 | n36809;
  assign n58051 = n36814 | ~n36815;
  assign n58052 = n36827 | ~n36828;
  assign n58053 = n36843 | ~n36844;
  assign n58054 = n36859 | ~n36860;
  assign n58055 = n36873 | n36874;
  assign n58056 = n36875 | n36876;
  assign n58057 = n36889 | n36890;
  assign n58058 = n36891 | n36892;
  assign n58059 = n36897 | ~n36898;
  assign n58060 = n36908 | n36909;
  assign n58061 = n36910 | n36911;
  assign n58062 = n36914 | n36915;
  assign n58063 = n36916 | n36917;
  assign n58064 = n36918 | ~n36919;
  assign n58065 = n36931 | ~n36932;
  assign n58066 = n36947 | ~n36948;
  assign n58067 = n36963 | ~n36964;
  assign n58068 = n36977 | n36978;
  assign n58069 = n36979 | n36980;
  assign n58070 = n36993 | ~n36994;
  assign n58071 = n37001 | ~n37002;
  assign n58072 = n37012 | n37013;
  assign n58073 = n37014 | n37015;
  assign n58074 = n37021 | n37022;
  assign n58075 = n37032 | ~n37033;
  assign n58076 = n37041 | n37042;
  assign n58077 = n37055 | n37056;
  assign n58078 = n37065 | ~n37066;
  assign n58079 = n37070 | n37071;
  assign n58080 = n37081 | n37082;
  assign n58081 = n37083 | n37084;
  assign n58082 = n37087 | n37088;
  assign n58083 = n37089 | n37090;
  assign n58084 = n37091 | ~n37092;
  assign n58085 = n37100 | n37101;
  assign n58086 = n37102 | n37103;
  assign n58087 = n37104 | ~n37105;
  assign n58088 = n37113 | n37114;
  assign n58089 = n37115 | n37116;
  assign n58090 = n37117 | ~n37118;
  assign n58091 = n37122 | n37123;
  assign n58092 = n37124 | n37125;
  assign n58093 = n37126 | ~n37127;
  assign n58094 = n37131 | n37132;
  assign n58095 = n37133 | n37134;
  assign n58096 = n37135 | ~n37136;
  assign n58097 = n37146 | ~n37147;
  assign n58098 = n37151 | n37152;
  assign n58099 = n37153 | n37154;
  assign n58100 = n37155 | ~n37156;
  assign n58101 = n37160 | n37161;
  assign n58102 = n37162 | n37163;
  assign n58103 = n37164 | ~n37165;
  assign n58104 = n37169 | n37170;
  assign n58105 = n37171 | n37172;
  assign n58106 = n37173 | ~n37174;
  assign n58107 = n37178 | n37179;
  assign n58108 = n37180 | n37181;
  assign n58109 = n37182 | ~n37183;
  assign n58110 = n37191 | n37192;
  assign n58111 = n37193 | n37194;
  assign n58112 = n37195 | ~n37196;
  assign n58113 = n37202 | ~n37203;
  assign n58114 = n37207 | n37208;
  assign n58115 = n37209 | n37210;
  assign n58116 = n37211 | ~n37212;
  assign n58117 = n37216 | n37217;
  assign n58118 = n37218 | n37219;
  assign n58119 = n37220 | ~n37221;
  assign n58120 = n37225 | n37226;
  assign n58121 = n37227 | n37228;
  assign n58122 = n37229 | ~n37230;
  assign n58123 = n37240 | ~n37241;
  assign n58124 = n37245 | n37246;
  assign n58125 = n37247 | n37248;
  assign n58126 = n37249 | ~n37250;
  assign n58127 = n37254 | n37255;
  assign n58128 = n37256 | n37257;
  assign n58129 = n37258 | ~n37259;
  assign n58130 = n37263 | n37264;
  assign n58131 = n37265 | n37266;
  assign n58132 = n37267 | ~n37268;
  assign n58133 = n37272 | n37273;
  assign n58134 = n37274 | n37275;
  assign n58135 = n37276 | ~n37277;
  assign n58136 = n37281 | n37282;
  assign n58137 = n37283 | n37284;
  assign n58138 = n37285 | ~n37286;
  assign n58139 = n37290 | n37291;
  assign n58140 = n37292 | n37293;
  assign n58141 = n37294 | ~n37295;
  assign n58142 = n37299 | n37300;
  assign n58143 = n37301 | n37302;
  assign n58144 = n37303 | ~n37304;
  assign n58145 = n37308 | n37309;
  assign n58146 = n37310 | n37311;
  assign n58147 = n37312 | ~n37313;
  assign n58148 = n37317 | n37318;
  assign n58149 = n37319 | n37320;
  assign n58150 = n37321 | ~n37322;
  assign n58151 = n37326 | n37327;
  assign n58152 = n37328 | n37329;
  assign n58153 = n37330 | ~n37331;
  assign n58154 = n37341 | ~n37342;
  assign n58155 = n37350 | n37351;
  assign n58156 = n37354 | n37355;
  assign n58157 = n37356 | n37357;
  assign n58158 = n37362 | n37363;
  assign n58159 = n37375 | n37376;
  assign n58160 = n37377 | n37378;
  assign n58161 = n37384 | n37385;
  assign n58162 = n37386 | n37387;
  assign n58163 = n37388 | ~n37389;
  assign n58164 = n37392 | n37393;
  assign n58165 = n37394 | n37395;
  assign n58166 = n37397 | ~n37398;
  assign n58167 = n37410 | n37411;
  assign n58168 = n37412 | n37413;
  assign n58169 = n37416 | n37417;
  assign n58170 = n37418 | n37419;
  assign n58171 = n37420 | ~n37421;
  assign n58172 = n37431 | n37432;
  assign n58173 = n37433 | n37434;
  assign n58174 = n37437 | n37438;
  assign n58175 = n37439 | n37440;
  assign n58176 = n37441 | ~n37442;
  assign n58177 = n37452 | n37453;
  assign n58178 = n37454 | n37455;
  assign n58179 = n37458 | n37459;
  assign n58180 = n37460 | n37461;
  assign n58181 = n37462 | ~n37463;
  assign n58182 = n37473 | n37474;
  assign n58183 = n37475 | n37476;
  assign n58184 = n37479 | n37480;
  assign n58185 = n37481 | n37482;
  assign n58186 = n37483 | ~n37484;
  assign n58187 = n37494 | n37495;
  assign n58188 = n37496 | n37497;
  assign n58189 = n37502 | ~n37503;
  assign n58190 = n37513 | n37514;
  assign n58191 = n37515 | n37516;
  assign n58192 = n37521 | ~n37522;
  assign n58193 = n37532 | n37533;
  assign n58194 = n37534 | n37535;
  assign n58195 = n37540 | ~n37541;
  assign n58196 = n37551 | n37552;
  assign n58197 = n37553 | n37554;
  assign n58198 = n37557 | n37558;
  assign n58199 = n37559 | n37560;
  assign n58200 = n37561 | ~n37562;
  assign n58201 = n37572 | n37573;
  assign n58202 = n37574 | n37575;
  assign n58203 = n37578 | n37579;
  assign n58204 = n37580 | n37581;
  assign n58205 = n37582 | ~n37583;
  assign n58206 = n37595 | ~n37596;
  assign n58207 = n37611 | ~n37612;
  assign n58208 = n37625 | n37626;
  assign n58209 = n37627 | n37628;
  assign n58210 = n37641 | n37642;
  assign n58211 = n37643 | n37644;
  assign n58212 = n37649 | ~n37650;
  assign n58213 = n37660 | n37661;
  assign n58214 = n37662 | n37663;
  assign n58215 = n37666 | n37667;
  assign n58216 = n37668 | n37669;
  assign n58217 = n37670 | ~n37671;
  assign n58218 = n37683 | ~n37684;
  assign n58219 = n37699 | ~n37700;
  assign n58220 = n37715 | ~n37716;
  assign n58221 = n37729 | n37730;
  assign n58222 = n37731 | n37732;
  assign n58223 = n37745 | n37746;
  assign n58224 = n37747 | n37748;
  assign n58225 = n37751 | n37752;
  assign n58226 = n37753 | n37754;
  assign n58227 = n37755 | ~n37756;
  assign n58228 = n37766 | n37767;
  assign n58229 = n37768 | n37769;
  assign n58230 = n37774 | ~n37775;
  assign n58231 = n37787 | ~n37788;
  assign n58232 = n37803 | ~n37804;
  assign n58233 = n37819 | ~n37820;
  assign n58234 = n37833 | n37834;
  assign n58235 = n37835 | n37836;
  assign n58236 = n37849 | n37850;
  assign n58237 = n37851 | n37852;
  assign n58238 = n37857 | ~n37858;
  assign n58239 = n37868 | n37869;
  assign n58240 = n37870 | n37871;
  assign n58241 = n37874 | n37875;
  assign n58242 = n37876 | n37877;
  assign n58243 = n37878 | ~n37879;
  assign n58244 = n37891 | ~n37892;
  assign n58245 = n37907 | ~n37908;
  assign n58246 = n37923 | ~n37924;
  assign n58247 = n37937 | n37938;
  assign n58248 = n37939 | n37940;
  assign n58249 = n37953 | ~n37954;
  assign n58250 = n37961 | ~n37962;
  assign n58251 = n37972 | n37973;
  assign n58252 = n37974 | n37975;
  assign n58253 = n37981 | n37982;
  assign n58254 = n37992 | ~n37993;
  assign n58255 = n38001 | n38002;
  assign n58256 = n38015 | n38016;
  assign n58257 = n38025 | ~n38026;
  assign n58258 = n38030 | n38031;
  assign n58259 = n38041 | n38042;
  assign n58260 = n38043 | n38044;
  assign n58261 = n38047 | n38048;
  assign n58262 = n38049 | n38050;
  assign n58263 = n38051 | ~n38052;
  assign n58264 = n38060 | n38061;
  assign n58265 = n38062 | n38063;
  assign n58266 = n38064 | ~n38065;
  assign n58267 = n38073 | n38074;
  assign n58268 = n38075 | n38076;
  assign n58269 = n38077 | ~n38078;
  assign n58270 = n38082 | n38083;
  assign n58271 = n38084 | n38085;
  assign n58272 = n38086 | ~n38087;
  assign n58273 = n38091 | n38092;
  assign n58274 = n38093 | n38094;
  assign n58275 = n38095 | ~n38096;
  assign n58276 = n38106 | ~n38107;
  assign n58277 = n38111 | n38112;
  assign n58278 = n38113 | n38114;
  assign n58279 = n38115 | ~n38116;
  assign n58280 = n38120 | n38121;
  assign n58281 = n38122 | n38123;
  assign n58282 = n38124 | ~n38125;
  assign n58283 = n38129 | n38130;
  assign n58284 = n38131 | n38132;
  assign n58285 = n38133 | ~n38134;
  assign n58286 = n38138 | n38139;
  assign n58287 = n38140 | n38141;
  assign n58288 = n38142 | ~n38143;
  assign n58289 = n38151 | n38152;
  assign n58290 = n38153 | n38154;
  assign n58291 = n38155 | ~n38156;
  assign n58292 = n38162 | ~n38163;
  assign n58293 = n38167 | n38168;
  assign n58294 = n38169 | n38170;
  assign n58295 = n38171 | ~n38172;
  assign n58296 = n38176 | n38177;
  assign n58297 = n38178 | n38179;
  assign n58298 = n38180 | ~n38181;
  assign n58299 = n38185 | n38186;
  assign n58300 = n38187 | n38188;
  assign n58301 = n38189 | ~n38190;
  assign n58302 = n38200 | ~n38201;
  assign n58303 = n38205 | n38206;
  assign n58304 = n38207 | n38208;
  assign n58305 = n38209 | ~n38210;
  assign n58306 = n38214 | n38215;
  assign n58307 = n38216 | n38217;
  assign n58308 = n38218 | ~n38219;
  assign n58309 = n38223 | n38224;
  assign n58310 = n38225 | n38226;
  assign n58311 = n38227 | ~n38228;
  assign n58312 = n38238 | ~n38239;
  assign n58313 = n38245 | ~n38246;
  assign n58314 = n38250 | n38251;
  assign n58315 = n38252 | n38253;
  assign n58316 = n38254 | ~n38255;
  assign n58317 = n38259 | n38260;
  assign n58318 = n38261 | n38262;
  assign n58319 = n38263 | ~n38264;
  assign n58320 = n38268 | n38269;
  assign n58321 = n38270 | n38271;
  assign n58322 = n38272 | ~n38273;
  assign n58323 = n38279 | ~n38280;
  assign n58324 = n38286 | ~n38287;
  assign n58325 = n38293 | ~n38294;
  assign n58326 = n38300 | ~n38301;
  assign n58327 = n38307 | ~n38308;
  assign n58328 = n38324 | n38325;
  assign n58329 = n38328 | ~n38329;
  assign n58330 = n38344 | ~n38345;
  assign n58331 = n38360 | ~n38361;
  assign n58332 = n38376 | ~n38377;
  assign n58333 = n38392 | ~n38393;
  assign n58334 = n38408 | ~n38409;
  assign n58335 = n38424 | ~n38425;
  assign n58336 = n38440 | ~n38441;
  assign n58337 = n38447 | n38448;
  assign n58338 = n38449 | n38450;
  assign n58339 = n38451 | ~n38452;
  assign n58340 = n38456 | n38457;
  assign n58341 = n38471 | ~n38472;
  assign n58342 = n38481 | n38482;
  assign n58343 = n38485 | n38486;
  assign n58344 = n38500 | ~n38501;
  assign n58345 = n38510 | n38511;
  assign n58346 = n38514 | n38515;
  assign n58347 = n38529 | ~n38530;
  assign n58348 = n38539 | n38540;
  assign n58349 = n38543 | n38544;
  assign n58350 = n38558 | ~n38559;
  assign n58351 = n38575 | ~n38576;
  assign n58352 = n38588 | n38589;
  assign n58353 = n38601 | ~n38602;
  assign n58354 = n38612 | ~n38613;
  assign n58355 = n38639 | n38647 | n38649 | n38650;
  assign n58356 = n38642 | n38643;
  assign n58357 = n38663 | ~n38664;
  assign n58358 = n38672 | n38673;
  assign n58359 = n38681 | ~n38682;
  assign n58360 = n38687 | ~n38688;
  assign n58361 = n38702 | ~n38703;
  assign n58362 = n38710 | ~n38711;
  assign n58363 = n38713 | n38714;
  assign n58364 = n38718 | ~n38719;
  assign n58365 = n38730 | ~n38731;
  assign n58366 = n38739 | ~n38740;
  assign n58367 = n38751 | ~n38752;
  assign n58368 = n38760 | ~n38761;
  assign n58369 = n38775 | ~n38776;
  assign n58370 = n38791 | ~n38792;
  assign n58371 = n38808 | ~n38809;
  assign n58372 = n38818 | ~n38819;
  assign n58373 = n38821 | n38822;
  assign n58374 = n38826 | ~n38827;
  assign n58375 = n38838 | ~n38839;
  assign n58376 = n38847 | ~n38848;
  assign n58377 = n38859 | ~n38860;
  assign n58378 = n38868 | ~n38869;
  assign n58379 = n38883 | ~n38884;
  assign n58380 = n38899 | ~n38900;
  assign n58381 = n38916 | ~n38917;
  assign n58382 = n38926 | ~n38927;
  assign n58383 = n38929 | n38930;
  assign n58384 = n38934 | ~n38935;
  assign n58385 = n38946 | ~n38947;
  assign n58386 = n38955 | ~n38956;
  assign n58387 = n38967 | ~n38968;
  assign n58388 = n38976 | ~n38977;
  assign n58389 = n38991 | ~n38992;
  assign n58390 = n39007 | ~n39008;
  assign n58391 = n39024 | ~n39025;
  assign n58392 = n39034 | ~n39035;
  assign n58393 = n39037 | n39038;
  assign n58394 = n39042 | ~n39043;
  assign n58395 = n39054 | ~n39055;
  assign n58396 = n39063 | ~n39064;
  assign n58397 = n39075 | ~n39076;
  assign n58398 = n39084 | ~n39085;
  assign n58399 = n39099 | ~n39100;
  assign n58400 = n39116 | ~n39117;
  assign n58401 = n39167 | n39168;
  assign n58402 = n39169 | n39170;
  assign n58403 = n39171 | ~n39172;
  assign n58404 = n39182 | n39183;
  assign n58405 = n39184 | n39185;
  assign n58406 = n39186 | ~n39187;
  assign n58407 = n39197 | n39198;
  assign n58408 = n39199 | n39200;
  assign n58409 = n39201 | ~n39202;
  assign n58410 = n39212 | n39213;
  assign n58411 = n39214 | n39215;
  assign n58412 = n39216 | ~n39217;
  assign n58413 = n39227 | n39228;
  assign n58414 = n39229 | n39230;
  assign n58415 = n39231 | ~n39232;
  assign n58416 = n39246 | n39247;
  assign n58417 = n39248 | n39249;
  assign n58418 = n39259 | n39260;
  assign n58419 = n39261 | n39262;
  assign n58420 = n39279 | n39280;
  assign n58421 = n39291 | n39292;
  assign n58422 = n39308 | n39301 | n39307;
  assign n58423 = n39325 | n39326;
  assign n58424 = n39346 | n39335 | n39345;
  assign n58425 = n39365 | n39366;
  assign n58426 = n39380 | ~n39381;
  assign n58427 = n39386 | n39387;
  assign n58428 = n39388 | n39389;
  assign n58429 = n39391 | ~n39392;
  assign n58430 = n39395 | n39396;
  assign n58431 = n39397 | n39398;
  assign n58432 = n39399 | ~n39400;
  assign n58433 = n39409 | n39410;
  assign n58434 = n39413 | n39414;
  assign n58435 = n39415 | n39416;
  assign n58436 = n39419 | n39420;
  assign n58437 = n39423 | n39424;
  assign n58438 = n39425 | n39426;
  assign n58439 = n39427 | ~n39428;
  assign n58440 = n39433 | n39434;
  assign n58441 = n39449 | n39446 | n39448;
  assign n58442 = n39452 | n39453;
  assign n58443 = n39454 | n39455;
  assign n58444 = n39466 | n39467;
  assign n58445 = n39468 | n39469;
  assign n58446 = n39483 | n39484;
  assign n58447 = n39489 | ~n39490;
  assign n58448 = n39502 | ~n39503;
  assign n58449 = n39511 | n39512;
  assign n58450 = n39517 | n39518;
  assign n58451 = n39519 | n39520;
  assign n58452 = n39522 | ~n39523;
  assign n58453 = n39529 | n39530;
  assign n58454 = n39531 | n39532;
  assign n58455 = n39533 | ~n39534;
  assign n58456 = n39539 | ~n39540;
  assign n58457 = n39630 | ~n39631;
  assign n58458 = n39636 | ~n39637;
  assign n58459 = n39663 | n39664;
  assign n58460 = n39681 | n39682;
  assign n58461 = n39687 | n39688;
  assign n58462 = n39697 | n39698;
  assign n58463 = n39703 | n39704;
  assign n58464 = n39713 | n39714;
  assign n58465 = n39719 | n39720;
  assign n58466 = n39729 | n39730;
  assign n58467 = n39735 | n39736;
  assign n58468 = n39745 | n39746;
  assign n58469 = n39751 | n39752;
  assign n58470 = n39761 | n39762;
  assign n58471 = n39767 | n39768;
  assign n58472 = n39771 | n39772 | n39774 | n39775;
  assign n58473 = n39780 | n39781;
  assign n58474 = n39794 | ~n39795;
  assign n58475 = n39810 | n39811;
  assign n58476 = n39829 | n39821 | n39828;
  assign n58477 = n39839 | n39840;
  assign n58478 = n39847 | n39843 | n39846;
  assign n58479 = n39850 | n39851;
  assign n58480 = n39868 | n39869;
  assign n58481 = n39874 | n39875;
  assign n58482 = n39880 | ~n39881;
  assign n58483 = n39891 | n39892;
  assign n58484 = n39893 | n39894;
  assign n58485 = n39895 | ~n39896;
  assign n58486 = n39911 | n39912;
  assign n58487 = n39913 | n39914;
  assign n58488 = n39920 | ~n39921;
  assign n58489 = n39926 | ~n39927;
  assign n58490 = n39929 | ~n39930;
  assign n58491 = n39952 | n39953;
  assign n58492 = n39954 | n39955;
  assign n58493 = n39960 | ~n39961;
  assign n58494 = n39970 | n39971;
  assign n58495 = n39972 | n39973;
  assign n58496 = n39985 | n39986;
  assign n58497 = n39987 | n39988;
  assign n58498 = n40000 | ~n40001;
  assign n58499 = n40015 | n40016;
  assign n58500 = n40017 | n40018;
  assign n58501 = n40035 | n40036;
  assign n58502 = n40048 | ~n40049;
  assign n58503 = n40053 | n40054;
  assign n58504 = n40057 | n40058;
  assign n58505 = n40059 | n40060;
  assign n58506 = n40061 | ~n40062;
  assign n58507 = n40067 | ~n40068;
  assign n58508 = n40080 | n40081;
  assign n58509 = n40082 | n40083;
  assign n58510 = n40089 | n40090;
  assign n58511 = n40102 | ~n40103;
  assign n58512 = n40111 | n40112;
  assign n58513 = n40125 | n40126;
  assign n58514 = n40135 | ~n40136;
  assign n58515 = n40140 | n40141;
  assign n58516 = n40151 | n40152;
  assign n58517 = n40153 | n40154;
  assign n58518 = n40157 | n40158;
  assign n58519 = n40159 | n40160;
  assign n58520 = n40161 | ~n40162;
  assign n58521 = n40170 | n40171;
  assign n58522 = n40172 | n40173;
  assign n58523 = n40174 | ~n40175;
  assign n58524 = n40192 | n40193;
  assign n58525 = n40194 | n40195;
  assign n58526 = n40206 | ~n40207;
  assign n58527 = n40224 | n40225;
  assign n58528 = n40227 | n40228;
  assign n58529 = n40237 | n40238;
  assign n58530 = n40239 | n40240;
  assign n58531 = n40241 | ~n40242;
  assign n58532 = n40256 | ~n40257;
  assign n58533 = n40267 | ~n40268;
  assign n58534 = n40277 | ~n40278;
  assign n58535 = n40295 | ~n40296;
  assign n58536 = n40309 | n40310;
  assign n58537 = n40311 | n40312;
  assign n58538 = n40325 | ~n40326;
  assign n58539 = n40333 | ~n40334;
  assign n58540 = n40344 | n40345;
  assign n58541 = n40346 | n40347;
  assign n58542 = n40353 | n40354;
  assign n58543 = n40364 | ~n40365;
  assign n58544 = n40373 | n40374;
  assign n58545 = n40387 | n40388;
  assign n58546 = n40397 | ~n40398;
  assign n58547 = n40402 | n40403;
  assign n58548 = n40413 | n40414;
  assign n58549 = n40415 | n40416;
  assign n58550 = n40419 | n40420;
  assign n58551 = n40421 | n40422;
  assign n58552 = n40423 | ~n40424;
  assign n58553 = n40432 | n40433;
  assign n58554 = n40434 | n40435;
  assign n58555 = n40436 | ~n40437;
  assign n58556 = n40445 | n40446;
  assign n58557 = n40447 | n40448;
  assign n58558 = n40449 | ~n40450;
  assign n58559 = n40454 | n40455;
  assign n58560 = n40456 | n40457;
  assign n58561 = n40458 | ~n40459;
  assign n58562 = n40463 | n40464;
  assign n58563 = n40465 | n40466;
  assign n58564 = n40467 | ~n40468;
  assign n58565 = n40485 | n40486;
  assign n58566 = n40487 | n40488;
  assign n58567 = n40500 | n40501;
  assign n58568 = n40502 | n40503;
  assign n58569 = n40514 | ~n40515;
  assign n58570 = n40521 | n40522;
  assign n58571 = n40524 | n40525;
  assign n58572 = n40528 | n40529;
  assign n58573 = n40530 | n40531;
  assign n58574 = n40532 | ~n40533;
  assign n58575 = n40545 | ~n40546;
  assign n58576 = n40552 | n40553;
  assign n58577 = n40554 | n40555;
  assign n58578 = n40556 | ~n40557;
  assign n58579 = n40560 | n40561;
  assign n58580 = n40562 | n40563;
  assign n58581 = n40564 | ~n40565;
  assign n58582 = n40570 | ~n40571;
  assign n58583 = n40578 | ~n40579;
  assign n58584 = n40588 | ~n40589;
  assign n58585 = n40597 | ~n40598;
  assign n58586 = n40607 | n40608;
  assign n58587 = n40609 | n40610;
  assign n58588 = n40625 | n40626;
  assign n58589 = n40627 | n40628;
  assign n58590 = n40633 | ~n40634;
  assign n58591 = n40644 | n40645;
  assign n58592 = n40646 | n40647;
  assign n58593 = n40650 | n40651;
  assign n58594 = n40652 | n40653;
  assign n58595 = n40654 | ~n40655;
  assign n58596 = n40667 | ~n40668;
  assign n58597 = n40683 | ~n40684;
  assign n58598 = n40699 | ~n40700;
  assign n58599 = n40713 | n40714;
  assign n58600 = n40715 | n40716;
  assign n58601 = n40729 | ~n40730;
  assign n58602 = n40737 | ~n40738;
  assign n58603 = n40748 | n40749;
  assign n58604 = n40750 | n40751;
  assign n58605 = n40757 | n40758;
  assign n58606 = n40768 | ~n40769;
  assign n58607 = n40777 | n40778;
  assign n58608 = n40791 | n40792;
  assign n58609 = n40801 | ~n40802;
  assign n58610 = n40806 | n40807;
  assign n58611 = n40817 | n40818;
  assign n58612 = n40819 | n40820;
  assign n58613 = n40823 | n40824;
  assign n58614 = n40825 | n40826;
  assign n58615 = n40827 | ~n40828;
  assign n58616 = n40836 | n40837;
  assign n58617 = n40838 | n40839;
  assign n58618 = n40840 | ~n40841;
  assign n58619 = n40849 | n40850;
  assign n58620 = n40851 | n40852;
  assign n58621 = n40853 | ~n40854;
  assign n58622 = n40858 | n40859;
  assign n58623 = n40860 | n40861;
  assign n58624 = n40862 | ~n40863;
  assign n58625 = n40867 | n40868;
  assign n58626 = n40869 | n40870;
  assign n58627 = n40871 | ~n40872;
  assign n58628 = n40882 | ~n40883;
  assign n58629 = n40887 | n40888;
  assign n58630 = n40889 | n40890;
  assign n58631 = n40891 | ~n40892;
  assign n58632 = n40896 | n40897;
  assign n58633 = n40898 | n40899;
  assign n58634 = n40900 | ~n40901;
  assign n58635 = n40905 | n40906;
  assign n58636 = n40907 | n40908;
  assign n58637 = n40909 | ~n40910;
  assign n58638 = n40922 | n40923;
  assign n58639 = n40924 | n40925;
  assign n58640 = n40937 | n40938;
  assign n58641 = n40939 | n40940;
  assign n58642 = n40950 | n40951;
  assign n58643 = n40952 | n40953;
  assign n58644 = n40960 | ~n40961;
  assign n58645 = n40967 | n40968;
  assign n58646 = n40969 | n40970;
  assign n58647 = n40971 | ~n40972;
  assign n58648 = n40984 | ~n40985;
  assign n58649 = n40997 | n40998;
  assign n58650 = n40999 | n41000;
  assign n58651 = n41001 | ~n41002;
  assign n58652 = n41016 | ~n41017;
  assign n58653 = n41031 | ~n41032;
  assign n58654 = n41041 | n41042;
  assign n58655 = n41043 | n41044;
  assign n58656 = n41049 | ~n41050;
  assign n58657 = n41057 | ~n41058;
  assign n58658 = n41067 | ~n41068;
  assign n58659 = n41083 | ~n41084;
  assign n58660 = n41099 | ~n41100;
  assign n58661 = n41113 | n41114;
  assign n58662 = n41115 | n41116;
  assign n58663 = n41129 | n41130;
  assign n58664 = n41131 | n41132;
  assign n58665 = n41137 | ~n41138;
  assign n58666 = n41148 | n41149;
  assign n58667 = n41150 | n41151;
  assign n58668 = n41154 | n41155;
  assign n58669 = n41156 | n41157;
  assign n58670 = n41158 | ~n41159;
  assign n58671 = n41171 | ~n41172;
  assign n58672 = n41187 | ~n41188;
  assign n58673 = n41203 | ~n41204;
  assign n58674 = n41217 | n41218;
  assign n58675 = n41219 | n41220;
  assign n58676 = n41233 | ~n41234;
  assign n58677 = n41241 | ~n41242;
  assign n58678 = n41252 | n41253;
  assign n58679 = n41254 | n41255;
  assign n58680 = n41261 | n41262;
  assign n58681 = n41272 | ~n41273;
  assign n58682 = n41281 | n41282;
  assign n58683 = n41295 | n41296;
  assign n58684 = n41305 | ~n41306;
  assign n58685 = n41310 | n41311;
  assign n58686 = n41321 | n41322;
  assign n58687 = n41323 | n41324;
  assign n58688 = n41327 | n41328;
  assign n58689 = n41329 | n41330;
  assign n58690 = n41331 | ~n41332;
  assign n58691 = n41340 | n41341;
  assign n58692 = n41342 | n41343;
  assign n58693 = n41344 | ~n41345;
  assign n58694 = n41353 | n41354;
  assign n58695 = n41355 | n41356;
  assign n58696 = n41357 | ~n41358;
  assign n58697 = n41362 | n41363;
  assign n58698 = n41364 | n41365;
  assign n58699 = n41366 | ~n41367;
  assign n58700 = n41371 | n41372;
  assign n58701 = n41373 | n41374;
  assign n58702 = n41375 | ~n41376;
  assign n58703 = n41386 | ~n41387;
  assign n58704 = n41391 | n41392;
  assign n58705 = n41393 | n41394;
  assign n58706 = n41395 | ~n41396;
  assign n58707 = n41400 | n41401;
  assign n58708 = n41402 | n41403;
  assign n58709 = n41404 | ~n41405;
  assign n58710 = n41409 | n41410;
  assign n58711 = n41411 | n41412;
  assign n58712 = n41413 | ~n41414;
  assign n58713 = n41418 | n41419;
  assign n58714 = n41420 | n41421;
  assign n58715 = n41422 | ~n41423;
  assign n58716 = n41431 | n41432;
  assign n58717 = n41433 | n41434;
  assign n58718 = n41435 | ~n41436;
  assign n58719 = n41440 | n41441;
  assign n58720 = n41442 | n41443;
  assign n58721 = n41444 | ~n41445;
  assign n58722 = n41457 | n41458;
  assign n58723 = n41459 | n41460;
  assign n58724 = n41472 | n41473;
  assign n58725 = n41474 | n41475;
  assign n58726 = n41486 | ~n41487;
  assign n58727 = n41500 | n41501;
  assign n58728 = n41502 | n41503;
  assign n58729 = n41509 | n41510;
  assign n58730 = n41524 | n41532 | n41541 | n41542;
  assign n58731 = n41545 | n41546;
  assign n58732 = n41574 | n41561 | n41573;
  assign n58733 = n41580 | n41581;
  assign n58734 = n41597 | n41598;
  assign n58735 = n41599 | n41600;
  assign n58736 = n41615 | n41616;
  assign n58737 = n41634 | n41635;
  assign n58738 = n41641 | n41642;
  assign n58739 = n41645 | n41646;
  assign n58740 = n41647 | n41648;
  assign n58741 = n41649 | ~n41650;
  assign n58742 = n41655 | ~n41656;
  assign n58743 = n41661 | ~n41662;
  assign n58744 = n41665 | n41666;
  assign n58745 = n41667 | n41668;
  assign n58746 = n41669 | ~n41670;
  assign n58747 = n41675 | ~n41676;
  assign n58748 = n41679 | n41680;
  assign n58749 = n41681 | n41682;
  assign n58750 = n41683 | ~n41684;
  assign n58751 = n41696 | ~n41697;
  assign n58752 = n41703 | n41704;
  assign n58753 = n41705 | n41706;
  assign n58754 = n41707 | ~n41708;
  assign n58755 = n41711 | n41712;
  assign n58756 = n41713 | n41714;
  assign n58757 = n41715 | ~n41716;
  assign n58758 = n41721 | ~n41722;
  assign n58759 = n41729 | ~n41730;
  assign n58760 = n41739 | ~n41740;
  assign n58761 = n41746 | n41747;
  assign n58762 = n41748 | n41749;
  assign n58763 = n41750 | ~n41751;
  assign n58764 = n41756 | ~n41757;
  assign n58765 = n41771 | ~n41772;
  assign n58766 = n41782 | ~n41783;
  assign n58767 = n41792 | ~n41793;
  assign n58768 = n41806 | n41807;
  assign n58769 = n41808 | n41809;
  assign n58770 = n41822 | n41823;
  assign n58771 = n41824 | n41825;
  assign n58772 = n41828 | n41829;
  assign n58773 = n41830 | n41831;
  assign n58774 = n41832 | ~n41833;
  assign n58775 = n41843 | n41844;
  assign n58776 = n41845 | n41846;
  assign n58777 = n41851 | ~n41852;
  assign n58778 = n41864 | ~n41865;
  assign n58779 = n41880 | ~n41881;
  assign n58780 = n41896 | ~n41897;
  assign n58781 = n41910 | n41911;
  assign n58782 = n41912 | n41913;
  assign n58783 = n41926 | n41927;
  assign n58784 = n41928 | n41929;
  assign n58785 = n41934 | ~n41935;
  assign n58786 = n41945 | n41946;
  assign n58787 = n41947 | n41948;
  assign n58788 = n41951 | n41952;
  assign n58789 = n41953 | n41954;
  assign n58790 = n41955 | ~n41956;
  assign n58791 = n41968 | ~n41969;
  assign n58792 = n41984 | ~n41985;
  assign n58793 = n42000 | ~n42001;
  assign n58794 = n42014 | n42015;
  assign n58795 = n42016 | n42017;
  assign n58796 = n42030 | ~n42031;
  assign n58797 = n42038 | ~n42039;
  assign n58798 = n42049 | n42050;
  assign n58799 = n42051 | n42052;
  assign n58800 = n42058 | n42059;
  assign n58801 = n42069 | ~n42070;
  assign n58802 = n42078 | n42079;
  assign n58803 = n42092 | n42093;
  assign n58804 = n42102 | ~n42103;
  assign n58805 = n42107 | n42108;
  assign n58806 = n42118 | n42119;
  assign n58807 = n42120 | n42121;
  assign n58808 = n42124 | n42125;
  assign n58809 = n42126 | n42127;
  assign n58810 = n42128 | ~n42129;
  assign n58811 = n42137 | n42138;
  assign n58812 = n42139 | n42140;
  assign n58813 = n42141 | ~n42142;
  assign n58814 = n42150 | n42151;
  assign n58815 = n42152 | n42153;
  assign n58816 = n42154 | ~n42155;
  assign n58817 = n42159 | n42160;
  assign n58818 = n42161 | n42162;
  assign n58819 = n42163 | ~n42164;
  assign n58820 = n42168 | n42169;
  assign n58821 = n42170 | n42171;
  assign n58822 = n42172 | ~n42173;
  assign n58823 = n42183 | ~n42184;
  assign n58824 = n42188 | n42189;
  assign n58825 = n42190 | n42191;
  assign n58826 = n42192 | ~n42193;
  assign n58827 = n42197 | n42198;
  assign n58828 = n42199 | n42200;
  assign n58829 = n42201 | ~n42202;
  assign n58830 = n42206 | n42207;
  assign n58831 = n42208 | n42209;
  assign n58832 = n42210 | ~n42211;
  assign n58833 = n42215 | n42216;
  assign n58834 = n42217 | n42218;
  assign n58835 = n42219 | ~n42220;
  assign n58836 = n42228 | n42229;
  assign n58837 = n42230 | n42231;
  assign n58838 = n42232 | ~n42233;
  assign n58839 = n42239 | ~n42240;
  assign n58840 = n42244 | n42245;
  assign n58841 = n42246 | n42247;
  assign n58842 = n42248 | ~n42249;
  assign n58843 = n42253 | n42254;
  assign n58844 = n42255 | n42256;
  assign n58845 = n42257 | ~n42258;
  assign n58846 = n42266 | n42267;
  assign n58847 = n42268 | n42269;
  assign n58848 = n42270 | ~n42271;
  assign n58849 = n42277 | ~n42278;
  assign n58850 = n42287 | n42288;
  assign n58851 = n42289 | n42290;
  assign n58852 = n42302 | n42303;
  assign n58853 = n42304 | n42305;
  assign n58854 = n42317 | n42318;
  assign n58855 = n42319 | n42320;
  assign n58856 = n42332 | n42333;
  assign n58857 = n42334 | n42335;
  assign n58858 = n42339 | n42340;
  assign n58859 = n42353 | n42350 | n42352;
  assign n58860 = n42362 | n42363;
  assign n58861 = n42372 | n42373;
  assign n58862 = n42392 | n42393;
  assign n58863 = n42408 | ~n42409;
  assign n58864 = n42414 | ~n42415;
  assign n58865 = n42427 | ~n42428;
  assign n58866 = n42434 | n42435;
  assign n58867 = n42436 | n42437;
  assign n58868 = n42438 | ~n42439;
  assign n58869 = n42444 | ~n42445;
  assign n58870 = n42448 | n42449;
  assign n58871 = n42450 | n42451;
  assign n58872 = n42452 | ~n42453;
  assign n58873 = n42465 | ~n42466;
  assign n58874 = n42472 | n42473;
  assign n58875 = n42474 | n42475;
  assign n58876 = n42476 | ~n42477;
  assign n58877 = n42480 | n42481;
  assign n58878 = n42482 | n42483;
  assign n58879 = n42484 | ~n42485;
  assign n58880 = n42490 | ~n42491;
  assign n58881 = n42503 | ~n42504;
  assign n58882 = n42510 | n42511;
  assign n58883 = n42512 | n42513;
  assign n58884 = n42514 | ~n42515;
  assign n58885 = n42520 | ~n42521;
  assign n58886 = n42524 | n42525;
  assign n58887 = n42526 | n42527;
  assign n58888 = n42528 | ~n42529;
  assign n58889 = n42536 | ~n42537;
  assign n58890 = n42546 | ~n42547;
  assign n58891 = n42557 | ~n42558;
  assign n58892 = n42567 | ~n42568;
  assign n58893 = n42583 | n42584;
  assign n58894 = n42585 | n42586;
  assign n58895 = n42599 | n42600;
  assign n58896 = n42601 | n42602;
  assign n58897 = n42605 | n42606;
  assign n58898 = n42607 | n42608;
  assign n58899 = n42609 | ~n42610;
  assign n58900 = n42622 | ~n42623;
  assign n58901 = n42638 | ~n42639;
  assign n58902 = n42654 | ~n42655;
  assign n58903 = n42668 | n42669;
  assign n58904 = n42670 | n42671;
  assign n58905 = n42684 | n42685;
  assign n58906 = n42686 | n42687;
  assign n58907 = n42690 | n42691;
  assign n58908 = n42692 | n42693;
  assign n58909 = n42694 | ~n42695;
  assign n58910 = n42705 | n42706;
  assign n58911 = n42707 | n42708;
  assign n58912 = n42713 | ~n42714;
  assign n58913 = n42726 | ~n42727;
  assign n58914 = n42742 | ~n42743;
  assign n58915 = n42758 | ~n42759;
  assign n58916 = n42772 | n42773;
  assign n58917 = n42774 | n42775;
  assign n58918 = n42788 | n42789;
  assign n58919 = n42790 | n42791;
  assign n58920 = n42796 | ~n42797;
  assign n58921 = n42807 | n42808;
  assign n58922 = n42809 | n42810;
  assign n58923 = n42813 | n42814;
  assign n58924 = n42815 | n42816;
  assign n58925 = n42817 | ~n42818;
  assign n58926 = n42830 | ~n42831;
  assign n58927 = n42846 | ~n42847;
  assign n58928 = n42862 | ~n42863;
  assign n58929 = n42876 | n42877;
  assign n58930 = n42878 | n42879;
  assign n58931 = n42892 | ~n42893;
  assign n58932 = n42900 | ~n42901;
  assign n58933 = n42911 | n42912;
  assign n58934 = n42913 | n42914;
  assign n58935 = n42920 | n42921;
  assign n58936 = n42931 | ~n42932;
  assign n58937 = n42940 | n42941;
  assign n58938 = n42954 | n42955;
  assign n58939 = n42964 | ~n42965;
  assign n58940 = n42969 | n42970;
  assign n58941 = n42980 | n42981;
  assign n58942 = n42982 | n42983;
  assign n58943 = n42986 | n42987;
  assign n58944 = n42988 | n42989;
  assign n58945 = n42990 | ~n42991;
  assign n58946 = n42999 | n43000;
  assign n58947 = n43001 | n43002;
  assign n58948 = n43003 | ~n43004;
  assign n58949 = n43012 | n43013;
  assign n58950 = n43014 | n43015;
  assign n58951 = n43016 | ~n43017;
  assign n58952 = n43021 | n43022;
  assign n58953 = n43023 | n43024;
  assign n58954 = n43025 | ~n43026;
  assign n58955 = n43030 | n43031;
  assign n58956 = n43032 | n43033;
  assign n58957 = n43034 | ~n43035;
  assign n58958 = n43045 | ~n43046;
  assign n58959 = n43050 | n43051;
  assign n58960 = n43052 | n43053;
  assign n58961 = n43054 | ~n43055;
  assign n58962 = n43059 | n43060;
  assign n58963 = n43061 | n43062;
  assign n58964 = n43063 | ~n43064;
  assign n58965 = n43068 | n43069;
  assign n58966 = n43070 | n43071;
  assign n58967 = n43072 | ~n43073;
  assign n58968 = n43077 | n43078;
  assign n58969 = n43079 | n43080;
  assign n58970 = n43081 | ~n43082;
  assign n58971 = n43090 | n43091;
  assign n58972 = n43092 | n43093;
  assign n58973 = n43094 | ~n43095;
  assign n58974 = n43101 | ~n43102;
  assign n58975 = n43106 | n43107;
  assign n58976 = n43108 | n43109;
  assign n58977 = n43110 | ~n43111;
  assign n58978 = n43115 | n43116;
  assign n58979 = n43117 | n43118;
  assign n58980 = n43119 | ~n43120;
  assign n58981 = n43124 | n43125;
  assign n58982 = n43126 | n43127;
  assign n58983 = n43128 | ~n43129;
  assign n58984 = n43139 | ~n43140;
  assign n58985 = n43144 | n43145;
  assign n58986 = n43146 | n43147;
  assign n58987 = n43148 | ~n43149;
  assign n58988 = n43153 | n43154;
  assign n58989 = n43155 | n43156;
  assign n58990 = n43157 | ~n43158;
  assign n58991 = n43162 | n43163;
  assign n58992 = n43164 | n43165;
  assign n58993 = n43166 | ~n43167;
  assign n58994 = n43179 | n43180;
  assign n58995 = n43181 | n43182;
  assign n58996 = n43194 | n43195;
  assign n58997 = n43196 | n43197;
  assign n58998 = n43209 | n43210;
  assign n58999 = n43211 | n43212;
  assign n59000 = n43224 | n43225;
  assign n59001 = n43226 | n43227;
  assign n59002 = n43230 | n43231;
  assign n59003 = n43239 | n43240;
  assign n59004 = n43248 | n43249;
  assign n59005 = n43265 | n43257 | n43264;
  assign n59006 = n43284 | n43285;
  assign n59007 = n43294 | n43295;
  assign n59008 = n43298 | n43299;
  assign n59009 = n43300 | n43301;
  assign n59010 = n43302 | ~n43303;
  assign n59011 = n43308 | ~n43309;
  assign n59012 = n43312 | n43313;
  assign n59013 = n43314 | n43315;
  assign n59014 = n43316 | ~n43317;
  assign n59015 = n43329 | ~n43330;
  assign n59016 = n43336 | n43337;
  assign n59017 = n43338 | n43339;
  assign n59018 = n43340 | ~n43341;
  assign n59019 = n43344 | n43345;
  assign n59020 = n43346 | n43347;
  assign n59021 = n43348 | ~n43349;
  assign n59022 = n43354 | ~n43355;
  assign n59023 = n43367 | ~n43368;
  assign n59024 = n43374 | n43375;
  assign n59025 = n43376 | n43377;
  assign n59026 = n43378 | ~n43379;
  assign n59027 = n43384 | ~n43385;
  assign n59028 = n43388 | n43389;
  assign n59029 = n43390 | n43391;
  assign n59030 = n43392 | ~n43393;
  assign n59031 = n43405 | ~n43406;
  assign n59032 = n43412 | n43413;
  assign n59033 = n43414 | n43415;
  assign n59034 = n43416 | ~n43417;
  assign n59035 = n43420 | n43421;
  assign n59036 = n43422 | n43423;
  assign n59037 = n43424 | ~n43425;
  assign n59038 = n43430 | ~n43431;
  assign n59039 = n43445 | ~n43446;
  assign n59040 = n43452 | n43453;
  assign n59041 = n43454 | n43455;
  assign n59042 = n43456 | ~n43457;
  assign n59043 = n43462 | ~n43463;
  assign n59044 = n43468 | ~n43469;
  assign n59045 = n43478 | n43479;
  assign n59046 = n43480 | n43481;
  assign n59047 = n43484 | n43485;
  assign n59048 = n43486 | n43487;
  assign n59049 = n43488 | ~n43489;
  assign n59050 = n43494 | ~n43495;
  assign n59051 = n43504 | n43505;
  assign n59052 = n43506 | n43507;
  assign n59053 = n43510 | n43511;
  assign n59054 = n43512 | n43513;
  assign n59055 = n43514 | ~n43515;
  assign n59056 = n43527 | ~n43528;
  assign n59057 = n43543 | ~n43544;
  assign n59058 = n43557 | n43558;
  assign n59059 = n43559 | n43560;
  assign n59060 = n43573 | n43574;
  assign n59061 = n43575 | n43576;
  assign n59062 = n43581 | ~n43582;
  assign n59063 = n43592 | n43593;
  assign n59064 = n43594 | n43595;
  assign n59065 = n43598 | n43599;
  assign n59066 = n43600 | n43601;
  assign n59067 = n43602 | ~n43603;
  assign n59068 = n43615 | ~n43616;
  assign n59069 = n43631 | ~n43632;
  assign n59070 = n43647 | ~n43648;
  assign n59071 = n43661 | n43662;
  assign n59072 = n43663 | n43664;
  assign n59073 = n43677 | n43678;
  assign n59074 = n43679 | n43680;
  assign n59075 = n43683 | n43684;
  assign n59076 = n43685 | n43686;
  assign n59077 = n43687 | ~n43688;
  assign n59078 = n43698 | n43699;
  assign n59079 = n43700 | n43701;
  assign n59080 = n43706 | ~n43707;
  assign n59081 = n43719 | ~n43720;
  assign n59082 = n43735 | ~n43736;
  assign n59083 = n43751 | ~n43752;
  assign n59084 = n43765 | n43766;
  assign n59085 = n43767 | n43768;
  assign n59086 = n43781 | n43782;
  assign n59087 = n43783 | n43784;
  assign n59088 = n43789 | ~n43790;
  assign n59089 = n43800 | n43801;
  assign n59090 = n43802 | n43803;
  assign n59091 = n43806 | n43807;
  assign n59092 = n43808 | n43809;
  assign n59093 = n43810 | ~n43811;
  assign n59094 = n43823 | ~n43824;
  assign n59095 = n43839 | ~n43840;
  assign n59096 = n43855 | ~n43856;
  assign n59097 = n43869 | n43870;
  assign n59098 = n43871 | n43872;
  assign n59099 = n43885 | ~n43886;
  assign n59100 = n43893 | ~n43894;
  assign n59101 = n43904 | n43905;
  assign n59102 = n43906 | n43907;
  assign n59103 = n43913 | n43914;
  assign n59104 = n43924 | ~n43925;
  assign n59105 = n43933 | n43934;
  assign n59106 = n43947 | n43948;
  assign n59107 = n43957 | ~n43958;
  assign n59108 = n43962 | n43963;
  assign n59109 = n43973 | n43974;
  assign n59110 = n43975 | n43976;
  assign n59111 = n43979 | n43980;
  assign n59112 = n43981 | n43982;
  assign n59113 = n43983 | ~n43984;
  assign n59114 = n43992 | n43993;
  assign n59115 = n43994 | n43995;
  assign n59116 = n43996 | ~n43997;
  assign n59117 = n44005 | n44006;
  assign n59118 = n44007 | n44008;
  assign n59119 = n44009 | ~n44010;
  assign n59120 = n44014 | n44015;
  assign n59121 = n44016 | n44017;
  assign n59122 = n44018 | ~n44019;
  assign n59123 = n44023 | n44024;
  assign n59124 = n44025 | n44026;
  assign n59125 = n44027 | ~n44028;
  assign n59126 = n44038 | ~n44039;
  assign n59127 = n44043 | n44044;
  assign n59128 = n44045 | n44046;
  assign n59129 = n44047 | ~n44048;
  assign n59130 = n44052 | n44053;
  assign n59131 = n44054 | n44055;
  assign n59132 = n44056 | ~n44057;
  assign n59133 = n44061 | n44062;
  assign n59134 = n44063 | n44064;
  assign n59135 = n44065 | ~n44066;
  assign n59136 = n44070 | n44071;
  assign n59137 = n44072 | n44073;
  assign n59138 = n44074 | ~n44075;
  assign n59139 = n44083 | n44084;
  assign n59140 = n44085 | n44086;
  assign n59141 = n44087 | ~n44088;
  assign n59142 = n44094 | ~n44095;
  assign n59143 = n44099 | n44100;
  assign n59144 = n44101 | n44102;
  assign n59145 = n44103 | ~n44104;
  assign n59146 = n44108 | n44109;
  assign n59147 = n44110 | n44111;
  assign n59148 = n44112 | ~n44113;
  assign n59149 = n44117 | n44118;
  assign n59150 = n44119 | n44120;
  assign n59151 = n44121 | ~n44122;
  assign n59152 = n44132 | ~n44133;
  assign n59153 = n44137 | n44138;
  assign n59154 = n44139 | n44140;
  assign n59155 = n44141 | ~n44142;
  assign n59156 = n44146 | n44147;
  assign n59157 = n44148 | n44149;
  assign n59158 = n44150 | ~n44151;
  assign n59159 = n44155 | n44156;
  assign n59160 = n44157 | n44158;
  assign n59161 = n44159 | ~n44160;
  assign n59162 = n44170 | ~n44171;
  assign n59163 = n44177 | ~n44178;
  assign n59164 = n44182 | n44183;
  assign n59165 = n44184 | n44185;
  assign n59166 = n44186 | ~n44187;
  assign n59167 = n44197 | n44198;
  assign n59168 = n44201 | n44202;
  assign n59169 = n44203 | n44204;
  assign n59170 = n44207 | ~n44208;
  assign n59171 = n44211 | n44212;
  assign n59172 = n44213 | n44214;
  assign n59173 = n44215 | ~n44216;
  assign n59174 = n44231 | n44232;
  assign n59175 = n44248 | n44239 | n44247;
  assign n59176 = n44267 | n44268;
  assign n59177 = n44289 | ~n44290;
  assign n59178 = n44302 | n44303;
  assign n59179 = n44304 | n44305;
  assign n59180 = n44311 | ~n44312;
  assign n59181 = n44317 | ~n44318;
  assign n59182 = n44320 | ~n44321;
  assign n59183 = n44332 | n44333;
  assign n59184 = n44338 | ~n44339;
  assign n59185 = n44348 | n44349;
  assign n59186 = n44350 | n44351;
  assign n59187 = n44363 | n44364;
  assign n59188 = n44365 | n44366;
  assign n59189 = n44378 | n44379;
  assign n59190 = n44380 | n44381;
  assign n59191 = n44393 | n44394;
  assign n59192 = n44395 | n44396;
  assign n59193 = n44408 | n44409;
  assign n59194 = n44410 | n44411;
  assign n59195 = n44445 | n44433 | n44444;
  assign n59196 = n44461 | n44462;
  assign n59197 = n44471 | n44472;
  assign n59198 = n44475 | n44476;
  assign n59199 = n44477 | n44478;
  assign n59200 = n44479 | ~n44480;
  assign n59201 = n44485 | ~n44486;
  assign n59202 = n44489 | n44490;
  assign n59203 = n44491 | n44492;
  assign n59204 = n44493 | ~n44494;
  assign n59205 = n44506 | ~n44507;
  assign n59206 = n44513 | n44514;
  assign n59207 = n44515 | n44516;
  assign n59208 = n44517 | ~n44518;
  assign n59209 = n44521 | n44522;
  assign n59210 = n44523 | n44524;
  assign n59211 = n44525 | ~n44526;
  assign n59212 = n44531 | ~n44532;
  assign n59213 = n44544 | ~n44545;
  assign n59214 = n44551 | n44552;
  assign n59215 = n44553 | n44554;
  assign n59216 = n44555 | ~n44556;
  assign n59217 = n44561 | ~n44562;
  assign n59218 = n44565 | n44566;
  assign n59219 = n44567 | n44568;
  assign n59220 = n44569 | ~n44570;
  assign n59221 = n44582 | ~n44583;
  assign n59222 = n44589 | n44590;
  assign n59223 = n44591 | n44592;
  assign n59224 = n44593 | ~n44594;
  assign n59225 = n44597 | n44598;
  assign n59226 = n44599 | n44600;
  assign n59227 = n44601 | ~n44602;
  assign n59228 = n44607 | ~n44608;
  assign n59229 = n44620 | ~n44621;
  assign n59230 = n44627 | n44628;
  assign n59231 = n44629 | n44630;
  assign n59232 = n44631 | ~n44632;
  assign n59233 = n44637 | ~n44638;
  assign n59234 = n44641 | n44642;
  assign n59235 = n44643 | n44644;
  assign n59236 = n44645 | ~n44646;
  assign n59237 = n44657 | n44654 | n44656;
  assign n59238 = n44660 | n44661;
  assign n59239 = n44662 | n44663;
  assign n59240 = n44673 | n44669 | n44672;
  assign n59241 = n44687 | n44682 | n44686;
  assign n59242 = n44693 | n44694;
  assign n59243 = n44698 | n44699;
  assign n59244 = n44713 | n44714;
  assign n59245 = n44726 | n44727;
  assign n59246 = n44732 | ~n44733;
  assign n59247 = n44745 | ~n44746;
  assign n59248 = n44754 | ~n44755;
  assign n59249 = n44761 | n44762;
  assign n59250 = n44763 | n44764;
  assign n59251 = n44765 | ~n44766;
  assign n59252 = n44771 | ~n44772;
  assign n59253 = n44787 | n44783 | n44786;
  assign n59254 = n44807 | n44804 | n44806;
  assign n59255 = n44819 | n44820;
  assign n59256 = n44825 | ~n44826;
  assign n59257 = n44834 | n44835;
  assign n59258 = n44845 | n44846;
  assign n59259 = n44847 | n44848;
  assign n59260 = n44852 | n44853;
  assign n59261 = n44854 | n44855;
  assign n59262 = n44856 | ~n44857;
  assign n59263 = ~n44865 | n44863 | n44864;
  assign n59264 = n44877 | n44878;
  assign n59265 = n44883 | n44884;
  assign n59266 = n44892 | n44893;
  assign n59267 = n44896 | n44897;
  assign n59268 = n44898 | n44899;
  assign n59269 = n44902 | n44903;
  assign n59270 = n44912 | n44913;
  assign n59271 = n44925 | n44926;
  assign n59272 = n44935 | ~n44936;
  assign n59273 = n44941 | ~n44942;
  assign n59274 = n44957 | n44958;
  assign n59275 = n44963 | ~n44964;
  assign n59276 = n44973 | ~n44974;
  assign n59277 = n44980 | n44981;
  assign n59278 = n44982 | n44983;
  assign n59279 = n44984 | ~n44985;
  assign n59280 = n44989 | ~n44990;
  assign n59281 = n44999 | ~n45000;
  assign n59282 = n45007 | ~n45008;
  assign n59283 = n45017 | ~n45018;
  assign n59284 = n45030 | ~n45031;
  assign n59285 = n45038 | n45039;
  assign n59286 = n45049 | ~n45050;
  assign n59287 = n45062 | ~n45063;
  assign n59288 = n45075 | ~n45076;
  assign n59289 = n45083 | n45084;
  assign n59290 = n45087 | n45088;
  assign n59291 = n45098 | ~n45099;
  assign n59292 = n45111 | ~n45112;
  assign n59293 = n45124 | ~n45125;
  assign n59294 = n45132 | n45133;
  assign n59295 = n45136 | n45137;
  assign n59296 = n45147 | ~n45148;
  assign n59297 = n45160 | ~n45161;
  assign n59298 = n45173 | ~n45174;
  assign n59299 = n45184 | n45181 | n45183;
  assign n59300 = n45187 | n45188;
  assign n59301 = n45198 | ~n45199;
  assign n59302 = n45211 | ~n45212;
  assign n59303 = n45224 | ~n45225;
  assign n59304 = n45239 | ~n45240;
  assign n59305 = n45248 | n45249;
  assign n59306 = n45258 | ~n45259;
  assign n59307 = n45285 | n45293 | n45295 | n45296;
  assign n59308 = n45288 | n45289;
  assign n59309 = n45309 | ~n45310;
  assign n59310 = n45318 | n45319;
  assign n59311 = n45335 | ~n45336;
  assign n59312 = n45358 | ~n45359;
  assign n59313 = n45393 | ~n45394;
  assign n59314 = n45410 | ~n45411;
  assign n59315 = n45427 | ~n45428;
  assign n59316 = n45462 | ~n45463;
  assign n59317 = n45479 | ~n45480;
  assign n59318 = n45496 | ~n45497;
  assign n59319 = n45531 | ~n45532;
  assign n59320 = n45548 | ~n45549;
  assign n59321 = n45565 | ~n45566;
  assign n59322 = n45600 | ~n45601;
  assign n59323 = n45617 | ~n45618;
  assign n59324 = n45650 | n45651;
  assign n59325 = n45652 | n45653;
  assign n59326 = n45665 | n45666;
  assign n59327 = n45667 | n45668;
  assign n59328 = n45680 | n45681;
  assign n59329 = n45682 | n45683;
  assign n59330 = n45695 | n45696;
  assign n59331 = n45697 | n45698;
  assign n59332 = n45710 | n45711;
  assign n59333 = n45712 | n45713;
  assign n59334 = n45733 | n45734;
  assign n59335 = n45749 | n45739 | n45748;
  assign n59336 = n45765 | n45766;
  assign n59337 = n45775 | n45776;
  assign n59338 = n45779 | n45780;
  assign n59339 = n45781 | n45782;
  assign n59340 = n45783 | ~n45784;
  assign n59341 = n45789 | ~n45790;
  assign n59342 = n45793 | n45794;
  assign n59343 = n45795 | n45796;
  assign n59344 = n45797 | ~n45798;
  assign n59345 = n45810 | ~n45811;
  assign n59346 = n45817 | n45818;
  assign n59347 = n45819 | n45820;
  assign n59348 = n45821 | ~n45822;
  assign n59349 = n45825 | n45826;
  assign n59350 = n45827 | n45828;
  assign n59351 = n45829 | ~n45830;
  assign n59352 = n45835 | ~n45836;
  assign n59353 = n45848 | ~n45849;
  assign n59354 = n45855 | n45856;
  assign n59355 = n45857 | n45858;
  assign n59356 = n45859 | ~n45860;
  assign n59357 = n45865 | ~n45866;
  assign n59358 = n45869 | n45870;
  assign n59359 = n45871 | n45872;
  assign n59360 = n45873 | ~n45874;
  assign n59361 = n45886 | ~n45887;
  assign n59362 = n45893 | n45894;
  assign n59363 = n45895 | n45896;
  assign n59364 = n45897 | ~n45898;
  assign n59365 = n45901 | n45902;
  assign n59366 = n45903 | n45904;
  assign n59367 = n45905 | ~n45906;
  assign n59368 = n45911 | ~n45912;
  assign n59369 = n45924 | ~n45925;
  assign n59370 = n45931 | n45932;
  assign n59371 = n45933 | n45934;
  assign n59372 = n45935 | ~n45936;
  assign n59373 = n45941 | ~n45942;
  assign n59374 = n45945 | n45946;
  assign n59375 = n45947 | n45948;
  assign n59376 = n45949 | ~n45950;
  assign n59377 = n45961 | n45962;
  assign n59378 = n45976 | ~n45977;
  assign n59379 = n45979 | ~n45980;
  assign n59380 = n45984 | ~n45985;
  assign n59381 = n45990 | n45987 | n45989;
  assign n59382 = n45991 | n45992 | n45993 | n45994;
  assign n59383 = n45996 | n45997;
  assign n59384 = n45998 | n45999;
  assign n59385 = n46014 | n46015;
  assign n59386 = n46020 | ~n46021;
  assign n59387 = n46030 | ~n46031;
  assign n59388 = n46042 | n46043;
  assign n59389 = n46044 | n46045;
  assign n59390 = n46046 | ~n46047;
  assign n59391 = n46052 | ~n46053;
  assign n59392 = n46064 | n46065;
  assign n59393 = n46066 | n46067;
  assign n59394 = n46079 | n46080;
  assign n59395 = n46081 | n46082;
  assign n59396 = n46094 | n46095;
  assign n59397 = n46096 | n46097;
  assign n59398 = n46109 | n46110;
  assign n59399 = n46111 | n46112;
  assign n59400 = n46124 | ~n46125;
  assign n59401 = n46136 | n46137;
  assign n59402 = n46173 | n46159 | n46172;
  assign n59403 = n46193 | n46194;
  assign n59404 = n46203 | n46204;
  assign n59405 = n46207 | n46208;
  assign n59406 = n46209 | n46210;
  assign n59407 = n46211 | ~n46212;
  assign n59408 = n46217 | ~n46218;
  assign n59409 = n46233 | ~n46234;
  assign n59410 = n46240 | n46241;
  assign n59411 = n46242 | n46243;
  assign n59412 = n46244 | ~n46245;
  assign n59413 = n46250 | ~n46251;
  assign n59414 = n46254 | n46255;
  assign n59415 = n46256 | n46257;
  assign n59416 = n46258 | ~n46259;
  assign n59417 = n46271 | ~n46272;
  assign n59418 = n46278 | n46279;
  assign n59419 = n46280 | n46281;
  assign n59420 = n46282 | ~n46283;
  assign n59421 = n46286 | n46287;
  assign n59422 = n46288 | n46289;
  assign n59423 = n46290 | ~n46291;
  assign n59424 = n46296 | ~n46297;
  assign n59425 = n46309 | ~n46310;
  assign n59426 = n46316 | n46317;
  assign n59427 = n46318 | n46319;
  assign n59428 = n46320 | ~n46321;
  assign n59429 = n46326 | ~n46327;
  assign n59430 = n46330 | n46331;
  assign n59431 = n46332 | n46333;
  assign n59432 = n46334 | ~n46335;
  assign n59433 = n46347 | ~n46348;
  assign n59434 = n46354 | n46355;
  assign n59435 = n46356 | n46357;
  assign n59436 = n46358 | ~n46359;
  assign n59437 = n46362 | n46363;
  assign n59438 = n46364 | n46365;
  assign n59439 = n46366 | ~n46367;
  assign n59440 = n46372 | ~n46373;
  assign n59441 = n46384 | ~n46385;
  assign n59442 = n46387 | n46388;
  assign n59443 = n46393 | ~n46394;
  assign n59444 = n46403 | n46404;
  assign n59445 = n46405 | n46406;
  assign n59446 = n46407 | ~n46408;
  assign n59447 = n46413 | ~n46414;
  assign n59448 = n46435 | ~n46436;
  assign n59449 = n46459 | n46460;
  assign n59450 = n46461 | n46462;
  assign n59451 = n46474 | n46475;
  assign n59452 = n46476 | n46477;
  assign n59453 = n46489 | n46490;
  assign n59454 = n46491 | n46492;
  assign n59455 = n46504 | n46505;
  assign n59456 = n46506 | n46507;
  assign n59457 = n46519 | ~n46520;
  assign n59458 = n46541 | n46535 | n46540;
  assign n59459 = n46548 | n46549;
  assign n59460 = n46573 | n46574;
  assign n59461 = n46583 | n46584;
  assign n59462 = n46587 | n46588;
  assign n59463 = n46589 | n46590;
  assign n59464 = n46591 | ~n46592;
  assign n59465 = n46597 | ~n46598;
  assign n59466 = n46613 | ~n46614;
  assign n59467 = n46620 | n46621;
  assign n59468 = n46622 | n46623;
  assign n59469 = n46624 | ~n46625;
  assign n59470 = n46630 | ~n46631;
  assign n59471 = n46634 | n46635;
  assign n59472 = n46636 | n46637;
  assign n59473 = n46638 | ~n46639;
  assign n59474 = n46651 | ~n46652;
  assign n59475 = n46658 | n46659;
  assign n59476 = n46660 | n46661;
  assign n59477 = n46662 | ~n46663;
  assign n59478 = n46666 | n46667;
  assign n59479 = n46668 | n46669;
  assign n59480 = n46670 | ~n46671;
  assign n59481 = n46676 | ~n46677;
  assign n59482 = n46689 | ~n46690;
  assign n59483 = n46696 | n46697;
  assign n59484 = n46698 | n46699;
  assign n59485 = n46700 | ~n46701;
  assign n59486 = n46706 | ~n46707;
  assign n59487 = n46710 | n46711;
  assign n59488 = n46712 | n46713;
  assign n59489 = n46714 | ~n46715;
  assign n59490 = n46727 | ~n46728;
  assign n59491 = n46734 | n46735;
  assign n59492 = n46736 | n46737;
  assign n59493 = n46738 | ~n46739;
  assign n59494 = n46742 | n46743;
  assign n59495 = n46744 | n46745;
  assign n59496 = n46746 | ~n46747;
  assign n59497 = n46752 | ~n46753;
  assign n59498 = n46769 | n46766 | n46768;
  assign n59499 = n46770 | n46771;
  assign n59500 = n46774 | n46775;
  assign n59501 = n46776 | n46777;
  assign n59502 = n46778 | ~n46779;
  assign n59503 = n46799 | n46800;
  assign n59504 = n46814 | ~n46815;
  assign n59505 = n46838 | n46839;
  assign n59506 = n46840 | n46841;
  assign n59507 = n46853 | n46854;
  assign n59508 = n46855 | n46856;
  assign n59509 = n46868 | n46869;
  assign n59510 = n46870 | n46871;
  assign n59511 = n46883 | n46884;
  assign n59512 = n46885 | n46886;
  assign n59513 = n46898 | ~n46899;
  assign n59514 = n46911 | n46912;
  assign n59515 = n46931 | n46922 | n46930;
  assign n59516 = n46947 | n46948;
  assign n59517 = n46957 | n46958;
  assign n59518 = n46961 | n46962;
  assign n59519 = n46963 | n46964;
  assign n59520 = n46965 | ~n46966;
  assign n59521 = n46971 | ~n46972;
  assign n59522 = n46987 | ~n46988;
  assign n59523 = n46994 | n46995;
  assign n59524 = n46996 | n46997;
  assign n59525 = n46998 | ~n46999;
  assign n59526 = n47004 | ~n47005;
  assign n59527 = n47008 | n47009;
  assign n59528 = n47010 | n47011;
  assign n59529 = n47012 | ~n47013;
  assign n59530 = n47025 | ~n47026;
  assign n59531 = n47032 | n47033;
  assign n59532 = n47034 | n47035;
  assign n59533 = n47036 | ~n47037;
  assign n59534 = n47040 | n47041;
  assign n59535 = n47042 | n47043;
  assign n59536 = n47044 | ~n47045;
  assign n59537 = n47050 | ~n47051;
  assign n59538 = n47063 | ~n47064;
  assign n59539 = n47070 | n47071;
  assign n59540 = n47072 | n47073;
  assign n59541 = n47074 | ~n47075;
  assign n59542 = n47080 | ~n47081;
  assign n59543 = n47084 | n47085;
  assign n59544 = n47086 | n47087;
  assign n59545 = n47088 | ~n47089;
  assign n59546 = n47101 | ~n47102;
  assign n59547 = n47108 | n47109;
  assign n59548 = n47110 | n47111;
  assign n59549 = n47112 | ~n47113;
  assign n59550 = n47116 | n47117;
  assign n59551 = n47118 | n47119;
  assign n59552 = n47120 | ~n47121;
  assign n59553 = n47126 | ~n47127;
  assign n59554 = n47137 | ~n47138;
  assign n59555 = n47147 | ~n47148;
  assign n59556 = n47171 | n47172;
  assign n59557 = n47173 | n47174;
  assign n59558 = n47186 | n47187;
  assign n59559 = n47188 | n47189;
  assign n59560 = n47201 | n47202;
  assign n59561 = n47203 | n47204;
  assign n59562 = n47216 | n47217;
  assign n59563 = n47218 | n47219;
  assign n59564 = n47231 | ~n47232;
  assign n59565 = n47280 | n47258 | n47272 | n47285 | n47286;
  assign n59566 = n47263 | n47264;
  assign n59567 = n47289 | n47290;
  assign n59568 = n47323 | n47306 | n47322;
  assign n59569 = n47342 | n47343;
  assign n59570 = n47352 | n47353;
  assign n59571 = n47356 | n47357;
  assign n59572 = n47358 | n47359;
  assign n59573 = n47360 | ~n47361;
  assign n59574 = n47366 | ~n47367;
  assign n59575 = n47382 | ~n47383;
  assign n59576 = n47389 | n47390;
  assign n59577 = n47391 | n47392;
  assign n59578 = n47393 | ~n47394;
  assign n59579 = n47399 | ~n47400;
  assign n59580 = n47403 | n47404;
  assign n59581 = n47405 | n47406;
  assign n59582 = n47407 | ~n47408;
  assign n59583 = n47420 | ~n47421;
  assign n59584 = n47427 | n47428;
  assign n59585 = n47429 | n47430;
  assign n59586 = n47431 | ~n47432;
  assign n59587 = n47435 | n47436;
  assign n59588 = n47437 | n47438;
  assign n59589 = n47439 | ~n47440;
  assign n59590 = n47445 | ~n47446;
  assign n59591 = n47458 | ~n47459;
  assign n59592 = n47465 | n47466;
  assign n59593 = n47467 | n47468;
  assign n59594 = n47469 | ~n47470;
  assign n59595 = n47475 | ~n47476;
  assign n59596 = n47479 | n47480;
  assign n59597 = n47481 | n47482;
  assign n59598 = n47483 | ~n47484;
  assign n59599 = n47496 | ~n47497;
  assign n59600 = n47503 | n47504;
  assign n59601 = n47505 | n47506;
  assign n59602 = n47507 | ~n47508;
  assign n59603 = n47511 | n47512;
  assign n59604 = n47513 | n47514;
  assign n59605 = n47515 | ~n47516;
  assign n59606 = n47521 | ~n47522;
  assign n59607 = n47533 | ~n47534;
  assign n59608 = n47557 | n47558;
  assign n59609 = n47559 | n47560;
  assign n59610 = n47572 | n47573;
  assign n59611 = n47574 | n47575;
  assign n59612 = n47587 | n47588;
  assign n59613 = n47589 | n47590;
  assign n59614 = n47602 | n47603;
  assign n59615 = n47604 | n47605;
  assign n59616 = n47617 | ~n47618;
  assign n59617 = n47644 | n47657 | n47671 | n47672;
  assign n59618 = n47691 | n47692;
  assign n59619 = n47701 | n47702;
  assign n59620 = n47705 | n47706;
  assign n59621 = n47707 | n47708;
  assign n59622 = n47709 | ~n47710;
  assign n59623 = n47715 | ~n47716;
  assign n59624 = n47731 | ~n47732;
  assign n59625 = n47738 | n47739;
  assign n59626 = n47740 | n47741;
  assign n59627 = n47742 | ~n47743;
  assign n59628 = n47748 | ~n47749;
  assign n59629 = n47752 | n47753;
  assign n59630 = n47754 | n47755;
  assign n59631 = n47756 | ~n47757;
  assign n59632 = n47769 | ~n47770;
  assign n59633 = n47776 | n47777;
  assign n59634 = n47778 | n47779;
  assign n59635 = n47780 | ~n47781;
  assign n59636 = n47784 | n47785;
  assign n59637 = n47786 | n47787;
  assign n59638 = n47788 | ~n47789;
  assign n59639 = n47794 | ~n47795;
  assign n59640 = n47807 | ~n47808;
  assign n59641 = n47814 | n47815;
  assign n59642 = n47816 | n47817;
  assign n59643 = n47818 | ~n47819;
  assign n59644 = n47824 | ~n47825;
  assign n59645 = n47828 | n47829;
  assign n59646 = n47830 | n47831;
  assign n59647 = n47832 | ~n47833;
  assign n59648 = n47845 | ~n47846;
  assign n59649 = n47852 | n47853;
  assign n59650 = n47854 | n47855;
  assign n59651 = n47856 | ~n47857;
  assign n59652 = n47860 | n47861;
  assign n59653 = n47862 | n47863;
  assign n59654 = n47864 | ~n47865;
  assign n59655 = n47870 | ~n47871;
  assign n59656 = n47895 | n47896;
  assign n59657 = n47897 | n47898;
  assign n59658 = n47910 | n47911;
  assign n59659 = n47912 | n47913;
  assign n59660 = n47925 | n47926;
  assign n59661 = n47927 | n47928;
  assign n59662 = n47940 | n47941;
  assign n59663 = n47942 | n47943;
  assign n59664 = n47955 | ~n47956;
  assign n59665 = n47972 | n47973;
  assign n59666 = n47977 | n47981 | n47984 | n47985;
  assign n59667 = n48001 | n48002;
  assign n59668 = n48033 | n48018 | n48032;
  assign n59669 = n48055 | n48056;
  assign n59670 = n48065 | n48066;
  assign n59671 = n48069 | n48070;
  assign n59672 = n48071 | n48072;
  assign n59673 = n48073 | ~n48074;
  assign n59674 = n48079 | ~n48080;
  assign n59675 = n48095 | ~n48096;
  assign n59676 = n48108 | n48109;
  assign n59677 = n48110 | n48111;
  assign n59678 = n48112 | ~n48113;
  assign n59679 = n48125 | ~n48126;
  assign n59680 = n48138 | n48139;
  assign n59681 = n48140 | n48141;
  assign n59682 = n48142 | ~n48143;
  assign n59683 = n48155 | ~n48156;
  assign n59684 = n48168 | n48169;
  assign n59685 = n48170 | n48171;
  assign n59686 = n48172 | ~n48173;
  assign n59687 = n48185 | ~n48186;
  assign n59688 = n48198 | n48199;
  assign n59689 = n48200 | n48201;
  assign n59690 = n48202 | ~n48203;
  assign n59691 = n48208 | ~n48209;
  assign n59692 = n48257 | n48245 | n48256;
  assign n59693 = n48260 | n48261;
  assign n59694 = n48281 | n48282;
  assign n59695 = n48298 | n48295 | n48297;
  assign n59696 = n48300 | n48301;
  assign n59697 = n48303 | ~n48304;
  assign n59698 = n48316 | ~n48317;
  assign n59699 = n48335 | n48336;
  assign n59700 = n48337 | n48338;
  assign n59701 = n48344 | ~n48345;
  assign n59702 = n48357 | n48358;
  assign n59703 = n48359 | n48360;
  assign n59704 = n48366 | ~n48367;
  assign n59705 = n48379 | n48380;
  assign n59706 = n48381 | n48382;
  assign n59707 = n48388 | ~n48389;
  assign n59708 = n48401 | n48402;
  assign n59709 = n48403 | n48404;
  assign n59710 = n48410 | ~n48411;
  assign n59711 = n48423 | n48424;
  assign n59712 = n48425 | n48426;
  assign n59713 = n48432 | ~n48433;
  assign n59714 = n48445 | n48446;
  assign n59715 = n48447 | n48448;
  assign n59716 = n48454 | ~n48455;
  assign n59717 = n48467 | n48468;
  assign n59718 = n48469 | n48470;
  assign n59719 = n48476 | ~n48477;
  assign n59720 = n48487 | n48488;
  assign n59721 = n48489 | n48490;
  assign n59722 = n48496 | ~n48497;
  assign n59723 = n48516 | n48517;
  assign n59724 = n48518 | n48519;
  assign n59725 = n48537 | n48538;
  assign n59726 = n48555 | n48544 | n48554;
  assign n59727 = n48558 | n48559;
  assign n59728 = n48564 | n48565;
  assign n59729 = n48586 | n48587;
  assign n59730 = n48592 | n48593;
  assign n59731 = n48598 | ~n48599;
  assign n59732 = n48609 | n48610;
  assign n59733 = n48611 | n48612;
  assign n59734 = n48613 | ~n48614;
  assign n59735 = n48626 | n48627;
  assign n59736 = n48628 | n48629;
  assign n59737 = n48633 | n48634;
  assign n59738 = n48635 | n48636;
  assign n59739 = n48637 | ~n48638;
  assign n59740 = n48641 | n48642;
  assign n59741 = n48643 | n48644;
  assign n59742 = n48645 | ~n48646;
  assign n59743 = n48648 | ~n48649;
  assign n59744 = n48661 | n48662;
  assign n59745 = n48663 | n48664;
  assign n59746 = n48670 | ~n48671;
  assign n59747 = n48673 | ~n48674;
  assign n59748 = n48686 | n48687;
  assign n59749 = n48688 | n48689;
  assign n59750 = n48695 | ~n48696;
  assign n59751 = n48698 | ~n48699;
  assign n59752 = n48711 | n48712;
  assign n59753 = n48713 | n48714;
  assign n59754 = n48720 | ~n48721;
  assign n59755 = n48723 | ~n48724;
  assign n59756 = n48736 | n48737;
  assign n59757 = n48738 | n48739;
  assign n59758 = n48745 | ~n48746;
  assign n59759 = n48748 | ~n48749;
  assign n59760 = n48761 | n48762;
  assign n59761 = n48763 | n48764;
  assign n59762 = n48770 | ~n48771;
  assign n59763 = n48773 | ~n48774;
  assign n59764 = n48786 | n48787;
  assign n59765 = n48788 | n48789;
  assign n59766 = n48795 | ~n48796;
  assign n59767 = n48798 | ~n48799;
  assign n59768 = n48805 | n48806;
  assign n59769 = n48807 | n48808;
  assign n59770 = n48814 | ~n48815;
  assign n59771 = n48817 | ~n48818;
  assign n59772 = n48830 | ~n48831;
  assign n59773 = n48844 | n48845;
  assign n59774 = n48846 | n48847;
  assign n59775 = n48857 | n48858;
  assign n59776 = n48869 | n48864 | n48868;
  assign n59777 = n48873 | n48874;
  assign n59778 = n48892 | n48893;
  assign n59779 = n48898 | n48899;
  assign n59780 = n48904 | ~n48905;
  assign n59781 = n48915 | n48916;
  assign n59782 = n48917 | n48918;
  assign n59783 = n48919 | ~n48920;
  assign n59784 = n48932 | n48933;
  assign n59785 = n48934 | n48935;
  assign n59786 = n48939 | n48940;
  assign n59787 = n48941 | n48942;
  assign n59788 = n48943 | ~n48944;
  assign n59789 = n48947 | n48948;
  assign n59790 = n48949 | n48950;
  assign n59791 = n48951 | ~n48952;
  assign n59792 = n48964 | n48965;
  assign n59793 = n48966 | n48967;
  assign n59794 = n48973 | ~n48974;
  assign n59795 = n48976 | ~n48977;
  assign n59796 = n48989 | n48990;
  assign n59797 = n48991 | n48992;
  assign n59798 = n48998 | ~n48999;
  assign n59799 = n49001 | ~n49002;
  assign n59800 = n49014 | n49015;
  assign n59801 = n49016 | n49017;
  assign n59802 = n49023 | ~n49024;
  assign n59803 = n49026 | ~n49027;
  assign n59804 = n49039 | n49040;
  assign n59805 = n49041 | n49042;
  assign n59806 = n49048 | ~n49049;
  assign n59807 = n49051 | ~n49052;
  assign n59808 = n49064 | n49065;
  assign n59809 = n49066 | n49067;
  assign n59810 = n49073 | ~n49074;
  assign n59811 = n49076 | ~n49077;
  assign n59812 = n49089 | n49090;
  assign n59813 = n49091 | n49092;
  assign n59814 = n49098 | ~n49099;
  assign n59815 = n49104 | ~n49105;
  assign n59816 = n49107 | ~n49108;
  assign n59817 = n49129 | n49130;
  assign n59818 = n49131 | n49132;
  assign n59819 = n49153 | n49154;
  assign n59820 = n49171 | n49172;
  assign n59821 = n49177 | ~n49178;
  assign n59822 = n49183 | ~n49184;
  assign n59823 = n49189 | ~n49190;
  assign n59824 = n49212 | n49213;
  assign n59825 = n49214 | n49215;
  assign n59826 = n49221 | ~n49222;
  assign n59827 = n49227 | ~n49228;
  assign n59828 = n49240 | n49241;
  assign n59829 = n49242 | n49243;
  assign n59830 = n49247 | n49248;
  assign n59831 = n49249 | n49250;
  assign n59832 = n49251 | ~n49252;
  assign n59833 = n49254 | ~n49255;
  assign n59834 = n49267 | n49268;
  assign n59835 = n49269 | n49270;
  assign n59836 = n49274 | n49275;
  assign n59837 = n49276 | n49277;
  assign n59838 = n49278 | ~n49279;
  assign n59839 = n49281 | ~n49282;
  assign n59840 = n49294 | n49295;
  assign n59841 = n49296 | n49297;
  assign n59842 = n49301 | n49302;
  assign n59843 = n49303 | n49304;
  assign n59844 = n49305 | ~n49306;
  assign n59845 = n49308 | ~n49309;
  assign n59846 = n49321 | n49322;
  assign n59847 = n49323 | n49324;
  assign n59848 = n49327 | ~n49328;
  assign n59849 = n49331 | n49332;
  assign n59850 = n49333 | n49334;
  assign n59851 = n49335 | ~n49336;
  assign n59852 = n49348 | n49349;
  assign n59853 = n49350 | n49351;
  assign n59854 = n49355 | n49356;
  assign n59855 = n49357 | n49358;
  assign n59856 = n49359 | ~n49360;
  assign n59857 = n49362 | ~n49363;
  assign n59858 = n49373 | n49374;
  assign n59859 = n49375 | n49376;
  assign n59860 = n49379 | ~n49380;
  assign n59861 = n49383 | n49384;
  assign n59862 = n49385 | n49386;
  assign n59863 = n49387 | ~n49388;
  assign n59864 = n49393 | ~n49394;
  assign n59865 = n49415 | n49416;
  assign n59866 = n49417 | n49418;
  assign n59867 = n49461 | n49448 | n49460;
  assign n59868 = n49480 | n49481;
  assign n59869 = n49510 | n49495 | n49509;
  assign n59870 = n49528 | n49529;
  assign n59871 = n49544 | ~n49545;
  assign n59872 = n49557 | ~n49558;
  assign n59873 = n49566 | ~n49567;
  assign n59874 = n49579 | n49580;
  assign n59875 = n49581 | n49582;
  assign n59876 = n49588 | ~n49589;
  assign n59877 = n49601 | n49602;
  assign n59878 = n49603 | n49604;
  assign n59879 = n49610 | ~n49611;
  assign n59880 = n49623 | n49624;
  assign n59881 = n49625 | n49626;
  assign n59882 = n49632 | ~n49633;
  assign n59883 = n49645 | n49646;
  assign n59884 = n49647 | n49648;
  assign n59885 = n49654 | ~n49655;
  assign n59886 = n49667 | n49668;
  assign n59887 = n49669 | n49670;
  assign n59888 = n49676 | ~n49677;
  assign n59889 = n49680 | n49681;
  assign n59890 = n49682 | n49683;
  assign n59891 = n49684 | ~n49685;
  assign n59892 = n49690 | ~n49691;
  assign n59893 = n49697 | n49698;
  assign n59894 = n49699 | n49700;
  assign n59895 = n49706 | ~n49707;
  assign n59896 = n49712 | ~n49713;
  assign n59897 = n49732 | n49733;
  assign n59898 = n49734 | n49735;
  assign n59899 = n49745 | n49746;
  assign n59900 = n49751 | n49752;
  assign n59901 = n49762 | n49763;
  assign n59902 = n49767 | n49768;
  assign n59903 = n49780 | n49781;
  assign n59904 = n49790 | n49791;
  assign n59905 = n49799 | n49806 | n49812 | n49813;
  assign n59906 = n49831 | n49823 | n49830;
  assign n59907 = n49828 | n49829;
  assign n59908 = n49851 | n49852;
  assign n59909 = n49857 | ~n49858;
  assign n59910 = n49860 | n49861;
  assign n59911 = n49866 | ~n49867;
  assign n59912 = n49877 | n49878;
  assign n59913 = n49879 | n49880;
  assign n59914 = n49881 | ~n49882;
  assign n59915 = n49894 | n49895;
  assign n59916 = n49896 | n49897;
  assign n59917 = n49901 | n49902;
  assign n59918 = n49903 | n49904;
  assign n59919 = n49905 | ~n49906;
  assign n59920 = n49909 | n49910;
  assign n59921 = n49911 | n49912;
  assign n59922 = n49913 | ~n49914;
  assign n59923 = n49916 | ~n49917;
  assign n59924 = n49929 | n49930;
  assign n59925 = n49931 | n49932;
  assign n59926 = n49938 | ~n49939;
  assign n59927 = n49941 | ~n49942;
  assign n59928 = n49954 | n49955;
  assign n59929 = n49956 | n49957;
  assign n59930 = n49963 | ~n49964;
  assign n59931 = n49966 | ~n49967;
  assign n59932 = n49979 | n49980;
  assign n59933 = n49981 | n49982;
  assign n59934 = n49988 | ~n49989;
  assign n59935 = n49991 | ~n49992;
  assign n59936 = n50004 | n50005;
  assign n59937 = n50006 | n50007;
  assign n59938 = n50013 | ~n50014;
  assign n59939 = n50016 | ~n50017;
  assign n59940 = n50029 | n50030;
  assign n59941 = n50031 | n50032;
  assign n59942 = n50038 | ~n50039;
  assign n59943 = n50044 | ~n50045;
  assign n59944 = n50047 | ~n50048;
  assign n59945 = n50070 | n50071;
  assign n59946 = n50072 | n50073;
  assign n59947 = n50086 | n50087;
  assign n59948 = n50094 | n50095;
  assign n59949 = n50111 | n50112;
  assign n59950 = n50133 | ~n50134;
  assign n59951 = n50139 | ~n50140;
  assign n59952 = n50152 | n50153;
  assign n59953 = n50154 | n50155;
  assign n59954 = n50159 | n50160;
  assign n59955 = n50161 | n50162;
  assign n59956 = n50163 | ~n50164;
  assign n59957 = n50176 | n50177;
  assign n59958 = n50178 | n50179;
  assign n59959 = n50183 | n50184;
  assign n59960 = n50185 | n50186;
  assign n59961 = n50187 | ~n50188;
  assign n59962 = n50190 | ~n50191;
  assign n59963 = n50203 | n50204;
  assign n59964 = n50205 | n50206;
  assign n59965 = n50210 | n50211;
  assign n59966 = n50212 | n50213;
  assign n59967 = n50214 | ~n50215;
  assign n59968 = n50217 | ~n50218;
  assign n59969 = n50230 | n50231;
  assign n59970 = n50232 | n50233;
  assign n59971 = n50236 | ~n50237;
  assign n59972 = n50240 | n50241;
  assign n59973 = n50242 | n50243;
  assign n59974 = n50244 | ~n50245;
  assign n59975 = n50257 | n50258;
  assign n59976 = n50259 | n50260;
  assign n59977 = n50264 | n50265;
  assign n59978 = n50266 | n50267;
  assign n59979 = n50268 | ~n50269;
  assign n59980 = n50271 | ~n50272;
  assign n59981 = n50282 | n50283;
  assign n59982 = n50284 | n50285;
  assign n59983 = n50288 | ~n50289;
  assign n59984 = n50292 | n50293;
  assign n59985 = n50294 | n50295;
  assign n59986 = n50296 | ~n50297;
  assign n59987 = n50302 | ~n50303;
  assign n59988 = n50324 | n50325;
  assign n59989 = n50326 | n50327;
  assign n59990 = n50337 | n50338;
  assign n59991 = n50346 | n50347;
  assign n59992 = n50357 | n50358;
  assign n59993 = n50375 | n50376;
  assign n59994 = n50391 | ~n50392;
  assign n59995 = n50394 | ~n50395;
  assign n59996 = n50407 | ~n50408;
  assign n59997 = n50426 | n50427;
  assign n59998 = n50428 | n50429;
  assign n59999 = n50435 | ~n50436;
  assign n60000 = n50448 | n50449;
  assign n60001 = n50450 | n50451;
  assign n60002 = n50457 | ~n50458;
  assign n60003 = n50470 | n50471;
  assign n60004 = n50472 | n50473;
  assign n60005 = n50479 | ~n50480;
  assign n60006 = n50492 | n50493;
  assign n60007 = n50494 | n50495;
  assign n60008 = n50501 | ~n50502;
  assign n60009 = n50505 | n50506;
  assign n60010 = n50507 | n50508;
  assign n60011 = n50509 | ~n50510;
  assign n60012 = n50515 | ~n50516;
  assign n60013 = n50522 | n50523;
  assign n60014 = n50524 | n50525;
  assign n60015 = n50531 | ~n50532;
  assign n60016 = n50537 | ~n50538;
  assign n60017 = n50558 | ~n50559;
  assign n60018 = n50565 | n50566;
  assign n60019 = n50595 | n50584 | n50594;
  assign n60020 = n50616 | n50617;
  assign n60021 = n50622 | ~n50623;
  assign n60022 = n50625 | n50626;
  assign n60023 = n50631 | ~n50632;
  assign n60024 = n50642 | n50643;
  assign n60025 = n50644 | n50645;
  assign n60026 = n50646 | ~n50647;
  assign n60027 = n50662 | n50663;
  assign n60028 = n50664 | n50665;
  assign n60029 = n50671 | ~n50672;
  assign n60030 = n50674 | ~n50675;
  assign n60031 = n50687 | n50688;
  assign n60032 = n50689 | n50690;
  assign n60033 = n50696 | ~n50697;
  assign n60034 = n50699 | ~n50700;
  assign n60035 = n50712 | n50713;
  assign n60036 = n50714 | n50715;
  assign n60037 = n50721 | ~n50722;
  assign n60038 = n50724 | ~n50725;
  assign n60039 = n50737 | n50738;
  assign n60040 = n50739 | n50740;
  assign n60041 = n50746 | ~n50747;
  assign n60042 = n50749 | ~n50750;
  assign n60043 = n50762 | n50763;
  assign n60044 = n50764 | n50765;
  assign n60045 = n50771 | ~n50772;
  assign n60046 = n50777 | ~n50778;
  assign n60047 = n50780 | ~n50781;
  assign n60048 = n50801 | n50802;
  assign n60049 = n50803 | n50804;
  assign n60050 = n50814 | n50815;
  assign n60051 = n50816 | n50817;
  assign n60052 = n50828 | n50824 | n50827;
  assign n60053 = n50845 | n50846;
  assign n60054 = n50864 | n50865;
  assign n60055 = n50881 | n50882;
  assign n60056 = n50883 | n50884;
  assign n60057 = n50885 | ~n50886;
  assign n60058 = n50889 | n50890;
  assign n60059 = n50891 | n50892;
  assign n60060 = n50893 | ~n50894;
  assign n60061 = n50899 | ~n50900;
  assign n60062 = n50905 | ~n50906;
  assign n60063 = n50909 | n50910;
  assign n60064 = n50911 | n50912;
  assign n60065 = n50913 | ~n50914;
  assign n60066 = n50916 | ~n50917;
  assign n60067 = n50929 | n50930;
  assign n60068 = n50931 | n50932;
  assign n60069 = n50936 | n50937;
  assign n60070 = n50938 | n50939;
  assign n60071 = n50940 | ~n50941;
  assign n60072 = n50943 | ~n50944;
  assign n60073 = n50956 | n50957;
  assign n60074 = n50958 | n50959;
  assign n60075 = n50962 | ~n50963;
  assign n60076 = n50966 | n50967;
  assign n60077 = n50968 | n50969;
  assign n60078 = n50970 | ~n50971;
  assign n60079 = n50983 | n50984;
  assign n60080 = n50985 | n50986;
  assign n60081 = n50990 | n50991;
  assign n60082 = n50992 | n50993;
  assign n60083 = n50994 | ~n50995;
  assign n60084 = n50997 | ~n50998;
  assign n60085 = n51008 | n51009;
  assign n60086 = n51010 | n51011;
  assign n60087 = n51014 | ~n51015;
  assign n60088 = n51018 | n51019;
  assign n60089 = n51020 | n51021;
  assign n60090 = n51022 | ~n51023;
  assign n60091 = n51028 | ~n51029;
  assign n60092 = n51050 | n51051;
  assign n60093 = n51052 | n51053;
  assign n60094 = n51065 | n51066;
  assign n60095 = n51081 | n51082;
  assign n60096 = n51085 | n51086;
  assign n60097 = n51105 | n51102 | n51104;
  assign n60098 = n51120 | ~n51121;
  assign n60099 = n51133 | ~n51134;
  assign n60100 = n51142 | ~n51143;
  assign n60101 = n51155 | n51156;
  assign n60102 = n51157 | n51158;
  assign n60103 = n51164 | ~n51165;
  assign n60104 = n51177 | n51178;
  assign n60105 = n51179 | n51180;
  assign n60106 = n51186 | ~n51187;
  assign n60107 = n51199 | n51200;
  assign n60108 = n51201 | n51202;
  assign n60109 = n51208 | ~n51209;
  assign n60110 = n51212 | n51213;
  assign n60111 = n51214 | n51215;
  assign n60112 = n51216 | ~n51217;
  assign n60113 = n51222 | ~n51223;
  assign n60114 = n51229 | n51230;
  assign n60115 = n51231 | n51232;
  assign n60116 = n51238 | ~n51239;
  assign n60117 = n51244 | ~n51245;
  assign n60118 = n51264 | n51265;
  assign n60119 = n51266 | n51267;
  assign n60120 = n51271 | n51272;
  assign n60121 = n51283 | n51284;
  assign n60122 = n51303 | n51295 | n51302;
  assign n60123 = n51304 | n51305;
  assign n60124 = n51326 | n51327;
  assign n60125 = n51339 | n51340;
  assign n60126 = n51345 | ~n51346;
  assign n60127 = n51348 | ~n51349;
  assign n60128 = n51365 | n51366;
  assign n60129 = n51367 | n51368;
  assign n60130 = n51372 | n51373;
  assign n60131 = n51374 | n51375;
  assign n60132 = n51376 | ~n51377;
  assign n60133 = n51382 | ~n51383;
  assign n60134 = n51385 | ~n51386;
  assign n60135 = n51398 | n51399;
  assign n60136 = n51400 | n51401;
  assign n60137 = n51407 | ~n51408;
  assign n60138 = n51410 | ~n51411;
  assign n60139 = n51423 | n51424;
  assign n60140 = n51425 | n51426;
  assign n60141 = n51432 | ~n51433;
  assign n60142 = n51435 | ~n51436;
  assign n60143 = n51448 | n51449;
  assign n60144 = n51450 | n51451;
  assign n60145 = n51457 | ~n51458;
  assign n60146 = n51463 | ~n51464;
  assign n60147 = n51466 | ~n51467;
  assign n60148 = n51489 | n51490;
  assign n60149 = n51491 | n51492;
  assign n60150 = n51497 | n51498;
  assign n60151 = n51517 | n51518;
  assign n60152 = n51539 | ~n51540;
  assign n60153 = n51545 | ~n51546;
  assign n60154 = n51558 | n51559;
  assign n60155 = n51560 | n51561;
  assign n60156 = n51565 | n51566;
  assign n60157 = n51567 | n51568;
  assign n60158 = n51569 | ~n51570;
  assign n60159 = n51582 | n51583;
  assign n60160 = n51584 | n51585;
  assign n60161 = n51588 | ~n51589;
  assign n60162 = n51592 | n51593;
  assign n60163 = n51594 | n51595;
  assign n60164 = n51596 | ~n51597;
  assign n60165 = n51609 | n51610;
  assign n60166 = n51611 | n51612;
  assign n60167 = n51616 | n51617;
  assign n60168 = n51618 | n51619;
  assign n60169 = n51620 | ~n51621;
  assign n60170 = n51623 | ~n51624;
  assign n60171 = n51634 | n51635;
  assign n60172 = n51636 | n51637;
  assign n60173 = n51640 | ~n51641;
  assign n60174 = n51644 | n51645;
  assign n60175 = n51646 | n51647;
  assign n60176 = n51648 | ~n51649;
  assign n60177 = n51654 | ~n51655;
  assign n60178 = n51676 | n51677;
  assign n60179 = n51678 | n51679;
  assign n60180 = n51690 | n51691;
  assign n60181 = n51695 | n51696;
  assign n60182 = n51711 | n51712;
  assign n60183 = n51731 | n51732;
  assign n60184 = n51747 | ~n51748;
  assign n60185 = n51750 | ~n51751;
  assign n60186 = n51763 | ~n51764;
  assign n60187 = n51782 | n51783;
  assign n60188 = n51784 | n51785;
  assign n60189 = n51791 | ~n51792;
  assign n60190 = n51804 | n51805;
  assign n60191 = n51806 | n51807;
  assign n60192 = n51813 | ~n51814;
  assign n60193 = n51817 | n51818;
  assign n60194 = n51819 | n51820;
  assign n60195 = n51821 | ~n51822;
  assign n60196 = n51827 | ~n51828;
  assign n60197 = n51834 | n51835;
  assign n60198 = n51836 | n51837;
  assign n60199 = n51843 | ~n51844;
  assign n60200 = n51849 | ~n51850;
  assign n60201 = n51870 | ~n51871;
  assign n60202 = n51877 | n51878;
  assign n60203 = n51883 | n51884;
  assign n60204 = n51901 | n51902;
  assign n60205 = n51920 | n51921;
  assign n60206 = n51926 | ~n51927;
  assign n60207 = n51929 | n51930;
  assign n60208 = n51935 | ~n51936;
  assign n60209 = n51946 | n51947;
  assign n60210 = n51948 | n51949;
  assign n60211 = n51950 | ~n51951;
  assign n60212 = n51966 | n51967;
  assign n60213 = n51968 | n51969;
  assign n60214 = n51975 | ~n51976;
  assign n60215 = n51978 | ~n51979;
  assign n60216 = n51991 | n51992;
  assign n60217 = n51993 | n51994;
  assign n60218 = n52000 | ~n52001;
  assign n60219 = n52003 | ~n52004;
  assign n60220 = n52016 | n52017;
  assign n60221 = n52018 | n52019;
  assign n60222 = n52025 | ~n52026;
  assign n60223 = n52031 | ~n52032;
  assign n60224 = n52034 | ~n52035;
  assign n60225 = n52055 | n52056;
  assign n60226 = n52057 | n52058;
  assign n60227 = n52068 | n52069;
  assign n60228 = n52070 | n52071;
  assign n60229 = n52074 | ~n52075;
  assign n60230 = n52078 | n52079;
  assign n60231 = n52080 | n52081;
  assign n60232 = n52082 | ~n52083;
  assign n60233 = n52092 | n52093;
  assign n60234 = n52094 | n52095;
  assign n60235 = n52100 | n52101;
  assign n60236 = n52105 | n52106;
  assign n60237 = n52111 | n52112;
  assign n60238 = n52127 | n52128;
  assign n60239 = n52144 | n52145;
  assign n60240 = n52146 | n52147;
  assign n60241 = n52148 | ~n52149;
  assign n60242 = n52152 | n52153;
  assign n60243 = n52154 | n52155;
  assign n60244 = n52156 | ~n52157;
  assign n60245 = n52162 | ~n52163;
  assign n60246 = n52168 | ~n52169;
  assign n60247 = n52174 | ~n52175;
  assign n60248 = n52180 | ~n52181;
  assign n60249 = n52191 | n52192;
  assign n60250 = n52193 | n52194;
  assign n60251 = n52197 | ~n52198;
  assign n60252 = n52201 | n52202;
  assign n60253 = n52203 | n52204;
  assign n60254 = n52205 | ~n52206;
  assign n60255 = n52211 | ~n52212;
  assign n60256 = n52233 | n52234;
  assign n60257 = n52235 | n52236;
  assign n60258 = n52257 | n52251 | n52256;
  assign n60259 = n52278 | n52279;
  assign n60260 = n52294 | ~n52295;
  assign n60261 = n52307 | ~n52308;
  assign n60262 = n52316 | ~n52317;
  assign n60263 = n52329 | n52330;
  assign n60264 = n52331 | n52332;
  assign n60265 = n52338 | ~n52339;
  assign n60266 = n52344 | ~n52345;
  assign n60267 = n52347 | n52348;
  assign n60268 = n52349 | n52350;
  assign n60269 = n52352 | ~n52353;
  assign n60270 = n52359 | n52360;
  assign n60271 = n52361 | n52362;
  assign n60272 = n52368 | ~n52369;
  assign n60273 = n52372 | n52373;
  assign n60274 = n52374 | n52375;
  assign n60275 = n52376 | ~n52377;
  assign n60276 = n52385 | ~n52386;
  assign n60277 = n52398 | n52399;
  assign n60278 = n52400 | n52401;
  assign n60279 = n52413 | n52414;
  assign n60280 = n52431 | n52432;
  assign n60281 = n52444 | n52445;
  assign n60282 = n52450 | ~n52451;
  assign n60283 = n52453 | ~n52454;
  assign n60284 = n52470 | n52471;
  assign n60285 = n52472 | n52473;
  assign n60286 = n52477 | n52478;
  assign n60287 = n52479 | n52480;
  assign n60288 = n52481 | ~n52482;
  assign n60289 = n52487 | ~n52488;
  assign n60290 = n52490 | ~n52491;
  assign n60291 = n52503 | n52504;
  assign n60292 = n52505 | n52506;
  assign n60293 = n52512 | ~n52513;
  assign n60294 = n52518 | ~n52519;
  assign n60295 = n52521 | ~n52522;
  assign n60296 = n52543 | n52544;
  assign n60297 = n52545 | n52546;
  assign n60298 = n52555 | n52556;
  assign n60299 = n52571 | n52562 | n52570;
  assign n60300 = n52579 | n52576 | n52578;
  assign n60301 = n52598 | n52599;
  assign n60302 = n52620 | ~n52621;
  assign n60303 = n52633 | n52634;
  assign n60304 = n52635 | n52636;
  assign n60305 = n52642 | ~n52643;
  assign n60306 = n52646 | n52647;
  assign n60307 = n52648 | n52649;
  assign n60308 = n52650 | ~n52651;
  assign n60309 = n52661 | n52662;
  assign n60310 = n52663 | n52664;
  assign n60311 = n52667 | ~n52668;
  assign n60312 = n52671 | n52672;
  assign n60313 = n52673 | n52674;
  assign n60314 = n52675 | ~n52676;
  assign n60315 = n52681 | ~n52682;
  assign n60316 = n52698 | n52699;
  assign n60317 = n52713 | n52714;
  assign n60318 = n52716 | n52717;
  assign n60319 = n52733 | n52734;
  assign n60320 = n52749 | ~n52750;
  assign n60321 = n52752 | ~n52753;
  assign n60322 = n52765 | ~n52766;
  assign n60323 = n52774 | ~n52775;
  assign n60324 = n52787 | n52788;
  assign n60325 = n52789 | n52790;
  assign n60326 = n52796 | ~n52797;
  assign n60327 = n52803 | n52804;
  assign n60328 = n52805 | n52806;
  assign n60329 = n52812 | ~n52813;
  assign n60330 = n52816 | n52817;
  assign n60331 = n52818 | n52819;
  assign n60332 = n52820 | ~n52821;
  assign n60333 = n52829 | ~n52830;
  assign n60334 = n52842 | n52843;
  assign n60335 = n52844 | n52845;
  assign n60336 = n52859 | n52855 | n52858;
  assign n60337 = n52875 | n52867 | n52874;
  assign n60338 = n52893 | n52894;
  assign n60339 = n52899 | ~n52900;
  assign n60340 = n52902 | n52903;
  assign n60341 = n52908 | ~n52909;
  assign n60342 = n52919 | n52920;
  assign n60343 = n52921 | n52922;
  assign n60344 = n52923 | ~n52924;
  assign n60345 = n52936 | n52937;
  assign n60346 = n52938 | n52939;
  assign n60347 = n52943 | n52944;
  assign n60348 = n52945 | n52946;
  assign n60349 = n52947 | ~n52948;
  assign n60350 = n52951 | n52952;
  assign n60351 = n52953 | n52954;
  assign n60352 = n52955 | ~n52956;
  assign n60353 = n52961 | ~n52962;
  assign n60354 = n52964 | ~n52965;
  assign n60355 = n52984 | n52985;
  assign n60356 = n52986 | n52987;
  assign n60357 = n52991 | n52992;
  assign n60358 = n52993 | n52994;
  assign n60359 = n52995 | ~n52996;
  assign n60360 = n53010 | n53019 | n53029 | n53030;
  assign n60361 = n53033 | n53034;
  assign n60362 = n53048 | n53049;
  assign n60363 = n53070 | ~n53071;
  assign n60364 = n53083 | n53084;
  assign n60365 = n53085 | n53086;
  assign n60366 = n53092 | ~n53093;
  assign n60367 = n53098 | ~n53099;
  assign n60368 = n53101 | ~n53102;
  assign n60369 = n53144 | n53134 | n53143;
  assign n60370 = n53147 | n53148;
  assign n60371 = n53165 | n53166;
  assign n60372 = n53181 | ~n53182;
  assign n60373 = n53184 | ~n53185;
  assign n60374 = n53197 | ~n53198;
  assign n60375 = n53206 | ~n53207;
  assign n60376 = n53213 | n53214;
  assign n60377 = n53215 | n53216;
  assign n60378 = n53222 | ~n53223;
  assign n60379 = n53228 | ~n53229;
  assign n60380 = n53241 | n53242;
  assign n60381 = n53245 | n53246;
  assign n60382 = n53248 | n53249;
  assign n60383 = n53257 | n53252 | n53256;
  assign n60384 = n53262 | n53263;
  assign n60385 = n53268 | ~n53269;
  assign n60386 = n53271 | n53272;
  assign n60387 = n53277 | ~n53278;
  assign n60388 = n53288 | n53289;
  assign n60389 = n53290 | n53291;
  assign n60390 = n53292 | ~n53293;
  assign n60391 = n53305 | n53306;
  assign n60392 = n53307 | n53308;
  assign n60393 = n53312 | n53313;
  assign n60394 = n53314 | n53315;
  assign n60395 = n53316 | ~n53317;
  assign n60396 = n53322 | ~n53323;
  assign n60397 = ~n53349 | n53345 | ~n53348;
  assign n60398 = n53365 | n53366;
  assign n60399 = n53389 | n53390;
  assign n60400 = ~n53420 | n53395 | ~n53419;
  assign n60401 = n53415 | n53416;
  assign n60402 = n53438 | n53431 | n53437;
  assign po0  = ~n59391;
  assign po31  = ~n60402;
endmodule
