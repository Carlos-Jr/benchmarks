module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n181, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n484, n486, n487, n488,
    n489, n490, n491, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673,
    n675, n676, n677;
  assign n23 = ~pi08 & ~pi10;
  assign n24 = pi04 & n23;
  assign n25 = pi08 & ~pi10;
  assign n26 = pi10 & ~pi11;
  assign n27 = ~pi09 & ~n26;
  assign n28 = ~n25 & n27;
  assign n29 = ~n24 & ~n28;
  assign n30 = pi09 & pi11;
  assign n31 = ~pi10 & ~n30;
  assign n32 = ~pi13 & n31;
  assign n33 = ~pi08 & n32;
  assign n34 = ~pi00 & n33;
  assign n35 = pi00 & ~pi04;
  assign n36 = ~pi00 & pi04;
  assign n37 = n26 & n36;
  assign n38 = ~n35 & ~n37;
  assign n39 = ~pi08 & pi09;
  assign n40 = pi13 & n39;
  assign n41 = ~n38 & n40;
  assign n42 = ~pi08 & ~pi09;
  assign n43 = pi08 & pi09;
  assign n44 = ~n42 & ~n43;
  assign n45 = ~pi10 & pi11;
  assign n46 = ~n44 & n45;
  assign n47 = pi13 & n46;
  assign n48 = ~pi08 & pi10;
  assign n49 = ~pi09 & ~pi11;
  assign n50 = n48 & n49;
  assign n51 = ~n47 & ~n50;
  assign n52 = pi00 & pi04;
  assign n53 = ~n51 & n52;
  assign n54 = ~pi00 & ~pi04;
  assign n55 = ~pi10 & ~pi11;
  assign n56 = ~pi13 & ~n55;
  assign n57 = pi08 & ~pi09;
  assign n58 = ~pi10 & pi13;
  assign n59 = n57 & ~n58;
  assign n60 = ~n56 & n59;
  assign n61 = ~n54 & n60;
  assign n62 = ~n26 & n40;
  assign n63 = n26 & n43;
  assign n64 = ~n62 & ~n63;
  assign n65 = ~pi09 & pi11;
  assign n66 = pi08 & pi10;
  assign n67 = ~pi13 & n66;
  assign n68 = n65 & n67;
  assign n69 = n64 & ~n68;
  assign n70 = ~pi04 & ~n69;
  assign n71 = ~n61 & ~n70;
  assign n72 = ~n53 & n71;
  assign n73 = ~n41 & n72;
  assign n74 = ~n34 & n73;
  assign n75 = ~n29 & ~n74;
  assign n76 = ~pi08 & n26;
  assign n77 = n54 & n76;
  assign n78 = pi00 & ~n73;
  assign n79 = n66 & n78;
  assign n80 = ~pi08 & pi11;
  assign n81 = pi04 & n80;
  assign n82 = ~pi11 & ~n48;
  assign n83 = n52 & ~n82;
  assign n84 = ~n81 & ~n83;
  assign n85 = ~n79 & n84;
  assign n86 = ~n77 & n85;
  assign n87 = pi09 & ~n86;
  assign n88 = pi08 & n55;
  assign n89 = ~n48 & ~n88;
  assign n90 = n74 & ~n89;
  assign n91 = pi08 & n26;
  assign n92 = ~pi04 & n91;
  assign n93 = pi04 & n25;
  assign n94 = ~pi00 & ~n93;
  assign n95 = ~n52 & ~n94;
  assign n96 = pi11 & n95;
  assign n97 = ~n92 & ~n96;
  assign n98 = ~n90 & n97;
  assign n99 = ~pi09 & ~n98;
  assign n100 = ~n87 & ~n99;
  assign n101 = ~n75 & n100;
  assign n102 = ~pi10 & ~n42;
  assign n103 = pi00 & pi11;
  assign n104 = ~n102 & n103;
  assign n105 = n101 & ~n104;
  assign n106 = ~pi13 & ~n105;
  assign n107 = ~pi11 & n43;
  assign n108 = n58 & n107;
  assign n109 = ~pi13 & n48;
  assign n110 = n65 & n109;
  assign n111 = ~n108 & ~n110;
  assign n112 = ~n106 & n111;
  assign n113 = ~pi00 & n74;
  assign n114 = ~pi08 & pi13;
  assign n115 = n30 & n114;
  assign n116 = ~n113 & n115;
  assign n117 = pi13 & n26;
  assign n118 = n52 & n57;
  assign n119 = n43 & n78;
  assign n120 = ~n118 & ~n119;
  assign n121 = n42 & n74;
  assign n122 = n120 & ~n121;
  assign n123 = n117 & ~n122;
  assign n124 = ~n116 & ~n123;
  assign n125 = n23 & n30;
  assign n126 = pi13 & n125;
  assign n127 = n52 & n126;
  assign n128 = n57 & n117;
  assign n129 = n124 & n128;
  assign n130 = ~n127 & ~n129;
  assign n131 = n125 & n130;
  assign n132 = ~pi00 & n50;
  assign n133 = ~n131 & ~n132;
  assign n134 = ~n124 & ~n133;
  assign n135 = pi09 & ~n74;
  assign n136 = ~pi00 & ~n135;
  assign n137 = ~pi09 & n74;
  assign n138 = pi11 & ~n137;
  assign n139 = n23 & ~n138;
  assign n140 = ~n136 & n139;
  assign n141 = pi11 & ~n102;
  assign n142 = ~pi00 & n141;
  assign n143 = n26 & n57;
  assign n144 = n130 & n143;
  assign n145 = ~n142 & ~n144;
  assign n146 = ~n74 & ~n145;
  assign n147 = n43 & n45;
  assign n148 = n26 & n39;
  assign n149 = ~n147 & ~n148;
  assign n150 = ~n43 & n103;
  assign n151 = pi08 & ~n130;
  assign n152 = n49 & n151;
  assign n153 = ~n150 & ~n152;
  assign n154 = pi10 & ~n153;
  assign n155 = n149 & ~n154;
  assign n156 = n74 & ~n155;
  assign n157 = pi00 & ~pi08;
  assign n158 = n124 & n157;
  assign n159 = ~n93 & ~n158;
  assign n160 = n49 & ~n159;
  assign n161 = n125 & ~n130;
  assign n162 = ~n63 & ~n161;
  assign n163 = n124 & ~n162;
  assign n164 = pi10 & n43;
  assign n165 = ~pi00 & n164;
  assign n166 = pi11 & n165;
  assign n167 = ~n163 & ~n166;
  assign n168 = ~n160 & n167;
  assign n169 = ~n156 & n168;
  assign n170 = ~n146 & n169;
  assign n171 = ~pi09 & n25;
  assign n172 = ~n52 & ~n54;
  assign n173 = n171 & n172;
  assign n174 = n170 & ~n173;
  assign n175 = ~n140 & n174;
  assign n176 = ~n134 & n175;
  assign n177 = pi13 & ~n176;
  assign n178 = pi12 & ~n177;
  assign n179 = ~pi12 & n177;
  assign n180 = ~n178 & ~n179;
  assign n181 = pi13 & n180;
  assign po0 = ~n112 | n181;
  assign n183 = ~pi01 & n33;
  assign n184 = ~pi05 & ~n69;
  assign n185 = pi01 & pi05;
  assign n186 = n37 & n114;
  assign n187 = ~pi09 & n26;
  assign n188 = ~n46 & ~n187;
  assign n189 = pi13 & ~n188;
  assign n190 = ~n50 & ~n189;
  assign n191 = ~n186 & n190;
  assign n192 = n185 & ~n191;
  assign n193 = ~pi09 & pi10;
  assign n194 = n103 & n193;
  assign n195 = ~pi01 & ~pi05;
  assign n196 = n36 & ~n195;
  assign n197 = pi09 & ~n196;
  assign n198 = pi01 & ~pi05;
  assign n199 = ~pi01 & pi05;
  assign n200 = n26 & n199;
  assign n201 = ~n36 & ~n200;
  assign n202 = ~n198 & n201;
  assign n203 = n197 & ~n202;
  assign n204 = ~n194 & ~n203;
  assign n205 = n114 & ~n204;
  assign n206 = n60 & ~n195;
  assign n207 = ~n205 & ~n206;
  assign n208 = ~n192 & n207;
  assign n209 = ~n184 & n208;
  assign n210 = ~n183 & n209;
  assign n211 = n164 & ~n210;
  assign n212 = ~n141 & ~n211;
  assign n213 = pi01 & ~n212;
  assign n214 = pi05 & n23;
  assign n215 = ~n28 & ~n214;
  assign n216 = ~n210 & ~n215;
  assign n217 = n76 & n195;
  assign n218 = pi01 & ~n82;
  assign n219 = ~n80 & ~n218;
  assign n220 = pi05 & ~n219;
  assign n221 = ~n217 & ~n220;
  assign n222 = pi09 & ~n221;
  assign n223 = ~n89 & n210;
  assign n224 = ~pi05 & n91;
  assign n225 = pi05 & n25;
  assign n226 = ~pi01 & ~n225;
  assign n227 = ~n185 & ~n226;
  assign n228 = pi11 & n227;
  assign n229 = ~n224 & ~n228;
  assign n230 = ~n223 & n229;
  assign n231 = ~pi09 & ~n230;
  assign n232 = ~n222 & ~n231;
  assign n233 = ~n216 & n232;
  assign n234 = ~n213 & n233;
  assign n235 = ~pi13 & ~n234;
  assign n236 = n111 & ~n235;
  assign n237 = pi10 & ~n43;
  assign n238 = ~n42 & ~n237;
  assign n239 = pi11 & ~n238;
  assign n240 = n78 & ~n210;
  assign n241 = ~n78 & n210;
  assign n242 = ~n240 & ~n241;
  assign n243 = n239 & n242;
  assign n244 = ~pi01 & n210;
  assign n245 = n115 & ~n244;
  assign n246 = ~pi05 & ~pi09;
  assign n247 = pi01 & ~n246;
  assign n248 = pi08 & ~n247;
  assign n249 = pi09 & n210;
  assign n250 = ~pi08 & ~n210;
  assign n251 = n117 & ~n250;
  assign n252 = ~n249 & n251;
  assign n253 = ~n248 & n252;
  assign n254 = ~n245 & ~n253;
  assign n255 = pi00 & ~n124;
  assign n256 = n254 & ~n255;
  assign n257 = ~n124 & ~n254;
  assign n258 = pi00 & n257;
  assign n259 = ~n256 & ~n258;
  assign n260 = n50 & n259;
  assign n261 = ~n243 & ~n260;
  assign n262 = ~pi01 & ~n261;
  assign n263 = n74 & n210;
  assign n264 = ~n149 & n263;
  assign n265 = n52 & n195;
  assign n266 = n171 & n265;
  assign n267 = ~pi00 & ~pi01;
  assign n268 = n164 & n267;
  assign n269 = ~n266 & ~n268;
  assign n270 = pi11 & ~n269;
  assign n271 = n103 & n164;
  assign n272 = ~pi05 & n171;
  assign n273 = ~n52 & n272;
  assign n274 = ~n26 & ~n238;
  assign n275 = ~n242 & n274;
  assign n276 = ~n43 & n55;
  assign n277 = ~n275 & ~n276;
  assign n278 = ~n273 & n277;
  assign n279 = ~n271 & n278;
  assign n280 = pi01 & ~n279;
  assign n281 = n124 & n254;
  assign n282 = ~n257 & ~n281;
  assign n283 = n164 & ~n282;
  assign n284 = pi09 & n23;
  assign n285 = ~n210 & n284;
  assign n286 = ~n283 & ~n285;
  assign n287 = ~pi11 & ~n286;
  assign n288 = ~n52 & ~n199;
  assign n289 = n52 & ~n185;
  assign n290 = n171 & ~n289;
  assign n291 = ~n288 & n290;
  assign n292 = ~pi11 & n39;
  assign n293 = ~n147 & ~n292;
  assign n294 = ~n74 & ~n210;
  assign n295 = ~n293 & n294;
  assign n296 = ~n291 & ~n295;
  assign n297 = ~n287 & n296;
  assign n298 = ~n280 & n297;
  assign n299 = n126 & n185;
  assign n300 = n128 & n254;
  assign n301 = ~n299 & ~n300;
  assign n302 = ~n124 & n127;
  assign n303 = ~n301 & n302;
  assign n304 = n301 & ~n302;
  assign n305 = ~n303 & ~n304;
  assign n306 = n254 & ~n305;
  assign n307 = ~n254 & n305;
  assign n308 = ~n306 & ~n307;
  assign n309 = n125 & n308;
  assign n310 = n298 & ~n309;
  assign n311 = ~n270 & n310;
  assign n312 = ~n74 & ~n130;
  assign n313 = ~n301 & n312;
  assign n314 = n301 & ~n312;
  assign n315 = ~n313 & ~n314;
  assign n316 = n210 & ~n315;
  assign n317 = ~n210 & n315;
  assign n318 = ~n316 & ~n317;
  assign n319 = n66 & n318;
  assign n320 = ~pi08 & ~n259;
  assign n321 = pi01 & n320;
  assign n322 = ~n225 & ~n321;
  assign n323 = ~n319 & n322;
  assign n324 = n49 & ~n323;
  assign n325 = n311 & ~n324;
  assign n326 = ~n264 & n325;
  assign n327 = ~n262 & n326;
  assign n328 = n179 & ~n327;
  assign n329 = ~n179 & n327;
  assign n330 = pi13 & ~n329;
  assign n331 = ~n328 & n330;
  assign po1 = ~n236 | n331;
  assign n333 = pi02 & pi11;
  assign n334 = ~pi06 & ~pi09;
  assign n335 = n102 & ~n334;
  assign n336 = n333 & ~n335;
  assign n337 = pi09 & n80;
  assign n338 = ~pi02 & n65;
  assign n339 = n25 & n338;
  assign n340 = ~n337 & ~n339;
  assign n341 = pi06 & ~n340;
  assign n342 = pi02 & pi06;
  assign n343 = ~n82 & n342;
  assign n344 = ~pi02 & ~pi06;
  assign n345 = n76 & n344;
  assign n346 = ~n343 & ~n345;
  assign n347 = pi09 & ~n346;
  assign n348 = ~pi06 & ~n69;
  assign n349 = n60 & ~n344;
  assign n350 = ~n36 & ~n199;
  assign n351 = ~n198 & ~n350;
  assign n352 = pi06 & n26;
  assign n353 = ~n351 & ~n352;
  assign n354 = ~pi02 & pi09;
  assign n355 = pi06 & n351;
  assign n356 = n354 & ~n355;
  assign n357 = ~n353 & n356;
  assign n358 = pi01 & n65;
  assign n359 = pi10 & n358;
  assign n360 = ~n357 & ~n359;
  assign n361 = ~pi06 & ~n351;
  assign n362 = n26 & n355;
  assign n363 = ~n361 & ~n362;
  assign n364 = ~n334 & ~n363;
  assign n365 = pi02 & n364;
  assign n366 = n360 & ~n365;
  assign n367 = n114 & ~n366;
  assign n368 = ~n190 & n342;
  assign n369 = ~pi02 & n33;
  assign n370 = ~n368 & ~n369;
  assign n371 = ~n367 & n370;
  assign n372 = ~n349 & n371;
  assign n373 = ~n348 & n372;
  assign n374 = ~n89 & n373;
  assign n375 = ~pi06 & n91;
  assign n376 = ~n374 & ~n375;
  assign n377 = ~pi09 & ~n376;
  assign n378 = ~n347 & ~n377;
  assign n379 = ~n341 & n378;
  assign n380 = pi06 & n23;
  assign n381 = pi02 & n164;
  assign n382 = ~n380 & ~n381;
  assign n383 = ~n28 & n382;
  assign n384 = ~n373 & ~n383;
  assign n385 = n379 & ~n384;
  assign n386 = ~n336 & n385;
  assign n387 = ~pi13 & ~n386;
  assign n388 = n111 & ~n387;
  assign n389 = ~pi02 & n373;
  assign n390 = n115 & ~n389;
  assign n391 = n42 & n373;
  assign n392 = pi09 & n373;
  assign n393 = pi02 & ~n392;
  assign n394 = ~n334 & n393;
  assign n395 = pi08 & n394;
  assign n396 = ~n391 & ~n395;
  assign n397 = n117 & ~n396;
  assign n398 = ~n390 & ~n397;
  assign n399 = pi01 & ~n256;
  assign n400 = ~n258 & ~n399;
  assign n401 = ~n398 & n400;
  assign n402 = n398 & ~n400;
  assign n403 = ~n401 & ~n402;
  assign n404 = n50 & ~n403;
  assign n405 = pi01 & ~n241;
  assign n406 = ~n240 & ~n405;
  assign n407 = n239 & ~n373;
  assign n408 = n406 & n407;
  assign n409 = ~n404 & ~n408;
  assign n410 = ~pi02 & ~n409;
  assign n411 = ~pi08 & n403;
  assign n412 = pi02 & n411;
  assign n413 = pi06 & n25;
  assign n414 = n126 & n342;
  assign n415 = n128 & n398;
  assign n416 = ~n414 & ~n415;
  assign n417 = n373 & n416;
  assign n418 = ~n373 & ~n416;
  assign n419 = ~n417 & ~n418;
  assign n420 = ~n210 & ~n314;
  assign n421 = ~n313 & ~n420;
  assign n422 = n419 & ~n421;
  assign n423 = ~n419 & n421;
  assign n424 = n66 & ~n423;
  assign n425 = ~n422 & n424;
  assign n426 = ~n413 & ~n425;
  assign n427 = ~n412 & n426;
  assign n428 = n49 & ~n427;
  assign n429 = ~n373 & ~n406;
  assign n430 = n274 & n429;
  assign n431 = ~n276 & ~n430;
  assign n432 = pi02 & ~n431;
  assign n433 = ~n267 & n333;
  assign n434 = n281 & n398;
  assign n435 = ~n281 & ~n398;
  assign n436 = ~n434 & ~n435;
  assign n437 = ~pi11 & ~n436;
  assign n438 = ~n433 & ~n437;
  assign n439 = ~pi02 & n267;
  assign n440 = pi11 & n439;
  assign n441 = n438 & ~n440;
  assign n442 = n164 & ~n441;
  assign n443 = ~pi10 & n292;
  assign n444 = n263 & ~n443;
  assign n445 = ~n293 & ~n444;
  assign n446 = ~n373 & n445;
  assign n447 = ~n442 & ~n446;
  assign n448 = ~n432 & n447;
  assign n449 = ~n428 & n448;
  assign n450 = ~n254 & ~n304;
  assign n451 = ~n303 & ~n450;
  assign n452 = n416 & n451;
  assign n453 = ~n416 & ~n451;
  assign n454 = ~n452 & ~n453;
  assign n455 = n398 & ~n454;
  assign n456 = ~n398 & n454;
  assign n457 = ~n455 & ~n456;
  assign n458 = n125 & n457;
  assign n459 = n449 & ~n458;
  assign n460 = ~n410 & n459;
  assign n461 = ~n52 & ~n185;
  assign n462 = ~n195 & ~n461;
  assign n463 = ~n342 & ~n344;
  assign n464 = ~n462 & ~n463;
  assign n465 = n171 & ~n464;
  assign n466 = pi11 & n344;
  assign n467 = ~n342 & ~n466;
  assign n468 = n462 & n467;
  assign n469 = n465 & ~n468;
  assign n470 = n460 & ~n469;
  assign n471 = n264 & n373;
  assign n472 = ~pi02 & n406;
  assign n473 = n274 & n406;
  assign n474 = ~pi02 & n239;
  assign n475 = ~n473 & ~n474;
  assign n476 = n373 & ~n475;
  assign n477 = ~n472 & n476;
  assign n478 = ~n471 & ~n477;
  assign n479 = n470 & n478;
  assign n480 = pi13 & ~n479;
  assign n481 = n328 & n480;
  assign n482 = ~n328 & ~n480;
  assign n483 = pi13 & ~n482;
  assign n484 = ~n481 & n483;
  assign po2 = ~n388 | n484;
  assign n486 = pi03 & pi11;
  assign n487 = ~pi07 & ~pi09;
  assign n488 = n102 & ~n487;
  assign n489 = n486 & ~n488;
  assign n490 = pi07 & n23;
  assign n491 = ~n28 & ~n490;
  assign po5 = pi03 & pi07;
  assign n493 = n189 & po5;
  assign n494 = ~pi03 & ~pi07;
  assign n495 = n60 & ~n494;
  assign n496 = pi02 & ~n355;
  assign n497 = ~n361 & ~n496;
  assign n498 = pi09 & ~n497;
  assign n499 = pi03 & n498;
  assign n500 = n114 & n499;
  assign n501 = n69 & ~n500;
  assign n502 = ~pi07 & ~n501;
  assign n503 = n117 & n497;
  assign n504 = ~n187 & ~n503;
  assign n505 = po5 & ~n504;
  assign n506 = pi07 & n498;
  assign n507 = n117 & n506;
  assign n508 = ~n32 & ~n507;
  assign n509 = ~pi03 & ~n508;
  assign n510 = n193 & n333;
  assign n511 = pi09 & n497;
  assign n512 = n494 & n511;
  assign n513 = ~n510 & ~n512;
  assign n514 = pi13 & ~n513;
  assign n515 = ~n509 & ~n514;
  assign n516 = ~n505 & n515;
  assign n517 = ~pi08 & ~n516;
  assign n518 = ~n502 & ~n517;
  assign n519 = ~n495 & n518;
  assign n520 = ~n493 & n519;
  assign n521 = ~n491 & ~n520;
  assign n522 = ~pi03 & n57;
  assign n523 = n45 & n522;
  assign n524 = ~n337 & ~n523;
  assign n525 = pi07 & ~n524;
  assign n526 = ~n89 & n520;
  assign n527 = ~pi07 & n91;
  assign n528 = ~n526 & ~n527;
  assign n529 = ~pi09 & ~n528;
  assign n530 = n76 & n494;
  assign n531 = ~n82 & po5;
  assign n532 = pi03 & ~n520;
  assign n533 = n66 & n532;
  assign n534 = ~n531 & ~n533;
  assign n535 = ~n530 & n534;
  assign n536 = pi09 & ~n535;
  assign n537 = ~n529 & ~n536;
  assign n538 = ~n525 & n537;
  assign n539 = ~n521 & n538;
  assign n540 = ~n489 & n539;
  assign n541 = ~pi13 & ~n540;
  assign n542 = n111 & ~n541;
  assign n543 = n263 & n373;
  assign n544 = ~n443 & n543;
  assign n545 = ~n293 & ~n544;
  assign n546 = ~n520 & n545;
  assign n547 = n471 & n520;
  assign n548 = n373 & n406;
  assign n549 = pi02 & ~n548;
  assign n550 = ~n429 & ~n549;
  assign n551 = ~n520 & n550;
  assign n552 = n520 & ~n550;
  assign n553 = ~n551 & ~n552;
  assign n554 = n239 & ~n553;
  assign n555 = ~n342 & ~n462;
  assign n556 = ~n344 & ~n555;
  assign n557 = pi07 & n171;
  assign n558 = ~n556 & n557;
  assign n559 = ~n554 & ~n558;
  assign n560 = ~pi03 & ~n559;
  assign n561 = pi07 & ~n556;
  assign n562 = ~pi07 & n556;
  assign n563 = pi03 & ~n562;
  assign n564 = n171 & n563;
  assign n565 = ~n561 & n564;
  assign n566 = n274 & n553;
  assign n567 = ~n276 & ~n566;
  assign n568 = pi03 & ~n567;
  assign n569 = ~n439 & n486;
  assign n570 = n164 & n569;
  assign n571 = ~n568 & ~n570;
  assign n572 = ~n565 & n571;
  assign n573 = ~pi03 & n519;
  assign n574 = n115 & ~n573;
  assign n575 = n57 & po5;
  assign n576 = ~n42 & ~n532;
  assign n577 = ~n43 & ~n520;
  assign n578 = ~n576 & ~n577;
  assign n579 = ~n575 & ~n578;
  assign n580 = n117 & ~n579;
  assign n581 = ~n574 & ~n580;
  assign n582 = n434 & n581;
  assign n583 = ~n434 & ~n581;
  assign n584 = ~n582 & ~n583;
  assign n585 = n164 & ~n584;
  assign n586 = ~pi02 & n398;
  assign n587 = ~n400 & ~n586;
  assign n588 = pi02 & ~n398;
  assign n589 = ~n587 & ~n588;
  assign n590 = ~n581 & ~n589;
  assign n591 = n581 & n589;
  assign n592 = ~n590 & ~n591;
  assign n593 = pi03 & ~n592;
  assign n594 = n42 & n593;
  assign n595 = ~n557 & ~n594;
  assign n596 = ~n585 & n595;
  assign n597 = ~pi11 & ~n596;
  assign n598 = n572 & ~n597;
  assign n599 = ~n560 & n598;
  assign n600 = n126 & po5;
  assign n601 = n128 & n581;
  assign n602 = ~n600 & ~n601;
  assign n603 = ~n398 & ~n452;
  assign n604 = ~n453 & ~n603;
  assign n605 = n602 & n604;
  assign n606 = ~n602 & ~n604;
  assign n607 = ~n605 & ~n606;
  assign n608 = ~n581 & n607;
  assign n609 = n581 & ~n607;
  assign n610 = n284 & ~n609;
  assign n611 = ~n608 & n610;
  assign n612 = ~pi03 & n439;
  assign n613 = n164 & n612;
  assign n614 = n171 & n556;
  assign n615 = n494 & n614;
  assign n616 = ~n613 & ~n615;
  assign n617 = ~n611 & n616;
  assign n618 = pi11 & ~n617;
  assign n619 = n599 & ~n618;
  assign n620 = ~pi03 & ~n590;
  assign n621 = ~n591 & n620;
  assign n622 = ~pi08 & ~n621;
  assign n623 = ~n417 & ~n421;
  assign n624 = ~n418 & ~n623;
  assign n625 = n520 & n624;
  assign n626 = ~n520 & ~n624;
  assign n627 = ~n625 & ~n626;
  assign n628 = ~n602 & ~n627;
  assign n629 = n602 & n627;
  assign n630 = ~n628 & ~n629;
  assign n631 = pi08 & n630;
  assign n632 = n187 & ~n631;
  assign n633 = ~n622 & n632;
  assign n634 = n619 & ~n633;
  assign n635 = ~n547 & n634;
  assign n636 = ~n546 & n635;
  assign n637 = n481 & ~n636;
  assign n638 = ~n481 & n636;
  assign n639 = pi13 & ~n638;
  assign n640 = ~n637 & n639;
  assign po3 = ~n542 | n640;
  assign po4 = po5 | n494;
  assign n643 = ~po5 & ~n556;
  assign n644 = ~n494 & ~n643;
  assign n645 = n171 & n644;
  assign n646 = ~n532 & n550;
  assign n647 = ~n238 & ~n573;
  assign n648 = ~n646 & n647;
  assign n649 = ~n613 & ~n648;
  assign n650 = ~n645 & n649;
  assign n651 = n581 & ~n606;
  assign n652 = ~n605 & ~n651;
  assign n653 = n284 & n652;
  assign n654 = n650 & ~n653;
  assign n655 = pi11 & ~n654;
  assign n656 = ~pi08 & ~n620;
  assign n657 = ~n591 & n656;
  assign n658 = n602 & ~n626;
  assign n659 = ~n625 & ~n658;
  assign n660 = pi08 & n659;
  assign n661 = ~n657 & ~n660;
  assign n662 = n193 & ~n661;
  assign n663 = pi10 & ~n582;
  assign n664 = n43 & ~n663;
  assign n665 = ~n662 & ~n664;
  assign n666 = ~pi11 & ~n665;
  assign n667 = ~n655 & ~n666;
  assign n668 = pi09 & n25;
  assign n669 = ~n148 & ~n668;
  assign n670 = n543 & ~n669;
  assign n671 = n520 & n670;
  assign n672 = ~n637 & ~n671;
  assign n673 = n667 & n672;
  assign po6 = pi13 & ~n673;
  assign n675 = ~n185 & ~n195;
  assign n676 = ~n463 & po4;
  assign n677 = ~n172 & n676;
  assign po7 = ~n675 & n677;
endmodule
