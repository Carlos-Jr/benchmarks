module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n329, n330, n331, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n475,
    n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489,
    n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n616,
    n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n627, n628, n629, n630, n631,
    n632, n633, n634, n635, n636, n637, n638,
    n639, n640, n641, n642, n643, n644, n645,
    n646, n647, n648, n649, n650, n651, n652,
    n654, n655;
  assign n23 = ~pi08 & ~pi10;
  assign n24 = pi04 & n23;
  assign n25 = pi10 & ~pi11;
  assign n26 = ~pi08 & ~pi09;
  assign n27 = ~pi10 & ~n26;
  assign n28 = pi08 & pi09;
  assign n29 = ~n27 & ~n28;
  assign n30 = ~n25 & n29;
  assign n31 = ~pi09 & n30;
  assign n32 = ~n24 & ~n31;
  assign n33 = pi09 & pi11;
  assign n34 = ~pi10 & ~n33;
  assign n35 = ~pi13 & n34;
  assign n36 = ~pi08 & n35;
  assign n37 = ~pi00 & n36;
  assign n38 = pi00 & pi04;
  assign n39 = ~pi08 & pi10;
  assign n40 = ~pi11 & ~n39;
  assign n41 = n38 & ~n40;
  assign n42 = ~pi09 & ~pi11;
  assign n43 = n39 & n42;
  assign n44 = ~pi09 & n25;
  assign n45 = ~pi09 & pi11;
  assign n46 = n23 & n45;
  assign n47 = ~pi10 & n28;
  assign n48 = pi11 & n47;
  assign n49 = ~n46 & ~n48;
  assign n50 = ~n44 & n49;
  assign n51 = pi13 & ~n50;
  assign n52 = ~n43 & ~n51;
  assign n53 = n41 & ~n52;
  assign n54 = ~pi08 & pi09;
  assign n55 = pi13 & n54;
  assign n56 = ~pi00 & ~n25;
  assign n57 = ~pi00 & ~pi04;
  assign n58 = ~n38 & ~n57;
  assign n59 = ~n56 & n58;
  assign n60 = n55 & n59;
  assign n61 = ~pi10 & ~pi11;
  assign n62 = ~pi13 & ~n61;
  assign n63 = pi08 & ~pi09;
  assign n64 = ~pi10 & pi13;
  assign n65 = n63 & ~n64;
  assign n66 = ~n62 & n65;
  assign n67 = ~n57 & n66;
  assign n68 = ~n25 & n55;
  assign n69 = n25 & n28;
  assign n70 = ~n68 & ~n69;
  assign n71 = pi08 & pi10;
  assign n72 = ~pi13 & n71;
  assign n73 = n45 & n72;
  assign n74 = n70 & ~n73;
  assign n75 = ~pi04 & ~n74;
  assign n76 = ~n67 & ~n75;
  assign n77 = ~n60 & n76;
  assign n78 = ~n53 & n77;
  assign n79 = ~n37 & n78;
  assign n80 = ~n32 & ~n79;
  assign n81 = ~pi08 & n25;
  assign n82 = n57 & n81;
  assign n83 = pi00 & ~n78;
  assign n84 = n71 & n83;
  assign n85 = ~pi08 & pi11;
  assign n86 = pi04 & n85;
  assign n87 = ~n41 & ~n86;
  assign n88 = ~n84 & n87;
  assign n89 = ~n82 & n88;
  assign n90 = pi09 & ~n89;
  assign n91 = pi08 & n61;
  assign n92 = ~n39 & ~n91;
  assign n93 = n79 & ~n92;
  assign n94 = pi08 & n25;
  assign n95 = ~pi04 & n94;
  assign n96 = pi08 & ~pi10;
  assign n97 = ~pi00 & ~n96;
  assign n98 = pi11 & ~n97;
  assign n99 = n58 & n98;
  assign n100 = ~n95 & ~n99;
  assign n101 = ~n93 & n100;
  assign n102 = ~pi09 & ~n101;
  assign n103 = ~n90 & ~n102;
  assign n104 = ~n80 & n103;
  assign n105 = pi00 & pi11;
  assign n106 = ~n27 & n105;
  assign n107 = n104 & ~n106;
  assign n108 = ~pi13 & ~n107;
  assign n109 = ~pi00 & n79;
  assign n110 = ~pi08 & pi13;
  assign n111 = n33 & n110;
  assign n112 = ~n109 & n111;
  assign n113 = pi13 & n25;
  assign n114 = n38 & n63;
  assign n115 = n28 & n83;
  assign n116 = ~n114 & ~n115;
  assign n117 = n26 & n79;
  assign n118 = n116 & ~n117;
  assign n119 = n113 & ~n118;
  assign n120 = ~n112 & ~n119;
  assign n121 = ~pi00 & n43;
  assign n122 = ~pi10 & n111;
  assign n123 = n38 & n122;
  assign n124 = n63 & n113;
  assign n125 = n120 & n124;
  assign n126 = ~n123 & ~n125;
  assign n127 = n23 & n33;
  assign n128 = n126 & n127;
  assign n129 = ~n121 & ~n128;
  assign n130 = ~n120 & ~n129;
  assign n131 = pi11 & ~n27;
  assign n132 = ~pi00 & n131;
  assign n133 = n28 & n132;
  assign n134 = ~pi09 & n96;
  assign n135 = n58 & n134;
  assign n136 = pi08 & n126;
  assign n137 = n44 & n136;
  assign n138 = ~n132 & ~n137;
  assign n139 = ~n79 & ~n138;
  assign n140 = n25 & n54;
  assign n141 = ~n48 & ~n140;
  assign n142 = ~n28 & n105;
  assign n143 = pi08 & ~n126;
  assign n144 = n42 & n143;
  assign n145 = ~n142 & ~n144;
  assign n146 = pi10 & ~n145;
  assign n147 = n141 & ~n146;
  assign n148 = n79 & ~n147;
  assign n149 = pi04 & n96;
  assign n150 = pi00 & ~pi08;
  assign n151 = n120 & n150;
  assign n152 = ~n149 & ~n151;
  assign n153 = n42 & ~n152;
  assign n154 = ~n126 & n127;
  assign n155 = ~n69 & ~n154;
  assign n156 = n120 & ~n155;
  assign n157 = ~n153 & ~n156;
  assign n158 = ~n148 & n157;
  assign n159 = ~n139 & n158;
  assign n160 = pi09 & ~n79;
  assign n161 = ~pi00 & ~n160;
  assign n162 = ~pi09 & n79;
  assign n163 = pi11 & ~n162;
  assign n164 = n23 & ~n163;
  assign n165 = ~n161 & n164;
  assign n166 = n159 & ~n165;
  assign n167 = ~n135 & n166;
  assign n168 = ~n133 & n167;
  assign n169 = ~n130 & n168;
  assign n170 = pi13 & ~n169;
  assign n171 = pi12 & ~n170;
  assign n172 = ~pi12 & n170;
  assign n173 = pi13 & ~n172;
  assign n174 = ~n171 & n173;
  assign n175 = ~pi11 & n28;
  assign n176 = n64 & n175;
  assign n177 = ~pi13 & n39;
  assign n178 = n45 & n177;
  assign n179 = ~n176 & ~n178;
  assign n180 = ~n174 & n179;
  assign po0 = n108 | ~n180;
  assign n182 = pi10 & n28;
  assign n183 = ~pi01 & n36;
  assign n184 = ~pi05 & ~n74;
  assign n185 = pi01 & pi05;
  assign n186 = ~pi00 & n60;
  assign n187 = n52 & ~n186;
  assign n188 = n185 & ~n187;
  assign n189 = ~pi09 & pi10;
  assign n190 = n105 & n189;
  assign n191 = ~pi00 & pi04;
  assign n192 = ~pi01 & ~pi05;
  assign n193 = n191 & ~n192;
  assign n194 = pi09 & ~n193;
  assign n195 = pi01 & ~pi05;
  assign n196 = ~pi01 & pi05;
  assign n197 = ~n191 & ~n196;
  assign n198 = ~n195 & ~n197;
  assign n199 = n25 & n198;
  assign n200 = ~n191 & ~n199;
  assign n201 = ~n195 & n200;
  assign n202 = n194 & ~n201;
  assign n203 = ~n190 & ~n202;
  assign n204 = n110 & ~n203;
  assign n205 = n66 & ~n192;
  assign n206 = ~n204 & ~n205;
  assign n207 = ~n188 & n206;
  assign n208 = ~n184 & n207;
  assign n209 = ~n183 & n208;
  assign n210 = n182 & ~n209;
  assign n211 = ~n131 & ~n210;
  assign n212 = pi01 & ~n211;
  assign n213 = pi05 & n23;
  assign n214 = ~n31 & ~n213;
  assign n215 = ~n209 & ~n214;
  assign n216 = n81 & n192;
  assign n217 = pi01 & ~n40;
  assign n218 = ~n85 & ~n217;
  assign n219 = pi05 & ~n218;
  assign n220 = ~n216 & ~n219;
  assign n221 = pi09 & ~n220;
  assign n222 = ~n92 & n209;
  assign n223 = ~pi05 & n94;
  assign n224 = ~n195 & ~n196;
  assign n225 = ~pi01 & ~n96;
  assign n226 = ~n224 & ~n225;
  assign n227 = pi11 & n226;
  assign n228 = ~n223 & ~n227;
  assign n229 = ~n222 & n228;
  assign n230 = ~pi09 & ~n229;
  assign n231 = ~n221 & ~n230;
  assign n232 = ~n215 & n231;
  assign n233 = ~n212 & n232;
  assign n234 = ~pi13 & ~n233;
  assign n235 = n83 & ~n209;
  assign n236 = ~n83 & n209;
  assign n237 = ~n235 & ~n236;
  assign n238 = pi11 & n29;
  assign n239 = n237 & n238;
  assign n240 = ~pi01 & n209;
  assign n241 = n111 & ~n240;
  assign n242 = ~pi05 & ~pi09;
  assign n243 = pi01 & ~n242;
  assign n244 = pi08 & ~n243;
  assign n245 = pi09 & n209;
  assign n246 = ~pi08 & ~n209;
  assign n247 = n113 & ~n246;
  assign n248 = ~n245 & n247;
  assign n249 = ~n244 & n248;
  assign n250 = ~n241 & ~n249;
  assign n251 = pi00 & ~n120;
  assign n252 = n250 & ~n251;
  assign n253 = ~n120 & ~n250;
  assign n254 = pi00 & n253;
  assign n255 = ~n252 & ~n254;
  assign n256 = n43 & n255;
  assign n257 = ~n239 & ~n256;
  assign n258 = ~pi01 & ~n257;
  assign n259 = n79 & n209;
  assign n260 = ~n141 & n259;
  assign n261 = ~pi08 & ~n255;
  assign n262 = pi01 & n261;
  assign n263 = pi05 & n96;
  assign n264 = ~n79 & ~n126;
  assign n265 = n122 & n185;
  assign n266 = n124 & n250;
  assign n267 = ~n265 & ~n266;
  assign n268 = n264 & ~n267;
  assign n269 = ~n264 & n267;
  assign n270 = ~n268 & ~n269;
  assign n271 = n209 & n270;
  assign n272 = ~n209 & ~n270;
  assign n273 = ~n271 & ~n272;
  assign n274 = n71 & ~n273;
  assign n275 = ~n263 & ~n274;
  assign n276 = ~n262 & n275;
  assign n277 = n42 & ~n276;
  assign n278 = ~pi00 & ~pi01;
  assign n279 = n182 & n278;
  assign n280 = n38 & n192;
  assign n281 = n134 & n280;
  assign n282 = ~n279 & ~n281;
  assign n283 = pi11 & ~n282;
  assign n284 = ~n120 & n123;
  assign n285 = ~n267 & n284;
  assign n286 = n267 & ~n284;
  assign n287 = ~n285 & ~n286;
  assign n288 = n250 & n287;
  assign n289 = ~n250 & ~n287;
  assign n290 = ~n288 & ~n289;
  assign n291 = n127 & ~n290;
  assign n292 = n105 & n182;
  assign n293 = ~pi05 & n134;
  assign n294 = ~n38 & n293;
  assign n295 = n30 & ~n237;
  assign n296 = ~n28 & n61;
  assign n297 = ~n295 & ~n296;
  assign n298 = ~n294 & n297;
  assign n299 = ~n292 & n298;
  assign n300 = pi01 & ~n299;
  assign n301 = n120 & n250;
  assign n302 = ~n253 & ~n301;
  assign n303 = n182 & ~n302;
  assign n304 = pi09 & n23;
  assign n305 = ~n209 & n304;
  assign n306 = ~n303 & ~n305;
  assign n307 = ~pi11 & ~n306;
  assign n308 = ~n38 & ~n196;
  assign n309 = n38 & ~n185;
  assign n310 = n134 & ~n309;
  assign n311 = ~n308 & n310;
  assign n312 = ~pi11 & n304;
  assign n313 = n141 & ~n312;
  assign n314 = ~n79 & ~n313;
  assign n315 = ~n209 & n314;
  assign n316 = ~n311 & ~n315;
  assign n317 = ~n307 & n316;
  assign n318 = ~n300 & n317;
  assign n319 = ~n291 & n318;
  assign n320 = ~n283 & n319;
  assign n321 = ~n277 & n320;
  assign n322 = ~n260 & n321;
  assign n323 = ~n258 & n322;
  assign n324 = n172 & n323;
  assign n325 = n173 & ~n323;
  assign n326 = n179 & ~n325;
  assign n327 = ~n324 & n326;
  assign po1 = n234 | ~n327;
  assign n329 = n172 & ~n323;
  assign n330 = pi02 & pi06;
  assign n331 = ~pi02 & ~pi06;
  assign n332 = pi11 & n331;
  assign n333 = ~n330 & ~n332;
  assign n334 = ~n38 & ~n185;
  assign n335 = ~n192 & ~n334;
  assign n336 = ~n333 & n335;
  assign n337 = ~n330 & ~n331;
  assign n338 = ~n335 & n337;
  assign n339 = ~n336 & ~n338;
  assign n340 = n134 & ~n339;
  assign n341 = ~pi06 & ~n74;
  assign n342 = n66 & ~n331;
  assign n343 = ~pi06 & n198;
  assign n344 = pi06 & ~n199;
  assign n345 = n25 & n344;
  assign n346 = ~n343 & ~n345;
  assign n347 = pi09 & ~n346;
  assign n348 = ~pi02 & n347;
  assign n349 = pi01 & n45;
  assign n350 = pi10 & n349;
  assign n351 = ~n348 & ~n350;
  assign n352 = ~pi06 & ~pi09;
  assign n353 = pi02 & ~n344;
  assign n354 = ~n352 & n353;
  assign n355 = ~n343 & n354;
  assign n356 = n351 & ~n355;
  assign n357 = n110 & ~n356;
  assign n358 = ~n52 & n330;
  assign n359 = ~pi02 & n36;
  assign n360 = ~n358 & ~n359;
  assign n361 = ~n357 & n360;
  assign n362 = ~n342 & n361;
  assign n363 = ~n341 & n362;
  assign n364 = ~pi02 & n363;
  assign n365 = n111 & ~n364;
  assign n366 = n26 & n363;
  assign n367 = pi09 & n363;
  assign n368 = pi02 & ~n367;
  assign n369 = ~n352 & n368;
  assign n370 = pi08 & n369;
  assign n371 = ~n366 & ~n370;
  assign n372 = n113 & ~n371;
  assign n373 = ~n365 & ~n372;
  assign n374 = pi01 & ~n252;
  assign n375 = ~n254 & ~n374;
  assign n376 = n373 & n375;
  assign n377 = ~n373 & ~n375;
  assign n378 = ~n376 & ~n377;
  assign n379 = n43 & n378;
  assign n380 = pi01 & ~n236;
  assign n381 = ~n235 & ~n380;
  assign n382 = n238 & ~n363;
  assign n383 = n381 & n382;
  assign n384 = ~n379 & ~n383;
  assign n385 = ~pi02 & ~n384;
  assign n386 = n122 & n330;
  assign n387 = n124 & n373;
  assign n388 = ~n386 & ~n387;
  assign n389 = ~n286 & ~n288;
  assign n390 = n373 & ~n389;
  assign n391 = ~n373 & n389;
  assign n392 = ~n390 & ~n391;
  assign n393 = n388 & n392;
  assign n394 = ~n388 & ~n392;
  assign n395 = ~n393 & ~n394;
  assign n396 = n127 & ~n395;
  assign n397 = ~pi08 & ~n378;
  assign n398 = pi02 & n397;
  assign n399 = pi06 & n96;
  assign n400 = n363 & n388;
  assign n401 = ~n363 & ~n388;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~n269 & ~n271;
  assign n404 = ~n402 & n403;
  assign n405 = n402 & ~n403;
  assign n406 = ~n404 & ~n405;
  assign n407 = n71 & ~n406;
  assign n408 = ~n399 & ~n407;
  assign n409 = ~n398 & n408;
  assign n410 = n42 & ~n409;
  assign n411 = ~n363 & ~n381;
  assign n412 = n30 & n411;
  assign n413 = ~n296 & ~n412;
  assign n414 = pi02 & ~n413;
  assign n415 = pi02 & pi11;
  assign n416 = ~n278 & n415;
  assign n417 = n301 & n373;
  assign n418 = ~n301 & ~n373;
  assign n419 = ~n417 & ~n418;
  assign n420 = ~pi11 & ~n419;
  assign n421 = ~n416 & ~n420;
  assign n422 = ~pi02 & n278;
  assign n423 = pi11 & n422;
  assign n424 = n421 & ~n423;
  assign n425 = n182 & ~n424;
  assign n426 = n259 & ~n312;
  assign n427 = ~n313 & ~n426;
  assign n428 = ~n363 & n427;
  assign n429 = ~n425 & ~n428;
  assign n430 = ~n414 & n429;
  assign n431 = ~n410 & n430;
  assign n432 = ~n396 & n431;
  assign n433 = ~n385 & n432;
  assign n434 = ~n340 & n433;
  assign n435 = n260 & n363;
  assign n436 = ~pi02 & n381;
  assign n437 = ~pi02 & n238;
  assign n438 = n30 & n381;
  assign n439 = ~n437 & ~n438;
  assign n440 = n363 & ~n439;
  assign n441 = ~n436 & n440;
  assign n442 = ~n435 & ~n441;
  assign n443 = n434 & n442;
  assign n444 = pi13 & ~n443;
  assign n445 = n329 & n444;
  assign n446 = ~n329 & ~n444;
  assign n447 = ~n445 & ~n446;
  assign n448 = n27 & ~n352;
  assign n449 = n415 & ~n448;
  assign n450 = pi09 & n85;
  assign n451 = ~pi02 & n45;
  assign n452 = n96 & n451;
  assign n453 = ~n450 & ~n452;
  assign n454 = pi06 & ~n453;
  assign n455 = ~n92 & n363;
  assign n456 = ~pi06 & n94;
  assign n457 = ~n455 & ~n456;
  assign n458 = ~pi09 & ~n457;
  assign n459 = ~n81 & ~n415;
  assign n460 = ~n337 & ~n459;
  assign n461 = pi09 & n460;
  assign n462 = ~n458 & ~n461;
  assign n463 = ~n454 & n462;
  assign n464 = pi06 & n23;
  assign n465 = pi02 & n182;
  assign n466 = ~n31 & ~n465;
  assign n467 = ~n464 & n466;
  assign n468 = ~n363 & ~n467;
  assign n469 = n463 & ~n468;
  assign n470 = ~n449 & n469;
  assign n471 = ~pi13 & ~n470;
  assign n472 = n179 & ~n471;
  assign po2 = n447 | ~n472;
  assign po5 = pi03 & pi07;
  assign n475 = n51 & po5;
  assign n476 = ~pi03 & ~pi07;
  assign n477 = n66 & ~n476;
  assign n478 = ~pi02 & pi06;
  assign n479 = ~n198 & ~n478;
  assign n480 = pi02 & ~pi06;
  assign n481 = ~n479 & ~n480;
  assign n482 = pi09 & ~n481;
  assign n483 = pi03 & n482;
  assign n484 = n110 & n483;
  assign n485 = n74 & ~n484;
  assign n486 = ~pi07 & ~n485;
  assign n487 = n113 & n481;
  assign n488 = ~n44 & ~n487;
  assign n489 = po5 & ~n488;
  assign n490 = pi07 & n482;
  assign n491 = n113 & n490;
  assign n492 = ~n35 & ~n491;
  assign n493 = ~pi03 & ~n492;
  assign n494 = n189 & n415;
  assign n495 = pi09 & n481;
  assign n496 = n476 & n495;
  assign n497 = ~n494 & ~n496;
  assign n498 = pi13 & ~n497;
  assign n499 = ~n493 & ~n498;
  assign n500 = ~n489 & n499;
  assign n501 = ~pi08 & ~n500;
  assign n502 = ~n486 & ~n501;
  assign n503 = ~n477 & n502;
  assign n504 = ~n475 & n503;
  assign n505 = n259 & n363;
  assign n506 = ~n312 & n505;
  assign n507 = ~n313 & ~n506;
  assign n508 = ~n504 & n507;
  assign n509 = n435 & n504;
  assign n510 = ~n400 & ~n405;
  assign n511 = n122 & po5;
  assign n512 = ~pi03 & n503;
  assign n513 = n111 & ~n512;
  assign n514 = n63 & po5;
  assign n515 = pi03 & ~n504;
  assign n516 = ~n26 & ~n515;
  assign n517 = ~n28 & ~n504;
  assign n518 = ~n516 & ~n517;
  assign n519 = ~n514 & ~n518;
  assign n520 = n113 & ~n519;
  assign n521 = ~n513 & ~n520;
  assign n522 = n124 & n521;
  assign n523 = ~n511 & ~n522;
  assign n524 = n504 & n523;
  assign n525 = ~n504 & ~n523;
  assign n526 = ~n524 & ~n525;
  assign n527 = n510 & ~n526;
  assign n528 = ~n510 & n526;
  assign n529 = ~n527 & ~n528;
  assign n530 = pi08 & ~n529;
  assign n531 = pi02 & ~n376;
  assign n532 = ~n377 & ~n531;
  assign n533 = n521 & n532;
  assign n534 = ~pi08 & ~n533;
  assign n535 = ~n521 & ~n532;
  assign n536 = ~pi03 & ~n535;
  assign n537 = n534 & n536;
  assign n538 = ~n530 & ~n537;
  assign n539 = n44 & ~n538;
  assign n540 = n363 & n381;
  assign n541 = pi02 & ~n540;
  assign n542 = ~n411 & ~n541;
  assign n543 = ~n504 & n542;
  assign n544 = n504 & ~n542;
  assign n545 = ~n543 & ~n544;
  assign n546 = n238 & ~n545;
  assign n547 = ~n331 & ~n338;
  assign n548 = pi07 & n134;
  assign n549 = ~n547 & n548;
  assign n550 = ~n546 & ~n549;
  assign n551 = ~pi03 & ~n550;
  assign n552 = po5 & n547;
  assign n553 = ~po5 & ~n547;
  assign n554 = pi03 & n553;
  assign n555 = ~n552 & ~n554;
  assign n556 = n134 & ~n555;
  assign n557 = n30 & n545;
  assign n558 = ~n296 & ~n557;
  assign n559 = pi03 & ~n558;
  assign n560 = pi03 & pi11;
  assign n561 = ~n422 & n560;
  assign n562 = n182 & n561;
  assign n563 = ~n559 & ~n562;
  assign n564 = ~n556 & n563;
  assign n565 = n417 & n521;
  assign n566 = ~n417 & ~n521;
  assign n567 = ~n565 & ~n566;
  assign n568 = n182 & ~n567;
  assign n569 = ~n533 & ~n535;
  assign n570 = pi03 & ~n569;
  assign n571 = n26 & n570;
  assign n572 = ~n548 & ~n571;
  assign n573 = ~n568 & n572;
  assign n574 = ~pi11 & ~n573;
  assign n575 = n564 & ~n574;
  assign n576 = ~n551 & n575;
  assign n577 = ~pi03 & n422;
  assign n578 = n182 & n577;
  assign n579 = ~n390 & ~n393;
  assign n580 = n521 & ~n579;
  assign n581 = ~n521 & n579;
  assign n582 = ~n580 & ~n581;
  assign n583 = n523 & n582;
  assign n584 = ~n523 & ~n582;
  assign n585 = ~n583 & ~n584;
  assign n586 = n304 & ~n585;
  assign n587 = n134 & n547;
  assign n588 = n476 & n587;
  assign n589 = ~n586 & ~n588;
  assign n590 = ~n578 & n589;
  assign n591 = pi11 & ~n590;
  assign n592 = n576 & ~n591;
  assign n593 = ~n539 & n592;
  assign n594 = ~n509 & n593;
  assign n595 = ~n508 & n594;
  assign n596 = pi13 & ~n595;
  assign n597 = ~n445 & ~n596;
  assign n598 = n445 & ~n595;
  assign n599 = ~n597 & ~n598;
  assign n600 = ~pi07 & ~pi09;
  assign n601 = n27 & ~n600;
  assign n602 = n560 & ~n601;
  assign n603 = pi07 & n23;
  assign n604 = ~n31 & ~n603;
  assign n605 = ~n504 & ~n604;
  assign n606 = ~pi03 & n45;
  assign n607 = n96 & n606;
  assign n608 = ~n450 & ~n607;
  assign n609 = pi07 & ~n608;
  assign n610 = ~n92 & n504;
  assign n611 = ~pi07 & n94;
  assign n612 = ~n610 & ~n611;
  assign n613 = ~pi09 & ~n612;
  assign n614 = n71 & n515;
  assign po4 = po5 | n476;
  assign n616 = ~n81 & ~n560;
  assign n617 = po4 & ~n616;
  assign n618 = ~n614 & ~n617;
  assign n619 = pi09 & ~n618;
  assign n620 = ~n613 & ~n619;
  assign n621 = ~n609 & n620;
  assign n622 = ~n605 & n621;
  assign n623 = ~n602 & n622;
  assign n624 = ~pi13 & ~n623;
  assign n625 = n179 & ~n624;
  assign po3 = n599 | ~n625;
  assign n627 = ~n476 & ~n553;
  assign n628 = n134 & n627;
  assign n629 = ~n512 & ~n542;
  assign n630 = ~n515 & ~n629;
  assign n631 = n29 & ~n630;
  assign n632 = ~n578 & ~n631;
  assign n633 = ~n628 & n632;
  assign n634 = ~n580 & ~n583;
  assign n635 = n304 & n634;
  assign n636 = n633 & ~n635;
  assign n637 = pi11 & ~n636;
  assign n638 = n534 & ~n536;
  assign n639 = ~n524 & ~n528;
  assign n640 = pi08 & n639;
  assign n641 = ~n638 & ~n640;
  assign n642 = n189 & ~n641;
  assign n643 = pi10 & ~n565;
  assign n644 = n28 & ~n643;
  assign n645 = ~n642 & ~n644;
  assign n646 = ~pi11 & ~n645;
  assign n647 = ~n637 & ~n646;
  assign n648 = ~n47 & ~n140;
  assign n649 = n505 & ~n648;
  assign n650 = n504 & n649;
  assign n651 = ~n598 & ~n650;
  assign n652 = n647 & n651;
  assign po6 = pi13 & ~n652;
  assign n654 = ~n337 & po4;
  assign n655 = ~n58 & n654;
  assign po7 = n224 & n655;
endmodule
