module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 ,
    pi5 , pi6 , pi7 , pi8 , pi9 ,
    pi10 , pi11 , pi12 , pi13 , pi14 ,
    pi15 , pi16 , pi17 , pi18 , pi19 ,
    pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 ,
    pi35 , pi36 , pi37 , pi38 , pi39 ,
    pi40 , pi41 , pi42 , pi43 , pi44 ,
    pi45 , pi46 , pi47 , pi48 , pi49 ,
    pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 ,
    po14 , po15 , po16 , po17 ,
    po18 , po19 , po20 , po21 ,
    po22 , po23 , po24 , po25 ,
    po26 , po27 , po28 , po29 ;
  wire n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n136, n137, n138, n139, n140,
    n141, n142, n143, n144, n145, n146, n147,
    n148, n149, n150, n151, n152, n153, n154,
    n155, n156, n157, n158, n159, n160, n161,
    n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183,
    n184, n185, n186, n187, n188, n189, n190,
    n191, n192, n193, n194, n195, n196, n197,
    n198, n199, n200, n201, n202, n203, n204,
    n205, n206, n207, n208, n209, n210, n211,
    n212, n213, n214, n215, n216, n217, n218,
    n219, n220, n221, n222, n223, n224, n225,
    n226, n227, n228, n229, n230, n231, n232,
    n233, n234, n235, n236, n237, n238, n239,
    n240, n241, n242, n243, n244, n245, n246,
    n247, n248, n249, n250, n251, n252, n253,
    n254, n255, n256, n257, n258, n259, n260,
    n261, n262, n263, n265, n266, n267;
  assign n92 = pi27  & pi28 ;
  assign n93 = pi29  & n92;
  assign n94 = ~pi9  & ~pi10 ;
  assign n95 = pi11  & ~n94;
  assign n96 = ~pi12  & ~pi13 ;
  assign n97 = ~n95 & n96;
  assign n98 = pi14  & ~n97;
  assign n99 = pi15  & n98;
  assign n100 = ~pi16  & ~n99;
  assign n101 = pi17  & ~n100;
  assign n102 = ~pi18  & ~n101;
  assign n103 = pi19  & pi20 ;
  assign n104 = ~n102 & n103;
  assign n105 = ~pi21  & ~pi22 ;
  assign n106 = ~n104 & n105;
  assign n107 = pi23  & ~n106;
  assign n108 = pi24  & n107;
  assign n109 = pi25  & n108;
  assign n110 = ~pi26  & ~n109;
  assign n111 = n93 & ~n110;
  assign n112 = pi16  & n99;
  assign n113 = ~pi22  & pi23 ;
  assign n114 = pi20  & ~pi21 ;
  assign n115 = ~pi12  & n95;
  assign n116 = ~pi11  & pi12 ;
  assign n117 = n94 & n116;
  assign n118 = ~n115 & ~n117;
  assign n119 = ~pi15  & ~n98;
  assign n120 = ~n99 & ~n119;
  assign n121 = ~pi1  & ~pi2 ;
  assign n122 = ~pi3  & ~pi4 ;
  assign n123 = ~pi5  & ~pi6 ;
  assign n124 = ~pi7  & ~pi8 ;
  assign n125 = pi9  & ~pi10 ;
  assign n126 = ~pi13  & pi14 ;
  assign n127 = ~pi18  & pi19 ;
  assign n128 = pi24  & pi25 ;
  assign n129 = ~pi26  & n128;
  assign n130 = n126 & n127;
  assign n131 = n124 & n125;
  assign n132 = n122 & n123;
  assign n133 = n113 & n121;
  assign n134 = n114 & n133;
  assign n135 = n131 & n132;
  assign n136 = n129 & n130;
  assign n137 = n135 & n136;
  assign n138 = n134 & n137;
  assign n139 = ~n118 & n138;
  assign n140 = ~n112 & n139;
  assign n141 = ~n120 & n140;
  assign n142 = n101 & n141;
  assign n143 = n111 & ~n142;
  assign n144 = ~pi24  & ~n107;
  assign n145 = ~pi17  & n100;
  assign n146 = ~pi14  & n97;
  assign n147 = pi0  & pi1 ;
  assign n148 = pi2  & pi3 ;
  assign n149 = pi4  & pi5 ;
  assign n150 = pi6  & pi7 ;
  assign n151 = pi8  & pi11 ;
  assign n152 = pi15  & ~pi16 ;
  assign n153 = pi19  & pi25 ;
  assign n154 = ~pi26  & n153;
  assign n155 = n96 & n152;
  assign n156 = n150 & n151;
  assign n157 = n148 & n149;
  assign n158 = n94 & n147;
  assign n159 = n113 & n114;
  assign n160 = n158 & n159;
  assign n161 = n156 & n157;
  assign n162 = n154 & n155;
  assign n163 = n93 & n162;
  assign n164 = n160 & n161;
  assign n165 = n163 & n164;
  assign n166 = ~n98 & ~n146;
  assign n167 = n165 & n166;
  assign n168 = ~n145 & n167;
  assign n169 = n102 & n168;
  assign n170 = ~n108 & n169;
  assign n171 = ~n144 & n170;
  assign n172 = ~n111 & ~n171;
  assign po0  = n143 | n172;
  assign n174 = pi57  & pi58 ;
  assign n175 = pi59  & n174;
  assign n176 = pi54  & pi55 ;
  assign n177 = ~pi39  & ~pi40 ;
  assign n178 = pi41  & ~n177;
  assign n179 = ~pi42  & ~n178;
  assign n180 = ~pi43  & n179;
  assign n181 = pi44  & ~n180;
  assign n182 = pi45  & n181;
  assign n183 = ~pi46  & ~n182;
  assign n184 = pi47  & ~n183;
  assign n185 = ~pi48  & ~n184;
  assign n186 = pi49  & pi50 ;
  assign n187 = ~n185 & n186;
  assign n188 = ~pi51  & ~pi52 ;
  assign n189 = ~n187 & n188;
  assign n190 = pi53  & n176;
  assign n191 = ~n189 & n190;
  assign n192 = ~pi56  & ~n191;
  assign n193 = n175 & ~n192;
  assign n194 = ~pi0  & ~pi51 ;
  assign n195 = ~n193 & ~n194;
  assign n196 = ~pi52  & pi53 ;
  assign n197 = ~n187 & ~n196;
  assign n198 = pi42  & n178;
  assign n199 = pi43  & n198;
  assign n200 = ~pi44  & ~n199;
  assign n201 = ~pi49  & n184;
  assign n202 = ~n185 & ~n201;
  assign n203 = ~pi45  & ~n181;
  assign n204 = ~pi48  & ~pi49 ;
  assign n205 = pi52  & ~pi53 ;
  assign n206 = n187 & ~n205;
  assign n207 = pi30  & pi31 ;
  assign n208 = pi32  & pi33 ;
  assign n209 = pi34  & pi35 ;
  assign n210 = pi36  & pi37 ;
  assign n211 = pi38  & pi41 ;
  assign n212 = ~pi46  & pi47 ;
  assign n213 = pi50  & ~pi56 ;
  assign n214 = n212 & n213;
  assign n215 = n210 & n211;
  assign n216 = n208 & n209;
  assign n217 = n176 & n207;
  assign n218 = n177 & ~n204;
  assign n219 = n217 & n218;
  assign n220 = n215 & n216;
  assign n221 = n175 & n214;
  assign n222 = n220 & n221;
  assign n223 = n219 & n222;
  assign n224 = ~n181 & n223;
  assign n225 = ~n200 & n224;
  assign n226 = ~n182 & ~n203;
  assign n227 = n225 & n226;
  assign n228 = ~n202 & n227;
  assign n229 = ~n197 & n228;
  assign n230 = ~n206 & n229;
  assign n231 = ~n195 & n230;
  assign n232 = pi47  & pi48 ;
  assign n233 = pi48  & n183;
  assign n234 = ~n184 & ~n233;
  assign n235 = ~pi31  & ~pi32 ;
  assign n236 = ~pi33  & ~pi34 ;
  assign n237 = ~pi35  & ~pi36 ;
  assign n238 = ~pi37  & ~pi38 ;
  assign n239 = pi39  & ~pi40 ;
  assign n240 = pi41  & ~pi43 ;
  assign n241 = pi44  & pi45 ;
  assign n242 = ~pi46  & ~pi51 ;
  assign n243 = ~pi56  & pi57 ;
  assign n244 = n242 & n243;
  assign n245 = n240 & n241;
  assign n246 = n238 & n239;
  assign n247 = n236 & n237;
  assign n248 = n176 & n235;
  assign n249 = n186 & n196;
  assign n250 = ~n232 & n249;
  assign n251 = n247 & n248;
  assign n252 = n245 & n246;
  assign n253 = n244 & n252;
  assign n254 = n250 & n251;
  assign n255 = ~n179 & ~n198;
  assign n256 = n254 & n255;
  assign n257 = n253 & n256;
  assign n258 = ~n234 & n257;
  assign n259 = ~pi0  & ~pi30 ;
  assign n260 = n258 & n259;
  assign n261 = n193 & ~n260;
  assign n262 = ~n231 & ~n261;
  assign n263 = ~n172 & ~n262;
  assign po1  = ~n143 & ~n263;
  assign n265 = pi0  & pi30 ;
  assign n266 = n258 & ~n265;
  assign n267 = n193 & ~n266;
  assign po2  = ~po0  & n267;
  assign po3  = 1'b0;
  assign po4  = 1'b0;
  assign po5  = 1'b0;
  assign po6  = 1'b0;
  assign po7  = 1'b0;
  assign po8  = 1'b0;
  assign po9  = 1'b0;
  assign po10  = 1'b0;
  assign po11  = 1'b0;
  assign po12  = 1'b0;
  assign po13  = 1'b0;
  assign po14  = 1'b0;
  assign po15  = 1'b0;
  assign po16  = 1'b0;
  assign po17  = 1'b0;
  assign po18  = 1'b0;
  assign po19  = 1'b0;
  assign po20  = 1'b0;
  assign po21  = 1'b0;
  assign po22  = 1'b0;
  assign po23  = 1'b0;
  assign po24  = 1'b0;
  assign po25  = 1'b0;
  assign po26  = 1'b0;
  assign po27  = 1'b0;
  assign po28  = 1'b0;
  assign po29  = 1'b0;
endmodule
