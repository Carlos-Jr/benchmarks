module mem_ctrl ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17,
    pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26,
    pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34, pi35,
    pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43, pi44,
    pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52, pi53,
    pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61, pi62,
    pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70, pi71,
    pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79, pi80,
    pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107,
    pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116,
    pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124, pi125,
    pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133, pi134,
    pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142, pi143,
    pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151, pi152,
    pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160, pi161,
    pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169, pi170,
    pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178, pi179,
    pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187, pi188,
    pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196, pi197,
    pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205, pi206,
    pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214, pi215,
    pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223, pi224,
    pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232, pi233,
    pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241, pi242,
    pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250, pi251,
    pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259, pi260,
    pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268, pi269,
    pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277, pi278,
    pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286, pi287,
    pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295, pi296,
    pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304, pi305,
    pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313, pi314,
    pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322, pi323,
    pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331, pi332,
    pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340, pi341,
    pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349, pi350,
    pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358, pi359,
    pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367, pi368,
    pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376, pi377,
    pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385, pi386,
    pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394, pi395,
    pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403, pi404,
    pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412, pi413,
    pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421, pi422,
    pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430, pi431,
    pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439, pi440,
    pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448, pi449,
    pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457, pi458,
    pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466, pi467,
    pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475, pi476,
    pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484, pi485,
    pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493, pi494,
    pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502, pi503,
    pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511, pi512,
    pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520, pi521,
    pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529, pi530,
    pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538, pi539,
    pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547, pi548,
    pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556, pi557,
    pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565, pi566,
    pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574, pi575,
    pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583, pi584,
    pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592, pi593,
    pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601, pi602,
    pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610, pi611,
    pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619, pi620,
    pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628, pi629,
    pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637, pi638,
    pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646, pi647,
    pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655, pi656,
    pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664, pi665,
    pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673, pi674,
    pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682, pi683,
    pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691, pi692,
    pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700, pi701,
    pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709, pi710,
    pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718, pi719,
    pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727, pi728,
    pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736, pi737,
    pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745, pi746,
    pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754, pi755,
    pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763, pi764,
    pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772, pi773,
    pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781, pi782,
    pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790, pi791,
    pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799, pi800,
    pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808, pi809,
    pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817, pi818,
    pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826, pi827,
    pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835, pi836,
    pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844, pi845,
    pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853, pi854,
    pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862, pi863,
    pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871, pi872,
    pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880, pi881,
    pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889, pi890,
    pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898, pi899,
    pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907, pi908,
    pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916, pi917,
    pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925, pi926,
    pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934, pi935,
    pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943, pi944,
    pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952, pi953,
    pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961, pi962,
    pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970, pi971,
    pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979, pi980,
    pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988, pi989,
    pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997, pi998,
    pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006, pi1007,
    pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015, pi1016,
    pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024, pi1025,
    pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033, pi1034,
    pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042, pi1043,
    pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051, pi1052,
    pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060, pi1061,
    pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069, pi1070,
    pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078, pi1079,
    pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087, pi1088,
    pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096, pi1097,
    pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105, pi1106,
    pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114, pi1115,
    pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123, pi1124,
    pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132, pi1133,
    pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141, pi1142,
    pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150, pi1151,
    pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159, pi1160,
    pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168, pi1169,
    pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177, pi1178,
    pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186, pi1187,
    pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195, pi1196,
    pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203,
    po0, po1, po2, po3, po4, po5, po6, po7, po8,
    po9, po10, po11, po12, po13, po14, po15, po16, po17,
    po18, po19, po20, po21, po22, po23, po24, po25, po26,
    po27, po28, po29, po30, po31, po32, po33, po34, po35,
    po36, po37, po38, po39, po40, po41, po42, po43, po44,
    po45, po46, po47, po48, po49, po50, po51, po52, po53,
    po54, po55, po56, po57, po58, po59, po60, po61, po62,
    po63, po64, po65, po66, po67, po68, po69, po70, po71,
    po72, po73, po74, po75, po76, po77, po78, po79, po80,
    po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98,
    po99, po100, po101, po102, po103, po104, po105, po106, po107,
    po108, po109, po110, po111, po112, po113, po114, po115, po116,
    po117, po118, po119, po120, po121, po122, po123, po124, po125,
    po126, po127, po128, po129, po130, po131, po132, po133, po134,
    po135, po136, po137, po138, po139, po140, po141, po142, po143,
    po144, po145, po146, po147, po148, po149, po150, po151, po152,
    po153, po154, po155, po156, po157, po158, po159, po160, po161,
    po162, po163, po164, po165, po166, po167, po168, po169, po170,
    po171, po172, po173, po174, po175, po176, po177, po178, po179,
    po180, po181, po182, po183, po184, po185, po186, po187, po188,
    po189, po190, po191, po192, po193, po194, po195, po196, po197,
    po198, po199, po200, po201, po202, po203, po204, po205, po206,
    po207, po208, po209, po210, po211, po212, po213, po214, po215,
    po216, po217, po218, po219, po220, po221, po222, po223, po224,
    po225, po226, po227, po228, po229, po230, po231, po232, po233,
    po234, po235, po236, po237, po238, po239, po240, po241, po242,
    po243, po244, po245, po246, po247, po248, po249, po250, po251,
    po252, po253, po254, po255, po256, po257, po258, po259, po260,
    po261, po262, po263, po264, po265, po266, po267, po268, po269,
    po270, po271, po272, po273, po274, po275, po276, po277, po278,
    po279, po280, po281, po282, po283, po284, po285, po286, po287,
    po288, po289, po290, po291, po292, po293, po294, po295, po296,
    po297, po298, po299, po300, po301, po302, po303, po304, po305,
    po306, po307, po308, po309, po310, po311, po312, po313, po314,
    po315, po316, po317, po318, po319, po320, po321, po322, po323,
    po324, po325, po326, po327, po328, po329, po330, po331, po332,
    po333, po334, po335, po336, po337, po338, po339, po340, po341,
    po342, po343, po344, po345, po346, po347, po348, po349, po350,
    po351, po352, po353, po354, po355, po356, po357, po358, po359,
    po360, po361, po362, po363, po364, po365, po366, po367, po368,
    po369, po370, po371, po372, po373, po374, po375, po376, po377,
    po378, po379, po380, po381, po382, po383, po384, po385, po386,
    po387, po388, po389, po390, po391, po392, po393, po394, po395,
    po396, po397, po398, po399, po400, po401, po402, po403, po404,
    po405, po406, po407, po408, po409, po410, po411, po412, po413,
    po414, po415, po416, po417, po418, po419, po420, po421, po422,
    po423, po424, po425, po426, po427, po428, po429, po430, po431,
    po432, po433, po434, po435, po436, po437, po438, po439, po440,
    po441, po442, po443, po444, po445, po446, po447, po448, po449,
    po450, po451, po452, po453, po454, po455, po456, po457, po458,
    po459, po460, po461, po462, po463, po464, po465, po466, po467,
    po468, po469, po470, po471, po472, po473, po474, po475, po476,
    po477, po478, po479, po480, po481, po482, po483, po484, po485,
    po486, po487, po488, po489, po490, po491, po492, po493, po494,
    po495, po496, po497, po498, po499, po500, po501, po502, po503,
    po504, po505, po506, po507, po508, po509, po510, po511, po512,
    po513, po514, po515, po516, po517, po518, po519, po520, po521,
    po522, po523, po524, po525, po526, po527, po528, po529, po530,
    po531, po532, po533, po534, po535, po536, po537, po538, po539,
    po540, po541, po542, po543, po544, po545, po546, po547, po548,
    po549, po550, po551, po552, po553, po554, po555, po556, po557,
    po558, po559, po560, po561, po562, po563, po564, po565, po566,
    po567, po568, po569, po570, po571, po572, po573, po574, po575,
    po576, po577, po578, po579, po580, po581, po582, po583, po584,
    po585, po586, po587, po588, po589, po590, po591, po592, po593,
    po594, po595, po596, po597, po598, po599, po600, po601, po602,
    po603, po604, po605, po606, po607, po608, po609, po610, po611,
    po612, po613, po614, po615, po616, po617, po618, po619, po620,
    po621, po622, po623, po624, po625, po626, po627, po628, po629,
    po630, po631, po632, po633, po634, po635, po636, po637, po638,
    po639, po640, po641, po642, po643, po644, po645, po646, po647,
    po648, po649, po650, po651, po652, po653, po654, po655, po656,
    po657, po658, po659, po660, po661, po662, po663, po664, po665,
    po666, po667, po668, po669, po670, po671, po672, po673, po674,
    po675, po676, po677, po678, po679, po680, po681, po682, po683,
    po684, po685, po686, po687, po688, po689, po690, po691, po692,
    po693, po694, po695, po696, po697, po698, po699, po700, po701,
    po702, po703, po704, po705, po706, po707, po708, po709, po710,
    po711, po712, po713, po714, po715, po716, po717, po718, po719,
    po720, po721, po722, po723, po724, po725, po726, po727, po728,
    po729, po730, po731, po732, po733, po734, po735, po736, po737,
    po738, po739, po740, po741, po742, po743, po744, po745, po746,
    po747, po748, po749, po750, po751, po752, po753, po754, po755,
    po756, po757, po758, po759, po760, po761, po762, po763, po764,
    po765, po766, po767, po768, po769, po770, po771, po772, po773,
    po774, po775, po776, po777, po778, po779, po780, po781, po782,
    po783, po784, po785, po786, po787, po788, po789, po790, po791,
    po792, po793, po794, po795, po796, po797, po798, po799, po800,
    po801, po802, po803, po804, po805, po806, po807, po808, po809,
    po810, po811, po812, po813, po814, po815, po816, po817, po818,
    po819, po820, po821, po822, po823, po824, po825, po826, po827,
    po828, po829, po830, po831, po832, po833, po834, po835, po836,
    po837, po838, po839, po840, po841, po842, po843, po844, po845,
    po846, po847, po848, po849, po850, po851, po852, po853, po854,
    po855, po856, po857, po858, po859, po860, po861, po862, po863,
    po864, po865, po866, po867, po868, po869, po870, po871, po872,
    po873, po874, po875, po876, po877, po878, po879, po880, po881,
    po882, po883, po884, po885, po886, po887, po888, po889, po890,
    po891, po892, po893, po894, po895, po896, po897, po898, po899,
    po900, po901, po902, po903, po904, po905, po906, po907, po908,
    po909, po910, po911, po912, po913, po914, po915, po916, po917,
    po918, po919, po920, po921, po922, po923, po924, po925, po926,
    po927, po928, po929, po930, po931, po932, po933, po934, po935,
    po936, po937, po938, po939, po940, po941, po942, po943, po944,
    po945, po946, po947, po948, po949, po950, po951, po952, po953,
    po954, po955, po956, po957, po958, po959, po960, po961, po962,
    po963, po964, po965, po966, po967, po968, po969, po970, po971,
    po972, po973, po974, po975, po976, po977, po978, po979, po980,
    po981, po982, po983, po984, po985, po986, po987, po988, po989,
    po990, po991, po992, po993, po994, po995, po996, po997, po998,
    po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006, po1007,
    po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015, po1016,
    po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024, po1025,
    po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033, po1034,
    po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042, po1043,
    po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051, po1052,
    po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060, po1061,
    po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069, po1070,
    po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078, po1079,
    po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087, po1088,
    po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096, po1097,
    po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105, po1106,
    po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114, po1115,
    po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123, po1124,
    po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132, po1133,
    po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141, po1142,
    po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150, po1151,
    po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159, po1160,
    po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168, po1169,
    po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177, po1178,
    po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186, po1187,
    po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195, po1196,
    po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204, po1205,
    po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213, po1214,
    po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222, po1223,
    po1224, po1225, po1226, po1227, po1228, po1229, po1230  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7,
    pi8, pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16,
    pi17, pi18, pi19, pi20, pi21, pi22, pi23, pi24, pi25,
    pi26, pi27, pi28, pi29, pi30, pi31, pi32, pi33, pi34,
    pi35, pi36, pi37, pi38, pi39, pi40, pi41, pi42, pi43,
    pi44, pi45, pi46, pi47, pi48, pi49, pi50, pi51, pi52,
    pi53, pi54, pi55, pi56, pi57, pi58, pi59, pi60, pi61,
    pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69, pi70,
    pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97,
    pi98, pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106,
    pi107, pi108, pi109, pi110, pi111, pi112, pi113, pi114, pi115,
    pi116, pi117, pi118, pi119, pi120, pi121, pi122, pi123, pi124,
    pi125, pi126, pi127, pi128, pi129, pi130, pi131, pi132, pi133,
    pi134, pi135, pi136, pi137, pi138, pi139, pi140, pi141, pi142,
    pi143, pi144, pi145, pi146, pi147, pi148, pi149, pi150, pi151,
    pi152, pi153, pi154, pi155, pi156, pi157, pi158, pi159, pi160,
    pi161, pi162, pi163, pi164, pi165, pi166, pi167, pi168, pi169,
    pi170, pi171, pi172, pi173, pi174, pi175, pi176, pi177, pi178,
    pi179, pi180, pi181, pi182, pi183, pi184, pi185, pi186, pi187,
    pi188, pi189, pi190, pi191, pi192, pi193, pi194, pi195, pi196,
    pi197, pi198, pi199, pi200, pi201, pi202, pi203, pi204, pi205,
    pi206, pi207, pi208, pi209, pi210, pi211, pi212, pi213, pi214,
    pi215, pi216, pi217, pi218, pi219, pi220, pi221, pi222, pi223,
    pi224, pi225, pi226, pi227, pi228, pi229, pi230, pi231, pi232,
    pi233, pi234, pi235, pi236, pi237, pi238, pi239, pi240, pi241,
    pi242, pi243, pi244, pi245, pi246, pi247, pi248, pi249, pi250,
    pi251, pi252, pi253, pi254, pi255, pi256, pi257, pi258, pi259,
    pi260, pi261, pi262, pi263, pi264, pi265, pi266, pi267, pi268,
    pi269, pi270, pi271, pi272, pi273, pi274, pi275, pi276, pi277,
    pi278, pi279, pi280, pi281, pi282, pi283, pi284, pi285, pi286,
    pi287, pi288, pi289, pi290, pi291, pi292, pi293, pi294, pi295,
    pi296, pi297, pi298, pi299, pi300, pi301, pi302, pi303, pi304,
    pi305, pi306, pi307, pi308, pi309, pi310, pi311, pi312, pi313,
    pi314, pi315, pi316, pi317, pi318, pi319, pi320, pi321, pi322,
    pi323, pi324, pi325, pi326, pi327, pi328, pi329, pi330, pi331,
    pi332, pi333, pi334, pi335, pi336, pi337, pi338, pi339, pi340,
    pi341, pi342, pi343, pi344, pi345, pi346, pi347, pi348, pi349,
    pi350, pi351, pi352, pi353, pi354, pi355, pi356, pi357, pi358,
    pi359, pi360, pi361, pi362, pi363, pi364, pi365, pi366, pi367,
    pi368, pi369, pi370, pi371, pi372, pi373, pi374, pi375, pi376,
    pi377, pi378, pi379, pi380, pi381, pi382, pi383, pi384, pi385,
    pi386, pi387, pi388, pi389, pi390, pi391, pi392, pi393, pi394,
    pi395, pi396, pi397, pi398, pi399, pi400, pi401, pi402, pi403,
    pi404, pi405, pi406, pi407, pi408, pi409, pi410, pi411, pi412,
    pi413, pi414, pi415, pi416, pi417, pi418, pi419, pi420, pi421,
    pi422, pi423, pi424, pi425, pi426, pi427, pi428, pi429, pi430,
    pi431, pi432, pi433, pi434, pi435, pi436, pi437, pi438, pi439,
    pi440, pi441, pi442, pi443, pi444, pi445, pi446, pi447, pi448,
    pi449, pi450, pi451, pi452, pi453, pi454, pi455, pi456, pi457,
    pi458, pi459, pi460, pi461, pi462, pi463, pi464, pi465, pi466,
    pi467, pi468, pi469, pi470, pi471, pi472, pi473, pi474, pi475,
    pi476, pi477, pi478, pi479, pi480, pi481, pi482, pi483, pi484,
    pi485, pi486, pi487, pi488, pi489, pi490, pi491, pi492, pi493,
    pi494, pi495, pi496, pi497, pi498, pi499, pi500, pi501, pi502,
    pi503, pi504, pi505, pi506, pi507, pi508, pi509, pi510, pi511,
    pi512, pi513, pi514, pi515, pi516, pi517, pi518, pi519, pi520,
    pi521, pi522, pi523, pi524, pi525, pi526, pi527, pi528, pi529,
    pi530, pi531, pi532, pi533, pi534, pi535, pi536, pi537, pi538,
    pi539, pi540, pi541, pi542, pi543, pi544, pi545, pi546, pi547,
    pi548, pi549, pi550, pi551, pi552, pi553, pi554, pi555, pi556,
    pi557, pi558, pi559, pi560, pi561, pi562, pi563, pi564, pi565,
    pi566, pi567, pi568, pi569, pi570, pi571, pi572, pi573, pi574,
    pi575, pi576, pi577, pi578, pi579, pi580, pi581, pi582, pi583,
    pi584, pi585, pi586, pi587, pi588, pi589, pi590, pi591, pi592,
    pi593, pi594, pi595, pi596, pi597, pi598, pi599, pi600, pi601,
    pi602, pi603, pi604, pi605, pi606, pi607, pi608, pi609, pi610,
    pi611, pi612, pi613, pi614, pi615, pi616, pi617, pi618, pi619,
    pi620, pi621, pi622, pi623, pi624, pi625, pi626, pi627, pi628,
    pi629, pi630, pi631, pi632, pi633, pi634, pi635, pi636, pi637,
    pi638, pi639, pi640, pi641, pi642, pi643, pi644, pi645, pi646,
    pi647, pi648, pi649, pi650, pi651, pi652, pi653, pi654, pi655,
    pi656, pi657, pi658, pi659, pi660, pi661, pi662, pi663, pi664,
    pi665, pi666, pi667, pi668, pi669, pi670, pi671, pi672, pi673,
    pi674, pi675, pi676, pi677, pi678, pi679, pi680, pi681, pi682,
    pi683, pi684, pi685, pi686, pi687, pi688, pi689, pi690, pi691,
    pi692, pi693, pi694, pi695, pi696, pi697, pi698, pi699, pi700,
    pi701, pi702, pi703, pi704, pi705, pi706, pi707, pi708, pi709,
    pi710, pi711, pi712, pi713, pi714, pi715, pi716, pi717, pi718,
    pi719, pi720, pi721, pi722, pi723, pi724, pi725, pi726, pi727,
    pi728, pi729, pi730, pi731, pi732, pi733, pi734, pi735, pi736,
    pi737, pi738, pi739, pi740, pi741, pi742, pi743, pi744, pi745,
    pi746, pi747, pi748, pi749, pi750, pi751, pi752, pi753, pi754,
    pi755, pi756, pi757, pi758, pi759, pi760, pi761, pi762, pi763,
    pi764, pi765, pi766, pi767, pi768, pi769, pi770, pi771, pi772,
    pi773, pi774, pi775, pi776, pi777, pi778, pi779, pi780, pi781,
    pi782, pi783, pi784, pi785, pi786, pi787, pi788, pi789, pi790,
    pi791, pi792, pi793, pi794, pi795, pi796, pi797, pi798, pi799,
    pi800, pi801, pi802, pi803, pi804, pi805, pi806, pi807, pi808,
    pi809, pi810, pi811, pi812, pi813, pi814, pi815, pi816, pi817,
    pi818, pi819, pi820, pi821, pi822, pi823, pi824, pi825, pi826,
    pi827, pi828, pi829, pi830, pi831, pi832, pi833, pi834, pi835,
    pi836, pi837, pi838, pi839, pi840, pi841, pi842, pi843, pi844,
    pi845, pi846, pi847, pi848, pi849, pi850, pi851, pi852, pi853,
    pi854, pi855, pi856, pi857, pi858, pi859, pi860, pi861, pi862,
    pi863, pi864, pi865, pi866, pi867, pi868, pi869, pi870, pi871,
    pi872, pi873, pi874, pi875, pi876, pi877, pi878, pi879, pi880,
    pi881, pi882, pi883, pi884, pi885, pi886, pi887, pi888, pi889,
    pi890, pi891, pi892, pi893, pi894, pi895, pi896, pi897, pi898,
    pi899, pi900, pi901, pi902, pi903, pi904, pi905, pi906, pi907,
    pi908, pi909, pi910, pi911, pi912, pi913, pi914, pi915, pi916,
    pi917, pi918, pi919, pi920, pi921, pi922, pi923, pi924, pi925,
    pi926, pi927, pi928, pi929, pi930, pi931, pi932, pi933, pi934,
    pi935, pi936, pi937, pi938, pi939, pi940, pi941, pi942, pi943,
    pi944, pi945, pi946, pi947, pi948, pi949, pi950, pi951, pi952,
    pi953, pi954, pi955, pi956, pi957, pi958, pi959, pi960, pi961,
    pi962, pi963, pi964, pi965, pi966, pi967, pi968, pi969, pi970,
    pi971, pi972, pi973, pi974, pi975, pi976, pi977, pi978, pi979,
    pi980, pi981, pi982, pi983, pi984, pi985, pi986, pi987, pi988,
    pi989, pi990, pi991, pi992, pi993, pi994, pi995, pi996, pi997,
    pi998, pi999, pi1000, pi1001, pi1002, pi1003, pi1004, pi1005, pi1006,
    pi1007, pi1008, pi1009, pi1010, pi1011, pi1012, pi1013, pi1014, pi1015,
    pi1016, pi1017, pi1018, pi1019, pi1020, pi1021, pi1022, pi1023, pi1024,
    pi1025, pi1026, pi1027, pi1028, pi1029, pi1030, pi1031, pi1032, pi1033,
    pi1034, pi1035, pi1036, pi1037, pi1038, pi1039, pi1040, pi1041, pi1042,
    pi1043, pi1044, pi1045, pi1046, pi1047, pi1048, pi1049, pi1050, pi1051,
    pi1052, pi1053, pi1054, pi1055, pi1056, pi1057, pi1058, pi1059, pi1060,
    pi1061, pi1062, pi1063, pi1064, pi1065, pi1066, pi1067, pi1068, pi1069,
    pi1070, pi1071, pi1072, pi1073, pi1074, pi1075, pi1076, pi1077, pi1078,
    pi1079, pi1080, pi1081, pi1082, pi1083, pi1084, pi1085, pi1086, pi1087,
    pi1088, pi1089, pi1090, pi1091, pi1092, pi1093, pi1094, pi1095, pi1096,
    pi1097, pi1098, pi1099, pi1100, pi1101, pi1102, pi1103, pi1104, pi1105,
    pi1106, pi1107, pi1108, pi1109, pi1110, pi1111, pi1112, pi1113, pi1114,
    pi1115, pi1116, pi1117, pi1118, pi1119, pi1120, pi1121, pi1122, pi1123,
    pi1124, pi1125, pi1126, pi1127, pi1128, pi1129, pi1130, pi1131, pi1132,
    pi1133, pi1134, pi1135, pi1136, pi1137, pi1138, pi1139, pi1140, pi1141,
    pi1142, pi1143, pi1144, pi1145, pi1146, pi1147, pi1148, pi1149, pi1150,
    pi1151, pi1152, pi1153, pi1154, pi1155, pi1156, pi1157, pi1158, pi1159,
    pi1160, pi1161, pi1162, pi1163, pi1164, pi1165, pi1166, pi1167, pi1168,
    pi1169, pi1170, pi1171, pi1172, pi1173, pi1174, pi1175, pi1176, pi1177,
    pi1178, pi1179, pi1180, pi1181, pi1182, pi1183, pi1184, pi1185, pi1186,
    pi1187, pi1188, pi1189, pi1190, pi1191, pi1192, pi1193, pi1194, pi1195,
    pi1196, pi1197, pi1198, pi1199, pi1200, pi1201, pi1202, pi1203;
  output po0, po1, po2, po3, po4, po5, po6, po7,
    po8, po9, po10, po11, po12, po13, po14, po15, po16,
    po17, po18, po19, po20, po21, po22, po23, po24, po25,
    po26, po27, po28, po29, po30, po31, po32, po33, po34,
    po35, po36, po37, po38, po39, po40, po41, po42, po43,
    po44, po45, po46, po47, po48, po49, po50, po51, po52,
    po53, po54, po55, po56, po57, po58, po59, po60, po61,
    po62, po63, po64, po65, po66, po67, po68, po69, po70,
    po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88,
    po89, po90, po91, po92, po93, po94, po95, po96, po97,
    po98, po99, po100, po101, po102, po103, po104, po105, po106,
    po107, po108, po109, po110, po111, po112, po113, po114, po115,
    po116, po117, po118, po119, po120, po121, po122, po123, po124,
    po125, po126, po127, po128, po129, po130, po131, po132, po133,
    po134, po135, po136, po137, po138, po139, po140, po141, po142,
    po143, po144, po145, po146, po147, po148, po149, po150, po151,
    po152, po153, po154, po155, po156, po157, po158, po159, po160,
    po161, po162, po163, po164, po165, po166, po167, po168, po169,
    po170, po171, po172, po173, po174, po175, po176, po177, po178,
    po179, po180, po181, po182, po183, po184, po185, po186, po187,
    po188, po189, po190, po191, po192, po193, po194, po195, po196,
    po197, po198, po199, po200, po201, po202, po203, po204, po205,
    po206, po207, po208, po209, po210, po211, po212, po213, po214,
    po215, po216, po217, po218, po219, po220, po221, po222, po223,
    po224, po225, po226, po227, po228, po229, po230, po231, po232,
    po233, po234, po235, po236, po237, po238, po239, po240, po241,
    po242, po243, po244, po245, po246, po247, po248, po249, po250,
    po251, po252, po253, po254, po255, po256, po257, po258, po259,
    po260, po261, po262, po263, po264, po265, po266, po267, po268,
    po269, po270, po271, po272, po273, po274, po275, po276, po277,
    po278, po279, po280, po281, po282, po283, po284, po285, po286,
    po287, po288, po289, po290, po291, po292, po293, po294, po295,
    po296, po297, po298, po299, po300, po301, po302, po303, po304,
    po305, po306, po307, po308, po309, po310, po311, po312, po313,
    po314, po315, po316, po317, po318, po319, po320, po321, po322,
    po323, po324, po325, po326, po327, po328, po329, po330, po331,
    po332, po333, po334, po335, po336, po337, po338, po339, po340,
    po341, po342, po343, po344, po345, po346, po347, po348, po349,
    po350, po351, po352, po353, po354, po355, po356, po357, po358,
    po359, po360, po361, po362, po363, po364, po365, po366, po367,
    po368, po369, po370, po371, po372, po373, po374, po375, po376,
    po377, po378, po379, po380, po381, po382, po383, po384, po385,
    po386, po387, po388, po389, po390, po391, po392, po393, po394,
    po395, po396, po397, po398, po399, po400, po401, po402, po403,
    po404, po405, po406, po407, po408, po409, po410, po411, po412,
    po413, po414, po415, po416, po417, po418, po419, po420, po421,
    po422, po423, po424, po425, po426, po427, po428, po429, po430,
    po431, po432, po433, po434, po435, po436, po437, po438, po439,
    po440, po441, po442, po443, po444, po445, po446, po447, po448,
    po449, po450, po451, po452, po453, po454, po455, po456, po457,
    po458, po459, po460, po461, po462, po463, po464, po465, po466,
    po467, po468, po469, po470, po471, po472, po473, po474, po475,
    po476, po477, po478, po479, po480, po481, po482, po483, po484,
    po485, po486, po487, po488, po489, po490, po491, po492, po493,
    po494, po495, po496, po497, po498, po499, po500, po501, po502,
    po503, po504, po505, po506, po507, po508, po509, po510, po511,
    po512, po513, po514, po515, po516, po517, po518, po519, po520,
    po521, po522, po523, po524, po525, po526, po527, po528, po529,
    po530, po531, po532, po533, po534, po535, po536, po537, po538,
    po539, po540, po541, po542, po543, po544, po545, po546, po547,
    po548, po549, po550, po551, po552, po553, po554, po555, po556,
    po557, po558, po559, po560, po561, po562, po563, po564, po565,
    po566, po567, po568, po569, po570, po571, po572, po573, po574,
    po575, po576, po577, po578, po579, po580, po581, po582, po583,
    po584, po585, po586, po587, po588, po589, po590, po591, po592,
    po593, po594, po595, po596, po597, po598, po599, po600, po601,
    po602, po603, po604, po605, po606, po607, po608, po609, po610,
    po611, po612, po613, po614, po615, po616, po617, po618, po619,
    po620, po621, po622, po623, po624, po625, po626, po627, po628,
    po629, po630, po631, po632, po633, po634, po635, po636, po637,
    po638, po639, po640, po641, po642, po643, po644, po645, po646,
    po647, po648, po649, po650, po651, po652, po653, po654, po655,
    po656, po657, po658, po659, po660, po661, po662, po663, po664,
    po665, po666, po667, po668, po669, po670, po671, po672, po673,
    po674, po675, po676, po677, po678, po679, po680, po681, po682,
    po683, po684, po685, po686, po687, po688, po689, po690, po691,
    po692, po693, po694, po695, po696, po697, po698, po699, po700,
    po701, po702, po703, po704, po705, po706, po707, po708, po709,
    po710, po711, po712, po713, po714, po715, po716, po717, po718,
    po719, po720, po721, po722, po723, po724, po725, po726, po727,
    po728, po729, po730, po731, po732, po733, po734, po735, po736,
    po737, po738, po739, po740, po741, po742, po743, po744, po745,
    po746, po747, po748, po749, po750, po751, po752, po753, po754,
    po755, po756, po757, po758, po759, po760, po761, po762, po763,
    po764, po765, po766, po767, po768, po769, po770, po771, po772,
    po773, po774, po775, po776, po777, po778, po779, po780, po781,
    po782, po783, po784, po785, po786, po787, po788, po789, po790,
    po791, po792, po793, po794, po795, po796, po797, po798, po799,
    po800, po801, po802, po803, po804, po805, po806, po807, po808,
    po809, po810, po811, po812, po813, po814, po815, po816, po817,
    po818, po819, po820, po821, po822, po823, po824, po825, po826,
    po827, po828, po829, po830, po831, po832, po833, po834, po835,
    po836, po837, po838, po839, po840, po841, po842, po843, po844,
    po845, po846, po847, po848, po849, po850, po851, po852, po853,
    po854, po855, po856, po857, po858, po859, po860, po861, po862,
    po863, po864, po865, po866, po867, po868, po869, po870, po871,
    po872, po873, po874, po875, po876, po877, po878, po879, po880,
    po881, po882, po883, po884, po885, po886, po887, po888, po889,
    po890, po891, po892, po893, po894, po895, po896, po897, po898,
    po899, po900, po901, po902, po903, po904, po905, po906, po907,
    po908, po909, po910, po911, po912, po913, po914, po915, po916,
    po917, po918, po919, po920, po921, po922, po923, po924, po925,
    po926, po927, po928, po929, po930, po931, po932, po933, po934,
    po935, po936, po937, po938, po939, po940, po941, po942, po943,
    po944, po945, po946, po947, po948, po949, po950, po951, po952,
    po953, po954, po955, po956, po957, po958, po959, po960, po961,
    po962, po963, po964, po965, po966, po967, po968, po969, po970,
    po971, po972, po973, po974, po975, po976, po977, po978, po979,
    po980, po981, po982, po983, po984, po985, po986, po987, po988,
    po989, po990, po991, po992, po993, po994, po995, po996, po997,
    po998, po999, po1000, po1001, po1002, po1003, po1004, po1005, po1006,
    po1007, po1008, po1009, po1010, po1011, po1012, po1013, po1014, po1015,
    po1016, po1017, po1018, po1019, po1020, po1021, po1022, po1023, po1024,
    po1025, po1026, po1027, po1028, po1029, po1030, po1031, po1032, po1033,
    po1034, po1035, po1036, po1037, po1038, po1039, po1040, po1041, po1042,
    po1043, po1044, po1045, po1046, po1047, po1048, po1049, po1050, po1051,
    po1052, po1053, po1054, po1055, po1056, po1057, po1058, po1059, po1060,
    po1061, po1062, po1063, po1064, po1065, po1066, po1067, po1068, po1069,
    po1070, po1071, po1072, po1073, po1074, po1075, po1076, po1077, po1078,
    po1079, po1080, po1081, po1082, po1083, po1084, po1085, po1086, po1087,
    po1088, po1089, po1090, po1091, po1092, po1093, po1094, po1095, po1096,
    po1097, po1098, po1099, po1100, po1101, po1102, po1103, po1104, po1105,
    po1106, po1107, po1108, po1109, po1110, po1111, po1112, po1113, po1114,
    po1115, po1116, po1117, po1118, po1119, po1120, po1121, po1122, po1123,
    po1124, po1125, po1126, po1127, po1128, po1129, po1130, po1131, po1132,
    po1133, po1134, po1135, po1136, po1137, po1138, po1139, po1140, po1141,
    po1142, po1143, po1144, po1145, po1146, po1147, po1148, po1149, po1150,
    po1151, po1152, po1153, po1154, po1155, po1156, po1157, po1158, po1159,
    po1160, po1161, po1162, po1163, po1164, po1165, po1166, po1167, po1168,
    po1169, po1170, po1171, po1172, po1173, po1174, po1175, po1176, po1177,
    po1178, po1179, po1180, po1181, po1182, po1183, po1184, po1185, po1186,
    po1187, po1188, po1189, po1190, po1191, po1192, po1193, po1194, po1195,
    po1196, po1197, po1198, po1199, po1200, po1201, po1202, po1203, po1204,
    po1205, po1206, po1207, po1208, po1209, po1210, po1211, po1212, po1213,
    po1214, po1215, po1216, po1217, po1218, po1219, po1220, po1221, po1222,
    po1223, po1224, po1225, po1226, po1227, po1228, po1229, po1230;
  wire n2437, n2438, n2439, n2440, n2441, n2442,
    n2443, n2444, n2445, n2446, n2447, n2448,
    n2449, n2450, n2451, n2452, n2453, n2454,
    n2455, n2456, n2457, n2458, n2459, n2460,
    n2461, n2462, n2463, n2464, n2465, n2466,
    n2467, n2468, n2469, n2470, n2471, n2472,
    n2473, n2474, n2475, n2476, n2477, n2478,
    n2479, n2480, n2481, n2482, n2483, n2484,
    n2485, n2486, n2487, n2488, n2489, n2490,
    n2491, n2492, n2493, n2494, n2495, n2496,
    n2497, n2498, n2499, n2500, n2501, n2502,
    n2503, n2504, n2505, n2506, n2507, n2508,
    n2509, n2510, n2511, n2512, n2513, n2514,
    n2515, n2516, n2517, n2518, n2519, n2520,
    n2521, n2522, n2523, n2524, n2525, n2526,
    n2527, n2528, n2529, n2530, n2531, n2532,
    n2533, n2534, n2535, n2536, n2537, n2538,
    n2539, n2540, n2541, n2542, n2543, n2544,
    n2545, n2546, n2547, n2548, n2549, n2550,
    n2551, n2552, n2553, n2554, n2555, n2556,
    n2557, n2558, n2559, n2560, n2561, n2562,
    n2563, n2564, n2565, n2566, n2567, n2568,
    n2569, n2570, n2571, n2572, n2573, n2574,
    n2575, n2576, n2577, n2578, n2579, n2580,
    n2581, n2582, n2583, n2584, n2585, n2586,
    n2587, n2588, n2589, n2590, n2591, n2592,
    n2593, n2594, n2595, n2596, n2597, n2598,
    n2599, n2600, n2601, n2602, n2603, n2604,
    n2605, n2606, n2607, n2608, n2609, n2610,
    n2611, n2612, n2613, n2614, n2615, n2616,
    n2617, n2618, n2619, n2620, n2621, n2622,
    n2623, n2624, n2625, n2626, n2627, n2628,
    n2629, n2630, n2631, n2632, n2633, n2634,
    n2635, n2636, n2637, n2638, n2639, n2640,
    n2641, n2642, n2643, n2644, n2645, n2646,
    n2647, n2648, n2649, n2650, n2651, n2652,
    n2653, n2654, n2655, n2656, n2657, n2658,
    n2659, n2660, n2661, n2662, n2663, n2664,
    n2665, n2666, n2667, n2668, n2669, n2670,
    n2671, n2672, n2673, n2674, n2675, n2676,
    n2677, n2678, n2679, n2680, n2681, n2682,
    n2683, n2684, n2685, n2686, n2687, n2688,
    n2689, n2690, n2691, n2692, n2693, n2694,
    n2695, n2696, n2697, n2698, n2699, n2700,
    n2701, n2702, n2703, n2704, n2705, n2706,
    n2707, n2708, n2709, n2710, n2711, n2712,
    n2713, n2714, n2715, n2716, n2717, n2718,
    n2719, n2720, n2721, n2722, n2723, n2724,
    n2725, n2726, n2727, n2728, n2729, n2730,
    n2731, n2732, n2733, n2734, n2735, n2736,
    n2737, n2738, n2739, n2740, n2741, n2742,
    n2743, n2744, n2745, n2746, n2747, n2748,
    n2749, n2750, n2751, n2752, n2753, n2754,
    n2755, n2756, n2757, n2758, n2759, n2760,
    n2761, n2762, n2763, n2764, n2765, n2766,
    n2767, n2768, n2769, n2770, n2771, n2772,
    n2773, n2774, n2775, n2776, n2777, n2778,
    n2779, n2780, n2781, n2782, n2783, n2784,
    n2785, n2786, n2787, n2788, n2789, n2790,
    n2791, n2792, n2793, n2794, n2795, n2796,
    n2797, n2798, n2799, n2800, n2801, n2802,
    n2803, n2804, n2805, n2806, n2807, n2808,
    n2809, n2810, n2811, n2812, n2813, n2814,
    n2815, n2816, n2817, n2818, n2819, n2820,
    n2821, n2822, n2823, n2824, n2825, n2826,
    n2827, n2828, n2829, n2830, n2831, n2832,
    n2833, n2834, n2835, n2836, n2837, n2838,
    n2839, n2840, n2841, n2842, n2843, n2844,
    n2845, n2846, n2847, n2848, n2849, n2850,
    n2851, n2852, n2853, n2854, n2855, n2856,
    n2857, n2858, n2859, n2860, n2861, n2862,
    n2863, n2864, n2865, n2866, n2867, n2868,
    n2869, n2870, n2871, n2872, n2873, n2874,
    n2875, n2876, n2877, n2878, n2879, n2880,
    n2881, n2882, n2883, n2884, n2885, n2886,
    n2887, n2888, n2889, n2890, n2891, n2892,
    n2893, n2894, n2895, n2896, n2897, n2898,
    n2899, n2900, n2901, n2902, n2903, n2904,
    n2905, n2906, n2907, n2908, n2909, n2910,
    n2911, n2912, n2913, n2914, n2915, n2916,
    n2917, n2918, n2919, n2920, n2921, n2922,
    n2923, n2924, n2925, n2926, n2927, n2928,
    n2929, n2930, n2931, n2932, n2933, n2934,
    n2935, n2936, n2937, n2938, n2939, n2940,
    n2941, n2942, n2943, n2944, n2945, n2946,
    n2947, n2948, n2949, n2950, n2951, n2952,
    n2953, n2954, n2955, n2956, n2957, n2958,
    n2959, n2960, n2961, n2962, n2963, n2964,
    n2965, n2966, n2967, n2968, n2969, n2970,
    n2971, n2972, n2973, n2974, n2975, n2976,
    n2977, n2978, n2979, n2980, n2981, n2982,
    n2983, n2984, n2985, n2986, n2987, n2988,
    n2989, n2990, n2991, n2992, n2993, n2994,
    n2995, n2996, n2997, n2998, n2999, n3000,
    n3001, n3002, n3003, n3004, n3005, n3006,
    n3007, n3008, n3009, n3010, n3011, n3012,
    n3013, n3014, n3015, n3016, n3017, n3018,
    n3019, n3020, n3021, n3022, n3023, n3024,
    n3025, n3026, n3027, n3028, n3029, n3030,
    n3031, n3032, n3033, n3034, n3035, n3036,
    n3037, n3038, n3039, n3040, n3041, n3042,
    n3043, n3044, n3045, n3046, n3047, n3048,
    n3049, n3050, n3051, n3052, n3053, n3054,
    n3055, n3056, n3057, n3058, n3059, n3060,
    n3061, n3062, n3063, n3064, n3065, n3066,
    n3067, n3068, n3069, n3070, n3071, n3072,
    n3073, n3074, n3075, n3076, n3077, n3078,
    n3079, n3080, n3081, n3082, n3083, n3084,
    n3085, n3086, n3087, n3088, n3089, n3090,
    n3091, n3092, n3093, n3094, n3095, n3096,
    n3097, n3098, n3099, n3100, n3101, n3102,
    n3103, n3104, n3105, n3106, n3107, n3108,
    n3109, n3110, n3111, n3112, n3113, n3114,
    n3115, n3116, n3117, n3118, n3119, n3120,
    n3121, n3122, n3123, n3124, n3125, n3126,
    n3127, n3128, n3129, n3130, n3131, n3132,
    n3133, n3134, n3135, n3136, n3137, n3138,
    n3139, n3140, n3141, n3142, n3143, n3144,
    n3145, n3146, n3147, n3148, n3149, n3150,
    n3151, n3152, n3153, n3154, n3155, n3156,
    n3157, n3158, n3159, n3160, n3161, n3162,
    n3163, n3164, n3165, n3166, n3167, n3168,
    n3169, n3170, n3171, n3172, n3173, n3174,
    n3175, n3176, n3177, n3178, n3179, n3180,
    n3181, n3182, n3183, n3184, n3185, n3186,
    n3187, n3188, n3189, n3190, n3191, n3192,
    n3193, n3194, n3195, n3196, n3197, n3198,
    n3199, n3200, n3201, n3202, n3203, n3204,
    n3205, n3206, n3207, n3208, n3209, n3210,
    n3211, n3212, n3213, n3214, n3215, n3216,
    n3217, n3218, n3219, n3220, n3221, n3222,
    n3223, n3224, n3225, n3226, n3227, n3228,
    n3229, n3230, n3231, n3232, n3233, n3234,
    n3235, n3236, n3237, n3238, n3239, n3240,
    n3241, n3242, n3243, n3244, n3245, n3246,
    n3247, n3248, n3249, n3250, n3251, n3252,
    n3253, n3254, n3255, n3256, n3257, n3258,
    n3259, n3260, n3261, n3262, n3263, n3264,
    n3265, n3266, n3267, n3268, n3269, n3270,
    n3271, n3272, n3273, n3274, n3275, n3276,
    n3277, n3278, n3279, n3280, n3281, n3282,
    n3283, n3284, n3285, n3286, n3287, n3288,
    n3289, n3291, n3292, n3293, n3294, n3295,
    n3296, n3297, n3298, n3299, n3300, n3301,
    n3302, n3303, n3304, n3305, n3306, n3307,
    n3308, n3309, n3310, n3311, n3312, n3313,
    n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325,
    n3326, n3327, n3328, n3329, n3330, n3331,
    n3332, n3333, n3334, n3335, n3336, n3337,
    n3338, n3339, n3340, n3341, n3342, n3343,
    n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355,
    n3356, n3357, n3358, n3359, n3360, n3361,
    n3362, n3363, n3364, n3365, n3366, n3367,
    n3368, n3369, n3370, n3371, n3372, n3373,
    n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385,
    n3386, n3387, n3388, n3389, n3390, n3391,
    n3392, n3393, n3394, n3395, n3396, n3397,
    n3398, n3399, n3400, n3401, n3402, n3403,
    n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415,
    n3416, n3417, n3418, n3419, n3420, n3421,
    n3422, n3423, n3424, n3425, n3426, n3427,
    n3428, n3429, n3430, n3431, n3432, n3433,
    n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445,
    n3446, n3447, n3448, n3449, n3450, n3451,
    n3452, n3453, n3454, n3455, n3456, n3457,
    n3458, n3459, n3460, n3461, n3462, n3463,
    n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475,
    n3476, n3477, n3478, n3479, n3480, n3481,
    n3482, n3483, n3484, n3485, n3486, n3487,
    n3488, n3489, n3490, n3491, n3492, n3493,
    n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3506,
    n3507, n3508, n3509, n3510, n3511, n3512,
    n3513, n3514, n3515, n3516, n3517, n3518,
    n3519, n3520, n3521, n3522, n3523, n3524,
    n3525, n3526, n3527, n3528, n3529, n3530,
    n3531, n3532, n3533, n3534, n3535, n3536,
    n3537, n3538, n3539, n3540, n3541, n3542,
    n3543, n3544, n3545, n3546, n3547, n3548,
    n3549, n3550, n3551, n3552, n3553, n3554,
    n3555, n3556, n3557, n3558, n3559, n3560,
    n3561, n3562, n3563, n3564, n3565, n3566,
    n3567, n3568, n3569, n3570, n3571, n3572,
    n3573, n3574, n3575, n3576, n3577, n3578,
    n3579, n3580, n3581, n3582, n3583, n3584,
    n3585, n3586, n3587, n3588, n3589, n3590,
    n3591, n3592, n3593, n3594, n3595, n3596,
    n3597, n3598, n3599, n3600, n3601, n3602,
    n3603, n3604, n3605, n3606, n3607, n3608,
    n3609, n3610, n3611, n3612, n3613, n3614,
    n3615, n3616, n3617, n3618, n3619, n3620,
    n3621, n3622, n3623, n3624, n3625, n3626,
    n3627, n3628, n3629, n3630, n3631, n3632,
    n3633, n3634, n3635, n3636, n3637, n3638,
    n3639, n3640, n3641, n3642, n3643, n3644,
    n3645, n3646, n3647, n3648, n3649, n3650,
    n3651, n3652, n3653, n3654, n3655, n3656,
    n3657, n3658, n3659, n3660, n3661, n3662,
    n3663, n3664, n3665, n3666, n3667, n3668,
    n3669, n3670, n3671, n3672, n3673, n3674,
    n3675, n3676, n3677, n3679, n3680, n3681,
    n3682, n3683, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3908, n3909, n3910,
    n3911, n3912, n3913, n3914, n3915, n3916,
    n3917, n3918, n3919, n3920, n3921, n3922,
    n3923, n3924, n3925, n3926, n3927, n3928,
    n3929, n3930, n3931, n3932, n3933, n3934,
    n3935, n3936, n3937, n3938, n3939, n3940,
    n3941, n3942, n3943, n3944, n3945, n3946,
    n3947, n3948, n3949, n3950, n3951, n3952,
    n3953, n3954, n3955, n3956, n3957, n3958,
    n3959, n3960, n3961, n3962, n3963, n3964,
    n3965, n3966, n3967, n3968, n3969, n3970,
    n3971, n3972, n3973, n3974, n3975, n3976,
    n3977, n3978, n3979, n3980, n3981, n3982,
    n3983, n3984, n3985, n3986, n3987, n3988,
    n3989, n3990, n3991, n3992, n3993, n3994,
    n3995, n3996, n3997, n3998, n3999, n4000,
    n4001, n4002, n4003, n4004, n4005, n4006,
    n4007, n4008, n4009, n4010, n4011, n4012,
    n4013, n4014, n4015, n4016, n4017, n4018,
    n4019, n4020, n4021, n4022, n4023, n4024,
    n4025, n4026, n4027, n4028, n4029, n4030,
    n4031, n4032, n4033, n4034, n4035, n4036,
    n4037, n4038, n4039, n4040, n4041, n4042,
    n4043, n4044, n4045, n4046, n4047, n4048,
    n4049, n4050, n4051, n4052, n4053, n4054,
    n4055, n4056, n4057, n4058, n4059, n4060,
    n4061, n4062, n4063, n4064, n4065, n4066,
    n4067, n4068, n4069, n4070, n4071, n4072,
    n4073, n4074, n4075, n4076, n4077, n4078,
    n4079, n4080, n4081, n4082, n4083, n4084,
    n4085, n4086, n4087, n4088, n4089, n4090,
    n4091, n4092, n4093, n4094, n4095, n4096,
    n4097, n4098, n4099, n4100, n4101, n4102,
    n4103, n4104, n4105, n4106, n4107, n4108,
    n4109, n4110, n4111, n4112, n4113, n4114,
    n4115, n4116, n4117, n4118, n4119, n4120,
    n4121, n4122, n4123, n4124, n4125, n4126,
    n4127, n4128, n4129, n4130, n4131, n4132,
    n4133, n4135, n4136, n4137, n4138, n4139,
    n4140, n4141, n4142, n4143, n4144, n4145,
    n4146, n4147, n4148, n4149, n4150, n4151,
    n4152, n4153, n4154, n4155, n4156, n4157,
    n4158, n4159, n4160, n4161, n4162, n4163,
    n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175,
    n4176, n4177, n4178, n4179, n4180, n4181,
    n4182, n4183, n4184, n4185, n4186, n4187,
    n4188, n4189, n4190, n4191, n4192, n4193,
    n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205,
    n4206, n4207, n4208, n4209, n4210, n4211,
    n4212, n4213, n4214, n4215, n4216, n4217,
    n4218, n4219, n4220, n4221, n4222, n4223,
    n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235,
    n4236, n4237, n4238, n4239, n4240, n4241,
    n4242, n4243, n4244, n4245, n4246, n4247,
    n4248, n4249, n4250, n4251, n4252, n4253,
    n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265,
    n4266, n4267, n4268, n4269, n4270, n4271,
    n4272, n4273, n4274, n4275, n4276, n4277,
    n4278, n4279, n4280, n4281, n4282, n4283,
    n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295,
    n4296, n4297, n4298, n4299, n4300, n4301,
    n4302, n4303, n4304, n4305, n4306, n4307,
    n4308, n4309, n4310, n4311, n4312, n4313,
    n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325,
    n4326, n4327, n4328, n4329, n4330, n4331,
    n4332, n4333, n4334, n4335, n4336, n4337,
    n4338, n4339, n4340, n4341, n4342, n4343,
    n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355,
    n4357, n4358, n4359, n4360, n4361, n4362,
    n4363, n4364, n4365, n4366, n4367, n4368,
    n4369, n4370, n4371, n4372, n4373, n4374,
    n4375, n4376, n4377, n4378, n4379, n4380,
    n4381, n4382, n4383, n4384, n4385, n4386,
    n4387, n4388, n4389, n4390, n4391, n4392,
    n4393, n4394, n4395, n4396, n4397, n4398,
    n4399, n4400, n4401, n4402, n4403, n4404,
    n4405, n4406, n4407, n4408, n4409, n4410,
    n4411, n4412, n4413, n4414, n4415, n4416,
    n4417, n4418, n4419, n4420, n4421, n4422,
    n4423, n4424, n4425, n4426, n4427, n4428,
    n4429, n4430, n4431, n4432, n4433, n4434,
    n4435, n4436, n4437, n4438, n4439, n4440,
    n4441, n4442, n4443, n4444, n4445, n4446,
    n4447, n4448, n4449, n4450, n4451, n4452,
    n4453, n4454, n4455, n4456, n4457, n4458,
    n4459, n4460, n4461, n4462, n4463, n4464,
    n4465, n4466, n4467, n4468, n4469, n4470,
    n4471, n4472, n4473, n4474, n4475, n4476,
    n4477, n4478, n4479, n4480, n4481, n4482,
    n4483, n4484, n4485, n4486, n4487, n4488,
    n4489, n4490, n4491, n4492, n4493, n4494,
    n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506,
    n4507, n4508, n4509, n4510, n4511, n4512,
    n4513, n4514, n4515, n4516, n4517, n4518,
    n4519, n4520, n4521, n4522, n4523, n4524,
    n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536,
    n4537, n4538, n4539, n4540, n4541, n4542,
    n4543, n4544, n4545, n4546, n4547, n4548,
    n4549, n4550, n4551, n4552, n4553, n4554,
    n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4579,
    n4580, n4581, n4582, n4583, n4584, n4585,
    n4586, n4587, n4588, n4589, n4590, n4591,
    n4592, n4593, n4594, n4595, n4596, n4597,
    n4598, n4599, n4600, n4601, n4602, n4603,
    n4604, n4605, n4606, n4607, n4608, n4609,
    n4610, n4611, n4612, n4613, n4614, n4615,
    n4616, n4617, n4618, n4619, n4620, n4621,
    n4622, n4623, n4624, n4625, n4626, n4627,
    n4628, n4629, n4630, n4631, n4632, n4633,
    n4634, n4635, n4636, n4637, n4638, n4639,
    n4640, n4641, n4642, n4643, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4720, n4721, n4722, n4723,
    n4724, n4725, n4726, n4727, n4728, n4729,
    n4730, n4731, n4732, n4733, n4734, n4735,
    n4736, n4737, n4738, n4739, n4740, n4741,
    n4742, n4743, n4744, n4745, n4746, n4747,
    n4748, n4749, n4750, n4751, n4752, n4753,
    n4754, n4755, n4756, n4757, n4758, n4759,
    n4760, n4761, n4762, n4763, n4764, n4765,
    n4766, n4767, n4768, n4769, n4770, n4771,
    n4772, n4773, n4774, n4775, n4776, n4777,
    n4778, n4779, n4780, n4781, n4782, n4783,
    n4784, n4785, n4786, n4787, n4788, n4789,
    n4790, n4791, n4792, n4793, n4794, n4795,
    n4796, n4797, n4798, n4799, n4800, n4801,
    n4803, n4804, n4805, n4806, n4807, n4808,
    n4809, n4810, n4811, n4812, n4813, n4814,
    n4815, n4816, n4817, n4818, n4819, n4820,
    n4821, n4822, n4823, n4824, n4825, n4826,
    n4827, n4828, n4829, n4830, n4831, n4832,
    n4833, n4834, n4835, n4836, n4837, n4838,
    n4839, n4840, n4841, n4842, n4843, n4844,
    n4845, n4846, n4847, n4848, n4849, n4850,
    n4851, n4852, n4853, n4854, n4855, n4856,
    n4857, n4858, n4859, n4860, n4861, n4862,
    n4863, n4864, n4865, n4866, n4867, n4868,
    n4869, n4870, n4871, n4872, n4873, n4874,
    n4875, n4876, n4877, n4878, n4879, n4880,
    n4881, n4882, n4883, n4884, n4885, n4886,
    n4887, n4888, n4889, n4890, n4891, n4892,
    n4893, n4894, n4895, n4896, n4897, n4898,
    n4899, n4900, n4901, n4902, n4903, n4904,
    n4905, n4906, n4907, n4908, n4909, n4910,
    n4911, n4912, n4913, n4914, n4915, n4916,
    n4917, n4918, n4919, n4920, n4921, n4922,
    n4923, n4924, n4925, n4926, n4927, n4928,
    n4929, n4930, n4931, n4932, n4933, n4934,
    n4935, n4936, n4937, n4938, n4939, n4940,
    n4941, n4942, n4943, n4944, n4945, n4946,
    n4947, n4948, n4949, n4950, n4951, n4952,
    n4953, n4954, n4955, n4956, n4957, n4958,
    n4959, n4960, n4961, n4962, n4963, n4964,
    n4965, n4966, n4967, n4968, n4969, n4970,
    n4971, n4972, n4973, n4974, n4975, n4976,
    n4977, n4978, n4979, n4980, n4981, n4982,
    n4983, n4984, n4985, n4986, n4987, n4988,
    n4989, n4990, n4991, n4992, n4993, n4994,
    n4995, n4996, n4997, n4998, n4999, n5000,
    n5001, n5002, n5003, n5004, n5005, n5006,
    n5007, n5008, n5009, n5010, n5011, n5012,
    n5013, n5014, n5015, n5016, n5017, n5018,
    n5019, n5020, n5021, n5022, n5024, n5025,
    n5026, n5027, n5028, n5029, n5030, n5031,
    n5032, n5033, n5034, n5035, n5036, n5037,
    n5038, n5039, n5040, n5041, n5042, n5043,
    n5044, n5045, n5046, n5047, n5048, n5049,
    n5050, n5051, n5052, n5053, n5054, n5055,
    n5056, n5057, n5058, n5059, n5060, n5061,
    n5062, n5063, n5064, n5065, n5066, n5067,
    n5068, n5069, n5070, n5071, n5072, n5073,
    n5074, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5094, n5095, n5096, n5097,
    n5098, n5099, n5100, n5101, n5102, n5103,
    n5104, n5105, n5106, n5107, n5108, n5109,
    n5110, n5111, n5112, n5113, n5114, n5115,
    n5116, n5117, n5118, n5119, n5120, n5121,
    n5122, n5123, n5124, n5125, n5126, n5127,
    n5128, n5129, n5130, n5131, n5132, n5133,
    n5134, n5135, n5136, n5137, n5138, n5139,
    n5140, n5141, n5142, n5143, n5144, n5145,
    n5146, n5147, n5148, n5149, n5150, n5151,
    n5152, n5153, n5154, n5155, n5156, n5157,
    n5158, n5159, n5160, n5161, n5162, n5163,
    n5164, n5165, n5166, n5167, n5168, n5169,
    n5170, n5171, n5172, n5173, n5174, n5175,
    n5176, n5177, n5178, n5179, n5180, n5181,
    n5182, n5183, n5184, n5185, n5186, n5187,
    n5188, n5189, n5190, n5191, n5192, n5193,
    n5194, n5195, n5196, n5197, n5198, n5199,
    n5200, n5201, n5202, n5203, n5204, n5205,
    n5206, n5207, n5208, n5209, n5210, n5211,
    n5212, n5213, n5214, n5215, n5216, n5217,
    n5218, n5219, n5220, n5221, n5222, n5223,
    n5224, n5225, n5226, n5227, n5228, n5229,
    n5230, n5231, n5232, n5233, n5234, n5235,
    n5236, n5237, n5238, n5239, n5240, n5241,
    n5242, n5243, n5245, n5246, n5247, n5248,
    n5249, n5250, n5251, n5252, n5253, n5254,
    n5255, n5256, n5257, n5258, n5259, n5260,
    n5261, n5262, n5263, n5264, n5265, n5266,
    n5267, n5268, n5269, n5270, n5271, n5272,
    n5273, n5274, n5275, n5276, n5277, n5278,
    n5279, n5280, n5281, n5282, n5283, n5284,
    n5285, n5286, n5287, n5288, n5289, n5290,
    n5291, n5292, n5293, n5294, n5295, n5296,
    n5297, n5298, n5299, n5300, n5301, n5302,
    n5303, n5304, n5305, n5306, n5307, n5308,
    n5309, n5310, n5311, n5312, n5313, n5314,
    n5315, n5316, n5317, n5318, n5319, n5320,
    n5321, n5322, n5323, n5324, n5325, n5326,
    n5327, n5328, n5329, n5330, n5331, n5332,
    n5333, n5334, n5335, n5336, n5337, n5338,
    n5339, n5340, n5341, n5342, n5343, n5344,
    n5345, n5346, n5347, n5348, n5349, n5350,
    n5351, n5352, n5353, n5354, n5355, n5356,
    n5357, n5358, n5359, n5360, n5361, n5362,
    n5363, n5364, n5365, n5366, n5367, n5368,
    n5369, n5370, n5371, n5372, n5373, n5374,
    n5375, n5376, n5377, n5378, n5379, n5380,
    n5381, n5382, n5383, n5384, n5385, n5386,
    n5387, n5388, n5389, n5390, n5391, n5392,
    n5393, n5394, n5395, n5396, n5397, n5398,
    n5399, n5400, n5401, n5402, n5403, n5404,
    n5405, n5406, n5407, n5408, n5409, n5410,
    n5411, n5412, n5413, n5414, n5415, n5416,
    n5417, n5418, n5419, n5420, n5421, n5422,
    n5423, n5424, n5425, n5426, n5427, n5428,
    n5429, n5430, n5431, n5432, n5433, n5434,
    n5435, n5436, n5437, n5438, n5439, n5440,
    n5441, n5442, n5443, n5444, n5445, n5446,
    n5447, n5448, n5449, n5450, n5451, n5452,
    n5453, n5454, n5455, n5456, n5457, n5458,
    n5459, n5460, n5461, n5462, n5463, n5464,
    n5465, n5466, n5467, n5468, n5469, n5470,
    n5471, n5472, n5473, n5474, n5475, n5476,
    n5477, n5479, n5480, n5481, n5482, n5483,
    n5484, n5485, n5486, n5487, n5488, n5489,
    n5490, n5491, n5492, n5493, n5494, n5495,
    n5496, n5497, n5498, n5499, n5500, n5501,
    n5502, n5503, n5504, n5505, n5506, n5507,
    n5508, n5509, n5510, n5511, n5512, n5513,
    n5514, n5515, n5516, n5517, n5518, n5519,
    n5520, n5521, n5522, n5523, n5524, n5525,
    n5526, n5527, n5528, n5529, n5530, n5531,
    n5532, n5533, n5534, n5535, n5536, n5537,
    n5538, n5539, n5540, n5541, n5542, n5543,
    n5544, n5545, n5546, n5547, n5548, n5549,
    n5550, n5551, n5552, n5553, n5554, n5555,
    n5556, n5557, n5558, n5559, n5560, n5561,
    n5562, n5563, n5564, n5565, n5566, n5567,
    n5568, n5569, n5570, n5571, n5572, n5573,
    n5574, n5575, n5576, n5577, n5578, n5579,
    n5580, n5581, n5582, n5583, n5584, n5585,
    n5586, n5587, n5588, n5589, n5590, n5591,
    n5592, n5593, n5594, n5595, n5596, n5597,
    n5598, n5599, n5600, n5601, n5602, n5603,
    n5604, n5605, n5606, n5607, n5608, n5609,
    n5610, n5611, n5612, n5613, n5614, n5615,
    n5616, n5617, n5618, n5619, n5620, n5621,
    n5622, n5623, n5624, n5625, n5626, n5627,
    n5628, n5629, n5630, n5631, n5632, n5633,
    n5634, n5635, n5636, n5637, n5638, n5639,
    n5640, n5641, n5642, n5643, n5644, n5645,
    n5646, n5647, n5648, n5649, n5650, n5651,
    n5652, n5653, n5654, n5655, n5656, n5657,
    n5658, n5659, n5660, n5661, n5662, n5663,
    n5664, n5665, n5666, n5667, n5668, n5669,
    n5670, n5671, n5672, n5673, n5674, n5675,
    n5676, n5677, n5678, n5679, n5680, n5681,
    n5682, n5683, n5684, n5685, n5686, n5687,
    n5688, n5689, n5690, n5691, n5692, n5693,
    n5694, n5695, n5696, n5697, n5698, n5699,
    n5700, n5701, n5702, n5703, n5704, n5705,
    n5706, n5707, n5708, n5709, n5710, n5712,
    n5713, n5714, n5715, n5716, n5717, n5718,
    n5719, n5720, n5721, n5722, n5723, n5724,
    n5725, n5726, n5727, n5728, n5729, n5730,
    n5731, n5732, n5733, n5734, n5735, n5736,
    n5737, n5738, n5739, n5740, n5741, n5742,
    n5743, n5744, n5745, n5746, n5747, n5748,
    n5749, n5750, n5751, n5752, n5753, n5754,
    n5755, n5756, n5757, n5758, n5759, n5760,
    n5761, n5762, n5763, n5764, n5765, n5766,
    n5767, n5768, n5769, n5770, n5771, n5772,
    n5773, n5774, n5775, n5776, n5777, n5778,
    n5779, n5780, n5781, n5782, n5783, n5784,
    n5785, n5786, n5787, n5788, n5789, n5790,
    n5791, n5792, n5793, n5794, n5795, n5796,
    n5797, n5798, n5799, n5800, n5801, n5802,
    n5803, n5804, n5805, n5806, n5807, n5808,
    n5809, n5810, n5811, n5812, n5813, n5814,
    n5815, n5816, n5817, n5818, n5819, n5820,
    n5821, n5822, n5823, n5824, n5825, n5826,
    n5827, n5828, n5829, n5830, n5831, n5832,
    n5833, n5834, n5835, n5836, n5837, n5838,
    n5839, n5840, n5841, n5842, n5843, n5844,
    n5845, n5846, n5847, n5848, n5849, n5850,
    n5851, n5852, n5853, n5854, n5855, n5856,
    n5857, n5858, n5859, n5860, n5861, n5862,
    n5863, n5864, n5865, n5866, n5867, n5868,
    n5869, n5870, n5871, n5872, n5873, n5874,
    n5875, n5876, n5877, n5878, n5879, n5880,
    n5881, n5882, n5883, n5884, n5885, n5886,
    n5887, n5888, n5889, n5890, n5891, n5892,
    n5893, n5894, n5895, n5896, n5897, n5898,
    n5899, n5900, n5901, n5902, n5903, n5904,
    n5905, n5906, n5907, n5908, n5909, n5910,
    n5911, n5912, n5913, n5914, n5915, n5916,
    n5917, n5918, n5919, n5920, n5921, n5922,
    n5923, n5924, n5925, n5926, n5927, n5928,
    n5929, n5930, n5931, n5932, n5933, n5934,
    n5935, n5936, n5937, n5938, n5939, n5940,
    n5941, n5942, n5943, n5944, n5945, n5946,
    n5947, n5948, n5949, n5950, n5951, n5952,
    n5953, n5954, n5955, n5956, n5957, n5958,
    n5959, n5960, n5961, n5962, n5963, n5964,
    n5965, n5966, n5967, n5968, n5969, n5970,
    n5971, n5972, n5973, n5974, n5975, n5976,
    n5977, n5978, n5979, n5980, n5981, n5982,
    n5983, n5984, n5985, n5986, n5987, n5988,
    n5989, n5990, n5991, n5992, n5993, n5994,
    n5995, n5996, n5997, n5998, n5999, n6000,
    n6001, n6002, n6003, n6004, n6005, n6006,
    n6007, n6008, n6009, n6010, n6011, n6012,
    n6013, n6014, n6015, n6016, n6017, n6018,
    n6019, n6020, n6021, n6022, n6023, n6024,
    n6025, n6026, n6027, n6028, n6029, n6030,
    n6031, n6032, n6033, n6034, n6035, n6036,
    n6037, n6038, n6039, n6040, n6041, n6042,
    n6043, n6044, n6045, n6046, n6047, n6048,
    n6049, n6050, n6051, n6052, n6053, n6054,
    n6055, n6056, n6057, n6058, n6059, n6060,
    n6061, n6062, n6063, n6064, n6065, n6066,
    n6068, n6069, n6070, n6071, n6072, n6073,
    n6074, n6075, n6076, n6077, n6078, n6079,
    n6080, n6081, n6082, n6083, n6084, n6085,
    n6086, n6087, n6088, n6089, n6090, n6091,
    n6092, n6093, n6094, n6095, n6096, n6097,
    n6098, n6099, n6101, n6102, n6103, n6104,
    n6106, n6107, n6108, n6109, n6110, n6111,
    n6112, n6113, n6114, n6115, n6116, n6117,
    n6118, n6119, n6120, n6121, n6122, n6123,
    n6124, n6125, n6126, n6127, n6128, n6129,
    n6130, n6131, n6132, n6133, n6134, n6135,
    n6136, n6137, n6138, n6139, n6140, n6141,
    n6142, n6143, n6144, n6145, n6146, n6147,
    n6148, n6149, n6150, n6151, n6152, n6153,
    n6154, n6155, n6156, n6157, n6158, n6159,
    n6160, n6161, n6162, n6163, n6164, n6166,
    n6167, n6168, n6169, n6170, n6171, n6172,
    n6173, n6174, n6175, n6176, n6177, n6178,
    n6179, n6180, n6181, n6182, n6183, n6184,
    n6185, n6186, n6187, n6188, n6189, n6190,
    n6191, n6192, n6193, n6194, n6195, n6196,
    n6197, n6198, n6199, n6200, n6201, n6202,
    n6203, n6204, n6205, n6206, n6207, n6208,
    n6209, n6210, n6211, n6212, n6213, n6214,
    n6215, n6216, n6217, n6218, n6219, n6220,
    n6221, n6222, n6223, n6224, n6225, n6226,
    n6227, n6228, n6229, n6230, n6231, n6232,
    n6233, n6234, n6235, n6236, n6237, n6238,
    n6239, n6240, n6241, n6242, n6243, n6244,
    n6245, n6246, n6247, n6248, n6249, n6250,
    n6251, n6252, n6253, n6254, n6255, n6257,
    n6258, n6259, n6260, n6261, n6262, n6263,
    n6264, n6265, n6266, n6267, n6268, n6269,
    n6270, n6271, n6272, n6273, n6274, n6275,
    n6276, n6277, n6278, n6279, n6280, n6281,
    n6282, n6283, n6284, n6285, n6286, n6287,
    n6288, n6289, n6290, n6291, n6292, n6293,
    n6294, n6295, n6296, n6297, n6298, n6299,
    n6300, n6301, n6302, n6303, n6304, n6305,
    n6306, n6307, n6308, n6309, n6310, n6311,
    n6312, n6313, n6314, n6315, n6316, n6317,
    n6318, n6319, n6320, n6321, n6322, n6323,
    n6324, n6325, n6326, n6327, n6328, n6329,
    n6330, n6331, n6332, n6333, n6334, n6335,
    n6336, n6337, n6338, n6339, n6340, n6341,
    n6342, n6343, n6344, n6345, n6346, n6347,
    n6348, n6349, n6350, n6351, n6352, n6353,
    n6354, n6355, n6356, n6357, n6358, n6359,
    n6360, n6361, n6362, n6363, n6364, n6365,
    n6366, n6367, n6368, n6369, n6370, n6371,
    n6372, n6373, n6374, n6375, n6376, n6377,
    n6378, n6379, n6380, n6381, n6382, n6383,
    n6384, n6385, n6386, n6387, n6389, n6390,
    n6391, n6392, n6393, n6394, n6395, n6396,
    n6397, n6398, n6399, n6400, n6401, n6402,
    n6403, n6404, n6405, n6406, n6407, n6408,
    n6409, n6410, n6411, n6412, n6413, n6414,
    n6415, n6416, n6417, n6418, n6419, n6420,
    n6421, n6422, n6423, n6424, n6425, n6426,
    n6427, n6428, n6429, n6430, n6431, n6432,
    n6433, n6434, n6435, n6436, n6437, n6438,
    n6439, n6440, n6441, n6442, n6443, n6444,
    n6445, n6446, n6447, n6448, n6449, n6450,
    n6451, n6452, n6453, n6454, n6455, n6456,
    n6457, n6458, n6459, n6460, n6461, n6462,
    n6463, n6464, n6465, n6466, n6467, n6468,
    n6469, n6470, n6471, n6472, n6473, n6474,
    n6475, n6476, n6477, n6478, n6479, n6480,
    n6481, n6482, n6483, n6484, n6485, n6486,
    n6487, n6488, n6489, n6490, n6491, n6492,
    n6493, n6494, n6495, n6496, n6497, n6498,
    n6499, n6500, n6501, n6502, n6503, n6504,
    n6505, n6506, n6507, n6508, n6509, n6510,
    n6511, n6512, n6513, n6514, n6515, n6516,
    n6517, n6518, n6519, n6520, n6521, n6522,
    n6524, n6525, n6526, n6527, n6528, n6529,
    n6530, n6531, n6532, n6533, n6534, n6535,
    n6536, n6537, n6538, n6539, n6540, n6541,
    n6542, n6543, n6544, n6545, n6546, n6547,
    n6548, n6549, n6550, n6551, n6552, n6553,
    n6554, n6555, n6556, n6557, n6558, n6559,
    n6560, n6561, n6562, n6563, n6564, n6565,
    n6566, n6567, n6568, n6569, n6570, n6571,
    n6572, n6573, n6574, n6575, n6576, n6577,
    n6578, n6579, n6580, n6581, n6582, n6583,
    n6584, n6585, n6586, n6587, n6588, n6589,
    n6590, n6591, n6592, n6593, n6594, n6595,
    n6596, n6597, n6598, n6599, n6600, n6601,
    n6602, n6603, n6604, n6605, n6606, n6607,
    n6608, n6609, n6610, n6611, n6612, n6613,
    n6614, n6615, n6616, n6617, n6618, n6619,
    n6620, n6621, n6622, n6623, n6624, n6625,
    n6626, n6627, n6628, n6629, n6630, n6631,
    n6632, n6633, n6634, n6635, n6636, n6637,
    n6638, n6639, n6640, n6641, n6642, n6643,
    n6644, n6645, n6647, n6648, n6649, n6650,
    n6651, n6652, n6653, n6654, n6655, n6656,
    n6657, n6658, n6659, n6660, n6661, n6662,
    n6663, n6664, n6665, n6666, n6667, n6668,
    n6669, n6670, n6671, n6672, n6673, n6674,
    n6675, n6676, n6677, n6678, n6679, n6680,
    n6681, n6682, n6683, n6684, n6685, n6686,
    n6687, n6688, n6689, n6690, n6691, n6692,
    n6693, n6694, n6695, n6696, n6697, n6698,
    n6699, n6700, n6701, n6702, n6703, n6704,
    n6705, n6706, n6707, n6708, n6709, n6710,
    n6711, n6712, n6713, n6714, n6715, n6716,
    n6717, n6718, n6719, n6720, n6721, n6722,
    n6723, n6724, n6725, n6726, n6727, n6728,
    n6729, n6730, n6731, n6732, n6733, n6734,
    n6735, n6736, n6737, n6738, n6739, n6740,
    n6741, n6742, n6743, n6744, n6745, n6746,
    n6747, n6748, n6749, n6750, n6751, n6752,
    n6753, n6754, n6755, n6756, n6757, n6758,
    n6759, n6760, n6761, n6762, n6763, n6764,
    n6765, n6766, n6767, n6768, n6769, n6770,
    n6771, n6773, n6774, n6775, n6776, n6777,
    n6778, n6779, n6780, n6781, n6782, n6783,
    n6784, n6785, n6786, n6787, n6788, n6789,
    n6790, n6791, n6792, n6793, n6794, n6795,
    n6796, n6797, n6798, n6799, n6800, n6801,
    n6802, n6803, n6804, n6805, n6806, n6807,
    n6808, n6809, n6810, n6811, n6812, n6813,
    n6814, n6815, n6816, n6817, n6818, n6819,
    n6820, n6821, n6822, n6823, n6824, n6825,
    n6826, n6827, n6828, n6829, n6830, n6831,
    n6832, n6833, n6834, n6835, n6836, n6837,
    n6838, n6839, n6840, n6841, n6842, n6843,
    n6844, n6845, n6846, n6847, n6848, n6849,
    n6850, n6851, n6852, n6853, n6854, n6855,
    n6856, n6857, n6858, n6859, n6860, n6861,
    n6862, n6864, n6865, n6866, n6867, n6868,
    n6869, n6870, n6871, n6872, n6873, n6874,
    n6875, n6876, n6877, n6878, n6879, n6880,
    n6881, n6882, n6883, n6884, n6885, n6886,
    n6887, n6888, n6889, n6890, n6891, n6892,
    n6893, n6894, n6895, n6896, n6897, n6898,
    n6899, n6900, n6901, n6902, n6903, n6904,
    n6905, n6906, n6907, n6908, n6909, n6910,
    n6911, n6912, n6913, n6914, n6915, n6916,
    n6917, n6918, n6919, n6920, n6921, n6922,
    n6923, n6924, n6925, n6926, n6927, n6928,
    n6929, n6930, n6931, n6932, n6933, n6934,
    n6935, n6936, n6937, n6938, n6939, n6940,
    n6941, n6942, n6943, n6944, n6945, n6946,
    n6947, n6948, n6949, n6950, n6951, n6952,
    n6953, n6955, n6956, n6957, n6958, n6959,
    n6960, n6961, n6962, n6963, n6964, n6965,
    n6966, n6967, n6968, n6969, n6970, n6971,
    n6972, n6973, n6974, n6975, n6976, n6977,
    n6978, n6979, n6980, n6981, n6982, n6983,
    n6984, n6985, n6986, n6987, n6988, n6989,
    n6990, n6991, n6992, n6993, n6994, n6995,
    n6996, n6997, n6998, n6999, n7000, n7001,
    n7002, n7003, n7004, n7005, n7006, n7007,
    n7008, n7009, n7010, n7011, n7012, n7013,
    n7014, n7015, n7016, n7017, n7018, n7019,
    n7020, n7021, n7022, n7023, n7024, n7025,
    n7026, n7027, n7028, n7029, n7030, n7031,
    n7032, n7033, n7034, n7035, n7036, n7037,
    n7038, n7039, n7040, n7041, n7042, n7043,
    n7044, n7046, n7047, n7048, n7049, n7050,
    n7051, n7052, n7053, n7054, n7055, n7056,
    n7057, n7058, n7059, n7060, n7061, n7062,
    n7063, n7064, n7065, n7066, n7067, n7068,
    n7069, n7070, n7071, n7072, n7073, n7074,
    n7075, n7076, n7077, n7078, n7079, n7080,
    n7081, n7082, n7083, n7084, n7085, n7086,
    n7087, n7088, n7089, n7090, n7091, n7092,
    n7093, n7094, n7095, n7096, n7097, n7098,
    n7099, n7100, n7101, n7102, n7103, n7104,
    n7105, n7106, n7107, n7108, n7109, n7110,
    n7111, n7112, n7113, n7114, n7115, n7116,
    n7117, n7118, n7119, n7120, n7121, n7122,
    n7123, n7124, n7125, n7126, n7127, n7128,
    n7129, n7130, n7131, n7132, n7133, n7134,
    n7135, n7137, n7138, n7139, n7140, n7141,
    n7142, n7143, n7144, n7145, n7146, n7147,
    n7148, n7149, n7150, n7151, n7152, n7153,
    n7154, n7155, n7156, n7157, n7158, n7159,
    n7160, n7161, n7162, n7163, n7164, n7165,
    n7166, n7167, n7168, n7169, n7170, n7171,
    n7172, n7173, n7174, n7175, n7176, n7177,
    n7178, n7179, n7180, n7181, n7182, n7183,
    n7184, n7185, n7186, n7187, n7188, n7189,
    n7190, n7191, n7192, n7193, n7194, n7195,
    n7196, n7197, n7198, n7199, n7200, n7201,
    n7202, n7203, n7204, n7205, n7206, n7207,
    n7208, n7209, n7210, n7211, n7212, n7213,
    n7214, n7215, n7216, n7217, n7218, n7219,
    n7220, n7221, n7222, n7223, n7224, n7225,
    n7226, n7228, n7229, n7230, n7231, n7232,
    n7233, n7234, n7235, n7236, n7237, n7238,
    n7239, n7240, n7241, n7242, n7243, n7244,
    n7245, n7246, n7247, n7248, n7249, n7250,
    n7251, n7252, n7253, n7254, n7255, n7256,
    n7257, n7258, n7259, n7260, n7261, n7262,
    n7263, n7264, n7265, n7266, n7267, n7268,
    n7269, n7270, n7271, n7272, n7273, n7274,
    n7275, n7276, n7277, n7278, n7279, n7280,
    n7281, n7283, n7284, n7286, n7287, n7288,
    n7289, n7290, n7291, n7292, n7293, n7294,
    n7295, n7296, n7297, n7298, n7299, n7300,
    n7301, n7302, n7303, n7304, n7305, n7306,
    n7307, n7308, n7309, n7310, n7311, n7312,
    n7313, n7314, n7315, n7316, n7317, n7318,
    n7319, n7320, n7321, n7322, n7323, n7324,
    n7325, n7326, n7327, n7328, n7329, n7330,
    n7331, n7332, n7333, n7334, n7335, n7337,
    n7338, n7339, n7340, n7342, n7344, n7346,
    n7348, n7349, n7350, n7351, n7352, n7353,
    n7354, n7355, n7356, n7358, n7359, n7360,
    n7361, n7362, n7363, n7364, n7365, n7366,
    n7367, n7368, n7369, n7370, n7371, n7372,
    n7373, n7374, n7375, n7376, n7377, n7378,
    n7379, n7380, n7381, n7382, n7383, n7384,
    n7385, n7386, n7387, n7388, n7389, n7390,
    n7391, n7392, n7393, n7394, n7395, n7396,
    n7397, n7398, n7399, n7400, n7401, n7402,
    n7403, n7404, n7405, n7406, n7407, n7408,
    n7409, n7410, n7411, n7412, n7413, n7414,
    n7415, n7416, n7417, n7418, n7419, n7420,
    n7421, n7422, n7423, n7424, n7425, n7426,
    n7427, n7428, n7429, n7430, n7431, n7432,
    n7433, n7434, n7435, n7436, n7437, n7438,
    n7439, n7440, n7441, n7442, n7443, n7444,
    n7445, n7446, n7447, n7448, n7449, n7450,
    n7451, n7452, n7453, n7454, n7455, n7456,
    n7457, n7458, n7459, n7460, n7461, n7462,
    n7463, n7464, n7465, n7466, n7467, n7468,
    n7469, n7470, n7471, n7472, n7473, n7474,
    n7475, n7476, n7477, n7478, n7479, n7480,
    n7481, n7482, n7483, n7484, n7485, n7486,
    n7487, n7488, n7489, n7490, n7491, n7492,
    n7493, n7494, n7495, n7496, n7497, n7498,
    n7499, n7500, n7501, n7502, n7503, n7504,
    n7505, n7506, n7507, n7508, n7509, n7510,
    n7511, n7512, n7513, n7514, n7515, n7516,
    n7517, n7518, n7519, n7520, n7521, n7522,
    n7523, n7524, n7525, n7526, n7527, n7528,
    n7529, n7530, n7531, n7532, n7533, n7534,
    n7535, n7536, n7537, n7538, n7539, n7540,
    n7541, n7542, n7543, n7544, n7545, n7546,
    n7547, n7548, n7549, n7550, n7551, n7552,
    n7553, n7554, n7555, n7556, n7557, n7558,
    n7559, n7560, n7561, n7562, n7563, n7564,
    n7565, n7566, n7567, n7568, n7569, n7570,
    n7571, n7572, n7573, n7574, n7575, n7576,
    n7577, n7578, n7579, n7580, n7581, n7582,
    n7583, n7584, n7585, n7586, n7587, n7588,
    n7589, n7590, n7591, n7592, n7593, n7594,
    n7595, n7596, n7597, n7598, n7599, n7600,
    n7601, n7602, n7603, n7604, n7605, n7606,
    n7607, n7608, n7609, n7610, n7611, n7612,
    n7613, n7614, n7615, n7616, n7617, n7618,
    n7619, n7620, n7621, n7622, n7623, n7624,
    n7625, n7626, n7627, n7628, n7629, n7630,
    n7631, n7632, n7633, n7634, n7635, n7636,
    n7637, n7638, n7639, n7640, n7641, n7642,
    n7643, n7644, n7645, n7646, n7647, n7648,
    n7649, n7650, n7651, n7652, n7653, n7654,
    n7655, n7656, n7657, n7658, n7659, n7660,
    n7661, n7662, n7663, n7664, n7665, n7666,
    n7667, n7668, n7669, n7670, n7671, n7672,
    n7673, n7674, n7675, n7676, n7677, n7678,
    n7679, n7680, n7681, n7682, n7683, n7684,
    n7685, n7686, n7687, n7688, n7689, n7690,
    n7691, n7692, n7693, n7694, n7695, n7696,
    n7697, n7698, n7699, n7700, n7701, n7702,
    n7703, n7704, n7705, n7706, n7707, n7708,
    n7709, n7710, n7711, n7712, n7713, n7714,
    n7715, n7716, n7717, n7718, n7719, n7720,
    n7721, n7722, n7723, n7724, n7725, n7726,
    n7727, n7728, n7729, n7730, n7731, n7732,
    n7733, n7734, n7735, n7736, n7737, n7738,
    n7739, n7740, n7741, n7742, n7743, n7744,
    n7745, n7746, n7747, n7748, n7749, n7750,
    n7751, n7752, n7753, n7754, n7755, n7756,
    n7757, n7758, n7759, n7760, n7761, n7762,
    n7763, n7764, n7765, n7766, n7767, n7768,
    n7769, n7770, n7771, n7772, n7773, n7774,
    n7775, n7776, n7777, n7778, n7779, n7780,
    n7781, n7782, n7783, n7784, n7785, n7786,
    n7787, n7788, n7789, n7790, n7791, n7792,
    n7793, n7794, n7795, n7796, n7797, n7798,
    n7799, n7800, n7801, n7802, n7803, n7804,
    n7805, n7806, n7807, n7808, n7809, n7810,
    n7811, n7812, n7813, n7814, n7815, n7816,
    n7817, n7818, n7819, n7820, n7821, n7822,
    n7823, n7824, n7825, n7826, n7827, n7828,
    n7829, n7830, n7831, n7832, n7833, n7834,
    n7835, n7836, n7837, n7838, n7839, n7840,
    n7841, n7842, n7843, n7844, n7845, n7846,
    n7847, n7848, n7849, n7850, n7851, n7852,
    n7853, n7854, n7855, n7856, n7857, n7858,
    n7859, n7860, n7861, n7862, n7863, n7864,
    n7865, n7866, n7867, n7868, n7869, n7870,
    n7871, n7872, n7873, n7874, n7875, n7876,
    n7877, n7878, n7879, n7880, n7881, n7882,
    n7883, n7884, n7885, n7886, n7887, n7888,
    n7889, n7890, n7891, n7892, n7893, n7894,
    n7895, n7896, n7897, n7898, n7899, n7900,
    n7901, n7902, n7903, n7904, n7905, n7906,
    n7907, n7908, n7909, n7910, n7911, n7912,
    n7913, n7914, n7915, n7916, n7917, n7918,
    n7919, n7920, n7921, n7922, n7923, n7924,
    n7925, n7926, n7927, n7928, n7929, n7930,
    n7931, n7932, n7933, n7934, n7935, n7936,
    n7937, n7938, n7939, n7940, n7941, n7942,
    n7943, n7944, n7945, n7946, n7947, n7948,
    n7949, n7950, n7951, n7952, n7953, n7954,
    n7955, n7956, n7957, n7958, n7959, n7960,
    n7961, n7962, n7963, n7964, n7965, n7966,
    n7967, n7968, n7969, n7970, n7971, n7972,
    n7973, n7974, n7975, n7976, n7977, n7978,
    n7979, n7980, n7981, n7982, n7983, n7984,
    n7985, n7986, n7987, n7988, n7989, n7990,
    n7991, n7992, n7993, n7994, n7995, n7996,
    n7997, n7998, n7999, n8000, n8001, n8002,
    n8003, n8004, n8005, n8006, n8007, n8008,
    n8009, n8010, n8011, n8012, n8013, n8014,
    n8015, n8016, n8017, n8018, n8019, n8020,
    n8021, n8022, n8023, n8024, n8025, n8026,
    n8027, n8028, n8029, n8030, n8031, n8032,
    n8033, n8034, n8035, n8036, n8037, n8038,
    n8039, n8040, n8041, n8042, n8043, n8044,
    n8045, n8046, n8047, n8048, n8049, n8050,
    n8051, n8052, n8053, n8054, n8055, n8056,
    n8057, n8058, n8059, n8060, n8061, n8062,
    n8063, n8064, n8065, n8066, n8067, n8068,
    n8069, n8070, n8071, n8072, n8073, n8074,
    n8075, n8076, n8077, n8078, n8079, n8080,
    n8081, n8082, n8083, n8084, n8085, n8086,
    n8087, n8088, n8089, n8090, n8091, n8092,
    n8093, n8094, n8095, n8096, n8097, n8098,
    n8099, n8100, n8101, n8102, n8103, n8104,
    n8105, n8106, n8107, n8108, n8109, n8110,
    n8111, n8112, n8113, n8114, n8115, n8116,
    n8117, n8118, n8119, n8120, n8121, n8122,
    n8123, n8124, n8125, n8126, n8127, n8128,
    n8129, n8130, n8131, n8132, n8133, n8134,
    n8135, n8136, n8137, n8138, n8139, n8140,
    n8141, n8142, n8143, n8144, n8145, n8146,
    n8147, n8148, n8149, n8150, n8151, n8152,
    n8153, n8154, n8155, n8156, n8157, n8158,
    n8159, n8160, n8161, n8162, n8163, n8164,
    n8165, n8166, n8167, n8168, n8169, n8170,
    n8171, n8172, n8173, n8174, n8175, n8176,
    n8177, n8178, n8179, n8180, n8181, n8182,
    n8183, n8184, n8185, n8186, n8187, n8188,
    n8189, n8190, n8191, n8192, n8193, n8194,
    n8195, n8196, n8197, n8198, n8199, n8200,
    n8201, n8202, n8203, n8204, n8205, n8206,
    n8207, n8208, n8209, n8210, n8211, n8212,
    n8213, n8214, n8215, n8216, n8217, n8218,
    n8219, n8220, n8221, n8222, n8223, n8224,
    n8225, n8226, n8227, n8228, n8229, n8230,
    n8231, n8232, n8233, n8234, n8235, n8236,
    n8237, n8238, n8239, n8240, n8241, n8242,
    n8243, n8244, n8245, n8246, n8247, n8248,
    n8249, n8250, n8251, n8252, n8253, n8254,
    n8255, n8256, n8257, n8258, n8259, n8260,
    n8261, n8262, n8263, n8264, n8265, n8266,
    n8267, n8268, n8269, n8270, n8271, n8272,
    n8273, n8274, n8275, n8276, n8277, n8278,
    n8279, n8280, n8281, n8282, n8283, n8284,
    n8285, n8286, n8287, n8288, n8289, n8290,
    n8291, n8292, n8293, n8294, n8295, n8296,
    n8297, n8298, n8299, n8300, n8301, n8302,
    n8303, n8304, n8305, n8306, n8307, n8308,
    n8309, n8310, n8311, n8312, n8313, n8314,
    n8315, n8316, n8317, n8318, n8319, n8320,
    n8321, n8322, n8323, n8324, n8325, n8326,
    n8327, n8328, n8329, n8330, n8331, n8332,
    n8333, n8334, n8335, n8336, n8337, n8338,
    n8339, n8340, n8341, n8342, n8343, n8344,
    n8345, n8346, n8347, n8348, n8349, n8350,
    n8351, n8352, n8353, n8354, n8355, n8356,
    n8357, n8358, n8359, n8360, n8361, n8362,
    n8363, n8364, n8365, n8366, n8367, n8368,
    n8369, n8370, n8371, n8372, n8373, n8374,
    n8375, n8376, n8377, n8378, n8379, n8380,
    n8381, n8382, n8383, n8384, n8385, n8386,
    n8387, n8388, n8389, n8390, n8391, n8392,
    n8393, n8394, n8395, n8396, n8397, n8398,
    n8399, n8400, n8401, n8402, n8403, n8404,
    n8405, n8406, n8407, n8408, n8409, n8410,
    n8411, n8412, n8413, n8414, n8415, n8416,
    n8417, n8418, n8419, n8420, n8421, n8422,
    n8423, n8424, n8425, n8426, n8427, n8428,
    n8429, n8430, n8431, n8432, n8433, n8434,
    n8435, n8436, n8437, n8438, n8439, n8440,
    n8441, n8442, n8443, n8444, n8445, n8446,
    n8447, n8448, n8449, n8450, n8451, n8452,
    n8453, n8454, n8455, n8456, n8457, n8458,
    n8459, n8460, n8461, n8462, n8463, n8464,
    n8465, n8466, n8467, n8468, n8469, n8470,
    n8471, n8472, n8473, n8474, n8475, n8476,
    n8477, n8478, n8479, n8480, n8481, n8482,
    n8483, n8484, n8485, n8486, n8487, n8488,
    n8489, n8490, n8491, n8492, n8493, n8494,
    n8495, n8496, n8497, n8498, n8499, n8500,
    n8501, n8502, n8503, n8504, n8505, n8506,
    n8507, n8508, n8509, n8510, n8511, n8512,
    n8513, n8514, n8515, n8516, n8517, n8518,
    n8519, n8520, n8521, n8522, n8523, n8524,
    n8525, n8526, n8527, n8528, n8529, n8530,
    n8531, n8532, n8533, n8534, n8535, n8536,
    n8537, n8538, n8539, n8540, n8541, n8542,
    n8543, n8544, n8545, n8546, n8547, n8548,
    n8549, n8550, n8551, n8552, n8553, n8554,
    n8555, n8556, n8557, n8558, n8559, n8560,
    n8561, n8562, n8563, n8564, n8565, n8566,
    n8567, n8568, n8569, n8570, n8571, n8572,
    n8573, n8574, n8575, n8576, n8577, n8578,
    n8579, n8580, n8581, n8582, n8583, n8584,
    n8585, n8586, n8587, n8588, n8589, n8590,
    n8591, n8592, n8593, n8594, n8595, n8597,
    n8598, n8599, n8600, n8601, n8602, n8603,
    n8604, n8605, n8606, n8607, n8608, n8609,
    n8610, n8611, n8612, n8613, n8614, n8615,
    n8616, n8617, n8618, n8620, n8621, n8622,
    n8623, n8624, n8625, n8626, n8627, n8628,
    n8629, n8630, n8631, n8632, n8633, n8634,
    n8635, n8636, n8637, n8638, n8639, n8640,
    n8641, n8642, n8643, n8644, n8645, n8646,
    n8647, n8648, n8649, n8650, n8651, n8652,
    n8653, n8654, n8655, n8656, n8657, n8658,
    n8659, n8660, n8661, n8662, n8663, n8664,
    n8665, n8666, n8667, n8668, n8669, n8670,
    n8671, n8672, n8673, n8674, n8675, n8676,
    n8677, n8679, n8680, n8681, n8682, n8683,
    n8684, n8685, n8686, n8687, n8688, n8689,
    n8690, n8691, n8692, n8693, n8694, n8695,
    n8696, n8697, n8698, n8699, n8700, n8701,
    n8702, n8703, n8704, n8705, n8706, n8707,
    n8708, n8709, n8710, n8711, n8712, n8713,
    n8714, n8715, n8716, n8717, n8718, n8719,
    n8720, n8721, n8722, n8723, n8724, n8725,
    n8726, n8727, n8728, n8729, n8730, n8731,
    n8732, n8733, n8734, n8735, n8736, n8737,
    n8738, n8739, n8740, n8741, n8742, n8743,
    n8744, n8745, n8746, n8747, n8748, n8749,
    n8750, n8751, n8752, n8753, n8754, n8755,
    n8756, n8757, n8758, n8759, n8760, n8761,
    n8762, n8763, n8764, n8765, n8766, n8767,
    n8768, n8769, n8770, n8771, n8772, n8773,
    n8774, n8775, n8776, n8777, n8778, n8779,
    n8780, n8781, n8782, n8783, n8784, n8785,
    n8786, n8787, n8788, n8789, n8790, n8791,
    n8792, n8793, n8794, n8795, n8796, n8797,
    n8798, n8799, n8800, n8801, n8802, n8803,
    n8804, n8805, n8806, n8807, n8808, n8809,
    n8810, n8811, n8812, n8813, n8814, n8815,
    n8816, n8817, n8818, n8819, n8820, n8821,
    n8822, n8823, n8824, n8825, n8826, n8827,
    n8828, n8829, n8830, n8831, n8832, n8833,
    n8834, n8835, n8836, n8837, n8838, n8839,
    n8840, n8841, n8842, n8843, n8844, n8845,
    n8846, n8847, n8848, n8849, n8850, n8851,
    n8852, n8853, n8854, n8855, n8856, n8857,
    n8858, n8859, n8860, n8861, n8862, n8863,
    n8864, n8865, n8866, n8867, n8868, n8869,
    n8870, n8871, n8872, n8873, n8874, n8875,
    n8876, n8877, n8878, n8879, n8880, n8881,
    n8882, n8883, n8884, n8885, n8886, n8887,
    n8888, n8889, n8890, n8891, n8892, n8893,
    n8894, n8895, n8896, n8897, n8898, n8899,
    n8900, n8901, n8902, n8903, n8904, n8905,
    n8906, n8907, n8908, n8909, n8910, n8911,
    n8912, n8913, n8914, n8915, n8916, n8917,
    n8918, n8919, n8920, n8921, n8922, n8923,
    n8924, n8925, n8926, n8927, n8928, n8929,
    n8930, n8931, n8932, n8933, n8934, n8935,
    n8936, n8937, n8938, n8939, n8940, n8941,
    n8942, n8943, n8944, n8945, n8946, n8947,
    n8948, n8949, n8950, n8951, n8952, n8953,
    n8954, n8955, n8956, n8957, n8958, n8959,
    n8960, n8961, n8962, n8963, n8964, n8965,
    n8966, n8967, n8968, n8969, n8970, n8971,
    n8972, n8973, n8974, n8975, n8976, n8977,
    n8978, n8979, n8980, n8981, n8982, n8983,
    n8984, n8985, n8986, n8987, n8988, n8989,
    n8990, n8991, n8992, n8993, n8994, n8995,
    n8996, n8997, n8998, n8999, n9000, n9001,
    n9002, n9003, n9004, n9005, n9006, n9007,
    n9008, n9009, n9010, n9011, n9012, n9013,
    n9014, n9015, n9016, n9017, n9018, n9019,
    n9020, n9021, n9022, n9023, n9024, n9025,
    n9026, n9027, n9028, n9029, n9030, n9031,
    n9032, n9033, n9034, n9035, n9036, n9037,
    n9038, n9039, n9040, n9041, n9042, n9043,
    n9044, n9045, n9046, n9047, n9048, n9049,
    n9050, n9051, n9052, n9053, n9054, n9055,
    n9056, n9057, n9058, n9059, n9060, n9061,
    n9062, n9063, n9064, n9065, n9066, n9067,
    n9068, n9069, n9070, n9071, n9072, n9073,
    n9074, n9075, n9076, n9077, n9078, n9079,
    n9080, n9081, n9082, n9083, n9084, n9085,
    n9086, n9087, n9088, n9089, n9090, n9091,
    n9092, n9093, n9094, n9095, n9096, n9097,
    n9098, n9099, n9100, n9101, n9102, n9103,
    n9104, n9105, n9106, n9107, n9108, n9109,
    n9110, n9111, n9112, n9113, n9114, n9115,
    n9116, n9117, n9118, n9119, n9120, n9121,
    n9122, n9123, n9124, n9125, n9126, n9127,
    n9128, n9129, n9130, n9131, n9132, n9133,
    n9134, n9135, n9136, n9137, n9138, n9139,
    n9140, n9141, n9142, n9143, n9144, n9145,
    n9146, n9147, n9148, n9149, n9150, n9151,
    n9152, n9153, n9154, n9155, n9156, n9157,
    n9158, n9159, n9160, n9161, n9162, n9163,
    n9164, n9165, n9166, n9167, n9168, n9169,
    n9170, n9171, n9172, n9173, n9174, n9175,
    n9176, n9177, n9178, n9179, n9180, n9181,
    n9182, n9183, n9184, n9185, n9186, n9187,
    n9188, n9189, n9190, n9191, n9192, n9193,
    n9194, n9195, n9196, n9197, n9198, n9199,
    n9200, n9201, n9202, n9203, n9204, n9205,
    n9206, n9207, n9208, n9209, n9210, n9211,
    n9212, n9213, n9214, n9215, n9216, n9217,
    n9218, n9219, n9220, n9221, n9222, n9223,
    n9224, n9225, n9226, n9227, n9228, n9229,
    n9230, n9231, n9232, n9233, n9234, n9235,
    n9236, n9237, n9238, n9239, n9240, n9241,
    n9242, n9243, n9244, n9245, n9246, n9247,
    n9248, n9249, n9250, n9251, n9252, n9253,
    n9254, n9255, n9256, n9257, n9258, n9259,
    n9260, n9261, n9262, n9263, n9264, n9265,
    n9266, n9267, n9268, n9269, n9270, n9271,
    n9272, n9273, n9274, n9275, n9276, n9277,
    n9278, n9279, n9280, n9281, n9282, n9283,
    n9284, n9285, n9286, n9287, n9288, n9289,
    n9290, n9291, n9292, n9293, n9294, n9295,
    n9296, n9297, n9298, n9299, n9300, n9301,
    n9302, n9303, n9304, n9305, n9306, n9307,
    n9308, n9309, n9310, n9311, n9312, n9313,
    n9314, n9315, n9316, n9317, n9318, n9319,
    n9320, n9321, n9322, n9323, n9324, n9325,
    n9326, n9327, n9328, n9329, n9330, n9331,
    n9332, n9333, n9334, n9335, n9336, n9337,
    n9338, n9339, n9340, n9341, n9342, n9343,
    n9344, n9345, n9346, n9347, n9348, n9349,
    n9350, n9351, n9352, n9354, n9355, n9356,
    n9357, n9358, n9359, n9360, n9361, n9362,
    n9363, n9364, n9365, n9366, n9367, n9368,
    n9369, n9370, n9371, n9372, n9373, n9374,
    n9375, n9376, n9377, n9378, n9379, n9380,
    n9381, n9382, n9383, n9384, n9385, n9386,
    n9387, n9388, n9389, n9390, n9391, n9392,
    n9393, n9394, n9395, n9396, n9397, n9398,
    n9399, n9400, n9401, n9402, n9403, n9404,
    n9405, n9406, n9407, n9408, n9409, n9410,
    n9411, n9412, n9413, n9414, n9415, n9416,
    n9417, n9418, n9419, n9420, n9421, n9422,
    n9423, n9424, n9425, n9426, n9427, n9428,
    n9429, n9430, n9431, n9432, n9433, n9434,
    n9435, n9436, n9437, n9438, n9439, n9440,
    n9441, n9442, n9443, n9444, n9445, n9446,
    n9447, n9448, n9449, n9450, n9451, n9452,
    n9453, n9454, n9455, n9456, n9457, n9458,
    n9459, n9460, n9461, n9462, n9463, n9464,
    n9465, n9466, n9467, n9468, n9469, n9470,
    n9471, n9472, n9473, n9474, n9475, n9476,
    n9477, n9478, n9479, n9480, n9481, n9482,
    n9483, n9484, n9485, n9486, n9487, n9488,
    n9489, n9490, n9491, n9492, n9493, n9494,
    n9495, n9496, n9497, n9498, n9499, n9500,
    n9501, n9502, n9503, n9504, n9505, n9506,
    n9507, n9508, n9509, n9510, n9511, n9512,
    n9513, n9514, n9515, n9516, n9517, n9518,
    n9519, n9520, n9521, n9522, n9523, n9524,
    n9525, n9526, n9527, n9528, n9529, n9530,
    n9531, n9532, n9533, n9534, n9535, n9536,
    n9537, n9538, n9539, n9540, n9541, n9542,
    n9543, n9544, n9545, n9546, n9547, n9548,
    n9549, n9550, n9551, n9552, n9553, n9554,
    n9555, n9556, n9557, n9558, n9559, n9560,
    n9561, n9562, n9563, n9564, n9565, n9566,
    n9567, n9568, n9569, n9570, n9571, n9572,
    n9573, n9574, n9575, n9576, n9577, n9578,
    n9579, n9580, n9581, n9582, n9583, n9584,
    n9585, n9586, n9587, n9588, n9589, n9590,
    n9591, n9592, n9593, n9594, n9595, n9596,
    n9597, n9598, n9599, n9600, n9601, n9602,
    n9603, n9604, n9605, n9606, n9607, n9608,
    n9609, n9610, n9611, n9612, n9613, n9614,
    n9615, n9616, n9617, n9618, n9619, n9620,
    n9621, n9622, n9623, n9624, n9625, n9626,
    n9627, n9628, n9629, n9630, n9631, n9632,
    n9633, n9634, n9635, n9636, n9637, n9638,
    n9639, n9640, n9641, n9642, n9643, n9644,
    n9645, n9646, n9647, n9648, n9649, n9650,
    n9651, n9652, n9653, n9654, n9655, n9656,
    n9657, n9658, n9659, n9660, n9661, n9662,
    n9663, n9664, n9665, n9666, n9667, n9668,
    n9669, n9670, n9671, n9672, n9673, n9674,
    n9675, n9676, n9677, n9678, n9679, n9680,
    n9681, n9682, n9683, n9684, n9685, n9686,
    n9687, n9688, n9689, n9690, n9691, n9692,
    n9693, n9694, n9695, n9696, n9697, n9698,
    n9699, n9700, n9701, n9702, n9704, n9705,
    n9706, n9707, n9708, n9709, n9710, n9711,
    n9712, n9713, n9714, n9715, n9716, n9717,
    n9718, n9719, n9720, n9721, n9722, n9723,
    n9724, n9725, n9726, n9727, n9728, n9729,
    n9730, n9731, n9732, n9733, n9734, n9735,
    n9736, n9737, n9738, n9739, n9740, n9741,
    n9742, n9743, n9744, n9745, n9746, n9747,
    n9748, n9749, n9750, n9751, n9752, n9753,
    n9754, n9755, n9756, n9757, n9758, n9759,
    n9760, n9761, n9762, n9763, n9764, n9765,
    n9766, n9767, n9768, n9769, n9770, n9771,
    n9772, n9773, n9774, n9775, n9776, n9778,
    n9779, n9780, n9781, n9782, n9783, n9784,
    n9785, n9786, n9787, n9788, n9789, n9790,
    n9791, n9792, n9793, n9794, n9795, n9796,
    n9797, n9798, n9799, n9801, n9802, n9803,
    n9804, n9805, n9806, n9807, n9808, n9809,
    n9810, n9811, n9812, n9813, n9814, n9815,
    n9816, n9817, n9818, n9819, n9820, n9821,
    n9822, n9823, n9824, n9825, n9826, n9827,
    n9828, n9829, n9830, n9831, n9833, n9834,
    n9835, n9836, n9837, n9838, n9839, n9840,
    n9841, n9842, n9843, n9844, n9845, n9846,
    n9847, n9848, n9849, n9850, n9851, n9852,
    n9853, n9854, n9855, n9856, n9857, n9858,
    n9859, n9860, n9861, n9862, n9863, n9864,
    n9865, n9866, n9867, n9868, n9869, n9870,
    n9871, n9872, n9873, n9874, n9875, n9876,
    n9877, n9878, n9879, n9880, n9881, n9882,
    n9883, n9884, n9885, n9886, n9887, n9888,
    n9889, n9890, n9891, n9892, n9893, n9894,
    n9895, n9896, n9897, n9898, n9899, n9900,
    n9901, n9902, n9903, n9904, n9905, n9906,
    n9907, n9908, n9909, n9910, n9911, n9912,
    n9914, n9915, n9916, n9917, n9918, n9919,
    n9920, n9921, n9922, n9923, n9924, n9925,
    n9927, n9928, n9929, n9930, n9931, n9932,
    n9933, n9934, n9935, n9936, n9937, n9938,
    n9939, n9940, n9941, n9942, n9943, n9944,
    n9945, n9946, n9947, n9948, n9949, n9950,
    n9951, n9952, n9953, n9954, n9955, n9956,
    n9957, n9958, n9959, n9960, n9961, n9962,
    n9963, n9964, n9965, n9966, n9967, n9968,
    n9969, n9970, n9971, n9972, n9973, n9974,
    n9975, n9976, n9977, n9978, n9979, n9980,
    n9981, n9982, n9983, n9984, n9985, n9986,
    n9987, n9988, n9989, n9990, n9991, n9992,
    n9993, n9994, n9995, n9996, n9997, n9998,
    n9999, n10000, n10001, n10002, n10003, n10004,
    n10005, n10006, n10007, n10008, n10009, n10010,
    n10011, n10012, n10013, n10014, n10015, n10016,
    n10017, n10018, n10019, n10020, n10021, n10022,
    n10023, n10024, n10025, n10026, n10027, n10028,
    n10029, n10030, n10031, n10032, n10033, n10034,
    n10035, n10036, n10037, n10038, n10039, n10040,
    n10041, n10042, n10043, n10044, n10045, n10046,
    n10047, n10048, n10049, n10050, n10051, n10052,
    n10053, n10054, n10055, n10056, n10057, n10058,
    n10059, n10060, n10061, n10062, n10063, n10064,
    n10065, n10066, n10067, n10068, n10069, n10070,
    n10071, n10072, n10073, n10074, n10075, n10076,
    n10077, n10078, n10079, n10080, n10081, n10082,
    n10083, n10084, n10085, n10086, n10087, n10088,
    n10089, n10090, n10091, n10092, n10093, n10094,
    n10095, n10096, n10098, n10099, n10100, n10101,
    n10102, n10103, n10104, n10105, n10106, n10107,
    n10108, n10109, n10110, n10111, n10112, n10113,
    n10114, n10115, n10116, n10117, n10118, n10119,
    n10120, n10121, n10122, n10123, n10124, n10125,
    n10126, n10127, n10128, n10129, n10130, n10131,
    n10132, n10133, n10134, n10135, n10136, n10137,
    n10138, n10139, n10140, n10141, n10142, n10143,
    n10144, n10145, n10146, n10147, n10148, n10149,
    n10150, n10151, n10152, n10153, n10154, n10155,
    n10156, n10157, n10158, n10159, n10160, n10161,
    n10162, n10163, n10164, n10165, n10166, n10167,
    n10168, n10169, n10170, n10171, n10172, n10173,
    n10174, n10175, n10176, n10177, n10178, n10179,
    n10180, n10181, n10182, n10183, n10184, n10185,
    n10186, n10187, n10188, n10189, n10190, n10191,
    n10192, n10193, n10194, n10195, n10196, n10197,
    n10198, n10199, n10200, n10201, n10202, n10203,
    n10204, n10205, n10206, n10207, n10208, n10209,
    n10210, n10211, n10212, n10213, n10214, n10215,
    n10216, n10217, n10218, n10219, n10220, n10221,
    n10222, n10223, n10224, n10225, n10226, n10227,
    n10228, n10229, n10230, n10231, n10232, n10233,
    n10234, n10235, n10236, n10237, n10238, n10239,
    n10240, n10241, n10242, n10243, n10244, n10245,
    n10246, n10247, n10248, n10249, n10250, n10251,
    n10252, n10253, n10254, n10255, n10256, n10257,
    n10258, n10259, n10260, n10261, n10262, n10263,
    n10264, n10265, n10266, n10267, n10268, n10269,
    n10270, n10271, n10272, n10273, n10274, n10275,
    n10276, n10277, n10278, n10279, n10280, n10281,
    n10282, n10283, n10284, n10285, n10286, n10287,
    n10288, n10289, n10290, n10291, n10292, n10293,
    n10294, n10295, n10296, n10297, n10298, n10299,
    n10300, n10301, n10302, n10303, n10304, n10305,
    n10306, n10307, n10308, n10309, n10310, n10311,
    n10312, n10313, n10314, n10315, n10316, n10317,
    n10318, n10319, n10320, n10321, n10322, n10323,
    n10324, n10325, n10326, n10327, n10328, n10329,
    n10330, n10332, n10333, n10334, n10335, n10336,
    n10337, n10338, n10339, n10340, n10341, n10342,
    n10343, n10344, n10345, n10346, n10347, n10348,
    n10349, n10350, n10351, n10352, n10353, n10354,
    n10355, n10356, n10357, n10358, n10359, n10360,
    n10361, n10362, n10363, n10364, n10365, n10366,
    n10367, n10368, n10369, n10370, n10371, n10372,
    n10373, n10374, n10375, n10376, n10377, n10378,
    n10379, n10380, n10381, n10382, n10383, n10384,
    n10385, n10386, n10387, n10388, n10389, n10390,
    n10391, n10392, n10393, n10394, n10395, n10396,
    n10397, n10398, n10399, n10400, n10401, n10402,
    n10403, n10404, n10405, n10406, n10407, n10408,
    n10409, n10410, n10411, n10412, n10413, n10414,
    n10415, n10416, n10417, n10418, n10419, n10420,
    n10421, n10422, n10423, n10424, n10425, n10426,
    n10427, n10428, n10429, n10430, n10431, n10432,
    n10433, n10434, n10435, n10436, n10437, n10438,
    n10439, n10440, n10441, n10442, n10443, n10444,
    n10445, n10446, n10447, n10448, n10449, n10450,
    n10451, n10452, n10453, n10454, n10455, n10456,
    n10457, n10458, n10459, n10460, n10461, n10462,
    n10463, n10464, n10465, n10466, n10467, n10468,
    n10469, n10470, n10471, n10472, n10473, n10474,
    n10475, n10476, n10477, n10478, n10479, n10480,
    n10481, n10482, n10483, n10484, n10485, n10486,
    n10487, n10488, n10489, n10490, n10491, n10492,
    n10493, n10494, n10495, n10496, n10497, n10498,
    n10499, n10500, n10501, n10502, n10503, n10504,
    n10505, n10506, n10507, n10508, n10509, n10511,
    n10512, n10513, n10514, n10515, n10516, n10517,
    n10518, n10519, n10520, n10521, n10522, n10523,
    n10524, n10525, n10526, n10527, n10528, n10529,
    n10530, n10531, n10532, n10533, n10534, n10535,
    n10536, n10537, n10538, n10539, n10540, n10541,
    n10542, n10543, n10544, n10545, n10546, n10547,
    n10548, n10549, n10550, n10551, n10552, n10553,
    n10554, n10555, n10556, n10557, n10558, n10559,
    n10560, n10561, n10562, n10563, n10564, n10565,
    n10566, n10567, n10568, n10569, n10570, n10571,
    n10572, n10573, n10574, n10575, n10576, n10577,
    n10578, n10579, n10580, n10581, n10582, n10584,
    n10585, n10586, n10588, n10589, n10590, n10591,
    n10592, n10593, n10594, n10595, n10596, n10597,
    n10598, n10599, n10600, n10601, n10602, n10603,
    n10604, n10605, n10607, n10608, n10609, n10610,
    n10611, n10612, n10613, n10614, n10615, n10616,
    n10617, n10618, n10619, n10620, n10621, n10622,
    n10623, n10624, n10625, n10626, n10627, n10628,
    n10629, n10630, n10631, n10632, n10633, n10634,
    n10635, n10636, n10637, n10638, n10639, n10640,
    n10641, n10642, n10643, n10644, n10645, n10646,
    n10647, n10648, n10649, n10650, n10652, n10653,
    n10654, n10656, n10657, n10658, n10659, n10660,
    n10661, n10662, n10663, n10664, n10665, n10666,
    n10667, n10668, n10669, n10670, n10671, n10672,
    n10673, n10674, n10675, n10676, n10678, n10679,
    n10680, n10681, n10682, n10683, n10684, n10685,
    n10686, n10687, n10688, n10689, n10690, n10691,
    n10692, n10693, n10694, n10695, n10696, n10697,
    n10698, n10699, n10700, n10701, n10702, n10704,
    n10705, n10706, n10707, n10708, n10709, n10710,
    n10712, n10713, n10714, n10715, n10716, n10717,
    n10718, n10719, n10720, n10721, n10722, n10723,
    n10724, n10725, n10726, n10727, n10728, n10729,
    n10730, n10731, n10732, n10733, n10734, n10735,
    n10736, n10737, n10738, n10739, n10740, n10741,
    n10742, n10743, n10744, n10745, n10746, n10747,
    n10748, n10749, n10750, n10751, n10752, n10753,
    n10754, n10755, n10756, n10757, n10758, n10759,
    n10760, n10761, n10762, n10763, n10764, n10765,
    n10766, n10767, n10768, n10769, n10770, n10771,
    n10772, n10773, n10774, n10775, n10776, n10777,
    n10778, n10779, n10780, n10781, n10782, n10783,
    n10784, n10785, n10786, n10787, n10788, n10789,
    n10790, n10791, n10792, n10793, n10794, n10795,
    n10796, n10797, n10798, n10799, n10800, n10801,
    n10802, n10803, n10804, n10805, n10806, n10807,
    n10808, n10809, n10810, n10811, n10812, n10813,
    n10814, n10815, n10816, n10817, n10818, n10819,
    n10820, n10821, n10822, n10823, n10824, n10825,
    n10826, n10827, n10828, n10829, n10830, n10831,
    n10832, n10833, n10834, n10835, n10836, n10837,
    n10838, n10839, n10840, n10841, n10842, n10843,
    n10844, n10845, n10846, n10848, n10849, n10850,
    n10851, n10852, n10853, n10854, n10855, n10856,
    n10857, n10858, n10860, n10861, n10862, n10863,
    n10864, n10865, n10866, n10867, n10868, n10869,
    n10870, n10871, n10872, n10873, n10874, n10875,
    n10876, n10877, n10878, n10880, n10881, n10882,
    n10883, n10884, n10885, n10886, n10887, n10888,
    n10889, n10890, n10891, n10892, n10894, n10895,
    n10896, n10897, n10898, n10899, n10900, n10902,
    n10903, n10904, n10905, n10906, n10907, n10908,
    n10909, n10910, n10912, n10913, n10915, n10916,
    n10917, n10918, n10919, n10921, n10922, n10923,
    n10924, n10925, n10926, n10927, n10928, n10930,
    n10931, n10932, n10933, n10935, n10936, n10937,
    n10938, n10940, n10941, n10942, n10943, n10944,
    n10946, n10947, n10948, n10949, n10950, n10951,
    n10952, n10954, n10955, n10957, n10958, n10959,
    n10960, n10961, n10962, n10963, n10964, n10965,
    n10966, n10967, n10968, n10969, n10970, n10971,
    n10972, n10973, n10974, n10976, n10977, n10978,
    n10979, n10981, n10982, n10983, n10984, n10985,
    n10986, n10987, n10989, n10990, n10991, n10992,
    n10993, n10994, n10995, n10996, n10997, n10998,
    n10999, n11000, n11002, n11003, n11004, n11005,
    n11006, n11007, n11008, n11009, n11010, n11011,
    n11012, n11013, n11014, n11015, n11016, n11017,
    n11018, n11019, n11020, n11021, n11022, n11023,
    n11024, n11025, n11026, n11028, n11029, n11030,
    n11031, n11032, n11033, n11034, n11035, n11036,
    n11037, n11038, n11039, n11040, n11041, n11042,
    n11043, n11044, n11045, n11046, n11047, n11049,
    n11050, n11051, n11052, n11053, n11054, n11055,
    n11056, n11057, n11058, n11059, n11060, n11061,
    n11063, n11064, n11065, n11066, n11067, n11068,
    n11069, n11070, n11071, n11072, n11073, n11075,
    n11076, n11077, n11078, n11079, n11080, n11081,
    n11082, n11083, n11084, n11085, n11086, n11087,
    n11088, n11089, n11090, n11092, n11093, n11094,
    n11095, n11096, n11097, n11098, n11100, n11101,
    n11102, n11103, n11104, n11105, n11106, n11107,
    n11108, n11109, n11110, n11111, n11112, n11113,
    n11114, n11115, n11116, n11117, n11118, n11119,
    n11120, n11121, n11122, n11123, n11124, n11125,
    n11126, n11127, n11128, n11129, n11130, n11131,
    n11132, n11133, n11134, n11135, n11136, n11137,
    n11138, n11139, n11140, n11141, n11142, n11143,
    n11144, n11145, n11146, n11147, n11148, n11149,
    n11150, n11151, n11152, n11153, n11154, n11155,
    n11156, n11157, n11158, n11159, n11160, n11161,
    n11162, n11163, n11164, n11165, n11166, n11167,
    n11168, n11169, n11170, n11171, n11172, n11173,
    n11174, n11175, n11176, n11177, n11178, n11179,
    n11180, n11181, n11182, n11183, n11184, n11185,
    n11186, n11187, n11188, n11189, n11190, n11191,
    n11192, n11193, n11194, n11195, n11196, n11197,
    n11198, n11199, n11200, n11201, n11202, n11203,
    n11204, n11205, n11206, n11207, n11208, n11209,
    n11210, n11211, n11212, n11213, n11214, n11215,
    n11216, n11217, n11218, n11219, n11220, n11221,
    n11222, n11223, n11224, n11225, n11226, n11227,
    n11228, n11229, n11230, n11231, n11232, n11233,
    n11234, n11235, n11236, n11237, n11238, n11239,
    n11240, n11241, n11242, n11243, n11244, n11245,
    n11246, n11247, n11248, n11249, n11250, n11252,
    n11253, n11254, n11255, n11256, n11257, n11258,
    n11259, n11260, n11262, n11264, n11265, n11266,
    n11267, n11268, n11269, n11270, n11271, n11272,
    n11273, n11274, n11275, n11276, n11277, n11278,
    n11279, n11280, n11281, n11282, n11283, n11284,
    n11285, n11286, n11287, n11288, n11289, n11290,
    n11291, n11292, n11293, n11294, n11295, n11296,
    n11297, n11298, n11299, n11300, n11301, n11302,
    n11303, n11304, n11305, n11306, n11307, n11308,
    n11309, n11310, n11311, n11312, n11313, n11314,
    n11315, n11316, n11317, n11318, n11319, n11320,
    n11321, n11322, n11323, n11324, n11325, n11326,
    n11327, n11328, n11329, n11330, n11331, n11332,
    n11333, n11334, n11335, n11336, n11337, n11338,
    n11339, n11340, n11341, n11342, n11343, n11344,
    n11345, n11346, n11347, n11348, n11349, n11350,
    n11351, n11352, n11353, n11354, n11355, n11356,
    n11357, n11358, n11359, n11360, n11361, n11362,
    n11363, n11364, n11365, n11366, n11367, n11368,
    n11369, n11370, n11371, n11372, n11373, n11374,
    n11375, n11376, n11377, n11378, n11379, n11380,
    n11381, n11382, n11383, n11384, n11385, n11386,
    n11387, n11388, n11389, n11390, n11391, n11392,
    n11393, n11394, n11395, n11396, n11397, n11398,
    n11399, n11400, n11401, n11402, n11403, n11404,
    n11405, n11406, n11407, n11408, n11409, n11410,
    n11411, n11412, n11413, n11414, n11415, n11416,
    n11417, n11418, n11419, n11420, n11421, n11422,
    n11423, n11424, n11425, n11426, n11427, n11428,
    n11429, n11430, n11431, n11432, n11433, n11434,
    n11435, n11436, n11437, n11438, n11439, n11440,
    n11441, n11442, n11443, n11444, n11445, n11446,
    n11447, n11448, n11449, n11450, n11451, n11452,
    n11453, n11454, n11455, n11456, n11457, n11458,
    n11459, n11460, n11461, n11462, n11463, n11464,
    n11465, n11466, n11467, n11468, n11469, n11470,
    n11471, n11472, n11473, n11474, n11475, n11476,
    n11477, n11478, n11479, n11480, n11481, n11482,
    n11483, n11484, n11485, n11486, n11487, n11488,
    n11489, n11490, n11491, n11492, n11493, n11494,
    n11495, n11496, n11497, n11498, n11499, n11500,
    n11501, n11502, n11503, n11504, n11505, n11506,
    n11507, n11508, n11509, n11510, n11511, n11512,
    n11513, n11514, n11515, n11516, n11517, n11518,
    n11519, n11520, n11521, n11522, n11523, n11524,
    n11525, n11526, n11527, n11528, n11529, n11530,
    n11531, n11532, n11533, n11534, n11535, n11536,
    n11537, n11538, n11539, n11540, n11541, n11542,
    n11543, n11544, n11545, n11546, n11547, n11548,
    n11549, n11550, n11551, n11552, n11553, n11554,
    n11555, n11556, n11557, n11558, n11559, n11560,
    n11561, n11562, n11563, n11564, n11565, n11566,
    n11567, n11568, n11569, n11570, n11571, n11572,
    n11573, n11574, n11575, n11576, n11577, n11578,
    n11579, n11580, n11581, n11582, n11583, n11584,
    n11585, n11586, n11587, n11588, n11589, n11590,
    n11591, n11592, n11593, n11594, n11595, n11596,
    n11597, n11598, n11599, n11600, n11601, n11602,
    n11603, n11604, n11605, n11606, n11607, n11608,
    n11609, n11610, n11611, n11612, n11613, n11614,
    n11615, n11616, n11617, n11618, n11619, n11620,
    n11621, n11622, n11623, n11624, n11625, n11626,
    n11627, n11628, n11629, n11630, n11631, n11632,
    n11633, n11634, n11635, n11636, n11637, n11638,
    n11639, n11640, n11641, n11642, n11643, n11644,
    n11645, n11646, n11647, n11648, n11649, n11650,
    n11651, n11652, n11653, n11654, n11655, n11656,
    n11657, n11658, n11659, n11660, n11661, n11662,
    n11663, n11664, n11665, n11666, n11667, n11668,
    n11669, n11670, n11671, n11672, n11673, n11674,
    n11675, n11676, n11677, n11678, n11679, n11680,
    n11681, n11682, n11683, n11684, n11685, n11686,
    n11687, n11688, n11689, n11690, n11691, n11692,
    n11693, n11694, n11695, n11696, n11697, n11698,
    n11699, n11700, n11701, n11702, n11703, n11704,
    n11705, n11706, n11707, n11708, n11709, n11710,
    n11711, n11712, n11713, n11714, n11715, n11716,
    n11717, n11719, n11720, n11721, n11722, n11723,
    n11724, n11725, n11726, n11727, n11728, n11729,
    n11730, n11731, n11732, n11733, n11734, n11735,
    n11736, n11737, n11738, n11739, n11740, n11741,
    n11742, n11743, n11744, n11745, n11746, n11747,
    n11748, n11749, n11750, n11751, n11752, n11753,
    n11754, n11755, n11756, n11757, n11758, n11759,
    n11760, n11761, n11762, n11763, n11764, n11765,
    n11766, n11767, n11768, n11769, n11770, n11771,
    n11772, n11773, n11774, n11775, n11776, n11777,
    n11778, n11779, n11780, n11781, n11782, n11783,
    n11784, n11785, n11786, n11787, n11788, n11789,
    n11790, n11791, n11792, n11793, n11794, n11795,
    n11796, n11797, n11798, n11799, n11800, n11801,
    n11802, n11803, n11804, n11805, n11806, n11807,
    n11808, n11809, n11810, n11811, n11812, n11813,
    n11814, n11815, n11816, n11817, n11818, n11819,
    n11820, n11821, n11822, n11823, n11824, n11825,
    n11826, n11827, n11828, n11829, n11830, n11831,
    n11832, n11833, n11834, n11835, n11836, n11837,
    n11838, n11839, n11840, n11841, n11842, n11843,
    n11844, n11845, n11846, n11847, n11848, n11849,
    n11850, n11851, n11852, n11853, n11854, n11855,
    n11856, n11857, n11858, n11859, n11860, n11861,
    n11862, n11863, n11864, n11865, n11866, n11867,
    n11868, n11869, n11870, n11871, n11872, n11873,
    n11874, n11875, n11876, n11877, n11878, n11879,
    n11880, n11881, n11882, n11883, n11884, n11885,
    n11886, n11887, n11888, n11889, n11890, n11891,
    n11892, n11893, n11894, n11895, n11896, n11897,
    n11898, n11899, n11900, n11901, n11902, n11903,
    n11904, n11905, n11906, n11907, n11908, n11909,
    n11910, n11911, n11912, n11913, n11914, n11915,
    n11916, n11917, n11918, n11919, n11920, n11921,
    n11922, n11923, n11924, n11925, n11926, n11927,
    n11928, n11929, n11930, n11931, n11932, n11933,
    n11934, n11935, n11936, n11937, n11938, n11939,
    n11940, n11941, n11942, n11943, n11944, n11945,
    n11946, n11947, n11948, n11949, n11950, n11951,
    n11952, n11953, n11954, n11955, n11956, n11957,
    n11958, n11959, n11960, n11961, n11962, n11963,
    n11964, n11965, n11966, n11967, n11968, n11969,
    n11970, n11971, n11972, n11973, n11974, n11975,
    n11976, n11977, n11978, n11979, n11980, n11981,
    n11982, n11983, n11984, n11985, n11986, n11987,
    n11988, n11989, n11990, n11991, n11992, n11993,
    n11994, n11995, n11996, n11997, n11998, n11999,
    n12000, n12001, n12002, n12003, n12004, n12005,
    n12006, n12007, n12008, n12009, n12010, n12011,
    n12012, n12013, n12014, n12015, n12016, n12017,
    n12018, n12019, n12020, n12021, n12022, n12023,
    n12024, n12025, n12026, n12027, n12028, n12029,
    n12030, n12031, n12032, n12033, n12034, n12035,
    n12036, n12037, n12038, n12039, n12040, n12041,
    n12042, n12043, n12044, n12045, n12046, n12047,
    n12048, n12049, n12050, n12051, n12052, n12053,
    n12054, n12055, n12056, n12057, n12058, n12059,
    n12060, n12061, n12062, n12063, n12064, n12065,
    n12066, n12067, n12068, n12069, n12070, n12071,
    n12072, n12073, n12074, n12075, n12076, n12077,
    n12078, n12079, n12080, n12081, n12082, n12083,
    n12084, n12085, n12086, n12087, n12088, n12089,
    n12090, n12091, n12092, n12093, n12094, n12095,
    n12096, n12097, n12098, n12099, n12100, n12101,
    n12102, n12103, n12104, n12105, n12106, n12107,
    n12108, n12109, n12110, n12111, n12112, n12113,
    n12114, n12115, n12116, n12117, n12118, n12119,
    n12120, n12121, n12122, n12123, n12124, n12125,
    n12126, n12127, n12128, n12129, n12130, n12131,
    n12132, n12133, n12134, n12135, n12136, n12137,
    n12138, n12139, n12140, n12141, n12142, n12143,
    n12144, n12145, n12146, n12147, n12148, n12149,
    n12150, n12151, n12152, n12153, n12154, n12155,
    n12156, n12157, n12158, n12159, n12160, n12161,
    n12162, n12163, n12164, n12165, n12166, n12167,
    n12168, n12169, n12170, n12171, n12172, n12173,
    n12174, n12175, n12176, n12177, n12178, n12179,
    n12180, n12181, n12182, n12183, n12184, n12185,
    n12186, n12187, n12188, n12189, n12190, n12191,
    n12192, n12193, n12194, n12195, n12196, n12197,
    n12198, n12199, n12200, n12201, n12202, n12203,
    n12204, n12205, n12206, n12207, n12208, n12209,
    n12210, n12211, n12212, n12213, n12214, n12215,
    n12216, n12217, n12218, n12219, n12220, n12221,
    n12222, n12223, n12224, n12225, n12226, n12227,
    n12228, n12229, n12230, n12231, n12232, n12233,
    n12234, n12235, n12236, n12237, n12238, n12239,
    n12240, n12241, n12242, n12243, n12244, n12245,
    n12246, n12247, n12248, n12249, n12250, n12251,
    n12252, n12253, n12254, n12255, n12256, n12257,
    n12258, n12259, n12260, n12261, n12262, n12263,
    n12264, n12265, n12266, n12267, n12268, n12269,
    n12270, n12271, n12272, n12273, n12274, n12275,
    n12276, n12277, n12278, n12279, n12280, n12281,
    n12282, n12283, n12284, n12285, n12286, n12287,
    n12288, n12289, n12290, n12291, n12292, n12293,
    n12294, n12295, n12296, n12297, n12298, n12299,
    n12300, n12301, n12302, n12303, n12304, n12305,
    n12306, n12308, n12309, n12310, n12311, n12312,
    n12313, n12314, n12315, n12316, n12318, n12319,
    n12320, n12321, n12322, n12323, n12324, n12325,
    n12327, n12328, n12329, n12330, n12331, n12332,
    n12333, n12334, n12335, n12336, n12337, n12338,
    n12339, n12341, n12342, n12343, n12344, n12345,
    n12347, n12348, n12349, n12350, n12352, n12353,
    n12354, n12356, n12357, n12358, n12359, n12361,
    n12362, n12363, n12364, n12365, n12366, n12367,
    n12368, n12369, n12370, n12371, n12372, n12373,
    n12374, n12375, n12376, n12377, n12379, n12380,
    n12381, n12382, n12383, n12384, n12385, n12387,
    n12388, n12389, n12390, n12392, n12393, n12394,
    n12395, n12396, n12397, n12398, n12399, n12400,
    n12401, n12403, n12404, n12405, n12406, n12407,
    n12408, n12409, n12410, n12411, n12412, n12413,
    n12414, n12416, n12417, n12418, n12419, n12420,
    n12421, n12422, n12424, n12425, n12426, n12427,
    n12428, n12429, n12430, n12431, n12432, n12433,
    n12434, n12435, n12436, n12437, n12438, n12439,
    n12440, n12442, n12443, n12444, n12445, n12446,
    n12447, n12448, n12449, n12450, n12452, n12453,
    n12454, n12455, n12456, n12457, n12458, n12459,
    n12460, n12461, n12462, n12463, n12465, n12466,
    n12467, n12468, n12469, n12470, n12471, n12472,
    n12473, n12474, n12476, n12477, n12478, n12479,
    n12481, n12482, n12483, n12484, n12485, n12486,
    n12487, n12488, n12489, n12490, n12491, n12492,
    n12493, n12494, n12495, n12496, n12497, n12498,
    n12499, n12500, n12501, n12502, n12503, n12504,
    n12505, n12506, n12507, n12508, n12509, n12510,
    n12511, n12512, n12513, n12514, n12515, n12516,
    n12517, n12518, n12519, n12520, n12521, n12522,
    n12523, n12524, n12525, n12526, n12527, n12528,
    n12529, n12530, n12531, n12532, n12533, n12534,
    n12535, n12536, n12537, n12538, n12539, n12540,
    n12541, n12542, n12543, n12544, n12545, n12546,
    n12547, n12548, n12549, n12550, n12551, n12552,
    n12553, n12554, n12555, n12557, n12558, n12559,
    n12560, n12561, n12562, n12563, n12564, n12565,
    n12566, n12568, n12569, n12570, n12571, n12572,
    n12573, n12574, n12575, n12576, n12577, n12578,
    n12579, n12580, n12581, n12582, n12583, n12584,
    n12585, n12586, n12587, n12588, n12589, n12590,
    n12591, n12592, n12593, n12594, n12595, n12596,
    n12597, n12598, n12599, n12600, n12601, n12602,
    n12603, n12604, n12605, n12606, n12607, n12608,
    n12609, n12610, n12611, n12612, n12613, n12614,
    n12615, n12616, n12617, n12618, n12619, n12620,
    n12621, n12622, n12623, n12624, n12625, n12626,
    n12627, n12628, n12629, n12630, n12631, n12632,
    n12633, n12634, n12635, n12636, n12637, n12638,
    n12639, n12640, n12641, n12642, n12643, n12645,
    n12647, n12648, n12649, n12650, n12651, n12652,
    n12653, n12655, n12656, n12657, n12658, n12659,
    n12660, n12661, n12662, n12663, n12664, n12665,
    n12666, n12668, n12669, n12670, n12671, n12672,
    n12673, n12674, n12675, n12676, n12678, n12680,
    n12681, n12682, n12683, n12684, n12685, n12686,
    n12687, n12688, n12689, n12690, n12691, n12692,
    n12693, n12694, n12695, n12696, n12698, n12700,
    n12701, n12702, n12703, n12704, n12705, n12706,
    n12707, n12709, n12710, n12711, n12712, n12713,
    n12716, n12717, n12718, n12719, n12720, n12721,
    n12722, n12723, n12724, n12725, n12726, n12727,
    n12728, n12729, n12730, n12731, n12732, n12733,
    n12734, n12735, n12736, n12737, n12738, n12739,
    n12740, n12741, n12742, n12743, n12744, n12745,
    n12746, n12747, n12748, n12749, n12750, n12751,
    n12752, n12753, n12754, n12755, n12756, n12757,
    n12758, n12759, n12760, n12761, n12762, n12764,
    n12765, n12766, n12767, n12768, n12769, n12770,
    n12771, n12772, n12773, n12774, n12775, n12776,
    n12777, n12778, n12779, n12780, n12781, n12782,
    n12783, n12784, n12785, n12786, n12787, n12788,
    n12789, n12790, n12791, n12792, n12793, n12794,
    n12795, n12796, n12797, n12798, n12799, n12800,
    n12801, n12802, n12803, n12804, n12805, n12806,
    n12807, n12808, n12809, n12811, n12812, n12813,
    n12814, n12815, n12816, n12817, n12818, n12819,
    n12820, n12821, n12822, n12823, n12824, n12825,
    n12826, n12827, n12828, n12829, n12830, n12831,
    n12832, n12833, n12834, n12835, n12836, n12837,
    n12838, n12839, n12840, n12841, n12842, n12843,
    n12844, n12845, n12846, n12847, n12848, n12849,
    n12850, n12851, n12853, n12854, n12855, n12856,
    n12857, n12858, n12859, n12860, n12861, n12862,
    n12863, n12864, n12865, n12866, n12867, n12868,
    n12869, n12870, n12871, n12872, n12873, n12874,
    n12875, n12876, n12877, n12878, n12879, n12880,
    n12881, n12882, n12883, n12884, n12885, n12886,
    n12887, n12888, n12889, n12890, n12891, n12892,
    n12893, n12894, n12895, n12896, n12897, n12898,
    n12899, n12900, n12901, n12903, n12904, n12905,
    n12906, n12907, n12908, n12909, n12910, n12911,
    n12912, n12913, n12914, n12915, n12916, n12917,
    n12919, n12920, n12921, n12922, n12923, n12924,
    n12925, n12926, n12927, n12928, n12929, n12930,
    n12931, n12932, n12933, n12934, n12935, n12936,
    n12937, n12938, n12939, n12940, n12941, n12942,
    n12943, n12944, n12945, n12946, n12947, n12948,
    n12949, n12950, n12951, n12952, n12953, n12954,
    n12955, n12956, n12957, n12958, n12959, n12960,
    n12961, n12962, n12963, n12964, n12965, n12966,
    n12967, n12968, n12969, n12970, n12971, n12972,
    n12973, n12974, n12975, n12976, n12977, n12978,
    n12979, n12980, n12981, n12982, n12983, n12984,
    n12985, n12986, n12987, n12988, n12989, n12990,
    n12991, n12992, n12993, n12994, n12995, n12996,
    n12997, n12998, n12999, n13000, n13001, n13002,
    n13003, n13004, n13005, n13006, n13007, n13008,
    n13009, n13010, n13011, n13012, n13013, n13014,
    n13015, n13016, n13017, n13018, n13019, n13020,
    n13021, n13022, n13023, n13024, n13025, n13026,
    n13027, n13028, n13029, n13030, n13031, n13032,
    n13033, n13034, n13035, n13036, n13037, n13038,
    n13039, n13040, n13041, n13042, n13043, n13044,
    n13045, n13046, n13047, n13048, n13049, n13050,
    n13051, n13052, n13053, n13054, n13055, n13056,
    n13057, n13058, n13059, n13060, n13061, n13062,
    n13063, n13064, n13065, n13066, n13067, n13068,
    n13069, n13070, n13071, n13072, n13073, n13074,
    n13075, n13076, n13077, n13078, n13079, n13080,
    n13081, n13082, n13083, n13084, n13085, n13086,
    n13087, n13088, n13089, n13090, n13091, n13092,
    n13093, n13094, n13095, n13096, n13097, n13098,
    n13099, n13100, n13101, n13102, n13103, n13104,
    n13105, n13106, n13107, n13108, n13109, n13110,
    n13111, n13112, n13113, n13114, n13115, n13116,
    n13117, n13118, n13119, n13120, n13121, n13122,
    n13123, n13124, n13125, n13126, n13127, n13128,
    n13129, n13130, n13131, n13132, n13133, n13134,
    n13135, n13136, n13137, n13138, n13139, n13140,
    n13141, n13142, n13143, n13144, n13145, n13146,
    n13147, n13148, n13149, n13150, n13151, n13152,
    n13153, n13154, n13155, n13156, n13157, n13158,
    n13159, n13160, n13161, n13162, n13163, n13164,
    n13165, n13166, n13167, n13168, n13169, n13170,
    n13171, n13172, n13173, n13174, n13175, n13176,
    n13177, n13178, n13179, n13180, n13181, n13182,
    n13183, n13184, n13185, n13186, n13187, n13188,
    n13189, n13190, n13191, n13192, n13193, n13194,
    n13195, n13196, n13197, n13198, n13199, n13200,
    n13201, n13202, n13203, n13204, n13205, n13207,
    n13208, n13209, n13210, n13211, n13212, n13213,
    n13214, n13215, n13216, n13217, n13218, n13219,
    n13220, n13221, n13222, n13223, n13224, n13225,
    n13226, n13227, n13228, n13229, n13230, n13231,
    n13232, n13233, n13234, n13235, n13236, n13237,
    n13238, n13239, n13240, n13241, n13242, n13243,
    n13244, n13245, n13246, n13247, n13248, n13249,
    n13250, n13251, n13252, n13253, n13254, n13255,
    n13256, n13257, n13258, n13260, n13261, n13262,
    n13263, n13264, n13265, n13266, n13267, n13268,
    n13269, n13270, n13271, n13272, n13273, n13274,
    n13275, n13276, n13277, n13278, n13279, n13280,
    n13281, n13282, n13283, n13284, n13285, n13286,
    n13287, n13288, n13289, n13290, n13291, n13292,
    n13293, n13294, n13295, n13296, n13297, n13298,
    n13299, n13300, n13301, n13302, n13303, n13304,
    n13305, n13306, n13307, n13308, n13309, n13310,
    n13311, n13312, n13313, n13314, n13315, n13316,
    n13317, n13318, n13319, n13320, n13321, n13322,
    n13323, n13324, n13325, n13326, n13327, n13328,
    n13329, n13330, n13331, n13332, n13333, n13334,
    n13335, n13336, n13337, n13338, n13339, n13340,
    n13341, n13342, n13343, n13344, n13345, n13346,
    n13347, n13348, n13349, n13350, n13351, n13352,
    n13353, n13354, n13355, n13356, n13357, n13358,
    n13359, n13360, n13361, n13362, n13363, n13364,
    n13365, n13366, n13367, n13368, n13369, n13370,
    n13371, n13372, n13373, n13374, n13375, n13376,
    n13377, n13378, n13379, n13380, n13381, n13382,
    n13383, n13384, n13385, n13386, n13387, n13388,
    n13389, n13390, n13391, n13392, n13393, n13394,
    n13395, n13396, n13397, n13398, n13399, n13400,
    n13401, n13402, n13403, n13404, n13405, n13406,
    n13407, n13408, n13409, n13410, n13411, n13412,
    n13413, n13414, n13415, n13416, n13417, n13418,
    n13419, n13420, n13421, n13422, n13423, n13424,
    n13425, n13426, n13427, n13428, n13429, n13430,
    n13431, n13432, n13433, n13434, n13435, n13436,
    n13437, n13438, n13439, n13440, n13441, n13442,
    n13443, n13444, n13445, n13446, n13447, n13448,
    n13449, n13450, n13451, n13452, n13453, n13454,
    n13455, n13456, n13457, n13458, n13459, n13460,
    n13461, n13462, n13463, n13464, n13465, n13466,
    n13467, n13468, n13469, n13470, n13471, n13472,
    n13473, n13474, n13475, n13476, n13477, n13478,
    n13479, n13480, n13481, n13482, n13483, n13484,
    n13485, n13486, n13487, n13488, n13489, n13490,
    n13491, n13492, n13493, n13494, n13495, n13496,
    n13497, n13498, n13499, n13500, n13501, n13502,
    n13503, n13504, n13505, n13506, n13507, n13508,
    n13509, n13510, n13511, n13512, n13513, n13514,
    n13515, n13516, n13517, n13518, n13519, n13520,
    n13521, n13522, n13523, n13524, n13525, n13526,
    n13527, n13528, n13529, n13530, n13531, n13532,
    n13533, n13534, n13535, n13536, n13537, n13538,
    n13539, n13540, n13541, n13542, n13543, n13544,
    n13545, n13546, n13547, n13548, n13549, n13550,
    n13551, n13552, n13553, n13554, n13555, n13556,
    n13557, n13558, n13559, n13560, n13561, n13562,
    n13563, n13564, n13565, n13566, n13567, n13568,
    n13569, n13570, n13571, n13572, n13573, n13574,
    n13575, n13576, n13577, n13578, n13579, n13580,
    n13581, n13582, n13583, n13584, n13585, n13586,
    n13587, n13588, n13589, n13590, n13591, n13592,
    n13593, n13594, n13595, n13596, n13597, n13598,
    n13599, n13600, n13601, n13603, n13604, n13605,
    n13606, n13607, n13608, n13609, n13610, n13611,
    n13612, n13613, n13614, n13615, n13616, n13617,
    n13618, n13619, n13620, n13621, n13622, n13623,
    n13624, n13625, n13626, n13627, n13628, n13629,
    n13630, n13631, n13632, n13633, n13634, n13635,
    n13636, n13637, n13638, n13639, n13640, n13641,
    n13642, n13643, n13644, n13645, n13646, n13647,
    n13648, n13649, n13650, n13651, n13652, n13653,
    n13654, n13655, n13656, n13657, n13658, n13659,
    n13660, n13661, n13662, n13663, n13664, n13665,
    n13666, n13667, n13668, n13669, n13670, n13671,
    n13672, n13673, n13674, n13675, n13676, n13677,
    n13678, n13679, n13680, n13681, n13682, n13683,
    n13684, n13685, n13686, n13687, n13688, n13689,
    n13690, n13691, n13692, n13693, n13694, n13695,
    n13696, n13697, n13698, n13699, n13700, n13701,
    n13702, n13703, n13704, n13705, n13706, n13707,
    n13708, n13709, n13710, n13711, n13712, n13713,
    n13714, n13715, n13716, n13717, n13718, n13719,
    n13720, n13721, n13722, n13723, n13724, n13725,
    n13726, n13727, n13728, n13729, n13730, n13731,
    n13732, n13733, n13734, n13735, n13736, n13737,
    n13738, n13739, n13740, n13741, n13742, n13743,
    n13744, n13745, n13746, n13747, n13748, n13749,
    n13750, n13751, n13752, n13753, n13754, n13755,
    n13756, n13757, n13758, n13759, n13760, n13761,
    n13762, n13763, n13764, n13765, n13766, n13767,
    n13768, n13769, n13770, n13771, n13772, n13773,
    n13774, n13775, n13776, n13777, n13778, n13779,
    n13780, n13781, n13782, n13783, n13784, n13785,
    n13786, n13787, n13788, n13789, n13790, n13791,
    n13792, n13793, n13794, n13795, n13796, n13797,
    n13798, n13799, n13800, n13801, n13802, n13803,
    n13804, n13805, n13806, n13807, n13808, n13809,
    n13810, n13811, n13812, n13813, n13814, n13815,
    n13816, n13817, n13818, n13819, n13820, n13821,
    n13822, n13823, n13824, n13825, n13826, n13827,
    n13828, n13829, n13830, n13831, n13832, n13833,
    n13834, n13835, n13836, n13837, n13838, n13839,
    n13840, n13841, n13842, n13843, n13844, n13845,
    n13846, n13847, n13848, n13849, n13850, n13851,
    n13852, n13853, n13854, n13855, n13856, n13857,
    n13858, n13859, n13860, n13861, n13862, n13863,
    n13864, n13865, n13866, n13867, n13868, n13869,
    n13870, n13871, n13872, n13873, n13874, n13875,
    n13876, n13877, n13878, n13879, n13880, n13881,
    n13882, n13883, n13884, n13885, n13886, n13887,
    n13888, n13889, n13890, n13891, n13892, n13893,
    n13894, n13895, n13896, n13897, n13898, n13899,
    n13900, n13901, n13902, n13903, n13904, n13905,
    n13906, n13907, n13908, n13909, n13910, n13911,
    n13912, n13913, n13914, n13915, n13916, n13917,
    n13918, n13919, n13920, n13921, n13922, n13923,
    n13924, n13925, n13926, n13927, n13928, n13929,
    n13930, n13931, n13932, n13933, n13934, n13935,
    n13936, n13937, n13938, n13939, n13940, n13941,
    n13942, n13943, n13944, n13945, n13946, n13947,
    n13948, n13949, n13950, n13951, n13952, n13953,
    n13954, n13955, n13956, n13957, n13958, n13959,
    n13960, n13961, n13962, n13963, n13964, n13965,
    n13966, n13967, n13968, n13969, n13970, n13971,
    n13972, n13973, n13974, n13975, n13976, n13977,
    n13978, n13979, n13980, n13981, n13982, n13983,
    n13984, n13985, n13986, n13987, n13988, n13989,
    n13990, n13991, n13992, n13993, n13994, n13995,
    n13996, n13997, n13998, n13999, n14000, n14001,
    n14002, n14003, n14004, n14005, n14007, n14008,
    n14009, n14010, n14011, n14012, n14013, n14015,
    n14016, n14017, n14018, n14019, n14020, n14021,
    n14022, n14023, n14024, n14025, n14026, n14027,
    n14028, n14029, n14030, n14031, n14032, n14033,
    n14034, n14035, n14036, n14037, n14038, n14039,
    n14040, n14041, n14042, n14043, n14044, n14045,
    n14046, n14047, n14048, n14049, n14050, n14051,
    n14052, n14053, n14054, n14055, n14056, n14057,
    n14058, n14059, n14060, n14061, n14062, n14063,
    n14064, n14065, n14066, n14067, n14069, n14070,
    n14071, n14072, n14073, n14074, n14075, n14076,
    n14077, n14078, n14079, n14080, n14081, n14082,
    n14083, n14084, n14085, n14086, n14087, n14088,
    n14089, n14090, n14091, n14092, n14093, n14094,
    n14095, n14096, n14097, n14098, n14099, n14100,
    n14101, n14102, n14103, n14104, n14105, n14106,
    n14107, n14108, n14109, n14110, n14111, n14112,
    n14113, n14114, n14115, n14116, n14117, n14118,
    n14119, n14120, n14121, n14122, n14123, n14124,
    n14125, n14126, n14127, n14128, n14129, n14130,
    n14131, n14132, n14133, n14134, n14135, n14136,
    n14137, n14138, n14139, n14140, n14141, n14142,
    n14143, n14144, n14145, n14146, n14147, n14148,
    n14149, n14150, n14151, n14152, n14153, n14154,
    n14155, n14156, n14157, n14158, n14159, n14160,
    n14161, n14162, n14163, n14164, n14165, n14166,
    n14167, n14168, n14169, n14170, n14171, n14172,
    n14173, n14174, n14175, n14176, n14177, n14178,
    n14179, n14180, n14181, n14182, n14183, n14184,
    n14185, n14186, n14187, n14188, n14189, n14190,
    n14191, n14192, n14193, n14194, n14195, n14196,
    n14197, n14198, n14199, n14200, n14201, n14202,
    n14203, n14204, n14205, n14206, n14207, n14208,
    n14209, n14210, n14211, n14212, n14213, n14214,
    n14215, n14216, n14217, n14218, n14219, n14220,
    n14221, n14222, n14223, n14224, n14225, n14226,
    n14227, n14228, n14229, n14230, n14231, n14232,
    n14233, n14234, n14235, n14236, n14237, n14238,
    n14239, n14240, n14241, n14242, n14243, n14244,
    n14245, n14246, n14247, n14248, n14249, n14250,
    n14251, n14252, n14253, n14254, n14255, n14256,
    n14257, n14258, n14259, n14260, n14261, n14262,
    n14263, n14264, n14265, n14266, n14267, n14268,
    n14269, n14270, n14271, n14272, n14273, n14274,
    n14275, n14276, n14277, n14278, n14279, n14280,
    n14281, n14282, n14283, n14284, n14285, n14286,
    n14287, n14288, n14289, n14290, n14291, n14292,
    n14293, n14294, n14295, n14296, n14297, n14298,
    n14299, n14300, n14301, n14302, n14303, n14304,
    n14305, n14306, n14307, n14308, n14309, n14310,
    n14311, n14312, n14313, n14314, n14315, n14316,
    n14317, n14318, n14319, n14320, n14321, n14322,
    n14323, n14324, n14325, n14326, n14327, n14328,
    n14329, n14330, n14331, n14332, n14333, n14334,
    n14335, n14336, n14337, n14338, n14339, n14340,
    n14341, n14342, n14343, n14344, n14345, n14346,
    n14347, n14348, n14349, n14350, n14351, n14352,
    n14353, n14354, n14355, n14356, n14357, n14358,
    n14359, n14360, n14361, n14362, n14363, n14364,
    n14365, n14366, n14367, n14368, n14369, n14370,
    n14371, n14372, n14373, n14374, n14375, n14376,
    n14377, n14378, n14379, n14380, n14381, n14382,
    n14383, n14384, n14385, n14386, n14387, n14388,
    n14389, n14390, n14391, n14392, n14393, n14394,
    n14395, n14396, n14397, n14398, n14399, n14400,
    n14401, n14402, n14403, n14404, n14405, n14406,
    n14407, n14408, n14409, n14410, n14411, n14412,
    n14413, n14414, n14415, n14416, n14417, n14418,
    n14419, n14420, n14421, n14422, n14423, n14424,
    n14425, n14426, n14427, n14428, n14429, n14430,
    n14431, n14432, n14433, n14434, n14435, n14436,
    n14437, n14438, n14439, n14440, n14441, n14442,
    n14443, n14444, n14445, n14446, n14447, n14448,
    n14449, n14450, n14451, n14453, n14454, n14455,
    n14456, n14457, n14458, n14459, n14460, n14461,
    n14462, n14463, n14464, n14465, n14466, n14467,
    n14468, n14469, n14470, n14471, n14472, n14473,
    n14474, n14475, n14476, n14477, n14478, n14479,
    n14480, n14481, n14482, n14483, n14484, n14485,
    n14486, n14487, n14488, n14489, n14490, n14491,
    n14492, n14493, n14494, n14495, n14496, n14497,
    n14498, n14499, n14500, n14501, n14502, n14503,
    n14504, n14505, n14506, n14507, n14508, n14509,
    n14510, n14511, n14512, n14513, n14514, n14515,
    n14516, n14517, n14518, n14519, n14520, n14521,
    n14522, n14523, n14524, n14525, n14526, n14527,
    n14528, n14529, n14530, n14531, n14532, n14533,
    n14534, n14535, n14536, n14537, n14538, n14539,
    n14540, n14541, n14542, n14543, n14544, n14545,
    n14546, n14547, n14548, n14549, n14550, n14551,
    n14552, n14553, n14554, n14555, n14556, n14557,
    n14558, n14559, n14560, n14561, n14562, n14563,
    n14564, n14565, n14566, n14567, n14568, n14569,
    n14570, n14571, n14572, n14573, n14574, n14575,
    n14576, n14577, n14578, n14579, n14580, n14581,
    n14582, n14583, n14584, n14585, n14586, n14587,
    n14588, n14589, n14590, n14591, n14592, n14593,
    n14594, n14595, n14596, n14597, n14598, n14599,
    n14600, n14601, n14602, n14603, n14604, n14605,
    n14606, n14607, n14608, n14609, n14610, n14611,
    n14612, n14613, n14614, n14615, n14616, n14617,
    n14618, n14619, n14620, n14621, n14622, n14623,
    n14624, n14625, n14626, n14627, n14628, n14629,
    n14630, n14631, n14632, n14633, n14634, n14635,
    n14636, n14637, n14638, n14639, n14640, n14641,
    n14642, n14643, n14644, n14645, n14646, n14647,
    n14648, n14649, n14650, n14651, n14652, n14653,
    n14654, n14655, n14656, n14657, n14658, n14659,
    n14660, n14661, n14662, n14663, n14664, n14665,
    n14666, n14667, n14668, n14669, n14670, n14671,
    n14672, n14673, n14674, n14675, n14676, n14677,
    n14678, n14679, n14680, n14681, n14682, n14683,
    n14684, n14685, n14686, n14687, n14688, n14689,
    n14690, n14691, n14692, n14693, n14694, n14695,
    n14696, n14697, n14698, n14699, n14700, n14701,
    n14702, n14703, n14704, n14705, n14706, n14707,
    n14708, n14709, n14710, n14711, n14712, n14713,
    n14714, n14715, n14716, n14717, n14718, n14719,
    n14720, n14721, n14722, n14723, n14724, n14725,
    n14726, n14727, n14728, n14729, n14730, n14731,
    n14732, n14733, n14734, n14735, n14736, n14737,
    n14738, n14739, n14740, n14741, n14742, n14743,
    n14744, n14745, n14746, n14747, n14748, n14749,
    n14751, n14752, n14753, n14754, n14755, n14756,
    n14757, n14758, n14759, n14760, n14761, n14762,
    n14763, n14764, n14765, n14766, n14767, n14768,
    n14769, n14770, n14771, n14772, n14773, n14774,
    n14775, n14776, n14777, n14778, n14779, n14780,
    n14781, n14782, n14783, n14784, n14785, n14786,
    n14787, n14788, n14789, n14790, n14791, n14792,
    n14793, n14794, n14795, n14796, n14797, n14798,
    n14799, n14800, n14801, n14802, n14803, n14804,
    n14805, n14806, n14807, n14808, n14809, n14810,
    n14811, n14812, n14813, n14814, n14815, n14816,
    n14817, n14818, n14819, n14820, n14821, n14822,
    n14823, n14824, n14825, n14826, n14827, n14828,
    n14829, n14831, n14832, n14833, n14834, n14835,
    n14836, n14837, n14838, n14839, n14840, n14841,
    n14842, n14843, n14844, n14845, n14846, n14847,
    n14848, n14849, n14850, n14851, n14852, n14853,
    n14854, n14856, n14857, n14858, n14859, n14860,
    n14861, n14862, n14863, n14864, n14865, n14866,
    n14867, n14868, n14869, n14870, n14871, n14872,
    n14873, n14874, n14875, n14876, n14877, n14878,
    n14879, n14880, n14881, n14882, n14883, n14884,
    n14885, n14886, n14887, n14888, n14889, n14890,
    n14891, n14892, n14893, n14894, n14895, n14896,
    n14897, n14898, n14899, n14900, n14901, n14902,
    n14903, n14904, n14905, n14906, n14907, n14908,
    n14909, n14910, n14911, n14912, n14913, n14914,
    n14915, n14916, n14917, n14918, n14919, n14920,
    n14921, n14922, n14923, n14924, n14925, n14926,
    n14927, n14928, n14929, n14930, n14931, n14932,
    n14933, n14934, n14935, n14936, n14937, n14938,
    n14939, n14940, n14941, n14942, n14943, n14944,
    n14945, n14946, n14947, n14948, n14949, n14950,
    n14951, n14952, n14953, n14954, n14955, n14956,
    n14957, n14958, n14959, n14960, n14961, n14962,
    n14963, n14964, n14965, n14966, n14967, n14968,
    n14969, n14970, n14971, n14972, n14973, n14974,
    n14975, n14976, n14977, n14978, n14980, n14981,
    n14982, n14983, n14984, n14985, n14987, n14988,
    n14989, n14990, n14991, n14992, n14993, n14994,
    n14995, n14996, n14997, n14998, n14999, n15000,
    n15001, n15002, n15003, n15004, n15005, n15006,
    n15007, n15008, n15009, n15010, n15011, n15012,
    n15013, n15014, n15015, n15016, n15017, n15018,
    n15019, n15020, n15021, n15022, n15023, n15024,
    n15025, n15026, n15027, n15028, n15029, n15030,
    n15031, n15032, n15033, n15034, n15035, n15036,
    n15037, n15038, n15039, n15040, n15041, n15042,
    n15043, n15044, n15045, n15046, n15047, n15048,
    n15049, n15050, n15051, n15052, n15053, n15054,
    n15055, n15056, n15057, n15058, n15059, n15060,
    n15061, n15062, n15063, n15064, n15065, n15066,
    n15067, n15068, n15069, n15070, n15071, n15072,
    n15073, n15074, n15075, n15076, n15077, n15078,
    n15079, n15080, n15081, n15082, n15083, n15084,
    n15085, n15086, n15087, n15088, n15089, n15090,
    n15091, n15092, n15093, n15094, n15095, n15096,
    n15097, n15098, n15099, n15100, n15101, n15102,
    n15103, n15104, n15105, n15106, n15107, n15108,
    n15109, n15110, n15111, n15112, n15113, n15114,
    n15115, n15116, n15117, n15118, n15119, n15120,
    n15121, n15122, n15123, n15124, n15125, n15126,
    n15127, n15128, n15129, n15130, n15131, n15132,
    n15133, n15134, n15135, n15136, n15137, n15138,
    n15139, n15140, n15141, n15142, n15143, n15144,
    n15145, n15146, n15147, n15148, n15149, n15150,
    n15151, n15152, n15153, n15154, n15155, n15156,
    n15157, n15158, n15159, n15160, n15161, n15162,
    n15163, n15164, n15165, n15166, n15167, n15168,
    n15169, n15170, n15171, n15172, n15173, n15174,
    n15175, n15176, n15177, n15178, n15179, n15180,
    n15181, n15182, n15183, n15184, n15185, n15186,
    n15187, n15188, n15189, n15190, n15191, n15192,
    n15193, n15194, n15195, n15197, n15198, n15199,
    n15200, n15201, n15202, n15203, n15204, n15205,
    n15206, n15207, n15208, n15209, n15210, n15211,
    n15212, n15213, n15214, n15215, n15216, n15217,
    n15218, n15219, n15220, n15221, n15222, n15223,
    n15224, n15225, n15226, n15227, n15228, n15229,
    n15230, n15231, n15232, n15233, n15234, n15235,
    n15236, n15237, n15238, n15239, n15240, n15241,
    n15242, n15243, n15244, n15245, n15246, n15247,
    n15248, n15249, n15250, n15251, n15253, n15254,
    n15255, n15256, n15257, n15258, n15259, n15260,
    n15261, n15262, n15263, n15264, n15265, n15266,
    n15267, n15268, n15269, n15270, n15271, n15272,
    n15273, n15274, n15275, n15276, n15277, n15278,
    n15279, n15280, n15281, n15282, n15283, n15284,
    n15285, n15286, n15287, n15288, n15289, n15290,
    n15291, n15292, n15293, n15294, n15295, n15296,
    n15297, n15298, n15299, n15300, n15301, n15302,
    n15303, n15304, n15305, n15306, n15307, n15308,
    n15309, n15310, n15311, n15312, n15313, n15314,
    n15315, n15316, n15317, n15318, n15319, n15320,
    n15321, n15322, n15323, n15324, n15325, n15326,
    n15327, n15328, n15329, n15330, n15331, n15332,
    n15333, n15334, n15335, n15336, n15337, n15338,
    n15339, n15340, n15341, n15342, n15343, n15344,
    n15345, n15346, n15347, n15348, n15349, n15350,
    n15351, n15352, n15353, n15354, n15355, n15356,
    n15357, n15358, n15359, n15360, n15361, n15362,
    n15363, n15364, n15366, n15367, n15368, n15369,
    n15370, n15371, n15372, n15373, n15374, n15375,
    n15376, n15377, n15378, n15379, n15380, n15381,
    n15382, n15383, n15384, n15385, n15386, n15387,
    n15388, n15389, n15390, n15391, n15392, n15393,
    n15394, n15395, n15396, n15397, n15398, n15399,
    n15400, n15401, n15402, n15403, n15404, n15405,
    n15406, n15407, n15408, n15409, n15410, n15411,
    n15412, n15413, n15414, n15415, n15416, n15417,
    n15418, n15419, n15420, n15421, n15422, n15423,
    n15424, n15425, n15426, n15427, n15428, n15429,
    n15430, n15431, n15432, n15433, n15434, n15435,
    n15436, n15437, n15438, n15439, n15440, n15441,
    n15442, n15443, n15444, n15445, n15446, n15447,
    n15448, n15449, n15450, n15451, n15452, n15453,
    n15454, n15455, n15456, n15457, n15458, n15459,
    n15460, n15461, n15462, n15463, n15464, n15465,
    n15466, n15467, n15468, n15469, n15470, n15471,
    n15472, n15473, n15474, n15475, n15476, n15477,
    n15478, n15479, n15480, n15481, n15482, n15483,
    n15485, n15486, n15487, n15488, n15489, n15490,
    n15491, n15492, n15493, n15494, n15495, n15496,
    n15497, n15498, n15499, n15500, n15501, n15502,
    n15503, n15504, n15505, n15506, n15507, n15508,
    n15509, n15510, n15511, n15512, n15513, n15514,
    n15515, n15516, n15517, n15518, n15519, n15520,
    n15521, n15522, n15523, n15524, n15525, n15526,
    n15527, n15528, n15529, n15530, n15531, n15532,
    n15533, n15534, n15535, n15536, n15537, n15538,
    n15539, n15540, n15541, n15542, n15543, n15544,
    n15545, n15546, n15547, n15548, n15549, n15550,
    n15551, n15552, n15553, n15554, n15555, n15556,
    n15557, n15558, n15559, n15560, n15561, n15562,
    n15563, n15564, n15565, n15566, n15567, n15568,
    n15570, n15571, n15572, n15573, n15574, n15575,
    n15576, n15577, n15578, n15579, n15580, n15581,
    n15583, n15584, n15585, n15586, n15587, n15588,
    n15589, n15590, n15591, n15592, n15593, n15594,
    n15595, n15596, n15597, n15598, n15599, n15600,
    n15601, n15602, n15603, n15604, n15605, n15606,
    n15607, n15608, n15609, n15610, n15611, n15612,
    n15613, n15614, n15615, n15616, n15617, n15618,
    n15619, n15620, n15621, n15622, n15623, n15624,
    n15625, n15626, n15627, n15628, n15629, n15630,
    n15631, n15632, n15633, n15634, n15635, n15636,
    n15637, n15638, n15639, n15640, n15641, n15642,
    n15643, n15644, n15645, n15646, n15647, n15648,
    n15649, n15650, n15651, n15652, n15653, n15654,
    n15655, n15656, n15657, n15658, n15659, n15660,
    n15661, n15662, n15663, n15665, n15666, n15667,
    n15668, n15669, n15670, n15671, n15672, n15673,
    n15674, n15675, n15676, n15677, n15678, n15679,
    n15680, n15681, n15682, n15683, n15684, n15685,
    n15686, n15687, n15688, n15689, n15690, n15691,
    n15692, n15693, n15694, n15695, n15696, n15697,
    n15698, n15699, n15700, n15701, n15702, n15703,
    n15704, n15705, n15706, n15707, n15708, n15709,
    n15710, n15711, n15712, n15713, n15714, n15715,
    n15716, n15717, n15718, n15719, n15720, n15722,
    n15723, n15724, n15725, n15726, n15727, n15728,
    n15729, n15730, n15731, n15732, n15733, n15734,
    n15735, n15736, n15737, n15738, n15739, n15740,
    n15741, n15742, n15743, n15744, n15745, n15746,
    n15747, n15748, n15749, n15750, n15751, n15752,
    n15753, n15754, n15755, n15756, n15757, n15758,
    n15759, n15760, n15761, n15762, n15763, n15764,
    n15765, n15766, n15767, n15768, n15769, n15770,
    n15771, n15772, n15773, n15774, n15775, n15776,
    n15777, n15778, n15779, n15780, n15781, n15782,
    n15783, n15784, n15785, n15786, n15787, n15788,
    n15789, n15790, n15791, n15792, n15793, n15794,
    n15795, n15796, n15797, n15798, n15799, n15800,
    n15801, n15802, n15803, n15804, n15805, n15806,
    n15807, n15808, n15809, n15810, n15811, n15812,
    n15813, n15814, n15815, n15816, n15817, n15818,
    n15819, n15820, n15821, n15822, n15823, n15824,
    n15825, n15826, n15827, n15828, n15829, n15830,
    n15831, n15832, n15833, n15834, n15835, n15836,
    n15837, n15838, n15839, n15840, n15841, n15842,
    n15843, n15844, n15845, n15846, n15847, n15848,
    n15849, n15850, n15851, n15852, n15853, n15854,
    n15855, n15856, n15857, n15858, n15859, n15860,
    n15861, n15862, n15863, n15864, n15865, n15866,
    n15867, n15868, n15869, n15870, n15871, n15872,
    n15873, n15874, n15875, n15876, n15877, n15878,
    n15879, n15880, n15881, n15882, n15883, n15884,
    n15885, n15886, n15887, n15888, n15889, n15890,
    n15891, n15892, n15893, n15894, n15895, n15896,
    n15897, n15898, n15899, n15900, n15901, n15902,
    n15903, n15904, n15905, n15906, n15907, n15908,
    n15909, n15910, n15911, n15912, n15913, n15914,
    n15915, n15916, n15917, n15918, n15919, n15920,
    n15921, n15922, n15923, n15924, n15925, n15926,
    n15927, n15928, n15929, n15930, n15931, n15932,
    n15933, n15934, n15935, n15936, n15937, n15938,
    n15939, n15940, n15941, n15942, n15943, n15944,
    n15945, n15946, n15947, n15948, n15949, n15950,
    n15951, n15952, n15953, n15954, n15955, n15956,
    n15957, n15958, n15959, n15960, n15961, n15962,
    n15963, n15964, n15965, n15966, n15967, n15968,
    n15969, n15970, n15971, n15972, n15973, n15974,
    n15975, n15976, n15977, n15978, n15979, n15980,
    n15981, n15982, n15983, n15984, n15985, n15986,
    n15987, n15988, n15989, n15990, n15991, n15992,
    n15993, n15994, n15995, n15996, n15997, n15998,
    n15999, n16000, n16001, n16002, n16003, n16004,
    n16005, n16006, n16007, n16008, n16009, n16010,
    n16011, n16012, n16013, n16014, n16015, n16016,
    n16017, n16018, n16019, n16020, n16021, n16022,
    n16023, n16024, n16025, n16026, n16027, n16028,
    n16029, n16030, n16031, n16032, n16033, n16034,
    n16035, n16036, n16037, n16038, n16039, n16040,
    n16041, n16042, n16043, n16044, n16045, n16046,
    n16047, n16048, n16049, n16050, n16051, n16052,
    n16053, n16054, n16055, n16056, n16057, n16058,
    n16059, n16060, n16061, n16062, n16063, n16064,
    n16065, n16066, n16067, n16068, n16069, n16070,
    n16071, n16072, n16073, n16074, n16075, n16076,
    n16077, n16078, n16079, n16080, n16081, n16082,
    n16083, n16084, n16085, n16086, n16087, n16088,
    n16089, n16090, n16091, n16092, n16093, n16094,
    n16095, n16096, n16097, n16098, n16099, n16100,
    n16101, n16102, n16103, n16104, n16105, n16106,
    n16107, n16108, n16109, n16110, n16111, n16112,
    n16113, n16114, n16115, n16116, n16117, n16118,
    n16119, n16120, n16121, n16122, n16123, n16124,
    n16125, n16126, n16127, n16128, n16129, n16130,
    n16131, n16132, n16133, n16134, n16135, n16136,
    n16137, n16138, n16139, n16140, n16141, n16142,
    n16143, n16144, n16145, n16146, n16147, n16148,
    n16149, n16150, n16151, n16152, n16153, n16154,
    n16155, n16156, n16157, n16158, n16159, n16160,
    n16161, n16162, n16163, n16164, n16165, n16166,
    n16167, n16168, n16169, n16170, n16171, n16172,
    n16173, n16174, n16175, n16176, n16177, n16178,
    n16179, n16180, n16181, n16182, n16183, n16184,
    n16185, n16186, n16187, n16188, n16189, n16190,
    n16191, n16192, n16193, n16194, n16195, n16196,
    n16197, n16198, n16199, n16200, n16201, n16202,
    n16203, n16204, n16205, n16206, n16207, n16208,
    n16209, n16210, n16211, n16212, n16213, n16214,
    n16215, n16216, n16217, n16218, n16219, n16220,
    n16221, n16222, n16223, n16224, n16225, n16226,
    n16227, n16228, n16229, n16230, n16231, n16232,
    n16233, n16234, n16235, n16236, n16237, n16238,
    n16239, n16240, n16241, n16242, n16243, n16244,
    n16245, n16246, n16247, n16248, n16249, n16250,
    n16251, n16252, n16253, n16254, n16255, n16256,
    n16257, n16258, n16259, n16260, n16261, n16262,
    n16263, n16264, n16265, n16266, n16267, n16268,
    n16269, n16270, n16271, n16272, n16273, n16274,
    n16275, n16276, n16277, n16278, n16279, n16280,
    n16281, n16282, n16283, n16284, n16285, n16286,
    n16287, n16288, n16289, n16290, n16291, n16292,
    n16293, n16294, n16295, n16296, n16297, n16298,
    n16299, n16300, n16301, n16302, n16303, n16304,
    n16305, n16306, n16307, n16308, n16309, n16310,
    n16311, n16312, n16313, n16314, n16315, n16316,
    n16317, n16318, n16319, n16320, n16321, n16322,
    n16323, n16324, n16325, n16326, n16327, n16328,
    n16329, n16330, n16331, n16332, n16333, n16334,
    n16335, n16336, n16337, n16338, n16339, n16340,
    n16341, n16342, n16343, n16344, n16345, n16346,
    n16347, n16348, n16349, n16350, n16351, n16352,
    n16353, n16354, n16355, n16356, n16357, n16358,
    n16359, n16360, n16361, n16362, n16363, n16364,
    n16365, n16366, n16367, n16368, n16369, n16370,
    n16371, n16372, n16373, n16374, n16375, n16376,
    n16377, n16378, n16379, n16380, n16381, n16382,
    n16383, n16384, n16385, n16386, n16387, n16388,
    n16389, n16390, n16391, n16392, n16393, n16394,
    n16395, n16396, n16397, n16398, n16399, n16400,
    n16401, n16402, n16403, n16404, n16405, n16406,
    n16407, n16408, n16409, n16410, n16411, n16412,
    n16413, n16414, n16415, n16416, n16417, n16418,
    n16419, n16420, n16421, n16422, n16423, n16424,
    n16425, n16426, n16427, n16428, n16429, n16430,
    n16431, n16432, n16433, n16434, n16435, n16436,
    n16437, n16438, n16439, n16440, n16441, n16442,
    n16443, n16444, n16445, n16446, n16447, n16448,
    n16449, n16450, n16451, n16452, n16453, n16454,
    n16455, n16456, n16457, n16458, n16459, n16460,
    n16461, n16462, n16463, n16464, n16465, n16466,
    n16467, n16468, n16469, n16470, n16471, n16472,
    n16473, n16474, n16475, n16476, n16477, n16478,
    n16479, n16480, n16481, n16482, n16483, n16484,
    n16485, n16486, n16487, n16488, n16489, n16490,
    n16491, n16492, n16493, n16494, n16495, n16496,
    n16497, n16498, n16499, n16500, n16501, n16502,
    n16503, n16504, n16505, n16506, n16507, n16508,
    n16509, n16510, n16511, n16512, n16513, n16514,
    n16515, n16516, n16517, n16518, n16519, n16520,
    n16521, n16522, n16523, n16524, n16525, n16526,
    n16527, n16528, n16529, n16530, n16531, n16532,
    n16533, n16534, n16535, n16536, n16537, n16538,
    n16539, n16540, n16541, n16542, n16543, n16544,
    n16545, n16546, n16547, n16548, n16549, n16550,
    n16551, n16552, n16553, n16554, n16555, n16556,
    n16557, n16558, n16559, n16560, n16561, n16562,
    n16563, n16564, n16565, n16566, n16567, n16568,
    n16569, n16570, n16571, n16572, n16573, n16574,
    n16575, n16576, n16577, n16578, n16579, n16580,
    n16581, n16582, n16583, n16584, n16585, n16586,
    n16587, n16588, n16589, n16590, n16591, n16592,
    n16593, n16594, n16595, n16596, n16597, n16598,
    n16599, n16600, n16601, n16602, n16603, n16604,
    n16605, n16606, n16607, n16608, n16609, n16610,
    n16611, n16612, n16613, n16614, n16615, n16616,
    n16617, n16618, n16619, n16620, n16621, n16622,
    n16623, n16624, n16625, n16626, n16627, n16628,
    n16629, n16630, n16631, n16632, n16633, n16634,
    n16635, n16636, n16637, n16638, n16639, n16640,
    n16641, n16642, n16643, n16644, n16645, n16646,
    n16647, n16648, n16649, n16650, n16651, n16652,
    n16653, n16654, n16655, n16656, n16657, n16658,
    n16659, n16660, n16661, n16662, n16663, n16664,
    n16665, n16666, n16667, n16668, n16669, n16670,
    n16671, n16672, n16673, n16674, n16675, n16676,
    n16677, n16678, n16679, n16680, n16681, n16682,
    n16683, n16684, n16685, n16686, n16687, n16688,
    n16689, n16690, n16691, n16692, n16693, n16694,
    n16695, n16696, n16697, n16698, n16699, n16700,
    n16701, n16702, n16703, n16704, n16705, n16706,
    n16707, n16708, n16709, n16710, n16711, n16712,
    n16713, n16714, n16715, n16716, n16717, n16718,
    n16719, n16720, n16721, n16722, n16723, n16724,
    n16725, n16726, n16727, n16728, n16729, n16730,
    n16731, n16732, n16733, n16734, n16735, n16736,
    n16737, n16738, n16739, n16740, n16741, n16742,
    n16743, n16744, n16745, n16746, n16747, n16748,
    n16749, n16750, n16751, n16752, n16753, n16754,
    n16755, n16756, n16757, n16758, n16759, n16760,
    n16761, n16762, n16763, n16764, n16765, n16766,
    n16767, n16768, n16769, n16770, n16771, n16772,
    n16773, n16774, n16775, n16776, n16777, n16778,
    n16779, n16780, n16781, n16782, n16783, n16784,
    n16785, n16786, n16787, n16788, n16789, n16790,
    n16791, n16792, n16793, n16794, n16795, n16796,
    n16797, n16798, n16799, n16800, n16801, n16802,
    n16803, n16804, n16805, n16806, n16807, n16808,
    n16809, n16810, n16811, n16812, n16813, n16814,
    n16815, n16816, n16817, n16818, n16819, n16820,
    n16821, n16822, n16823, n16824, n16825, n16826,
    n16827, n16828, n16829, n16830, n16831, n16832,
    n16833, n16834, n16835, n16836, n16837, n16838,
    n16839, n16840, n16841, n16842, n16843, n16844,
    n16845, n16846, n16847, n16848, n16849, n16850,
    n16851, n16852, n16853, n16854, n16855, n16856,
    n16857, n16858, n16859, n16860, n16861, n16862,
    n16863, n16864, n16865, n16866, n16867, n16868,
    n16869, n16870, n16871, n16872, n16873, n16874,
    n16875, n16876, n16877, n16878, n16879, n16880,
    n16881, n16882, n16883, n16884, n16885, n16886,
    n16887, n16888, n16889, n16890, n16891, n16892,
    n16893, n16894, n16895, n16896, n16897, n16898,
    n16899, n16900, n16901, n16902, n16903, n16904,
    n16905, n16906, n16907, n16908, n16909, n16910,
    n16911, n16912, n16913, n16914, n16915, n16916,
    n16917, n16918, n16919, n16920, n16921, n16922,
    n16923, n16924, n16925, n16926, n16927, n16928,
    n16929, n16930, n16931, n16932, n16933, n16934,
    n16935, n16936, n16937, n16938, n16939, n16940,
    n16941, n16942, n16943, n16944, n16945, n16946,
    n16947, n16948, n16949, n16950, n16951, n16952,
    n16953, n16954, n16955, n16956, n16957, n16958,
    n16959, n16960, n16961, n16962, n16963, n16964,
    n16965, n16966, n16967, n16968, n16969, n16970,
    n16971, n16972, n16973, n16974, n16975, n16976,
    n16977, n16978, n16979, n16980, n16981, n16982,
    n16983, n16984, n16985, n16986, n16987, n16988,
    n16989, n16990, n16991, n16992, n16993, n16994,
    n16995, n16996, n16997, n16998, n16999, n17000,
    n17001, n17002, n17003, n17004, n17005, n17006,
    n17007, n17008, n17009, n17010, n17011, n17012,
    n17013, n17014, n17015, n17016, n17017, n17018,
    n17019, n17020, n17021, n17022, n17023, n17024,
    n17025, n17026, n17027, n17028, n17029, n17030,
    n17031, n17032, n17033, n17034, n17035, n17036,
    n17037, n17038, n17039, n17040, n17041, n17042,
    n17043, n17044, n17045, n17046, n17047, n17048,
    n17049, n17050, n17051, n17052, n17053, n17054,
    n17055, n17056, n17057, n17058, n17059, n17060,
    n17061, n17063, n17064, n17065, n17066, n17067,
    n17068, n17069, n17070, n17071, n17072, n17073,
    n17074, n17075, n17076, n17077, n17078, n17079,
    n17080, n17081, n17082, n17083, n17084, n17085,
    n17086, n17087, n17088, n17089, n17090, n17091,
    n17092, n17093, n17094, n17095, n17096, n17097,
    n17098, n17099, n17100, n17101, n17102, n17103,
    n17104, n17105, n17106, n17107, n17108, n17109,
    n17110, n17111, n17112, n17113, n17114, n17115,
    n17116, n17117, n17118, n17119, n17120, n17121,
    n17122, n17123, n17124, n17125, n17126, n17127,
    n17128, n17129, n17130, n17131, n17132, n17133,
    n17134, n17135, n17136, n17137, n17138, n17139,
    n17140, n17141, n17142, n17143, n17144, n17145,
    n17146, n17147, n17148, n17149, n17150, n17151,
    n17152, n17153, n17154, n17155, n17156, n17157,
    n17158, n17159, n17160, n17161, n17162, n17163,
    n17164, n17165, n17166, n17167, n17168, n17169,
    n17170, n17171, n17172, n17173, n17174, n17175,
    n17176, n17177, n17178, n17179, n17180, n17181,
    n17182, n17183, n17184, n17185, n17186, n17187,
    n17188, n17189, n17190, n17191, n17192, n17193,
    n17194, n17195, n17196, n17197, n17198, n17199,
    n17200, n17201, n17202, n17203, n17204, n17205,
    n17206, n17207, n17208, n17209, n17210, n17211,
    n17212, n17213, n17214, n17215, n17216, n17217,
    n17218, n17219, n17220, n17221, n17222, n17223,
    n17224, n17225, n17226, n17227, n17228, n17229,
    n17230, n17231, n17232, n17233, n17234, n17235,
    n17236, n17237, n17238, n17239, n17240, n17241,
    n17242, n17243, n17244, n17245, n17246, n17247,
    n17248, n17249, n17250, n17251, n17252, n17253,
    n17254, n17255, n17256, n17257, n17258, n17259,
    n17260, n17261, n17262, n17263, n17264, n17265,
    n17266, n17267, n17268, n17269, n17270, n17271,
    n17272, n17273, n17274, n17275, n17276, n17277,
    n17278, n17279, n17280, n17281, n17282, n17283,
    n17284, n17285, n17286, n17287, n17288, n17289,
    n17290, n17291, n17292, n17293, n17294, n17295,
    n17296, n17297, n17298, n17299, n17300, n17301,
    n17302, n17303, n17304, n17305, n17306, n17307,
    n17308, n17309, n17310, n17311, n17312, n17313,
    n17314, n17315, n17316, n17317, n17318, n17319,
    n17320, n17321, n17322, n17323, n17324, n17325,
    n17326, n17327, n17328, n17329, n17330, n17331,
    n17332, n17333, n17334, n17335, n17336, n17337,
    n17338, n17339, n17340, n17341, n17342, n17343,
    n17344, n17345, n17346, n17347, n17348, n17349,
    n17350, n17351, n17352, n17353, n17354, n17355,
    n17356, n17357, n17358, n17359, n17360, n17361,
    n17362, n17363, n17364, n17365, n17366, n17367,
    n17368, n17369, n17370, n17371, n17372, n17373,
    n17374, n17375, n17376, n17377, n17378, n17379,
    n17380, n17381, n17382, n17383, n17384, n17385,
    n17386, n17387, n17388, n17389, n17390, n17391,
    n17392, n17393, n17394, n17395, n17396, n17397,
    n17398, n17399, n17400, n17401, n17402, n17403,
    n17404, n17405, n17406, n17407, n17408, n17409,
    n17410, n17411, n17412, n17413, n17414, n17415,
    n17416, n17417, n17418, n17419, n17420, n17421,
    n17422, n17423, n17424, n17425, n17426, n17427,
    n17428, n17429, n17430, n17431, n17432, n17433,
    n17434, n17435, n17436, n17437, n17438, n17439,
    n17440, n17441, n17442, n17443, n17444, n17445,
    n17446, n17447, n17448, n17449, n17450, n17451,
    n17452, n17453, n17454, n17455, n17456, n17457,
    n17458, n17459, n17460, n17461, n17462, n17463,
    n17464, n17465, n17466, n17467, n17468, n17469,
    n17470, n17471, n17472, n17473, n17474, n17475,
    n17476, n17477, n17478, n17479, n17480, n17481,
    n17482, n17483, n17484, n17485, n17486, n17487,
    n17488, n17489, n17490, n17491, n17492, n17493,
    n17494, n17495, n17496, n17497, n17498, n17499,
    n17500, n17501, n17502, n17503, n17504, n17505,
    n17506, n17507, n17508, n17509, n17510, n17511,
    n17512, n17513, n17514, n17515, n17516, n17517,
    n17518, n17519, n17520, n17521, n17522, n17523,
    n17524, n17525, n17526, n17527, n17528, n17529,
    n17530, n17531, n17532, n17533, n17534, n17535,
    n17536, n17537, n17538, n17539, n17540, n17541,
    n17542, n17543, n17544, n17545, n17546, n17547,
    n17548, n17549, n17550, n17551, n17552, n17553,
    n17554, n17555, n17556, n17557, n17558, n17559,
    n17560, n17561, n17562, n17563, n17564, n17565,
    n17566, n17567, n17568, n17569, n17570, n17571,
    n17572, n17573, n17574, n17576, n17577, n17578,
    n17579, n17580, n17581, n17582, n17583, n17584,
    n17585, n17586, n17587, n17588, n17589, n17590,
    n17591, n17592, n17593, n17594, n17595, n17596,
    n17597, n17598, n17599, n17600, n17601, n17602,
    n17603, n17604, n17605, n17606, n17607, n17608,
    n17609, n17610, n17611, n17612, n17613, n17614,
    n17615, n17616, n17617, n17618, n17619, n17620,
    n17621, n17622, n17623, n17624, n17625, n17626,
    n17627, n17628, n17629, n17630, n17631, n17632,
    n17633, n17634, n17635, n17636, n17637, n17638,
    n17639, n17640, n17641, n17642, n17643, n17644,
    n17645, n17646, n17647, n17648, n17649, n17650,
    n17651, n17652, n17653, n17654, n17655, n17656,
    n17657, n17658, n17659, n17660, n17661, n17662,
    n17663, n17664, n17665, n17666, n17667, n17668,
    n17669, n17670, n17671, n17672, n17673, n17674,
    n17675, n17676, n17677, n17678, n17679, n17680,
    n17681, n17682, n17683, n17684, n17685, n17686,
    n17687, n17688, n17689, n17690, n17691, n17692,
    n17693, n17694, n17695, n17696, n17697, n17698,
    n17699, n17700, n17701, n17702, n17703, n17704,
    n17705, n17706, n17707, n17708, n17709, n17710,
    n17711, n17712, n17713, n17714, n17715, n17716,
    n17717, n17718, n17719, n17720, n17721, n17722,
    n17723, n17724, n17725, n17726, n17727, n17728,
    n17729, n17730, n17731, n17732, n17733, n17734,
    n17735, n17736, n17737, n17738, n17739, n17740,
    n17741, n17742, n17743, n17744, n17745, n17746,
    n17747, n17748, n17749, n17750, n17751, n17752,
    n17753, n17754, n17755, n17756, n17757, n17758,
    n17759, n17760, n17761, n17762, n17763, n17764,
    n17765, n17766, n17767, n17768, n17769, n17770,
    n17771, n17772, n17773, n17774, n17775, n17776,
    n17777, n17778, n17779, n17780, n17781, n17782,
    n17783, n17784, n17785, n17786, n17787, n17788,
    n17789, n17790, n17791, n17792, n17793, n17794,
    n17795, n17796, n17797, n17798, n17799, n17800,
    n17801, n17802, n17803, n17804, n17805, n17806,
    n17807, n17808, n17809, n17810, n17811, n17812,
    n17813, n17814, n17815, n17816, n17817, n17818,
    n17819, n17820, n17821, n17822, n17823, n17824,
    n17825, n17826, n17827, n17828, n17829, n17830,
    n17831, n17832, n17833, n17834, n17835, n17836,
    n17837, n17838, n17839, n17840, n17841, n17842,
    n17843, n17844, n17845, n17846, n17847, n17848,
    n17849, n17850, n17851, n17852, n17853, n17854,
    n17855, n17856, n17857, n17858, n17859, n17860,
    n17861, n17862, n17863, n17864, n17865, n17866,
    n17867, n17868, n17869, n17870, n17871, n17872,
    n17873, n17874, n17875, n17876, n17877, n17878,
    n17879, n17880, n17881, n17882, n17883, n17884,
    n17885, n17886, n17887, n17888, n17889, n17890,
    n17891, n17892, n17893, n17894, n17895, n17896,
    n17897, n17898, n17899, n17900, n17901, n17902,
    n17903, n17904, n17905, n17906, n17907, n17908,
    n17909, n17910, n17911, n17912, n17913, n17914,
    n17915, n17916, n17917, n17918, n17919, n17920,
    n17921, n17922, n17923, n17924, n17925, n17926,
    n17927, n17928, n17929, n17930, n17931, n17932,
    n17933, n17934, n17935, n17936, n17937, n17938,
    n17939, n17940, n17941, n17942, n17943, n17944,
    n17945, n17946, n17947, n17948, n17949, n17950,
    n17951, n17952, n17953, n17954, n17955, n17956,
    n17957, n17958, n17959, n17960, n17961, n17962,
    n17963, n17964, n17965, n17966, n17967, n17968,
    n17969, n17970, n17971, n17972, n17973, n17974,
    n17975, n17976, n17977, n17978, n17979, n17980,
    n17981, n17982, n17983, n17984, n17985, n17986,
    n17987, n17988, n17989, n17990, n17991, n17992,
    n17993, n17994, n17995, n17996, n17997, n17998,
    n17999, n18000, n18001, n18002, n18003, n18004,
    n18005, n18006, n18007, n18008, n18009, n18010,
    n18011, n18012, n18013, n18014, n18015, n18016,
    n18017, n18018, n18019, n18020, n18021, n18022,
    n18023, n18024, n18025, n18026, n18027, n18028,
    n18029, n18030, n18031, n18032, n18033, n18034,
    n18035, n18036, n18037, n18038, n18039, n18040,
    n18041, n18042, n18043, n18044, n18045, n18046,
    n18047, n18048, n18049, n18050, n18051, n18052,
    n18053, n18054, n18055, n18056, n18057, n18058,
    n18059, n18060, n18061, n18062, n18063, n18064,
    n18065, n18066, n18067, n18068, n18069, n18070,
    n18071, n18072, n18073, n18074, n18075, n18076,
    n18077, n18078, n18079, n18080, n18081, n18082,
    n18083, n18084, n18085, n18086, n18087, n18088,
    n18089, n18090, n18091, n18092, n18093, n18094,
    n18095, n18096, n18097, n18098, n18099, n18100,
    n18101, n18102, n18103, n18104, n18105, n18106,
    n18107, n18108, n18109, n18110, n18111, n18112,
    n18113, n18114, n18115, n18116, n18117, n18118,
    n18119, n18120, n18121, n18122, n18123, n18124,
    n18125, n18126, n18127, n18128, n18129, n18130,
    n18131, n18132, n18133, n18134, n18135, n18136,
    n18137, n18138, n18139, n18140, n18141, n18142,
    n18143, n18144, n18145, n18146, n18147, n18148,
    n18149, n18150, n18151, n18152, n18153, n18154,
    n18155, n18156, n18157, n18158, n18159, n18160,
    n18161, n18162, n18163, n18164, n18165, n18166,
    n18167, n18168, n18169, n18170, n18171, n18172,
    n18173, n18174, n18175, n18176, n18177, n18178,
    n18179, n18180, n18181, n18182, n18183, n18184,
    n18185, n18186, n18187, n18188, n18189, n18190,
    n18191, n18192, n18193, n18194, n18195, n18196,
    n18197, n18198, n18199, n18200, n18201, n18202,
    n18203, n18204, n18205, n18206, n18207, n18208,
    n18209, n18210, n18211, n18212, n18213, n18214,
    n18215, n18216, n18217, n18218, n18219, n18220,
    n18221, n18222, n18223, n18224, n18225, n18226,
    n18227, n18228, n18229, n18230, n18231, n18232,
    n18233, n18234, n18235, n18236, n18237, n18238,
    n18239, n18240, n18241, n18242, n18243, n18244,
    n18245, n18246, n18247, n18248, n18249, n18250,
    n18251, n18252, n18253, n18254, n18255, n18256,
    n18257, n18258, n18259, n18260, n18261, n18262,
    n18263, n18264, n18265, n18266, n18267, n18268,
    n18269, n18270, n18271, n18272, n18273, n18274,
    n18275, n18276, n18277, n18278, n18279, n18280,
    n18281, n18282, n18283, n18284, n18285, n18286,
    n18287, n18288, n18289, n18290, n18291, n18292,
    n18293, n18294, n18295, n18296, n18297, n18298,
    n18299, n18300, n18301, n18302, n18303, n18304,
    n18305, n18306, n18307, n18308, n18309, n18310,
    n18311, n18312, n18313, n18314, n18315, n18316,
    n18317, n18318, n18319, n18320, n18321, n18322,
    n18323, n18324, n18325, n18326, n18328, n18329,
    n18330, n18331, n18332, n18333, n18334, n18335,
    n18336, n18337, n18338, n18339, n18340, n18341,
    n18342, n18343, n18344, n18345, n18346, n18347,
    n18348, n18349, n18350, n18351, n18352, n18353,
    n18354, n18355, n18356, n18357, n18358, n18359,
    n18360, n18361, n18362, n18363, n18364, n18365,
    n18366, n18367, n18368, n18369, n18370, n18371,
    n18372, n18373, n18374, n18375, n18376, n18377,
    n18378, n18379, n18380, n18381, n18382, n18383,
    n18384, n18385, n18386, n18387, n18388, n18389,
    n18390, n18391, n18392, n18393, n18394, n18395,
    n18396, n18397, n18398, n18399, n18400, n18401,
    n18402, n18403, n18404, n18405, n18406, n18407,
    n18408, n18409, n18410, n18411, n18412, n18413,
    n18414, n18415, n18416, n18417, n18418, n18419,
    n18420, n18421, n18422, n18423, n18424, n18425,
    n18426, n18427, n18428, n18429, n18430, n18431,
    n18432, n18433, n18434, n18435, n18436, n18437,
    n18438, n18439, n18440, n18441, n18442, n18443,
    n18444, n18445, n18446, n18447, n18448, n18449,
    n18450, n18451, n18452, n18453, n18454, n18455,
    n18456, n18457, n18458, n18459, n18460, n18461,
    n18462, n18463, n18464, n18465, n18466, n18467,
    n18468, n18469, n18470, n18471, n18472, n18473,
    n18474, n18475, n18476, n18477, n18478, n18479,
    n18480, n18481, n18482, n18483, n18484, n18485,
    n18486, n18487, n18488, n18489, n18490, n18491,
    n18492, n18493, n18494, n18495, n18496, n18497,
    n18498, n18499, n18500, n18501, n18502, n18503,
    n18504, n18505, n18506, n18507, n18508, n18509,
    n18510, n18511, n18512, n18513, n18514, n18515,
    n18516, n18517, n18518, n18519, n18520, n18521,
    n18522, n18523, n18524, n18525, n18526, n18527,
    n18528, n18529, n18530, n18531, n18532, n18533,
    n18534, n18535, n18536, n18537, n18538, n18539,
    n18540, n18541, n18542, n18543, n18544, n18545,
    n18546, n18547, n18548, n18549, n18550, n18551,
    n18552, n18553, n18554, n18555, n18556, n18557,
    n18558, n18559, n18560, n18561, n18562, n18563,
    n18564, n18565, n18566, n18567, n18568, n18569,
    n18570, n18571, n18572, n18573, n18574, n18575,
    n18576, n18577, n18578, n18579, n18580, n18581,
    n18582, n18583, n18584, n18585, n18586, n18587,
    n18588, n18589, n18590, n18591, n18592, n18593,
    n18594, n18595, n18596, n18597, n18598, n18599,
    n18600, n18601, n18602, n18603, n18604, n18605,
    n18606, n18607, n18608, n18609, n18610, n18611,
    n18612, n18613, n18614, n18615, n18616, n18617,
    n18618, n18619, n18620, n18621, n18622, n18623,
    n18624, n18625, n18626, n18627, n18628, n18629,
    n18630, n18631, n18632, n18633, n18634, n18635,
    n18636, n18637, n18638, n18639, n18640, n18641,
    n18642, n18643, n18644, n18645, n18646, n18647,
    n18648, n18649, n18650, n18651, n18652, n18653,
    n18654, n18655, n18656, n18657, n18658, n18659,
    n18660, n18661, n18662, n18663, n18664, n18665,
    n18666, n18667, n18668, n18669, n18670, n18671,
    n18672, n18673, n18674, n18675, n18676, n18677,
    n18678, n18679, n18680, n18681, n18682, n18683,
    n18684, n18685, n18686, n18687, n18688, n18689,
    n18690, n18691, n18692, n18693, n18694, n18695,
    n18696, n18697, n18698, n18699, n18700, n18701,
    n18702, n18703, n18704, n18705, n18706, n18707,
    n18708, n18709, n18710, n18711, n18712, n18713,
    n18714, n18715, n18716, n18717, n18718, n18719,
    n18720, n18721, n18722, n18723, n18724, n18725,
    n18726, n18727, n18728, n18729, n18730, n18731,
    n18732, n18733, n18734, n18735, n18736, n18737,
    n18738, n18739, n18740, n18741, n18742, n18743,
    n18744, n18745, n18746, n18747, n18748, n18749,
    n18750, n18751, n18752, n18753, n18754, n18755,
    n18756, n18757, n18758, n18759, n18760, n18761,
    n18762, n18763, n18764, n18765, n18766, n18767,
    n18768, n18769, n18770, n18771, n18772, n18773,
    n18774, n18775, n18776, n18777, n18778, n18779,
    n18780, n18781, n18782, n18783, n18784, n18785,
    n18786, n18787, n18788, n18789, n18790, n18791,
    n18792, n18793, n18794, n18795, n18796, n18797,
    n18798, n18799, n18800, n18801, n18802, n18803,
    n18804, n18805, n18806, n18807, n18808, n18809,
    n18810, n18811, n18812, n18813, n18814, n18815,
    n18816, n18817, n18818, n18819, n18820, n18821,
    n18822, n18823, n18824, n18825, n18826, n18827,
    n18828, n18829, n18830, n18831, n18832, n18833,
    n18834, n18835, n18836, n18837, n18838, n18839,
    n18841, n18842, n18843, n18844, n18845, n18846,
    n18847, n18848, n18849, n18850, n18851, n18852,
    n18853, n18854, n18855, n18856, n18857, n18858,
    n18859, n18860, n18861, n18862, n18863, n18864,
    n18865, n18866, n18867, n18868, n18869, n18870,
    n18871, n18872, n18873, n18874, n18875, n18876,
    n18877, n18878, n18879, n18880, n18881, n18882,
    n18883, n18884, n18885, n18886, n18887, n18888,
    n18889, n18890, n18891, n18892, n18893, n18894,
    n18895, n18896, n18897, n18898, n18899, n18900,
    n18901, n18902, n18903, n18904, n18905, n18906,
    n18907, n18908, n18909, n18910, n18911, n18912,
    n18913, n18914, n18915, n18916, n18917, n18918,
    n18919, n18920, n18921, n18922, n18923, n18924,
    n18925, n18926, n18927, n18928, n18929, n18930,
    n18931, n18932, n18933, n18934, n18935, n18936,
    n18937, n18938, n18939, n18940, n18941, n18942,
    n18943, n18944, n18945, n18946, n18947, n18948,
    n18949, n18950, n18951, n18952, n18953, n18954,
    n18955, n18956, n18957, n18958, n18959, n18960,
    n18961, n18962, n18963, n18964, n18965, n18966,
    n18967, n18968, n18969, n18970, n18971, n18972,
    n18973, n18974, n18975, n18976, n18977, n18978,
    n18979, n18980, n18981, n18982, n18983, n18984,
    n18985, n18986, n18987, n18988, n18989, n18990,
    n18991, n18992, n18993, n18994, n18995, n18996,
    n18997, n18998, n18999, n19000, n19001, n19002,
    n19003, n19004, n19005, n19006, n19007, n19008,
    n19009, n19010, n19011, n19012, n19013, n19014,
    n19015, n19016, n19017, n19018, n19019, n19020,
    n19021, n19022, n19023, n19024, n19025, n19026,
    n19027, n19028, n19029, n19030, n19031, n19032,
    n19033, n19034, n19035, n19036, n19037, n19038,
    n19039, n19040, n19041, n19042, n19043, n19044,
    n19045, n19046, n19047, n19048, n19049, n19050,
    n19051, n19052, n19053, n19054, n19055, n19056,
    n19057, n19058, n19059, n19060, n19061, n19062,
    n19063, n19064, n19065, n19066, n19067, n19068,
    n19069, n19070, n19071, n19072, n19073, n19074,
    n19075, n19076, n19077, n19078, n19079, n19080,
    n19081, n19082, n19083, n19084, n19085, n19086,
    n19087, n19088, n19089, n19090, n19091, n19092,
    n19093, n19094, n19095, n19096, n19097, n19098,
    n19099, n19100, n19101, n19102, n19103, n19104,
    n19105, n19106, n19107, n19108, n19109, n19110,
    n19111, n19112, n19113, n19114, n19115, n19116,
    n19117, n19118, n19119, n19120, n19121, n19122,
    n19123, n19124, n19125, n19126, n19127, n19128,
    n19129, n19130, n19131, n19132, n19133, n19134,
    n19135, n19136, n19137, n19138, n19139, n19140,
    n19141, n19142, n19143, n19144, n19145, n19146,
    n19147, n19148, n19149, n19150, n19151, n19152,
    n19153, n19154, n19155, n19156, n19157, n19158,
    n19159, n19160, n19161, n19162, n19163, n19164,
    n19165, n19166, n19167, n19168, n19169, n19170,
    n19171, n19172, n19173, n19174, n19175, n19176,
    n19177, n19178, n19179, n19180, n19181, n19182,
    n19183, n19184, n19185, n19186, n19187, n19188,
    n19189, n19190, n19191, n19192, n19193, n19194,
    n19195, n19196, n19197, n19198, n19199, n19200,
    n19201, n19202, n19203, n19204, n19205, n19206,
    n19207, n19208, n19209, n19210, n19211, n19212,
    n19213, n19214, n19215, n19216, n19217, n19218,
    n19219, n19220, n19221, n19222, n19223, n19224,
    n19225, n19226, n19227, n19228, n19229, n19230,
    n19231, n19232, n19233, n19234, n19235, n19236,
    n19237, n19238, n19239, n19240, n19241, n19242,
    n19243, n19244, n19245, n19246, n19247, n19248,
    n19249, n19250, n19251, n19252, n19253, n19254,
    n19255, n19256, n19257, n19258, n19259, n19260,
    n19261, n19262, n19263, n19264, n19265, n19266,
    n19267, n19268, n19269, n19270, n19271, n19272,
    n19273, n19274, n19275, n19276, n19277, n19278,
    n19279, n19280, n19281, n19282, n19283, n19284,
    n19285, n19286, n19287, n19288, n19289, n19290,
    n19291, n19292, n19293, n19294, n19295, n19296,
    n19297, n19298, n19299, n19300, n19301, n19302,
    n19303, n19304, n19305, n19306, n19307, n19308,
    n19309, n19310, n19311, n19312, n19313, n19314,
    n19315, n19316, n19317, n19318, n19319, n19320,
    n19321, n19322, n19323, n19324, n19325, n19326,
    n19327, n19328, n19329, n19330, n19331, n19332,
    n19333, n19334, n19335, n19336, n19337, n19338,
    n19339, n19341, n19342, n19343, n19344, n19345,
    n19346, n19347, n19348, n19349, n19350, n19351,
    n19352, n19353, n19354, n19355, n19356, n19357,
    n19358, n19359, n19360, n19361, n19362, n19363,
    n19364, n19365, n19366, n19367, n19368, n19369,
    n19370, n19371, n19372, n19373, n19374, n19375,
    n19376, n19377, n19378, n19379, n19380, n19381,
    n19382, n19383, n19384, n19385, n19386, n19387,
    n19388, n19389, n19390, n19391, n19392, n19393,
    n19394, n19395, n19396, n19397, n19398, n19399,
    n19400, n19401, n19402, n19403, n19404, n19405,
    n19406, n19407, n19408, n19409, n19410, n19411,
    n19412, n19413, n19414, n19415, n19416, n19417,
    n19418, n19419, n19420, n19421, n19422, n19423,
    n19424, n19425, n19426, n19427, n19428, n19429,
    n19430, n19431, n19432, n19433, n19434, n19435,
    n19436, n19437, n19438, n19439, n19440, n19441,
    n19442, n19443, n19444, n19445, n19446, n19447,
    n19448, n19449, n19450, n19451, n19452, n19453,
    n19454, n19455, n19456, n19457, n19458, n19459,
    n19460, n19461, n19462, n19463, n19464, n19465,
    n19466, n19467, n19468, n19469, n19470, n19471,
    n19472, n19473, n19474, n19475, n19476, n19477,
    n19478, n19479, n19480, n19481, n19482, n19483,
    n19484, n19485, n19486, n19487, n19488, n19489,
    n19490, n19491, n19492, n19493, n19494, n19495,
    n19496, n19497, n19498, n19499, n19500, n19501,
    n19502, n19503, n19504, n19505, n19506, n19507,
    n19508, n19509, n19510, n19511, n19512, n19513,
    n19514, n19515, n19516, n19517, n19518, n19519,
    n19520, n19521, n19522, n19523, n19524, n19525,
    n19526, n19527, n19528, n19529, n19530, n19531,
    n19532, n19533, n19534, n19535, n19536, n19537,
    n19538, n19539, n19540, n19541, n19542, n19543,
    n19544, n19545, n19546, n19547, n19548, n19549,
    n19550, n19551, n19552, n19553, n19554, n19555,
    n19556, n19557, n19558, n19559, n19560, n19561,
    n19562, n19563, n19564, n19565, n19566, n19567,
    n19568, n19569, n19570, n19571, n19572, n19573,
    n19574, n19575, n19576, n19577, n19578, n19579,
    n19580, n19581, n19582, n19583, n19584, n19585,
    n19586, n19587, n19588, n19589, n19590, n19591,
    n19592, n19593, n19594, n19595, n19596, n19597,
    n19598, n19599, n19600, n19601, n19602, n19603,
    n19604, n19605, n19606, n19607, n19608, n19609,
    n19610, n19611, n19612, n19613, n19614, n19615,
    n19616, n19617, n19618, n19619, n19620, n19621,
    n19622, n19623, n19624, n19625, n19626, n19627,
    n19628, n19629, n19630, n19631, n19632, n19633,
    n19634, n19635, n19636, n19637, n19638, n19639,
    n19640, n19641, n19642, n19643, n19644, n19645,
    n19646, n19647, n19648, n19649, n19650, n19651,
    n19652, n19653, n19654, n19655, n19656, n19657,
    n19658, n19659, n19660, n19661, n19662, n19663,
    n19664, n19665, n19666, n19667, n19668, n19669,
    n19670, n19671, n19672, n19673, n19674, n19675,
    n19676, n19677, n19678, n19679, n19680, n19681,
    n19682, n19683, n19684, n19685, n19686, n19687,
    n19688, n19689, n19690, n19691, n19692, n19693,
    n19694, n19695, n19696, n19697, n19698, n19699,
    n19700, n19701, n19702, n19703, n19704, n19705,
    n19706, n19707, n19708, n19709, n19710, n19711,
    n19712, n19713, n19714, n19715, n19716, n19717,
    n19718, n19719, n19720, n19721, n19722, n19723,
    n19724, n19725, n19726, n19727, n19728, n19729,
    n19730, n19731, n19732, n19733, n19734, n19735,
    n19736, n19737, n19738, n19739, n19740, n19741,
    n19742, n19743, n19744, n19745, n19746, n19747,
    n19748, n19749, n19750, n19751, n19752, n19753,
    n19754, n19755, n19756, n19757, n19758, n19759,
    n19760, n19761, n19762, n19763, n19764, n19765,
    n19766, n19767, n19768, n19769, n19770, n19771,
    n19772, n19773, n19774, n19775, n19776, n19777,
    n19778, n19779, n19780, n19781, n19782, n19783,
    n19784, n19785, n19786, n19787, n19788, n19789,
    n19790, n19791, n19792, n19793, n19794, n19796,
    n19797, n19798, n19799, n19800, n19801, n19802,
    n19803, n19804, n19805, n19806, n19807, n19808,
    n19809, n19810, n19811, n19812, n19813, n19814,
    n19815, n19816, n19817, n19818, n19819, n19820,
    n19821, n19822, n19823, n19824, n19825, n19826,
    n19827, n19828, n19829, n19830, n19831, n19832,
    n19833, n19834, n19835, n19836, n19837, n19838,
    n19839, n19840, n19841, n19842, n19843, n19844,
    n19845, n19846, n19847, n19848, n19849, n19850,
    n19851, n19852, n19853, n19854, n19855, n19856,
    n19857, n19858, n19859, n19860, n19861, n19862,
    n19863, n19864, n19865, n19867, n19868, n19869,
    n19870, n19871, n19872, n19873, n19874, n19875,
    n19876, n19877, n19878, n19879, n19880, n19881,
    n19882, n19883, n19884, n19885, n19886, n19887,
    n19888, n19889, n19890, n19891, n19892, n19893,
    n19894, n19895, n19896, n19897, n19898, n19899,
    n19900, n19901, n19902, n19903, n19904, n19905,
    n19906, n19907, n19908, n19909, n19910, n19911,
    n19912, n19913, n19914, n19915, n19916, n19917,
    n19918, n19919, n19920, n19921, n19922, n19923,
    n19924, n19925, n19926, n19927, n19928, n19929,
    n19930, n19931, n19932, n19933, n19934, n19935,
    n19936, n19937, n19938, n19939, n19940, n19941,
    n19942, n19943, n19944, n19945, n19946, n19947,
    n19948, n19949, n19950, n19951, n19952, n19953,
    n19954, n19955, n19956, n19957, n19958, n19959,
    n19960, n19961, n19962, n19963, n19964, n19965,
    n19966, n19967, n19968, n19969, n19970, n19971,
    n19972, n19973, n19974, n19975, n19976, n19977,
    n19978, n19979, n19980, n19981, n19982, n19983,
    n19984, n19985, n19986, n19987, n19988, n19989,
    n19990, n19991, n19992, n19993, n19994, n19995,
    n19996, n19997, n19998, n19999, n20000, n20001,
    n20002, n20004, n20005, n20006, n20007, n20008,
    n20009, n20010, n20011, n20012, n20013, n20014,
    n20015, n20016, n20017, n20018, n20019, n20020,
    n20021, n20022, n20023, n20024, n20025, n20026,
    n20027, n20028, n20029, n20030, n20031, n20032,
    n20033, n20034, n20035, n20036, n20037, n20038,
    n20039, n20040, n20041, n20042, n20043, n20044,
    n20045, n20046, n20047, n20048, n20049, n20050,
    n20051, n20052, n20053, n20054, n20055, n20056,
    n20057, n20058, n20059, n20060, n20061, n20062,
    n20063, n20064, n20065, n20066, n20068, n20069,
    n20070, n20071, n20072, n20073, n20074, n20075,
    n20076, n20077, n20078, n20079, n20080, n20081,
    n20082, n20083, n20084, n20085, n20086, n20087,
    n20088, n20089, n20090, n20091, n20092, n20093,
    n20094, n20095, n20096, n20097, n20098, n20099,
    n20100, n20101, n20102, n20103, n20104, n20105,
    n20106, n20107, n20108, n20109, n20110, n20111,
    n20112, n20113, n20114, n20115, n20116, n20117,
    n20118, n20119, n20120, n20121, n20122, n20123,
    n20125, n20126, n20127, n20128, n20129, n20130,
    n20131, n20132, n20133, n20134, n20135, n20136,
    n20137, n20138, n20139, n20140, n20141, n20142,
    n20143, n20144, n20145, n20146, n20147, n20148,
    n20149, n20150, n20151, n20152, n20153, n20154,
    n20155, n20156, n20157, n20158, n20159, n20160,
    n20161, n20162, n20163, n20164, n20165, n20166,
    n20167, n20168, n20169, n20170, n20171, n20172,
    n20173, n20174, n20175, n20176, n20177, n20178,
    n20180, n20181, n20182, n20183, n20184, n20185,
    n20186, n20187, n20188, n20189, n20190, n20191,
    n20192, n20193, n20194, n20195, n20196, n20197,
    n20198, n20199, n20200, n20201, n20202, n20203,
    n20204, n20205, n20206, n20207, n20208, n20209,
    n20210, n20211, n20212, n20213, n20214, n20215,
    n20216, n20217, n20218, n20219, n20220, n20221,
    n20222, n20223, n20224, n20225, n20226, n20227,
    n20228, n20229, n20230, n20231, n20232, n20233,
    n20234, n20235, n20236, n20237, n20238, n20239,
    n20240, n20241, n20242, n20243, n20244, n20245,
    n20246, n20247, n20248, n20249, n20250, n20251,
    n20252, n20253, n20254, n20255, n20256, n20257,
    n20259, n20260, n20261, n20262, n20263, n20264,
    n20265, n20266, n20267, n20268, n20269, n20270,
    n20271, n20272, n20273, n20274, n20275, n20276,
    n20277, n20278, n20279, n20280, n20281, n20282,
    n20283, n20284, n20285, n20286, n20287, n20288,
    n20289, n20290, n20291, n20292, n20293, n20294,
    n20295, n20296, n20297, n20298, n20299, n20300,
    n20301, n20302, n20303, n20304, n20305, n20306,
    n20307, n20308, n20309, n20310, n20311, n20312,
    n20313, n20314, n20315, n20316, n20317, n20318,
    n20319, n20320, n20321, n20322, n20323, n20324,
    n20325, n20326, n20327, n20328, n20329, n20330,
    n20331, n20332, n20333, n20334, n20335, n20336,
    n20337, n20338, n20339, n20340, n20341, n20342,
    n20343, n20344, n20345, n20346, n20347, n20348,
    n20349, n20350, n20351, n20352, n20353, n20354,
    n20355, n20356, n20357, n20358, n20359, n20360,
    n20361, n20363, n20364, n20365, n20366, n20367,
    n20368, n20369, n20370, n20371, n20372, n20373,
    n20374, n20375, n20376, n20377, n20378, n20379,
    n20380, n20381, n20382, n20383, n20384, n20385,
    n20386, n20387, n20388, n20389, n20390, n20391,
    n20392, n20393, n20394, n20395, n20396, n20397,
    n20398, n20399, n20400, n20401, n20402, n20403,
    n20404, n20405, n20406, n20407, n20408, n20409,
    n20410, n20411, n20412, n20413, n20414, n20415,
    n20416, n20417, n20418, n20419, n20420, n20421,
    n20422, n20423, n20424, n20425, n20426, n20427,
    n20428, n20429, n20430, n20431, n20432, n20433,
    n20434, n20435, n20436, n20437, n20438, n20439,
    n20440, n20442, n20443, n20444, n20445, n20446,
    n20447, n20448, n20449, n20450, n20451, n20452,
    n20453, n20454, n20455, n20456, n20457, n20458,
    n20459, n20460, n20461, n20462, n20463, n20464,
    n20465, n20466, n20467, n20468, n20469, n20470,
    n20471, n20472, n20473, n20474, n20475, n20476,
    n20477, n20478, n20479, n20480, n20481, n20482,
    n20483, n20484, n20485, n20486, n20487, n20488,
    n20489, n20490, n20491, n20492, n20494, n20495,
    n20496, n20497, n20498, n20499, n20500, n20501,
    n20502, n20503, n20504, n20505, n20506, n20507,
    n20508, n20509, n20510, n20511, n20512, n20513,
    n20514, n20515, n20516, n20517, n20518, n20519,
    n20520, n20521, n20522, n20523, n20524, n20525,
    n20526, n20527, n20528, n20529, n20530, n20531,
    n20532, n20533, n20535, n20536, n20537, n20538,
    n20539, n20540, n20541, n20542, n20543, n20544,
    n20545, n20546, n20547, n20548, n20549, n20550,
    n20551, n20552, n20553, n20554, n20555, n20556,
    n20557, n20558, n20559, n20560, n20561, n20562,
    n20563, n20565, n20566, n20567, n20568, n20569,
    n20570, n20571, n20572, n20573, n20574, n20575,
    n20576, n20577, n20578, n20579, n20580, n20581,
    n20582, n20583, n20584, n20585, n20586, n20587,
    n20588, n20589, n20590, n20591, n20592, n20593,
    n20594, n20595, n20596, n20597, n20598, n20599,
    n20600, n20601, n20602, n20603, n20604, n20605,
    n20606, n20607, n20608, n20609, n20610, n20611,
    n20612, n20613, n20614, n20615, n20616, n20617,
    n20618, n20619, n20621, n20622, n20623, n20624,
    n20625, n20626, n20627, n20628, n20629, n20630,
    n20631, n20632, n20633, n20634, n20635, n20636,
    n20637, n20638, n20639, n20640, n20641, n20642,
    n20643, n20644, n20645, n20646, n20647, n20648,
    n20649, n20650, n20651, n20652, n20653, n20654,
    n20655, n20656, n20657, n20658, n20659, n20660,
    n20661, n20662, n20663, n20664, n20665, n20666,
    n20667, n20668, n20669, n20670, n20671, n20672,
    n20673, n20674, n20676, n20677, n20678, n20679,
    n20680, n20681, n20682, n20683, n20684, n20685,
    n20686, n20687, n20688, n20689, n20690, n20691,
    n20692, n20693, n20694, n20695, n20696, n20697,
    n20698, n20699, n20700, n20701, n20702, n20703,
    n20704, n20705, n20706, n20707, n20708, n20709,
    n20710, n20711, n20712, n20713, n20714, n20715,
    n20716, n20717, n20718, n20719, n20720, n20721,
    n20722, n20723, n20724, n20725, n20726, n20727,
    n20728, n20729, n20731, n20732, n20733, n20734,
    n20735, n20736, n20737, n20738, n20739, n20740,
    n20741, n20742, n20743, n20744, n20745, n20746,
    n20747, n20748, n20749, n20750, n20751, n20752,
    n20753, n20754, n20755, n20756, n20757, n20758,
    n20759, n20760, n20761, n20762, n20763, n20764,
    n20765, n20766, n20767, n20768, n20769, n20770,
    n20771, n20772, n20773, n20774, n20775, n20776,
    n20777, n20778, n20779, n20780, n20781, n20782,
    n20783, n20784, n20785, n20786, n20787, n20789,
    n20790, n20791, n20792, n20793, n20794, n20795,
    n20796, n20797, n20798, n20799, n20800, n20801,
    n20802, n20803, n20804, n20805, n20806, n20807,
    n20808, n20809, n20810, n20811, n20812, n20813,
    n20814, n20815, n20816, n20817, n20818, n20819,
    n20820, n20821, n20822, n20823, n20824, n20825,
    n20826, n20827, n20828, n20829, n20830, n20831,
    n20832, n20833, n20834, n20835, n20836, n20837,
    n20838, n20839, n20840, n20841, n20842, n20843,
    n20844, n20845, n20846, n20847, n20848, n20849,
    n20850, n20851, n20852, n20853, n20854, n20855,
    n20856, n20857, n20858, n20859, n20860, n20861,
    n20862, n20863, n20864, n20865, n20866, n20867,
    n20868, n20869, n20870, n20871, n20872, n20873,
    n20874, n20875, n20876, n20877, n20878, n20879,
    n20881, n20882, n20883, n20884, n20885, n20886,
    n20887, n20888, n20889, n20890, n20891, n20892,
    n20893, n20894, n20895, n20896, n20897, n20898,
    n20899, n20900, n20901, n20902, n20903, n20904,
    n20905, n20906, n20907, n20908, n20909, n20910,
    n20911, n20912, n20913, n20914, n20915, n20916,
    n20917, n20918, n20919, n20920, n20921, n20922,
    n20923, n20924, n20925, n20926, n20927, n20928,
    n20929, n20930, n20931, n20932, n20933, n20935,
    n20936, n20937, n20938, n20939, n20940, n20941,
    n20942, n20943, n20944, n20945, n20946, n20947,
    n20948, n20949, n20950, n20951, n20952, n20953,
    n20954, n20955, n20956, n20957, n20958, n20959,
    n20960, n20961, n20962, n20963, n20964, n20965,
    n20966, n20967, n20968, n20969, n20970, n20971,
    n20972, n20973, n20974, n20975, n20976, n20977,
    n20978, n20979, n20980, n20981, n20982, n20983,
    n20984, n20985, n20986, n20987, n20988, n20989,
    n20990, n20992, n20993, n20994, n20995, n20996,
    n20997, n20998, n20999, n21000, n21001, n21002,
    n21003, n21004, n21005, n21006, n21007, n21008,
    n21009, n21010, n21011, n21012, n21013, n21014,
    n21015, n21016, n21017, n21018, n21019, n21020,
    n21021, n21022, n21023, n21024, n21025, n21026,
    n21027, n21028, n21029, n21030, n21032, n21033,
    n21034, n21035, n21036, n21037, n21038, n21039,
    n21040, n21041, n21042, n21043, n21044, n21045,
    n21046, n21047, n21048, n21049, n21050, n21051,
    n21052, n21053, n21054, n21055, n21056, n21057,
    n21058, n21059, n21060, n21061, n21062, n21063,
    n21064, n21065, n21066, n21067, n21068, n21069,
    n21070, n21072, n21073, n21074, n21075, n21076,
    n21077, n21078, n21079, n21080, n21081, n21082,
    n21083, n21084, n21085, n21086, n21087, n21088,
    n21089, n21090, n21091, n21092, n21093, n21094,
    n21095, n21096, n21097, n21098, n21099, n21100,
    n21101, n21102, n21103, n21104, n21105, n21106,
    n21107, n21108, n21109, n21110, n21111, n21112,
    n21113, n21114, n21115, n21116, n21117, n21118,
    n21119, n21120, n21121, n21122, n21123, n21124,
    n21125, n21126, n21127, n21128, n21129, n21130,
    n21131, n21132, n21133, n21134, n21135, n21136,
    n21137, n21138, n21139, n21140, n21141, n21142,
    n21143, n21144, n21145, n21146, n21147, n21148,
    n21149, n21150, n21151, n21152, n21153, n21154,
    n21155, n21156, n21157, n21158, n21159, n21160,
    n21161, n21162, n21163, n21164, n21165, n21167,
    n21168, n21169, n21170, n21171, n21172, n21173,
    n21174, n21175, n21176, n21177, n21178, n21179,
    n21180, n21181, n21182, n21183, n21184, n21185,
    n21186, n21187, n21188, n21189, n21190, n21191,
    n21192, n21193, n21194, n21195, n21196, n21197,
    n21198, n21199, n21200, n21201, n21202, n21203,
    n21204, n21205, n21206, n21207, n21208, n21210,
    n21211, n21212, n21213, n21214, n21215, n21216,
    n21217, n21218, n21219, n21220, n21221, n21222,
    n21223, n21224, n21225, n21226, n21227, n21228,
    n21229, n21230, n21231, n21232, n21233, n21234,
    n21235, n21236, n21237, n21238, n21239, n21240,
    n21241, n21242, n21243, n21244, n21245, n21246,
    n21247, n21248, n21249, n21250, n21251, n21252,
    n21253, n21254, n21255, n21256, n21257, n21258,
    n21259, n21260, n21261, n21262, n21263, n21264,
    n21265, n21266, n21267, n21268, n21269, n21270,
    n21271, n21272, n21273, n21274, n21275, n21276,
    n21277, n21278, n21279, n21280, n21281, n21282,
    n21283, n21284, n21285, n21286, n21287, n21289,
    n21290, n21291, n21292, n21293, n21294, n21295,
    n21296, n21297, n21298, n21299, n21300, n21301,
    n21302, n21303, n21304, n21305, n21306, n21307,
    n21308, n21309, n21310, n21311, n21312, n21313,
    n21314, n21315, n21316, n21317, n21318, n21319,
    n21320, n21321, n21322, n21323, n21324, n21325,
    n21326, n21327, n21328, n21329, n21330, n21331,
    n21332, n21333, n21334, n21335, n21336, n21337,
    n21338, n21339, n21340, n21341, n21342, n21343,
    n21344, n21345, n21346, n21347, n21348, n21349,
    n21350, n21351, n21352, n21353, n21354, n21355,
    n21356, n21357, n21358, n21359, n21360, n21361,
    n21362, n21363, n21364, n21365, n21366, n21368,
    n21369, n21370, n21371, n21372, n21373, n21374,
    n21375, n21376, n21377, n21378, n21379, n21380,
    n21381, n21382, n21383, n21384, n21385, n21386,
    n21387, n21388, n21389, n21390, n21391, n21392,
    n21393, n21394, n21395, n21396, n21397, n21398,
    n21399, n21400, n21401, n21402, n21403, n21404,
    n21405, n21406, n21407, n21408, n21409, n21410,
    n21411, n21412, n21413, n21414, n21415, n21416,
    n21417, n21418, n21419, n21420, n21421, n21422,
    n21423, n21424, n21425, n21426, n21427, n21428,
    n21429, n21430, n21431, n21432, n21433, n21434,
    n21435, n21436, n21437, n21438, n21439, n21440,
    n21441, n21442, n21443, n21444, n21445, n21447,
    n21448, n21449, n21450, n21451, n21452, n21453,
    n21454, n21455, n21456, n21457, n21458, n21459,
    n21460, n21461, n21462, n21463, n21464, n21465,
    n21466, n21467, n21468, n21469, n21470, n21471,
    n21472, n21473, n21474, n21475, n21476, n21477,
    n21478, n21479, n21480, n21481, n21482, n21483,
    n21484, n21485, n21486, n21487, n21488, n21489,
    n21490, n21491, n21492, n21493, n21494, n21495,
    n21496, n21497, n21498, n21499, n21500, n21501,
    n21502, n21503, n21504, n21505, n21506, n21507,
    n21508, n21509, n21510, n21511, n21512, n21513,
    n21514, n21515, n21516, n21517, n21518, n21519,
    n21520, n21521, n21522, n21523, n21524, n21526,
    n21527, n21528, n21529, n21530, n21531, n21532,
    n21533, n21534, n21535, n21536, n21537, n21538,
    n21539, n21540, n21541, n21542, n21543, n21544,
    n21545, n21546, n21547, n21548, n21549, n21550,
    n21551, n21552, n21553, n21554, n21555, n21556,
    n21557, n21558, n21559, n21560, n21561, n21562,
    n21563, n21564, n21565, n21566, n21567, n21568,
    n21569, n21570, n21571, n21572, n21573, n21574,
    n21575, n21576, n21577, n21578, n21579, n21580,
    n21581, n21582, n21583, n21584, n21585, n21586,
    n21587, n21588, n21589, n21590, n21591, n21592,
    n21593, n21594, n21595, n21596, n21597, n21598,
    n21599, n21600, n21601, n21602, n21603, n21605,
    n21606, n21607, n21608, n21609, n21610, n21611,
    n21612, n21613, n21614, n21615, n21616, n21617,
    n21618, n21619, n21620, n21621, n21622, n21623,
    n21624, n21625, n21626, n21627, n21628, n21629,
    n21630, n21631, n21632, n21633, n21634, n21635,
    n21636, n21637, n21638, n21639, n21640, n21641,
    n21642, n21643, n21644, n21645, n21646, n21647,
    n21648, n21649, n21650, n21651, n21652, n21653,
    n21654, n21655, n21656, n21657, n21658, n21659,
    n21660, n21661, n21662, n21663, n21664, n21665,
    n21666, n21667, n21668, n21669, n21670, n21671,
    n21672, n21673, n21674, n21675, n21676, n21677,
    n21678, n21679, n21680, n21681, n21682, n21683,
    n21684, n21685, n21686, n21687, n21688, n21689,
    n21690, n21691, n21692, n21693, n21694, n21695,
    n21696, n21697, n21698, n21699, n21700, n21701,
    n21702, n21703, n21704, n21705, n21706, n21707,
    n21708, n21709, n21710, n21711, n21712, n21713,
    n21714, n21715, n21716, n21717, n21718, n21719,
    n21720, n21721, n21722, n21723, n21724, n21725,
    n21726, n21727, n21728, n21729, n21730, n21731,
    n21732, n21733, n21734, n21735, n21736, n21737,
    n21738, n21739, n21740, n21741, n21742, n21743,
    n21744, n21745, n21746, n21747, n21748, n21749,
    n21750, n21751, n21752, n21753, n21754, n21755,
    n21756, n21757, n21758, n21759, n21760, n21761,
    n21762, n21763, n21764, n21765, n21766, n21767,
    n21768, n21769, n21770, n21771, n21772, n21773,
    n21774, n21775, n21776, n21777, n21778, n21779,
    n21780, n21781, n21782, n21783, n21784, n21785,
    n21786, n21787, n21788, n21789, n21790, n21791,
    n21792, n21793, n21794, n21795, n21796, n21797,
    n21798, n21799, n21800, n21801, n21802, n21803,
    n21804, n21805, n21806, n21807, n21808, n21809,
    n21810, n21811, n21812, n21813, n21814, n21815,
    n21816, n21817, n21818, n21819, n21820, n21821,
    n21822, n21823, n21824, n21825, n21826, n21827,
    n21828, n21829, n21830, n21831, n21832, n21833,
    n21834, n21835, n21836, n21837, n21838, n21839,
    n21840, n21841, n21842, n21843, n21844, n21845,
    n21846, n21847, n21848, n21849, n21850, n21851,
    n21852, n21853, n21854, n21855, n21856, n21857,
    n21858, n21859, n21860, n21861, n21862, n21863,
    n21864, n21865, n21866, n21867, n21868, n21869,
    n21870, n21871, n21872, n21873, n21874, n21875,
    n21876, n21877, n21878, n21879, n21880, n21881,
    n21882, n21883, n21884, n21885, n21886, n21887,
    n21888, n21889, n21890, n21891, n21892, n21893,
    n21894, n21895, n21896, n21897, n21898, n21899,
    n21900, n21901, n21902, n21903, n21904, n21905,
    n21906, n21907, n21908, n21909, n21910, n21911,
    n21912, n21913, n21914, n21915, n21916, n21917,
    n21918, n21919, n21920, n21921, n21922, n21923,
    n21924, n21925, n21926, n21927, n21928, n21929,
    n21930, n21931, n21932, n21933, n21934, n21935,
    n21936, n21937, n21938, n21939, n21940, n21941,
    n21942, n21943, n21944, n21945, n21946, n21947,
    n21948, n21949, n21950, n21951, n21952, n21953,
    n21954, n21955, n21956, n21957, n21958, n21959,
    n21960, n21961, n21962, n21963, n21964, n21965,
    n21966, n21967, n21968, n21969, n21970, n21971,
    n21972, n21973, n21974, n21975, n21976, n21977,
    n21978, n21979, n21980, n21981, n21982, n21983,
    n21984, n21985, n21986, n21987, n21988, n21989,
    n21990, n21991, n21992, n21993, n21994, n21995,
    n21996, n21997, n21998, n21999, n22000, n22001,
    n22002, n22003, n22004, n22005, n22006, n22007,
    n22008, n22009, n22010, n22011, n22012, n22013,
    n22014, n22015, n22016, n22017, n22018, n22019,
    n22020, n22021, n22022, n22023, n22024, n22025,
    n22026, n22027, n22028, n22029, n22030, n22031,
    n22032, n22033, n22034, n22035, n22036, n22037,
    n22038, n22039, n22040, n22041, n22042, n22043,
    n22044, n22046, n22047, n22048, n22049, n22050,
    n22051, n22052, n22053, n22054, n22055, n22056,
    n22057, n22058, n22059, n22060, n22061, n22062,
    n22063, n22064, n22065, n22066, n22067, n22068,
    n22069, n22070, n22071, n22072, n22073, n22074,
    n22075, n22076, n22077, n22078, n22079, n22080,
    n22081, n22082, n22083, n22084, n22085, n22086,
    n22087, n22088, n22089, n22090, n22091, n22092,
    n22093, n22094, n22095, n22096, n22097, n22098,
    n22099, n22100, n22101, n22102, n22103, n22104,
    n22105, n22106, n22107, n22108, n22109, n22110,
    n22111, n22112, n22113, n22114, n22115, n22116,
    n22117, n22118, n22119, n22120, n22121, n22122,
    n22123, n22124, n22125, n22126, n22127, n22128,
    n22129, n22130, n22131, n22132, n22133, n22134,
    n22135, n22136, n22137, n22138, n22139, n22140,
    n22141, n22142, n22143, n22144, n22145, n22146,
    n22147, n22148, n22149, n22150, n22151, n22152,
    n22153, n22154, n22155, n22156, n22157, n22158,
    n22159, n22160, n22161, n22162, n22163, n22164,
    n22165, n22166, n22167, n22168, n22169, n22170,
    n22171, n22172, n22173, n22174, n22175, n22176,
    n22177, n22178, n22179, n22180, n22181, n22182,
    n22183, n22184, n22185, n22186, n22187, n22188,
    n22189, n22190, n22191, n22192, n22193, n22194,
    n22195, n22196, n22197, n22198, n22199, n22200,
    n22201, n22202, n22203, n22204, n22205, n22206,
    n22207, n22208, n22209, n22210, n22211, n22212,
    n22213, n22214, n22215, n22216, n22217, n22218,
    n22219, n22220, n22221, n22222, n22223, n22224,
    n22225, n22226, n22227, n22228, n22229, n22230,
    n22231, n22232, n22233, n22234, n22235, n22236,
    n22237, n22238, n22239, n22240, n22241, n22242,
    n22243, n22244, n22245, n22246, n22247, n22248,
    n22249, n22250, n22251, n22252, n22253, n22254,
    n22255, n22256, n22257, n22258, n22259, n22260,
    n22261, n22262, n22263, n22264, n22265, n22266,
    n22267, n22268, n22269, n22270, n22271, n22272,
    n22273, n22274, n22275, n22276, n22277, n22278,
    n22279, n22280, n22281, n22282, n22283, n22284,
    n22285, n22286, n22287, n22288, n22289, n22290,
    n22291, n22292, n22293, n22294, n22295, n22296,
    n22297, n22298, n22299, n22300, n22301, n22302,
    n22303, n22304, n22305, n22306, n22307, n22308,
    n22309, n22310, n22311, n22312, n22313, n22314,
    n22315, n22316, n22317, n22318, n22319, n22320,
    n22321, n22322, n22323, n22324, n22325, n22326,
    n22327, n22328, n22329, n22330, n22331, n22332,
    n22333, n22334, n22335, n22336, n22337, n22338,
    n22339, n22340, n22341, n22342, n22343, n22344,
    n22345, n22346, n22347, n22348, n22349, n22350,
    n22351, n22352, n22353, n22354, n22355, n22356,
    n22357, n22358, n22359, n22360, n22361, n22362,
    n22363, n22364, n22365, n22366, n22367, n22368,
    n22369, n22370, n22371, n22372, n22373, n22374,
    n22375, n22376, n22377, n22378, n22379, n22380,
    n22381, n22382, n22383, n22384, n22385, n22386,
    n22387, n22388, n22389, n22390, n22391, n22392,
    n22393, n22394, n22395, n22396, n22397, n22398,
    n22399, n22400, n22401, n22402, n22403, n22404,
    n22405, n22406, n22407, n22408, n22409, n22410,
    n22411, n22412, n22413, n22414, n22415, n22416,
    n22417, n22418, n22419, n22420, n22421, n22422,
    n22423, n22424, n22425, n22426, n22427, n22428,
    n22429, n22430, n22431, n22432, n22433, n22434,
    n22435, n22436, n22437, n22438, n22439, n22440,
    n22441, n22442, n22443, n22444, n22445, n22446,
    n22447, n22448, n22449, n22450, n22451, n22452,
    n22453, n22454, n22455, n22456, n22457, n22458,
    n22459, n22460, n22461, n22462, n22463, n22464,
    n22465, n22466, n22467, n22468, n22469, n22470,
    n22471, n22472, n22473, n22474, n22475, n22476,
    n22477, n22478, n22479, n22480, n22481, n22482,
    n22483, n22484, n22485, n22486, n22487, n22488,
    n22489, n22490, n22491, n22492, n22493, n22494,
    n22495, n22496, n22497, n22498, n22499, n22500,
    n22501, n22502, n22504, n22505, n22506, n22507,
    n22508, n22509, n22510, n22511, n22512, n22513,
    n22514, n22515, n22516, n22517, n22518, n22519,
    n22520, n22521, n22522, n22523, n22524, n22525,
    n22526, n22527, n22528, n22529, n22530, n22531,
    n22532, n22533, n22534, n22535, n22536, n22537,
    n22538, n22539, n22540, n22541, n22542, n22543,
    n22544, n22545, n22546, n22547, n22548, n22549,
    n22550, n22551, n22552, n22553, n22554, n22555,
    n22556, n22557, n22558, n22559, n22560, n22561,
    n22562, n22563, n22564, n22565, n22566, n22567,
    n22568, n22569, n22570, n22571, n22572, n22573,
    n22574, n22575, n22576, n22577, n22578, n22579,
    n22580, n22581, n22582, n22583, n22584, n22585,
    n22586, n22587, n22588, n22589, n22590, n22591,
    n22592, n22593, n22594, n22595, n22596, n22597,
    n22598, n22599, n22600, n22601, n22602, n22603,
    n22604, n22605, n22606, n22607, n22608, n22609,
    n22610, n22611, n22612, n22613, n22614, n22615,
    n22616, n22617, n22618, n22619, n22620, n22621,
    n22622, n22623, n22624, n22625, n22626, n22627,
    n22628, n22629, n22630, n22631, n22632, n22633,
    n22634, n22635, n22636, n22637, n22638, n22639,
    n22640, n22641, n22642, n22643, n22644, n22645,
    n22646, n22647, n22648, n22649, n22650, n22651,
    n22652, n22653, n22654, n22655, n22656, n22657,
    n22658, n22659, n22660, n22661, n22662, n22663,
    n22664, n22665, n22666, n22667, n22668, n22669,
    n22670, n22671, n22672, n22673, n22674, n22675,
    n22676, n22677, n22678, n22679, n22680, n22681,
    n22682, n22683, n22684, n22685, n22686, n22687,
    n22688, n22689, n22690, n22691, n22692, n22693,
    n22694, n22695, n22696, n22697, n22698, n22699,
    n22700, n22701, n22702, n22703, n22704, n22705,
    n22706, n22707, n22708, n22709, n22710, n22711,
    n22712, n22713, n22714, n22715, n22716, n22717,
    n22718, n22719, n22720, n22721, n22722, n22723,
    n22724, n22725, n22726, n22727, n22728, n22729,
    n22730, n22731, n22732, n22733, n22734, n22735,
    n22736, n22737, n22738, n22739, n22740, n22741,
    n22742, n22743, n22744, n22745, n22746, n22747,
    n22748, n22749, n22750, n22751, n22752, n22753,
    n22754, n22755, n22756, n22757, n22758, n22759,
    n22760, n22761, n22762, n22763, n22764, n22765,
    n22766, n22767, n22768, n22769, n22770, n22771,
    n22772, n22773, n22774, n22775, n22776, n22777,
    n22778, n22779, n22780, n22781, n22782, n22783,
    n22784, n22785, n22786, n22787, n22788, n22789,
    n22790, n22791, n22792, n22793, n22794, n22795,
    n22796, n22797, n22798, n22799, n22800, n22801,
    n22802, n22803, n22804, n22805, n22806, n22807,
    n22808, n22809, n22810, n22811, n22812, n22813,
    n22814, n22815, n22816, n22817, n22818, n22819,
    n22820, n22821, n22822, n22823, n22824, n22825,
    n22826, n22827, n22828, n22829, n22830, n22831,
    n22832, n22833, n22834, n22835, n22836, n22837,
    n22838, n22839, n22840, n22841, n22842, n22843,
    n22844, n22845, n22846, n22847, n22848, n22849,
    n22850, n22851, n22852, n22853, n22854, n22855,
    n22856, n22857, n22858, n22859, n22860, n22861,
    n22862, n22863, n22864, n22865, n22866, n22867,
    n22868, n22869, n22870, n22871, n22872, n22873,
    n22874, n22875, n22876, n22877, n22878, n22879,
    n22880, n22881, n22882, n22883, n22884, n22885,
    n22886, n22887, n22888, n22889, n22890, n22891,
    n22892, n22893, n22894, n22895, n22896, n22897,
    n22898, n22899, n22900, n22901, n22902, n22903,
    n22904, n22905, n22906, n22907, n22908, n22909,
    n22910, n22911, n22912, n22913, n22914, n22915,
    n22916, n22917, n22918, n22919, n22920, n22921,
    n22922, n22923, n22924, n22925, n22926, n22927,
    n22928, n22929, n22930, n22931, n22932, n22933,
    n22934, n22935, n22936, n22937, n22938, n22939,
    n22940, n22941, n22942, n22943, n22944, n22945,
    n22946, n22947, n22948, n22949, n22950, n22951,
    n22952, n22953, n22954, n22955, n22956, n22957,
    n22958, n22959, n22961, n22962, n22963, n22964,
    n22965, n22966, n22967, n22968, n22969, n22970,
    n22971, n22972, n22973, n22974, n22975, n22976,
    n22977, n22978, n22979, n22980, n22981, n22982,
    n22983, n22984, n22985, n22986, n22987, n22988,
    n22989, n22990, n22991, n22992, n22993, n22994,
    n22995, n22996, n22997, n22998, n22999, n23000,
    n23001, n23002, n23003, n23004, n23005, n23006,
    n23007, n23008, n23009, n23010, n23011, n23012,
    n23013, n23014, n23015, n23016, n23017, n23018,
    n23019, n23020, n23021, n23022, n23023, n23024,
    n23025, n23026, n23027, n23028, n23029, n23030,
    n23031, n23032, n23033, n23034, n23035, n23036,
    n23037, n23038, n23039, n23040, n23041, n23042,
    n23043, n23044, n23045, n23046, n23047, n23048,
    n23049, n23050, n23051, n23052, n23053, n23054,
    n23055, n23056, n23057, n23058, n23059, n23060,
    n23061, n23062, n23063, n23064, n23065, n23066,
    n23067, n23068, n23069, n23070, n23071, n23072,
    n23073, n23074, n23075, n23076, n23077, n23078,
    n23079, n23080, n23081, n23082, n23083, n23084,
    n23085, n23086, n23087, n23088, n23089, n23090,
    n23091, n23092, n23093, n23094, n23095, n23096,
    n23097, n23098, n23099, n23100, n23101, n23102,
    n23103, n23104, n23105, n23106, n23107, n23108,
    n23109, n23110, n23111, n23112, n23113, n23114,
    n23115, n23116, n23117, n23118, n23119, n23120,
    n23121, n23122, n23123, n23124, n23125, n23126,
    n23127, n23128, n23129, n23130, n23131, n23132,
    n23133, n23134, n23135, n23136, n23137, n23138,
    n23139, n23140, n23141, n23142, n23143, n23144,
    n23145, n23146, n23147, n23148, n23149, n23150,
    n23151, n23152, n23153, n23154, n23155, n23156,
    n23157, n23158, n23159, n23160, n23161, n23162,
    n23163, n23164, n23165, n23166, n23167, n23168,
    n23169, n23170, n23171, n23172, n23173, n23174,
    n23175, n23176, n23177, n23178, n23179, n23180,
    n23181, n23182, n23183, n23184, n23185, n23186,
    n23187, n23188, n23189, n23190, n23191, n23192,
    n23193, n23194, n23195, n23196, n23197, n23198,
    n23199, n23200, n23201, n23202, n23203, n23204,
    n23205, n23206, n23207, n23208, n23209, n23210,
    n23211, n23212, n23213, n23214, n23215, n23216,
    n23217, n23218, n23219, n23220, n23221, n23222,
    n23223, n23224, n23225, n23226, n23227, n23228,
    n23229, n23230, n23231, n23232, n23233, n23234,
    n23235, n23236, n23237, n23238, n23239, n23240,
    n23241, n23242, n23243, n23244, n23245, n23246,
    n23247, n23248, n23249, n23250, n23251, n23252,
    n23253, n23254, n23255, n23256, n23257, n23258,
    n23259, n23260, n23261, n23262, n23263, n23264,
    n23265, n23266, n23267, n23268, n23269, n23270,
    n23271, n23272, n23273, n23274, n23275, n23276,
    n23277, n23278, n23279, n23280, n23281, n23282,
    n23283, n23284, n23285, n23286, n23287, n23288,
    n23289, n23290, n23291, n23292, n23293, n23294,
    n23295, n23296, n23297, n23298, n23299, n23300,
    n23301, n23302, n23303, n23304, n23305, n23306,
    n23307, n23308, n23309, n23310, n23311, n23312,
    n23313, n23314, n23315, n23316, n23317, n23318,
    n23319, n23320, n23321, n23322, n23323, n23324,
    n23325, n23326, n23327, n23328, n23329, n23330,
    n23331, n23332, n23333, n23334, n23335, n23336,
    n23337, n23338, n23339, n23340, n23341, n23342,
    n23343, n23344, n23345, n23346, n23347, n23348,
    n23349, n23350, n23351, n23352, n23353, n23354,
    n23355, n23356, n23357, n23358, n23359, n23360,
    n23361, n23362, n23363, n23364, n23365, n23366,
    n23367, n23368, n23369, n23370, n23371, n23372,
    n23373, n23374, n23375, n23376, n23377, n23378,
    n23379, n23380, n23381, n23382, n23383, n23384,
    n23385, n23386, n23387, n23388, n23389, n23390,
    n23391, n23392, n23393, n23395, n23396, n23397,
    n23398, n23399, n23400, n23401, n23402, n23403,
    n23404, n23405, n23406, n23407, n23408, n23409,
    n23410, n23411, n23412, n23413, n23414, n23415,
    n23416, n23417, n23418, n23419, n23420, n23421,
    n23422, n23423, n23424, n23425, n23426, n23427,
    n23428, n23429, n23430, n23431, n23432, n23433,
    n23434, n23435, n23436, n23437, n23438, n23439,
    n23440, n23441, n23442, n23443, n23444, n23445,
    n23446, n23447, n23448, n23449, n23450, n23451,
    n23452, n23453, n23454, n23455, n23456, n23457,
    n23458, n23459, n23460, n23461, n23462, n23463,
    n23464, n23465, n23466, n23467, n23468, n23469,
    n23470, n23471, n23472, n23473, n23474, n23475,
    n23476, n23477, n23478, n23479, n23480, n23481,
    n23482, n23483, n23484, n23485, n23486, n23487,
    n23488, n23489, n23490, n23491, n23492, n23493,
    n23494, n23495, n23496, n23497, n23498, n23499,
    n23500, n23501, n23502, n23503, n23504, n23505,
    n23506, n23507, n23508, n23509, n23510, n23511,
    n23512, n23513, n23514, n23515, n23516, n23517,
    n23518, n23519, n23520, n23521, n23522, n23523,
    n23524, n23525, n23526, n23527, n23528, n23529,
    n23530, n23531, n23532, n23533, n23534, n23535,
    n23536, n23537, n23538, n23539, n23540, n23541,
    n23542, n23543, n23544, n23545, n23546, n23547,
    n23548, n23549, n23550, n23551, n23552, n23553,
    n23554, n23555, n23556, n23557, n23558, n23559,
    n23560, n23561, n23562, n23563, n23564, n23565,
    n23566, n23567, n23568, n23569, n23570, n23571,
    n23572, n23573, n23574, n23575, n23576, n23577,
    n23578, n23579, n23580, n23581, n23582, n23583,
    n23584, n23585, n23586, n23587, n23588, n23589,
    n23590, n23591, n23592, n23593, n23594, n23595,
    n23596, n23597, n23598, n23599, n23600, n23601,
    n23602, n23603, n23604, n23605, n23606, n23607,
    n23608, n23609, n23610, n23611, n23612, n23613,
    n23614, n23615, n23616, n23617, n23618, n23619,
    n23620, n23621, n23622, n23623, n23624, n23625,
    n23626, n23627, n23628, n23629, n23630, n23631,
    n23632, n23633, n23634, n23635, n23636, n23637,
    n23638, n23639, n23640, n23641, n23642, n23643,
    n23644, n23645, n23646, n23647, n23648, n23649,
    n23650, n23651, n23652, n23653, n23654, n23655,
    n23656, n23657, n23658, n23659, n23660, n23661,
    n23662, n23663, n23664, n23665, n23666, n23667,
    n23668, n23669, n23670, n23671, n23672, n23673,
    n23674, n23675, n23676, n23677, n23678, n23679,
    n23680, n23681, n23682, n23683, n23684, n23685,
    n23686, n23687, n23688, n23689, n23690, n23691,
    n23692, n23693, n23694, n23695, n23696, n23697,
    n23698, n23699, n23700, n23701, n23702, n23703,
    n23704, n23705, n23706, n23707, n23708, n23709,
    n23710, n23711, n23712, n23713, n23714, n23715,
    n23716, n23717, n23718, n23719, n23720, n23721,
    n23722, n23723, n23724, n23725, n23726, n23727,
    n23728, n23729, n23730, n23731, n23732, n23733,
    n23734, n23735, n23736, n23737, n23738, n23739,
    n23740, n23741, n23742, n23743, n23744, n23745,
    n23746, n23747, n23748, n23749, n23750, n23751,
    n23752, n23753, n23754, n23755, n23756, n23757,
    n23758, n23759, n23760, n23761, n23762, n23763,
    n23764, n23765, n23766, n23767, n23768, n23769,
    n23770, n23771, n23772, n23773, n23774, n23775,
    n23776, n23777, n23778, n23779, n23780, n23781,
    n23782, n23783, n23784, n23785, n23786, n23787,
    n23788, n23789, n23790, n23791, n23792, n23793,
    n23794, n23795, n23796, n23797, n23798, n23799,
    n23800, n23801, n23802, n23803, n23804, n23805,
    n23806, n23807, n23808, n23809, n23810, n23811,
    n23812, n23813, n23814, n23815, n23816, n23817,
    n23818, n23819, n23820, n23821, n23822, n23823,
    n23824, n23825, n23826, n23827, n23828, n23829,
    n23830, n23831, n23832, n23833, n23834, n23835,
    n23836, n23837, n23838, n23839, n23840, n23841,
    n23842, n23843, n23844, n23845, n23846, n23847,
    n23848, n23850, n23851, n23852, n23853, n23854,
    n23855, n23856, n23857, n23858, n23859, n23860,
    n23861, n23862, n23863, n23864, n23865, n23866,
    n23867, n23868, n23869, n23870, n23871, n23872,
    n23873, n23874, n23875, n23876, n23877, n23878,
    n23879, n23880, n23881, n23882, n23883, n23884,
    n23885, n23886, n23887, n23888, n23889, n23890,
    n23891, n23892, n23893, n23894, n23895, n23896,
    n23897, n23898, n23899, n23900, n23901, n23902,
    n23903, n23904, n23905, n23906, n23907, n23908,
    n23909, n23910, n23911, n23912, n23913, n23914,
    n23915, n23916, n23917, n23918, n23919, n23920,
    n23921, n23922, n23923, n23924, n23925, n23926,
    n23927, n23928, n23929, n23930, n23931, n23932,
    n23933, n23934, n23935, n23936, n23937, n23938,
    n23939, n23940, n23941, n23942, n23943, n23944,
    n23945, n23946, n23947, n23948, n23949, n23950,
    n23951, n23952, n23953, n23954, n23955, n23956,
    n23957, n23958, n23959, n23960, n23961, n23962,
    n23963, n23964, n23965, n23966, n23967, n23968,
    n23969, n23970, n23971, n23972, n23973, n23974,
    n23975, n23976, n23977, n23978, n23979, n23980,
    n23981, n23982, n23983, n23984, n23985, n23986,
    n23987, n23988, n23989, n23990, n23991, n23992,
    n23993, n23994, n23995, n23996, n23997, n23998,
    n23999, n24000, n24001, n24002, n24003, n24004,
    n24005, n24006, n24007, n24008, n24009, n24010,
    n24011, n24012, n24013, n24014, n24015, n24016,
    n24017, n24018, n24019, n24020, n24021, n24022,
    n24023, n24024, n24025, n24026, n24027, n24028,
    n24029, n24030, n24031, n24032, n24033, n24034,
    n24035, n24036, n24037, n24038, n24039, n24040,
    n24041, n24042, n24043, n24044, n24045, n24046,
    n24047, n24048, n24049, n24050, n24051, n24052,
    n24053, n24054, n24055, n24056, n24057, n24058,
    n24059, n24060, n24061, n24062, n24063, n24064,
    n24065, n24066, n24067, n24068, n24069, n24070,
    n24071, n24072, n24073, n24074, n24075, n24076,
    n24077, n24078, n24079, n24080, n24081, n24082,
    n24083, n24084, n24085, n24086, n24087, n24088,
    n24089, n24090, n24091, n24092, n24093, n24094,
    n24095, n24096, n24097, n24098, n24099, n24100,
    n24101, n24102, n24103, n24104, n24105, n24106,
    n24107, n24108, n24109, n24110, n24111, n24112,
    n24113, n24114, n24115, n24116, n24117, n24118,
    n24119, n24120, n24121, n24122, n24123, n24124,
    n24125, n24126, n24127, n24128, n24129, n24130,
    n24131, n24132, n24133, n24134, n24135, n24136,
    n24137, n24138, n24139, n24140, n24141, n24142,
    n24143, n24144, n24145, n24146, n24147, n24148,
    n24149, n24150, n24151, n24152, n24153, n24154,
    n24155, n24156, n24157, n24158, n24159, n24160,
    n24161, n24162, n24163, n24164, n24165, n24166,
    n24167, n24168, n24169, n24170, n24171, n24172,
    n24173, n24174, n24175, n24176, n24177, n24178,
    n24179, n24180, n24181, n24182, n24183, n24184,
    n24185, n24186, n24187, n24188, n24189, n24190,
    n24191, n24192, n24193, n24194, n24195, n24196,
    n24197, n24198, n24199, n24200, n24201, n24202,
    n24203, n24204, n24205, n24206, n24207, n24208,
    n24209, n24210, n24211, n24212, n24213, n24214,
    n24215, n24216, n24217, n24218, n24219, n24220,
    n24221, n24222, n24223, n24224, n24225, n24226,
    n24227, n24228, n24229, n24230, n24231, n24232,
    n24233, n24234, n24235, n24236, n24237, n24238,
    n24239, n24240, n24241, n24242, n24243, n24244,
    n24245, n24246, n24247, n24248, n24249, n24250,
    n24251, n24252, n24253, n24254, n24255, n24256,
    n24257, n24258, n24259, n24260, n24261, n24262,
    n24263, n24264, n24265, n24266, n24267, n24268,
    n24269, n24270, n24271, n24272, n24273, n24274,
    n24275, n24276, n24277, n24278, n24279, n24280,
    n24281, n24282, n24283, n24284, n24285, n24286,
    n24287, n24288, n24289, n24290, n24291, n24292,
    n24293, n24294, n24295, n24296, n24297, n24298,
    n24299, n24300, n24301, n24303, n24304, n24305,
    n24306, n24307, n24308, n24309, n24310, n24311,
    n24312, n24313, n24314, n24315, n24316, n24317,
    n24318, n24319, n24320, n24321, n24322, n24323,
    n24324, n24325, n24326, n24327, n24328, n24329,
    n24330, n24331, n24332, n24333, n24334, n24335,
    n24336, n24337, n24338, n24339, n24340, n24341,
    n24342, n24343, n24344, n24345, n24346, n24347,
    n24348, n24349, n24350, n24351, n24352, n24353,
    n24354, n24355, n24356, n24357, n24358, n24359,
    n24360, n24361, n24362, n24363, n24364, n24365,
    n24366, n24367, n24368, n24369, n24370, n24371,
    n24372, n24373, n24374, n24375, n24376, n24377,
    n24378, n24379, n24380, n24381, n24382, n24383,
    n24384, n24385, n24386, n24387, n24388, n24389,
    n24390, n24391, n24392, n24393, n24394, n24395,
    n24396, n24397, n24398, n24399, n24400, n24401,
    n24402, n24403, n24404, n24405, n24406, n24407,
    n24408, n24409, n24410, n24411, n24412, n24413,
    n24414, n24415, n24416, n24417, n24418, n24419,
    n24420, n24421, n24422, n24423, n24424, n24425,
    n24426, n24427, n24428, n24429, n24430, n24431,
    n24432, n24433, n24434, n24435, n24436, n24437,
    n24438, n24439, n24440, n24441, n24442, n24443,
    n24444, n24445, n24446, n24447, n24448, n24449,
    n24450, n24451, n24452, n24453, n24454, n24455,
    n24456, n24457, n24458, n24459, n24460, n24461,
    n24462, n24463, n24464, n24465, n24466, n24467,
    n24468, n24469, n24470, n24471, n24472, n24473,
    n24474, n24475, n24476, n24477, n24478, n24479,
    n24480, n24481, n24482, n24483, n24484, n24485,
    n24486, n24487, n24488, n24489, n24490, n24491,
    n24492, n24493, n24494, n24495, n24496, n24497,
    n24498, n24499, n24500, n24501, n24502, n24503,
    n24504, n24505, n24506, n24507, n24508, n24509,
    n24510, n24511, n24512, n24513, n24514, n24515,
    n24516, n24517, n24518, n24519, n24520, n24521,
    n24522, n24523, n24524, n24525, n24526, n24527,
    n24528, n24529, n24530, n24531, n24532, n24533,
    n24534, n24535, n24536, n24537, n24538, n24539,
    n24540, n24541, n24542, n24543, n24544, n24545,
    n24546, n24547, n24548, n24549, n24550, n24551,
    n24552, n24553, n24554, n24555, n24556, n24557,
    n24558, n24559, n24560, n24561, n24562, n24563,
    n24564, n24565, n24566, n24567, n24568, n24569,
    n24570, n24571, n24572, n24573, n24574, n24575,
    n24576, n24577, n24578, n24579, n24580, n24581,
    n24582, n24583, n24584, n24585, n24586, n24587,
    n24588, n24589, n24590, n24591, n24592, n24593,
    n24594, n24595, n24596, n24597, n24598, n24599,
    n24600, n24601, n24602, n24603, n24604, n24605,
    n24606, n24607, n24608, n24609, n24610, n24611,
    n24612, n24613, n24614, n24615, n24616, n24617,
    n24618, n24619, n24620, n24621, n24622, n24623,
    n24624, n24625, n24626, n24627, n24628, n24629,
    n24630, n24631, n24632, n24633, n24634, n24635,
    n24636, n24637, n24638, n24639, n24640, n24641,
    n24642, n24643, n24644, n24645, n24646, n24647,
    n24648, n24649, n24650, n24651, n24652, n24653,
    n24654, n24655, n24656, n24657, n24658, n24659,
    n24660, n24661, n24662, n24663, n24664, n24665,
    n24666, n24667, n24668, n24669, n24670, n24671,
    n24672, n24673, n24674, n24675, n24676, n24677,
    n24678, n24679, n24680, n24681, n24682, n24683,
    n24684, n24685, n24686, n24687, n24688, n24689,
    n24690, n24691, n24692, n24693, n24694, n24695,
    n24696, n24697, n24698, n24699, n24700, n24701,
    n24702, n24703, n24704, n24705, n24706, n24707,
    n24708, n24709, n24710, n24711, n24712, n24713,
    n24714, n24715, n24716, n24717, n24718, n24719,
    n24720, n24721, n24722, n24723, n24724, n24725,
    n24726, n24727, n24728, n24729, n24730, n24731,
    n24732, n24733, n24734, n24735, n24736, n24737,
    n24738, n24739, n24740, n24741, n24742, n24743,
    n24744, n24745, n24746, n24747, n24748, n24749,
    n24750, n24751, n24753, n24754, n24755, n24756,
    n24757, n24758, n24759, n24760, n24761, n24762,
    n24763, n24764, n24765, n24766, n24767, n24768,
    n24769, n24770, n24771, n24772, n24773, n24774,
    n24775, n24776, n24777, n24778, n24779, n24780,
    n24781, n24782, n24783, n24784, n24785, n24786,
    n24787, n24788, n24789, n24790, n24791, n24792,
    n24793, n24794, n24795, n24796, n24797, n24798,
    n24799, n24800, n24801, n24802, n24803, n24804,
    n24805, n24806, n24807, n24808, n24809, n24810,
    n24811, n24812, n24813, n24814, n24815, n24816,
    n24817, n24818, n24819, n24820, n24821, n24822,
    n24823, n24824, n24825, n24826, n24827, n24828,
    n24829, n24830, n24831, n24832, n24833, n24834,
    n24835, n24836, n24837, n24838, n24839, n24840,
    n24841, n24842, n24843, n24844, n24845, n24846,
    n24847, n24848, n24849, n24850, n24851, n24852,
    n24853, n24854, n24855, n24856, n24857, n24858,
    n24859, n24860, n24861, n24862, n24863, n24864,
    n24865, n24866, n24867, n24868, n24869, n24870,
    n24871, n24872, n24873, n24874, n24875, n24876,
    n24877, n24878, n24879, n24880, n24881, n24882,
    n24883, n24884, n24885, n24886, n24887, n24888,
    n24889, n24890, n24891, n24892, n24893, n24894,
    n24895, n24896, n24897, n24898, n24899, n24900,
    n24901, n24902, n24903, n24904, n24905, n24906,
    n24907, n24908, n24909, n24910, n24911, n24912,
    n24913, n24914, n24915, n24916, n24917, n24918,
    n24919, n24920, n24921, n24922, n24923, n24924,
    n24925, n24926, n24927, n24928, n24929, n24930,
    n24931, n24932, n24933, n24934, n24935, n24936,
    n24937, n24938, n24939, n24940, n24941, n24942,
    n24943, n24944, n24945, n24946, n24947, n24948,
    n24949, n24950, n24951, n24952, n24953, n24954,
    n24955, n24956, n24957, n24958, n24959, n24960,
    n24961, n24962, n24963, n24964, n24965, n24966,
    n24967, n24968, n24969, n24970, n24971, n24972,
    n24973, n24974, n24975, n24976, n24977, n24978,
    n24979, n24980, n24981, n24982, n24983, n24984,
    n24985, n24986, n24987, n24988, n24989, n24990,
    n24991, n24992, n24993, n24994, n24995, n24996,
    n24997, n24998, n24999, n25000, n25001, n25002,
    n25003, n25004, n25005, n25006, n25007, n25008,
    n25009, n25010, n25011, n25012, n25013, n25014,
    n25015, n25016, n25017, n25018, n25019, n25020,
    n25021, n25022, n25023, n25024, n25025, n25026,
    n25027, n25028, n25029, n25030, n25031, n25032,
    n25033, n25034, n25035, n25036, n25037, n25038,
    n25039, n25040, n25041, n25042, n25043, n25044,
    n25045, n25046, n25047, n25048, n25049, n25050,
    n25051, n25052, n25053, n25054, n25055, n25056,
    n25057, n25058, n25059, n25060, n25061, n25062,
    n25063, n25064, n25065, n25066, n25067, n25068,
    n25069, n25070, n25071, n25072, n25073, n25074,
    n25075, n25076, n25077, n25078, n25079, n25080,
    n25081, n25082, n25083, n25084, n25085, n25086,
    n25087, n25088, n25089, n25090, n25091, n25092,
    n25093, n25094, n25095, n25096, n25097, n25098,
    n25099, n25100, n25101, n25102, n25103, n25104,
    n25105, n25106, n25107, n25108, n25109, n25110,
    n25111, n25112, n25113, n25114, n25115, n25116,
    n25117, n25118, n25119, n25120, n25121, n25122,
    n25123, n25124, n25125, n25126, n25127, n25128,
    n25129, n25130, n25131, n25132, n25133, n25134,
    n25135, n25136, n25137, n25138, n25139, n25140,
    n25141, n25142, n25143, n25144, n25145, n25146,
    n25147, n25148, n25149, n25150, n25151, n25152,
    n25153, n25154, n25155, n25156, n25157, n25158,
    n25159, n25160, n25161, n25162, n25163, n25164,
    n25165, n25166, n25167, n25168, n25169, n25170,
    n25171, n25172, n25173, n25174, n25175, n25176,
    n25177, n25178, n25179, n25180, n25181, n25182,
    n25183, n25184, n25185, n25186, n25187, n25188,
    n25189, n25190, n25191, n25192, n25193, n25194,
    n25195, n25196, n25197, n25198, n25199, n25200,
    n25201, n25202, n25204, n25205, n25206, n25207,
    n25208, n25209, n25210, n25211, n25212, n25213,
    n25214, n25215, n25216, n25217, n25218, n25219,
    n25220, n25221, n25222, n25223, n25224, n25225,
    n25226, n25227, n25228, n25229, n25230, n25231,
    n25232, n25233, n25234, n25235, n25236, n25237,
    n25238, n25239, n25240, n25241, n25242, n25243,
    n25244, n25245, n25246, n25247, n25248, n25249,
    n25250, n25251, n25252, n25253, n25254, n25255,
    n25256, n25257, n25258, n25259, n25260, n25261,
    n25262, n25263, n25264, n25265, n25266, n25267,
    n25268, n25269, n25270, n25271, n25272, n25273,
    n25274, n25275, n25276, n25277, n25278, n25279,
    n25280, n25281, n25282, n25283, n25284, n25285,
    n25286, n25287, n25288, n25289, n25290, n25291,
    n25292, n25293, n25294, n25295, n25296, n25297,
    n25298, n25299, n25300, n25301, n25302, n25303,
    n25304, n25305, n25306, n25307, n25308, n25309,
    n25310, n25311, n25312, n25313, n25314, n25315,
    n25316, n25317, n25318, n25319, n25320, n25321,
    n25322, n25323, n25324, n25325, n25326, n25327,
    n25328, n25329, n25330, n25331, n25332, n25333,
    n25334, n25335, n25336, n25337, n25338, n25339,
    n25340, n25341, n25342, n25343, n25344, n25345,
    n25346, n25347, n25348, n25349, n25350, n25351,
    n25352, n25353, n25354, n25355, n25356, n25357,
    n25358, n25359, n25360, n25361, n25362, n25363,
    n25364, n25365, n25366, n25367, n25368, n25369,
    n25370, n25371, n25372, n25373, n25374, n25375,
    n25376, n25377, n25378, n25379, n25380, n25381,
    n25382, n25383, n25384, n25385, n25386, n25387,
    n25388, n25389, n25390, n25391, n25392, n25393,
    n25394, n25395, n25396, n25397, n25398, n25399,
    n25400, n25401, n25402, n25403, n25404, n25405,
    n25406, n25407, n25408, n25409, n25410, n25411,
    n25412, n25413, n25414, n25415, n25416, n25417,
    n25418, n25419, n25420, n25421, n25422, n25423,
    n25424, n25425, n25426, n25427, n25428, n25429,
    n25430, n25431, n25432, n25433, n25434, n25435,
    n25436, n25437, n25438, n25439, n25440, n25441,
    n25442, n25443, n25444, n25445, n25446, n25447,
    n25448, n25449, n25450, n25451, n25452, n25453,
    n25454, n25455, n25456, n25457, n25458, n25459,
    n25460, n25461, n25462, n25463, n25464, n25465,
    n25466, n25467, n25468, n25469, n25470, n25471,
    n25472, n25473, n25474, n25475, n25476, n25477,
    n25478, n25479, n25480, n25481, n25482, n25483,
    n25484, n25485, n25486, n25487, n25488, n25489,
    n25490, n25491, n25492, n25493, n25494, n25495,
    n25496, n25497, n25498, n25499, n25500, n25501,
    n25502, n25503, n25504, n25505, n25506, n25507,
    n25508, n25509, n25510, n25511, n25512, n25513,
    n25514, n25515, n25516, n25517, n25518, n25519,
    n25520, n25521, n25522, n25523, n25524, n25525,
    n25526, n25527, n25528, n25529, n25530, n25531,
    n25532, n25533, n25534, n25535, n25536, n25537,
    n25538, n25539, n25540, n25541, n25542, n25543,
    n25544, n25545, n25546, n25547, n25548, n25549,
    n25550, n25551, n25552, n25553, n25554, n25555,
    n25556, n25557, n25558, n25559, n25560, n25561,
    n25562, n25563, n25564, n25565, n25566, n25567,
    n25568, n25569, n25570, n25571, n25572, n25573,
    n25574, n25575, n25576, n25577, n25578, n25579,
    n25580, n25581, n25582, n25583, n25584, n25585,
    n25586, n25587, n25588, n25589, n25590, n25591,
    n25592, n25593, n25594, n25595, n25596, n25597,
    n25598, n25599, n25600, n25601, n25602, n25603,
    n25604, n25605, n25606, n25607, n25608, n25609,
    n25610, n25611, n25612, n25613, n25614, n25615,
    n25616, n25617, n25618, n25619, n25620, n25621,
    n25622, n25623, n25624, n25625, n25626, n25627,
    n25628, n25629, n25630, n25631, n25632, n25633,
    n25634, n25635, n25636, n25637, n25638, n25639,
    n25640, n25641, n25642, n25643, n25644, n25645,
    n25646, n25647, n25648, n25649, n25650, n25651,
    n25652, n25653, n25655, n25656, n25657, n25658,
    n25659, n25660, n25661, n25662, n25663, n25664,
    n25665, n25666, n25667, n25668, n25669, n25670,
    n25671, n25672, n25673, n25674, n25675, n25676,
    n25677, n25678, n25679, n25680, n25681, n25682,
    n25683, n25684, n25685, n25686, n25687, n25688,
    n25689, n25690, n25691, n25692, n25693, n25694,
    n25695, n25696, n25697, n25698, n25699, n25700,
    n25701, n25702, n25703, n25704, n25705, n25706,
    n25707, n25708, n25709, n25710, n25711, n25712,
    n25713, n25714, n25715, n25716, n25717, n25718,
    n25719, n25720, n25721, n25722, n25723, n25724,
    n25725, n25726, n25727, n25728, n25729, n25730,
    n25731, n25732, n25733, n25734, n25735, n25736,
    n25737, n25738, n25739, n25740, n25741, n25742,
    n25743, n25744, n25745, n25746, n25747, n25748,
    n25749, n25750, n25751, n25752, n25753, n25754,
    n25755, n25756, n25757, n25758, n25759, n25760,
    n25761, n25762, n25763, n25764, n25765, n25766,
    n25767, n25768, n25769, n25770, n25771, n25772,
    n25773, n25774, n25775, n25776, n25777, n25778,
    n25779, n25780, n25781, n25782, n25783, n25784,
    n25785, n25786, n25787, n25788, n25789, n25790,
    n25791, n25792, n25793, n25794, n25795, n25796,
    n25797, n25798, n25799, n25800, n25801, n25802,
    n25803, n25804, n25805, n25806, n25807, n25808,
    n25809, n25810, n25811, n25812, n25813, n25814,
    n25815, n25816, n25817, n25818, n25819, n25820,
    n25821, n25822, n25823, n25824, n25825, n25826,
    n25827, n25828, n25829, n25830, n25831, n25832,
    n25833, n25834, n25835, n25836, n25837, n25838,
    n25839, n25840, n25841, n25842, n25843, n25844,
    n25845, n25846, n25847, n25848, n25849, n25850,
    n25851, n25852, n25853, n25854, n25855, n25856,
    n25857, n25858, n25859, n25860, n25861, n25862,
    n25863, n25864, n25865, n25866, n25867, n25868,
    n25869, n25870, n25871, n25872, n25873, n25874,
    n25875, n25876, n25877, n25878, n25879, n25880,
    n25881, n25882, n25883, n25884, n25885, n25886,
    n25887, n25888, n25889, n25890, n25891, n25892,
    n25893, n25894, n25895, n25896, n25897, n25898,
    n25899, n25900, n25901, n25902, n25903, n25904,
    n25905, n25906, n25907, n25908, n25909, n25910,
    n25911, n25912, n25913, n25914, n25915, n25916,
    n25917, n25918, n25919, n25920, n25921, n25922,
    n25923, n25924, n25925, n25926, n25927, n25928,
    n25929, n25930, n25931, n25932, n25933, n25934,
    n25935, n25936, n25937, n25938, n25939, n25940,
    n25941, n25942, n25943, n25944, n25945, n25946,
    n25947, n25948, n25949, n25950, n25951, n25952,
    n25953, n25954, n25955, n25956, n25957, n25958,
    n25959, n25960, n25961, n25962, n25963, n25964,
    n25965, n25966, n25967, n25968, n25969, n25970,
    n25971, n25972, n25973, n25974, n25975, n25976,
    n25977, n25978, n25979, n25980, n25981, n25982,
    n25983, n25984, n25985, n25986, n25987, n25988,
    n25989, n25990, n25991, n25992, n25993, n25994,
    n25995, n25996, n25997, n25998, n25999, n26000,
    n26001, n26002, n26003, n26004, n26005, n26006,
    n26007, n26008, n26009, n26010, n26011, n26012,
    n26013, n26014, n26015, n26016, n26017, n26018,
    n26019, n26020, n26021, n26022, n26023, n26024,
    n26025, n26026, n26027, n26028, n26029, n26030,
    n26031, n26032, n26033, n26034, n26035, n26036,
    n26037, n26038, n26039, n26040, n26041, n26042,
    n26043, n26044, n26045, n26046, n26047, n26048,
    n26049, n26050, n26051, n26052, n26053, n26054,
    n26055, n26056, n26057, n26058, n26059, n26060,
    n26061, n26062, n26063, n26064, n26065, n26066,
    n26067, n26068, n26069, n26070, n26071, n26072,
    n26073, n26074, n26075, n26076, n26077, n26078,
    n26079, n26080, n26081, n26082, n26083, n26084,
    n26085, n26086, n26087, n26088, n26089, n26090,
    n26091, n26092, n26093, n26094, n26095, n26096,
    n26097, n26098, n26099, n26100, n26101, n26102,
    n26103, n26104, n26105, n26106, n26108, n26109,
    n26110, n26111, n26112, n26113, n26114, n26115,
    n26116, n26117, n26118, n26119, n26120, n26121,
    n26122, n26123, n26124, n26125, n26126, n26127,
    n26128, n26129, n26130, n26131, n26132, n26133,
    n26134, n26135, n26136, n26137, n26138, n26139,
    n26140, n26141, n26142, n26143, n26144, n26145,
    n26146, n26147, n26148, n26149, n26150, n26151,
    n26152, n26153, n26154, n26155, n26156, n26157,
    n26158, n26159, n26160, n26161, n26162, n26163,
    n26164, n26165, n26166, n26167, n26168, n26169,
    n26170, n26171, n26172, n26173, n26174, n26175,
    n26176, n26177, n26178, n26179, n26180, n26181,
    n26182, n26183, n26184, n26185, n26186, n26187,
    n26188, n26189, n26190, n26191, n26192, n26193,
    n26194, n26195, n26196, n26197, n26198, n26199,
    n26200, n26201, n26202, n26203, n26204, n26205,
    n26206, n26207, n26208, n26209, n26210, n26211,
    n26212, n26213, n26214, n26215, n26216, n26217,
    n26218, n26219, n26220, n26221, n26222, n26223,
    n26224, n26225, n26226, n26227, n26228, n26229,
    n26230, n26231, n26232, n26233, n26234, n26235,
    n26236, n26237, n26238, n26239, n26240, n26241,
    n26242, n26243, n26244, n26245, n26246, n26247,
    n26248, n26249, n26250, n26251, n26252, n26253,
    n26254, n26255, n26256, n26257, n26258, n26259,
    n26260, n26261, n26262, n26263, n26264, n26265,
    n26266, n26267, n26268, n26269, n26270, n26271,
    n26272, n26273, n26274, n26275, n26276, n26277,
    n26278, n26279, n26280, n26281, n26282, n26283,
    n26284, n26285, n26286, n26287, n26288, n26289,
    n26290, n26291, n26292, n26293, n26294, n26295,
    n26296, n26297, n26298, n26299, n26300, n26301,
    n26302, n26303, n26304, n26305, n26306, n26307,
    n26308, n26309, n26310, n26311, n26312, n26313,
    n26314, n26315, n26316, n26317, n26318, n26319,
    n26320, n26321, n26322, n26323, n26324, n26325,
    n26326, n26327, n26328, n26329, n26330, n26331,
    n26332, n26333, n26334, n26335, n26336, n26337,
    n26338, n26339, n26340, n26341, n26342, n26343,
    n26344, n26345, n26346, n26347, n26348, n26349,
    n26350, n26351, n26352, n26353, n26354, n26355,
    n26356, n26357, n26358, n26359, n26360, n26361,
    n26362, n26363, n26364, n26365, n26366, n26367,
    n26368, n26369, n26370, n26371, n26372, n26373,
    n26374, n26375, n26376, n26377, n26378, n26379,
    n26380, n26381, n26382, n26383, n26384, n26385,
    n26386, n26387, n26388, n26389, n26390, n26391,
    n26392, n26393, n26394, n26395, n26396, n26397,
    n26398, n26399, n26400, n26401, n26402, n26403,
    n26404, n26405, n26406, n26407, n26408, n26409,
    n26410, n26411, n26412, n26413, n26414, n26415,
    n26416, n26417, n26418, n26419, n26420, n26421,
    n26422, n26423, n26424, n26425, n26426, n26427,
    n26428, n26429, n26430, n26431, n26432, n26433,
    n26434, n26435, n26436, n26437, n26438, n26439,
    n26440, n26441, n26442, n26443, n26444, n26445,
    n26446, n26447, n26448, n26449, n26450, n26451,
    n26452, n26453, n26454, n26455, n26456, n26457,
    n26458, n26459, n26460, n26461, n26462, n26463,
    n26464, n26465, n26466, n26467, n26468, n26469,
    n26470, n26471, n26472, n26473, n26474, n26475,
    n26476, n26477, n26478, n26479, n26480, n26481,
    n26482, n26483, n26484, n26485, n26486, n26487,
    n26488, n26489, n26490, n26491, n26492, n26493,
    n26494, n26495, n26496, n26497, n26498, n26499,
    n26500, n26501, n26502, n26503, n26504, n26505,
    n26506, n26507, n26508, n26509, n26510, n26511,
    n26512, n26513, n26514, n26515, n26516, n26517,
    n26518, n26519, n26520, n26521, n26522, n26523,
    n26524, n26525, n26526, n26527, n26528, n26529,
    n26530, n26531, n26532, n26533, n26534, n26535,
    n26536, n26537, n26538, n26539, n26540, n26541,
    n26542, n26543, n26544, n26545, n26546, n26547,
    n26548, n26549, n26550, n26551, n26552, n26553,
    n26554, n26555, n26556, n26557, n26558, n26559,
    n26561, n26562, n26563, n26564, n26565, n26566,
    n26567, n26568, n26569, n26570, n26571, n26572,
    n26573, n26574, n26575, n26576, n26577, n26578,
    n26579, n26580, n26581, n26582, n26583, n26584,
    n26585, n26586, n26587, n26588, n26589, n26590,
    n26591, n26592, n26593, n26594, n26595, n26596,
    n26597, n26598, n26599, n26600, n26601, n26602,
    n26603, n26604, n26605, n26606, n26607, n26608,
    n26609, n26610, n26611, n26612, n26613, n26614,
    n26615, n26616, n26617, n26618, n26619, n26620,
    n26621, n26622, n26623, n26624, n26625, n26626,
    n26627, n26628, n26629, n26630, n26631, n26632,
    n26633, n26634, n26635, n26636, n26637, n26638,
    n26639, n26640, n26641, n26642, n26643, n26644,
    n26645, n26646, n26647, n26648, n26649, n26650,
    n26651, n26652, n26653, n26654, n26655, n26656,
    n26657, n26658, n26659, n26660, n26661, n26662,
    n26663, n26664, n26665, n26666, n26667, n26668,
    n26669, n26670, n26671, n26672, n26673, n26674,
    n26675, n26676, n26677, n26678, n26679, n26680,
    n26681, n26682, n26683, n26684, n26685, n26686,
    n26687, n26688, n26689, n26690, n26691, n26692,
    n26693, n26694, n26695, n26696, n26697, n26698,
    n26699, n26700, n26701, n26702, n26703, n26704,
    n26705, n26706, n26707, n26708, n26709, n26710,
    n26711, n26712, n26713, n26714, n26715, n26716,
    n26717, n26718, n26719, n26720, n26721, n26722,
    n26723, n26724, n26725, n26726, n26727, n26728,
    n26729, n26730, n26731, n26732, n26733, n26734,
    n26735, n26736, n26737, n26738, n26739, n26740,
    n26741, n26742, n26743, n26744, n26745, n26746,
    n26747, n26748, n26749, n26750, n26751, n26752,
    n26753, n26754, n26755, n26756, n26757, n26758,
    n26759, n26760, n26761, n26762, n26763, n26764,
    n26765, n26766, n26767, n26768, n26769, n26770,
    n26771, n26772, n26773, n26774, n26775, n26776,
    n26777, n26778, n26779, n26780, n26781, n26782,
    n26783, n26784, n26785, n26786, n26787, n26788,
    n26789, n26790, n26791, n26792, n26793, n26794,
    n26795, n26796, n26797, n26798, n26799, n26800,
    n26801, n26802, n26803, n26804, n26805, n26806,
    n26807, n26808, n26809, n26810, n26811, n26812,
    n26813, n26814, n26815, n26816, n26817, n26818,
    n26819, n26820, n26821, n26822, n26823, n26824,
    n26825, n26826, n26827, n26828, n26829, n26830,
    n26831, n26832, n26833, n26834, n26835, n26836,
    n26837, n26838, n26839, n26840, n26841, n26842,
    n26843, n26844, n26845, n26846, n26847, n26848,
    n26849, n26850, n26851, n26852, n26853, n26854,
    n26855, n26856, n26857, n26858, n26859, n26860,
    n26861, n26862, n26863, n26864, n26865, n26866,
    n26867, n26868, n26869, n26870, n26871, n26872,
    n26873, n26874, n26875, n26876, n26877, n26878,
    n26879, n26880, n26881, n26882, n26883, n26884,
    n26885, n26886, n26887, n26888, n26889, n26890,
    n26891, n26892, n26893, n26894, n26895, n26896,
    n26897, n26898, n26899, n26900, n26901, n26902,
    n26903, n26904, n26905, n26906, n26907, n26908,
    n26909, n26910, n26911, n26912, n26913, n26914,
    n26915, n26916, n26917, n26918, n26919, n26920,
    n26921, n26922, n26923, n26924, n26925, n26926,
    n26927, n26928, n26929, n26930, n26931, n26932,
    n26933, n26934, n26935, n26936, n26937, n26938,
    n26939, n26940, n26941, n26942, n26943, n26944,
    n26945, n26946, n26947, n26948, n26949, n26950,
    n26951, n26952, n26953, n26954, n26955, n26956,
    n26957, n26958, n26959, n26960, n26961, n26962,
    n26963, n26964, n26965, n26966, n26967, n26968,
    n26969, n26970, n26971, n26972, n26973, n26974,
    n26975, n26976, n26977, n26978, n26979, n26980,
    n26981, n26982, n26983, n26984, n26985, n26986,
    n26987, n26988, n26989, n26990, n26991, n26992,
    n26993, n26994, n26995, n26996, n26997, n26998,
    n26999, n27000, n27001, n27002, n27003, n27004,
    n27005, n27006, n27007, n27008, n27009, n27010,
    n27011, n27012, n27014, n27015, n27016, n27017,
    n27018, n27019, n27020, n27021, n27022, n27023,
    n27024, n27025, n27026, n27027, n27028, n27029,
    n27030, n27031, n27032, n27033, n27034, n27035,
    n27036, n27037, n27038, n27039, n27040, n27041,
    n27042, n27043, n27044, n27045, n27046, n27047,
    n27048, n27049, n27050, n27051, n27052, n27053,
    n27054, n27055, n27056, n27057, n27058, n27059,
    n27060, n27061, n27062, n27063, n27064, n27065,
    n27066, n27067, n27068, n27069, n27070, n27071,
    n27072, n27073, n27074, n27075, n27076, n27077,
    n27078, n27079, n27080, n27081, n27082, n27083,
    n27084, n27085, n27086, n27087, n27088, n27089,
    n27090, n27091, n27092, n27093, n27094, n27095,
    n27096, n27097, n27098, n27099, n27100, n27101,
    n27102, n27103, n27104, n27105, n27106, n27107,
    n27108, n27109, n27110, n27111, n27112, n27113,
    n27114, n27115, n27116, n27117, n27118, n27119,
    n27120, n27121, n27122, n27123, n27124, n27125,
    n27126, n27127, n27128, n27129, n27130, n27131,
    n27132, n27133, n27134, n27135, n27136, n27137,
    n27138, n27139, n27140, n27141, n27142, n27143,
    n27144, n27145, n27146, n27147, n27148, n27149,
    n27150, n27151, n27152, n27153, n27154, n27155,
    n27156, n27157, n27158, n27159, n27160, n27161,
    n27162, n27163, n27164, n27165, n27166, n27167,
    n27168, n27169, n27170, n27171, n27172, n27173,
    n27174, n27175, n27176, n27177, n27178, n27179,
    n27180, n27181, n27182, n27183, n27184, n27185,
    n27186, n27187, n27188, n27189, n27190, n27191,
    n27192, n27193, n27194, n27195, n27196, n27197,
    n27198, n27199, n27200, n27201, n27202, n27203,
    n27204, n27205, n27206, n27207, n27208, n27209,
    n27210, n27211, n27212, n27213, n27214, n27215,
    n27216, n27217, n27218, n27219, n27220, n27221,
    n27222, n27223, n27224, n27225, n27226, n27227,
    n27228, n27229, n27230, n27231, n27232, n27233,
    n27234, n27235, n27236, n27237, n27238, n27239,
    n27240, n27241, n27242, n27243, n27244, n27245,
    n27246, n27247, n27248, n27249, n27250, n27251,
    n27252, n27253, n27254, n27255, n27256, n27257,
    n27258, n27259, n27260, n27261, n27262, n27263,
    n27264, n27265, n27266, n27267, n27268, n27269,
    n27270, n27271, n27272, n27273, n27274, n27275,
    n27276, n27277, n27278, n27279, n27280, n27281,
    n27282, n27283, n27284, n27285, n27286, n27287,
    n27288, n27289, n27290, n27291, n27292, n27293,
    n27294, n27295, n27296, n27297, n27298, n27299,
    n27300, n27301, n27302, n27303, n27304, n27305,
    n27306, n27307, n27308, n27309, n27310, n27311,
    n27312, n27313, n27314, n27315, n27316, n27317,
    n27318, n27319, n27320, n27321, n27322, n27323,
    n27324, n27325, n27326, n27327, n27328, n27329,
    n27330, n27331, n27332, n27333, n27334, n27335,
    n27336, n27337, n27338, n27339, n27340, n27341,
    n27342, n27343, n27344, n27345, n27346, n27347,
    n27348, n27349, n27350, n27351, n27352, n27353,
    n27354, n27355, n27356, n27357, n27358, n27359,
    n27360, n27361, n27362, n27363, n27364, n27365,
    n27366, n27367, n27368, n27369, n27370, n27371,
    n27372, n27373, n27374, n27375, n27376, n27377,
    n27378, n27379, n27380, n27381, n27382, n27383,
    n27384, n27385, n27386, n27387, n27388, n27389,
    n27390, n27391, n27392, n27393, n27394, n27395,
    n27396, n27397, n27398, n27399, n27400, n27401,
    n27402, n27403, n27404, n27405, n27406, n27407,
    n27408, n27409, n27410, n27411, n27412, n27413,
    n27414, n27415, n27416, n27417, n27418, n27419,
    n27420, n27421, n27422, n27423, n27424, n27425,
    n27426, n27427, n27428, n27429, n27430, n27431,
    n27432, n27433, n27434, n27435, n27436, n27437,
    n27438, n27439, n27440, n27441, n27442, n27443,
    n27444, n27445, n27446, n27447, n27448, n27449,
    n27450, n27451, n27452, n27453, n27454, n27455,
    n27456, n27457, n27458, n27459, n27460, n27461,
    n27462, n27463, n27465, n27466, n27467, n27468,
    n27469, n27470, n27471, n27472, n27473, n27474,
    n27475, n27476, n27477, n27478, n27479, n27480,
    n27481, n27482, n27483, n27484, n27485, n27486,
    n27487, n27488, n27489, n27490, n27491, n27492,
    n27493, n27494, n27495, n27496, n27497, n27498,
    n27499, n27500, n27501, n27502, n27503, n27504,
    n27505, n27506, n27507, n27508, n27509, n27510,
    n27511, n27512, n27513, n27514, n27515, n27516,
    n27517, n27518, n27519, n27520, n27521, n27522,
    n27523, n27524, n27525, n27526, n27527, n27528,
    n27529, n27530, n27531, n27532, n27533, n27534,
    n27535, n27536, n27537, n27538, n27539, n27540,
    n27541, n27542, n27543, n27544, n27545, n27546,
    n27547, n27548, n27549, n27550, n27551, n27552,
    n27553, n27554, n27555, n27556, n27557, n27558,
    n27559, n27560, n27561, n27562, n27563, n27564,
    n27565, n27566, n27567, n27568, n27569, n27570,
    n27571, n27572, n27573, n27574, n27575, n27576,
    n27577, n27578, n27579, n27580, n27581, n27582,
    n27583, n27584, n27585, n27586, n27587, n27588,
    n27589, n27590, n27591, n27592, n27593, n27594,
    n27595, n27596, n27597, n27598, n27599, n27600,
    n27601, n27602, n27603, n27604, n27605, n27606,
    n27607, n27608, n27609, n27610, n27611, n27612,
    n27613, n27614, n27615, n27616, n27617, n27618,
    n27619, n27620, n27621, n27622, n27623, n27624,
    n27625, n27626, n27627, n27628, n27629, n27630,
    n27631, n27632, n27633, n27634, n27635, n27636,
    n27637, n27638, n27639, n27640, n27641, n27642,
    n27643, n27644, n27645, n27646, n27647, n27648,
    n27649, n27650, n27651, n27652, n27653, n27654,
    n27655, n27656, n27657, n27658, n27659, n27660,
    n27661, n27662, n27663, n27664, n27665, n27666,
    n27667, n27668, n27669, n27670, n27671, n27672,
    n27673, n27674, n27675, n27676, n27677, n27678,
    n27679, n27680, n27681, n27682, n27683, n27684,
    n27685, n27686, n27687, n27688, n27689, n27690,
    n27691, n27692, n27693, n27694, n27695, n27696,
    n27697, n27698, n27699, n27700, n27701, n27702,
    n27703, n27704, n27705, n27706, n27707, n27708,
    n27709, n27710, n27711, n27712, n27713, n27714,
    n27715, n27716, n27717, n27718, n27719, n27720,
    n27721, n27722, n27723, n27724, n27725, n27726,
    n27727, n27728, n27729, n27730, n27731, n27732,
    n27733, n27734, n27735, n27736, n27737, n27738,
    n27739, n27740, n27741, n27742, n27743, n27744,
    n27745, n27746, n27747, n27748, n27749, n27750,
    n27751, n27752, n27753, n27754, n27755, n27756,
    n27757, n27758, n27759, n27760, n27761, n27762,
    n27763, n27764, n27765, n27766, n27767, n27768,
    n27769, n27770, n27771, n27772, n27773, n27774,
    n27775, n27776, n27777, n27778, n27779, n27780,
    n27781, n27782, n27783, n27784, n27785, n27786,
    n27787, n27788, n27789, n27790, n27791, n27792,
    n27793, n27794, n27795, n27796, n27797, n27798,
    n27799, n27800, n27801, n27802, n27803, n27804,
    n27805, n27806, n27807, n27808, n27809, n27810,
    n27811, n27812, n27813, n27814, n27815, n27816,
    n27817, n27818, n27819, n27820, n27821, n27822,
    n27823, n27824, n27825, n27826, n27827, n27828,
    n27829, n27830, n27831, n27832, n27833, n27834,
    n27835, n27836, n27837, n27838, n27839, n27840,
    n27841, n27842, n27843, n27844, n27845, n27846,
    n27847, n27848, n27849, n27850, n27851, n27852,
    n27853, n27854, n27855, n27856, n27857, n27858,
    n27859, n27860, n27861, n27862, n27863, n27864,
    n27865, n27866, n27867, n27868, n27869, n27870,
    n27871, n27872, n27873, n27874, n27875, n27876,
    n27877, n27878, n27879, n27880, n27881, n27882,
    n27883, n27884, n27885, n27886, n27887, n27888,
    n27889, n27890, n27891, n27892, n27893, n27894,
    n27895, n27896, n27897, n27898, n27899, n27900,
    n27901, n27902, n27903, n27904, n27905, n27906,
    n27907, n27908, n27909, n27910, n27911, n27912,
    n27914, n27915, n27916, n27917, n27918, n27919,
    n27920, n27921, n27922, n27923, n27924, n27925,
    n27926, n27927, n27928, n27929, n27930, n27931,
    n27932, n27933, n27934, n27935, n27936, n27937,
    n27938, n27939, n27940, n27941, n27942, n27943,
    n27944, n27945, n27946, n27947, n27948, n27949,
    n27950, n27951, n27952, n27953, n27954, n27955,
    n27956, n27957, n27958, n27959, n27960, n27961,
    n27962, n27963, n27964, n27965, n27966, n27967,
    n27968, n27969, n27970, n27971, n27972, n27973,
    n27974, n27975, n27976, n27977, n27978, n27979,
    n27980, n27981, n27982, n27983, n27984, n27985,
    n27986, n27987, n27988, n27989, n27990, n27991,
    n27992, n27993, n27994, n27995, n27996, n27997,
    n27998, n27999, n28000, n28001, n28002, n28003,
    n28004, n28005, n28006, n28007, n28008, n28009,
    n28010, n28011, n28012, n28013, n28014, n28015,
    n28016, n28017, n28018, n28019, n28020, n28021,
    n28022, n28023, n28024, n28025, n28026, n28027,
    n28028, n28029, n28030, n28031, n28032, n28033,
    n28034, n28035, n28036, n28037, n28038, n28039,
    n28040, n28041, n28042, n28043, n28044, n28045,
    n28046, n28047, n28048, n28049, n28050, n28051,
    n28052, n28053, n28054, n28055, n28056, n28057,
    n28058, n28059, n28060, n28061, n28062, n28063,
    n28064, n28065, n28066, n28067, n28068, n28069,
    n28070, n28071, n28072, n28073, n28074, n28075,
    n28076, n28077, n28078, n28079, n28080, n28081,
    n28082, n28083, n28084, n28085, n28086, n28087,
    n28088, n28089, n28090, n28091, n28092, n28093,
    n28094, n28095, n28096, n28097, n28098, n28099,
    n28100, n28101, n28102, n28103, n28104, n28105,
    n28106, n28107, n28108, n28109, n28110, n28111,
    n28112, n28113, n28114, n28115, n28116, n28117,
    n28118, n28119, n28120, n28121, n28122, n28123,
    n28124, n28125, n28126, n28127, n28128, n28129,
    n28130, n28131, n28132, n28133, n28134, n28135,
    n28136, n28137, n28138, n28139, n28140, n28141,
    n28142, n28143, n28144, n28145, n28146, n28147,
    n28148, n28149, n28150, n28151, n28152, n28153,
    n28154, n28155, n28156, n28157, n28158, n28159,
    n28160, n28161, n28162, n28163, n28164, n28165,
    n28166, n28167, n28168, n28169, n28170, n28171,
    n28172, n28173, n28174, n28175, n28176, n28177,
    n28178, n28179, n28180, n28181, n28182, n28183,
    n28184, n28185, n28186, n28187, n28188, n28189,
    n28190, n28191, n28192, n28193, n28194, n28195,
    n28196, n28197, n28198, n28199, n28200, n28201,
    n28202, n28203, n28204, n28205, n28206, n28207,
    n28208, n28209, n28210, n28211, n28212, n28213,
    n28214, n28215, n28216, n28217, n28218, n28219,
    n28220, n28221, n28222, n28223, n28224, n28225,
    n28226, n28227, n28228, n28229, n28230, n28231,
    n28232, n28233, n28234, n28235, n28236, n28237,
    n28238, n28239, n28240, n28241, n28242, n28243,
    n28244, n28245, n28246, n28247, n28248, n28249,
    n28250, n28251, n28252, n28253, n28254, n28255,
    n28256, n28257, n28258, n28259, n28260, n28261,
    n28262, n28263, n28264, n28265, n28266, n28267,
    n28268, n28269, n28270, n28271, n28272, n28273,
    n28274, n28275, n28276, n28277, n28278, n28279,
    n28280, n28281, n28282, n28283, n28284, n28285,
    n28286, n28287, n28288, n28289, n28290, n28291,
    n28292, n28293, n28294, n28295, n28296, n28297,
    n28298, n28299, n28300, n28301, n28302, n28303,
    n28304, n28305, n28306, n28307, n28308, n28309,
    n28310, n28311, n28312, n28313, n28314, n28315,
    n28316, n28317, n28318, n28319, n28320, n28321,
    n28322, n28323, n28324, n28325, n28326, n28327,
    n28328, n28329, n28330, n28331, n28332, n28333,
    n28334, n28335, n28336, n28337, n28338, n28339,
    n28340, n28341, n28342, n28343, n28344, n28345,
    n28346, n28347, n28348, n28349, n28350, n28351,
    n28352, n28353, n28354, n28355, n28356, n28357,
    n28358, n28359, n28360, n28362, n28363, n28364,
    n28365, n28366, n28367, n28368, n28369, n28370,
    n28371, n28372, n28373, n28374, n28375, n28376,
    n28377, n28378, n28379, n28380, n28381, n28382,
    n28383, n28384, n28385, n28386, n28387, n28388,
    n28389, n28390, n28391, n28392, n28393, n28394,
    n28395, n28396, n28397, n28398, n28399, n28400,
    n28401, n28402, n28403, n28404, n28405, n28406,
    n28407, n28408, n28409, n28410, n28411, n28412,
    n28413, n28414, n28415, n28416, n28417, n28418,
    n28419, n28420, n28421, n28422, n28423, n28424,
    n28425, n28426, n28427, n28428, n28429, n28430,
    n28431, n28432, n28433, n28434, n28435, n28436,
    n28437, n28438, n28439, n28440, n28441, n28442,
    n28443, n28444, n28445, n28446, n28447, n28448,
    n28449, n28450, n28451, n28452, n28453, n28454,
    n28455, n28456, n28457, n28458, n28459, n28460,
    n28461, n28462, n28463, n28464, n28465, n28466,
    n28467, n28468, n28469, n28470, n28471, n28472,
    n28473, n28474, n28475, n28476, n28477, n28478,
    n28479, n28480, n28481, n28482, n28483, n28484,
    n28485, n28486, n28487, n28488, n28489, n28490,
    n28491, n28492, n28493, n28494, n28495, n28496,
    n28497, n28498, n28499, n28500, n28501, n28502,
    n28503, n28504, n28505, n28506, n28507, n28508,
    n28509, n28510, n28511, n28512, n28513, n28514,
    n28515, n28516, n28517, n28518, n28519, n28520,
    n28521, n28522, n28523, n28524, n28525, n28526,
    n28527, n28528, n28529, n28530, n28531, n28532,
    n28533, n28534, n28535, n28536, n28537, n28538,
    n28539, n28540, n28541, n28542, n28543, n28544,
    n28545, n28546, n28547, n28548, n28549, n28550,
    n28551, n28552, n28553, n28554, n28555, n28556,
    n28557, n28558, n28559, n28560, n28561, n28562,
    n28563, n28564, n28565, n28566, n28567, n28568,
    n28569, n28570, n28571, n28572, n28573, n28574,
    n28575, n28576, n28577, n28578, n28579, n28580,
    n28581, n28582, n28583, n28584, n28585, n28586,
    n28587, n28588, n28589, n28590, n28591, n28592,
    n28593, n28594, n28595, n28596, n28597, n28598,
    n28599, n28600, n28601, n28602, n28603, n28604,
    n28605, n28606, n28607, n28608, n28609, n28610,
    n28611, n28612, n28613, n28614, n28615, n28616,
    n28617, n28618, n28619, n28620, n28621, n28622,
    n28623, n28624, n28625, n28626, n28627, n28628,
    n28629, n28630, n28631, n28632, n28633, n28634,
    n28635, n28636, n28637, n28638, n28639, n28640,
    n28641, n28642, n28643, n28644, n28645, n28646,
    n28647, n28648, n28649, n28650, n28651, n28652,
    n28653, n28654, n28655, n28656, n28657, n28658,
    n28659, n28660, n28661, n28662, n28663, n28664,
    n28665, n28666, n28667, n28668, n28669, n28670,
    n28671, n28672, n28673, n28674, n28675, n28676,
    n28677, n28678, n28679, n28680, n28681, n28682,
    n28683, n28684, n28685, n28686, n28687, n28688,
    n28689, n28690, n28691, n28692, n28693, n28694,
    n28695, n28696, n28697, n28698, n28699, n28700,
    n28701, n28702, n28703, n28704, n28705, n28706,
    n28707, n28708, n28709, n28710, n28711, n28712,
    n28713, n28714, n28715, n28716, n28717, n28718,
    n28719, n28720, n28721, n28722, n28723, n28724,
    n28725, n28726, n28727, n28728, n28729, n28730,
    n28731, n28732, n28733, n28734, n28735, n28736,
    n28737, n28738, n28739, n28740, n28741, n28742,
    n28743, n28744, n28745, n28746, n28747, n28748,
    n28749, n28750, n28751, n28752, n28753, n28754,
    n28755, n28756, n28757, n28758, n28759, n28760,
    n28761, n28762, n28763, n28764, n28765, n28766,
    n28767, n28768, n28769, n28770, n28771, n28772,
    n28773, n28774, n28775, n28776, n28777, n28778,
    n28779, n28780, n28781, n28782, n28783, n28784,
    n28785, n28786, n28787, n28788, n28789, n28790,
    n28791, n28792, n28793, n28794, n28795, n28796,
    n28797, n28798, n28799, n28800, n28801, n28802,
    n28803, n28804, n28805, n28806, n28807, n28808,
    n28809, n28811, n28812, n28813, n28814, n28815,
    n28816, n28817, n28818, n28819, n28820, n28821,
    n28822, n28823, n28824, n28825, n28826, n28827,
    n28828, n28829, n28830, n28831, n28832, n28833,
    n28834, n28835, n28836, n28837, n28838, n28839,
    n28840, n28841, n28842, n28843, n28844, n28845,
    n28846, n28847, n28848, n28849, n28850, n28851,
    n28852, n28853, n28854, n28855, n28856, n28857,
    n28858, n28859, n28860, n28861, n28862, n28863,
    n28864, n28865, n28866, n28867, n28868, n28869,
    n28870, n28871, n28872, n28873, n28874, n28875,
    n28876, n28877, n28878, n28879, n28880, n28881,
    n28882, n28883, n28884, n28885, n28886, n28887,
    n28888, n28889, n28890, n28891, n28892, n28893,
    n28894, n28895, n28896, n28897, n28898, n28899,
    n28900, n28901, n28902, n28903, n28904, n28905,
    n28906, n28907, n28908, n28909, n28910, n28911,
    n28912, n28913, n28914, n28915, n28916, n28917,
    n28918, n28919, n28920, n28921, n28922, n28923,
    n28924, n28925, n28926, n28927, n28928, n28929,
    n28930, n28931, n28932, n28933, n28934, n28935,
    n28936, n28937, n28938, n28939, n28940, n28941,
    n28942, n28943, n28944, n28945, n28946, n28947,
    n28948, n28949, n28950, n28951, n28952, n28953,
    n28954, n28955, n28956, n28957, n28958, n28959,
    n28960, n28961, n28962, n28963, n28964, n28965,
    n28966, n28967, n28968, n28969, n28970, n28971,
    n28972, n28973, n28974, n28975, n28976, n28977,
    n28978, n28979, n28980, n28981, n28982, n28983,
    n28984, n28985, n28986, n28987, n28988, n28989,
    n28990, n28991, n28992, n28993, n28994, n28995,
    n28996, n28997, n28998, n28999, n29000, n29001,
    n29002, n29003, n29004, n29005, n29006, n29007,
    n29008, n29009, n29010, n29011, n29012, n29013,
    n29014, n29015, n29016, n29017, n29018, n29019,
    n29020, n29021, n29022, n29023, n29024, n29025,
    n29026, n29027, n29028, n29029, n29030, n29031,
    n29032, n29033, n29034, n29035, n29036, n29037,
    n29038, n29039, n29040, n29041, n29042, n29043,
    n29044, n29045, n29046, n29047, n29048, n29049,
    n29050, n29051, n29052, n29053, n29054, n29055,
    n29056, n29057, n29058, n29059, n29060, n29061,
    n29062, n29063, n29064, n29065, n29066, n29067,
    n29068, n29069, n29070, n29071, n29072, n29073,
    n29074, n29075, n29076, n29077, n29078, n29079,
    n29080, n29081, n29082, n29083, n29084, n29085,
    n29086, n29087, n29088, n29089, n29090, n29091,
    n29092, n29093, n29094, n29095, n29096, n29097,
    n29098, n29099, n29100, n29101, n29102, n29103,
    n29104, n29105, n29106, n29107, n29108, n29109,
    n29110, n29111, n29112, n29113, n29114, n29115,
    n29116, n29117, n29118, n29119, n29120, n29121,
    n29122, n29123, n29124, n29125, n29126, n29127,
    n29128, n29129, n29130, n29131, n29132, n29133,
    n29134, n29135, n29136, n29137, n29138, n29139,
    n29140, n29141, n29142, n29143, n29144, n29145,
    n29146, n29147, n29148, n29149, n29150, n29151,
    n29152, n29153, n29154, n29155, n29156, n29157,
    n29158, n29159, n29160, n29161, n29162, n29163,
    n29164, n29165, n29166, n29167, n29168, n29169,
    n29170, n29171, n29172, n29173, n29174, n29175,
    n29176, n29177, n29178, n29179, n29180, n29181,
    n29182, n29183, n29184, n29185, n29186, n29187,
    n29188, n29189, n29190, n29191, n29192, n29193,
    n29194, n29195, n29196, n29197, n29198, n29199,
    n29200, n29201, n29202, n29203, n29204, n29205,
    n29206, n29207, n29208, n29209, n29210, n29211,
    n29212, n29213, n29214, n29215, n29216, n29217,
    n29218, n29219, n29220, n29221, n29222, n29223,
    n29224, n29225, n29226, n29227, n29228, n29229,
    n29230, n29231, n29232, n29233, n29234, n29235,
    n29236, n29237, n29238, n29239, n29240, n29241,
    n29242, n29243, n29244, n29245, n29246, n29247,
    n29248, n29249, n29250, n29251, n29252, n29253,
    n29254, n29255, n29256, n29257, n29258, n29259,
    n29260, n29261, n29262, n29263, n29265, n29266,
    n29267, n29268, n29269, n29270, n29271, n29272,
    n29273, n29274, n29275, n29276, n29277, n29278,
    n29279, n29280, n29281, n29282, n29283, n29284,
    n29285, n29286, n29287, n29288, n29289, n29290,
    n29291, n29292, n29293, n29294, n29295, n29296,
    n29297, n29298, n29299, n29300, n29301, n29302,
    n29303, n29304, n29305, n29306, n29307, n29308,
    n29309, n29310, n29311, n29312, n29313, n29314,
    n29315, n29316, n29317, n29318, n29319, n29320,
    n29321, n29322, n29323, n29324, n29325, n29326,
    n29327, n29328, n29329, n29330, n29331, n29332,
    n29333, n29334, n29335, n29336, n29337, n29338,
    n29339, n29340, n29341, n29342, n29343, n29344,
    n29345, n29346, n29347, n29348, n29349, n29350,
    n29351, n29352, n29353, n29354, n29355, n29356,
    n29357, n29358, n29359, n29360, n29361, n29362,
    n29363, n29364, n29365, n29366, n29367, n29368,
    n29369, n29370, n29371, n29372, n29373, n29374,
    n29375, n29376, n29377, n29378, n29379, n29380,
    n29381, n29382, n29383, n29384, n29385, n29386,
    n29387, n29388, n29389, n29390, n29391, n29392,
    n29393, n29394, n29395, n29396, n29397, n29398,
    n29399, n29400, n29401, n29402, n29403, n29404,
    n29405, n29406, n29407, n29408, n29409, n29410,
    n29411, n29412, n29413, n29414, n29415, n29416,
    n29417, n29418, n29419, n29420, n29421, n29422,
    n29423, n29424, n29425, n29426, n29427, n29428,
    n29429, n29430, n29431, n29432, n29433, n29434,
    n29435, n29436, n29437, n29438, n29439, n29440,
    n29441, n29442, n29443, n29444, n29445, n29446,
    n29447, n29448, n29449, n29450, n29451, n29452,
    n29453, n29454, n29455, n29456, n29457, n29458,
    n29459, n29460, n29461, n29462, n29463, n29464,
    n29465, n29466, n29467, n29468, n29469, n29470,
    n29471, n29472, n29473, n29474, n29475, n29476,
    n29477, n29478, n29479, n29480, n29481, n29482,
    n29483, n29484, n29485, n29486, n29487, n29488,
    n29489, n29490, n29491, n29492, n29493, n29494,
    n29495, n29496, n29497, n29498, n29499, n29500,
    n29501, n29502, n29503, n29504, n29505, n29506,
    n29507, n29508, n29509, n29510, n29511, n29512,
    n29513, n29514, n29515, n29516, n29517, n29518,
    n29519, n29520, n29521, n29522, n29523, n29524,
    n29525, n29526, n29527, n29528, n29529, n29530,
    n29531, n29532, n29533, n29534, n29535, n29536,
    n29537, n29538, n29539, n29540, n29541, n29542,
    n29543, n29544, n29545, n29546, n29547, n29548,
    n29549, n29550, n29551, n29552, n29553, n29554,
    n29555, n29556, n29557, n29558, n29559, n29560,
    n29561, n29562, n29563, n29564, n29565, n29566,
    n29567, n29568, n29569, n29570, n29571, n29572,
    n29573, n29574, n29575, n29576, n29577, n29578,
    n29579, n29580, n29581, n29582, n29583, n29584,
    n29585, n29586, n29587, n29588, n29589, n29590,
    n29591, n29592, n29593, n29594, n29595, n29596,
    n29597, n29598, n29599, n29600, n29601, n29602,
    n29603, n29604, n29605, n29606, n29607, n29608,
    n29609, n29610, n29611, n29612, n29613, n29614,
    n29615, n29616, n29617, n29618, n29619, n29620,
    n29621, n29622, n29623, n29624, n29625, n29626,
    n29627, n29628, n29629, n29630, n29631, n29632,
    n29633, n29634, n29635, n29636, n29637, n29638,
    n29639, n29640, n29641, n29642, n29643, n29644,
    n29645, n29646, n29647, n29648, n29649, n29650,
    n29651, n29652, n29653, n29654, n29655, n29656,
    n29657, n29658, n29659, n29660, n29661, n29662,
    n29663, n29664, n29665, n29666, n29667, n29668,
    n29669, n29670, n29671, n29672, n29673, n29674,
    n29675, n29676, n29677, n29678, n29679, n29680,
    n29681, n29682, n29683, n29684, n29685, n29686,
    n29687, n29688, n29689, n29690, n29691, n29692,
    n29693, n29694, n29695, n29696, n29697, n29698,
    n29699, n29700, n29701, n29702, n29703, n29704,
    n29705, n29706, n29707, n29708, n29709, n29710,
    n29711, n29712, n29713, n29714, n29715, n29716,
    n29717, n29718, n29720, n29721, n29722, n29723,
    n29724, n29725, n29726, n29727, n29728, n29729,
    n29730, n29731, n29732, n29733, n29734, n29735,
    n29736, n29737, n29738, n29739, n29740, n29741,
    n29742, n29743, n29744, n29745, n29746, n29747,
    n29748, n29749, n29750, n29751, n29752, n29753,
    n29754, n29755, n29756, n29757, n29758, n29759,
    n29760, n29761, n29762, n29763, n29764, n29765,
    n29766, n29767, n29768, n29769, n29770, n29771,
    n29772, n29773, n29774, n29775, n29776, n29777,
    n29778, n29779, n29780, n29781, n29782, n29783,
    n29784, n29785, n29786, n29787, n29788, n29789,
    n29790, n29791, n29792, n29793, n29794, n29795,
    n29796, n29797, n29798, n29799, n29800, n29801,
    n29802, n29803, n29804, n29805, n29806, n29807,
    n29808, n29809, n29810, n29811, n29812, n29813,
    n29814, n29815, n29816, n29817, n29818, n29819,
    n29820, n29821, n29822, n29823, n29824, n29825,
    n29826, n29827, n29828, n29829, n29830, n29831,
    n29832, n29833, n29834, n29835, n29836, n29837,
    n29838, n29839, n29840, n29841, n29842, n29843,
    n29844, n29845, n29846, n29847, n29848, n29849,
    n29850, n29851, n29852, n29853, n29854, n29855,
    n29856, n29857, n29858, n29859, n29860, n29861,
    n29862, n29863, n29864, n29865, n29866, n29867,
    n29868, n29869, n29870, n29871, n29872, n29873,
    n29874, n29875, n29876, n29877, n29878, n29879,
    n29880, n29881, n29882, n29883, n29884, n29885,
    n29886, n29887, n29888, n29889, n29890, n29891,
    n29892, n29893, n29894, n29895, n29896, n29897,
    n29898, n29899, n29900, n29901, n29902, n29903,
    n29904, n29905, n29906, n29907, n29908, n29909,
    n29910, n29911, n29912, n29913, n29914, n29915,
    n29916, n29917, n29918, n29919, n29920, n29921,
    n29922, n29923, n29924, n29925, n29926, n29927,
    n29928, n29929, n29930, n29931, n29932, n29933,
    n29934, n29935, n29936, n29937, n29938, n29939,
    n29940, n29941, n29942, n29943, n29944, n29945,
    n29946, n29947, n29948, n29949, n29950, n29951,
    n29952, n29953, n29954, n29955, n29956, n29957,
    n29958, n29959, n29960, n29961, n29962, n29963,
    n29964, n29965, n29966, n29967, n29968, n29969,
    n29970, n29971, n29972, n29973, n29974, n29975,
    n29976, n29977, n29978, n29979, n29980, n29981,
    n29982, n29983, n29984, n29985, n29986, n29987,
    n29988, n29989, n29990, n29991, n29992, n29993,
    n29994, n29995, n29996, n29997, n29998, n29999,
    n30000, n30001, n30002, n30003, n30004, n30005,
    n30006, n30007, n30008, n30009, n30010, n30011,
    n30012, n30013, n30014, n30015, n30016, n30017,
    n30018, n30019, n30020, n30021, n30022, n30023,
    n30024, n30025, n30026, n30027, n30028, n30029,
    n30030, n30031, n30032, n30033, n30034, n30035,
    n30036, n30037, n30038, n30039, n30040, n30041,
    n30042, n30043, n30044, n30045, n30046, n30047,
    n30048, n30049, n30050, n30051, n30052, n30053,
    n30054, n30055, n30056, n30057, n30058, n30059,
    n30060, n30061, n30062, n30063, n30064, n30065,
    n30066, n30067, n30068, n30069, n30070, n30071,
    n30072, n30073, n30074, n30075, n30076, n30077,
    n30078, n30079, n30080, n30081, n30082, n30083,
    n30084, n30085, n30086, n30087, n30088, n30089,
    n30090, n30091, n30092, n30093, n30094, n30095,
    n30096, n30097, n30098, n30099, n30100, n30101,
    n30102, n30103, n30104, n30105, n30106, n30107,
    n30108, n30109, n30110, n30111, n30112, n30113,
    n30114, n30115, n30116, n30117, n30118, n30119,
    n30120, n30121, n30122, n30123, n30124, n30125,
    n30126, n30127, n30128, n30129, n30130, n30131,
    n30132, n30133, n30134, n30135, n30136, n30137,
    n30138, n30139, n30140, n30141, n30142, n30143,
    n30144, n30145, n30146, n30147, n30148, n30149,
    n30150, n30151, n30152, n30153, n30154, n30155,
    n30156, n30157, n30158, n30159, n30160, n30161,
    n30162, n30163, n30164, n30165, n30166, n30167,
    n30168, n30169, n30170, n30171, n30172, n30173,
    n30175, n30176, n30177, n30178, n30179, n30180,
    n30181, n30182, n30183, n30184, n30185, n30186,
    n30187, n30188, n30189, n30190, n30191, n30192,
    n30193, n30194, n30195, n30196, n30197, n30198,
    n30199, n30200, n30201, n30202, n30203, n30204,
    n30205, n30206, n30207, n30208, n30209, n30210,
    n30211, n30212, n30213, n30214, n30215, n30216,
    n30217, n30218, n30219, n30220, n30221, n30222,
    n30223, n30224, n30225, n30226, n30227, n30228,
    n30229, n30230, n30231, n30232, n30233, n30234,
    n30235, n30236, n30237, n30238, n30239, n30240,
    n30241, n30242, n30243, n30244, n30245, n30246,
    n30247, n30248, n30249, n30250, n30251, n30252,
    n30253, n30254, n30255, n30256, n30257, n30258,
    n30259, n30260, n30261, n30262, n30263, n30264,
    n30265, n30266, n30267, n30268, n30269, n30270,
    n30271, n30272, n30273, n30274, n30275, n30276,
    n30277, n30278, n30279, n30280, n30281, n30282,
    n30283, n30284, n30285, n30286, n30287, n30288,
    n30289, n30290, n30291, n30292, n30293, n30294,
    n30295, n30296, n30297, n30298, n30299, n30300,
    n30301, n30302, n30303, n30304, n30305, n30306,
    n30307, n30308, n30309, n30310, n30311, n30312,
    n30313, n30314, n30315, n30316, n30317, n30318,
    n30319, n30320, n30321, n30322, n30323, n30324,
    n30325, n30326, n30327, n30328, n30329, n30330,
    n30331, n30332, n30333, n30334, n30335, n30336,
    n30337, n30338, n30339, n30340, n30341, n30342,
    n30343, n30344, n30345, n30346, n30347, n30348,
    n30349, n30350, n30351, n30352, n30353, n30354,
    n30355, n30356, n30357, n30358, n30359, n30360,
    n30361, n30362, n30363, n30364, n30365, n30366,
    n30367, n30368, n30369, n30370, n30371, n30372,
    n30373, n30374, n30375, n30376, n30377, n30378,
    n30379, n30380, n30381, n30382, n30383, n30384,
    n30385, n30386, n30387, n30388, n30389, n30390,
    n30391, n30392, n30393, n30394, n30395, n30396,
    n30397, n30398, n30399, n30400, n30401, n30402,
    n30403, n30404, n30405, n30406, n30407, n30408,
    n30409, n30410, n30411, n30412, n30413, n30414,
    n30415, n30416, n30417, n30418, n30419, n30420,
    n30421, n30422, n30423, n30424, n30425, n30426,
    n30427, n30428, n30429, n30430, n30431, n30432,
    n30433, n30434, n30435, n30436, n30437, n30438,
    n30439, n30440, n30441, n30442, n30443, n30444,
    n30445, n30446, n30447, n30448, n30449, n30450,
    n30451, n30452, n30453, n30454, n30455, n30456,
    n30457, n30458, n30459, n30460, n30461, n30462,
    n30463, n30464, n30465, n30466, n30467, n30468,
    n30469, n30470, n30471, n30472, n30473, n30474,
    n30475, n30476, n30477, n30478, n30479, n30480,
    n30481, n30482, n30483, n30484, n30485, n30486,
    n30487, n30488, n30489, n30490, n30491, n30492,
    n30493, n30494, n30495, n30496, n30497, n30498,
    n30499, n30500, n30501, n30502, n30503, n30504,
    n30505, n30506, n30507, n30508, n30509, n30510,
    n30511, n30512, n30513, n30514, n30515, n30516,
    n30517, n30518, n30519, n30520, n30521, n30522,
    n30523, n30524, n30525, n30526, n30527, n30528,
    n30529, n30530, n30531, n30532, n30533, n30534,
    n30535, n30536, n30537, n30538, n30539, n30540,
    n30541, n30542, n30543, n30544, n30545, n30546,
    n30547, n30548, n30549, n30550, n30551, n30552,
    n30553, n30554, n30555, n30556, n30557, n30558,
    n30559, n30560, n30561, n30562, n30563, n30564,
    n30565, n30566, n30567, n30568, n30569, n30570,
    n30571, n30572, n30573, n30574, n30575, n30576,
    n30577, n30578, n30579, n30580, n30581, n30582,
    n30583, n30584, n30585, n30586, n30587, n30588,
    n30589, n30590, n30591, n30592, n30593, n30594,
    n30595, n30596, n30597, n30598, n30599, n30600,
    n30601, n30602, n30603, n30604, n30605, n30606,
    n30607, n30608, n30609, n30610, n30611, n30612,
    n30613, n30614, n30615, n30616, n30617, n30618,
    n30619, n30620, n30621, n30622, n30623, n30624,
    n30625, n30626, n30627, n30628, n30630, n30631,
    n30632, n30633, n30634, n30635, n30636, n30637,
    n30638, n30639, n30640, n30641, n30642, n30643,
    n30644, n30645, n30646, n30647, n30648, n30649,
    n30650, n30651, n30652, n30653, n30654, n30655,
    n30656, n30657, n30658, n30659, n30660, n30661,
    n30662, n30663, n30664, n30665, n30666, n30667,
    n30668, n30669, n30670, n30671, n30672, n30673,
    n30674, n30675, n30676, n30677, n30678, n30679,
    n30680, n30681, n30682, n30683, n30684, n30685,
    n30686, n30687, n30688, n30689, n30690, n30691,
    n30692, n30693, n30694, n30695, n30696, n30697,
    n30698, n30699, n30700, n30701, n30702, n30703,
    n30704, n30705, n30706, n30707, n30708, n30709,
    n30710, n30711, n30712, n30713, n30714, n30715,
    n30716, n30717, n30718, n30719, n30720, n30721,
    n30722, n30723, n30724, n30725, n30726, n30727,
    n30728, n30729, n30730, n30731, n30732, n30733,
    n30734, n30735, n30736, n30737, n30738, n30739,
    n30740, n30741, n30742, n30743, n30744, n30745,
    n30746, n30747, n30748, n30749, n30750, n30751,
    n30752, n30753, n30754, n30755, n30756, n30757,
    n30758, n30759, n30760, n30761, n30762, n30763,
    n30764, n30765, n30766, n30767, n30768, n30769,
    n30770, n30771, n30772, n30773, n30774, n30775,
    n30776, n30777, n30778, n30779, n30780, n30781,
    n30782, n30783, n30784, n30785, n30786, n30787,
    n30788, n30789, n30790, n30791, n30792, n30793,
    n30794, n30795, n30796, n30797, n30798, n30799,
    n30800, n30801, n30802, n30803, n30804, n30805,
    n30806, n30807, n30808, n30809, n30810, n30811,
    n30812, n30813, n30814, n30815, n30816, n30817,
    n30818, n30819, n30820, n30821, n30822, n30823,
    n30824, n30825, n30826, n30827, n30828, n30829,
    n30830, n30831, n30832, n30833, n30834, n30835,
    n30836, n30837, n30838, n30839, n30840, n30841,
    n30842, n30843, n30844, n30845, n30846, n30847,
    n30848, n30849, n30850, n30851, n30852, n30853,
    n30854, n30855, n30856, n30857, n30858, n30859,
    n30860, n30861, n30862, n30863, n30864, n30865,
    n30866, n30867, n30868, n30869, n30870, n30871,
    n30872, n30873, n30874, n30875, n30876, n30877,
    n30878, n30879, n30880, n30881, n30882, n30883,
    n30884, n30885, n30886, n30887, n30888, n30889,
    n30890, n30891, n30892, n30893, n30894, n30895,
    n30896, n30897, n30898, n30899, n30900, n30901,
    n30902, n30903, n30904, n30905, n30906, n30907,
    n30908, n30909, n30910, n30911, n30912, n30913,
    n30914, n30915, n30916, n30917, n30918, n30919,
    n30920, n30921, n30922, n30923, n30924, n30925,
    n30926, n30927, n30928, n30929, n30930, n30931,
    n30932, n30933, n30934, n30935, n30936, n30937,
    n30938, n30939, n30940, n30941, n30942, n30943,
    n30944, n30945, n30946, n30947, n30948, n30949,
    n30950, n30951, n30952, n30953, n30954, n30955,
    n30956, n30957, n30958, n30959, n30960, n30961,
    n30962, n30963, n30964, n30965, n30966, n30967,
    n30968, n30969, n30970, n30971, n30972, n30973,
    n30974, n30975, n30976, n30977, n30978, n30979,
    n30980, n30981, n30982, n30983, n30984, n30985,
    n30986, n30987, n30988, n30989, n30990, n30991,
    n30992, n30993, n30994, n30995, n30996, n30997,
    n30998, n30999, n31000, n31001, n31002, n31003,
    n31004, n31005, n31006, n31007, n31008, n31009,
    n31010, n31011, n31012, n31013, n31014, n31015,
    n31016, n31017, n31018, n31019, n31020, n31021,
    n31022, n31023, n31024, n31025, n31026, n31027,
    n31028, n31029, n31030, n31031, n31032, n31033,
    n31034, n31035, n31036, n31037, n31038, n31039,
    n31040, n31041, n31042, n31043, n31044, n31045,
    n31046, n31047, n31048, n31049, n31050, n31051,
    n31052, n31053, n31054, n31055, n31056, n31057,
    n31058, n31059, n31060, n31061, n31062, n31063,
    n31064, n31065, n31066, n31067, n31068, n31069,
    n31070, n31071, n31072, n31073, n31074, n31075,
    n31077, n31078, n31079, n31080, n31081, n31082,
    n31083, n31084, n31085, n31086, n31087, n31088,
    n31089, n31090, n31091, n31092, n31093, n31094,
    n31095, n31096, n31097, n31098, n31099, n31100,
    n31101, n31102, n31103, n31104, n31105, n31106,
    n31107, n31108, n31109, n31110, n31111, n31112,
    n31113, n31114, n31115, n31116, n31117, n31118,
    n31119, n31120, n31121, n31122, n31123, n31124,
    n31125, n31126, n31127, n31128, n31129, n31130,
    n31131, n31132, n31133, n31134, n31135, n31136,
    n31137, n31138, n31139, n31140, n31141, n31142,
    n31143, n31144, n31145, n31146, n31147, n31148,
    n31149, n31150, n31151, n31152, n31153, n31154,
    n31155, n31156, n31157, n31158, n31159, n31160,
    n31161, n31162, n31163, n31164, n31165, n31166,
    n31167, n31168, n31169, n31170, n31171, n31172,
    n31173, n31174, n31175, n31176, n31177, n31178,
    n31179, n31180, n31181, n31182, n31183, n31184,
    n31185, n31186, n31187, n31188, n31189, n31190,
    n31191, n31192, n31193, n31194, n31195, n31196,
    n31197, n31198, n31199, n31200, n31201, n31202,
    n31203, n31204, n31205, n31206, n31207, n31208,
    n31209, n31210, n31211, n31212, n31213, n31214,
    n31215, n31216, n31217, n31218, n31219, n31220,
    n31221, n31222, n31223, n31224, n31225, n31226,
    n31227, n31228, n31229, n31230, n31231, n31232,
    n31233, n31234, n31235, n31236, n31237, n31238,
    n31239, n31240, n31241, n31242, n31243, n31244,
    n31245, n31246, n31247, n31248, n31249, n31250,
    n31251, n31252, n31253, n31254, n31255, n31256,
    n31257, n31258, n31259, n31260, n31261, n31262,
    n31263, n31264, n31265, n31266, n31267, n31268,
    n31269, n31270, n31271, n31272, n31273, n31274,
    n31275, n31276, n31277, n31278, n31279, n31280,
    n31281, n31282, n31283, n31284, n31285, n31286,
    n31287, n31288, n31289, n31290, n31291, n31292,
    n31293, n31294, n31295, n31296, n31297, n31298,
    n31299, n31300, n31301, n31302, n31303, n31304,
    n31305, n31306, n31307, n31308, n31309, n31310,
    n31311, n31312, n31313, n31314, n31315, n31316,
    n31317, n31318, n31319, n31320, n31321, n31322,
    n31323, n31324, n31325, n31326, n31327, n31328,
    n31329, n31330, n31331, n31332, n31333, n31334,
    n31335, n31336, n31337, n31338, n31339, n31340,
    n31341, n31342, n31343, n31344, n31345, n31346,
    n31347, n31348, n31349, n31350, n31351, n31352,
    n31353, n31354, n31355, n31356, n31357, n31358,
    n31359, n31360, n31361, n31362, n31363, n31364,
    n31365, n31366, n31367, n31368, n31369, n31370,
    n31371, n31372, n31373, n31374, n31375, n31376,
    n31377, n31378, n31379, n31380, n31381, n31382,
    n31383, n31384, n31385, n31386, n31387, n31388,
    n31389, n31390, n31391, n31392, n31393, n31394,
    n31395, n31396, n31397, n31398, n31399, n31400,
    n31401, n31402, n31403, n31404, n31405, n31406,
    n31407, n31408, n31409, n31410, n31411, n31412,
    n31413, n31414, n31415, n31416, n31417, n31418,
    n31419, n31420, n31421, n31422, n31423, n31424,
    n31425, n31426, n31427, n31428, n31429, n31430,
    n31431, n31432, n31433, n31434, n31435, n31436,
    n31437, n31438, n31439, n31440, n31441, n31442,
    n31443, n31444, n31445, n31446, n31447, n31448,
    n31449, n31450, n31451, n31452, n31453, n31454,
    n31455, n31456, n31457, n31458, n31459, n31460,
    n31461, n31462, n31463, n31464, n31465, n31466,
    n31467, n31468, n31469, n31470, n31471, n31472,
    n31473, n31474, n31475, n31476, n31477, n31478,
    n31479, n31480, n31481, n31482, n31483, n31484,
    n31485, n31486, n31487, n31488, n31489, n31490,
    n31491, n31492, n31493, n31494, n31495, n31496,
    n31497, n31498, n31499, n31500, n31501, n31502,
    n31503, n31504, n31505, n31506, n31507, n31508,
    n31509, n31510, n31511, n31512, n31513, n31514,
    n31515, n31516, n31517, n31519, n31520, n31521,
    n31522, n31523, n31524, n31525, n31526, n31527,
    n31528, n31529, n31530, n31531, n31532, n31533,
    n31534, n31535, n31536, n31537, n31538, n31539,
    n31540, n31541, n31542, n31543, n31544, n31545,
    n31546, n31547, n31548, n31549, n31550, n31551,
    n31552, n31553, n31554, n31555, n31556, n31557,
    n31558, n31559, n31560, n31561, n31562, n31563,
    n31564, n31565, n31566, n31567, n31569, n31570,
    n31571, n31572, n31573, n31574, n31575, n31576,
    n31577, n31578, n31579, n31580, n31581, n31582,
    n31583, n31584, n31585, n31586, n31587, n31588,
    n31589, n31590, n31591, n31592, n31593, n31594,
    n31595, n31596, n31597, n31598, n31599, n31600,
    n31601, n31602, n31603, n31604, n31605, n31606,
    n31607, n31608, n31609, n31610, n31611, n31612,
    n31613, n31614, n31615, n31616, n31617, n31618,
    n31619, n31620, n31621, n31622, n31623, n31624,
    n31625, n31626, n31627, n31628, n31629, n31630,
    n31631, n31632, n31633, n31634, n31635, n31636,
    n31638, n31639, n31640, n31641, n31642, n31643,
    n31644, n31645, n31646, n31647, n31648, n31649,
    n31650, n31651, n31652, n31653, n31654, n31655,
    n31656, n31657, n31658, n31659, n31660, n31661,
    n31662, n31663, n31664, n31665, n31666, n31667,
    n31668, n31669, n31670, n31671, n31672, n31673,
    n31674, n31675, n31676, n31677, n31678, n31679,
    n31680, n31681, n31682, n31683, n31684, n31685,
    n31686, n31687, n31688, n31689, n31690, n31691,
    n31692, n31693, n31694, n31695, n31696, n31698,
    n31699, n31700, n31701, n31702, n31703, n31704,
    n31705, n31706, n31707, n31708, n31709, n31710,
    n31711, n31712, n31713, n31714, n31715, n31716,
    n31717, n31718, n31719, n31720, n31721, n31722,
    n31723, n31724, n31725, n31726, n31727, n31728,
    n31729, n31730, n31731, n31732, n31733, n31734,
    n31735, n31736, n31737, n31738, n31739, n31740,
    n31741, n31742, n31743, n31744, n31745, n31746,
    n31747, n31748, n31749, n31750, n31751, n31752,
    n31753, n31754, n31755, n31756, n31757, n31758,
    n31759, n31760, n31761, n31762, n31763, n31764,
    n31765, n31766, n31767, n31768, n31769, n31770,
    n31771, n31772, n31773, n31774, n31775, n31776,
    n31777, n31778, n31779, n31780, n31781, n31782,
    n31783, n31784, n31785, n31786, n31787, n31788,
    n31789, n31790, n31791, n31792, n31793, n31794,
    n31795, n31796, n31797, n31798, n31799, n31800,
    n31801, n31802, n31803, n31804, n31805, n31806,
    n31807, n31808, n31809, n31810, n31811, n31812,
    n31813, n31814, n31815, n31816, n31817, n31818,
    n31819, n31820, n31821, n31822, n31823, n31824,
    n31825, n31826, n31827, n31828, n31829, n31830,
    n31831, n31832, n31833, n31834, n31835, n31836,
    n31837, n31838, n31839, n31840, n31841, n31842,
    n31843, n31844, n31845, n31846, n31847, n31848,
    n31849, n31850, n31851, n31852, n31853, n31854,
    n31855, n31856, n31857, n31858, n31859, n31860,
    n31861, n31862, n31863, n31864, n31865, n31866,
    n31867, n31868, n31869, n31870, n31871, n31872,
    n31873, n31874, n31875, n31876, n31877, n31878,
    n31879, n31880, n31881, n31882, n31883, n31884,
    n31885, n31886, n31887, n31888, n31889, n31890,
    n31891, n31892, n31893, n31894, n31895, n31896,
    n31897, n31898, n31899, n31900, n31901, n31902,
    n31903, n31904, n31905, n31906, n31907, n31908,
    n31909, n31910, n31911, n31912, n31913, n31914,
    n31915, n31916, n31917, n31918, n31919, n31920,
    n31921, n31922, n31923, n31924, n31925, n31926,
    n31927, n31928, n31929, n31930, n31931, n31932,
    n31933, n31934, n31935, n31936, n31937, n31938,
    n31939, n31940, n31941, n31942, n31943, n31944,
    n31945, n31946, n31947, n31948, n31949, n31950,
    n31951, n31952, n31953, n31954, n31955, n31956,
    n31957, n31958, n31959, n31960, n31961, n31962,
    n31963, n31964, n31965, n31966, n31967, n31968,
    n31969, n31970, n31971, n31972, n31973, n31974,
    n31975, n31976, n31977, n31978, n31979, n31980,
    n31981, n31982, n31983, n31984, n31985, n31986,
    n31987, n31988, n31989, n31990, n31991, n31992,
    n31993, n31994, n31995, n31996, n31997, n31998,
    n31999, n32000, n32001, n32002, n32003, n32004,
    n32005, n32006, n32007, n32008, n32009, n32010,
    n32011, n32012, n32013, n32014, n32015, n32016,
    n32017, n32018, n32019, n32020, n32021, n32022,
    n32023, n32024, n32025, n32026, n32027, n32028,
    n32029, n32030, n32031, n32032, n32033, n32034,
    n32035, n32036, n32037, n32038, n32039, n32040,
    n32041, n32042, n32043, n32044, n32045, n32046,
    n32047, n32048, n32049, n32050, n32051, n32052,
    n32053, n32054, n32055, n32056, n32057, n32058,
    n32059, n32060, n32061, n32062, n32063, n32064,
    n32065, n32066, n32067, n32068, n32069, n32070,
    n32071, n32072, n32073, n32074, n32075, n32076,
    n32077, n32078, n32079, n32080, n32081, n32082,
    n32083, n32084, n32085, n32086, n32087, n32088,
    n32089, n32090, n32091, n32092, n32093, n32094,
    n32095, n32096, n32097, n32098, n32099, n32100,
    n32101, n32102, n32103, n32104, n32105, n32106,
    n32107, n32108, n32109, n32110, n32111, n32112,
    n32113, n32114, n32115, n32116, n32117, n32118,
    n32119, n32120, n32121, n32122, n32123, n32124,
    n32125, n32126, n32127, n32128, n32129, n32130,
    n32131, n32132, n32133, n32134, n32135, n32136,
    n32137, n32138, n32139, n32140, n32141, n32142,
    n32143, n32144, n32145, n32146, n32147, n32148,
    n32149, n32150, n32151, n32152, n32153, n32154,
    n32155, n32156, n32157, n32158, n32159, n32160,
    n32161, n32162, n32163, n32164, n32165, n32166,
    n32167, n32168, n32169, n32170, n32171, n32172,
    n32173, n32174, n32175, n32176, n32177, n32178,
    n32179, n32180, n32181, n32182, n32183, n32184,
    n32185, n32186, n32187, n32188, n32189, n32190,
    n32191, n32192, n32193, n32194, n32195, n32196,
    n32197, n32198, n32199, n32200, n32201, n32202,
    n32203, n32204, n32205, n32206, n32207, n32208,
    n32209, n32210, n32211, n32212, n32213, n32214,
    n32215, n32216, n32217, n32218, n32219, n32220,
    n32221, n32222, n32223, n32224, n32225, n32226,
    n32227, n32228, n32229, n32230, n32231, n32232,
    n32233, n32234, n32235, n32236, n32237, n32238,
    n32239, n32240, n32241, n32242, n32243, n32244,
    n32245, n32246, n32247, n32248, n32249, n32250,
    n32251, n32252, n32253, n32254, n32255, n32256,
    n32257, n32258, n32259, n32260, n32261, n32262,
    n32263, n32264, n32265, n32266, n32267, n32268,
    n32269, n32270, n32271, n32272, n32273, n32274,
    n32275, n32276, n32277, n32278, n32279, n32280,
    n32281, n32282, n32283, n32284, n32285, n32286,
    n32287, n32288, n32289, n32290, n32291, n32292,
    n32293, n32294, n32295, n32296, n32297, n32298,
    n32299, n32300, n32301, n32302, n32303, n32304,
    n32305, n32306, n32307, n32308, n32309, n32311,
    n32312, n32313, n32314, n32315, n32316, n32317,
    n32318, n32319, n32320, n32321, n32322, n32323,
    n32324, n32325, n32326, n32327, n32328, n32329,
    n32330, n32331, n32332, n32333, n32334, n32335,
    n32336, n32337, n32338, n32339, n32340, n32341,
    n32342, n32343, n32344, n32345, n32346, n32347,
    n32348, n32349, n32350, n32351, n32352, n32353,
    n32354, n32355, n32356, n32357, n32358, n32359,
    n32360, n32361, n32362, n32363, n32364, n32365,
    n32366, n32367, n32368, n32369, n32370, n32371,
    n32372, n32373, n32374, n32375, n32376, n32377,
    n32378, n32379, n32380, n32381, n32382, n32383,
    n32384, n32385, n32386, n32387, n32388, n32389,
    n32390, n32391, n32392, n32393, n32394, n32395,
    n32396, n32397, n32398, n32399, n32400, n32401,
    n32402, n32403, n32404, n32405, n32406, n32407,
    n32408, n32409, n32410, n32411, n32412, n32413,
    n32414, n32415, n32416, n32417, n32418, n32419,
    n32420, n32421, n32422, n32423, n32424, n32425,
    n32426, n32427, n32428, n32429, n32430, n32431,
    n32432, n32433, n32434, n32435, n32436, n32437,
    n32438, n32439, n32440, n32441, n32442, n32443,
    n32444, n32445, n32446, n32447, n32448, n32449,
    n32450, n32451, n32452, n32453, n32454, n32455,
    n32456, n32457, n32458, n32459, n32460, n32461,
    n32462, n32463, n32464, n32465, n32466, n32467,
    n32468, n32469, n32470, n32471, n32472, n32473,
    n32474, n32475, n32476, n32477, n32478, n32479,
    n32480, n32481, n32482, n32483, n32484, n32485,
    n32486, n32487, n32488, n32489, n32490, n32491,
    n32492, n32493, n32494, n32495, n32496, n32497,
    n32498, n32499, n32500, n32501, n32502, n32503,
    n32504, n32505, n32506, n32507, n32508, n32509,
    n32510, n32511, n32512, n32513, n32514, n32515,
    n32516, n32517, n32518, n32519, n32520, n32521,
    n32522, n32523, n32524, n32525, n32526, n32527,
    n32528, n32529, n32530, n32531, n32532, n32533,
    n32534, n32535, n32536, n32537, n32538, n32539,
    n32540, n32541, n32542, n32543, n32544, n32545,
    n32546, n32547, n32548, n32549, n32550, n32551,
    n32552, n32553, n32554, n32555, n32556, n32557,
    n32558, n32559, n32560, n32561, n32562, n32563,
    n32564, n32565, n32566, n32567, n32568, n32569,
    n32570, n32571, n32572, n32573, n32574, n32575,
    n32576, n32577, n32578, n32579, n32580, n32581,
    n32583, n32584, n32585, n32586, n32587, n32588,
    n32589, n32590, n32591, n32592, n32593, n32594,
    n32595, n32596, n32597, n32598, n32599, n32600,
    n32601, n32602, n32603, n32604, n32605, n32606,
    n32607, n32608, n32609, n32610, n32611, n32612,
    n32613, n32614, n32615, n32616, n32617, n32618,
    n32619, n32620, n32621, n32622, n32623, n32624,
    n32625, n32626, n32627, n32628, n32629, n32630,
    n32631, n32632, n32633, n32634, n32635, n32636,
    n32637, n32638, n32639, n32640, n32641, n32642,
    n32643, n32644, n32645, n32646, n32647, n32648,
    n32649, n32650, n32651, n32652, n32653, n32654,
    n32655, n32656, n32657, n32658, n32659, n32660,
    n32661, n32662, n32663, n32664, n32665, n32666,
    n32667, n32668, n32669, n32670, n32671, n32672,
    n32673, n32674, n32675, n32676, n32677, n32678,
    n32679, n32680, n32681, n32682, n32683, n32684,
    n32685, n32686, n32687, n32688, n32689, n32690,
    n32691, n32692, n32693, n32694, n32695, n32696,
    n32697, n32698, n32699, n32700, n32701, n32702,
    n32703, n32704, n32705, n32706, n32707, n32708,
    n32709, n32710, n32711, n32712, n32713, n32714,
    n32715, n32716, n32717, n32718, n32719, n32720,
    n32721, n32722, n32723, n32724, n32725, n32726,
    n32727, n32728, n32729, n32730, n32731, n32732,
    n32733, n32734, n32735, n32736, n32737, n32738,
    n32739, n32740, n32741, n32742, n32743, n32744,
    n32745, n32746, n32747, n32748, n32749, n32750,
    n32751, n32752, n32753, n32754, n32755, n32756,
    n32757, n32758, n32759, n32760, n32761, n32762,
    n32763, n32764, n32765, n32766, n32767, n32768,
    n32769, n32770, n32771, n32772, n32773, n32774,
    n32775, n32776, n32777, n32778, n32779, n32780,
    n32781, n32782, n32783, n32784, n32785, n32786,
    n32787, n32788, n32789, n32790, n32791, n32792,
    n32793, n32794, n32795, n32796, n32797, n32798,
    n32799, n32800, n32801, n32802, n32803, n32804,
    n32805, n32806, n32807, n32808, n32809, n32810,
    n32811, n32812, n32813, n32814, n32815, n32816,
    n32817, n32818, n32819, n32820, n32821, n32822,
    n32823, n32824, n32825, n32826, n32827, n32828,
    n32829, n32830, n32831, n32832, n32833, n32834,
    n32835, n32836, n32837, n32838, n32839, n32840,
    n32841, n32842, n32843, n32844, n32845, n32846,
    n32847, n32848, n32850, n32851, n32852, n32853,
    n32854, n32855, n32856, n32857, n32858, n32859,
    n32860, n32861, n32862, n32863, n32864, n32865,
    n32866, n32867, n32868, n32869, n32870, n32871,
    n32872, n32873, n32874, n32875, n32876, n32877,
    n32878, n32879, n32880, n32881, n32882, n32883,
    n32884, n32885, n32886, n32887, n32888, n32889,
    n32890, n32891, n32892, n32893, n32894, n32895,
    n32896, n32897, n32898, n32899, n32900, n32901,
    n32902, n32903, n32904, n32905, n32906, n32907,
    n32908, n32909, n32910, n32911, n32912, n32913,
    n32914, n32915, n32916, n32917, n32918, n32919,
    n32920, n32921, n32922, n32923, n32924, n32925,
    n32926, n32927, n32928, n32929, n32930, n32931,
    n32932, n32933, n32934, n32935, n32936, n32937,
    n32938, n32939, n32940, n32941, n32942, n32943,
    n32944, n32945, n32946, n32947, n32948, n32949,
    n32950, n32951, n32952, n32953, n32954, n32955,
    n32956, n32957, n32958, n32959, n32960, n32961,
    n32962, n32963, n32964, n32965, n32966, n32967,
    n32968, n32969, n32970, n32971, n32972, n32973,
    n32974, n32975, n32976, n32977, n32978, n32979,
    n32980, n32981, n32982, n32983, n32984, n32985,
    n32986, n32987, n32988, n32989, n32990, n32991,
    n32992, n32993, n32994, n32995, n32996, n32997,
    n32998, n32999, n33000, n33001, n33002, n33003,
    n33004, n33005, n33006, n33007, n33008, n33009,
    n33010, n33011, n33012, n33013, n33014, n33015,
    n33016, n33017, n33018, n33019, n33020, n33021,
    n33022, n33023, n33024, n33025, n33026, n33027,
    n33028, n33029, n33030, n33031, n33032, n33033,
    n33034, n33035, n33037, n33038, n33039, n33040,
    n33041, n33042, n33043, n33045, n33046, n33047,
    n33048, n33049, n33050, n33051, n33053, n33054,
    n33055, n33056, n33057, n33058, n33059, n33060,
    n33061, n33062, n33063, n33064, n33065, n33066,
    n33067, n33068, n33069, n33070, n33071, n33072,
    n33073, n33074, n33075, n33076, n33077, n33078,
    n33079, n33080, n33081, n33082, n33083, n33084,
    n33085, n33086, n33087, n33088, n33089, n33090,
    n33091, n33092, n33093, n33094, n33095, n33096,
    n33097, n33098, n33099, n33100, n33101, n33102,
    n33103, n33104, n33105, n33106, n33107, n33108,
    n33109, n33110, n33111, n33112, n33113, n33114,
    n33115, n33116, n33117, n33118, n33119, n33120,
    n33121, n33122, n33123, n33124, n33125, n33126,
    n33127, n33128, n33129, n33130, n33131, n33132,
    n33133, n33134, n33135, n33136, n33137, n33138,
    n33139, n33140, n33141, n33142, n33143, n33144,
    n33145, n33146, n33147, n33148, n33149, n33150,
    n33151, n33152, n33153, n33154, n33155, n33157,
    n33158, n33159, n33160, n33161, n33162, n33164,
    n33165, n33166, n33167, n33168, n33169, n33170,
    n33172, n33173, n33174, n33175, n33176, n33177,
    n33178, n33179, n33180, n33181, n33182, n33183,
    n33184, n33185, n33186, n33187, n33188, n33189,
    n33190, n33191, n33192, n33193, n33194, n33195,
    n33196, n33197, n33198, n33199, n33200, n33201,
    n33202, n33203, n33204, n33205, n33206, n33207,
    n33208, n33209, n33210, n33211, n33212, n33213,
    n33214, n33215, n33216, n33217, n33218, n33219,
    n33220, n33221, n33222, n33223, n33224, n33225,
    n33226, n33227, n33228, n33229, n33230, n33231,
    n33232, n33233, n33234, n33235, n33236, n33237,
    n33238, n33239, n33240, n33241, n33242, n33243,
    n33244, n33245, n33246, n33247, n33248, n33249,
    n33250, n33251, n33252, n33253, n33254, n33255,
    n33256, n33257, n33258, n33259, n33260, n33261,
    n33262, n33263, n33264, n33265, n33266, n33267,
    n33268, n33269, n33270, n33271, n33272, n33273,
    n33274, n33275, n33276, n33277, n33278, n33279,
    n33280, n33281, n33282, n33283, n33284, n33285,
    n33286, n33287, n33288, n33289, n33290, n33291,
    n33292, n33293, n33294, n33295, n33296, n33297,
    n33298, n33299, n33300, n33301, n33302, n33303,
    n33304, n33305, n33306, n33307, n33308, n33309,
    n33310, n33311, n33312, n33313, n33314, n33315,
    n33316, n33317, n33318, n33319, n33320, n33321,
    n33322, n33323, n33324, n33325, n33326, n33327,
    n33328, n33329, n33330, n33331, n33332, n33333,
    n33334, n33335, n33336, n33337, n33338, n33339,
    n33340, n33341, n33342, n33343, n33344, n33345,
    n33346, n33347, n33348, n33349, n33350, n33351,
    n33352, n33353, n33354, n33355, n33356, n33357,
    n33358, n33359, n33360, n33361, n33362, n33363,
    n33364, n33365, n33366, n33367, n33368, n33369,
    n33370, n33371, n33372, n33373, n33374, n33375,
    n33376, n33377, n33378, n33379, n33380, n33381,
    n33382, n33383, n33384, n33385, n33386, n33387,
    n33388, n33389, n33390, n33391, n33392, n33393,
    n33394, n33395, n33396, n33397, n33398, n33399,
    n33400, n33401, n33402, n33403, n33404, n33405,
    n33406, n33407, n33408, n33409, n33410, n33411,
    n33412, n33413, n33414, n33415, n33416, n33417,
    n33418, n33419, n33420, n33421, n33422, n33423,
    n33424, n33425, n33426, n33427, n33428, n33429,
    n33430, n33431, n33432, n33433, n33434, n33435,
    n33436, n33437, n33438, n33439, n33440, n33441,
    n33442, n33443, n33444, n33445, n33446, n33447,
    n33448, n33449, n33450, n33451, n33452, n33453,
    n33454, n33455, n33456, n33457, n33458, n33459,
    n33460, n33461, n33462, n33463, n33464, n33465,
    n33466, n33467, n33468, n33469, n33470, n33471,
    n33472, n33473, n33474, n33475, n33476, n33477,
    n33478, n33479, n33480, n33481, n33482, n33483,
    n33484, n33485, n33486, n33487, n33488, n33489,
    n33490, n33491, n33492, n33493, n33494, n33495,
    n33496, n33497, n33498, n33499, n33500, n33501,
    n33502, n33503, n33504, n33505, n33506, n33507,
    n33508, n33509, n33510, n33511, n33512, n33513,
    n33514, n33515, n33516, n33517, n33518, n33519,
    n33520, n33521, n33522, n33523, n33524, n33525,
    n33526, n33527, n33528, n33529, n33530, n33531,
    n33532, n33533, n33534, n33535, n33536, n33537,
    n33538, n33539, n33540, n33541, n33542, n33543,
    n33544, n33545, n33546, n33547, n33548, n33549,
    n33550, n33551, n33552, n33553, n33554, n33555,
    n33556, n33557, n33558, n33559, n33560, n33561,
    n33562, n33563, n33564, n33565, n33566, n33567,
    n33568, n33569, n33570, n33571, n33572, n33573,
    n33574, n33575, n33576, n33577, n33578, n33579,
    n33580, n33581, n33582, n33583, n33584, n33585,
    n33586, n33587, n33588, n33589, n33590, n33591,
    n33592, n33593, n33594, n33595, n33596, n33597,
    n33598, n33599, n33600, n33601, n33602, n33603,
    n33604, n33605, n33606, n33607, n33608, n33609,
    n33610, n33611, n33612, n33613, n33614, n33615,
    n33616, n33617, n33618, n33619, n33620, n33621,
    n33622, n33623, n33624, n33625, n33626, n33627,
    n33628, n33629, n33630, n33631, n33632, n33633,
    n33634, n33635, n33636, n33637, n33638, n33639,
    n33641, n33642, n33643, n33644, n33645, n33646,
    n33647, n33648, n33649, n33650, n33651, n33652,
    n33653, n33654, n33655, n33656, n33657, n33658,
    n33659, n33660, n33661, n33662, n33663, n33664,
    n33665, n33666, n33667, n33668, n33669, n33670,
    n33671, n33672, n33673, n33674, n33675, n33676,
    n33677, n33678, n33679, n33680, n33681, n33682,
    n33683, n33684, n33685, n33686, n33687, n33688,
    n33689, n33690, n33691, n33692, n33693, n33694,
    n33695, n33696, n33697, n33698, n33699, n33700,
    n33701, n33702, n33703, n33704, n33705, n33706,
    n33707, n33708, n33709, n33710, n33711, n33712,
    n33713, n33714, n33716, n33717, n33718, n33719,
    n33720, n33721, n33722, n33723, n33724, n33725,
    n33726, n33727, n33728, n33729, n33730, n33731,
    n33732, n33733, n33734, n33735, n33736, n33737,
    n33738, n33739, n33740, n33741, n33742, n33743,
    n33744, n33745, n33746, n33747, n33748, n33749,
    n33750, n33751, n33752, n33753, n33754, n33755,
    n33756, n33757, n33758, n33759, n33760, n33761,
    n33762, n33763, n33764, n33765, n33766, n33767,
    n33768, n33769, n33770, n33771, n33772, n33773,
    n33774, n33775, n33776, n33777, n33778, n33779,
    n33780, n33781, n33782, n33783, n33784, n33785,
    n33786, n33787, n33788, n33789, n33790, n33791,
    n33792, n33793, n33794, n33795, n33796, n33797,
    n33798, n33799, n33800, n33801, n33802, n33803,
    n33804, n33805, n33806, n33807, n33808, n33809,
    n33810, n33811, n33812, n33813, n33814, n33815,
    n33816, n33817, n33818, n33819, n33820, n33821,
    n33822, n33823, n33824, n33825, n33826, n33827,
    n33828, n33829, n33830, n33831, n33832, n33833,
    n33834, n33835, n33836, n33837, n33838, n33839,
    n33840, n33841, n33842, n33843, n33844, n33845,
    n33846, n33847, n33848, n33849, n33850, n33851,
    n33852, n33853, n33854, n33855, n33856, n33857,
    n33858, n33859, n33860, n33862, n33863, n33864,
    n33865, n33866, n33867, n33868, n33869, n33870,
    n33871, n33872, n33873, n33874, n33875, n33876,
    n33877, n33878, n33879, n33880, n33881, n33882,
    n33883, n33884, n33885, n33886, n33887, n33888,
    n33889, n33890, n33891, n33892, n33893, n33894,
    n33895, n33896, n33897, n33898, n33899, n33900,
    n33901, n33902, n33903, n33904, n33905, n33906,
    n33907, n33908, n33909, n33910, n33911, n33912,
    n33913, n33914, n33915, n33916, n33917, n33918,
    n33919, n33920, n33921, n33922, n33923, n33924,
    n33925, n33926, n33927, n33928, n33929, n33930,
    n33931, n33932, n33933, n33934, n33935, n33936,
    n33937, n33938, n33939, n33940, n33941, n33942,
    n33943, n33944, n33945, n33946, n33947, n33948,
    n33949, n33950, n33951, n33952, n33953, n33954,
    n33955, n33956, n33957, n33958, n33959, n33960,
    n33961, n33962, n33963, n33964, n33965, n33966,
    n33967, n33968, n33969, n33970, n33971, n33972,
    n33973, n33974, n33975, n33976, n33977, n33978,
    n33979, n33980, n33981, n33982, n33983, n33984,
    n33985, n33986, n33988, n33989, n33990, n33991,
    n33992, n33993, n33994, n33995, n33996, n33997,
    n33998, n33999, n34000, n34001, n34002, n34003,
    n34004, n34005, n34006, n34007, n34008, n34009,
    n34010, n34011, n34012, n34013, n34015, n34016,
    n34017, n34018, n34019, n34020, n34021, n34022,
    n34023, n34024, n34025, n34026, n34027, n34028,
    n34029, n34030, n34031, n34032, n34033, n34034,
    n34036, n34037, n34038, n34039, n34040, n34041,
    n34042, n34043, n34044, n34045, n34046, n34047,
    n34048, n34049, n34050, n34051, n34052, n34053,
    n34054, n34055, n34057, n34058, n34059, n34060,
    n34061, n34062, n34063, n34064, n34065, n34066,
    n34067, n34068, n34069, n34070, n34071, n34072,
    n34073, n34074, n34075, n34076, n34078, n34079,
    n34080, n34081, n34082, n34083, n34084, n34085,
    n34086, n34087, n34088, n34089, n34090, n34091,
    n34092, n34093, n34094, n34095, n34096, n34097,
    n34098, n34099, n34100, n34101, n34102, n34103,
    n34104, n34105, n34106, n34107, n34108, n34109,
    n34110, n34111, n34112, n34113, n34114, n34115,
    n34116, n34117, n34118, n34119, n34120, n34121,
    n34122, n34123, n34124, n34125, n34126, n34127,
    n34128, n34129, n34130, n34131, n34132, n34133,
    n34134, n34135, n34136, n34137, n34138, n34139,
    n34140, n34141, n34142, n34143, n34144, n34145,
    n34146, n34147, n34148, n34149, n34150, n34151,
    n34152, n34153, n34154, n34155, n34156, n34157,
    n34158, n34159, n34160, n34161, n34162, n34163,
    n34164, n34165, n34166, n34167, n34168, n34169,
    n34170, n34171, n34172, n34173, n34174, n34175,
    n34176, n34177, n34178, n34179, n34180, n34181,
    n34182, n34183, n34184, n34185, n34186, n34187,
    n34188, n34190, n34191, n34192, n34193, n34194,
    n34195, n34196, n34197, n34198, n34199, n34200,
    n34201, n34202, n34203, n34204, n34205, n34206,
    n34207, n34208, n34209, n34210, n34211, n34212,
    n34213, n34214, n34215, n34216, n34217, n34218,
    n34219, n34220, n34221, n34222, n34223, n34224,
    n34225, n34226, n34227, n34228, n34229, n34230,
    n34231, n34232, n34233, n34234, n34235, n34236,
    n34237, n34238, n34239, n34240, n34241, n34242,
    n34243, n34244, n34245, n34246, n34247, n34248,
    n34249, n34250, n34251, n34252, n34253, n34254,
    n34255, n34256, n34257, n34258, n34259, n34260,
    n34261, n34262, n34263, n34264, n34265, n34266,
    n34267, n34268, n34269, n34270, n34271, n34272,
    n34273, n34274, n34275, n34276, n34277, n34278,
    n34279, n34280, n34281, n34282, n34283, n34284,
    n34285, n34286, n34287, n34289, n34290, n34291,
    n34292, n34293, n34294, n34295, n34296, n34297,
    n34298, n34299, n34300, n34301, n34302, n34303,
    n34304, n34305, n34306, n34308, n34309, n34310,
    n34311, n34312, n34313, n34315, n34316, n34317,
    n34318, n34319, n34320, n34321, n34322, n34323,
    n34324, n34325, n34326, n34327, n34328, n34329,
    n34330, n34331, n34332, n34333, n34334, n34336,
    n34337, n34338, n34339, n34340, n34341, n34343,
    n34344, n34345, n34346, n34347, n34348, n34349,
    n34350, n34351, n34352, n34353, n34354, n34355,
    n34356, n34357, n34358, n34359, n34360, n34361,
    n34362, n34363, n34364, n34365, n34366, n34367,
    n34368, n34369, n34370, n34371, n34372, n34373,
    n34374, n34375, n34376, n34377, n34378, n34379,
    n34380, n34381, n34382, n34383, n34384, n34385,
    n34386, n34387, n34388, n34389, n34390, n34391,
    n34392, n34393, n34394, n34395, n34396, n34397,
    n34398, n34399, n34400, n34401, n34402, n34403,
    n34404, n34405, n34406, n34407, n34408, n34409,
    n34410, n34411, n34412, n34413, n34414, n34415,
    n34416, n34417, n34418, n34419, n34420, n34421,
    n34422, n34423, n34424, n34425, n34426, n34427,
    n34428, n34429, n34430, n34431, n34432, n34433,
    n34434, n34435, n34436, n34437, n34438, n34439,
    n34440, n34441, n34442, n34443, n34444, n34445,
    n34446, n34448, n34449, n34450, n34451, n34452,
    n34453, n34454, n34455, n34456, n34457, n34458,
    n34459, n34460, n34461, n34462, n34463, n34464,
    n34465, n34466, n34467, n34468, n34469, n34470,
    n34471, n34472, n34473, n34474, n34475, n34476,
    n34477, n34478, n34479, n34480, n34481, n34482,
    n34483, n34484, n34485, n34486, n34487, n34488,
    n34489, n34490, n34491, n34492, n34493, n34494,
    n34495, n34496, n34497, n34498, n34499, n34500,
    n34501, n34502, n34503, n34504, n34505, n34506,
    n34507, n34508, n34509, n34510, n34511, n34512,
    n34513, n34514, n34515, n34516, n34517, n34518,
    n34519, n34520, n34521, n34522, n34523, n34524,
    n34525, n34526, n34527, n34528, n34529, n34530,
    n34531, n34532, n34533, n34534, n34535, n34536,
    n34537, n34538, n34539, n34540, n34541, n34542,
    n34543, n34544, n34545, n34546, n34547, n34548,
    n34549, n34550, n34551, n34552, n34553, n34554,
    n34555, n34556, n34557, n34558, n34559, n34560,
    n34561, n34562, n34563, n34564, n34565, n34566,
    n34567, n34568, n34569, n34570, n34571, n34572,
    n34573, n34574, n34575, n34576, n34577, n34578,
    n34579, n34580, n34581, n34582, n34583, n34584,
    n34585, n34586, n34587, n34588, n34589, n34590,
    n34591, n34592, n34593, n34594, n34595, n34596,
    n34597, n34598, n34599, n34600, n34601, n34602,
    n34603, n34604, n34605, n34606, n34607, n34608,
    n34609, n34610, n34611, n34612, n34613, n34614,
    n34615, n34616, n34617, n34618, n34619, n34620,
    n34621, n34622, n34623, n34624, n34625, n34626,
    n34627, n34628, n34629, n34630, n34631, n34632,
    n34633, n34634, n34635, n34636, n34637, n34638,
    n34639, n34640, n34641, n34642, n34643, n34644,
    n34645, n34646, n34647, n34648, n34649, n34650,
    n34651, n34652, n34653, n34654, n34655, n34656,
    n34657, n34658, n34659, n34660, n34661, n34662,
    n34663, n34664, n34665, n34666, n34667, n34668,
    n34669, n34670, n34671, n34672, n34673, n34674,
    n34675, n34676, n34677, n34678, n34679, n34680,
    n34681, n34682, n34683, n34684, n34685, n34686,
    n34687, n34688, n34689, n34690, n34691, n34692,
    n34693, n34694, n34695, n34696, n34697, n34698,
    n34699, n34700, n34701, n34702, n34703, n34704,
    n34705, n34706, n34707, n34708, n34709, n34710,
    n34711, n34712, n34713, n34714, n34715, n34716,
    n34717, n34718, n34719, n34720, n34721, n34722,
    n34723, n34724, n34725, n34726, n34727, n34728,
    n34729, n34730, n34731, n34732, n34733, n34734,
    n34735, n34736, n34737, n34738, n34739, n34740,
    n34741, n34742, n34743, n34744, n34745, n34746,
    n34747, n34748, n34749, n34750, n34751, n34752,
    n34753, n34754, n34755, n34756, n34757, n34758,
    n34759, n34760, n34761, n34762, n34763, n34764,
    n34765, n34766, n34767, n34768, n34769, n34770,
    n34771, n34772, n34773, n34774, n34775, n34776,
    n34777, n34778, n34779, n34780, n34781, n34782,
    n34783, n34784, n34785, n34786, n34787, n34788,
    n34789, n34790, n34791, n34792, n34793, n34794,
    n34795, n34796, n34797, n34798, n34799, n34800,
    n34801, n34802, n34803, n34804, n34805, n34806,
    n34807, n34808, n34809, n34810, n34811, n34812,
    n34813, n34814, n34815, n34816, n34817, n34818,
    n34819, n34820, n34821, n34822, n34823, n34824,
    n34825, n34826, n34827, n34828, n34829, n34830,
    n34831, n34832, n34833, n34834, n34835, n34836,
    n34837, n34838, n34839, n34840, n34841, n34842,
    n34843, n34844, n34845, n34846, n34847, n34848,
    n34849, n34850, n34851, n34852, n34853, n34854,
    n34855, n34856, n34857, n34858, n34859, n34860,
    n34861, n34862, n34863, n34864, n34865, n34866,
    n34867, n34868, n34869, n34870, n34871, n34872,
    n34873, n34874, n34875, n34876, n34877, n34878,
    n34879, n34880, n34881, n34882, n34883, n34884,
    n34885, n34886, n34887, n34888, n34889, n34890,
    n34891, n34892, n34893, n34894, n34895, n34896,
    n34897, n34898, n34899, n34900, n34901, n34902,
    n34903, n34904, n34905, n34906, n34907, n34908,
    n34909, n34910, n34911, n34912, n34913, n34914,
    n34915, n34916, n34917, n34918, n34919, n34920,
    n34921, n34922, n34923, n34924, n34925, n34926,
    n34927, n34928, n34929, n34930, n34931, n34932,
    n34933, n34934, n34935, n34936, n34937, n34938,
    n34939, n34940, n34941, n34942, n34943, n34944,
    n34945, n34946, n34947, n34948, n34949, n34950,
    n34951, n34952, n34953, n34954, n34955, n34956,
    n34957, n34958, n34959, n34960, n34961, n34962,
    n34963, n34964, n34965, n34966, n34967, n34968,
    n34969, n34970, n34971, n34972, n34973, n34974,
    n34975, n34976, n34977, n34978, n34979, n34980,
    n34981, n34982, n34983, n34984, n34985, n34986,
    n34987, n34988, n34989, n34990, n34991, n34992,
    n34993, n34994, n34995, n34996, n34997, n34998,
    n34999, n35000, n35001, n35002, n35003, n35004,
    n35005, n35006, n35007, n35008, n35009, n35010,
    n35011, n35012, n35013, n35014, n35015, n35016,
    n35017, n35018, n35019, n35020, n35021, n35022,
    n35023, n35024, n35025, n35026, n35027, n35028,
    n35029, n35030, n35031, n35032, n35033, n35034,
    n35035, n35036, n35037, n35038, n35039, n35040,
    n35041, n35042, n35043, n35044, n35045, n35046,
    n35047, n35048, n35050, n35051, n35052, n35053,
    n35054, n35055, n35056, n35057, n35058, n35059,
    n35060, n35061, n35062, n35063, n35064, n35065,
    n35066, n35067, n35068, n35069, n35070, n35071,
    n35072, n35073, n35074, n35075, n35076, n35077,
    n35078, n35079, n35080, n35081, n35082, n35083,
    n35084, n35085, n35086, n35087, n35088, n35089,
    n35090, n35091, n35092, n35093, n35094, n35095,
    n35096, n35097, n35098, n35099, n35100, n35101,
    n35102, n35103, n35104, n35105, n35106, n35107,
    n35108, n35109, n35110, n35111, n35112, n35113,
    n35114, n35115, n35116, n35117, n35118, n35119,
    n35120, n35121, n35122, n35123, n35124, n35125,
    n35126, n35127, n35128, n35129, n35130, n35131,
    n35132, n35133, n35134, n35135, n35136, n35137,
    n35138, n35139, n35140, n35141, n35142, n35143,
    n35144, n35145, n35146, n35147, n35148, n35149,
    n35150, n35151, n35152, n35153, n35154, n35155,
    n35156, n35157, n35158, n35159, n35160, n35161,
    n35162, n35163, n35164, n35165, n35166, n35167,
    n35168, n35169, n35170, n35171, n35172, n35173,
    n35174, n35175, n35176, n35177, n35178, n35179,
    n35180, n35181, n35182, n35183, n35184, n35185,
    n35186, n35187, n35188, n35189, n35190, n35191,
    n35192, n35193, n35194, n35195, n35196, n35197,
    n35198, n35199, n35200, n35201, n35202, n35203,
    n35204, n35205, n35206, n35207, n35208, n35209,
    n35210, n35211, n35212, n35213, n35214, n35215,
    n35216, n35217, n35218, n35219, n35220, n35221,
    n35222, n35223, n35224, n35225, n35226, n35227,
    n35228, n35229, n35230, n35231, n35232, n35233,
    n35234, n35235, n35236, n35237, n35238, n35239,
    n35240, n35241, n35242, n35243, n35244, n35245,
    n35246, n35247, n35248, n35249, n35250, n35251,
    n35252, n35253, n35254, n35255, n35256, n35257,
    n35258, n35259, n35260, n35261, n35262, n35263,
    n35264, n35265, n35266, n35267, n35268, n35269,
    n35270, n35271, n35272, n35273, n35274, n35275,
    n35276, n35277, n35278, n35279, n35280, n35281,
    n35282, n35283, n35284, n35285, n35286, n35287,
    n35288, n35289, n35290, n35291, n35292, n35293,
    n35294, n35295, n35296, n35297, n35298, n35299,
    n35300, n35301, n35302, n35303, n35304, n35305,
    n35306, n35307, n35308, n35309, n35310, n35311,
    n35312, n35313, n35314, n35315, n35316, n35317,
    n35318, n35319, n35320, n35321, n35322, n35323,
    n35324, n35325, n35326, n35327, n35328, n35329,
    n35330, n35331, n35332, n35333, n35334, n35335,
    n35336, n35337, n35338, n35339, n35340, n35341,
    n35342, n35343, n35344, n35345, n35346, n35347,
    n35348, n35349, n35350, n35351, n35352, n35353,
    n35354, n35355, n35356, n35357, n35358, n35359,
    n35360, n35361, n35362, n35363, n35364, n35365,
    n35366, n35367, n35368, n35369, n35370, n35371,
    n35372, n35373, n35374, n35375, n35376, n35377,
    n35378, n35379, n35380, n35381, n35382, n35383,
    n35384, n35385, n35386, n35387, n35388, n35389,
    n35390, n35391, n35392, n35393, n35394, n35395,
    n35396, n35397, n35398, n35399, n35400, n35401,
    n35402, n35403, n35404, n35405, n35406, n35407,
    n35408, n35409, n35410, n35411, n35412, n35413,
    n35414, n35415, n35416, n35417, n35418, n35419,
    n35420, n35421, n35422, n35423, n35424, n35425,
    n35426, n35427, n35428, n35429, n35430, n35431,
    n35432, n35433, n35434, n35435, n35436, n35437,
    n35438, n35439, n35440, n35441, n35442, n35443,
    n35444, n35445, n35446, n35447, n35448, n35449,
    n35450, n35451, n35452, n35453, n35454, n35455,
    n35456, n35457, n35458, n35459, n35460, n35461,
    n35462, n35463, n35464, n35465, n35466, n35467,
    n35468, n35469, n35470, n35471, n35472, n35473,
    n35474, n35475, n35476, n35477, n35478, n35479,
    n35480, n35481, n35482, n35483, n35484, n35485,
    n35486, n35487, n35488, n35489, n35490, n35491,
    n35492, n35493, n35494, n35495, n35496, n35497,
    n35498, n35499, n35500, n35501, n35502, n35503,
    n35504, n35505, n35506, n35507, n35508, n35509,
    n35510, n35511, n35512, n35513, n35514, n35515,
    n35516, n35517, n35518, n35519, n35520, n35521,
    n35522, n35523, n35524, n35525, n35526, n35527,
    n35528, n35529, n35530, n35531, n35532, n35533,
    n35534, n35535, n35536, n35537, n35538, n35539,
    n35540, n35541, n35542, n35543, n35544, n35545,
    n35546, n35547, n35548, n35549, n35550, n35551,
    n35552, n35553, n35554, n35555, n35556, n35557,
    n35558, n35559, n35560, n35561, n35562, n35563,
    n35564, n35565, n35566, n35567, n35568, n35569,
    n35570, n35571, n35572, n35573, n35574, n35575,
    n35576, n35577, n35578, n35579, n35580, n35581,
    n35582, n35583, n35584, n35585, n35586, n35587,
    n35588, n35589, n35590, n35591, n35592, n35593,
    n35594, n35595, n35596, n35597, n35598, n35599,
    n35600, n35601, n35602, n35603, n35604, n35605,
    n35606, n35607, n35608, n35610, n35611, n35612,
    n35613, n35614, n35615, n35616, n35617, n35618,
    n35619, n35620, n35621, n35622, n35623, n35624,
    n35625, n35626, n35627, n35628, n35629, n35630,
    n35631, n35632, n35633, n35634, n35635, n35636,
    n35637, n35638, n35639, n35640, n35641, n35642,
    n35643, n35644, n35645, n35646, n35647, n35648,
    n35649, n35650, n35651, n35652, n35653, n35654,
    n35655, n35656, n35657, n35658, n35659, n35660,
    n35661, n35662, n35663, n35664, n35665, n35666,
    n35667, n35668, n35669, n35670, n35671, n35672,
    n35673, n35674, n35675, n35676, n35677, n35678,
    n35679, n35680, n35681, n35682, n35683, n35684,
    n35685, n35686, n35687, n35688, n35689, n35690,
    n35691, n35692, n35693, n35694, n35695, n35696,
    n35697, n35698, n35699, n35700, n35701, n35702,
    n35703, n35704, n35705, n35706, n35707, n35708,
    n35709, n35710, n35711, n35712, n35713, n35714,
    n35715, n35716, n35717, n35718, n35719, n35720,
    n35721, n35722, n35723, n35724, n35725, n35726,
    n35727, n35728, n35729, n35730, n35731, n35732,
    n35733, n35734, n35735, n35736, n35737, n35738,
    n35739, n35740, n35741, n35742, n35743, n35744,
    n35745, n35746, n35747, n35748, n35749, n35750,
    n35751, n35752, n35753, n35754, n35755, n35756,
    n35757, n35758, n35759, n35760, n35761, n35762,
    n35763, n35764, n35765, n35766, n35767, n35768,
    n35769, n35770, n35771, n35772, n35773, n35774,
    n35775, n35776, n35777, n35778, n35779, n35780,
    n35781, n35782, n35783, n35784, n35785, n35786,
    n35787, n35788, n35789, n35790, n35791, n35792,
    n35793, n35794, n35795, n35796, n35797, n35798,
    n35799, n35800, n35801, n35802, n35803, n35804,
    n35805, n35806, n35807, n35808, n35809, n35810,
    n35811, n35812, n35813, n35814, n35815, n35816,
    n35817, n35818, n35819, n35820, n35821, n35822,
    n35823, n35824, n35825, n35826, n35827, n35828,
    n35829, n35830, n35831, n35832, n35833, n35834,
    n35835, n35836, n35837, n35838, n35839, n35840,
    n35841, n35842, n35843, n35844, n35845, n35846,
    n35847, n35848, n35849, n35850, n35851, n35852,
    n35853, n35854, n35855, n35856, n35857, n35858,
    n35859, n35860, n35861, n35862, n35863, n35864,
    n35865, n35866, n35867, n35868, n35869, n35870,
    n35871, n35872, n35873, n35874, n35875, n35876,
    n35877, n35878, n35879, n35880, n35881, n35882,
    n35883, n35884, n35885, n35886, n35887, n35888,
    n35889, n35890, n35891, n35892, n35893, n35894,
    n35895, n35896, n35897, n35898, n35899, n35900,
    n35901, n35902, n35903, n35904, n35905, n35906,
    n35907, n35908, n35909, n35910, n35911, n35912,
    n35913, n35914, n35915, n35916, n35917, n35918,
    n35919, n35920, n35921, n35922, n35923, n35924,
    n35925, n35926, n35927, n35928, n35929, n35930,
    n35931, n35932, n35933, n35934, n35935, n35936,
    n35937, n35938, n35939, n35940, n35941, n35942,
    n35943, n35944, n35945, n35946, n35947, n35948,
    n35949, n35950, n35951, n35952, n35953, n35954,
    n35955, n35956, n35957, n35958, n35959, n35960,
    n35961, n35962, n35963, n35964, n35965, n35966,
    n35967, n35968, n35969, n35970, n35971, n35972,
    n35973, n35974, n35975, n35976, n35977, n35978,
    n35979, n35980, n35981, n35982, n35983, n35984,
    n35985, n35986, n35987, n35988, n35989, n35990,
    n35991, n35992, n35993, n35994, n35995, n35996,
    n35997, n35998, n35999, n36000, n36001, n36002,
    n36003, n36004, n36005, n36006, n36007, n36008,
    n36009, n36010, n36011, n36012, n36013, n36014,
    n36015, n36016, n36017, n36018, n36019, n36020,
    n36021, n36022, n36023, n36024, n36025, n36026,
    n36027, n36028, n36029, n36030, n36031, n36032,
    n36033, n36034, n36035, n36036, n36037, n36038,
    n36039, n36040, n36041, n36042, n36043, n36044,
    n36045, n36046, n36047, n36048, n36049, n36050,
    n36051, n36052, n36053, n36054, n36055, n36056,
    n36057, n36058, n36059, n36060, n36061, n36062,
    n36063, n36064, n36065, n36066, n36067, n36068,
    n36069, n36070, n36071, n36072, n36073, n36074,
    n36075, n36076, n36077, n36078, n36079, n36080,
    n36081, n36082, n36083, n36084, n36085, n36086,
    n36087, n36088, n36089, n36090, n36091, n36092,
    n36093, n36094, n36095, n36096, n36097, n36098,
    n36099, n36100, n36101, n36102, n36103, n36104,
    n36105, n36106, n36107, n36108, n36109, n36110,
    n36111, n36112, n36113, n36114, n36115, n36116,
    n36117, n36118, n36119, n36120, n36121, n36122,
    n36123, n36124, n36125, n36126, n36127, n36128,
    n36129, n36130, n36131, n36132, n36133, n36134,
    n36135, n36136, n36137, n36138, n36139, n36140,
    n36141, n36142, n36143, n36144, n36145, n36146,
    n36147, n36148, n36150, n36151, n36152, n36153,
    n36154, n36155, n36156, n36157, n36158, n36159,
    n36160, n36161, n36162, n36163, n36164, n36165,
    n36166, n36167, n36168, n36169, n36170, n36171,
    n36172, n36173, n36174, n36175, n36176, n36177,
    n36178, n36179, n36180, n36181, n36182, n36183,
    n36184, n36185, n36186, n36187, n36188, n36189,
    n36190, n36191, n36192, n36193, n36194, n36195,
    n36196, n36197, n36198, n36199, n36200, n36201,
    n36202, n36203, n36204, n36205, n36206, n36207,
    n36208, n36209, n36210, n36211, n36212, n36213,
    n36214, n36215, n36216, n36217, n36218, n36219,
    n36220, n36221, n36222, n36223, n36224, n36225,
    n36226, n36227, n36228, n36229, n36230, n36231,
    n36232, n36233, n36234, n36235, n36236, n36237,
    n36238, n36239, n36240, n36241, n36242, n36243,
    n36244, n36245, n36246, n36247, n36248, n36249,
    n36250, n36251, n36252, n36253, n36254, n36255,
    n36256, n36257, n36258, n36259, n36260, n36261,
    n36262, n36263, n36264, n36265, n36266, n36267,
    n36268, n36269, n36270, n36271, n36272, n36274,
    n36275, n36276, n36277, n36278, n36279, n36280,
    n36281, n36282, n36283, n36284, n36285, n36286,
    n36287, n36288, n36289, n36290, n36291, n36292,
    n36293, n36294, n36295, n36296, n36297, n36298,
    n36299, n36300, n36301, n36302, n36303, n36304,
    n36305, n36306, n36307, n36308, n36309, n36310,
    n36311, n36312, n36313, n36314, n36315, n36316,
    n36317, n36318, n36319, n36320, n36321, n36322,
    n36323, n36324, n36325, n36326, n36328, n36329,
    n36330, n36331, n36332, n36333, n36334, n36335,
    n36336, n36337, n36338, n36339, n36340, n36341,
    n36342, n36343, n36344, n36345, n36346, n36347,
    n36348, n36349, n36350, n36351, n36352, n36353,
    n36354, n36355, n36356, n36358, n36359, n36360,
    n36361, n36362, n36363, n36364, n36365, n36367,
    n36368, n36369, n36370, n36371, n36372, n36373,
    n36374, n36375, n36376, n36377, n36378, n36379,
    n36380, n36381, n36382, n36383, n36384, n36385,
    n36386, n36387, n36388, n36389, n36390, n36391,
    n36392, n36393, n36394, n36395, n36396, n36397,
    n36398, n36399, n36400, n36401, n36402, n36403,
    n36404, n36405, n36406, n36407, n36408, n36409,
    n36410, n36411, n36412, n36413, n36414, n36415,
    n36416, n36417, n36418, n36419, n36420, n36421,
    n36422, n36423, n36424, n36425, n36426, n36427,
    n36428, n36429, n36430, n36431, n36432, n36433,
    n36434, n36435, n36436, n36437, n36438, n36439,
    n36440, n36441, n36442, n36444, n36445, n36446,
    n36447, n36448, n36449, n36450, n36451, n36452,
    n36453, n36454, n36455, n36456, n36457, n36458,
    n36459, n36460, n36461, n36462, n36463, n36464,
    n36465, n36466, n36467, n36468, n36469, n36470,
    n36471, n36472, n36473, n36474, n36475, n36476,
    n36477, n36478, n36480, n36481, n36482, n36483,
    n36484, n36485, n36486, n36487, n36488, n36489,
    n36490, n36491, n36492, n36493, n36494, n36495,
    n36496, n36497, n36498, n36499, n36500, n36501,
    n36502, n36504, n36505, n36506, n36507, n36508,
    n36509, n36510, n36511, n36512, n36513, n36514,
    n36515, n36516, n36517, n36518, n36519, n36520,
    n36521, n36522, n36523, n36524, n36525, n36526,
    n36527, n36528, n36529, n36530, n36531, n36532,
    n36533, n36534, n36535, n36536, n36537, n36538,
    n36539, n36540, n36541, n36542, n36543, n36544,
    n36545, n36546, n36547, n36548, n36549, n36550,
    n36551, n36552, n36553, n36554, n36555, n36556,
    n36557, n36558, n36559, n36560, n36561, n36562,
    n36563, n36564, n36565, n36566, n36567, n36568,
    n36569, n36570, n36571, n36572, n36573, n36574,
    n36575, n36576, n36577, n36578, n36579, n36580,
    n36581, n36582, n36583, n36584, n36585, n36586,
    n36587, n36588, n36589, n36590, n36591, n36592,
    n36593, n36594, n36595, n36596, n36597, n36598,
    n36599, n36600, n36601, n36602, n36603, n36604,
    n36605, n36606, n36607, n36608, n36609, n36610,
    n36611, n36612, n36613, n36614, n36615, n36616,
    n36617, n36618, n36619, n36620, n36621, n36622,
    n36623, n36624, n36625, n36626, n36627, n36628,
    n36629, n36630, n36631, n36632, n36633, n36634,
    n36635, n36636, n36637, n36638, n36639, n36640,
    n36641, n36642, n36643, n36644, n36645, n36646,
    n36647, n36648, n36649, n36650, n36651, n36652,
    n36653, n36654, n36655, n36656, n36657, n36658,
    n36659, n36660, n36661, n36662, n36663, n36664,
    n36665, n36666, n36667, n36668, n36669, n36670,
    n36671, n36672, n36673, n36674, n36675, n36676,
    n36677, n36678, n36679, n36680, n36681, n36682,
    n36683, n36684, n36685, n36686, n36687, n36688,
    n36689, n36690, n36691, n36692, n36693, n36694,
    n36695, n36696, n36697, n36698, n36699, n36700,
    n36701, n36702, n36703, n36704, n36705, n36706,
    n36707, n36708, n36709, n36710, n36711, n36712,
    n36713, n36714, n36715, n36716, n36717, n36718,
    n36719, n36720, n36721, n36722, n36723, n36724,
    n36725, n36726, n36727, n36728, n36729, n36730,
    n36731, n36732, n36733, n36734, n36735, n36736,
    n36737, n36738, n36739, n36740, n36741, n36742,
    n36743, n36744, n36745, n36746, n36747, n36748,
    n36749, n36750, n36751, n36752, n36753, n36754,
    n36755, n36756, n36757, n36758, n36759, n36760,
    n36761, n36762, n36763, n36764, n36765, n36766,
    n36767, n36768, n36769, n36770, n36771, n36772,
    n36773, n36774, n36775, n36776, n36777, n36778,
    n36779, n36780, n36781, n36782, n36783, n36784,
    n36785, n36786, n36787, n36788, n36789, n36790,
    n36791, n36792, n36793, n36794, n36795, n36796,
    n36797, n36798, n36799, n36800, n36801, n36802,
    n36803, n36804, n36805, n36806, n36807, n36808,
    n36809, n36810, n36811, n36812, n36813, n36814,
    n36815, n36816, n36817, n36818, n36819, n36820,
    n36821, n36822, n36823, n36824, n36825, n36826,
    n36827, n36828, n36829, n36830, n36831, n36832,
    n36833, n36834, n36835, n36836, n36837, n36838,
    n36839, n36840, n36841, n36842, n36843, n36844,
    n36845, n36846, n36847, n36848, n36849, n36850,
    n36851, n36852, n36853, n36854, n36855, n36856,
    n36857, n36858, n36859, n36860, n36861, n36862,
    n36863, n36864, n36865, n36866, n36867, n36868,
    n36870, n36871, n36872, n36873, n36874, n36875,
    n36876, n36877, n36878, n36879, n36880, n36881,
    n36882, n36883, n36884, n36885, n36886, n36887,
    n36888, n36889, n36890, n36891, n36892, n36893,
    n36894, n36895, n36896, n36897, n36898, n36899,
    n36900, n36901, n36902, n36903, n36904, n36905,
    n36906, n36907, n36908, n36909, n36910, n36911,
    n36912, n36913, n36914, n36915, n36916, n36917,
    n36918, n36919, n36920, n36921, n36922, n36923,
    n36924, n36925, n36926, n36927, n36928, n36929,
    n36930, n36931, n36932, n36933, n36934, n36935,
    n36936, n36937, n36938, n36939, n36940, n36941,
    n36942, n36943, n36944, n36945, n36946, n36947,
    n36948, n36949, n36950, n36951, n36952, n36953,
    n36954, n36955, n36956, n36957, n36958, n36959,
    n36960, n36961, n36962, n36963, n36964, n36965,
    n36966, n36967, n36968, n36969, n36970, n36971,
    n36972, n36973, n36974, n36975, n36976, n36977,
    n36978, n36979, n36980, n36981, n36982, n36983,
    n36984, n36985, n36986, n36987, n36988, n36989,
    n36990, n36991, n36992, n36993, n36994, n36995,
    n36996, n36997, n36998, n36999, n37000, n37001,
    n37002, n37003, n37004, n37005, n37006, n37007,
    n37008, n37009, n37010, n37011, n37012, n37013,
    n37014, n37015, n37016, n37017, n37018, n37019,
    n37020, n37021, n37022, n37023, n37024, n37025,
    n37026, n37027, n37028, n37029, n37030, n37031,
    n37032, n37033, n37034, n37035, n37036, n37037,
    n37038, n37039, n37040, n37041, n37042, n37043,
    n37044, n37045, n37046, n37047, n37048, n37049,
    n37050, n37051, n37052, n37053, n37054, n37055,
    n37056, n37057, n37058, n37059, n37060, n37061,
    n37062, n37063, n37064, n37065, n37066, n37067,
    n37068, n37069, n37070, n37071, n37072, n37073,
    n37074, n37075, n37076, n37077, n37078, n37079,
    n37080, n37081, n37082, n37083, n37084, n37085,
    n37086, n37087, n37088, n37089, n37090, n37091,
    n37092, n37093, n37094, n37095, n37096, n37097,
    n37098, n37099, n37100, n37101, n37102, n37103,
    n37104, n37105, n37106, n37107, n37108, n37109,
    n37110, n37111, n37112, n37113, n37114, n37115,
    n37116, n37117, n37118, n37119, n37120, n37121,
    n37122, n37123, n37124, n37125, n37127, n37128,
    n37129, n37130, n37131, n37132, n37133, n37134,
    n37135, n37136, n37137, n37138, n37139, n37140,
    n37141, n37142, n37143, n37144, n37145, n37146,
    n37147, n37148, n37149, n37150, n37151, n37152,
    n37153, n37154, n37155, n37156, n37157, n37158,
    n37159, n37160, n37161, n37162, n37163, n37164,
    n37165, n37166, n37167, n37168, n37169, n37170,
    n37171, n37172, n37173, n37174, n37175, n37176,
    n37177, n37178, n37179, n37180, n37181, n37182,
    n37183, n37184, n37185, n37186, n37187, n37188,
    n37189, n37190, n37191, n37192, n37193, n37194,
    n37195, n37196, n37197, n37198, n37199, n37200,
    n37201, n37202, n37203, n37204, n37205, n37206,
    n37207, n37208, n37209, n37210, n37211, n37212,
    n37213, n37214, n37215, n37216, n37217, n37218,
    n37219, n37220, n37221, n37222, n37223, n37224,
    n37225, n37226, n37227, n37228, n37229, n37230,
    n37231, n37232, n37233, n37234, n37235, n37236,
    n37237, n37238, n37239, n37240, n37241, n37242,
    n37243, n37244, n37245, n37246, n37247, n37248,
    n37249, n37250, n37251, n37252, n37253, n37254,
    n37255, n37256, n37257, n37258, n37259, n37260,
    n37261, n37262, n37263, n37264, n37265, n37266,
    n37267, n37268, n37269, n37270, n37271, n37272,
    n37273, n37274, n37275, n37276, n37277, n37278,
    n37279, n37280, n37281, n37282, n37283, n37284,
    n37285, n37286, n37287, n37288, n37289, n37290,
    n37291, n37292, n37293, n37294, n37295, n37296,
    n37298, n37299, n37300, n37301, n37302, n37303,
    n37304, n37305, n37306, n37307, n37308, n37309,
    n37311, n37312, n37313, n37314, n37315, n37316,
    n37317, n37318, n37319, n37320, n37321, n37322,
    n37323, n37324, n37325, n37326, n37327, n37328,
    n37329, n37330, n37331, n37332, n37333, n37334,
    n37335, n37336, n37337, n37338, n37339, n37340,
    n37341, n37342, n37343, n37344, n37345, n37346,
    n37347, n37348, n37349, n37350, n37351, n37352,
    n37353, n37354, n37355, n37356, n37357, n37358,
    n37359, n37360, n37361, n37362, n37363, n37364,
    n37365, n37366, n37367, n37368, n37369, n37370,
    n37371, n37372, n37373, n37374, n37375, n37376,
    n37377, n37378, n37379, n37380, n37381, n37382,
    n37383, n37384, n37385, n37386, n37387, n37388,
    n37389, n37390, n37391, n37392, n37393, n37394,
    n37395, n37396, n37397, n37398, n37399, n37400,
    n37401, n37402, n37403, n37404, n37405, n37406,
    n37407, n37408, n37409, n37410, n37411, n37412,
    n37413, n37414, n37415, n37416, n37417, n37418,
    n37419, n37420, n37421, n37422, n37423, n37424,
    n37425, n37426, n37427, n37428, n37429, n37430,
    n37431, n37432, n37433, n37434, n37435, n37436,
    n37437, n37438, n37439, n37440, n37441, n37442,
    n37443, n37444, n37445, n37446, n37447, n37448,
    n37449, n37450, n37451, n37452, n37453, n37454,
    n37455, n37456, n37457, n37458, n37459, n37460,
    n37461, n37462, n37463, n37464, n37465, n37466,
    n37467, n37468, n37469, n37470, n37471, n37472,
    n37473, n37474, n37475, n37476, n37477, n37478,
    n37479, n37480, n37481, n37482, n37483, n37484,
    n37485, n37486, n37487, n37488, n37489, n37490,
    n37491, n37492, n37493, n37494, n37495, n37496,
    n37497, n37498, n37499, n37500, n37501, n37502,
    n37503, n37504, n37505, n37506, n37507, n37508,
    n37509, n37510, n37511, n37512, n37513, n37514,
    n37515, n37516, n37517, n37518, n37519, n37520,
    n37521, n37522, n37523, n37524, n37525, n37526,
    n37527, n37528, n37529, n37530, n37531, n37532,
    n37533, n37534, n37535, n37536, n37537, n37538,
    n37539, n37540, n37541, n37542, n37543, n37544,
    n37545, n37546, n37547, n37548, n37549, n37550,
    n37551, n37552, n37553, n37554, n37555, n37556,
    n37558, n37559, n37560, n37561, n37562, n37563,
    n37564, n37565, n37566, n37567, n37568, n37569,
    n37570, n37571, n37572, n37573, n37574, n37575,
    n37576, n37577, n37578, n37579, n37580, n37581,
    n37582, n37583, n37584, n37585, n37586, n37587,
    n37588, n37589, n37590, n37591, n37592, n37593,
    n37594, n37595, n37596, n37597, n37598, n37599,
    n37600, n37601, n37602, n37603, n37604, n37605,
    n37606, n37607, n37608, n37609, n37610, n37611,
    n37612, n37613, n37614, n37615, n37616, n37617,
    n37618, n37619, n37620, n37621, n37622, n37623,
    n37624, n37625, n37626, n37627, n37628, n37629,
    n37630, n37631, n37632, n37633, n37634, n37635,
    n37636, n37637, n37638, n37639, n37640, n37641,
    n37642, n37643, n37644, n37645, n37646, n37647,
    n37648, n37649, n37650, n37651, n37652, n37653,
    n37654, n37655, n37656, n37657, n37658, n37659,
    n37660, n37661, n37662, n37663, n37664, n37665,
    n37666, n37667, n37668, n37669, n37670, n37671,
    n37672, n37673, n37674, n37675, n37676, n37677,
    n37678, n37679, n37680, n37681, n37682, n37683,
    n37684, n37685, n37686, n37687, n37688, n37689,
    n37690, n37691, n37692, n37693, n37694, n37695,
    n37696, n37697, n37698, n37699, n37700, n37701,
    n37702, n37703, n37704, n37705, n37706, n37707,
    n37708, n37709, n37710, n37711, n37712, n37713,
    n37714, n37715, n37716, n37717, n37718, n37719,
    n37720, n37721, n37722, n37723, n37724, n37725,
    n37726, n37727, n37728, n37729, n37730, n37731,
    n37732, n37733, n37734, n37735, n37736, n37737,
    n37738, n37739, n37740, n37741, n37742, n37743,
    n37744, n37745, n37746, n37747, n37748, n37749,
    n37750, n37751, n37752, n37753, n37754, n37755,
    n37756, n37757, n37758, n37759, n37760, n37761,
    n37762, n37763, n37764, n37765, n37766, n37767,
    n37768, n37769, n37770, n37771, n37772, n37773,
    n37774, n37775, n37776, n37777, n37778, n37779,
    n37780, n37781, n37782, n37783, n37784, n37785,
    n37786, n37787, n37788, n37789, n37790, n37791,
    n37792, n37793, n37794, n37795, n37796, n37797,
    n37798, n37799, n37800, n37801, n37802, n37803,
    n37804, n37805, n37806, n37807, n37808, n37809,
    n37810, n37811, n37812, n37813, n37814, n37815,
    n37816, n37817, n37818, n37819, n37820, n37821,
    n37822, n37823, n37824, n37825, n37826, n37827,
    n37828, n37829, n37830, n37831, n37832, n37833,
    n37834, n37835, n37836, n37837, n37838, n37839,
    n37840, n37841, n37842, n37843, n37844, n37845,
    n37846, n37847, n37848, n37849, n37850, n37851,
    n37853, n37854, n37855, n37856, n37857, n37858,
    n37859, n37860, n37861, n37862, n37863, n37864,
    n37865, n37866, n37867, n37868, n37869, n37870,
    n37871, n37872, n37873, n37874, n37875, n37876,
    n37877, n37878, n37879, n37880, n37881, n37882,
    n37883, n37884, n37885, n37886, n37887, n37888,
    n37889, n37890, n37891, n37892, n37893, n37894,
    n37895, n37896, n37897, n37898, n37899, n37900,
    n37901, n37902, n37903, n37904, n37905, n37906,
    n37907, n37908, n37909, n37910, n37911, n37912,
    n37913, n37914, n37915, n37916, n37917, n37918,
    n37919, n37920, n37921, n37922, n37923, n37924,
    n37925, n37926, n37927, n37928, n37929, n37930,
    n37931, n37932, n37933, n37934, n37935, n37936,
    n37938, n37939, n37940, n37941, n37942, n37943,
    n37944, n37945, n37946, n37947, n37948, n37949,
    n37950, n37951, n37952, n37953, n37954, n37955,
    n37956, n37957, n37958, n37959, n37960, n37961,
    n37962, n37963, n37964, n37965, n37966, n37967,
    n37968, n37969, n37970, n37971, n37972, n37973,
    n37974, n37975, n37976, n37977, n37978, n37979,
    n37980, n37981, n37982, n37983, n37984, n37985,
    n37986, n37987, n37988, n37989, n37990, n37991,
    n37992, n37993, n37994, n37995, n37996, n37997,
    n37998, n37999, n38000, n38001, n38002, n38003,
    n38004, n38005, n38006, n38007, n38008, n38009,
    n38010, n38011, n38012, n38013, n38014, n38015,
    n38016, n38017, n38018, n38019, n38020, n38021,
    n38022, n38023, n38024, n38025, n38026, n38027,
    n38028, n38029, n38030, n38031, n38032, n38033,
    n38034, n38035, n38036, n38037, n38038, n38039,
    n38040, n38041, n38042, n38043, n38044, n38045,
    n38046, n38047, n38048, n38049, n38050, n38051,
    n38052, n38053, n38054, n38055, n38056, n38057,
    n38058, n38059, n38060, n38061, n38062, n38063,
    n38064, n38065, n38066, n38067, n38068, n38069,
    n38070, n38071, n38072, n38073, n38074, n38075,
    n38076, n38077, n38078, n38079, n38080, n38081,
    n38082, n38083, n38084, n38085, n38086, n38087,
    n38088, n38089, n38090, n38091, n38092, n38093,
    n38094, n38095, n38096, n38097, n38098, n38099,
    n38100, n38101, n38102, n38103, n38104, n38105,
    n38106, n38107, n38108, n38109, n38110, n38111,
    n38112, n38113, n38114, n38115, n38116, n38117,
    n38118, n38119, n38120, n38121, n38122, n38123,
    n38124, n38125, n38126, n38127, n38128, n38129,
    n38130, n38131, n38132, n38133, n38134, n38135,
    n38136, n38137, n38138, n38139, n38140, n38141,
    n38142, n38143, n38144, n38145, n38146, n38147,
    n38148, n38149, n38150, n38151, n38152, n38153,
    n38154, n38155, n38156, n38157, n38158, n38159,
    n38160, n38161, n38162, n38163, n38164, n38165,
    n38166, n38167, n38168, n38169, n38170, n38171,
    n38172, n38173, n38174, n38175, n38176, n38177,
    n38178, n38179, n38180, n38181, n38182, n38183,
    n38184, n38185, n38186, n38187, n38188, n38189,
    n38190, n38191, n38192, n38193, n38194, n38195,
    n38196, n38197, n38198, n38199, n38200, n38201,
    n38202, n38203, n38204, n38205, n38206, n38207,
    n38208, n38209, n38210, n38211, n38212, n38213,
    n38214, n38215, n38216, n38217, n38218, n38219,
    n38220, n38221, n38222, n38223, n38224, n38225,
    n38226, n38227, n38228, n38229, n38230, n38231,
    n38232, n38233, n38234, n38235, n38236, n38237,
    n38238, n38239, n38240, n38241, n38242, n38243,
    n38244, n38245, n38246, n38247, n38248, n38249,
    n38250, n38251, n38252, n38253, n38254, n38255,
    n38256, n38257, n38258, n38259, n38260, n38261,
    n38262, n38263, n38264, n38265, n38266, n38267,
    n38268, n38269, n38270, n38271, n38272, n38273,
    n38274, n38275, n38276, n38277, n38278, n38279,
    n38281, n38282, n38283, n38284, n38285, n38286,
    n38287, n38288, n38289, n38290, n38291, n38292,
    n38293, n38294, n38295, n38296, n38297, n38298,
    n38299, n38300, n38301, n38302, n38303, n38304,
    n38305, n38306, n38307, n38308, n38309, n38310,
    n38311, n38312, n38313, n38314, n38315, n38316,
    n38317, n38318, n38319, n38320, n38321, n38322,
    n38323, n38324, n38325, n38326, n38327, n38328,
    n38329, n38330, n38331, n38332, n38333, n38334,
    n38335, n38336, n38337, n38338, n38339, n38340,
    n38341, n38342, n38343, n38344, n38345, n38346,
    n38347, n38348, n38349, n38350, n38351, n38352,
    n38353, n38354, n38355, n38356, n38357, n38358,
    n38359, n38360, n38361, n38362, n38363, n38364,
    n38365, n38366, n38367, n38368, n38369, n38370,
    n38371, n38372, n38373, n38374, n38375, n38376,
    n38377, n38378, n38379, n38380, n38381, n38382,
    n38383, n38384, n38385, n38386, n38387, n38388,
    n38389, n38390, n38391, n38392, n38393, n38394,
    n38395, n38396, n38397, n38398, n38399, n38400,
    n38401, n38402, n38403, n38404, n38405, n38406,
    n38407, n38408, n38409, n38410, n38411, n38412,
    n38413, n38414, n38415, n38416, n38417, n38418,
    n38419, n38420, n38421, n38422, n38423, n38424,
    n38425, n38426, n38427, n38428, n38429, n38430,
    n38431, n38432, n38433, n38434, n38435, n38436,
    n38437, n38438, n38439, n38440, n38441, n38442,
    n38443, n38444, n38445, n38446, n38447, n38448,
    n38449, n38450, n38451, n38452, n38453, n38454,
    n38455, n38456, n38457, n38458, n38459, n38460,
    n38461, n38462, n38463, n38464, n38465, n38466,
    n38467, n38468, n38469, n38470, n38471, n38472,
    n38473, n38474, n38475, n38476, n38477, n38478,
    n38479, n38480, n38481, n38482, n38483, n38484,
    n38485, n38486, n38487, n38488, n38489, n38490,
    n38491, n38492, n38493, n38494, n38495, n38496,
    n38497, n38498, n38499, n38500, n38501, n38502,
    n38503, n38504, n38505, n38506, n38507, n38508,
    n38509, n38510, n38511, n38512, n38513, n38514,
    n38515, n38516, n38517, n38518, n38519, n38520,
    n38521, n38522, n38523, n38524, n38525, n38526,
    n38527, n38528, n38529, n38530, n38531, n38532,
    n38533, n38534, n38535, n38536, n38537, n38538,
    n38539, n38540, n38541, n38542, n38543, n38544,
    n38545, n38546, n38547, n38548, n38549, n38551,
    n38552, n38553, n38554, n38555, n38556, n38557,
    n38558, n38559, n38560, n38561, n38562, n38563,
    n38564, n38565, n38566, n38567, n38568, n38569,
    n38570, n38571, n38572, n38573, n38574, n38575,
    n38576, n38577, n38578, n38579, n38580, n38581,
    n38582, n38583, n38584, n38585, n38586, n38587,
    n38588, n38589, n38590, n38591, n38592, n38593,
    n38594, n38595, n38596, n38597, n38598, n38599,
    n38600, n38601, n38602, n38603, n38604, n38605,
    n38606, n38607, n38608, n38609, n38610, n38611,
    n38612, n38613, n38614, n38615, n38616, n38618,
    n38619, n38620, n38621, n38622, n38623, n38624,
    n38625, n38626, n38627, n38628, n38629, n38630,
    n38631, n38632, n38633, n38634, n38635, n38636,
    n38637, n38638, n38639, n38640, n38641, n38642,
    n38643, n38644, n38645, n38646, n38647, n38648,
    n38649, n38650, n38651, n38652, n38653, n38654,
    n38655, n38656, n38657, n38658, n38659, n38660,
    n38661, n38662, n38663, n38664, n38665, n38666,
    n38667, n38668, n38669, n38670, n38671, n38672,
    n38673, n38674, n38675, n38676, n38677, n38678,
    n38679, n38680, n38681, n38682, n38683, n38684,
    n38685, n38686, n38687, n38688, n38689, n38690,
    n38691, n38692, n38693, n38694, n38695, n38696,
    n38697, n38698, n38699, n38700, n38701, n38702,
    n38703, n38704, n38705, n38706, n38707, n38708,
    n38709, n38710, n38711, n38712, n38713, n38714,
    n38715, n38716, n38717, n38718, n38719, n38720,
    n38721, n38722, n38723, n38724, n38725, n38726,
    n38727, n38728, n38729, n38730, n38731, n38732,
    n38733, n38734, n38735, n38736, n38737, n38738,
    n38739, n38740, n38741, n38742, n38743, n38744,
    n38745, n38746, n38747, n38748, n38749, n38750,
    n38751, n38752, n38753, n38754, n38755, n38756,
    n38757, n38758, n38759, n38760, n38761, n38762,
    n38763, n38764, n38765, n38766, n38767, n38768,
    n38769, n38770, n38771, n38772, n38773, n38774,
    n38775, n38776, n38777, n38778, n38779, n38780,
    n38781, n38782, n38783, n38784, n38785, n38786,
    n38787, n38788, n38789, n38790, n38791, n38792,
    n38793, n38794, n38795, n38796, n38797, n38798,
    n38799, n38800, n38801, n38802, n38803, n38804,
    n38805, n38806, n38807, n38808, n38809, n38810,
    n38811, n38812, n38813, n38814, n38815, n38816,
    n38817, n38818, n38819, n38820, n38821, n38822,
    n38823, n38824, n38825, n38826, n38827, n38828,
    n38829, n38830, n38831, n38832, n38833, n38834,
    n38835, n38836, n38837, n38838, n38839, n38840,
    n38841, n38842, n38843, n38844, n38845, n38846,
    n38847, n38848, n38849, n38850, n38851, n38852,
    n38853, n38854, n38855, n38856, n38857, n38858,
    n38859, n38860, n38861, n38862, n38863, n38864,
    n38865, n38866, n38867, n38868, n38869, n38870,
    n38871, n38872, n38873, n38874, n38875, n38876,
    n38877, n38878, n38879, n38880, n38881, n38882,
    n38883, n38884, n38885, n38886, n38887, n38888,
    n38889, n38890, n38891, n38892, n38893, n38894,
    n38895, n38896, n38897, n38898, n38899, n38900,
    n38901, n38902, n38903, n38904, n38905, n38906,
    n38907, n38908, n38909, n38910, n38911, n38912,
    n38913, n38914, n38915, n38916, n38917, n38918,
    n38919, n38920, n38921, n38923, n38924, n38925,
    n38926, n38927, n38928, n38929, n38930, n38931,
    n38932, n38933, n38934, n38935, n38936, n38937,
    n38938, n38939, n38940, n38941, n38942, n38943,
    n38944, n38945, n38946, n38947, n38948, n38949,
    n38950, n38951, n38952, n38953, n38954, n38955,
    n38956, n38957, n38958, n38959, n38960, n38961,
    n38962, n38963, n38964, n38965, n38966, n38967,
    n38969, n38970, n38971, n38972, n38973, n38974,
    n38975, n38976, n38977, n38978, n38979, n38980,
    n38981, n38982, n38983, n38984, n38985, n38986,
    n38987, n38988, n38989, n38990, n38991, n38992,
    n38993, n38994, n38995, n38996, n38997, n38998,
    n38999, n39000, n39001, n39002, n39003, n39004,
    n39005, n39006, n39007, n39008, n39009, n39010,
    n39011, n39012, n39013, n39014, n39015, n39016,
    n39017, n39018, n39019, n39020, n39021, n39022,
    n39023, n39024, n39025, n39026, n39027, n39028,
    n39029, n39030, n39031, n39032, n39033, n39034,
    n39035, n39036, n39037, n39038, n39039, n39040,
    n39041, n39042, n39043, n39044, n39045, n39046,
    n39047, n39048, n39049, n39050, n39051, n39052,
    n39053, n39054, n39055, n39056, n39057, n39058,
    n39059, n39060, n39061, n39062, n39063, n39064,
    n39065, n39066, n39067, n39068, n39069, n39070,
    n39071, n39072, n39073, n39074, n39075, n39076,
    n39077, n39078, n39079, n39080, n39081, n39082,
    n39083, n39084, n39085, n39086, n39087, n39088,
    n39089, n39090, n39091, n39092, n39093, n39094,
    n39095, n39096, n39097, n39098, n39099, n39100,
    n39101, n39102, n39103, n39104, n39105, n39106,
    n39107, n39108, n39109, n39110, n39111, n39112,
    n39113, n39114, n39115, n39116, n39117, n39118,
    n39119, n39120, n39121, n39122, n39123, n39124,
    n39125, n39126, n39127, n39128, n39129, n39130,
    n39131, n39132, n39133, n39134, n39135, n39136,
    n39137, n39138, n39139, n39140, n39141, n39142,
    n39143, n39144, n39145, n39146, n39147, n39148,
    n39149, n39150, n39151, n39152, n39153, n39154,
    n39155, n39156, n39157, n39158, n39159, n39160,
    n39161, n39162, n39163, n39164, n39165, n39166,
    n39167, n39168, n39169, n39170, n39172, n39173,
    n39174, n39175, n39176, n39177, n39178, n39179,
    n39180, n39181, n39182, n39183, n39184, n39185,
    n39186, n39187, n39188, n39189, n39190, n39191,
    n39192, n39193, n39194, n39195, n39196, n39197,
    n39198, n39199, n39200, n39201, n39202, n39203,
    n39204, n39205, n39206, n39207, n39208, n39209,
    n39210, n39211, n39212, n39213, n39214, n39215,
    n39216, n39217, n39218, n39219, n39220, n39221,
    n39222, n39223, n39224, n39225, n39226, n39227,
    n39228, n39229, n39230, n39231, n39232, n39233,
    n39234, n39235, n39236, n39237, n39238, n39239,
    n39240, n39241, n39242, n39243, n39244, n39245,
    n39246, n39247, n39248, n39249, n39250, n39251,
    n39252, n39253, n39254, n39255, n39256, n39257,
    n39258, n39259, n39260, n39261, n39262, n39263,
    n39264, n39265, n39266, n39267, n39268, n39269,
    n39270, n39271, n39272, n39273, n39274, n39275,
    n39276, n39277, n39278, n39279, n39280, n39281,
    n39282, n39283, n39284, n39285, n39286, n39287,
    n39288, n39289, n39290, n39291, n39292, n39293,
    n39294, n39295, n39296, n39297, n39298, n39299,
    n39300, n39301, n39302, n39303, n39304, n39305,
    n39306, n39307, n39308, n39309, n39310, n39311,
    n39312, n39313, n39314, n39315, n39316, n39317,
    n39318, n39319, n39320, n39321, n39322, n39323,
    n39324, n39325, n39326, n39327, n39328, n39329,
    n39330, n39331, n39332, n39333, n39334, n39335,
    n39336, n39337, n39338, n39339, n39340, n39341,
    n39342, n39343, n39344, n39345, n39346, n39347,
    n39348, n39349, n39350, n39351, n39352, n39353,
    n39354, n39355, n39356, n39357, n39358, n39359,
    n39360, n39361, n39362, n39363, n39364, n39365,
    n39366, n39367, n39368, n39369, n39370, n39371,
    n39372, n39373, n39374, n39375, n39376, n39377,
    n39378, n39379, n39380, n39381, n39382, n39383,
    n39384, n39385, n39386, n39387, n39388, n39389,
    n39390, n39391, n39392, n39393, n39394, n39395,
    n39396, n39397, n39398, n39399, n39400, n39401,
    n39402, n39404, n39405, n39406, n39407, n39408,
    n39409, n39410, n39411, n39412, n39413, n39414,
    n39415, n39416, n39417, n39418, n39419, n39420,
    n39421, n39422, n39423, n39424, n39425, n39426,
    n39427, n39428, n39429, n39430, n39431, n39432,
    n39433, n39434, n39435, n39436, n39437, n39438,
    n39439, n39440, n39441, n39442, n39443, n39444,
    n39445, n39446, n39447, n39448, n39449, n39450,
    n39451, n39452, n39453, n39454, n39455, n39456,
    n39457, n39458, n39459, n39460, n39461, n39462,
    n39463, n39464, n39465, n39466, n39467, n39468,
    n39469, n39470, n39471, n39472, n39473, n39474,
    n39475, n39476, n39477, n39478, n39479, n39480,
    n39481, n39482, n39483, n39484, n39485, n39486,
    n39487, n39488, n39489, n39490, n39491, n39492,
    n39493, n39494, n39495, n39496, n39497, n39498,
    n39499, n39500, n39501, n39502, n39503, n39504,
    n39505, n39506, n39507, n39508, n39509, n39510,
    n39511, n39512, n39513, n39514, n39515, n39516,
    n39517, n39518, n39519, n39520, n39521, n39522,
    n39523, n39524, n39525, n39526, n39527, n39528,
    n39529, n39530, n39531, n39532, n39533, n39534,
    n39535, n39536, n39537, n39538, n39539, n39540,
    n39541, n39542, n39543, n39544, n39545, n39546,
    n39547, n39548, n39549, n39550, n39551, n39552,
    n39553, n39554, n39555, n39556, n39557, n39558,
    n39559, n39560, n39561, n39562, n39563, n39564,
    n39565, n39566, n39567, n39568, n39569, n39570,
    n39571, n39572, n39573, n39574, n39575, n39576,
    n39577, n39578, n39579, n39580, n39581, n39582,
    n39583, n39584, n39585, n39586, n39587, n39588,
    n39589, n39590, n39591, n39592, n39593, n39594,
    n39595, n39596, n39597, n39598, n39599, n39600,
    n39601, n39602, n39603, n39604, n39605, n39606,
    n39607, n39608, n39609, n39610, n39611, n39612,
    n39613, n39614, n39615, n39616, n39617, n39618,
    n39619, n39620, n39621, n39622, n39624, n39625,
    n39626, n39627, n39628, n39629, n39630, n39631,
    n39632, n39633, n39634, n39635, n39636, n39637,
    n39638, n39639, n39640, n39641, n39642, n39643,
    n39644, n39645, n39646, n39647, n39648, n39649,
    n39650, n39651, n39652, n39653, n39654, n39655,
    n39656, n39657, n39658, n39659, n39660, n39661,
    n39662, n39663, n39664, n39665, n39666, n39667,
    n39668, n39669, n39670, n39671, n39672, n39673,
    n39674, n39675, n39676, n39677, n39678, n39679,
    n39680, n39681, n39682, n39683, n39684, n39685,
    n39686, n39687, n39688, n39689, n39690, n39691,
    n39692, n39693, n39694, n39695, n39696, n39697,
    n39698, n39699, n39700, n39701, n39702, n39703,
    n39704, n39705, n39706, n39707, n39708, n39709,
    n39710, n39711, n39712, n39713, n39714, n39715,
    n39716, n39717, n39718, n39719, n39720, n39721,
    n39722, n39723, n39724, n39725, n39726, n39727,
    n39728, n39729, n39730, n39731, n39732, n39733,
    n39734, n39735, n39736, n39737, n39738, n39739,
    n39740, n39741, n39742, n39743, n39744, n39745,
    n39746, n39747, n39748, n39749, n39750, n39751,
    n39752, n39753, n39754, n39755, n39756, n39757,
    n39758, n39759, n39760, n39761, n39762, n39763,
    n39764, n39765, n39766, n39767, n39768, n39769,
    n39770, n39771, n39772, n39773, n39774, n39775,
    n39776, n39777, n39778, n39779, n39780, n39781,
    n39782, n39783, n39785, n39786, n39787, n39788,
    n39789, n39790, n39791, n39792, n39793, n39794,
    n39795, n39796, n39797, n39798, n39799, n39800,
    n39801, n39802, n39803, n39804, n39805, n39806,
    n39807, n39808, n39809, n39810, n39811, n39812,
    n39813, n39814, n39815, n39816, n39817, n39818,
    n39819, n39820, n39821, n39822, n39823, n39824,
    n39825, n39826, n39827, n39828, n39829, n39830,
    n39831, n39832, n39833, n39834, n39835, n39836,
    n39837, n39838, n39839, n39840, n39841, n39842,
    n39843, n39844, n39845, n39846, n39847, n39848,
    n39849, n39850, n39851, n39852, n39853, n39854,
    n39855, n39856, n39857, n39858, n39859, n39860,
    n39861, n39862, n39863, n39864, n39865, n39866,
    n39867, n39868, n39869, n39870, n39871, n39872,
    n39873, n39874, n39875, n39876, n39877, n39878,
    n39879, n39880, n39881, n39882, n39883, n39884,
    n39885, n39886, n39887, n39888, n39889, n39890,
    n39891, n39892, n39893, n39894, n39895, n39896,
    n39897, n39898, n39899, n39900, n39901, n39902,
    n39903, n39904, n39905, n39906, n39907, n39908,
    n39909, n39910, n39911, n39912, n39913, n39914,
    n39915, n39916, n39917, n39918, n39919, n39920,
    n39921, n39922, n39923, n39924, n39925, n39926,
    n39927, n39928, n39929, n39930, n39931, n39932,
    n39933, n39934, n39935, n39936, n39937, n39938,
    n39940, n39941, n39942, n39943, n39944, n39945,
    n39946, n39948, n39949, n39950, n39951, n39952,
    n39953, n39954, n39955, n39956, n39958, n39959,
    n39960, n39961, n39962, n39963, n39964, n39965,
    n39966, n39967, n39968, n39969, n39970, n39971,
    n39972, n39973, n39974, n39975, n39976, n39977,
    n39978, n39979, n39980, n39981, n39982, n39983,
    n39984, n39985, n39986, n39987, n39988, n39989,
    n39990, n39991, n39992, n39993, n39994, n39995,
    n39996, n39997, n39998, n40000, n40001, n40002,
    n40003, n40004, n40005, n40006, n40007, n40008,
    n40009, n40010, n40011, n40012, n40013, n40014,
    n40015, n40016, n40017, n40018, n40019, n40020,
    n40021, n40022, n40023, n40024, n40025, n40026,
    n40027, n40028, n40029, n40030, n40031, n40032,
    n40033, n40034, n40035, n40036, n40037, n40038,
    n40039, n40040, n40041, n40042, n40043, n40044,
    n40045, n40046, n40047, n40048, n40049, n40050,
    n40051, n40052, n40053, n40054, n40055, n40056,
    n40057, n40058, n40059, n40060, n40061, n40062,
    n40063, n40064, n40065, n40066, n40067, n40068,
    n40069, n40070, n40071, n40072, n40073, n40074,
    n40075, n40076, n40077, n40078, n40079, n40080,
    n40081, n40082, n40083, n40084, n40085, n40086,
    n40087, n40088, n40089, n40090, n40091, n40092,
    n40093, n40094, n40095, n40096, n40097, n40098,
    n40099, n40100, n40101, n40102, n40103, n40104,
    n40105, n40106, n40107, n40108, n40109, n40110,
    n40111, n40112, n40113, n40114, n40115, n40116,
    n40117, n40118, n40119, n40120, n40121, n40122,
    n40123, n40124, n40125, n40126, n40127, n40128,
    n40129, n40130, n40131, n40132, n40133, n40134,
    n40135, n40136, n40137, n40138, n40139, n40140,
    n40141, n40142, n40143, n40144, n40145, n40146,
    n40147, n40148, n40149, n40150, n40151, n40152,
    n40153, n40154, n40155, n40156, n40157, n40158,
    n40159, n40160, n40161, n40162, n40163, n40164,
    n40165, n40166, n40167, n40168, n40169, n40170,
    n40171, n40172, n40173, n40174, n40175, n40176,
    n40177, n40178, n40179, n40180, n40181, n40182,
    n40183, n40184, n40185, n40186, n40187, n40188,
    n40189, n40190, n40191, n40192, n40193, n40194,
    n40195, n40196, n40197, n40198, n40199, n40200,
    n40201, n40202, n40203, n40204, n40205, n40206,
    n40207, n40208, n40209, n40210, n40211, n40212,
    n40213, n40214, n40215, n40216, n40217, n40219,
    n40220, n40221, n40222, n40223, n40224, n40225,
    n40226, n40227, n40228, n40229, n40230, n40231,
    n40232, n40233, n40234, n40235, n40236, n40237,
    n40238, n40239, n40240, n40241, n40242, n40243,
    n40244, n40245, n40246, n40247, n40248, n40249,
    n40250, n40251, n40252, n40253, n40254, n40255,
    n40256, n40257, n40258, n40259, n40260, n40261,
    n40262, n40263, n40264, n40265, n40266, n40267,
    n40268, n40269, n40270, n40271, n40272, n40273,
    n40274, n40275, n40276, n40277, n40278, n40279,
    n40280, n40281, n40282, n40283, n40284, n40285,
    n40286, n40287, n40288, n40289, n40290, n40291,
    n40292, n40293, n40294, n40295, n40296, n40297,
    n40298, n40299, n40300, n40301, n40302, n40303,
    n40304, n40305, n40306, n40307, n40308, n40309,
    n40310, n40311, n40312, n40313, n40314, n40315,
    n40316, n40317, n40318, n40319, n40320, n40321,
    n40322, n40323, n40324, n40325, n40326, n40327,
    n40328, n40329, n40330, n40331, n40332, n40333,
    n40334, n40335, n40336, n40337, n40338, n40339,
    n40340, n40341, n40342, n40343, n40344, n40345,
    n40346, n40347, n40348, n40349, n40350, n40351,
    n40352, n40353, n40354, n40355, n40356, n40357,
    n40358, n40359, n40360, n40361, n40362, n40363,
    n40364, n40365, n40366, n40367, n40368, n40369,
    n40370, n40371, n40372, n40373, n40374, n40375,
    n40376, n40377, n40378, n40379, n40380, n40381,
    n40382, n40383, n40384, n40385, n40386, n40387,
    n40388, n40389, n40390, n40391, n40392, n40393,
    n40394, n40395, n40396, n40397, n40398, n40399,
    n40400, n40401, n40402, n40403, n40404, n40405,
    n40406, n40407, n40408, n40409, n40410, n40411,
    n40412, n40413, n40414, n40415, n40416, n40417,
    n40418, n40419, n40420, n40421, n40423, n40424,
    n40425, n40426, n40427, n40429, n40430, n40431,
    n40432, n40433, n40435, n40436, n40437, n40438,
    n40439, n40441, n40442, n40443, n40444, n40445,
    n40447, n40448, n40449, n40450, n40451, n40453,
    n40454, n40455, n40456, n40457, n40458, n40460,
    n40461, n40462, n40463, n40464, n40465, n40467,
    n40468, n40469, n40470, n40471, n40472, n40473,
    n40474, n40475, n40476, n40477, n40478, n40479,
    n40480, n40481, n40482, n40483, n40484, n40485,
    n40486, n40487, n40488, n40489, n40490, n40491,
    n40492, n40493, n40494, n40495, n40497, n40498,
    n40499, n40500, n40501, n40502, n40503, n40504,
    n40505, n40506, n40507, n40508, n40509, n40510,
    n40511, n40512, n40513, n40514, n40515, n40516,
    n40517, n40518, n40519, n40520, n40521, n40522,
    n40523, n40524, n40525, n40526, n40527, n40528,
    n40529, n40530, n40531, n40532, n40533, n40534,
    n40535, n40536, n40537, n40538, n40539, n40540,
    n40541, n40542, n40543, n40544, n40545, n40546,
    n40547, n40548, n40549, n40550, n40551, n40552,
    n40553, n40554, n40555, n40556, n40557, n40558,
    n40559, n40560, n40561, n40562, n40563, n40564,
    n40565, n40566, n40567, n40568, n40569, n40570,
    n40571, n40572, n40573, n40574, n40575, n40576,
    n40577, n40578, n40579, n40580, n40581, n40582,
    n40583, n40584, n40585, n40586, n40587, n40588,
    n40589, n40590, n40591, n40592, n40593, n40594,
    n40595, n40596, n40597, n40598, n40599, n40600,
    n40601, n40602, n40603, n40604, n40605, n40606,
    n40607, n40608, n40609, n40610, n40611, n40612,
    n40613, n40614, n40615, n40616, n40617, n40618,
    n40619, n40620, n40621, n40622, n40623, n40624,
    n40625, n40626, n40627, n40628, n40629, n40630,
    n40631, n40632, n40633, n40634, n40635, n40636,
    n40637, n40638, n40639, n40640, n40641, n40642,
    n40643, n40644, n40645, n40646, n40647, n40648,
    n40649, n40650, n40651, n40652, n40653, n40654,
    n40655, n40656, n40657, n40658, n40659, n40660,
    n40661, n40662, n40663, n40664, n40665, n40666,
    n40667, n40668, n40669, n40670, n40671, n40672,
    n40673, n40674, n40675, n40676, n40677, n40678,
    n40679, n40680, n40681, n40682, n40683, n40684,
    n40686, n40687, n40688, n40689, n40690, n40691,
    n40692, n40693, n40694, n40695, n40696, n40697,
    n40698, n40699, n40700, n40701, n40702, n40703,
    n40704, n40705, n40706, n40707, n40708, n40709,
    n40710, n40711, n40712, n40713, n40714, n40715,
    n40716, n40717, n40718, n40719, n40720, n40721,
    n40722, n40723, n40724, n40725, n40726, n40727,
    n40728, n40729, n40731, n40732, n40733, n40734,
    n40735, n40736, n40737, n40738, n40739, n40740,
    n40741, n40742, n40743, n40744, n40745, n40746,
    n40747, n40748, n40749, n40750, n40751, n40752,
    n40753, n40754, n40755, n40756, n40757, n40758,
    n40759, n40760, n40761, n40762, n40763, n40764,
    n40765, n40766, n40767, n40768, n40769, n40771,
    n40772, n40773, n40774, n40775, n40776, n40777,
    n40778, n40779, n40780, n40781, n40782, n40783,
    n40784, n40785, n40786, n40787, n40788, n40789,
    n40790, n40791, n40792, n40793, n40794, n40795,
    n40796, n40797, n40798, n40799, n40800, n40801,
    n40802, n40803, n40804, n40805, n40806, n40807,
    n40808, n40809, n40810, n40811, n40812, n40813,
    n40814, n40815, n40816, n40817, n40818, n40819,
    n40820, n40821, n40822, n40823, n40824, n40825,
    n40826, n40827, n40828, n40829, n40830, n40831,
    n40832, n40833, n40834, n40835, n40836, n40838,
    n40839, n40840, n40841, n40842, n40843, n40844,
    n40845, n40846, n40847, n40848, n40849, n40850,
    n40851, n40852, n40853, n40854, n40855, n40856,
    n40857, n40858, n40859, n40860, n40861, n40862,
    n40863, n40864, n40865, n40866, n40867, n40868,
    n40869, n40870, n40871, n40872, n40873, n40874,
    n40875, n40876, n40877, n40878, n40879, n40880,
    n40881, n40882, n40883, n40884, n40885, n40886,
    n40887, n40888, n40889, n40890, n40891, n40892,
    n40893, n40894, n40895, n40896, n40897, n40898,
    n40899, n40900, n40901, n40902, n40903, n40904,
    n40905, n40906, n40907, n40908, n40909, n40910,
    n40911, n40912, n40913, n40914, n40915, n40916,
    n40917, n40918, n40919, n40920, n40921, n40922,
    n40923, n40924, n40925, n40926, n40927, n40928,
    n40929, n40930, n40931, n40932, n40933, n40934,
    n40935, n40936, n40937, n40938, n40939, n40940,
    n40941, n40942, n40943, n40944, n40945, n40946,
    n40947, n40948, n40949, n40950, n40951, n40952,
    n40953, n40954, n40955, n40956, n40957, n40958,
    n40959, n40960, n40961, n40962, n40963, n40964,
    n40965, n40966, n40967, n40968, n40969, n40970,
    n40971, n40972, n40973, n40974, n40975, n40976,
    n40977, n40978, n40979, n40980, n40981, n40982,
    n40983, n40984, n40985, n40986, n40987, n40988,
    n40989, n40990, n40991, n40992, n40993, n40994,
    n40995, n40996, n40997, n40998, n40999, n41000,
    n41001, n41002, n41003, n41004, n41005, n41006,
    n41007, n41008, n41009, n41010, n41011, n41012,
    n41013, n41014, n41015, n41016, n41017, n41018,
    n41019, n41020, n41021, n41022, n41023, n41024,
    n41025, n41027, n41028, n41029, n41030, n41031,
    n41032, n41033, n41034, n41035, n41036, n41037,
    n41038, n41039, n41040, n41041, n41042, n41043,
    n41044, n41045, n41046, n41047, n41048, n41049,
    n41050, n41051, n41052, n41053, n41054, n41055,
    n41056, n41057, n41058, n41059, n41060, n41061,
    n41062, n41063, n41064, n41065, n41066, n41067,
    n41068, n41069, n41070, n41071, n41072, n41073,
    n41074, n41075, n41076, n41077, n41078, n41079,
    n41080, n41081, n41082, n41083, n41084, n41085,
    n41086, n41087, n41088, n41089, n41090, n41091,
    n41092, n41093, n41094, n41095, n41096, n41097,
    n41098, n41099, n41100, n41101, n41102, n41103,
    n41104, n41105, n41106, n41107, n41108, n41109,
    n41110, n41111, n41112, n41113, n41114, n41115,
    n41116, n41117, n41118, n41119, n41120, n41121,
    n41122, n41123, n41124, n41125, n41126, n41127,
    n41128, n41129, n41130, n41131, n41132, n41133,
    n41134, n41135, n41136, n41137, n41138, n41139,
    n41140, n41141, n41142, n41143, n41144, n41145,
    n41146, n41147, n41148, n41149, n41150, n41151,
    n41152, n41153, n41154, n41155, n41156, n41157,
    n41158, n41159, n41160, n41161, n41162, n41163,
    n41164, n41165, n41166, n41167, n41168, n41169,
    n41170, n41171, n41173, n41174, n41175, n41176,
    n41177, n41178, n41179, n41180, n41181, n41182,
    n41183, n41184, n41185, n41186, n41187, n41188,
    n41189, n41190, n41191, n41192, n41193, n41194,
    n41195, n41196, n41197, n41198, n41199, n41200,
    n41201, n41202, n41203, n41204, n41205, n41206,
    n41207, n41208, n41209, n41210, n41211, n41212,
    n41213, n41214, n41215, n41216, n41218, n41219,
    n41220, n41221, n41222, n41223, n41224, n41225,
    n41226, n41227, n41228, n41229, n41230, n41231,
    n41232, n41233, n41234, n41235, n41236, n41237,
    n41238, n41239, n41240, n41241, n41242, n41243,
    n41244, n41245, n41246, n41247, n41248, n41249,
    n41250, n41251, n41252, n41253, n41254, n41255,
    n41256, n41257, n41258, n41259, n41261, n41262,
    n41263, n41264, n41265, n41266, n41267, n41268,
    n41269, n41270, n41271, n41272, n41273, n41274,
    n41275, n41276, n41277, n41278, n41279, n41280,
    n41281, n41282, n41283, n41284, n41285, n41286,
    n41287, n41288, n41289, n41290, n41291, n41292,
    n41293, n41294, n41295, n41296, n41297, n41298,
    n41299, n41300, n41301, n41302, n41303, n41304,
    n41305, n41306, n41308, n41309, n41310, n41311,
    n41312, n41313, n41314, n41315, n41316, n41317,
    n41318, n41319, n41320, n41321, n41322, n41323,
    n41324, n41325, n41326, n41327, n41328, n41329,
    n41330, n41331, n41332, n41333, n41334, n41335,
    n41336, n41337, n41338, n41339, n41340, n41341,
    n41342, n41343, n41344, n41345, n41346, n41347,
    n41348, n41349, n41350, n41351, n41352, n41353,
    n41354, n41355, n41356, n41357, n41358, n41359,
    n41360, n41361, n41362, n41363, n41364, n41365,
    n41366, n41367, n41368, n41369, n41370, n41371,
    n41372, n41373, n41374, n41375, n41376, n41377,
    n41378, n41380, n41381, n41382, n41383, n41384,
    n41385, n41386, n41387, n41388, n41389, n41390,
    n41391, n41392, n41393, n41394, n41395, n41396,
    n41397, n41398, n41399, n41400, n41401, n41402,
    n41403, n41404, n41405, n41406, n41407, n41408,
    n41409, n41410, n41411, n41412, n41413, n41414,
    n41415, n41416, n41417, n41418, n41419, n41420,
    n41421, n41422, n41423, n41424, n41425, n41426,
    n41427, n41428, n41429, n41431, n41432, n41433,
    n41434, n41435, n41436, n41437, n41438, n41439,
    n41440, n41441, n41442, n41443, n41444, n41445,
    n41446, n41447, n41448, n41449, n41450, n41451,
    n41452, n41453, n41454, n41455, n41456, n41457,
    n41458, n41459, n41460, n41461, n41462, n41463,
    n41464, n41465, n41466, n41467, n41468, n41469,
    n41470, n41472, n41473, n41474, n41475, n41476,
    n41477, n41478, n41479, n41480, n41481, n41482,
    n41483, n41484, n41485, n41486, n41487, n41488,
    n41489, n41490, n41491, n41492, n41493, n41494,
    n41495, n41496, n41497, n41498, n41499, n41500,
    n41501, n41502, n41503, n41504, n41505, n41506,
    n41507, n41508, n41509, n41510, n41511, n41512,
    n41513, n41514, n41515, n41516, n41517, n41518,
    n41519, n41520, n41521, n41522, n41523, n41524,
    n41525, n41526, n41527, n41528, n41529, n41530,
    n41531, n41532, n41533, n41534, n41535, n41536,
    n41537, n41538, n41539, n41540, n41541, n41542,
    n41544, n41545, n41546, n41547, n41548, n41549,
    n41550, n41551, n41552, n41553, n41554, n41555,
    n41556, n41557, n41558, n41559, n41560, n41561,
    n41562, n41563, n41564, n41565, n41566, n41567,
    n41568, n41569, n41570, n41571, n41572, n41574,
    n41575, n41576, n41577, n41578, n41579, n41580,
    n41581, n41582, n41583, n41584, n41585, n41586,
    n41587, n41588, n41589, n41590, n41591, n41592,
    n41593, n41594, n41595, n41596, n41597, n41598,
    n41599, n41600, n41601, n41602, n41603, n41604,
    n41605, n41606, n41607, n41608, n41609, n41610,
    n41611, n41612, n41613, n41614, n41615, n41617,
    n41618, n41619, n41620, n41621, n41622, n41623,
    n41624, n41625, n41626, n41627, n41628, n41629,
    n41630, n41631, n41632, n41633, n41634, n41635,
    n41636, n41637, n41638, n41639, n41640, n41641,
    n41642, n41643, n41644, n41645, n41646, n41647,
    n41648, n41649, n41650, n41651, n41652, n41653,
    n41654, n41655, n41656, n41657, n41658, n41659,
    n41660, n41661, n41662, n41663, n41664, n41665,
    n41666, n41667, n41668, n41669, n41670, n41671,
    n41672, n41673, n41674, n41675, n41676, n41677,
    n41678, n41679, n41680, n41681, n41683, n41684,
    n41685, n41686, n41687, n41688, n41689, n41690,
    n41691, n41692, n41693, n41694, n41695, n41696,
    n41697, n41698, n41699, n41700, n41701, n41702,
    n41703, n41704, n41705, n41706, n41707, n41708,
    n41709, n41710, n41711, n41712, n41713, n41714,
    n41715, n41716, n41717, n41718, n41719, n41720,
    n41721, n41722, n41723, n41724, n41725, n41726,
    n41727, n41728, n41729, n41730, n41731, n41732,
    n41733, n41734, n41735, n41736, n41737, n41738,
    n41739, n41740, n41742, n41743, n41744, n41745,
    n41746, n41747, n41748, n41749, n41750, n41751,
    n41752, n41753, n41754, n41755, n41756, n41757,
    n41758, n41759, n41760, n41761, n41762, n41763,
    n41764, n41765, n41766, n41767, n41768, n41769,
    n41770, n41771, n41772, n41773, n41774, n41775,
    n41776, n41777, n41778, n41779, n41780, n41781,
    n41782, n41783, n41784, n41786, n41787, n41788,
    n41789, n41790, n41791, n41792, n41793, n41794,
    n41795, n41796, n41797, n41798, n41799, n41800,
    n41801, n41802, n41803, n41804, n41805, n41806,
    n41807, n41808, n41809, n41810, n41811, n41812,
    n41813, n41814, n41815, n41816, n41817, n41818,
    n41819, n41820, n41821, n41822, n41823, n41825,
    n41826, n41827, n41828, n41829, n41830, n41831,
    n41832, n41833, n41834, n41835, n41836, n41837,
    n41838, n41839, n41840, n41841, n41842, n41843,
    n41844, n41845, n41846, n41847, n41848, n41849,
    n41850, n41851, n41852, n41853, n41854, n41855,
    n41856, n41857, n41858, n41859, n41860, n41861,
    n41862, n41864, n41865, n41866, n41867, n41868,
    n41869, n41870, n41871, n41872, n41873, n41874,
    n41875, n41876, n41877, n41878, n41879, n41880,
    n41881, n41882, n41883, n41884, n41885, n41886,
    n41887, n41888, n41889, n41890, n41891, n41892,
    n41893, n41894, n41895, n41896, n41897, n41898,
    n41899, n41900, n41901, n41902, n41903, n41904,
    n41905, n41906, n41907, n41908, n41909, n41910,
    n41911, n41912, n41913, n41914, n41915, n41916,
    n41917, n41918, n41919, n41920, n41921, n41923,
    n41924, n41925, n41927, n41929, n41930, n41931,
    n41932, n41933, n41934, n41935, n41936, n41937,
    n41938, n41939, n41940, n41941, n41942, n41943,
    n41944, n41946, n41947, n41948, n41949, n41950,
    n41951, n41952, n41953, n41954, n41955, n41956,
    n41957, n41958, n41959, n41960, n41961, n41962,
    n41964, n41966, n41967, n41968, n41969, n41970,
    n41972, n41973, n41974, n41975, n41976, n41977,
    n41978, n41979, n41980, n41981, n41982, n41983,
    n41985, n41986, n41988, n41989, n41991, n41992,
    n41994, n41995, n41997, n41998, n42000, n42001,
    n42003, n42004, n42006, n42007, n42009, n42010,
    n42012, n42013, n42014, n42015, n42016, n42017,
    n42018, n42020, n42021, n42022, n42023, n42024,
    n42025, n42027, n42028, n42029, n42030, n42032,
    n42033, n42034, n42035, n42036, n42037, n42038,
    n42039, n42040, n42041, n42042, n42043, n42044,
    n42045, n42046, n42047, n42048, n42049, n42050,
    n42051, n42053, n42054, n42056, n42057, n42059,
    n42060, n42062, n42063, n42065, n42066, n42068,
    n42069, n42071, n42072, n42074, n42075, n42076,
    n42077, n42078, n42079, n42080, n42081, n42082,
    n42083, n42084, n42085, n42086, n42087, n42088,
    n42089, n42090, n42091, n42092, n42094, n42095,
    n42096, n42098, n42099, n42101, n42102, n42103,
    n42105, n42106, n42108, n42109, n42110, n42111,
    n42112, n42113, n42114, n42115, n42116, n42117,
    n42118, n42120, n42121, n42122, n42123, n42125,
    n42126, n42128, n42129, n42130, n42132, n42133,
    n42134, n42135, n42137, n42138, n42140, n42141,
    n42143, n42144, n42146, n42147, n42149, n42150,
    n42152, n42153, n42155, n42156, n42158, n42159,
    n42161, n42162, n42164, n42165, n42167, n42168,
    n42170, n42171, n42172, n42173, n42174, n42175,
    n42176, n42178, n42179, n42180, n42181, n42183,
    n42184, n42185, n42186, n42187, n42188, n42189,
    n42190, n42191, n42192, n42193, n42195, n42196,
    n42198, n42199, n42201, n42202, n42204, n42205,
    n42207, n42208, n42210, n42211, n42213, n42214,
    n42216, n42217, n42218, n42219, n42220, n42222,
    n42223, n42225, n42226, n42228, n42229, n42231,
    n42232, n42234, n42235, n42237, n42238, n42240,
    n42241, n42243, n42244, n42246, n42247, n42249,
    n42250, n42252, n42253, n42255, n42256, n42258,
    n42259, n42261, n42262, n42264, n42265, n42267,
    n42268, n42270, n42271, n42273, n42274, n42276,
    n42277, n42279, n42280, n42282, n42283, n42285,
    n42286, n42288, n42289, n42291, n42292, n42294,
    n42295, n42297, n42298, n42300, n42301, n42303,
    n42304, n42306, n42307, n42309, n42310, n42312,
    n42313, n42315, n42316, n42318, n42319, n42321,
    n42322, n42324, n42325, n42327, n42328, n42330,
    n42331, n42333, n42334, n42336, n42337, n42339,
    n42340, n42342, n42343, n42345, n42346, n42348,
    n42349, n42351, n42352, n42354, n42355, n42357,
    n42358, n42360, n42361, n42363, n42364, n42366,
    n42367, n42369, n42370, n42372, n42373, n42375,
    n42376, n42378, n42379, n42381, n42382, n42384,
    n42385, n42387, n42388, n42390, n42391, n42393,
    n42394, n42396, n42397, n42399, n42400, n42402,
    n42403, n42405, n42406, n42408, n42409, n42411,
    n42412, n42414, n42415, n42417, n42418, n42420,
    n42421, n42423, n42424, n42426, n42427, n42429,
    n42430, n42432, n42433, n42435, n42436, n42438,
    n42439, n42441, n42442, n42443, n42445, n42446,
    n42448, n42449, n42451, n42452, n42454, n42455,
    n42457, n42458, n42460, n42461, n42463, n42464,
    n42466, n42467, n42469, n42470, n42472, n42473,
    n42475, n42476, n42478, n42479, n42481, n42482,
    n42484, n42485, n42487, n42488, n42490, n42491,
    n42493, n42494, n42496, n42497, n42499, n42500,
    n42502, n42503, n42505, n42506, n42508, n42509,
    n42511, n42512, n42514, n42515, n42517, n42518,
    n42520, n42521, n42523, n42524, n42526, n42527,
    n42529, n42530, n42532, n42533, n42535, n42536,
    n42538, n42539, n42541, n42542, n42544, n42545,
    n42547, n42548, n42550, n42551, n42553, n42554,
    n42556, n42557, n42559, n42560, n42562, n42563,
    n42565, n42566, n42568, n42569, n42571, n42572,
    n42573, n42574, n42575, n42576, n42577, n42578,
    n42579, n42580, n42581, n42582, n42583, n42584,
    n42585, n42586, n42587, n42588, n42589, n42590,
    n42591, n42592, n42593, n42595, n42596, n42598,
    n42599, n42601, n42602, n42604, n42605, n42607,
    n42608, n42610, n42611, n42613, n42614, n42616,
    n42617, n42618, n42619, n42620, n42621, n42622,
    n42623, n42624, n42625, n42626, n42627, n42628,
    n42629, n42630, n42631, n42632, n42633, n42634,
    n42635, n42636, n42637, n42638, n42640, n42641,
    n42642, n42643, n42644, n42645, n42646, n42647,
    n42648, n42649, n42650, n42651, n42652, n42653,
    n42654, n42655, n42656, n42658, n42659, n42660,
    n42661, n42662, n42663, n42664, n42665, n42666,
    n42667, n42668, n42669, n42670, n42671, n42672,
    n42673, n42674, n42675, n42676, n42677, n42678,
    n42679, n42680, n42681, n42682, n42683, n42684,
    n42685, n42687, n42688, n42689, n42690, n42692,
    n42693, n42694, n42695, n42696, n42697, n42698,
    n42699, n42700, n42701, n42702, n42703, n42704,
    n42705, n42706, n42707, n42708, n42709, n42711,
    n42712, n42713, n42714, n42715, n42716, n42717,
    n42718, n42719, n42720, n42721, n42722, n42723,
    n42724, n42725, n42726, n42727, n42728, n42730,
    n42731, n42732, n42733, n42734, n42735, n42736,
    n42737, n42738, n42739, n42740, n42741, n42742,
    n42743, n42744, n42745, n42746, n42747, n42749,
    n42750, n42751, n42752, n42753, n42754, n42755,
    n42756, n42757, n42758, n42759, n42760, n42761,
    n42762, n42763, n42764, n42765, n42766, n42768,
    n42769, n42770, n42771, n42772, n42773, n42774,
    n42775, n42776, n42778, n42779, n42780, n42781,
    n42782, n42783, n42784, n42785, n42786, n42788,
    n42789, n42790, n42791, n42792, n42793, n42794,
    n42795, n42796, n42798, n42799, n42800, n42801,
    n42802, n42803, n42804, n42805, n42806, n42807,
    n42810, n42811, n42813, n42814, n42816, n42817,
    n42819, n42820, n42822, n42823, n42825, n42826,
    n42828, n42829, n42831, n42832, n42834, n42835,
    n42837, n42838, n42840, n42841, n42843, n42844,
    n42846, n42847, n42849, n42850, n42852, n42853,
    n42855, n42856, n42858, n42859, n42861, n42862,
    n42864, n42865, n42867, n42868, n42870, n42871,
    n42873, n42874, n42876, n42877, n42879, n42880,
    n42882, n42883, n42884, n42886, n42887, n42889,
    n42890, n42892, n42893, n42895, n42896, n42898,
    n42899, n42901, n42902, n42903, n42904, n42905,
    n42907, n42908, n42910, n42911, n42913, n42914,
    n42916, n42917, n42919, n42920, n42922, n42923,
    n42925, n42926, n42927, n42929, n42930, n42932,
    n42933, n42935, n42936, n42938, n42939, n42941,
    n42942, n42944, n42945, n42947, n42948, n42950,
    n42951, n42953, n42954, n42956, n42957, n42959,
    n42960, n42962, n42963, n42965, n42966, n42968,
    n42969, n42971, n42972, n42974, n42975, n42977,
    n42978, n42980, n42981, n42983, n42984, n42986,
    n42987, n42989, n42990, n42992, n42993, n42995,
    n42996, n42998, n42999, n43001, n43002, n43004,
    n43005, n43007, n43008, n43010, n43011, n43013,
    n43014, n43016, n43017, n43019, n43020, n43022,
    n43023, n43025, n43026, n43028, n43029, n43031,
    n43032, n43034, n43035, n43037, n43038, n43040,
    n43041, n43043, n43044, n43046, n43047, n43049,
    n43050, n43052, n43053, n43055, n43056, n43058,
    n43059, n43061, n43062, n43064, n43065, n43067,
    n43068, n43070, n43071, n43073, n43074, n43075,
    n43076, n43077, n43078, n43079, n43080, n43081,
    n43082, n43083, n43084, n43085, n43086, n43087,
    n43088, n43089, n43090, n43091, n43092, n43093,
    n43094, n43095, n43096, n43097, n43098, n43099,
    n43100, n43101, n43102, n43103, n43104, n43105,
    n43106, n43107, n43108, n43109, n43110, n43111,
    n43112, n43113, n43114, n43115, n43116, n43117,
    n43118, n43119, n43120, n43121, n43122, n43123,
    n43124, n43125, n43126, n43127, n43128, n43129,
    n43130, n43131, n43132, n43133, n43134, n43135,
    n43136, n43137, n43138, n43139, n43140, n43141,
    n43142, n43143, n43144, n43145, n43146, n43147,
    n43148, n43149, n43150, n43151, n43152, n43153,
    n43154, n43155, n43156, n43157, n43158, n43159,
    n43160, n43161, n43162, n43163, n43164, n43165,
    n43167, n43168, n43170, n43171, n43173, n43174,
    n43176, n43177, n43179, n43180, n43182, n43183,
    n43185, n43186, n43188, n43189, n43191, n43192,
    n43194, n43195, n43197, n43198, n43200, n43201,
    n43203, n43204, n43206, n43207, n43209, n43210,
    n43212, n43213, n43215, n43216, n43218, n43219,
    n43221, n43222, n43223, n43224, n43225, n43227,
    n43228, n43229, n43230, n43232, n43233, n43234,
    n43235, n43236, n43237, n43238, n43239, n43240,
    n43241, n43242, n43243, n43244, n43245, n43246,
    n43247, n43248, n43249, n43250, n43251, n43252,
    n43253, n43255, n43256, n43257, n43259, n43260,
    n43261, n43263, n43264, n43265, n43267, n43268,
    n43269, n43270, n43271, n43272, n43273, n43274,
    n43275, n43276, n43277, n43278, n43279, n43280,
    n43281, n43282, n43283, n43284, n43285, n43286,
    n43287, n43288, n43289, n43290, n43291, n43292,
    n43293, n43294, n43295, n43296, n43297, n43298,
    n43299, n43300, n43301, n43302, n43303, n43304,
    n43305, n43306, n43307, n43308, n43309, n43310,
    n43311, n43312, n43313, n43314, n43315, n43316,
    n43317, n43318, n43319, n43320, n43321, n43322,
    n43323, n43324, n43325, n43326, n43327, n43328,
    n43329, n43330, n43331, n43332, n43333, n43334,
    n43335, n43336, n43337, n43338, n43339, n43340,
    n43341, n43342, n43343, n43344, n43345, n43346,
    n43347, n43348, n43349, n43350, n43351, n43352,
    n43353, n43354, n43355, n43356, n43357, n43358,
    n43359, n43360, n43361, n43362, n43363, n43364,
    n43365, n43366, n43367, n43368, n43369, n43370,
    n43371, n43372, n43373, n43374, n43375, n43376,
    n43377, n43378, n43379, n43380, n43381, n43382,
    n43383, n43384, n43385, n43386, n43387, n43388,
    n43389, n43390, n43391, n43392, n43393, n43394,
    n43395, n43396, n43397, n43398, n43399, n43400,
    n43401, n43402, n43403, n43404, n43405, n43406,
    n43407, n43408, n43409, n43410, n43411, n43412,
    n43413, n43414, n43415, n43416, n43417, n43418,
    n43419, n43420, n43421, n43422, n43423, n43424,
    n43425, n43426, n43427, n43428, n43429, n43430,
    n43431, n43432, n43433, n43434, n43435, n43436,
    n43437, n43438, n43439, n43440, n43441, n43442,
    n43443, n43444, n43445, n43446, n43447, n43448,
    n43449, n43450, n43451, n43452, n43453, n43454,
    n43455, n43456, n43457, n43458, n43459, n43460,
    n43461, n43462, n43463, n43464, n43465, n43466,
    n43467, n43468, n43469, n43470, n43471, n43472,
    n43473, n43474, n43475, n43476, n43477, n43478,
    n43479, n43480, n43481, n43482, n43483, n43484,
    n43485, n43486, n43487, n43488, n43489, n43490,
    n43491, n43492, n43493, n43494, n43495, n43496,
    n43497, n43498, n43499, n43500, n43501, n43502,
    n43503, n43504, n43505, n43506, n43507, n43508,
    n43509, n43510, n43511, n43512, n43513, n43514,
    n43515, n43516, n43517, n43518, n43519, n43520,
    n43521, n43522, n43523, n43524, n43525, n43526,
    n43527, n43528, n43529, n43530, n43531, n43532,
    n43533, n43534, n43535, n43536, n43537, n43538,
    n43539, n43540, n43541, n43542, n43543, n43544,
    n43545, n43546, n43547, n43548, n43549, n43550,
    n43551, n43552, n43553, n43554, n43555, n43556,
    n43557, n43558, n43559, n43560, n43561, n43562,
    n43563, n43564, n43565, n43566, n43567, n43568,
    n43569, n43570, n43571, n43572, n43573, n43574,
    n43575, n43576, n43577, n43578, n43579, n43580,
    n43581, n43582, n43583, n43584, n43585, n43586,
    n43587, n43588, n43589, n43590, n43591, n43592,
    n43593, n43594, n43595, n43596, n43597, n43598,
    n43599, n43600, n43601, n43602, n43603, n43604,
    n43605, n43606, n43607, n43608, n43609, n43610,
    n43611, n43612, n43613, n43614, n43615, n43616,
    n43617, n43618, n43619, n43620, n43621, n43622,
    n43623, n43624, n43625, n43626, n43627, n43628,
    n43629, n43630, n43631, n43632, n43633, n43634,
    n43635, n43636, n43637, n43638, n43639, n43640,
    n43641, n43642, n43643, n43644, n43645, n43646,
    n43647, n43648, n43649, n43650, n43651, n43652,
    n43653, n43654, n43655, n43656, n43657, n43658,
    n43659, n43660, n43661, n43662, n43663, n43664,
    n43665, n43666, n43667, n43668, n43669, n43670,
    n43671, n43672, n43673, n43674, n43675, n43676,
    n43677, n43678, n43679, n43680, n43681, n43682,
    n43683, n43684, n43685, n43686, n43687, n43688,
    n43689, n43690, n43691, n43692, n43693, n43694,
    n43695, n43696, n43697, n43698, n43699, n43700,
    n43701, n43702, n43703, n43704, n43705, n43706,
    n43707, n43708, n43709, n43710, n43711, n43712,
    n43713, n43714, n43715, n43716, n43717, n43718,
    n43719, n43720, n43721, n43722, n43723, n43724,
    n43725, n43726, n43727, n43728, n43729, n43730,
    n43731, n43732, n43733, n43734, n43735, n43736,
    n43737, n43738, n43739, n43740, n43741, n43742,
    n43743, n43744, n43745, n43746, n43747, n43748,
    n43749, n43750, n43751, n43752, n43753, n43754,
    n43755, n43756, n43757, n43758, n43759, n43760,
    n43761, n43762, n43763, n43764, n43765, n43766,
    n43767, n43768, n43769, n43770, n43771, n43772,
    n43773, n43774, n43775, n43776, n43777, n43778,
    n43779, n43780, n43781, n43782, n43783, n43784,
    n43785, n43786, n43787, n43788, n43789, n43790,
    n43791, n43792, n43793, n43794, n43795, n43796,
    n43797, n43798, n43799, n43800, n43801, n43802,
    n43803, n43804, n43805, n43806, n43807, n43808,
    n43809, n43810, n43811, n43812, n43813, n43814,
    n43815, n43816, n43817, n43818, n43819, n43820,
    n43821, n43822, n43823, n43824, n43825, n43826,
    n43827, n43828, n43829, n43830, n43831, n43832,
    n43833, n43834, n43835, n43836, n43837, n43838,
    n43839, n43840, n43841, n43842, n43843, n43844,
    n43845, n43846, n43848, n43849, n43850, n43851,
    n43852, n43853, n43855, n43856, n43857, n43858,
    n43859, n43861, n43862, n43863, n43864, n43865,
    n43867, n43868, n43869, n43871, n43872, n43873,
    n43874, n43875, n43877, n43878, n43879, n43881,
    n43882, n43884, n43885, n43886, n43888, n43889,
    n43890, n43891, n43892, n43893, n43894, n43895,
    n43896, n43897, n43898, n43900, n43901, n43902,
    n43903, n43904, n43905, n43906, n43907, n43909,
    n43910, n43911, n43912, n43914, n43915, n43916,
    n43917, n43918, n43919, n43921, n43922, n43924,
    n43925, n43926, n43927, n43928, n43930, n43931,
    n43932, n43934, n43935, n43936, n43938, n43939,
    n43940, n43942, n43943, n43944, n43946, n43947,
    n43948, n43950, n43951, n43952, n43954, n43955,
    n43956, n43958, n43959, n43960, n43961, n43963,
    n43964, n43965, n43966, n43968, n43969, n43970,
    n43971, n43973, n43974, n43975, n43976, n43977,
    n43979, n43980, n43981, n43983, n43984, n43985,
    n43987, n43988, n43989, n43991, n43992, n43993,
    n43995, n43996, n43997, n43999, n44000, n44001,
    n44003, n44004, n44005, n44006, n44007, n44009,
    n44010, n44011, n44012, n44014, n44015, n44016,
    n44018, n44019, n44020, n44022, n44023, n44024,
    n44026, n44027, n44028, n44030, n44031, n44032,
    n44034, n44035, n44036, n44038, n44039, n44040,
    n44042, n44043, n44044, n44046, n44047, n44048,
    n44050, n44051, n44052, n44054, n44055, n44056,
    n44058, n44059, n44060, n44062, n44063, n44064,
    n44066, n44067, n44068, n44070, n44071, n44072,
    n44074, n44075, n44076, n44078, n44079, n44080,
    n44082, n44083, n44084, n44086, n44087, n44088,
    n44090, n44091, n44092, n44094, n44095, n44096,
    n44098, n44099, n44100, n44102, n44103, n44104,
    n44106, n44107, n44108, n44110, n44111, n44112,
    n44114, n44115, n44116, n44118, n44119, n44120,
    n44122, n44123, n44124, n44126, n44127, n44128,
    n44130, n44131, n44132, n44134, n44135, n44136,
    n44138, n44139, n44140, n44142, n44143, n44144,
    n44146, n44147, n44148, n44150, n44151, n44152,
    n44153, n44154, n44155, n44156, n44157, n44158,
    n44160, n44162, n44163, n44164, n44166, n44167,
    n44168, n44170, n44171, n44172, n44174, n44175,
    n44176, n44177, n44178, n44179, n44180, n44181,
    n44182, n44183, n44184, n44185, n44186, n44187,
    n44188, n44189, n44190, n44191, n44192, n44193,
    n44194, n44195, n44196, n44197, n44198, n44199,
    n44200, n44201, n44202, n44203, n44204, n44205,
    n44206, n44207, n44208, n44209, n44210, n44211,
    n44212, n44213, n44214, n44215, n44216, n44217,
    n44218, n44219, n44220, n44222, n44223, n44224,
    n44225, n44226, n44227, n44228, n44229, n44230,
    n44231, n44232, n44233, n44234, n44235, n44236,
    n44237, n44238, n44239, n44240, n44241, n44242,
    n44243, n44244, n44245, n44246, n44247, n44248,
    n44249, n44250, n44251, n44252, n44253, n44254,
    n44255, n44256, n44257, n44258, n44259, n44260,
    n44261, n44262, n44264, n44265, n44266, n44268,
    n44269, n44270, n44271, n44272, n44273, n44274,
    n44275, n44276, n44277, n44278, n44279, n44280,
    n44281, n44282, n44283, n44284, n44285, n44286,
    n44287, n44288, n44289, n44290, n44291, n44292,
    n44293, n44294, n44295, n44296, n44297, n44298,
    n44299, n44300, n44301, n44302, n44304, n44305,
    n44306, n44307, n44308, n44309, n44310, n44311,
    n44312, n44313, n44314, n44315, n44316, n44317,
    n44318, n44319, n44320, n44321, n44322, n44323,
    n44324, n44325, n44326, n44327, n44328, n44329,
    n44330, n44331, n44332, n44333, n44334, n44335,
    n44336, n44337, n44338, n44339, n44341, n44342,
    n44343, n44344, n44345, n44346, n44347, n44348,
    n44349, n44350, n44351, n44352, n44353, n44354,
    n44355, n44356, n44357, n44358, n44359, n44360,
    n44361, n44362, n44363, n44364, n44365, n44366,
    n44367, n44368, n44369, n44370, n44371, n44372,
    n44373, n44374, n44375, n44377, n44378, n44379,
    n44381, n44382, n44383, n44384, n44385, n44386,
    n44387, n44388, n44389, n44390, n44391, n44392,
    n44393, n44394, n44395, n44396, n44397, n44398,
    n44399, n44400, n44401, n44402, n44403, n44404,
    n44405, n44406, n44407, n44408, n44409, n44410,
    n44411, n44412, n44414, n44415, n44416, n44417,
    n44418, n44419, n44420, n44421, n44422, n44423,
    n44424, n44425, n44426, n44427, n44428, n44429,
    n44430, n44431, n44432, n44433, n44434, n44435,
    n44436, n44437, n44438, n44439, n44440, n44441,
    n44442, n44443, n44444, n44446, n44447, n44448,
    n44449, n44450, n44451, n44452, n44453, n44454,
    n44455, n44456, n44457, n44458, n44459, n44460,
    n44461, n44462, n44463, n44464, n44465, n44466,
    n44467, n44468, n44469, n44470, n44471, n44472,
    n44473, n44474, n44475, n44476, n44477, n44478,
    n44479, n44480, n44482, n44483, n44484, n44485,
    n44486, n44487, n44488, n44489, n44490, n44491,
    n44492, n44493, n44494, n44495, n44496, n44497,
    n44498, n44499, n44500, n44501, n44502, n44503,
    n44504, n44505, n44506, n44507, n44508, n44509,
    n44510, n44511, n44512, n44513, n44514, n44515,
    n44516, n44518, n44519, n44520, n44521, n44522,
    n44523, n44524, n44525, n44526, n44527, n44528,
    n44529, n44530, n44531, n44532, n44533, n44534,
    n44535, n44536, n44537, n44538, n44539, n44540,
    n44541, n44542, n44543, n44544, n44545, n44546,
    n44547, n44548, n44549, n44550, n44551, n44552,
    n44553, n44554, n44556, n44557, n44558, n44559,
    n44560, n44561, n44562, n44563, n44564, n44565,
    n44566, n44567, n44568, n44569, n44570, n44571,
    n44572, n44573, n44574, n44575, n44576, n44577,
    n44578, n44579, n44580, n44581, n44582, n44583,
    n44584, n44585, n44586, n44587, n44588, n44589,
    n44590, n44592, n44593, n44594, n44595, n44596,
    n44597, n44598, n44599, n44600, n44601, n44602,
    n44603, n44604, n44605, n44606, n44607, n44608,
    n44609, n44610, n44611, n44612, n44613, n44614,
    n44615, n44616, n44617, n44618, n44619, n44620,
    n44621, n44622, n44623, n44624, n44625, n44626,
    n44628, n44629, n44630, n44631, n44632, n44633,
    n44634, n44635, n44636, n44637, n44638, n44639,
    n44640, n44641, n44642, n44643, n44644, n44645,
    n44646, n44647, n44648, n44649, n44650, n44651,
    n44652, n44653, n44654, n44655, n44656, n44657,
    n44658, n44660, n44661, n44662, n44663, n44664,
    n44665, n44666, n44667, n44668, n44669, n44670,
    n44671, n44672, n44673, n44674, n44675, n44676,
    n44677, n44678, n44679, n44680, n44681, n44682,
    n44683, n44684, n44685, n44686, n44687, n44688,
    n44689, n44690, n44692, n44693, n44694, n44695,
    n44696, n44697, n44698, n44699, n44700, n44701,
    n44702, n44703, n44704, n44705, n44706, n44707,
    n44708, n44709, n44710, n44711, n44712, n44713,
    n44714, n44715, n44716, n44717, n44718, n44719,
    n44720, n44721, n44722, n44723, n44724, n44725,
    n44726, n44727, n44729, n44730, n44731, n44733,
    n44734, n44735, n44737, n44738, n44739, n44740,
    n44741, n44742, n44743, n44744, n44745, n44746,
    n44747, n44748, n44749, n44750, n44751, n44752,
    n44753, n44754, n44755, n44756, n44757, n44758,
    n44759, n44760, n44761, n44762, n44763, n44764,
    n44765, n44766, n44767, n44770, n44771, n44772,
    n44774, n44775, n44776, n44777, n44778, n44779,
    n44780, n44781, n44782, n44783, n44784, n44785,
    n44786, n44787, n44788, n44789, n44790, n44791,
    n44792, n44793, n44794, n44795, n44796, n44797,
    n44798, n44799, n44800, n44801, n44802, n44803,
    n44804, n44805, n44806, n44807, n44808, n44809,
    n44810, n44811, n44813, n44814, n44815, n44817,
    n44818, n44819, n44821, n44822, n44823, n44825,
    n44826, n44827, n44828, n44829, n44830, n44831,
    n44832, n44833, n44834, n44835, n44836, n44837,
    n44838, n44839, n44840, n44841, n44842, n44843,
    n44844, n44845, n44846, n44847, n44848, n44849,
    n44850, n44851, n44852, n44853, n44854, n44855,
    n44856, n44857, n44859, n44860, n44861, n44863,
    n44864, n44865, n44867, n44868, n44869, n44870,
    n44871, n44872, n44873, n44874, n44875, n44876,
    n44877, n44878, n44879, n44880, n44881, n44882,
    n44883, n44884, n44885, n44886, n44887, n44888,
    n44889, n44890, n44891, n44892, n44893, n44894,
    n44895, n44896, n44897, n44898, n44899, n44900,
    n44902, n44903, n44904, n44906, n44907, n44908,
    n44910, n44911, n44912, n44914, n44915, n44916,
    n44918, n44919, n44920, n44922, n44923, n44924,
    n44926, n44927, n44928, n44930, n44931, n44932,
    n44934, n44935, n44936, n44938, n44939, n44940,
    n44942, n44943, n44944, n44946, n44947, n44948,
    n44950, n44951, n44952, n44954, n44955, n44956,
    n44958, n44959, n44960, n44961, n44962, n44963,
    n44964, n44965, n44966, n44967, n44968, n44969,
    n44970, n44971, n44972, n44973, n44974, n44975,
    n44976, n44977, n44978, n44979, n44980, n44981,
    n44982, n44983, n44984, n44985, n44986, n44987,
    n44988, n44989, n44990, n44991, n44992, n44994,
    n44995, n44996, n44997, n44998, n44999, n45000,
    n45001, n45002, n45003, n45004, n45005, n45006,
    n45007, n45008, n45009, n45010, n45011, n45012,
    n45013, n45014, n45015, n45016, n45017, n45018,
    n45019, n45020, n45021, n45022, n45023, n45024,
    n45025, n45026, n45027, n45028, n45029, n45030,
    n45032, n45033, n45034, n45036, n45037, n45038,
    n45040, n45041, n45042, n45043, n45044, n45045,
    n45046, n45047, n45048, n45049, n45050, n45051,
    n45052, n45053, n45054, n45055, n45056, n45057,
    n45058, n45059, n45060, n45061, n45062, n45063,
    n45064, n45065, n45066, n45067, n45068, n45069,
    n45070, n45071, n45072, n45074, n45075, n45076,
    n45077, n45078, n45079, n45080, n45081, n45082,
    n45083, n45084, n45085, n45086, n45087, n45088,
    n45089, n45090, n45091, n45092, n45093, n45094,
    n45095, n45096, n45097, n45098, n45099, n45100,
    n45101, n45102, n45103, n45104, n45105, n45106,
    n45108, n45109, n45110, n45111, n45112, n45113,
    n45114, n45115, n45116, n45117, n45118, n45119,
    n45120, n45121, n45122, n45123, n45124, n45125,
    n45126, n45127, n45128, n45129, n45130, n45131,
    n45132, n45133, n45134, n45135, n45136, n45137,
    n45138, n45139, n45140, n45142, n45143, n45144,
    n45145, n45146, n45147, n45148, n45149, n45150,
    n45151, n45152, n45153, n45154, n45155, n45156,
    n45157, n45158, n45159, n45160, n45161, n45162,
    n45163, n45164, n45165, n45166, n45167, n45168,
    n45169, n45170, n45171, n45172, n45173, n45174,
    n45175, n45177, n45178, n45179, n45181, n45182,
    n45183, n45184, n45185, n45186, n45187, n45188,
    n45189, n45190, n45191, n45192, n45193, n45194,
    n45195, n45196, n45197, n45198, n45199, n45200,
    n45201, n45202, n45203, n45204, n45205, n45206,
    n45207, n45208, n45209, n45210, n45211, n45212,
    n45213, n45214, n45216, n45217, n45218, n45219,
    n45220, n45221, n45222, n45223, n45224, n45225,
    n45226, n45227, n45228, n45229, n45230, n45231,
    n45232, n45233, n45234, n45235, n45236, n45237,
    n45238, n45239, n45240, n45241, n45242, n45243,
    n45244, n45245, n45246, n45247, n45249, n45250,
    n45251, n45252, n45253, n45254, n45255, n45256,
    n45257, n45258, n45259, n45260, n45261, n45262,
    n45263, n45264, n45265, n45266, n45267, n45268,
    n45269, n45270, n45271, n45272, n45273, n45274,
    n45275, n45276, n45277, n45278, n45279, n45280,
    n45281, n45282, n45284, n45285, n45286, n45287,
    n45288, n45289, n45290, n45291, n45292, n45293,
    n45294, n45295, n45296, n45297, n45298, n45299,
    n45300, n45301, n45302, n45303, n45304, n45305,
    n45306, n45307, n45308, n45309, n45310, n45311,
    n45312, n45313, n45314, n45315, n45317, n45318,
    n45319, n45320, n45321, n45322, n45323, n45324,
    n45325, n45326, n45327, n45328, n45329, n45330,
    n45331, n45332, n45333, n45334, n45335, n45336,
    n45337, n45338, n45339, n45340, n45341, n45342,
    n45343, n45344, n45345, n45346, n45347, n45348,
    n45349, n45350, n45352, n45353, n45354, n45355,
    n45356, n45357, n45358, n45359, n45360, n45361,
    n45362, n45363, n45364, n45365, n45366, n45367,
    n45368, n45369, n45370, n45371, n45372, n45373,
    n45374, n45375, n45376, n45377, n45378, n45379,
    n45380, n45381, n45382, n45383, n45384, n45385,
    n45386, n45387, n45388, n45389, n45390, n45391,
    n45392, n45393, n45394, n45395, n45396, n45397,
    n45398, n45399, n45400, n45401, n45402, n45403,
    n45404, n45405, n45407, n45408, n45409, n45411,
    n45412, n45413, n45414, n45415, n45416, n45417,
    n45418, n45419, n45420, n45421, n45422, n45423,
    n45424, n45425, n45426, n45427, n45428, n45429,
    n45430, n45431, n45432, n45433, n45434, n45435,
    n45436, n45437, n45438, n45439, n45440, n45441,
    n45442, n45443, n45444, n45446, n45447, n45448,
    n45450, n45451, n45452, n45454, n45455, n45456,
    n45458, n45459, n45460, n45462, n45463, n45464,
    n45466, n45467, n45468, n45470, n45471, n45472,
    n45474, n45475, n45476, n45478, n45479, n45480,
    n45481, n45482, n45483, n45484, n45485, n45486,
    n45488, n45489, n45490, n45492, n45493, n45494,
    n45495, n45496, n45497, n45498, n45499, n45500,
    n45501, n45502, n45503, n45504, n45505, n45506,
    n45507, n45508, n45509, n45510, n45511, n45512,
    n45513, n45514, n45515, n45516, n45517, n45518,
    n45519, n45520, n45521, n45522, n45523, n45524,
    n45525, n45527, n45528, n45529, n45531, n45532,
    n45533, n45535, n45536, n45537, n45539, n45540,
    n45541, n45543, n45544, n45545, n45547, n45548,
    n45550, n45551, n45552, n45554, n45555, n45556,
    n45558, n45559, n45560, n45562, n45563, n45564,
    n45566, n45567, n45568, n45570, n45571, n45572,
    n45574, n45575, n45576, n45578, n45579, n45580,
    n45581, n45582, n45583, n45584, n45585, n45586,
    n45588, n45589, n45590, n45592, n45593, n45594,
    n45596, n45597, n45598, n45600, n45601, n45602,
    n45604, n45605, n45606, n45608, n45609, n45610,
    n45612, n45613, n45614, n45616, n45617, n45618,
    n45620, n45621, n45622, n45624, n45625, n45626,
    n45628, n45629, n45630, n45632, n45633, n45634,
    n45636, n45637, n45638, n45640, n45641, n45642,
    n45644, n45645, n45646, n45648, n45649, n45650,
    n45652, n45653, n45654, n45656, n45657, n45658,
    n45659, n45660, n45661, n45662, n45663, n45664,
    n45665, n45667, n45668, n45670, n45671, n45672,
    n45674, n45675, n45676, n45678, n45679, n45680,
    n45682, n45683, n45684, n45685, n45686, n45687,
    n45688, n45689, n45690, n45691, n45692, n45693,
    n45694, n45695, n45696, n45698, n45699, n45700,
    n45702, n45703, n45705, n45706, n45707, n45709,
    n45710, n45711, n45712, n45714, n45715, n45716,
    n45718, n45719, n45720, n45721, n45722, n45723,
    n45724, n45725, n45726, n45727, n45728, n45729,
    n45730, n45731, n45732, n45733, n45734, n45736,
    n45737, n45738, n45740, n45741, n45742, n45744,
    n45745, n45746, n45747, n45748, n45749, n45750,
    n45754, n45755, n45757, n45759, n45760, n45762,
    n45763, n45765, n45766, n45768, n45769, n45771,
    n45772, n45774, n45775, n45777, n45778, n45780,
    n45781, n45783, n45784, n45786, n45787, n45789,
    n45790, n45791, n45793, n45794, n45796, n45797,
    n45798, n45799, n45800, n45801, n45802, n45803,
    n45805, n45806, n45808, n45809, n45811, n45812,
    n45814, n45815, n45817, n45818, n45820, n45821,
    n45823, n45824, n45825, n45827, n45828, n45830,
    n45831, n45833, n45834, n45836, n45837, n45839,
    n45840, n45842, n45843, n45845, n45846, n45848,
    n45849, n45851, n45852, n45854, n45855, n45857,
    n45859, n45861, n45863, n45866, n45867, n45868,
    n45870, n45871, n45872, n45873, n45874, n45875,
    n45876, n45877, n45878, n45879, n45880, n45881,
    n45882, n45883, n45884, n45885, n45886, n45887,
    n45888, n45889, n45890, n45891, n45892, n45893,
    n45894, n45895, n45896, n45897, n45899, n45900,
    n45901, n45902, n45903, n45904, n45905, n45906,
    n45907, n45908, n45909, n45910, n45911, n45912,
    n45913, n45914, n45915, n45916, n45917, n45918,
    n45919, n45920, n45921, n45922, n45923, n45924,
    n45925, n45927, n45928, n45929, n45930, n45931,
    n45932, n45933, n45934, n45935, n45936, n45937,
    n45938, n45939, n45940, n45941, n45942, n45943,
    n45944, n45945, n45946, n45947, n45948, n45949,
    n45950, n45951, n45952, n45953, n45955, n45956,
    n45957, n45958, n45959, n45960, n45961, n45962,
    n45963, n45964, n45965, n45966, n45967, n45968,
    n45969, n45970, n45971, n45972, n45973, n45974,
    n45975, n45976, n45977, n45978, n45979, n45980,
    n45981, n45983, n45984, n45986, n45988, n45989,
    n45991, n45992, n45995, n45997, n45998, n46000,
    n46001, n46003, n46004, n46006, n46007, n46010,
    n46011, n46013, n46014, n46016, n46017, n46019,
    n46020, n46022, n46023, n46025, n46026, n46028,
    n46029, n46031, n46032, n46034, n46035, n46037,
    n46038, n46040, n46041, n46043, n46044, n46046,
    n46047, n46049, n46050, n46052, n46053, n46055,
    n46056, n46058, n46059, n46061, n46062, n46064,
    n46065, n46067, n46068, n46069, n46070, n46071,
    n46072, n46073, n46074, n46076, n46077, n46079,
    n46080, n46082, n46083, n46085, n46086, n46088,
    n46089, n46091, n46092, n46094, n46095, n46097,
    n46098, n46099, n46100, n46101, n46102, n46103,
    n46104, n46106, n46107, n46109, n46110, n46112,
    n46113, n46115, n46116, n46118, n46119, n46121,
    n46122, n46123, n46124, n46125, n46126, n46127,
    n46128, n46130, n46131, n46133, n46134, n46135,
    n46136, n46137, n46138, n46139, n46140, n46142,
    n46143, n46144, n46145, n46146, n46147, n46148,
    n46149, n46151, n46152, n46153, n46154, n46155,
    n46156, n46157, n46158, n46160, n46161, n46163,
    n46164, n46166, n46168, n46169, n46171, n46172,
    n46174, n46175, n46177, n46179, n46180, n46182,
    n46183, n46185, n46186, n46188, n46189, n46191,
    n46192, n46194, n46195, n46197, n46198, n46200,
    n46201, n46203, n46204, n46206, n46208, n46209,
    n46211, n46212, n46214, n46215, n46217, n46219,
    n46221, n46222, n46224, n46225, n46226, n46227,
    n46228, n46229, n46230, n46231, n46232, n46233,
    n46235, n46237, n46238, n46240, n46241, n46243,
    n46244, n46246, n46248, n46249, n46251, n46253,
    n46254, n46256, n46258, n46259, n46261, n46262,
    n46264, n46265, n46267, n46268, n46270, n46272,
    n46273, n46275, n46276, n46278, n46280, n46281,
    n46283, n46284, n46286, n46287, n46289, n46291,
    n46292, n46294, n46295, n46297, n46298, n46300,
    n46302, n46304, n46305, n46307, n46309, n46310,
    n46312, n46313, n46315, n46317, n46318, n46320,
    n46322, n46323, n46325, n46326, n46328, n46329,
    n46331, n46332, n46335, n46337, n46339, n46340,
    n46344;
  assign n2437 = ~pi332 & ~pi1144;
  assign n2438 = pi215 & ~n2437;
  assign n2439 = pi265 & ~pi332;
  assign n2440 = pi216 & ~n2439;
  assign n2441 = pi105 & pi228;
  assign n2442 = pi95 & ~pi479;
  assign n2443 = pi234 & n2442;
  assign n2444 = ~pi332 & ~n2443;
  assign n2445 = n2441 & n2444;
  assign n2446 = pi153 & ~pi332;
  assign n2447 = ~n2441 & n2446;
  assign n2448 = ~pi216 & ~n2447;
  assign n2449 = ~n2445 & n2448;
  assign n2450 = ~n2440 & ~n2449;
  assign n2451 = ~pi221 & ~n2450;
  assign n2452 = ~pi216 & pi833;
  assign n2453 = pi1144 & ~n2452;
  assign n2454 = pi929 & n2452;
  assign n2455 = ~pi332 & ~n2453;
  assign n2456 = ~n2454 & n2455;
  assign n2457 = pi221 & ~n2456;
  assign n2458 = ~n2451 & ~n2457;
  assign n2459 = ~pi215 & ~n2458;
  assign n2460 = ~n2438 & ~n2459;
  assign n2461 = ~pi215 & ~pi221;
  assign n2462 = ~pi32 & ~pi40;
  assign n2463 = ~pi58 & ~pi90;
  assign n2464 = ~pi88 & ~pi98;
  assign n2465 = ~pi77 & n2464;
  assign n2466 = ~pi50 & n2465;
  assign n2467 = ~pi102 & n2466;
  assign n2468 = ~pi65 & ~pi71;
  assign n2469 = ~pi61 & ~pi76;
  assign n2470 = ~pi85 & ~pi106;
  assign n2471 = n2469 & n2470;
  assign n2472 = ~pi48 & n2471;
  assign n2473 = ~pi89 & n2472;
  assign n2474 = ~pi49 & n2473;
  assign n2475 = ~pi104 & n2474;
  assign n2476 = ~pi45 & n2475;
  assign n2477 = ~pi68 & ~pi84;
  assign n2478 = ~pi82 & ~pi111;
  assign n2479 = ~pi36 & n2478;
  assign n2480 = n2477 & n2479;
  assign n2481 = ~pi66 & ~pi73;
  assign n2482 = n2480 & n2481;
  assign n2483 = n2476 & n2482;
  assign n2484 = ~pi69 & ~pi83;
  assign n2485 = ~pi67 & ~pi103;
  assign n2486 = n2484 & n2485;
  assign n2487 = n2483 & n2486;
  assign n2488 = n2468 & n2487;
  assign n2489 = ~pi63 & ~pi107;
  assign n2490 = n2488 & n2489;
  assign n2491 = ~pi64 & n2490;
  assign n2492 = ~pi81 & n2491;
  assign n2493 = n2467 & n2492;
  assign n2494 = ~pi53 & ~pi60;
  assign n2495 = ~pi86 & n2494;
  assign n2496 = ~pi109 & ~pi110;
  assign n2497 = ~pi46 & ~pi97;
  assign n2498 = ~pi108 & n2497;
  assign n2499 = n2496 & n2498;
  assign n2500 = ~pi94 & n2499;
  assign n2501 = n2495 & n2500;
  assign n2502 = ~pi47 & ~pi91;
  assign n2503 = n2501 & n2502;
  assign n2504 = n2493 & n2503;
  assign n2505 = n2463 & n2504;
  assign n2506 = ~pi93 & n2505;
  assign n2507 = ~pi72 & ~pi96;
  assign n2508 = ~pi35 & ~pi70;
  assign n2509 = ~pi51 & n2508;
  assign n2510 = n2507 & n2509;
  assign n2511 = n2506 & n2510;
  assign n2512 = n2462 & n2511;
  assign n2513 = ~pi95 & n2512;
  assign n2514 = ~n2442 & ~n2513;
  assign n2515 = pi234 & ~n2514;
  assign n2516 = ~pi35 & ~pi93;
  assign n2517 = n2505 & n2516;
  assign n2518 = ~pi32 & ~pi95;
  assign n2519 = ~pi51 & ~pi70;
  assign n2520 = n2507 & n2519;
  assign n2521 = ~pi40 & n2520;
  assign n2522 = n2518 & n2521;
  assign n2523 = n2517 & n2522;
  assign n2524 = ~pi234 & n2523;
  assign n2525 = ~n2515 & ~n2524;
  assign n2526 = pi137 & ~n2525;
  assign n2527 = n2444 & ~n2526;
  assign n2528 = n2448 & n2461;
  assign n2529 = ~n2527 & n2528;
  assign n2530 = ~pi56 & ~pi62;
  assign n2531 = ~pi38 & ~pi39;
  assign n2532 = ~pi100 & n2531;
  assign n2533 = ~pi54 & ~pi74;
  assign n2534 = ~pi75 & ~pi87;
  assign n2535 = ~pi92 & n2534;
  assign n2536 = n2533 & n2535;
  assign n2537 = ~pi55 & n2536;
  assign n2538 = n2532 & n2537;
  assign n2539 = n2530 & n2538;
  assign n2540 = n2529 & n2539;
  assign n2541 = ~pi59 & n2540;
  assign n2542 = n2460 & ~n2541;
  assign n2543 = pi57 & ~n2542;
  assign n2544 = pi59 & n2460;
  assign n2545 = ~n2540 & n2544;
  assign n2546 = n2460 & ~n2538;
  assign n2547 = ~pi105 & ~n2446;
  assign n2548 = pi105 & ~n2527;
  assign n2549 = ~n2547 & ~n2548;
  assign n2550 = pi228 & ~n2549;
  assign n2551 = ~pi137 & ~pi153;
  assign n2552 = ~pi332 & n2551;
  assign n2553 = n2513 & n2552;
  assign n2554 = pi137 & n2523;
  assign n2555 = n2446 & ~n2554;
  assign n2556 = ~pi228 & ~n2555;
  assign n2557 = ~n2553 & n2556;
  assign n2558 = ~n2550 & ~n2557;
  assign n2559 = ~pi216 & ~n2558;
  assign n2560 = ~n2440 & ~n2559;
  assign n2561 = ~pi221 & ~n2560;
  assign n2562 = ~n2457 & ~n2561;
  assign n2563 = ~pi215 & ~n2562;
  assign n2564 = ~n2438 & ~n2563;
  assign n2565 = n2538 & n2564;
  assign n2566 = ~n2546 & ~n2565;
  assign n2567 = ~pi56 & ~n2566;
  assign n2568 = pi56 & n2460;
  assign n2569 = pi62 & ~n2568;
  assign n2570 = ~n2567 & n2569;
  assign n2571 = pi56 & ~n2566;
  assign n2572 = ~pi75 & ~pi92;
  assign n2573 = ~pi87 & ~pi100;
  assign n2574 = ~pi38 & n2573;
  assign n2575 = n2572 & n2574;
  assign n2576 = n2533 & n2575;
  assign n2577 = ~pi39 & n2576;
  assign n2578 = n2460 & ~n2577;
  assign n2579 = pi228 & ~n2547;
  assign n2580 = ~pi332 & n2525;
  assign n2581 = pi105 & ~n2580;
  assign n2582 = n2579 & ~n2581;
  assign n2583 = ~pi228 & n2446;
  assign n2584 = ~n2523 & n2583;
  assign n2585 = ~pi216 & ~n2584;
  assign n2586 = ~n2582 & n2585;
  assign n2587 = ~n2440 & ~n2586;
  assign n2588 = ~pi221 & ~n2587;
  assign n2589 = ~n2457 & ~n2588;
  assign n2590 = ~pi215 & ~n2589;
  assign n2591 = ~n2438 & n2577;
  assign n2592 = ~n2590 & n2591;
  assign n2593 = pi55 & ~n2578;
  assign n2594 = ~n2592 & n2593;
  assign n2595 = pi299 & n2460;
  assign n2596 = ~pi224 & pi833;
  assign n2597 = pi222 & ~n2596;
  assign n2598 = ~pi223 & ~n2597;
  assign n2599 = n2437 & ~n2598;
  assign n2600 = pi224 & ~n2439;
  assign n2601 = ~pi222 & ~n2600;
  assign n2602 = ~pi332 & ~pi929;
  assign n2603 = n2596 & n2602;
  assign n2604 = ~n2601 & ~n2603;
  assign n2605 = ~pi223 & ~n2604;
  assign n2606 = ~n2599 & ~n2605;
  assign n2607 = ~pi299 & ~n2606;
  assign n2608 = ~pi222 & ~pi224;
  assign n2609 = ~pi223 & n2608;
  assign n2610 = ~n2444 & n2609;
  assign n2611 = n2607 & ~n2610;
  assign n2612 = ~n2595 & ~n2611;
  assign n2613 = ~pi38 & ~pi100;
  assign n2614 = ~pi39 & ~pi87;
  assign n2615 = n2613 & n2614;
  assign n2616 = n2572 & n2615;
  assign n2617 = n2612 & ~n2616;
  assign n2618 = ~n2527 & n2609;
  assign n2619 = ~n2606 & ~n2618;
  assign n2620 = ~pi299 & ~n2619;
  assign n2621 = n2460 & ~n2529;
  assign n2622 = pi299 & ~n2621;
  assign n2623 = ~n2620 & ~n2622;
  assign n2624 = ~pi39 & ~n2623;
  assign n2625 = n2575 & n2624;
  assign n2626 = ~n2617 & ~n2625;
  assign n2627 = pi54 & n2626;
  assign n2628 = ~pi39 & n2613;
  assign n2629 = ~n2612 & ~n2628;
  assign n2630 = pi299 & ~n2564;
  assign n2631 = ~n2620 & ~n2630;
  assign n2632 = n2628 & n2631;
  assign n2633 = ~n2629 & ~n2632;
  assign n2634 = n2534 & ~n2633;
  assign n2635 = ~n2534 & ~n2612;
  assign n2636 = pi92 & ~n2635;
  assign n2637 = ~n2634 & n2636;
  assign n2638 = pi87 & ~n2633;
  assign n2639 = ~n2531 & ~n2612;
  assign n2640 = ~pi144 & ~pi174;
  assign n2641 = ~pi189 & n2640;
  assign n2642 = ~pi223 & ~n2641;
  assign n2643 = pi142 & ~pi198;
  assign n2644 = ~pi137 & ~n2643;
  assign n2645 = ~n2525 & ~n2644;
  assign n2646 = n2444 & ~n2645;
  assign n2647 = n2642 & ~n2646;
  assign n2648 = ~pi234 & ~pi332;
  assign n2649 = ~pi137 & pi198;
  assign n2650 = n2523 & ~n2649;
  assign n2651 = n2648 & ~n2650;
  assign n2652 = ~pi223 & n2641;
  assign n2653 = pi234 & ~pi332;
  assign n2654 = ~pi95 & n2649;
  assign n2655 = ~n2514 & ~n2654;
  assign n2656 = n2653 & ~n2655;
  assign n2657 = ~n2651 & n2652;
  assign n2658 = ~n2656 & n2657;
  assign n2659 = ~n2647 & ~n2658;
  assign n2660 = n2608 & ~n2659;
  assign n2661 = ~n2606 & ~n2660;
  assign n2662 = ~pi299 & ~n2661;
  assign n2663 = pi95 & pi234;
  assign n2664 = ~pi152 & ~pi161;
  assign n2665 = ~pi166 & n2664;
  assign n2666 = ~pi146 & ~n2665;
  assign n2667 = ~pi210 & ~n2666;
  assign n2668 = ~pi137 & ~n2667;
  assign n2669 = ~n2663 & n2668;
  assign n2670 = ~n2525 & ~n2669;
  assign n2671 = ~pi332 & ~n2670;
  assign n2672 = pi105 & ~n2671;
  assign n2673 = n2579 & ~n2672;
  assign n2674 = n2554 & n2666;
  assign n2675 = ~pi252 & ~n2666;
  assign n2676 = n2513 & n2675;
  assign n2677 = pi153 & ~n2674;
  assign n2678 = ~n2676 & n2677;
  assign n2679 = pi252 & ~n2666;
  assign n2680 = n2668 & ~n2679;
  assign n2681 = n2513 & n2680;
  assign n2682 = ~n2678 & ~n2681;
  assign n2683 = ~pi228 & ~pi332;
  assign n2684 = ~n2682 & n2683;
  assign n2685 = ~pi216 & ~n2684;
  assign n2686 = ~n2673 & n2685;
  assign n2687 = ~n2440 & ~n2686;
  assign n2688 = ~pi221 & ~n2687;
  assign n2689 = ~n2457 & ~n2688;
  assign n2690 = ~pi215 & ~n2689;
  assign n2691 = ~n2438 & ~n2690;
  assign n2692 = pi299 & ~n2691;
  assign n2693 = n2531 & ~n2662;
  assign n2694 = ~n2692 & n2693;
  assign n2695 = pi100 & ~n2639;
  assign n2696 = ~n2694 & n2695;
  assign n2697 = pi39 & n2612;
  assign n2698 = pi38 & ~n2697;
  assign n2699 = ~n2624 & n2698;
  assign n2700 = pi39 & ~n2631;
  assign n2701 = ~pi40 & ~pi72;
  assign n2702 = ~pi94 & n2498;
  assign n2703 = n2495 & n2702;
  assign n2704 = n2493 & n2703;
  assign n2705 = ~pi58 & ~pi91;
  assign n2706 = ~pi47 & n2705;
  assign n2707 = n2496 & n2706;
  assign n2708 = n2704 & n2707;
  assign n2709 = ~pi90 & ~pi93;
  assign n2710 = ~pi96 & n2509;
  assign n2711 = n2709 & n2710;
  assign n2712 = n2708 & n2711;
  assign n2713 = n2701 & n2712;
  assign n2714 = pi225 & n2713;
  assign n2715 = pi32 & ~n2714;
  assign n2716 = ~pi95 & ~n2715;
  assign n2717 = n2498 & n2707;
  assign n2718 = pi60 & n2493;
  assign n2719 = ~pi53 & ~n2718;
  assign n2720 = ~pi86 & ~pi94;
  assign n2721 = ~pi60 & n2493;
  assign n2722 = pi53 & ~n2721;
  assign n2723 = n2720 & ~n2722;
  assign n2724 = ~n2719 & n2723;
  assign n2725 = n2709 & n2717;
  assign n2726 = n2724 & n2725;
  assign n2727 = ~pi35 & ~n2726;
  assign n2728 = pi35 & ~n2506;
  assign n2729 = pi35 & n2506;
  assign n2730 = ~pi225 & n2729;
  assign n2731 = ~pi70 & ~n2730;
  assign n2732 = ~pi51 & n2731;
  assign n2733 = ~n2728 & n2732;
  assign n2734 = ~n2727 & n2733;
  assign n2735 = ~pi40 & n2507;
  assign n2736 = n2734 & n2735;
  assign n2737 = ~pi32 & ~n2736;
  assign n2738 = n2716 & ~n2737;
  assign n2739 = ~pi137 & ~n2738;
  assign n2740 = pi95 & ~n2512;
  assign n2741 = ~n2442 & ~n2740;
  assign n2742 = pi40 & n2511;
  assign n2743 = ~pi32 & ~n2742;
  assign n2744 = pi72 & ~n2712;
  assign n2745 = ~pi40 & ~n2744;
  assign n2746 = ~pi70 & n2517;
  assign n2747 = pi51 & ~n2746;
  assign n2748 = ~pi96 & ~n2747;
  assign n2749 = ~pi51 & pi70;
  assign n2750 = n2748 & ~n2749;
  assign n2751 = ~n2728 & ~n2730;
  assign n2752 = pi93 & n2505;
  assign n2753 = ~pi35 & ~n2752;
  assign n2754 = ~pi47 & n2501;
  assign n2755 = n2493 & n2754;
  assign n2756 = pi91 & n2755;
  assign n2757 = n2463 & ~n2756;
  assign n2758 = ~pi109 & n2704;
  assign n2759 = pi110 & ~n2758;
  assign n2760 = pi47 & n2493;
  assign n2761 = n2501 & n2760;
  assign n2762 = pi47 & ~n2761;
  assign n2763 = ~pi91 & ~n2759;
  assign n2764 = ~n2762 & n2763;
  assign n2765 = ~pi47 & ~pi110;
  assign n2766 = pi109 & ~n2704;
  assign n2767 = ~pi50 & n2494;
  assign n2768 = ~pi102 & n2492;
  assign n2769 = n2465 & n2768;
  assign n2770 = n2767 & n2769;
  assign n2771 = n2720 & n2770;
  assign n2772 = ~pi97 & n2771;
  assign n2773 = pi108 & ~n2772;
  assign n2774 = ~pi46 & ~n2773;
  assign n2775 = pi97 & ~n2771;
  assign n2776 = ~pi86 & pi94;
  assign n2777 = n2770 & n2776;
  assign n2778 = ~pi97 & ~n2777;
  assign n2779 = pi86 & ~n2770;
  assign n2780 = ~pi94 & ~n2779;
  assign n2781 = pi77 & n2464;
  assign n2782 = n2768 & n2781;
  assign n2783 = ~pi50 & ~n2782;
  assign n2784 = pi81 & ~n2491;
  assign n2785 = pi102 & ~n2492;
  assign n2786 = ~n2784 & ~n2785;
  assign n2787 = pi64 & ~n2490;
  assign n2788 = pi71 & ~n2487;
  assign n2789 = ~pi65 & ~n2788;
  assign n2790 = ~pi67 & n2483;
  assign n2791 = pi69 & ~n2790;
  assign n2792 = ~pi67 & ~pi69;
  assign n2793 = n2483 & n2792;
  assign n2794 = pi83 & ~n2793;
  assign n2795 = ~pi103 & ~n2794;
  assign n2796 = ~n2791 & n2795;
  assign n2797 = pi67 & ~n2483;
  assign n2798 = n2476 & n2481;
  assign n2799 = ~pi84 & n2798;
  assign n2800 = ~pi68 & n2799;
  assign n2801 = n2478 & n2800;
  assign n2802 = pi36 & ~n2801;
  assign n2803 = ~pi36 & ~pi67;
  assign n2804 = ~pi68 & ~pi111;
  assign n2805 = pi82 & n2804;
  assign n2806 = n2799 & n2805;
  assign n2807 = pi111 & ~n2800;
  assign n2808 = ~pi82 & ~n2807;
  assign n2809 = pi84 & ~n2798;
  assign n2810 = pi104 & ~n2474;
  assign n2811 = pi85 & pi106;
  assign n2812 = n2469 & ~n2811;
  assign n2813 = pi61 & pi76;
  assign n2814 = n2470 & ~n2813;
  assign n2815 = ~n2812 & ~n2814;
  assign n2816 = ~pi48 & ~n2815;
  assign n2817 = ~n2471 & ~n2816;
  assign n2818 = pi89 & ~n2472;
  assign n2819 = ~pi49 & ~n2818;
  assign n2820 = ~n2817 & n2819;
  assign n2821 = ~n2473 & ~n2820;
  assign n2822 = ~pi45 & ~n2810;
  assign n2823 = ~n2821 & n2822;
  assign n2824 = ~n2475 & ~n2823;
  assign n2825 = ~n2476 & ~n2824;
  assign n2826 = n2481 & ~n2825;
  assign n2827 = pi66 & pi73;
  assign n2828 = ~n2476 & ~n2481;
  assign n2829 = ~n2827 & ~n2828;
  assign n2830 = ~n2826 & n2829;
  assign n2831 = ~pi84 & ~n2830;
  assign n2832 = ~n2809 & ~n2831;
  assign n2833 = n2804 & ~n2832;
  assign n2834 = pi68 & ~n2799;
  assign n2835 = n2808 & ~n2834;
  assign n2836 = ~n2833 & n2835;
  assign n2837 = n2803 & ~n2806;
  assign n2838 = ~n2836 & n2837;
  assign n2839 = ~n2797 & ~n2802;
  assign n2840 = ~n2838 & n2839;
  assign n2841 = n2484 & ~n2840;
  assign n2842 = n2796 & ~n2841;
  assign n2843 = ~pi83 & pi103;
  assign n2844 = n2793 & n2843;
  assign n2845 = ~pi71 & ~n2844;
  assign n2846 = ~n2842 & n2845;
  assign n2847 = n2789 & ~n2846;
  assign n2848 = ~pi107 & ~n2847;
  assign n2849 = ~pi63 & pi107;
  assign n2850 = n2488 & n2849;
  assign n2851 = ~n2489 & ~n2850;
  assign n2852 = ~n2848 & ~n2851;
  assign n2853 = pi65 & ~pi71;
  assign n2854 = n2487 & n2853;
  assign n2855 = ~n2851 & n2854;
  assign n2856 = ~pi64 & ~n2855;
  assign n2857 = ~n2852 & n2856;
  assign n2858 = ~n2787 & ~n2857;
  assign n2859 = ~pi81 & ~pi102;
  assign n2860 = ~n2858 & n2859;
  assign n2861 = pi63 & ~pi107;
  assign n2862 = n2488 & n2861;
  assign n2863 = ~pi64 & ~n2862;
  assign n2864 = ~n2852 & n2863;
  assign n2865 = ~n2787 & ~n2864;
  assign n2866 = n2860 & ~n2865;
  assign n2867 = n2786 & ~n2866;
  assign n2868 = n2464 & ~n2867;
  assign n2869 = pi98 & ~n2768;
  assign n2870 = ~pi98 & n2768;
  assign n2871 = pi88 & ~n2870;
  assign n2872 = ~pi77 & ~n2869;
  assign n2873 = ~n2871 & n2872;
  assign n2874 = ~n2868 & n2873;
  assign n2875 = n2783 & ~n2874;
  assign n2876 = pi50 & ~n2769;
  assign n2877 = ~pi60 & ~n2876;
  assign n2878 = ~n2875 & n2877;
  assign n2879 = n2719 & ~n2878;
  assign n2880 = ~n2722 & ~n2879;
  assign n2881 = ~pi86 & ~n2880;
  assign n2882 = n2780 & ~n2881;
  assign n2883 = n2778 & ~n2882;
  assign n2884 = ~n2775 & ~n2883;
  assign n2885 = ~pi108 & ~n2884;
  assign n2886 = n2774 & ~n2885;
  assign n2887 = ~pi108 & n2771;
  assign n2888 = pi46 & ~pi97;
  assign n2889 = n2887 & n2888;
  assign n2890 = ~pi109 & ~n2889;
  assign n2891 = ~n2886 & n2890;
  assign n2892 = ~n2766 & ~n2891;
  assign n2893 = n2765 & ~n2892;
  assign n2894 = n2764 & ~n2893;
  assign n2895 = n2757 & ~n2894;
  assign n2896 = pi58 & ~n2504;
  assign n2897 = pi90 & ~n2708;
  assign n2898 = ~pi93 & ~n2897;
  assign n2899 = ~n2896 & n2898;
  assign n2900 = ~n2895 & n2899;
  assign n2901 = n2753 & ~n2900;
  assign n2902 = n2751 & ~n2901;
  assign n2903 = ~pi51 & ~n2902;
  assign n2904 = n2750 & ~n2903;
  assign n2905 = ~pi72 & ~n2904;
  assign n2906 = n2745 & ~n2905;
  assign n2907 = n2743 & ~n2906;
  assign n2908 = ~n2715 & ~n2907;
  assign n2909 = ~pi95 & ~n2908;
  assign n2910 = n2741 & ~n2909;
  assign n2911 = pi137 & ~n2910;
  assign n2912 = ~n2739 & ~n2911;
  assign n2913 = pi210 & ~n2912;
  assign n2914 = pi841 & n2505;
  assign n2915 = ~pi93 & n2914;
  assign n2916 = ~pi35 & n2521;
  assign n2917 = n2915 & n2916;
  assign n2918 = pi225 & n2917;
  assign n2919 = pi32 & ~n2918;
  assign n2920 = ~pi95 & ~n2919;
  assign n2921 = ~pi833 & pi957;
  assign n2922 = pi1091 & ~n2921;
  assign n2923 = pi1092 & pi1093;
  assign n2924 = pi829 & pi950;
  assign n2925 = n2923 & n2924;
  assign n2926 = n2922 & n2925;
  assign n2927 = ~pi46 & ~pi109;
  assign n2928 = n2502 & n2927;
  assign n2929 = ~pi108 & ~n2775;
  assign n2930 = ~pi110 & n2929;
  assign n2931 = ~pi93 & n2463;
  assign n2932 = ~pi97 & ~n2724;
  assign n2933 = n2928 & n2931;
  assign n2934 = ~n2932 & n2933;
  assign n2935 = n2930 & n2934;
  assign n2936 = ~pi35 & ~n2935;
  assign n2937 = n2926 & n2936;
  assign n2938 = n2727 & ~n2926;
  assign n2939 = n2521 & n2751;
  assign n2940 = ~n2938 & n2939;
  assign n2941 = ~n2937 & n2940;
  assign n2942 = ~pi32 & ~n2941;
  assign n2943 = n2920 & ~n2942;
  assign n2944 = ~pi137 & ~n2943;
  assign n2945 = ~n2907 & ~n2919;
  assign n2946 = ~pi95 & ~n2945;
  assign n2947 = n2741 & ~n2946;
  assign n2948 = pi137 & ~n2947;
  assign n2949 = ~n2944 & ~n2948;
  assign n2950 = ~pi210 & ~n2949;
  assign n2951 = ~n2913 & ~n2950;
  assign n2952 = ~pi234 & n2951;
  assign n2953 = ~pi96 & ~n2734;
  assign n2954 = ~pi91 & n2509;
  assign n2955 = n2931 & n2954;
  assign n2956 = n2755 & n2955;
  assign n2957 = pi96 & ~n2956;
  assign n2958 = n2701 & ~n2957;
  assign n2959 = ~n2953 & n2958;
  assign n2960 = ~pi32 & ~n2959;
  assign n2961 = n2716 & ~n2960;
  assign n2962 = ~n2442 & ~n2961;
  assign n2963 = ~pi137 & n2962;
  assign n2964 = pi96 & n2956;
  assign n2965 = ~pi51 & n2506;
  assign n2966 = ~pi35 & n2965;
  assign n2967 = n2701 & n2966;
  assign n2968 = n2964 & n2967;
  assign n2969 = n2907 & ~n2968;
  assign n2970 = ~n2715 & ~n2969;
  assign n2971 = ~pi95 & ~n2970;
  assign n2972 = pi479 & n2740;
  assign n2973 = ~n2971 & ~n2972;
  assign n2974 = pi137 & ~n2973;
  assign n2975 = ~n2963 & ~n2974;
  assign n2976 = pi210 & ~n2975;
  assign n2977 = ~n2919 & ~n2969;
  assign n2978 = ~pi95 & ~n2977;
  assign n2979 = ~n2972 & ~n2978;
  assign n2980 = pi137 & ~n2979;
  assign n2981 = n2733 & ~n2936;
  assign n2982 = ~pi96 & ~n2981;
  assign n2983 = n2958 & ~n2982;
  assign n2984 = ~pi32 & ~n2983;
  assign n2985 = n2920 & ~n2984;
  assign n2986 = ~n2442 & ~n2985;
  assign n2987 = n2926 & ~n2986;
  assign n2988 = n2920 & ~n2960;
  assign n2989 = ~n2442 & ~n2988;
  assign n2990 = ~n2926 & ~n2989;
  assign n2991 = ~pi137 & ~n2990;
  assign n2992 = ~n2987 & n2991;
  assign n2993 = ~n2980 & ~n2992;
  assign n2994 = ~pi210 & ~n2993;
  assign n2995 = ~n2976 & ~n2994;
  assign n2996 = pi234 & n2995;
  assign n2997 = n2665 & ~n2952;
  assign n2998 = ~n2996 & n2997;
  assign n2999 = ~n2666 & n2995;
  assign n3000 = ~pi137 & n2989;
  assign n3001 = ~n2980 & ~n3000;
  assign n3002 = ~pi210 & ~n3001;
  assign n3003 = ~pi146 & ~n2976;
  assign n3004 = ~n3002 & n3003;
  assign n3005 = pi234 & ~n2999;
  assign n3006 = ~n3004 & n3005;
  assign n3007 = ~n2998 & ~n3006;
  assign n3008 = ~pi332 & ~n3007;
  assign n3009 = pi146 & n2951;
  assign n3010 = ~n2737 & n2920;
  assign n3011 = ~pi137 & ~n3010;
  assign n3012 = ~n2948 & ~n3011;
  assign n3013 = ~pi210 & ~n3012;
  assign n3014 = ~pi146 & ~n2913;
  assign n3015 = ~n3013 & n3014;
  assign n3016 = n2648 & ~n2665;
  assign n3017 = ~n3009 & n3016;
  assign n3018 = ~n3015 & n3017;
  assign n3019 = pi105 & ~n3018;
  assign n3020 = ~n3008 & n3019;
  assign n3021 = n2579 & ~n3020;
  assign n3022 = ~pi109 & ~n2886;
  assign n3023 = ~n2766 & ~n3022;
  assign n3024 = n2765 & ~n3023;
  assign n3025 = n2764 & ~n3024;
  assign n3026 = n2757 & ~n3025;
  assign n3027 = n2899 & ~n3026;
  assign n3028 = n2753 & ~n3027;
  assign n3029 = n2751 & ~n3028;
  assign n3030 = ~pi51 & ~n3029;
  assign n3031 = n2750 & ~n3030;
  assign n3032 = ~pi72 & ~n3031;
  assign n3033 = n2745 & ~n3032;
  assign n3034 = n2743 & ~n3033;
  assign n3035 = ~n2919 & ~n3034;
  assign n3036 = ~pi95 & ~n3035;
  assign n3037 = n2741 & ~n3036;
  assign n3038 = pi137 & ~n3037;
  assign n3039 = n2666 & n3011;
  assign n3040 = ~n2666 & n2944;
  assign n3041 = ~pi210 & ~pi234;
  assign n3042 = ~n3039 & n3041;
  assign n3043 = ~n3040 & n3042;
  assign n3044 = ~n3038 & n3043;
  assign n3045 = ~n2715 & ~n3034;
  assign n3046 = ~pi95 & ~n3045;
  assign n3047 = n2741 & ~n3046;
  assign n3048 = pi137 & ~n3047;
  assign n3049 = pi210 & ~n2739;
  assign n3050 = ~n3048 & n3049;
  assign n3051 = ~pi95 & pi137;
  assign n3052 = ~n2968 & n3034;
  assign n3053 = ~n2919 & ~n3052;
  assign n3054 = n3051 & ~n3053;
  assign n3055 = ~n2666 & n2987;
  assign n3056 = n2666 & ~n2989;
  assign n3057 = n2991 & ~n3056;
  assign n3058 = ~n3055 & n3057;
  assign n3059 = ~n2740 & ~n3058;
  assign n3060 = ~n3054 & n3059;
  assign n3061 = ~pi210 & ~n3060;
  assign n3062 = pi234 & ~n3061;
  assign n3063 = ~n3044 & ~n3050;
  assign n3064 = ~n3062 & n3063;
  assign n3065 = ~pi137 & ~n2740;
  assign n3066 = ~n2962 & n3065;
  assign n3067 = ~n2715 & ~n3052;
  assign n3068 = ~pi95 & ~n3067;
  assign n3069 = pi137 & ~n2740;
  assign n3070 = ~n3068 & n3069;
  assign n3071 = pi210 & pi234;
  assign n3072 = ~n3066 & n3071;
  assign n3073 = ~n3070 & n3072;
  assign n3074 = ~n3064 & ~n3073;
  assign n3075 = n2446 & ~n3074;
  assign n3076 = pi225 & pi841;
  assign n3077 = n2713 & ~n3076;
  assign n3078 = pi32 & ~n3077;
  assign n3079 = ~pi95 & ~n3078;
  assign n3080 = ~pi51 & ~pi96;
  assign n3081 = pi70 & ~n2517;
  assign n3082 = n3080 & ~n3081;
  assign n3083 = n2701 & n3082;
  assign n3084 = ~n2731 & n3083;
  assign n3085 = ~pi32 & ~n3084;
  assign n3086 = n3079 & ~n3085;
  assign n3087 = pi137 & ~n3086;
  assign n3088 = pi93 & ~n2505;
  assign n3089 = ~pi35 & ~n3088;
  assign n3090 = ~n2896 & ~n2897;
  assign n3091 = ~pi53 & n2878;
  assign n3092 = ~pi86 & ~n3091;
  assign n3093 = n2780 & ~n3092;
  assign n3094 = n2778 & ~n3093;
  assign n3095 = ~n2775 & ~n3094;
  assign n3096 = ~pi108 & ~n3095;
  assign n3097 = n2774 & ~n3096;
  assign n3098 = ~pi109 & ~n3097;
  assign n3099 = ~n2766 & ~n3098;
  assign n3100 = n2765 & ~n3099;
  assign n3101 = n2764 & ~n3100;
  assign n3102 = n2757 & ~n3101;
  assign n3103 = n3090 & ~n3102;
  assign n3104 = ~pi93 & ~n3103;
  assign n3105 = n3089 & ~n3104;
  assign n3106 = n2732 & ~n3105;
  assign n3107 = n2748 & ~n3081;
  assign n3108 = ~n3106 & n3107;
  assign n3109 = ~pi72 & ~n3108;
  assign n3110 = n2745 & ~n3109;
  assign n3111 = n2743 & ~n3110;
  assign n3112 = ~n2926 & n3111;
  assign n3113 = n2743 & n2926;
  assign n3114 = ~pi97 & ~n3094;
  assign n3115 = ~pi108 & ~n3114;
  assign n3116 = n2774 & ~n3115;
  assign n3117 = ~pi109 & ~n3116;
  assign n3118 = ~n2766 & ~n3117;
  assign n3119 = n2765 & ~n3118;
  assign n3120 = n2764 & ~n3119;
  assign n3121 = n2757 & ~n3120;
  assign n3122 = n3090 & ~n3121;
  assign n3123 = ~pi93 & ~n3122;
  assign n3124 = n3089 & ~n3123;
  assign n3125 = n2732 & ~n3124;
  assign n3126 = n3107 & ~n3125;
  assign n3127 = ~pi72 & ~n3126;
  assign n3128 = n2745 & ~n3127;
  assign n3129 = n3113 & ~n3128;
  assign n3130 = ~n3078 & ~n3129;
  assign n3131 = ~n3112 & n3130;
  assign n3132 = ~pi95 & ~n3131;
  assign n3133 = n2741 & ~n3132;
  assign n3134 = ~pi137 & ~n3133;
  assign n3135 = ~n3087 & ~n3134;
  assign n3136 = ~pi210 & ~n3135;
  assign n3137 = ~pi225 & n2713;
  assign n3138 = pi32 & ~n3137;
  assign n3139 = ~n3111 & ~n3138;
  assign n3140 = ~pi95 & ~n3139;
  assign n3141 = ~pi137 & n2741;
  assign n3142 = ~n3140 & n3141;
  assign n3143 = ~n3085 & ~n3138;
  assign n3144 = n3051 & n3143;
  assign n3145 = pi210 & ~n3144;
  assign n3146 = ~n3142 & n3145;
  assign n3147 = n2653 & ~n3146;
  assign n3148 = ~n3136 & n3147;
  assign n3149 = ~pi72 & ~n2964;
  assign n3150 = ~n3108 & n3149;
  assign n3151 = n2745 & ~n3150;
  assign n3152 = n2743 & ~n3151;
  assign n3153 = ~n2926 & n3152;
  assign n3154 = ~n3126 & n3149;
  assign n3155 = n2745 & ~n3154;
  assign n3156 = n3113 & ~n3155;
  assign n3157 = ~n3078 & ~n3156;
  assign n3158 = ~n3153 & n3157;
  assign n3159 = ~pi95 & ~n3158;
  assign n3160 = ~n2740 & ~n3159;
  assign n3161 = ~pi137 & ~n3160;
  assign n3162 = n2442 & n2512;
  assign n3163 = ~pi72 & n2462;
  assign n3164 = n2964 & n3163;
  assign n3165 = n3085 & ~n3164;
  assign n3166 = n3079 & ~n3165;
  assign n3167 = pi137 & ~n3162;
  assign n3168 = ~n3166 & n3167;
  assign n3169 = ~n3161 & ~n3168;
  assign n3170 = ~pi210 & ~n3169;
  assign n3171 = ~n3138 & ~n3152;
  assign n3172 = ~pi95 & ~n3171;
  assign n3173 = n3065 & ~n3172;
  assign n3174 = n2518 & n2701;
  assign n3175 = n2964 & n3174;
  assign n3176 = ~n2442 & ~n3175;
  assign n3177 = ~n2740 & ~n3176;
  assign n3178 = ~pi95 & n3143;
  assign n3179 = ~n3177 & ~n3178;
  assign n3180 = pi137 & ~n3179;
  assign n3181 = pi210 & ~n3180;
  assign n3182 = ~n3173 & n3181;
  assign n3183 = n2648 & ~n3182;
  assign n3184 = ~n3170 & n3183;
  assign n3185 = n2665 & ~n3148;
  assign n3186 = ~n3184 & n3185;
  assign n3187 = pi146 & n3170;
  assign n3188 = ~pi146 & ~pi210;
  assign n3189 = ~n3078 & ~n3152;
  assign n3190 = ~pi95 & ~n3189;
  assign n3191 = ~n2740 & ~n3190;
  assign n3192 = ~pi137 & ~n3191;
  assign n3193 = ~n3168 & ~n3192;
  assign n3194 = n3188 & ~n3193;
  assign n3195 = n3183 & ~n3194;
  assign n3196 = ~n3187 & n3195;
  assign n3197 = ~n3078 & ~n3111;
  assign n3198 = ~pi95 & ~n3197;
  assign n3199 = n2741 & ~n3198;
  assign n3200 = ~pi137 & ~n3199;
  assign n3201 = ~n3087 & ~n3200;
  assign n3202 = n3188 & ~n3201;
  assign n3203 = pi146 & n3136;
  assign n3204 = n3147 & ~n3202;
  assign n3205 = ~n3203 & n3204;
  assign n3206 = ~n2665 & ~n3196;
  assign n3207 = ~n3205 & n3206;
  assign n3208 = ~pi153 & ~n3186;
  assign n3209 = ~n3207 & n3208;
  assign n3210 = ~n3075 & ~n3209;
  assign n3211 = ~pi228 & ~n3210;
  assign n3212 = ~pi216 & ~n3211;
  assign n3213 = ~n3021 & n3212;
  assign n3214 = ~n2440 & ~n3213;
  assign n3215 = ~pi221 & ~n3214;
  assign n3216 = ~n2457 & ~n3215;
  assign n3217 = ~pi215 & ~n3216;
  assign n3218 = pi299 & ~n2438;
  assign n3219 = ~n3217 & n3218;
  assign n3220 = pi198 & ~n2975;
  assign n3221 = ~pi198 & ~n2993;
  assign n3222 = ~n3220 & ~n3221;
  assign n3223 = pi234 & n3222;
  assign n3224 = pi198 & ~n2912;
  assign n3225 = ~pi198 & ~n2949;
  assign n3226 = ~n3224 & ~n3225;
  assign n3227 = ~pi234 & n3226;
  assign n3228 = ~pi332 & ~n3227;
  assign n3229 = ~n3223 & n3228;
  assign n3230 = n2652 & ~n3229;
  assign n3231 = pi142 & n3222;
  assign n3232 = ~pi198 & ~n3001;
  assign n3233 = ~pi142 & ~n3220;
  assign n3234 = ~n3232 & n3233;
  assign n3235 = n2653 & ~n3231;
  assign n3236 = ~n3234 & n3235;
  assign n3237 = pi142 & n3226;
  assign n3238 = ~pi198 & ~n3012;
  assign n3239 = ~pi142 & ~n3224;
  assign n3240 = ~n3238 & n3239;
  assign n3241 = n2648 & ~n3237;
  assign n3242 = ~n3240 & n3241;
  assign n3243 = n2642 & ~n3242;
  assign n3244 = ~n3236 & n3243;
  assign n3245 = ~n3230 & ~n3244;
  assign n3246 = n2608 & ~n3245;
  assign n3247 = n2607 & ~n3246;
  assign n3248 = ~pi39 & ~n3247;
  assign n3249 = ~n3219 & n3248;
  assign n3250 = ~pi38 & ~n2700;
  assign n3251 = ~n3249 & n3250;
  assign n3252 = ~pi100 & ~n2699;
  assign n3253 = ~n3251 & n3252;
  assign n3254 = ~pi87 & ~n2696;
  assign n3255 = ~n3253 & n3254;
  assign n3256 = ~pi75 & ~n2638;
  assign n3257 = ~n3255 & n3256;
  assign n3258 = ~n2612 & ~n2615;
  assign n3259 = n2448 & ~n2673;
  assign n3260 = ~n2440 & ~n3259;
  assign n3261 = ~pi221 & ~n3260;
  assign n3262 = ~n2457 & ~n3261;
  assign n3263 = ~pi215 & ~n3262;
  assign n3264 = ~n2438 & ~n3263;
  assign n3265 = pi299 & ~n3264;
  assign n3266 = n2615 & ~n2662;
  assign n3267 = ~n3265 & n3266;
  assign n3268 = pi75 & ~n3258;
  assign n3269 = ~n3267 & n3268;
  assign n3270 = ~n3257 & ~n3269;
  assign n3271 = ~pi92 & ~n3270;
  assign n3272 = ~pi54 & ~n2637;
  assign n3273 = ~n3271 & n3272;
  assign n3274 = ~pi74 & ~n2627;
  assign n3275 = ~n3273 & n3274;
  assign n3276 = pi54 & ~n2612;
  assign n3277 = ~pi54 & n2626;
  assign n3278 = pi74 & ~n3276;
  assign n3279 = ~n3277 & n3278;
  assign n3280 = ~n3275 & ~n3279;
  assign n3281 = ~pi55 & ~n3280;
  assign n3282 = ~pi56 & ~n2594;
  assign n3283 = ~n3281 & n3282;
  assign n3284 = ~pi62 & ~n2571;
  assign n3285 = ~n3283 & n3284;
  assign n3286 = ~pi59 & ~n2570;
  assign n3287 = ~n3285 & n3286;
  assign n3288 = ~pi57 & ~n2545;
  assign n3289 = ~n3287 & n3288;
  assign po153 = n2543 | n3289;
  assign n3291 = ~pi57 & ~pi59;
  assign n3292 = pi215 & pi1146;
  assign n3293 = pi216 & ~pi221;
  assign n3294 = pi276 & n3293;
  assign n3295 = ~pi1146 & ~n2452;
  assign n3296 = ~pi939 & n2452;
  assign n3297 = pi221 & ~n3295;
  assign n3298 = ~n3296 & n3297;
  assign n3299 = ~n3294 & ~n3298;
  assign n3300 = ~pi215 & ~n3299;
  assign n3301 = ~n3292 & ~n3300;
  assign n3302 = ~pi216 & ~pi221;
  assign n3303 = ~pi215 & n3302;
  assign n3304 = ~n2441 & n3303;
  assign n3305 = ~pi154 & n3304;
  assign n3306 = n3301 & ~n3305;
  assign n3307 = ~n3291 & n3306;
  assign n3308 = ~pi216 & ~pi228;
  assign n3309 = ~n3292 & n3308;
  assign n3310 = ~n3298 & n3309;
  assign n3311 = n2523 & n3310;
  assign n3312 = pi154 & ~n3301;
  assign n3313 = n3311 & ~n3312;
  assign n3314 = ~pi55 & n2577;
  assign n3315 = ~n3313 & n3314;
  assign n3316 = ~pi56 & n2537;
  assign n3317 = n2532 & n3316;
  assign n3318 = ~n3315 & n3317;
  assign n3319 = pi62 & ~n3306;
  assign n3320 = ~n3318 & n3319;
  assign n3321 = ~n2538 & ~n3306;
  assign n3322 = ~n3306 & n3315;
  assign n3323 = pi56 & ~n3321;
  assign n3324 = ~n3322 & n3323;
  assign n3325 = n2577 & n3313;
  assign n3326 = pi55 & ~n3306;
  assign n3327 = ~n3325 & n3326;
  assign n3328 = ~pi222 & pi224;
  assign n3329 = pi276 & n3328;
  assign n3330 = ~pi1146 & ~n2596;
  assign n3331 = ~pi939 & n2596;
  assign n3332 = pi222 & ~n3330;
  assign n3333 = ~n3331 & n3332;
  assign n3334 = ~pi223 & ~n3333;
  assign n3335 = ~n3329 & n3334;
  assign n3336 = pi223 & ~pi1146;
  assign n3337 = ~pi299 & ~n3336;
  assign n3338 = ~n3335 & n3337;
  assign n3339 = pi299 & ~n3306;
  assign n3340 = ~n3338 & ~n3339;
  assign n3341 = ~n2533 & n3340;
  assign n3342 = pi299 & ~n3301;
  assign n3343 = ~n3338 & ~n3342;
  assign n3344 = pi154 & ~n3343;
  assign n3345 = n3301 & ~n3304;
  assign n3346 = pi299 & ~n3345;
  assign n3347 = ~n3311 & n3346;
  assign n3348 = ~n3338 & ~n3347;
  assign n3349 = ~pi154 & ~n3348;
  assign n3350 = n2532 & ~n3344;
  assign n3351 = ~n3349 & n3350;
  assign n3352 = n2534 & n3351;
  assign n3353 = n2532 & n2534;
  assign n3354 = n3340 & ~n3353;
  assign n3355 = pi92 & ~n3354;
  assign n3356 = ~n3352 & n3355;
  assign n3357 = pi75 & n3340;
  assign n3358 = ~n2628 & n3340;
  assign n3359 = ~n3351 & ~n3358;
  assign n3360 = pi87 & ~n3359;
  assign n3361 = ~pi154 & pi299;
  assign n3362 = pi146 & pi252;
  assign n3363 = n2523 & ~n3362;
  assign n3364 = pi152 & ~n3363;
  assign n3365 = ~pi252 & n2523;
  assign n3366 = ~pi161 & ~pi166;
  assign n3367 = n3365 & n3366;
  assign n3368 = n3363 & ~n3366;
  assign n3369 = ~pi152 & ~n3367;
  assign n3370 = ~n3368 & n3369;
  assign n3371 = ~n3364 & ~n3370;
  assign n3372 = n2531 & n3361;
  assign n3373 = n3310 & n3372;
  assign n3374 = n3371 & n3373;
  assign n3375 = pi100 & ~n3340;
  assign n3376 = ~n3374 & n3375;
  assign n3377 = pi38 & n3340;
  assign n3378 = pi39 & ~n2523;
  assign n3379 = ~pi70 & n3028;
  assign n3380 = ~n2728 & ~n3081;
  assign n3381 = ~n3379 & n3380;
  assign n3382 = ~pi51 & ~n3381;
  assign n3383 = n2748 & ~n3382;
  assign n3384 = n3149 & ~n3383;
  assign n3385 = ~n2744 & ~n3384;
  assign n3386 = n2462 & ~n3385;
  assign n3387 = pi40 & ~n2511;
  assign n3388 = pi32 & ~n2713;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = ~n3386 & n3389;
  assign n3391 = ~pi95 & ~n3390;
  assign n3392 = ~n2740 & ~n3391;
  assign n3393 = ~pi39 & ~n3392;
  assign n3394 = ~n3378 & ~n3393;
  assign n3395 = n3310 & n3394;
  assign n3396 = n3346 & ~n3395;
  assign n3397 = ~n3338 & ~n3396;
  assign n3398 = ~pi154 & ~n3397;
  assign n3399 = ~pi38 & ~n3344;
  assign n3400 = ~n3398 & n3399;
  assign n3401 = ~pi100 & ~n3377;
  assign n3402 = ~n3400 & n3401;
  assign n3403 = ~pi87 & ~n3376;
  assign n3404 = ~n3402 & n3403;
  assign n3405 = ~n3360 & ~n3404;
  assign n3406 = ~pi75 & ~n3405;
  assign n3407 = ~pi92 & ~n3357;
  assign n3408 = ~n3406 & n3407;
  assign n3409 = n2533 & ~n3356;
  assign n3410 = ~n3408 & n3409;
  assign n3411 = ~pi55 & ~n3341;
  assign n3412 = ~n3410 & n3411;
  assign n3413 = ~pi56 & ~n3327;
  assign n3414 = ~n3412 & n3413;
  assign n3415 = ~pi62 & ~n3324;
  assign n3416 = ~n3414 & n3415;
  assign n3417 = n3291 & ~n3320;
  assign n3418 = ~n3416 & n3417;
  assign n3419 = ~pi239 & ~n3307;
  assign n3420 = ~n3418 & n3419;
  assign n3421 = n2441 & n2442;
  assign n3422 = n3303 & n3421;
  assign n3423 = n3306 & ~n3422;
  assign n3424 = ~n3291 & n3423;
  assign n3425 = ~n3317 & ~n3423;
  assign n3426 = n3301 & ~n3422;
  assign n3427 = pi154 & ~n3426;
  assign n3428 = n3311 & ~n3427;
  assign n3429 = ~n3423 & ~n3428;
  assign n3430 = n3314 & n3429;
  assign n3431 = ~pi56 & n3430;
  assign n3432 = ~n3425 & ~n3431;
  assign n3433 = pi62 & ~n3432;
  assign n3434 = ~n2538 & ~n3423;
  assign n3435 = pi56 & ~n3434;
  assign n3436 = ~n3430 & n3435;
  assign n3437 = n2577 & n3428;
  assign n3438 = pi55 & ~n3423;
  assign n3439 = ~n3437 & n3438;
  assign n3440 = n2442 & n2609;
  assign n3441 = ~pi299 & n3440;
  assign n3442 = pi299 & ~n3423;
  assign n3443 = ~n3338 & ~n3441;
  assign n3444 = ~n3442 & n3443;
  assign n3445 = ~n2533 & n3444;
  assign n3446 = pi299 & ~n3429;
  assign n3447 = n2628 & n3446;
  assign n3448 = n2534 & n3447;
  assign n3449 = pi92 & ~n3444;
  assign n3450 = ~n3448 & n3449;
  assign n3451 = pi75 & n3444;
  assign n3452 = pi87 & ~n3444;
  assign n3453 = ~n3447 & n3452;
  assign n3454 = ~n3444 & ~n3446;
  assign n3455 = pi39 & ~n3454;
  assign n3456 = ~pi224 & n3176;
  assign n3457 = ~n2608 & ~n3329;
  assign n3458 = ~n3456 & ~n3457;
  assign n3459 = n3334 & ~n3458;
  assign n3460 = n3337 & ~n3459;
  assign n3461 = ~pi72 & ~n3383;
  assign n3462 = ~n2744 & ~n3461;
  assign n3463 = n2462 & ~n3462;
  assign n3464 = n3389 & ~n3463;
  assign n3465 = ~pi95 & ~n3464;
  assign n3466 = n2741 & ~n3465;
  assign n3467 = ~pi228 & n3466;
  assign n3468 = n2441 & n3176;
  assign n3469 = ~n3467 & ~n3468;
  assign n3470 = ~pi154 & ~n3469;
  assign n3471 = pi105 & ~n3176;
  assign n3472 = pi228 & ~n3471;
  assign n3473 = ~pi228 & ~n3177;
  assign n3474 = ~n3472 & ~n3473;
  assign n3475 = pi154 & ~n3474;
  assign n3476 = n3303 & ~n3475;
  assign n3477 = ~n3470 & n3476;
  assign n3478 = n3301 & ~n3477;
  assign n3479 = pi299 & ~n3478;
  assign n3480 = ~pi39 & ~n3460;
  assign n3481 = ~n3479 & n3480;
  assign n3482 = n2613 & ~n3455;
  assign n3483 = ~n3481 & n3482;
  assign n3484 = pi100 & n3374;
  assign n3485 = ~n2613 & ~n3444;
  assign n3486 = ~n3484 & n3485;
  assign n3487 = ~n3483 & ~n3486;
  assign n3488 = ~pi87 & ~n3487;
  assign n3489 = ~pi75 & ~n3453;
  assign n3490 = ~n3488 & n3489;
  assign n3491 = ~pi92 & ~n3451;
  assign n3492 = ~n3490 & n3491;
  assign n3493 = n2533 & ~n3450;
  assign n3494 = ~n3492 & n3493;
  assign n3495 = ~pi55 & ~n3445;
  assign n3496 = ~n3494 & n3495;
  assign n3497 = ~pi56 & ~n3439;
  assign n3498 = ~n3496 & n3497;
  assign n3499 = ~pi62 & ~n3436;
  assign n3500 = ~n3498 & n3499;
  assign n3501 = n3291 & ~n3433;
  assign n3502 = ~n3500 & n3501;
  assign n3503 = pi239 & ~n3424;
  assign n3504 = ~n3502 & n3503;
  assign po154 = n3420 | n3504;
  assign n3506 = pi215 & pi1145;
  assign n3507 = pi216 & pi274;
  assign n3508 = ~pi221 & ~n3507;
  assign n3509 = ~pi151 & ~n2441;
  assign n3510 = ~pi216 & ~n3509;
  assign n3511 = n3508 & ~n3510;
  assign n3512 = ~pi1145 & ~n2452;
  assign n3513 = ~pi927 & n2452;
  assign n3514 = pi221 & ~n3512;
  assign n3515 = ~n3513 & n3514;
  assign n3516 = ~n3511 & ~n3515;
  assign n3517 = ~pi215 & ~n3516;
  assign n3518 = ~n3506 & ~n3517;
  assign n3519 = n2461 & n3421;
  assign n3520 = ~n3507 & n3519;
  assign n3521 = n3518 & ~n3520;
  assign n3522 = ~n3317 & n3521;
  assign n3523 = ~n3421 & ~n3509;
  assign n3524 = ~pi228 & n2523;
  assign n3525 = ~pi151 & n3524;
  assign n3526 = ~n3523 & ~n3525;
  assign n3527 = ~pi216 & ~n3526;
  assign n3528 = n3508 & ~n3527;
  assign n3529 = ~n3515 & ~n3528;
  assign n3530 = ~pi215 & ~n3529;
  assign n3531 = ~n3506 & ~n3530;
  assign n3532 = n3317 & n3531;
  assign n3533 = pi62 & ~n3522;
  assign n3534 = ~n3532 & n3533;
  assign n3535 = n2538 & ~n3531;
  assign n3536 = ~n2538 & ~n3521;
  assign n3537 = pi56 & ~n3536;
  assign n3538 = ~n3535 & n3537;
  assign n3539 = ~n2577 & n3521;
  assign n3540 = n2577 & n3531;
  assign n3541 = pi55 & ~n3539;
  assign n3542 = ~n3540 & n3541;
  assign n3543 = pi223 & pi1145;
  assign n3544 = ~pi1145 & ~n2596;
  assign n3545 = ~pi927 & n2596;
  assign n3546 = pi222 & ~n3544;
  assign n3547 = ~n3545 & n3546;
  assign n3548 = pi224 & pi274;
  assign n3549 = n3328 & ~n3548;
  assign n3550 = ~n3547 & ~n3549;
  assign n3551 = ~pi223 & ~n3550;
  assign n3552 = ~n3543 & ~n3551;
  assign n3553 = ~pi299 & ~n3552;
  assign n3554 = ~n3441 & ~n3553;
  assign n3555 = pi299 & ~n3521;
  assign n3556 = n3554 & ~n3555;
  assign n3557 = ~n2533 & n3556;
  assign n3558 = ~n2628 & n3556;
  assign n3559 = pi299 & ~n3531;
  assign n3560 = n3554 & ~n3559;
  assign n3561 = n2628 & n3560;
  assign n3562 = ~n3558 & ~n3561;
  assign n3563 = n2534 & ~n3562;
  assign n3564 = ~n2534 & n3556;
  assign n3565 = pi92 & ~n3564;
  assign n3566 = ~n3563 & n3565;
  assign n3567 = pi75 & n3556;
  assign n3568 = pi87 & n3562;
  assign n3569 = pi38 & n3556;
  assign n3570 = pi39 & ~n3560;
  assign n3571 = ~pi222 & ~n3548;
  assign n3572 = ~n3456 & n3571;
  assign n3573 = ~n3547 & ~n3572;
  assign n3574 = ~pi223 & ~n3573;
  assign n3575 = ~pi299 & ~n3543;
  assign n3576 = ~n3574 & n3575;
  assign n3577 = pi151 & n3474;
  assign n3578 = ~pi151 & n3469;
  assign n3579 = ~pi216 & ~n3577;
  assign n3580 = ~n3578 & n3579;
  assign n3581 = n3508 & ~n3580;
  assign n3582 = ~n3515 & ~n3581;
  assign n3583 = ~pi215 & ~n3582;
  assign n3584 = pi299 & ~n3506;
  assign n3585 = ~n3583 & n3584;
  assign n3586 = ~pi39 & ~n3576;
  assign n3587 = ~n3585 & n3586;
  assign n3588 = ~pi38 & ~n3570;
  assign n3589 = ~n3587 & n3588;
  assign n3590 = ~pi100 & ~n3569;
  assign n3591 = ~n3589 & n3590;
  assign n3592 = ~n2531 & n3556;
  assign n3593 = ~pi228 & n3371;
  assign n3594 = n2441 & ~n2442;
  assign n3595 = ~n3593 & ~n3594;
  assign n3596 = ~pi151 & n3595;
  assign n3597 = n3527 & ~n3596;
  assign n3598 = n3508 & ~n3597;
  assign n3599 = ~n3515 & ~n3598;
  assign n3600 = ~pi215 & ~n3599;
  assign n3601 = ~n3506 & ~n3600;
  assign n3602 = pi299 & ~n3601;
  assign n3603 = n2531 & n3554;
  assign n3604 = ~n3602 & n3603;
  assign n3605 = pi100 & ~n3592;
  assign n3606 = ~n3604 & n3605;
  assign n3607 = ~n3591 & ~n3606;
  assign n3608 = ~pi87 & ~n3607;
  assign n3609 = ~pi75 & ~n3568;
  assign n3610 = ~n3608 & n3609;
  assign n3611 = ~pi92 & ~n3567;
  assign n3612 = ~n3610 & n3611;
  assign n3613 = n2533 & ~n3566;
  assign n3614 = ~n3612 & n3613;
  assign n3615 = ~pi55 & ~n3557;
  assign n3616 = ~n3614 & n3615;
  assign n3617 = ~pi56 & ~n3542;
  assign n3618 = ~n3616 & n3617;
  assign n3619 = ~pi62 & ~n3538;
  assign n3620 = ~n3618 & n3619;
  assign n3621 = pi235 & n3291;
  assign n3622 = ~n3534 & n3621;
  assign n3623 = ~n3620 & n3622;
  assign n3624 = n3308 & ~n3506;
  assign n3625 = ~n3515 & n3624;
  assign n3626 = n2523 & n3625;
  assign n3627 = n3317 & n3626;
  assign n3628 = pi62 & ~n3518;
  assign n3629 = ~n3627 & n3628;
  assign n3630 = n2538 & n3626;
  assign n3631 = ~n3518 & ~n3630;
  assign n3632 = pi56 & ~n3631;
  assign n3633 = n2577 & n3626;
  assign n3634 = pi55 & ~n3518;
  assign n3635 = ~n3633 & n3634;
  assign n3636 = pi299 & ~n3518;
  assign n3637 = ~n3553 & ~n3636;
  assign n3638 = ~n2533 & n3637;
  assign n3639 = ~n3626 & n3636;
  assign n3640 = n2532 & ~n3553;
  assign n3641 = ~n3639 & n3640;
  assign n3642 = n2534 & n3641;
  assign n3643 = ~n3353 & n3637;
  assign n3644 = pi92 & ~n3643;
  assign n3645 = ~n3642 & n3644;
  assign n3646 = pi75 & n3637;
  assign n3647 = ~n2628 & n3637;
  assign n3648 = ~n3641 & ~n3647;
  assign n3649 = pi87 & ~n3648;
  assign n3650 = ~pi100 & n3394;
  assign n3651 = ~pi39 & pi100;
  assign n3652 = n3371 & n3651;
  assign n3653 = ~n3650 & ~n3652;
  assign n3654 = ~pi38 & n3625;
  assign n3655 = ~n3653 & n3654;
  assign n3656 = n3636 & ~n3655;
  assign n3657 = ~pi87 & ~n3553;
  assign n3658 = ~n3656 & n3657;
  assign n3659 = ~n3649 & ~n3658;
  assign n3660 = ~pi75 & ~n3659;
  assign n3661 = ~pi92 & ~n3646;
  assign n3662 = ~n3660 & n3661;
  assign n3663 = n2533 & ~n3645;
  assign n3664 = ~n3662 & n3663;
  assign n3665 = ~pi55 & ~n3638;
  assign n3666 = ~n3664 & n3665;
  assign n3667 = ~pi56 & ~n3635;
  assign n3668 = ~n3666 & n3667;
  assign n3669 = ~pi62 & ~n3632;
  assign n3670 = ~n3668 & n3669;
  assign n3671 = ~pi235 & n3291;
  assign n3672 = ~n3629 & n3671;
  assign n3673 = ~n3670 & n3672;
  assign n3674 = pi235 & n3520;
  assign n3675 = ~n3291 & ~n3674;
  assign n3676 = n3518 & n3675;
  assign n3677 = ~n3673 & ~n3676;
  assign po155 = ~n3623 & n3677;
  assign n3679 = pi215 & pi1143;
  assign n3680 = pi216 & pi264;
  assign n3681 = ~pi221 & ~n3680;
  assign n3682 = ~pi105 & pi146;
  assign n3683 = pi284 & ~n2442;
  assign n3684 = pi105 & ~n3683;
  assign n3685 = pi228 & ~n3682;
  assign n3686 = ~n3684 & n3685;
  assign n3687 = ~n3421 & ~n3686;
  assign n3688 = ~pi146 & ~pi228;
  assign n3689 = n3687 & ~n3688;
  assign n3690 = ~pi216 & ~n3689;
  assign n3691 = n3681 & ~n3690;
  assign n3692 = ~pi1143 & ~n2452;
  assign n3693 = ~pi944 & n2452;
  assign n3694 = pi221 & ~n3692;
  assign n3695 = ~n3693 & n3694;
  assign n3696 = ~n3691 & ~n3695;
  assign n3697 = ~pi215 & ~n3696;
  assign n3698 = ~n3679 & ~n3697;
  assign n3699 = ~n3317 & n3698;
  assign n3700 = ~pi284 & n2523;
  assign n3701 = ~n3524 & ~n3688;
  assign n3702 = ~n3700 & ~n3701;
  assign n3703 = n3687 & ~n3702;
  assign n3704 = ~pi216 & ~n3703;
  assign n3705 = n3681 & ~n3704;
  assign n3706 = ~n3695 & ~n3705;
  assign n3707 = ~pi215 & ~n3706;
  assign n3708 = ~n3679 & ~n3707;
  assign n3709 = n3317 & n3708;
  assign n3710 = pi62 & ~n3699;
  assign n3711 = ~n3709 & n3710;
  assign n3712 = n2538 & ~n3708;
  assign n3713 = ~n2538 & ~n3698;
  assign n3714 = pi56 & ~n3713;
  assign n3715 = ~n3712 & n3714;
  assign n3716 = ~n2577 & n3698;
  assign n3717 = n2577 & n3708;
  assign n3718 = pi55 & ~n3716;
  assign n3719 = ~n3717 & n3718;
  assign n3720 = pi223 & pi1143;
  assign n3721 = pi224 & pi264;
  assign n3722 = ~pi222 & ~n3721;
  assign n3723 = ~pi224 & n3683;
  assign n3724 = n3722 & ~n3723;
  assign n3725 = ~pi1143 & ~n2596;
  assign n3726 = ~pi944 & n2596;
  assign n3727 = pi222 & ~n3725;
  assign n3728 = ~n3726 & n3727;
  assign n3729 = ~n3724 & ~n3728;
  assign n3730 = ~pi223 & ~n3729;
  assign n3731 = ~n3720 & ~n3730;
  assign n3732 = ~pi299 & ~n3731;
  assign n3733 = ~n3440 & n3732;
  assign n3734 = pi299 & ~n3698;
  assign n3735 = ~n3733 & ~n3734;
  assign n3736 = ~n2533 & n3735;
  assign n3737 = ~n2628 & n3735;
  assign n3738 = pi299 & ~n3708;
  assign n3739 = ~n3733 & ~n3738;
  assign n3740 = n2628 & n3739;
  assign n3741 = ~n3737 & ~n3740;
  assign n3742 = n2534 & ~n3741;
  assign n3743 = ~n2534 & n3735;
  assign n3744 = pi92 & ~n3743;
  assign n3745 = ~n3742 & n3744;
  assign n3746 = pi75 & n3735;
  assign n3747 = pi87 & n3741;
  assign n3748 = pi38 & n3735;
  assign n3749 = pi39 & ~n3739;
  assign n3750 = ~pi299 & ~n3720;
  assign n3751 = ~pi284 & n3176;
  assign n3752 = ~pi224 & ~n3751;
  assign n3753 = n3722 & ~n3752;
  assign n3754 = ~n3728 & ~n3753;
  assign n3755 = n3750 & n3754;
  assign n3756 = pi299 & ~n3679;
  assign n3757 = n2441 & ~n3176;
  assign n3758 = pi146 & ~n3392;
  assign n3759 = pi284 & ~n3758;
  assign n3760 = pi146 & ~n3177;
  assign n3761 = ~pi146 & n3466;
  assign n3762 = ~pi284 & ~n3760;
  assign n3763 = ~n3761 & n3762;
  assign n3764 = ~n3759 & ~n3763;
  assign n3765 = ~pi228 & ~n3764;
  assign n3766 = ~n3686 & ~n3757;
  assign n3767 = ~n3765 & n3766;
  assign n3768 = ~pi216 & ~n3767;
  assign n3769 = n3681 & ~n3768;
  assign n3770 = ~n3695 & ~n3769;
  assign n3771 = ~pi215 & ~n3770;
  assign n3772 = n3756 & ~n3771;
  assign n3773 = ~n3176 & n3722;
  assign n3774 = n3754 & ~n3773;
  assign n3775 = ~pi223 & ~n3774;
  assign n3776 = n3750 & ~n3775;
  assign n3777 = ~pi39 & ~n3776;
  assign n3778 = ~n3755 & n3777;
  assign n3779 = ~n3772 & n3778;
  assign n3780 = ~pi38 & ~n3749;
  assign n3781 = ~n3779 & n3780;
  assign n3782 = ~pi100 & ~n3748;
  assign n3783 = ~n3781 & n3782;
  assign n3784 = ~n2531 & n3735;
  assign n3785 = pi252 & n2665;
  assign n3786 = n3700 & ~n3785;
  assign n3787 = pi146 & ~n3365;
  assign n3788 = ~pi228 & ~n3786;
  assign n3789 = ~n3787 & n3788;
  assign n3790 = n3687 & ~n3789;
  assign n3791 = ~pi216 & ~n3790;
  assign n3792 = n3681 & ~n3791;
  assign n3793 = ~n3695 & ~n3792;
  assign n3794 = ~pi215 & ~n3793;
  assign n3795 = ~n3679 & ~n3794;
  assign n3796 = pi299 & ~n3795;
  assign n3797 = n2531 & ~n3733;
  assign n3798 = ~n3796 & n3797;
  assign n3799 = pi100 & ~n3784;
  assign n3800 = ~n3798 & n3799;
  assign n3801 = ~n3783 & ~n3800;
  assign n3802 = ~pi87 & ~n3801;
  assign n3803 = ~pi75 & ~n3747;
  assign n3804 = ~n3802 & n3803;
  assign n3805 = ~pi92 & ~n3746;
  assign n3806 = ~n3804 & n3805;
  assign n3807 = n2533 & ~n3745;
  assign n3808 = ~n3806 & n3807;
  assign n3809 = ~pi55 & ~n3736;
  assign n3810 = ~n3808 & n3809;
  assign n3811 = ~pi56 & ~n3719;
  assign n3812 = ~n3810 & n3811;
  assign n3813 = ~pi62 & ~n3715;
  assign n3814 = ~n3812 & n3813;
  assign n3815 = ~pi238 & n3291;
  assign n3816 = ~n3711 & n3815;
  assign n3817 = ~n3814 & n3816;
  assign n3818 = ~n3686 & ~n3702;
  assign n3819 = ~pi216 & ~n3818;
  assign n3820 = n3681 & ~n3819;
  assign n3821 = ~n3695 & ~n3820;
  assign n3822 = ~pi215 & ~n3821;
  assign n3823 = ~n3679 & ~n3822;
  assign n3824 = n3317 & n3823;
  assign n3825 = n3519 & ~n3680;
  assign n3826 = n3698 & ~n3825;
  assign n3827 = ~n3317 & n3826;
  assign n3828 = pi62 & ~n3827;
  assign n3829 = ~n3824 & n3828;
  assign n3830 = n2538 & ~n3823;
  assign n3831 = ~n2538 & ~n3826;
  assign n3832 = pi56 & ~n3831;
  assign n3833 = ~n3830 & n3832;
  assign n3834 = ~n2577 & n3826;
  assign n3835 = n2577 & n3823;
  assign n3836 = pi55 & ~n3834;
  assign n3837 = ~n3835 & n3836;
  assign n3838 = pi299 & ~n3826;
  assign n3839 = ~n3732 & ~n3838;
  assign n3840 = ~n2533 & n3839;
  assign n3841 = ~n2628 & n3839;
  assign n3842 = pi299 & ~n3823;
  assign n3843 = ~n3732 & ~n3842;
  assign n3844 = n2628 & n3843;
  assign n3845 = ~n3841 & ~n3844;
  assign n3846 = n2534 & ~n3845;
  assign n3847 = ~n2534 & n3839;
  assign n3848 = pi92 & ~n3847;
  assign n3849 = ~n3846 & n3848;
  assign n3850 = pi75 & n3839;
  assign n3851 = pi87 & n3845;
  assign n3852 = pi38 & n3839;
  assign n3853 = pi39 & ~n3843;
  assign n3854 = ~n3471 & n3686;
  assign n3855 = ~pi146 & n3177;
  assign n3856 = pi146 & ~n3466;
  assign n3857 = pi284 & ~n3855;
  assign n3858 = ~n3856 & n3857;
  assign n3859 = ~pi146 & ~pi284;
  assign n3860 = ~n3392 & n3859;
  assign n3861 = ~n3858 & ~n3860;
  assign n3862 = ~pi228 & ~n3861;
  assign n3863 = ~n3854 & ~n3862;
  assign n3864 = ~pi216 & ~n3863;
  assign n3865 = n3681 & ~n3864;
  assign n3866 = ~n3695 & ~n3865;
  assign n3867 = ~pi215 & ~n3866;
  assign n3868 = n3756 & ~n3867;
  assign n3869 = n3777 & ~n3868;
  assign n3870 = ~pi38 & ~n3853;
  assign n3871 = ~n3869 & n3870;
  assign n3872 = ~pi100 & ~n3852;
  assign n3873 = ~n3871 & n3872;
  assign n3874 = ~n2531 & n3839;
  assign n3875 = ~n3686 & ~n3789;
  assign n3876 = ~pi216 & ~n3875;
  assign n3877 = n3681 & ~n3876;
  assign n3878 = ~n3695 & ~n3877;
  assign n3879 = ~pi215 & ~n3878;
  assign n3880 = ~n3679 & ~n3879;
  assign n3881 = pi299 & ~n3880;
  assign n3882 = n2531 & ~n3732;
  assign n3883 = ~n3881 & n3882;
  assign n3884 = pi100 & ~n3874;
  assign n3885 = ~n3883 & n3884;
  assign n3886 = ~n3873 & ~n3885;
  assign n3887 = ~pi87 & ~n3886;
  assign n3888 = ~pi75 & ~n3851;
  assign n3889 = ~n3887 & n3888;
  assign n3890 = ~pi92 & ~n3850;
  assign n3891 = ~n3889 & n3890;
  assign n3892 = n2533 & ~n3849;
  assign n3893 = ~n3891 & n3892;
  assign n3894 = ~pi55 & ~n3840;
  assign n3895 = ~n3893 & n3894;
  assign n3896 = ~pi56 & ~n3837;
  assign n3897 = ~n3895 & n3896;
  assign n3898 = ~pi62 & ~n3833;
  assign n3899 = ~n3897 & n3898;
  assign n3900 = pi238 & n3291;
  assign n3901 = ~n3829 & n3900;
  assign n3902 = ~n3899 & n3901;
  assign n3903 = pi238 & n3825;
  assign n3904 = ~n3291 & ~n3903;
  assign n3905 = n3698 & n3904;
  assign n3906 = ~n3817 & ~n3905;
  assign po156 = ~n3902 & n3906;
  assign n3908 = pi215 & pi1142;
  assign n3909 = pi216 & pi277;
  assign n3910 = ~pi221 & ~n3909;
  assign n3911 = pi172 & ~pi228;
  assign n3912 = pi262 & ~n2442;
  assign n3913 = pi105 & n3912;
  assign n3914 = ~pi105 & pi172;
  assign n3915 = ~n3913 & ~n3914;
  assign n3916 = pi228 & ~n3915;
  assign n3917 = ~n3911 & ~n3916;
  assign n3918 = ~pi216 & ~n3917;
  assign n3919 = n3910 & ~n3918;
  assign n3920 = ~pi1142 & ~n2452;
  assign n3921 = ~pi932 & n2452;
  assign n3922 = pi221 & ~n3920;
  assign n3923 = ~n3921 & n3922;
  assign n3924 = ~n3919 & ~n3923;
  assign n3925 = ~pi215 & ~n3924;
  assign n3926 = ~n3908 & ~n3925;
  assign n3927 = ~n3422 & ~n3926;
  assign n3928 = ~n3291 & ~n3927;
  assign n3929 = ~pi262 & n2523;
  assign n3930 = ~n3524 & ~n3911;
  assign n3931 = ~n3929 & ~n3930;
  assign n3932 = ~n3421 & ~n3916;
  assign n3933 = ~n3931 & n3932;
  assign n3934 = ~pi216 & ~n3933;
  assign n3935 = n3910 & ~n3934;
  assign n3936 = ~n3923 & ~n3935;
  assign n3937 = ~pi215 & ~n3936;
  assign n3938 = ~n3908 & ~n3937;
  assign n3939 = n2538 & ~n3938;
  assign n3940 = ~pi56 & n3939;
  assign n3941 = ~n3317 & n3927;
  assign n3942 = ~n3940 & ~n3941;
  assign n3943 = pi62 & ~n3942;
  assign n3944 = ~n2538 & n3927;
  assign n3945 = pi56 & ~n3944;
  assign n3946 = ~n3939 & n3945;
  assign n3947 = ~n2577 & ~n3927;
  assign n3948 = n2577 & n3938;
  assign n3949 = pi55 & ~n3947;
  assign n3950 = ~n3948 & n3949;
  assign n3951 = pi223 & pi1142;
  assign n3952 = pi224 & pi277;
  assign n3953 = ~pi222 & ~n3952;
  assign n3954 = ~pi224 & n3912;
  assign n3955 = n3953 & ~n3954;
  assign n3956 = ~pi1142 & ~n2596;
  assign n3957 = ~pi932 & n2596;
  assign n3958 = pi222 & ~n3956;
  assign n3959 = ~n3957 & n3958;
  assign n3960 = ~n3955 & ~n3959;
  assign n3961 = ~pi223 & ~n3960;
  assign n3962 = ~n3951 & ~n3961;
  assign n3963 = ~pi299 & ~n3962;
  assign n3964 = ~n3440 & n3963;
  assign n3965 = pi299 & n3927;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = ~n2533 & n3966;
  assign n3968 = ~n2628 & n3966;
  assign n3969 = pi299 & ~n3938;
  assign n3970 = ~n3964 & ~n3969;
  assign n3971 = n2628 & n3970;
  assign n3972 = ~n3968 & ~n3971;
  assign n3973 = n2534 & ~n3972;
  assign n3974 = ~n2534 & n3966;
  assign n3975 = pi92 & ~n3974;
  assign n3976 = ~n3973 & n3975;
  assign n3977 = pi75 & n3966;
  assign n3978 = pi87 & n3972;
  assign n3979 = pi38 & n3966;
  assign n3980 = pi39 & ~n3970;
  assign n3981 = ~pi299 & ~n3951;
  assign n3982 = ~pi262 & n3176;
  assign n3983 = ~pi224 & ~n3982;
  assign n3984 = n3953 & ~n3983;
  assign n3985 = ~n3959 & ~n3984;
  assign n3986 = n3981 & n3985;
  assign n3987 = ~n3176 & n3953;
  assign n3988 = n3985 & ~n3987;
  assign n3989 = ~pi223 & ~n3988;
  assign n3990 = n3981 & ~n3989;
  assign n3991 = ~pi39 & ~n3990;
  assign n3992 = pi299 & ~n3908;
  assign n3993 = ~pi262 & n3466;
  assign n3994 = pi172 & ~n3993;
  assign n3995 = pi262 & n3391;
  assign n3996 = ~pi172 & ~n2740;
  assign n3997 = ~n3982 & n3996;
  assign n3998 = ~n3995 & n3997;
  assign n3999 = ~pi228 & ~n3998;
  assign n4000 = ~n3994 & n3999;
  assign n4001 = ~n3175 & n3913;
  assign n4002 = pi228 & ~n3914;
  assign n4003 = ~n4001 & n4002;
  assign n4004 = ~n3471 & n4003;
  assign n4005 = ~pi216 & ~n4004;
  assign n4006 = ~n4000 & n4005;
  assign n4007 = n3910 & ~n4006;
  assign n4008 = ~n3923 & ~n4007;
  assign n4009 = ~pi215 & ~n4008;
  assign n4010 = n3992 & ~n4009;
  assign n4011 = ~n3986 & n3991;
  assign n4012 = ~n4010 & n4011;
  assign n4013 = ~pi38 & ~n3980;
  assign n4014 = ~n4012 & n4013;
  assign n4015 = ~pi100 & ~n3979;
  assign n4016 = ~n4014 & n4015;
  assign n4017 = ~n2531 & n3966;
  assign n4018 = ~pi262 & n3371;
  assign n4019 = ~n3593 & ~n3911;
  assign n4020 = ~n4018 & ~n4019;
  assign n4021 = n3932 & ~n4020;
  assign n4022 = ~pi216 & ~n4021;
  assign n4023 = n3910 & ~n4022;
  assign n4024 = ~n3923 & ~n4023;
  assign n4025 = ~pi215 & ~n4024;
  assign n4026 = ~n3908 & ~n4025;
  assign n4027 = pi299 & ~n4026;
  assign n4028 = n2531 & ~n3964;
  assign n4029 = ~n4027 & n4028;
  assign n4030 = pi100 & ~n4017;
  assign n4031 = ~n4029 & n4030;
  assign n4032 = ~n4016 & ~n4031;
  assign n4033 = ~pi87 & ~n4032;
  assign n4034 = ~pi75 & ~n3978;
  assign n4035 = ~n4033 & n4034;
  assign n4036 = ~pi92 & ~n3977;
  assign n4037 = ~n4035 & n4036;
  assign n4038 = n2533 & ~n3976;
  assign n4039 = ~n4037 & n4038;
  assign n4040 = ~pi55 & ~n3967;
  assign n4041 = ~n4039 & n4040;
  assign n4042 = ~pi56 & ~n3950;
  assign n4043 = ~n4041 & n4042;
  assign n4044 = ~pi62 & ~n3946;
  assign n4045 = ~n4043 & n4044;
  assign n4046 = n3291 & ~n3943;
  assign n4047 = ~n4045 & n4046;
  assign n4048 = ~pi249 & ~n3928;
  assign n4049 = ~n4047 & n4048;
  assign n4050 = ~n3291 & n3926;
  assign n4051 = ~n3317 & ~n3926;
  assign n4052 = ~n3916 & ~n3931;
  assign n4053 = ~pi216 & ~n4052;
  assign n4054 = n3910 & ~n4053;
  assign n4055 = ~n3923 & ~n4054;
  assign n4056 = ~pi215 & ~n4055;
  assign n4057 = ~n3908 & ~n4056;
  assign n4058 = n2538 & ~n4057;
  assign n4059 = ~pi56 & n4058;
  assign n4060 = ~n4051 & ~n4059;
  assign n4061 = pi62 & ~n4060;
  assign n4062 = ~n2538 & ~n3926;
  assign n4063 = pi56 & ~n4062;
  assign n4064 = ~n4058 & n4063;
  assign n4065 = ~n2577 & n3926;
  assign n4066 = n2577 & n4057;
  assign n4067 = pi55 & ~n4065;
  assign n4068 = ~n4066 & n4067;
  assign n4069 = pi299 & ~n3926;
  assign n4070 = ~n3963 & ~n4069;
  assign n4071 = ~n2533 & n4070;
  assign n4072 = ~n2628 & n4070;
  assign n4073 = pi299 & ~n4057;
  assign n4074 = ~n3963 & ~n4073;
  assign n4075 = n2628 & n4074;
  assign n4076 = ~n4072 & ~n4075;
  assign n4077 = n2534 & ~n4076;
  assign n4078 = ~n2534 & n4070;
  assign n4079 = pi92 & ~n4078;
  assign n4080 = ~n4077 & n4079;
  assign n4081 = pi75 & n4070;
  assign n4082 = pi87 & n4076;
  assign n4083 = pi38 & n4070;
  assign n4084 = pi39 & ~n4074;
  assign n4085 = pi262 & n3466;
  assign n4086 = ~pi172 & ~n4085;
  assign n4087 = ~pi262 & ~n3392;
  assign n4088 = pi262 & ~n3177;
  assign n4089 = pi172 & ~n4088;
  assign n4090 = ~n4087 & n4089;
  assign n4091 = ~n4086 & ~n4090;
  assign n4092 = ~pi228 & ~n4091;
  assign n4093 = ~pi216 & ~n4003;
  assign n4094 = ~n4092 & n4093;
  assign n4095 = n3910 & ~n4094;
  assign n4096 = ~n3923 & ~n4095;
  assign n4097 = ~pi215 & ~n4096;
  assign n4098 = n3992 & ~n4097;
  assign n4099 = n3991 & ~n4098;
  assign n4100 = ~pi38 & ~n4084;
  assign n4101 = ~n4099 & n4100;
  assign n4102 = ~pi100 & ~n4083;
  assign n4103 = ~n4101 & n4102;
  assign n4104 = ~n2531 & n4070;
  assign n4105 = ~n3916 & ~n4020;
  assign n4106 = ~pi216 & ~n4105;
  assign n4107 = n3910 & ~n4106;
  assign n4108 = ~n3923 & ~n4107;
  assign n4109 = ~pi215 & ~n4108;
  assign n4110 = ~n3908 & ~n4109;
  assign n4111 = pi299 & ~n4110;
  assign n4112 = n2531 & ~n3963;
  assign n4113 = ~n4111 & n4112;
  assign n4114 = pi100 & ~n4104;
  assign n4115 = ~n4113 & n4114;
  assign n4116 = ~n4103 & ~n4115;
  assign n4117 = ~pi87 & ~n4116;
  assign n4118 = ~pi75 & ~n4082;
  assign n4119 = ~n4117 & n4118;
  assign n4120 = ~pi92 & ~n4081;
  assign n4121 = ~n4119 & n4120;
  assign n4122 = n2533 & ~n4080;
  assign n4123 = ~n4121 & n4122;
  assign n4124 = ~pi55 & ~n4071;
  assign n4125 = ~n4123 & n4124;
  assign n4126 = ~pi56 & ~n4068;
  assign n4127 = ~n4125 & n4126;
  assign n4128 = ~pi62 & ~n4064;
  assign n4129 = ~n4127 & n4128;
  assign n4130 = n3291 & ~n4061;
  assign n4131 = ~n4129 & n4130;
  assign n4132 = pi249 & ~n4050;
  assign n4133 = ~n4131 & n4132;
  assign po157 = n4049 | n4133;
  assign n4135 = pi215 & pi1141;
  assign n4136 = pi216 & pi270;
  assign n4137 = ~pi221 & ~n4136;
  assign n4138 = ~pi105 & pi171;
  assign n4139 = pi861 & ~n2442;
  assign n4140 = pi105 & ~n4139;
  assign n4141 = pi228 & ~n4138;
  assign n4142 = ~n4140 & n4141;
  assign n4143 = ~pi216 & ~n4142;
  assign n4144 = ~pi171 & ~pi228;
  assign n4145 = n4143 & ~n4144;
  assign n4146 = n4137 & ~n4145;
  assign n4147 = ~pi1141 & ~n2452;
  assign n4148 = ~pi935 & n2452;
  assign n4149 = pi221 & ~n4147;
  assign n4150 = ~n4148 & n4149;
  assign n4151 = ~n4146 & ~n4150;
  assign n4152 = ~pi215 & ~n4151;
  assign n4153 = ~n4135 & ~n4152;
  assign n4154 = ~n3317 & n4153;
  assign n4155 = ~pi861 & n2523;
  assign n4156 = pi171 & ~n2523;
  assign n4157 = ~pi228 & ~n4155;
  assign n4158 = ~n4156 & n4157;
  assign n4159 = n4143 & ~n4158;
  assign n4160 = n4137 & ~n4159;
  assign n4161 = ~n4150 & ~n4160;
  assign n4162 = ~pi215 & ~n4161;
  assign n4163 = ~n4135 & ~n4162;
  assign n4164 = n3317 & n4163;
  assign n4165 = pi62 & ~n4154;
  assign n4166 = ~n4164 & n4165;
  assign n4167 = n2538 & ~n4163;
  assign n4168 = ~n2538 & ~n4153;
  assign n4169 = pi56 & ~n4168;
  assign n4170 = ~n4167 & n4169;
  assign n4171 = ~n2577 & n4153;
  assign n4172 = n2577 & n4163;
  assign n4173 = pi55 & ~n4171;
  assign n4174 = ~n4172 & n4173;
  assign n4175 = pi223 & pi1141;
  assign n4176 = pi224 & pi270;
  assign n4177 = ~pi222 & ~n4176;
  assign n4178 = ~pi224 & ~n4139;
  assign n4179 = n4177 & ~n4178;
  assign n4180 = ~pi1141 & ~n2596;
  assign n4181 = ~pi935 & n2596;
  assign n4182 = pi222 & ~n4180;
  assign n4183 = ~n4181 & n4182;
  assign n4184 = ~n4179 & ~n4183;
  assign n4185 = ~pi223 & ~n4184;
  assign n4186 = ~n4175 & ~n4185;
  assign n4187 = ~pi299 & ~n4186;
  assign n4188 = pi299 & ~n4153;
  assign n4189 = ~n4187 & ~n4188;
  assign n4190 = ~n2533 & n4189;
  assign n4191 = ~n2628 & n4189;
  assign n4192 = pi299 & ~n4163;
  assign n4193 = ~n4187 & ~n4192;
  assign n4194 = n2628 & n4193;
  assign n4195 = ~n4191 & ~n4194;
  assign n4196 = n2534 & ~n4195;
  assign n4197 = ~n2534 & n4189;
  assign n4198 = pi92 & ~n4197;
  assign n4199 = ~n4196 & n4198;
  assign n4200 = pi75 & n4189;
  assign n4201 = pi87 & n4195;
  assign n4202 = pi38 & n4189;
  assign n4203 = pi39 & ~n4193;
  assign n4204 = ~pi299 & ~n4175;
  assign n4205 = pi861 & n3176;
  assign n4206 = ~pi224 & ~n4205;
  assign n4207 = n4177 & ~n4206;
  assign n4208 = ~n4183 & ~n4207;
  assign n4209 = n4204 & n4208;
  assign n4210 = ~n3176 & n4177;
  assign n4211 = n4208 & ~n4210;
  assign n4212 = ~pi223 & ~n4211;
  assign n4213 = n4204 & ~n4212;
  assign n4214 = ~pi39 & ~n4213;
  assign n4215 = pi299 & ~n4135;
  assign n4216 = ~pi861 & n3391;
  assign n4217 = ~n2740 & ~n4205;
  assign n4218 = ~n4216 & n4217;
  assign n4219 = ~pi171 & ~n4218;
  assign n4220 = pi171 & pi861;
  assign n4221 = n3466 & n4220;
  assign n4222 = ~n4219 & ~n4221;
  assign n4223 = ~pi228 & ~n4222;
  assign n4224 = ~n3471 & n4142;
  assign n4225 = ~pi216 & ~n4224;
  assign n4226 = ~n4223 & n4225;
  assign n4227 = n4137 & ~n4226;
  assign n4228 = ~n4150 & ~n4227;
  assign n4229 = ~pi215 & ~n4228;
  assign n4230 = n4215 & ~n4229;
  assign n4231 = ~n4209 & n4214;
  assign n4232 = ~n4230 & n4231;
  assign n4233 = ~pi38 & ~n4203;
  assign n4234 = ~n4232 & n4233;
  assign n4235 = ~pi100 & ~n4202;
  assign n4236 = ~n4234 & n4235;
  assign n4237 = ~n2531 & n4189;
  assign n4238 = ~pi861 & n3371;
  assign n4239 = ~n3593 & ~n4144;
  assign n4240 = ~n4238 & ~n4239;
  assign n4241 = n4143 & ~n4240;
  assign n4242 = n4137 & ~n4241;
  assign n4243 = ~n4150 & ~n4242;
  assign n4244 = ~pi215 & ~n4243;
  assign n4245 = ~n4135 & ~n4244;
  assign n4246 = pi299 & ~n4245;
  assign n4247 = n2531 & ~n4187;
  assign n4248 = ~n4246 & n4247;
  assign n4249 = pi100 & ~n4237;
  assign n4250 = ~n4248 & n4249;
  assign n4251 = ~n4236 & ~n4250;
  assign n4252 = ~pi87 & ~n4251;
  assign n4253 = ~pi75 & ~n4201;
  assign n4254 = ~n4252 & n4253;
  assign n4255 = ~pi92 & ~n4200;
  assign n4256 = ~n4254 & n4255;
  assign n4257 = n2533 & ~n4199;
  assign n4258 = ~n4256 & n4257;
  assign n4259 = ~pi55 & ~n4190;
  assign n4260 = ~n4258 & n4259;
  assign n4261 = ~pi56 & ~n4174;
  assign n4262 = ~n4260 & n4261;
  assign n4263 = ~pi62 & ~n4170;
  assign n4264 = ~n4262 & n4263;
  assign n4265 = ~pi241 & n3291;
  assign n4266 = ~n4166 & n4265;
  assign n4267 = ~n4264 & n4266;
  assign n4268 = ~n3421 & n4143;
  assign n4269 = ~n4158 & n4268;
  assign n4270 = n4137 & ~n4269;
  assign n4271 = ~n4150 & ~n4270;
  assign n4272 = ~pi215 & ~n4271;
  assign n4273 = ~n4135 & ~n4272;
  assign n4274 = n3317 & n4273;
  assign n4275 = n3519 & ~n4136;
  assign n4276 = n4153 & ~n4275;
  assign n4277 = ~n3317 & n4276;
  assign n4278 = pi62 & ~n4277;
  assign n4279 = ~n4274 & n4278;
  assign n4280 = n2538 & ~n4273;
  assign n4281 = ~n2538 & ~n4276;
  assign n4282 = pi56 & ~n4281;
  assign n4283 = ~n4280 & n4282;
  assign n4284 = ~n2577 & n4276;
  assign n4285 = n2577 & n4273;
  assign n4286 = pi55 & ~n4284;
  assign n4287 = ~n4285 & n4286;
  assign n4288 = ~n3441 & ~n4187;
  assign n4289 = pi299 & ~n4276;
  assign n4290 = n4288 & ~n4289;
  assign n4291 = ~n2533 & n4290;
  assign n4292 = ~n2628 & n4290;
  assign n4293 = pi299 & ~n4273;
  assign n4294 = n4288 & ~n4293;
  assign n4295 = n2628 & n4294;
  assign n4296 = ~n4292 & ~n4295;
  assign n4297 = n2534 & ~n4296;
  assign n4298 = ~n2534 & n4290;
  assign n4299 = pi92 & ~n4298;
  assign n4300 = ~n4297 & n4299;
  assign n4301 = pi75 & n4290;
  assign n4302 = pi87 & n4296;
  assign n4303 = pi38 & n4290;
  assign n4304 = pi39 & ~n4294;
  assign n4305 = ~pi861 & n3466;
  assign n4306 = ~pi171 & ~n4305;
  assign n4307 = pi861 & ~n3392;
  assign n4308 = ~pi861 & ~n3177;
  assign n4309 = pi171 & ~n4308;
  assign n4310 = ~n4307 & n4309;
  assign n4311 = ~n4306 & ~n4310;
  assign n4312 = ~pi228 & ~n4311;
  assign n4313 = ~n3757 & n4143;
  assign n4314 = ~n4312 & n4313;
  assign n4315 = n4137 & ~n4314;
  assign n4316 = ~n4150 & ~n4315;
  assign n4317 = ~pi215 & ~n4316;
  assign n4318 = n4215 & ~n4317;
  assign n4319 = n4214 & ~n4318;
  assign n4320 = ~pi38 & ~n4304;
  assign n4321 = ~n4319 & n4320;
  assign n4322 = ~pi100 & ~n4303;
  assign n4323 = ~n4321 & n4322;
  assign n4324 = ~n2531 & n4290;
  assign n4325 = ~n4240 & n4268;
  assign n4326 = n4137 & ~n4325;
  assign n4327 = ~n4150 & ~n4326;
  assign n4328 = ~pi215 & ~n4327;
  assign n4329 = ~n4135 & ~n4328;
  assign n4330 = pi299 & ~n4329;
  assign n4331 = n2531 & n4288;
  assign n4332 = ~n4330 & n4331;
  assign n4333 = pi100 & ~n4324;
  assign n4334 = ~n4332 & n4333;
  assign n4335 = ~n4323 & ~n4334;
  assign n4336 = ~pi87 & ~n4335;
  assign n4337 = ~pi75 & ~n4302;
  assign n4338 = ~n4336 & n4337;
  assign n4339 = ~pi92 & ~n4301;
  assign n4340 = ~n4338 & n4339;
  assign n4341 = n2533 & ~n4300;
  assign n4342 = ~n4340 & n4341;
  assign n4343 = ~pi55 & ~n4291;
  assign n4344 = ~n4342 & n4343;
  assign n4345 = ~pi56 & ~n4287;
  assign n4346 = ~n4344 & n4345;
  assign n4347 = ~pi62 & ~n4283;
  assign n4348 = ~n4346 & n4347;
  assign n4349 = pi241 & n3291;
  assign n4350 = ~n4279 & n4349;
  assign n4351 = ~n4348 & n4350;
  assign n4352 = pi241 & n4275;
  assign n4353 = ~n3291 & ~n4352;
  assign n4354 = n4153 & n4353;
  assign n4355 = ~n4267 & ~n4354;
  assign po158 = ~n4351 & n4355;
  assign n4357 = pi215 & pi1140;
  assign n4358 = pi216 & pi282;
  assign n4359 = ~pi221 & ~n4358;
  assign n4360 = ~pi105 & pi170;
  assign n4361 = pi869 & ~n2442;
  assign n4362 = pi105 & ~n4361;
  assign n4363 = pi228 & ~n4360;
  assign n4364 = ~n4362 & n4363;
  assign n4365 = ~pi216 & ~n4364;
  assign n4366 = ~pi170 & ~pi228;
  assign n4367 = n4365 & ~n4366;
  assign n4368 = n4359 & ~n4367;
  assign n4369 = ~pi1140 & ~n2452;
  assign n4370 = ~pi921 & n2452;
  assign n4371 = pi221 & ~n4369;
  assign n4372 = ~n4370 & n4371;
  assign n4373 = ~n4368 & ~n4372;
  assign n4374 = ~pi215 & ~n4373;
  assign n4375 = ~n4357 & ~n4374;
  assign n4376 = ~n3317 & n4375;
  assign n4377 = ~pi869 & n2523;
  assign n4378 = pi170 & ~n2523;
  assign n4379 = ~pi228 & ~n4377;
  assign n4380 = ~n4378 & n4379;
  assign n4381 = n4365 & ~n4380;
  assign n4382 = n4359 & ~n4381;
  assign n4383 = ~n4372 & ~n4382;
  assign n4384 = ~pi215 & ~n4383;
  assign n4385 = ~n4357 & ~n4384;
  assign n4386 = n3317 & n4385;
  assign n4387 = pi62 & ~n4376;
  assign n4388 = ~n4386 & n4387;
  assign n4389 = n2538 & ~n4385;
  assign n4390 = ~n2538 & ~n4375;
  assign n4391 = pi56 & ~n4390;
  assign n4392 = ~n4389 & n4391;
  assign n4393 = ~n2577 & n4375;
  assign n4394 = n2577 & n4385;
  assign n4395 = pi55 & ~n4393;
  assign n4396 = ~n4394 & n4395;
  assign n4397 = pi223 & pi1140;
  assign n4398 = pi224 & pi282;
  assign n4399 = ~pi222 & ~n4398;
  assign n4400 = ~pi224 & ~n4361;
  assign n4401 = n4399 & ~n4400;
  assign n4402 = ~pi1140 & ~n2596;
  assign n4403 = ~pi921 & n2596;
  assign n4404 = pi222 & ~n4402;
  assign n4405 = ~n4403 & n4404;
  assign n4406 = ~n4401 & ~n4405;
  assign n4407 = ~pi223 & ~n4406;
  assign n4408 = ~n4397 & ~n4407;
  assign n4409 = ~pi299 & ~n4408;
  assign n4410 = pi299 & ~n4375;
  assign n4411 = ~n4409 & ~n4410;
  assign n4412 = ~n2533 & n4411;
  assign n4413 = ~n2628 & n4411;
  assign n4414 = pi299 & ~n4385;
  assign n4415 = ~n4409 & ~n4414;
  assign n4416 = n2628 & n4415;
  assign n4417 = ~n4413 & ~n4416;
  assign n4418 = n2534 & ~n4417;
  assign n4419 = ~n2534 & n4411;
  assign n4420 = pi92 & ~n4419;
  assign n4421 = ~n4418 & n4420;
  assign n4422 = pi75 & n4411;
  assign n4423 = pi87 & n4417;
  assign n4424 = pi38 & n4411;
  assign n4425 = pi39 & ~n4415;
  assign n4426 = ~pi299 & ~n4397;
  assign n4427 = pi869 & n3176;
  assign n4428 = ~pi224 & ~n4427;
  assign n4429 = n4399 & ~n4428;
  assign n4430 = ~n4405 & ~n4429;
  assign n4431 = n4426 & n4430;
  assign n4432 = ~n3176 & n4399;
  assign n4433 = n4430 & ~n4432;
  assign n4434 = ~pi223 & ~n4433;
  assign n4435 = n4426 & ~n4434;
  assign n4436 = ~pi39 & ~n4435;
  assign n4437 = pi299 & ~n4357;
  assign n4438 = ~pi869 & n3391;
  assign n4439 = ~n2740 & ~n4427;
  assign n4440 = ~n4438 & n4439;
  assign n4441 = ~pi170 & ~n4440;
  assign n4442 = pi170 & pi869;
  assign n4443 = n3466 & n4442;
  assign n4444 = ~n4441 & ~n4443;
  assign n4445 = ~pi228 & ~n4444;
  assign n4446 = ~n3471 & n4364;
  assign n4447 = ~pi216 & ~n4446;
  assign n4448 = ~n4445 & n4447;
  assign n4449 = n4359 & ~n4448;
  assign n4450 = ~n4372 & ~n4449;
  assign n4451 = ~pi215 & ~n4450;
  assign n4452 = n4437 & ~n4451;
  assign n4453 = ~n4431 & n4436;
  assign n4454 = ~n4452 & n4453;
  assign n4455 = ~pi38 & ~n4425;
  assign n4456 = ~n4454 & n4455;
  assign n4457 = ~pi100 & ~n4424;
  assign n4458 = ~n4456 & n4457;
  assign n4459 = ~n2531 & n4411;
  assign n4460 = ~pi869 & n3371;
  assign n4461 = ~n3593 & ~n4366;
  assign n4462 = ~n4460 & ~n4461;
  assign n4463 = n4365 & ~n4462;
  assign n4464 = n4359 & ~n4463;
  assign n4465 = ~n4372 & ~n4464;
  assign n4466 = ~pi215 & ~n4465;
  assign n4467 = ~n4357 & ~n4466;
  assign n4468 = pi299 & ~n4467;
  assign n4469 = n2531 & ~n4409;
  assign n4470 = ~n4468 & n4469;
  assign n4471 = pi100 & ~n4459;
  assign n4472 = ~n4470 & n4471;
  assign n4473 = ~n4458 & ~n4472;
  assign n4474 = ~pi87 & ~n4473;
  assign n4475 = ~pi75 & ~n4423;
  assign n4476 = ~n4474 & n4475;
  assign n4477 = ~pi92 & ~n4422;
  assign n4478 = ~n4476 & n4477;
  assign n4479 = n2533 & ~n4421;
  assign n4480 = ~n4478 & n4479;
  assign n4481 = ~pi55 & ~n4412;
  assign n4482 = ~n4480 & n4481;
  assign n4483 = ~pi56 & ~n4396;
  assign n4484 = ~n4482 & n4483;
  assign n4485 = ~pi62 & ~n4392;
  assign n4486 = ~n4484 & n4485;
  assign n4487 = ~pi248 & n3291;
  assign n4488 = ~n4388 & n4487;
  assign n4489 = ~n4486 & n4488;
  assign n4490 = ~n3421 & n4365;
  assign n4491 = ~n4380 & n4490;
  assign n4492 = n4359 & ~n4491;
  assign n4493 = ~n4372 & ~n4492;
  assign n4494 = ~pi215 & ~n4493;
  assign n4495 = ~n4357 & ~n4494;
  assign n4496 = n3317 & n4495;
  assign n4497 = n3519 & ~n4358;
  assign n4498 = n4375 & ~n4497;
  assign n4499 = ~n3317 & n4498;
  assign n4500 = pi62 & ~n4499;
  assign n4501 = ~n4496 & n4500;
  assign n4502 = n2538 & ~n4495;
  assign n4503 = ~n2538 & ~n4498;
  assign n4504 = pi56 & ~n4503;
  assign n4505 = ~n4502 & n4504;
  assign n4506 = ~n2577 & n4498;
  assign n4507 = n2577 & n4495;
  assign n4508 = pi55 & ~n4506;
  assign n4509 = ~n4507 & n4508;
  assign n4510 = ~n3441 & ~n4409;
  assign n4511 = pi299 & ~n4498;
  assign n4512 = n4510 & ~n4511;
  assign n4513 = ~n2533 & n4512;
  assign n4514 = ~n2628 & n4512;
  assign n4515 = pi299 & ~n4495;
  assign n4516 = n4510 & ~n4515;
  assign n4517 = n2628 & n4516;
  assign n4518 = ~n4514 & ~n4517;
  assign n4519 = n2534 & ~n4518;
  assign n4520 = ~n2534 & n4512;
  assign n4521 = pi92 & ~n4520;
  assign n4522 = ~n4519 & n4521;
  assign n4523 = pi75 & n4512;
  assign n4524 = pi87 & n4518;
  assign n4525 = pi38 & n4512;
  assign n4526 = pi39 & ~n4516;
  assign n4527 = ~pi869 & n3466;
  assign n4528 = ~pi170 & ~n4527;
  assign n4529 = pi869 & ~n3392;
  assign n4530 = ~pi869 & ~n3177;
  assign n4531 = pi170 & ~n4530;
  assign n4532 = ~n4529 & n4531;
  assign n4533 = ~n4528 & ~n4532;
  assign n4534 = ~pi228 & ~n4533;
  assign n4535 = ~n3757 & n4365;
  assign n4536 = ~n4534 & n4535;
  assign n4537 = n4359 & ~n4536;
  assign n4538 = ~n4372 & ~n4537;
  assign n4539 = ~pi215 & ~n4538;
  assign n4540 = n4437 & ~n4539;
  assign n4541 = n4436 & ~n4540;
  assign n4542 = ~pi38 & ~n4526;
  assign n4543 = ~n4541 & n4542;
  assign n4544 = ~pi100 & ~n4525;
  assign n4545 = ~n4543 & n4544;
  assign n4546 = ~n2531 & n4512;
  assign n4547 = ~n4462 & n4490;
  assign n4548 = n4359 & ~n4547;
  assign n4549 = ~n4372 & ~n4548;
  assign n4550 = ~pi215 & ~n4549;
  assign n4551 = ~n4357 & ~n4550;
  assign n4552 = pi299 & ~n4551;
  assign n4553 = n2531 & n4510;
  assign n4554 = ~n4552 & n4553;
  assign n4555 = pi100 & ~n4546;
  assign n4556 = ~n4554 & n4555;
  assign n4557 = ~n4545 & ~n4556;
  assign n4558 = ~pi87 & ~n4557;
  assign n4559 = ~pi75 & ~n4524;
  assign n4560 = ~n4558 & n4559;
  assign n4561 = ~pi92 & ~n4523;
  assign n4562 = ~n4560 & n4561;
  assign n4563 = n2533 & ~n4522;
  assign n4564 = ~n4562 & n4563;
  assign n4565 = ~pi55 & ~n4513;
  assign n4566 = ~n4564 & n4565;
  assign n4567 = ~pi56 & ~n4509;
  assign n4568 = ~n4566 & n4567;
  assign n4569 = ~pi62 & ~n4505;
  assign n4570 = ~n4568 & n4569;
  assign n4571 = pi248 & n3291;
  assign n4572 = ~n4501 & n4571;
  assign n4573 = ~n4570 & n4572;
  assign n4574 = pi248 & n4497;
  assign n4575 = ~n3291 & ~n4574;
  assign n4576 = n4375 & n4575;
  assign n4577 = ~n4489 & ~n4576;
  assign po159 = ~n4573 & n4577;
  assign n4579 = pi215 & pi1139;
  assign n4580 = pi216 & pi281;
  assign n4581 = ~pi221 & ~n4580;
  assign n4582 = ~pi216 & ~pi862;
  assign n4583 = n3594 & n4582;
  assign n4584 = n4581 & ~n4583;
  assign n4585 = ~pi1139 & ~n2452;
  assign n4586 = ~pi920 & n2452;
  assign n4587 = pi221 & ~n4585;
  assign n4588 = ~n4586 & n4587;
  assign n4589 = ~n4584 & ~n4588;
  assign n4590 = ~pi216 & ~n4588;
  assign n4591 = pi148 & ~n2441;
  assign n4592 = n4590 & n4591;
  assign n4593 = ~pi215 & ~n4592;
  assign n4594 = ~n4589 & n4593;
  assign n4595 = ~n4579 & ~n4594;
  assign n4596 = ~n3422 & ~n4595;
  assign n4597 = ~n3291 & ~n4596;
  assign n4598 = ~pi148 & ~pi215;
  assign n4599 = ~n2441 & ~n3524;
  assign n4600 = pi862 & ~n3421;
  assign n4601 = ~pi216 & ~n4600;
  assign n4602 = ~n4599 & n4601;
  assign n4603 = n4581 & ~n4602;
  assign n4604 = ~n4588 & ~n4603;
  assign n4605 = n4598 & ~n4604;
  assign n4606 = ~n3524 & ~n3594;
  assign n4607 = n4590 & n4606;
  assign n4608 = n4582 & ~n4606;
  assign n4609 = n4581 & ~n4608;
  assign n4610 = ~n4588 & ~n4609;
  assign n4611 = pi148 & ~pi215;
  assign n4612 = ~n4610 & n4611;
  assign n4613 = ~n4607 & n4612;
  assign n4614 = ~n4579 & ~n4613;
  assign n4615 = ~n4605 & n4614;
  assign n4616 = n2538 & ~n4615;
  assign n4617 = ~pi56 & n4616;
  assign n4618 = ~n3317 & n4596;
  assign n4619 = ~n4617 & ~n4618;
  assign n4620 = pi62 & ~n4619;
  assign n4621 = ~n2538 & n4596;
  assign n4622 = pi56 & ~n4621;
  assign n4623 = ~n4616 & n4622;
  assign n4624 = ~n2577 & ~n4596;
  assign n4625 = n2577 & n4615;
  assign n4626 = pi55 & ~n4624;
  assign n4627 = ~n4625 & n4626;
  assign n4628 = pi223 & pi1139;
  assign n4629 = ~pi1139 & ~n2596;
  assign n4630 = ~pi920 & n2596;
  assign n4631 = pi222 & ~n4629;
  assign n4632 = ~n4630 & n4631;
  assign n4633 = ~pi224 & ~n4628;
  assign n4634 = ~n4632 & n4633;
  assign n4635 = ~pi862 & n4634;
  assign n4636 = pi224 & pi281;
  assign n4637 = ~pi222 & ~n4636;
  assign n4638 = ~n4632 & ~n4637;
  assign n4639 = ~pi223 & ~n4638;
  assign n4640 = ~n4628 & ~n4639;
  assign n4641 = ~pi299 & ~n4640;
  assign n4642 = ~n4635 & n4641;
  assign n4643 = ~n3440 & n4642;
  assign n4644 = pi299 & n4596;
  assign n4645 = ~n4643 & ~n4644;
  assign n4646 = ~n2533 & n4645;
  assign n4647 = ~n2628 & n4645;
  assign n4648 = pi299 & ~n4615;
  assign n4649 = ~n4643 & ~n4648;
  assign n4650 = n2628 & n4649;
  assign n4651 = ~n4647 & ~n4650;
  assign n4652 = n2534 & ~n4651;
  assign n4653 = ~n2534 & n4645;
  assign n4654 = pi92 & ~n4653;
  assign n4655 = ~n4652 & n4654;
  assign n4656 = pi75 & n4645;
  assign n4657 = pi87 & n4651;
  assign n4658 = ~n2531 & n4645;
  assign n4659 = ~n2441 & ~n3593;
  assign n4660 = n4581 & n4659;
  assign n4661 = n4604 & ~n4660;
  assign n4662 = n4598 & ~n4661;
  assign n4663 = n3595 & n4590;
  assign n4664 = n4612 & ~n4663;
  assign n4665 = ~n4579 & ~n4664;
  assign n4666 = ~n4662 & n4665;
  assign n4667 = pi299 & ~n4666;
  assign n4668 = n2531 & ~n4643;
  assign n4669 = ~n4667 & n4668;
  assign n4670 = pi100 & ~n4658;
  assign n4671 = ~n4669 & n4670;
  assign n4672 = pi38 & n4645;
  assign n4673 = pi39 & ~n4649;
  assign n4674 = ~n3176 & n4634;
  assign n4675 = ~n4635 & ~n4640;
  assign n4676 = ~n4674 & n4675;
  assign n4677 = ~pi299 & ~n4676;
  assign n4678 = n3469 & n4590;
  assign n4679 = ~n3469 & n4582;
  assign n4680 = n4581 & ~n4679;
  assign n4681 = ~n4588 & ~n4680;
  assign n4682 = n4611 & ~n4678;
  assign n4683 = ~n4681 & n4682;
  assign n4684 = pi862 & ~n3474;
  assign n4685 = ~pi228 & n3392;
  assign n4686 = ~n2441 & ~n4685;
  assign n4687 = ~pi862 & n4686;
  assign n4688 = ~pi216 & ~n4684;
  assign n4689 = ~n4687 & n4688;
  assign n4690 = n4581 & ~n4689;
  assign n4691 = ~n4588 & ~n4690;
  assign n4692 = n4598 & ~n4691;
  assign n4693 = pi299 & ~n4579;
  assign n4694 = ~n4683 & n4693;
  assign n4695 = ~n4692 & n4694;
  assign n4696 = ~pi39 & ~n4677;
  assign n4697 = ~n4695 & n4696;
  assign n4698 = ~pi38 & ~n4673;
  assign n4699 = ~n4697 & n4698;
  assign n4700 = ~pi100 & ~n4672;
  assign n4701 = ~n4699 & n4700;
  assign n4702 = ~n4671 & ~n4701;
  assign n4703 = ~pi87 & ~n4702;
  assign n4704 = ~pi75 & ~n4657;
  assign n4705 = ~n4703 & n4704;
  assign n4706 = ~pi92 & ~n4656;
  assign n4707 = ~n4705 & n4706;
  assign n4708 = n2533 & ~n4655;
  assign n4709 = ~n4707 & n4708;
  assign n4710 = ~pi55 & ~n4646;
  assign n4711 = ~n4709 & n4710;
  assign n4712 = ~pi56 & ~n4627;
  assign n4713 = ~n4711 & n4712;
  assign n4714 = ~pi62 & ~n4623;
  assign n4715 = ~n4713 & n4714;
  assign n4716 = n3291 & ~n4620;
  assign n4717 = ~n4715 & n4716;
  assign n4718 = ~pi247 & ~n4597;
  assign n4719 = ~n4717 & n4718;
  assign n4720 = ~n3291 & n4595;
  assign n4721 = ~n3317 & ~n4595;
  assign n4722 = n4593 & ~n4610;
  assign n4723 = n4614 & ~n4722;
  assign n4724 = n2538 & ~n4723;
  assign n4725 = ~pi56 & n4724;
  assign n4726 = ~n4721 & ~n4725;
  assign n4727 = pi62 & ~n4726;
  assign n4728 = ~n2538 & ~n4595;
  assign n4729 = pi56 & ~n4728;
  assign n4730 = ~n4724 & n4729;
  assign n4731 = ~n2577 & n4595;
  assign n4732 = n2577 & n4723;
  assign n4733 = pi55 & ~n4731;
  assign n4734 = ~n4732 & n4733;
  assign n4735 = ~n3441 & ~n4642;
  assign n4736 = pi299 & ~n4595;
  assign n4737 = n4735 & ~n4736;
  assign n4738 = ~n2533 & n4737;
  assign n4739 = ~n2628 & n4737;
  assign n4740 = pi299 & ~n4723;
  assign n4741 = n4735 & ~n4740;
  assign n4742 = n2628 & n4741;
  assign n4743 = ~n4739 & ~n4742;
  assign n4744 = n2534 & ~n4743;
  assign n4745 = ~n2534 & n4737;
  assign n4746 = pi92 & ~n4745;
  assign n4747 = ~n4744 & n4746;
  assign n4748 = pi75 & n4737;
  assign n4749 = pi87 & n4743;
  assign n4750 = ~n2531 & n4737;
  assign n4751 = n3595 & n4581;
  assign n4752 = n4610 & ~n4751;
  assign n4753 = n4598 & ~n4752;
  assign n4754 = n4590 & n4659;
  assign n4755 = n4612 & ~n4754;
  assign n4756 = ~n4579 & ~n4755;
  assign n4757 = ~n4753 & n4756;
  assign n4758 = pi299 & ~n4757;
  assign n4759 = n2531 & n4735;
  assign n4760 = ~n4758 & n4759;
  assign n4761 = pi100 & ~n4750;
  assign n4762 = ~n4760 & n4761;
  assign n4763 = pi38 & n4737;
  assign n4764 = pi39 & ~n4741;
  assign n4765 = n3176 & n4635;
  assign n4766 = n4641 & ~n4765;
  assign n4767 = pi862 & ~n4686;
  assign n4768 = ~pi862 & n3474;
  assign n4769 = ~pi216 & ~n4768;
  assign n4770 = ~n4767 & n4769;
  assign n4771 = n4581 & ~n4770;
  assign n4772 = ~n4588 & ~n4771;
  assign n4773 = n4611 & ~n4772;
  assign n4774 = n4598 & ~n4681;
  assign n4775 = ~n4579 & ~n4774;
  assign n4776 = ~n4773 & n4775;
  assign n4777 = pi299 & ~n4776;
  assign n4778 = ~n4766 & ~n4777;
  assign n4779 = ~pi39 & ~n4778;
  assign n4780 = ~pi38 & ~n4764;
  assign n4781 = ~n4779 & n4780;
  assign n4782 = ~pi100 & ~n4763;
  assign n4783 = ~n4781 & n4782;
  assign n4784 = ~n4762 & ~n4783;
  assign n4785 = ~pi87 & ~n4784;
  assign n4786 = ~pi75 & ~n4749;
  assign n4787 = ~n4785 & n4786;
  assign n4788 = ~pi92 & ~n4748;
  assign n4789 = ~n4787 & n4788;
  assign n4790 = n2533 & ~n4747;
  assign n4791 = ~n4789 & n4790;
  assign n4792 = ~pi55 & ~n4738;
  assign n4793 = ~n4791 & n4792;
  assign n4794 = ~pi56 & ~n4734;
  assign n4795 = ~n4793 & n4794;
  assign n4796 = ~pi62 & ~n4730;
  assign n4797 = ~n4795 & n4796;
  assign n4798 = n3291 & ~n4727;
  assign n4799 = ~n4797 & n4798;
  assign n4800 = pi247 & ~n4720;
  assign n4801 = ~n4799 & n4800;
  assign po160 = n4719 | n4801;
  assign n4803 = pi215 & pi1138;
  assign n4804 = pi216 & pi269;
  assign n4805 = ~pi221 & ~n4804;
  assign n4806 = ~pi105 & pi169;
  assign n4807 = pi877 & ~n2442;
  assign n4808 = pi105 & ~n4807;
  assign n4809 = pi228 & ~n4806;
  assign n4810 = ~n4808 & n4809;
  assign n4811 = ~pi216 & ~n4810;
  assign n4812 = ~pi169 & ~pi228;
  assign n4813 = n4811 & ~n4812;
  assign n4814 = n4805 & ~n4813;
  assign n4815 = ~pi1138 & ~n2452;
  assign n4816 = ~pi940 & n2452;
  assign n4817 = pi221 & ~n4815;
  assign n4818 = ~n4816 & n4817;
  assign n4819 = ~n4814 & ~n4818;
  assign n4820 = ~pi215 & ~n4819;
  assign n4821 = ~n4803 & ~n4820;
  assign n4822 = ~n3317 & n4821;
  assign n4823 = ~pi877 & n2523;
  assign n4824 = ~n3524 & ~n4812;
  assign n4825 = ~n4823 & ~n4824;
  assign n4826 = n4811 & ~n4825;
  assign n4827 = n4805 & ~n4826;
  assign n4828 = ~n4818 & ~n4827;
  assign n4829 = ~pi215 & ~n4828;
  assign n4830 = ~n4803 & ~n4829;
  assign n4831 = n3317 & n4830;
  assign n4832 = pi62 & ~n4822;
  assign n4833 = ~n4831 & n4832;
  assign n4834 = n2538 & ~n4830;
  assign n4835 = ~n2538 & ~n4821;
  assign n4836 = pi56 & ~n4835;
  assign n4837 = ~n4834 & n4836;
  assign n4838 = ~n2577 & n4821;
  assign n4839 = n2577 & n4830;
  assign n4840 = pi55 & ~n4838;
  assign n4841 = ~n4839 & n4840;
  assign n4842 = pi223 & pi1138;
  assign n4843 = pi224 & pi269;
  assign n4844 = ~pi222 & ~n4843;
  assign n4845 = ~pi224 & ~n4807;
  assign n4846 = n4844 & ~n4845;
  assign n4847 = ~pi1138 & ~n2596;
  assign n4848 = ~pi940 & n2596;
  assign n4849 = pi222 & ~n4847;
  assign n4850 = ~n4848 & n4849;
  assign n4851 = ~n4846 & ~n4850;
  assign n4852 = ~pi223 & ~n4851;
  assign n4853 = ~n4842 & ~n4852;
  assign n4854 = ~pi299 & ~n4853;
  assign n4855 = pi299 & ~n4821;
  assign n4856 = ~n4854 & ~n4855;
  assign n4857 = ~n2533 & n4856;
  assign n4858 = ~n2628 & n4856;
  assign n4859 = pi299 & ~n4830;
  assign n4860 = ~n4854 & ~n4859;
  assign n4861 = n2628 & n4860;
  assign n4862 = ~n4858 & ~n4861;
  assign n4863 = n2534 & ~n4862;
  assign n4864 = ~n2534 & n4856;
  assign n4865 = pi92 & ~n4864;
  assign n4866 = ~n4863 & n4865;
  assign n4867 = pi75 & n4856;
  assign n4868 = pi87 & n4862;
  assign n4869 = pi38 & n4856;
  assign n4870 = pi39 & ~n4860;
  assign n4871 = ~pi299 & ~n4842;
  assign n4872 = pi877 & n3176;
  assign n4873 = ~pi224 & ~n4872;
  assign n4874 = n4844 & ~n4873;
  assign n4875 = ~n4850 & ~n4874;
  assign n4876 = n4871 & n4875;
  assign n4877 = ~n3176 & n4844;
  assign n4878 = n4875 & ~n4877;
  assign n4879 = ~pi223 & ~n4878;
  assign n4880 = n4871 & ~n4879;
  assign n4881 = ~pi39 & ~n4880;
  assign n4882 = pi299 & ~n4803;
  assign n4883 = ~pi877 & n3391;
  assign n4884 = ~n2740 & ~n4872;
  assign n4885 = ~n4883 & n4884;
  assign n4886 = ~pi169 & ~n4885;
  assign n4887 = pi169 & pi877;
  assign n4888 = n3466 & n4887;
  assign n4889 = ~n4886 & ~n4888;
  assign n4890 = ~pi228 & ~n4889;
  assign n4891 = ~n3471 & n4810;
  assign n4892 = ~pi216 & ~n4891;
  assign n4893 = ~n4890 & n4892;
  assign n4894 = n4805 & ~n4893;
  assign n4895 = ~n4818 & ~n4894;
  assign n4896 = ~pi215 & ~n4895;
  assign n4897 = n4882 & ~n4896;
  assign n4898 = ~n4876 & n4881;
  assign n4899 = ~n4897 & n4898;
  assign n4900 = ~pi38 & ~n4870;
  assign n4901 = ~n4899 & n4900;
  assign n4902 = ~pi100 & ~n4869;
  assign n4903 = ~n4901 & n4902;
  assign n4904 = ~n2531 & n4856;
  assign n4905 = ~pi877 & n3371;
  assign n4906 = ~n3593 & ~n4812;
  assign n4907 = ~n4905 & ~n4906;
  assign n4908 = n4811 & ~n4907;
  assign n4909 = n4805 & ~n4908;
  assign n4910 = ~n4818 & ~n4909;
  assign n4911 = ~pi215 & ~n4910;
  assign n4912 = ~n4803 & ~n4911;
  assign n4913 = pi299 & ~n4912;
  assign n4914 = n2531 & ~n4854;
  assign n4915 = ~n4913 & n4914;
  assign n4916 = pi100 & ~n4904;
  assign n4917 = ~n4915 & n4916;
  assign n4918 = ~n4903 & ~n4917;
  assign n4919 = ~pi87 & ~n4918;
  assign n4920 = ~pi75 & ~n4868;
  assign n4921 = ~n4919 & n4920;
  assign n4922 = ~pi92 & ~n4867;
  assign n4923 = ~n4921 & n4922;
  assign n4924 = n2533 & ~n4866;
  assign n4925 = ~n4923 & n4924;
  assign n4926 = ~pi55 & ~n4857;
  assign n4927 = ~n4925 & n4926;
  assign n4928 = ~pi56 & ~n4841;
  assign n4929 = ~n4927 & n4928;
  assign n4930 = ~pi62 & ~n4837;
  assign n4931 = ~n4929 & n4930;
  assign n4932 = ~pi246 & n3291;
  assign n4933 = ~n4833 & n4932;
  assign n4934 = ~n4931 & n4933;
  assign n4935 = ~n3421 & n4811;
  assign n4936 = ~n4825 & n4935;
  assign n4937 = n4805 & ~n4936;
  assign n4938 = ~n4818 & ~n4937;
  assign n4939 = ~pi215 & ~n4938;
  assign n4940 = ~n4803 & ~n4939;
  assign n4941 = n3317 & n4940;
  assign n4942 = n3519 & ~n4804;
  assign n4943 = n4821 & ~n4942;
  assign n4944 = ~n3317 & n4943;
  assign n4945 = pi62 & ~n4944;
  assign n4946 = ~n4941 & n4945;
  assign n4947 = n2538 & ~n4940;
  assign n4948 = ~n2538 & ~n4943;
  assign n4949 = pi56 & ~n4948;
  assign n4950 = ~n4947 & n4949;
  assign n4951 = ~n2577 & n4943;
  assign n4952 = n2577 & n4940;
  assign n4953 = pi55 & ~n4951;
  assign n4954 = ~n4952 & n4953;
  assign n4955 = ~n3441 & ~n4854;
  assign n4956 = pi299 & ~n4943;
  assign n4957 = n4955 & ~n4956;
  assign n4958 = ~n2533 & n4957;
  assign n4959 = ~n2628 & n4957;
  assign n4960 = pi299 & ~n4940;
  assign n4961 = n4955 & ~n4960;
  assign n4962 = n2628 & n4961;
  assign n4963 = ~n4959 & ~n4962;
  assign n4964 = n2534 & ~n4963;
  assign n4965 = ~n2534 & n4957;
  assign n4966 = pi92 & ~n4965;
  assign n4967 = ~n4964 & n4966;
  assign n4968 = pi75 & n4957;
  assign n4969 = pi87 & n4963;
  assign n4970 = pi38 & n4957;
  assign n4971 = pi39 & ~n4961;
  assign n4972 = ~pi877 & n3466;
  assign n4973 = ~pi169 & ~n4972;
  assign n4974 = pi877 & ~n3392;
  assign n4975 = ~pi877 & ~n3177;
  assign n4976 = pi169 & ~n4975;
  assign n4977 = ~n4974 & n4976;
  assign n4978 = ~n4973 & ~n4977;
  assign n4979 = ~pi228 & ~n4978;
  assign n4980 = ~n3757 & n4811;
  assign n4981 = ~n4979 & n4980;
  assign n4982 = n4805 & ~n4981;
  assign n4983 = ~n4818 & ~n4982;
  assign n4984 = ~pi215 & ~n4983;
  assign n4985 = n4882 & ~n4984;
  assign n4986 = n4881 & ~n4985;
  assign n4987 = ~pi38 & ~n4971;
  assign n4988 = ~n4986 & n4987;
  assign n4989 = ~pi100 & ~n4970;
  assign n4990 = ~n4988 & n4989;
  assign n4991 = ~n2531 & n4957;
  assign n4992 = ~n4907 & n4935;
  assign n4993 = n4805 & ~n4992;
  assign n4994 = ~n4818 & ~n4993;
  assign n4995 = ~pi215 & ~n4994;
  assign n4996 = ~n4803 & ~n4995;
  assign n4997 = pi299 & ~n4996;
  assign n4998 = n2531 & n4955;
  assign n4999 = ~n4997 & n4998;
  assign n5000 = pi100 & ~n4991;
  assign n5001 = ~n4999 & n5000;
  assign n5002 = ~n4990 & ~n5001;
  assign n5003 = ~pi87 & ~n5002;
  assign n5004 = ~pi75 & ~n4969;
  assign n5005 = ~n5003 & n5004;
  assign n5006 = ~pi92 & ~n4968;
  assign n5007 = ~n5005 & n5006;
  assign n5008 = n2533 & ~n4967;
  assign n5009 = ~n5007 & n5008;
  assign n5010 = ~pi55 & ~n4958;
  assign n5011 = ~n5009 & n5010;
  assign n5012 = ~pi56 & ~n4954;
  assign n5013 = ~n5011 & n5012;
  assign n5014 = ~pi62 & ~n4950;
  assign n5015 = ~n5013 & n5014;
  assign n5016 = pi246 & n3291;
  assign n5017 = ~n4946 & n5016;
  assign n5018 = ~n5015 & n5017;
  assign n5019 = pi246 & n4942;
  assign n5020 = ~n3291 & ~n5019;
  assign n5021 = n4821 & n5020;
  assign n5022 = ~n4934 & ~n5021;
  assign po161 = ~n5018 & n5022;
  assign n5024 = pi215 & pi1137;
  assign n5025 = pi216 & pi280;
  assign n5026 = ~pi221 & ~n5025;
  assign n5027 = ~pi105 & pi168;
  assign n5028 = pi878 & ~n2442;
  assign n5029 = pi105 & ~n5028;
  assign n5030 = pi228 & ~n5027;
  assign n5031 = ~n5029 & n5030;
  assign n5032 = ~pi216 & ~n5031;
  assign n5033 = ~pi168 & ~pi228;
  assign n5034 = n5032 & ~n5033;
  assign n5035 = n5026 & ~n5034;
  assign n5036 = ~pi1137 & ~n2452;
  assign n5037 = ~pi933 & n2452;
  assign n5038 = pi221 & ~n5036;
  assign n5039 = ~n5037 & n5038;
  assign n5040 = ~n5035 & ~n5039;
  assign n5041 = ~pi215 & ~n5040;
  assign n5042 = ~n5024 & ~n5041;
  assign n5043 = ~n3317 & n5042;
  assign n5044 = ~pi878 & n2523;
  assign n5045 = ~n3524 & ~n5033;
  assign n5046 = ~n5044 & ~n5045;
  assign n5047 = n5032 & ~n5046;
  assign n5048 = n5026 & ~n5047;
  assign n5049 = ~n5039 & ~n5048;
  assign n5050 = ~pi215 & ~n5049;
  assign n5051 = ~n5024 & ~n5050;
  assign n5052 = n3317 & n5051;
  assign n5053 = pi62 & ~n5043;
  assign n5054 = ~n5052 & n5053;
  assign n5055 = n2538 & ~n5051;
  assign n5056 = ~n2538 & ~n5042;
  assign n5057 = pi56 & ~n5056;
  assign n5058 = ~n5055 & n5057;
  assign n5059 = ~n2577 & n5042;
  assign n5060 = n2577 & n5051;
  assign n5061 = pi55 & ~n5059;
  assign n5062 = ~n5060 & n5061;
  assign n5063 = pi223 & pi1137;
  assign n5064 = pi224 & pi280;
  assign n5065 = ~pi222 & ~n5064;
  assign n5066 = ~pi224 & ~n5028;
  assign n5067 = n5065 & ~n5066;
  assign n5068 = ~pi1137 & ~n2596;
  assign n5069 = ~pi933 & n2596;
  assign n5070 = pi222 & ~n5068;
  assign n5071 = ~n5069 & n5070;
  assign n5072 = ~n5067 & ~n5071;
  assign n5073 = ~pi223 & ~n5072;
  assign n5074 = ~n5063 & ~n5073;
  assign n5075 = ~pi299 & ~n5074;
  assign n5076 = pi299 & ~n5042;
  assign n5077 = ~n5075 & ~n5076;
  assign n5078 = ~n2533 & n5077;
  assign n5079 = ~n2628 & n5077;
  assign n5080 = pi299 & ~n5051;
  assign n5081 = ~n5075 & ~n5080;
  assign n5082 = n2628 & n5081;
  assign n5083 = ~n5079 & ~n5082;
  assign n5084 = n2534 & ~n5083;
  assign n5085 = ~n2534 & n5077;
  assign n5086 = pi92 & ~n5085;
  assign n5087 = ~n5084 & n5086;
  assign n5088 = pi75 & n5077;
  assign n5089 = pi87 & n5083;
  assign n5090 = pi38 & n5077;
  assign n5091 = pi39 & ~n5081;
  assign n5092 = ~pi299 & ~n5063;
  assign n5093 = pi878 & n3176;
  assign n5094 = ~pi224 & ~n5093;
  assign n5095 = n5065 & ~n5094;
  assign n5096 = ~n5071 & ~n5095;
  assign n5097 = n5092 & n5096;
  assign n5098 = ~n3176 & n5065;
  assign n5099 = n5096 & ~n5098;
  assign n5100 = ~pi223 & ~n5099;
  assign n5101 = n5092 & ~n5100;
  assign n5102 = ~pi39 & ~n5101;
  assign n5103 = pi299 & ~n5024;
  assign n5104 = ~pi878 & n3391;
  assign n5105 = ~n2740 & ~n5093;
  assign n5106 = ~n5104 & n5105;
  assign n5107 = ~pi168 & ~n5106;
  assign n5108 = pi168 & pi878;
  assign n5109 = n3466 & n5108;
  assign n5110 = ~n5107 & ~n5109;
  assign n5111 = ~pi228 & ~n5110;
  assign n5112 = ~n3471 & n5031;
  assign n5113 = ~pi216 & ~n5112;
  assign n5114 = ~n5111 & n5113;
  assign n5115 = n5026 & ~n5114;
  assign n5116 = ~n5039 & ~n5115;
  assign n5117 = ~pi215 & ~n5116;
  assign n5118 = n5103 & ~n5117;
  assign n5119 = ~n5097 & n5102;
  assign n5120 = ~n5118 & n5119;
  assign n5121 = ~pi38 & ~n5091;
  assign n5122 = ~n5120 & n5121;
  assign n5123 = ~pi100 & ~n5090;
  assign n5124 = ~n5122 & n5123;
  assign n5125 = ~n2531 & n5077;
  assign n5126 = ~pi878 & n3371;
  assign n5127 = ~n3593 & ~n5033;
  assign n5128 = ~n5126 & ~n5127;
  assign n5129 = n5032 & ~n5128;
  assign n5130 = n5026 & ~n5129;
  assign n5131 = ~n5039 & ~n5130;
  assign n5132 = ~pi215 & ~n5131;
  assign n5133 = ~n5024 & ~n5132;
  assign n5134 = pi299 & ~n5133;
  assign n5135 = n2531 & ~n5075;
  assign n5136 = ~n5134 & n5135;
  assign n5137 = pi100 & ~n5125;
  assign n5138 = ~n5136 & n5137;
  assign n5139 = ~n5124 & ~n5138;
  assign n5140 = ~pi87 & ~n5139;
  assign n5141 = ~pi75 & ~n5089;
  assign n5142 = ~n5140 & n5141;
  assign n5143 = ~pi92 & ~n5088;
  assign n5144 = ~n5142 & n5143;
  assign n5145 = n2533 & ~n5087;
  assign n5146 = ~n5144 & n5145;
  assign n5147 = ~pi55 & ~n5078;
  assign n5148 = ~n5146 & n5147;
  assign n5149 = ~pi56 & ~n5062;
  assign n5150 = ~n5148 & n5149;
  assign n5151 = ~pi62 & ~n5058;
  assign n5152 = ~n5150 & n5151;
  assign n5153 = ~pi240 & n3291;
  assign n5154 = ~n5054 & n5153;
  assign n5155 = ~n5152 & n5154;
  assign n5156 = ~n3421 & n5032;
  assign n5157 = ~n5046 & n5156;
  assign n5158 = n5026 & ~n5157;
  assign n5159 = ~n5039 & ~n5158;
  assign n5160 = ~pi215 & ~n5159;
  assign n5161 = ~n5024 & ~n5160;
  assign n5162 = n3317 & n5161;
  assign n5163 = n3519 & ~n5025;
  assign n5164 = n5042 & ~n5163;
  assign n5165 = ~n3317 & n5164;
  assign n5166 = pi62 & ~n5165;
  assign n5167 = ~n5162 & n5166;
  assign n5168 = n2538 & ~n5161;
  assign n5169 = ~n2538 & ~n5164;
  assign n5170 = pi56 & ~n5169;
  assign n5171 = ~n5168 & n5170;
  assign n5172 = ~n2577 & n5164;
  assign n5173 = n2577 & n5161;
  assign n5174 = pi55 & ~n5172;
  assign n5175 = ~n5173 & n5174;
  assign n5176 = ~n3441 & ~n5075;
  assign n5177 = pi299 & ~n5164;
  assign n5178 = n5176 & ~n5177;
  assign n5179 = ~n2533 & n5178;
  assign n5180 = ~n2628 & n5178;
  assign n5181 = pi299 & ~n5161;
  assign n5182 = n5176 & ~n5181;
  assign n5183 = n2628 & n5182;
  assign n5184 = ~n5180 & ~n5183;
  assign n5185 = n2534 & ~n5184;
  assign n5186 = ~n2534 & n5178;
  assign n5187 = pi92 & ~n5186;
  assign n5188 = ~n5185 & n5187;
  assign n5189 = pi75 & n5178;
  assign n5190 = pi87 & n5184;
  assign n5191 = pi38 & n5178;
  assign n5192 = pi39 & ~n5182;
  assign n5193 = ~pi878 & n3466;
  assign n5194 = ~pi168 & ~n5193;
  assign n5195 = pi878 & ~n3392;
  assign n5196 = ~pi878 & ~n3177;
  assign n5197 = pi168 & ~n5196;
  assign n5198 = ~n5195 & n5197;
  assign n5199 = ~n5194 & ~n5198;
  assign n5200 = ~pi228 & ~n5199;
  assign n5201 = ~n3757 & n5032;
  assign n5202 = ~n5200 & n5201;
  assign n5203 = n5026 & ~n5202;
  assign n5204 = ~n5039 & ~n5203;
  assign n5205 = ~pi215 & ~n5204;
  assign n5206 = n5103 & ~n5205;
  assign n5207 = n5102 & ~n5206;
  assign n5208 = ~pi38 & ~n5192;
  assign n5209 = ~n5207 & n5208;
  assign n5210 = ~pi100 & ~n5191;
  assign n5211 = ~n5209 & n5210;
  assign n5212 = ~n2531 & n5178;
  assign n5213 = ~n5128 & n5156;
  assign n5214 = n5026 & ~n5213;
  assign n5215 = ~n5039 & ~n5214;
  assign n5216 = ~pi215 & ~n5215;
  assign n5217 = ~n5024 & ~n5216;
  assign n5218 = pi299 & ~n5217;
  assign n5219 = n2531 & n5176;
  assign n5220 = ~n5218 & n5219;
  assign n5221 = pi100 & ~n5212;
  assign n5222 = ~n5220 & n5221;
  assign n5223 = ~n5211 & ~n5222;
  assign n5224 = ~pi87 & ~n5223;
  assign n5225 = ~pi75 & ~n5190;
  assign n5226 = ~n5224 & n5225;
  assign n5227 = ~pi92 & ~n5189;
  assign n5228 = ~n5226 & n5227;
  assign n5229 = n2533 & ~n5188;
  assign n5230 = ~n5228 & n5229;
  assign n5231 = ~pi55 & ~n5179;
  assign n5232 = ~n5230 & n5231;
  assign n5233 = ~pi56 & ~n5175;
  assign n5234 = ~n5232 & n5233;
  assign n5235 = ~pi62 & ~n5171;
  assign n5236 = ~n5234 & n5235;
  assign n5237 = pi240 & n3291;
  assign n5238 = ~n5167 & n5237;
  assign n5239 = ~n5236 & n5238;
  assign n5240 = pi240 & n5163;
  assign n5241 = ~n3291 & ~n5240;
  assign n5242 = n5042 & n5241;
  assign n5243 = ~n5155 & ~n5242;
  assign po162 = ~n5239 & n5243;
  assign n5245 = pi215 & pi1136;
  assign n5246 = pi216 & pi266;
  assign n5247 = ~pi105 & pi166;
  assign n5248 = pi105 & ~n2442;
  assign n5249 = pi875 & n5248;
  assign n5250 = ~n5247 & ~n5249;
  assign n5251 = pi228 & ~n5250;
  assign n5252 = pi166 & ~pi228;
  assign n5253 = ~n5251 & ~n5252;
  assign n5254 = ~pi216 & ~n5253;
  assign n5255 = ~n5246 & ~n5254;
  assign n5256 = ~pi221 & ~n5255;
  assign n5257 = ~pi1136 & ~n2452;
  assign n5258 = ~pi928 & n2452;
  assign n5259 = pi221 & ~n5257;
  assign n5260 = ~n5258 & n5259;
  assign n5261 = ~n5256 & ~n5260;
  assign n5262 = ~pi215 & ~n5261;
  assign n5263 = ~n5245 & ~n5262;
  assign n5264 = ~n3291 & n5263;
  assign n5265 = ~n3317 & ~n5263;
  assign n5266 = ~pi875 & n2523;
  assign n5267 = ~n3524 & ~n5252;
  assign n5268 = ~n5266 & ~n5267;
  assign n5269 = ~n5251 & ~n5268;
  assign n5270 = ~pi216 & ~n5269;
  assign n5271 = ~n5246 & ~n5270;
  assign n5272 = ~pi221 & ~n5271;
  assign n5273 = ~n5260 & ~n5272;
  assign n5274 = ~pi215 & ~n5273;
  assign n5275 = ~n5245 & ~n5274;
  assign n5276 = n2538 & ~n5275;
  assign n5277 = ~pi56 & n5276;
  assign n5278 = ~n5265 & ~n5277;
  assign n5279 = pi62 & ~n5278;
  assign n5280 = ~n2538 & ~n5263;
  assign n5281 = pi56 & ~n5280;
  assign n5282 = ~n5276 & n5281;
  assign n5283 = ~n2577 & n5263;
  assign n5284 = n2577 & n5275;
  assign n5285 = pi55 & ~n5283;
  assign n5286 = ~n5284 & n5285;
  assign n5287 = pi223 & pi1136;
  assign n5288 = ~pi224 & ~pi875;
  assign n5289 = ~n2442 & n5288;
  assign n5290 = pi224 & ~pi266;
  assign n5291 = ~pi222 & ~n5290;
  assign n5292 = ~n5289 & n5291;
  assign n5293 = ~pi1136 & ~n2596;
  assign n5294 = ~pi928 & n2596;
  assign n5295 = pi222 & ~n5293;
  assign n5296 = ~n5294 & n5295;
  assign n5297 = ~n5292 & ~n5296;
  assign n5298 = ~pi223 & ~n5297;
  assign n5299 = ~n5287 & ~n5298;
  assign n5300 = ~pi299 & ~n5299;
  assign n5301 = ~n3440 & n5300;
  assign n5302 = pi299 & ~n5263;
  assign n5303 = ~n5301 & ~n5302;
  assign n5304 = ~n2533 & n5303;
  assign n5305 = ~n2628 & n5303;
  assign n5306 = pi299 & ~n5275;
  assign n5307 = ~n5301 & ~n5306;
  assign n5308 = n2628 & n5307;
  assign n5309 = ~n5305 & ~n5308;
  assign n5310 = n2534 & ~n5309;
  assign n5311 = ~n2534 & n5303;
  assign n5312 = pi92 & ~n5311;
  assign n5313 = ~n5310 & n5312;
  assign n5314 = pi75 & n5303;
  assign n5315 = pi87 & n5309;
  assign n5316 = pi38 & n5303;
  assign n5317 = pi39 & ~n5307;
  assign n5318 = n2608 & ~n3176;
  assign n5319 = n5292 & ~n5318;
  assign n5320 = ~pi299 & ~n5287;
  assign n5321 = ~n5296 & n5320;
  assign n5322 = ~n5319 & n5321;
  assign n5323 = n3472 & n5250;
  assign n5324 = ~pi216 & ~n5323;
  assign n5325 = pi166 & n3177;
  assign n5326 = ~pi166 & ~n3466;
  assign n5327 = pi875 & ~n5325;
  assign n5328 = ~n5326 & n5327;
  assign n5329 = pi166 & ~pi875;
  assign n5330 = ~n3392 & n5329;
  assign n5331 = ~n5328 & ~n5330;
  assign n5332 = ~pi228 & ~n5331;
  assign n5333 = ~n3472 & ~n5332;
  assign n5334 = n5324 & ~n5333;
  assign n5335 = ~n5246 & ~n5334;
  assign n5336 = ~pi221 & ~n5335;
  assign n5337 = ~n5260 & ~n5336;
  assign n5338 = ~pi215 & ~n5337;
  assign n5339 = pi299 & ~n5245;
  assign n5340 = ~n5338 & n5339;
  assign n5341 = n5297 & ~n5318;
  assign n5342 = ~pi223 & ~n5341;
  assign n5343 = n5320 & ~n5342;
  assign n5344 = ~pi39 & ~n5343;
  assign n5345 = ~n5322 & n5344;
  assign n5346 = ~n5340 & n5345;
  assign n5347 = ~pi38 & ~n5317;
  assign n5348 = ~n5346 & n5347;
  assign n5349 = ~pi100 & ~n5316;
  assign n5350 = ~n5348 & n5349;
  assign n5351 = ~n2531 & n5303;
  assign n5352 = ~pi875 & n3363;
  assign n5353 = pi166 & ~n5352;
  assign n5354 = n2664 & ~n3365;
  assign n5355 = ~n2664 & ~n3363;
  assign n5356 = pi875 & ~n5354;
  assign n5357 = ~n5355 & n5356;
  assign n5358 = ~n5353 & ~n5357;
  assign n5359 = ~pi228 & ~n5358;
  assign n5360 = ~n5251 & ~n5359;
  assign n5361 = ~pi216 & ~n5360;
  assign n5362 = ~n5246 & ~n5361;
  assign n5363 = ~pi221 & ~n5362;
  assign n5364 = ~n5260 & ~n5363;
  assign n5365 = ~pi215 & ~n5364;
  assign n5366 = ~n5245 & ~n5365;
  assign n5367 = pi299 & ~n5366;
  assign n5368 = n2531 & ~n5301;
  assign n5369 = ~n5367 & n5368;
  assign n5370 = pi100 & ~n5351;
  assign n5371 = ~n5369 & n5370;
  assign n5372 = ~n5350 & ~n5371;
  assign n5373 = ~pi87 & ~n5372;
  assign n5374 = ~pi75 & ~n5315;
  assign n5375 = ~n5373 & n5374;
  assign n5376 = ~pi92 & ~n5314;
  assign n5377 = ~n5375 & n5376;
  assign n5378 = n2533 & ~n5313;
  assign n5379 = ~n5377 & n5378;
  assign n5380 = ~pi55 & ~n5304;
  assign n5381 = ~n5379 & n5380;
  assign n5382 = ~pi56 & ~n5286;
  assign n5383 = ~n5381 & n5382;
  assign n5384 = ~pi62 & ~n5282;
  assign n5385 = ~n5383 & n5384;
  assign n5386 = n3291 & ~n5279;
  assign n5387 = ~n5385 & n5386;
  assign n5388 = ~pi245 & ~n5264;
  assign n5389 = ~n5387 & n5388;
  assign n5390 = ~n3422 & n5263;
  assign n5391 = ~n3291 & n5390;
  assign n5392 = ~n3317 & ~n5390;
  assign n5393 = ~n3421 & ~n5251;
  assign n5394 = ~n5268 & n5393;
  assign n5395 = ~pi216 & ~n5394;
  assign n5396 = ~n5246 & ~n5395;
  assign n5397 = ~pi221 & ~n5396;
  assign n5398 = ~n5260 & ~n5397;
  assign n5399 = ~pi215 & ~n5398;
  assign n5400 = ~n5245 & ~n5399;
  assign n5401 = n2538 & ~n5400;
  assign n5402 = ~pi56 & n5401;
  assign n5403 = ~n5392 & ~n5402;
  assign n5404 = pi62 & ~n5403;
  assign n5405 = ~n2538 & ~n5390;
  assign n5406 = pi56 & ~n5405;
  assign n5407 = ~n5401 & n5406;
  assign n5408 = ~n2577 & n5390;
  assign n5409 = n2577 & n5400;
  assign n5410 = pi55 & ~n5408;
  assign n5411 = ~n5409 & n5410;
  assign n5412 = pi299 & ~n5390;
  assign n5413 = ~n5300 & ~n5412;
  assign n5414 = ~n2533 & n5413;
  assign n5415 = ~n2628 & n5413;
  assign n5416 = pi299 & ~n5400;
  assign n5417 = ~n5300 & ~n5416;
  assign n5418 = n2628 & n5417;
  assign n5419 = ~n5415 & ~n5418;
  assign n5420 = n2534 & ~n5419;
  assign n5421 = ~n2534 & n5413;
  assign n5422 = pi92 & ~n5421;
  assign n5423 = ~n5420 & n5422;
  assign n5424 = pi75 & n5413;
  assign n5425 = pi87 & n5419;
  assign n5426 = pi38 & n5413;
  assign n5427 = pi39 & ~n5417;
  assign n5428 = ~pi166 & ~n3177;
  assign n5429 = pi166 & n3466;
  assign n5430 = ~pi875 & ~n5428;
  assign n5431 = ~n5429 & n5430;
  assign n5432 = ~pi166 & ~n3392;
  assign n5433 = pi875 & ~n5432;
  assign n5434 = ~pi228 & ~n5431;
  assign n5435 = ~n5433 & n5434;
  assign n5436 = n5324 & ~n5435;
  assign n5437 = ~n5246 & ~n5436;
  assign n5438 = ~pi221 & ~n5437;
  assign n5439 = ~n5260 & ~n5438;
  assign n5440 = ~pi215 & ~n5439;
  assign n5441 = n5339 & ~n5440;
  assign n5442 = n5344 & ~n5441;
  assign n5443 = ~pi38 & ~n5427;
  assign n5444 = ~n5442 & n5443;
  assign n5445 = ~pi100 & ~n5426;
  assign n5446 = ~n5444 & n5445;
  assign n5447 = ~n2531 & n5413;
  assign n5448 = ~n5359 & n5393;
  assign n5449 = ~pi216 & ~n5448;
  assign n5450 = ~n5246 & ~n5449;
  assign n5451 = ~pi221 & ~n5450;
  assign n5452 = ~n5260 & ~n5451;
  assign n5453 = ~pi215 & ~n5452;
  assign n5454 = ~n5245 & ~n5453;
  assign n5455 = pi299 & ~n5454;
  assign n5456 = n2531 & ~n5300;
  assign n5457 = ~n5455 & n5456;
  assign n5458 = pi100 & ~n5447;
  assign n5459 = ~n5457 & n5458;
  assign n5460 = ~n5446 & ~n5459;
  assign n5461 = ~pi87 & ~n5460;
  assign n5462 = ~pi75 & ~n5425;
  assign n5463 = ~n5461 & n5462;
  assign n5464 = ~pi92 & ~n5424;
  assign n5465 = ~n5463 & n5464;
  assign n5466 = n2533 & ~n5423;
  assign n5467 = ~n5465 & n5466;
  assign n5468 = ~pi55 & ~n5414;
  assign n5469 = ~n5467 & n5468;
  assign n5470 = ~pi56 & ~n5411;
  assign n5471 = ~n5469 & n5470;
  assign n5472 = ~pi62 & ~n5407;
  assign n5473 = ~n5471 & n5472;
  assign n5474 = n3291 & ~n5404;
  assign n5475 = ~n5473 & n5474;
  assign n5476 = pi245 & ~n5391;
  assign n5477 = ~n5475 & n5476;
  assign po163 = n5389 | n5477;
  assign n5479 = pi215 & pi1135;
  assign n5480 = pi216 & pi279;
  assign n5481 = ~pi105 & pi161;
  assign n5482 = pi879 & n5248;
  assign n5483 = ~n5481 & ~n5482;
  assign n5484 = pi228 & ~n5483;
  assign n5485 = pi161 & ~pi228;
  assign n5486 = ~n5484 & ~n5485;
  assign n5487 = ~pi216 & ~n5486;
  assign n5488 = ~n5480 & ~n5487;
  assign n5489 = ~pi221 & ~n5488;
  assign n5490 = ~pi1135 & ~n2452;
  assign n5491 = ~pi938 & n2452;
  assign n5492 = pi221 & ~n5490;
  assign n5493 = ~n5491 & n5492;
  assign n5494 = ~n5489 & ~n5493;
  assign n5495 = ~pi215 & ~n5494;
  assign n5496 = ~n5479 & ~n5495;
  assign n5497 = ~n3291 & n5496;
  assign n5498 = ~n3317 & ~n5496;
  assign n5499 = ~pi879 & n2523;
  assign n5500 = ~n3524 & ~n5485;
  assign n5501 = ~n5499 & ~n5500;
  assign n5502 = ~n5484 & ~n5501;
  assign n5503 = ~pi216 & ~n5502;
  assign n5504 = ~n5480 & ~n5503;
  assign n5505 = ~pi221 & ~n5504;
  assign n5506 = ~n5493 & ~n5505;
  assign n5507 = ~pi215 & ~n5506;
  assign n5508 = ~n5479 & ~n5507;
  assign n5509 = n2538 & ~n5508;
  assign n5510 = ~pi56 & n5509;
  assign n5511 = ~n5498 & ~n5510;
  assign n5512 = pi62 & ~n5511;
  assign n5513 = ~n2538 & ~n5496;
  assign n5514 = pi56 & ~n5513;
  assign n5515 = ~n5509 & n5514;
  assign n5516 = ~n2577 & n5496;
  assign n5517 = n2577 & n5508;
  assign n5518 = pi55 & ~n5516;
  assign n5519 = ~n5517 & n5518;
  assign n5520 = pi223 & pi1135;
  assign n5521 = ~pi1135 & ~n2596;
  assign n5522 = ~pi938 & n2596;
  assign n5523 = pi222 & ~n5521;
  assign n5524 = ~n5522 & n5523;
  assign n5525 = pi224 & ~pi279;
  assign n5526 = ~pi224 & ~pi879;
  assign n5527 = ~n2442 & n5526;
  assign n5528 = ~pi222 & ~n5525;
  assign n5529 = ~n5527 & n5528;
  assign n5530 = ~n5524 & ~n5529;
  assign n5531 = ~pi223 & ~n5530;
  assign n5532 = ~n5520 & ~n5531;
  assign n5533 = ~pi299 & ~n5532;
  assign n5534 = ~n3440 & n5533;
  assign n5535 = pi299 & ~n5496;
  assign n5536 = ~n5534 & ~n5535;
  assign n5537 = ~n2533 & n5536;
  assign n5538 = ~n2628 & n5536;
  assign n5539 = pi299 & ~n5508;
  assign n5540 = ~n5534 & ~n5539;
  assign n5541 = n2628 & n5540;
  assign n5542 = ~n5538 & ~n5541;
  assign n5543 = n2534 & ~n5542;
  assign n5544 = ~n2534 & n5536;
  assign n5545 = pi92 & ~n5544;
  assign n5546 = ~n5543 & n5545;
  assign n5547 = pi75 & n5536;
  assign n5548 = pi87 & n5542;
  assign n5549 = pi38 & n5536;
  assign n5550 = pi39 & ~n5540;
  assign n5551 = ~pi299 & ~n5520;
  assign n5552 = n5318 & ~n5524;
  assign n5553 = n5531 & ~n5552;
  assign n5554 = n5551 & ~n5553;
  assign n5555 = n3472 & n5483;
  assign n5556 = ~pi216 & ~n5555;
  assign n5557 = pi161 & n3177;
  assign n5558 = ~pi161 & ~n3466;
  assign n5559 = pi879 & ~n5557;
  assign n5560 = ~n5558 & n5559;
  assign n5561 = pi161 & ~pi879;
  assign n5562 = ~n3392 & n5561;
  assign n5563 = ~n5560 & ~n5562;
  assign n5564 = ~pi228 & ~n5563;
  assign n5565 = ~n3472 & ~n5564;
  assign n5566 = n5556 & ~n5565;
  assign n5567 = ~n5480 & ~n5566;
  assign n5568 = ~pi221 & ~n5567;
  assign n5569 = ~n5493 & ~n5568;
  assign n5570 = ~pi215 & ~n5569;
  assign n5571 = pi299 & ~n5479;
  assign n5572 = ~n5570 & n5571;
  assign n5573 = ~pi39 & ~n5554;
  assign n5574 = ~n5572 & n5573;
  assign n5575 = ~pi38 & ~n5550;
  assign n5576 = ~n5574 & n5575;
  assign n5577 = ~pi100 & ~n5549;
  assign n5578 = ~n5576 & n5577;
  assign n5579 = ~n2531 & n5536;
  assign n5580 = ~pi879 & n3363;
  assign n5581 = pi161 & ~n5580;
  assign n5582 = ~pi152 & ~pi166;
  assign n5583 = ~n3365 & n5582;
  assign n5584 = ~n3363 & ~n5582;
  assign n5585 = pi879 & ~n5583;
  assign n5586 = ~n5584 & n5585;
  assign n5587 = ~n5581 & ~n5586;
  assign n5588 = ~pi228 & ~n5587;
  assign n5589 = ~n5484 & ~n5588;
  assign n5590 = ~pi216 & ~n5589;
  assign n5591 = ~n5480 & ~n5590;
  assign n5592 = ~pi221 & ~n5591;
  assign n5593 = ~n5493 & ~n5592;
  assign n5594 = ~pi215 & ~n5593;
  assign n5595 = ~n5479 & ~n5594;
  assign n5596 = pi299 & ~n5595;
  assign n5597 = n2531 & ~n5534;
  assign n5598 = ~n5596 & n5597;
  assign n5599 = pi100 & ~n5579;
  assign n5600 = ~n5598 & n5599;
  assign n5601 = ~n5578 & ~n5600;
  assign n5602 = ~pi87 & ~n5601;
  assign n5603 = ~pi75 & ~n5548;
  assign n5604 = ~n5602 & n5603;
  assign n5605 = ~pi92 & ~n5547;
  assign n5606 = ~n5604 & n5605;
  assign n5607 = n2533 & ~n5546;
  assign n5608 = ~n5606 & n5607;
  assign n5609 = ~pi55 & ~n5537;
  assign n5610 = ~n5608 & n5609;
  assign n5611 = ~pi56 & ~n5519;
  assign n5612 = ~n5610 & n5611;
  assign n5613 = ~pi62 & ~n5515;
  assign n5614 = ~n5612 & n5613;
  assign n5615 = n3291 & ~n5512;
  assign n5616 = ~n5614 & n5615;
  assign n5617 = ~pi244 & ~n5497;
  assign n5618 = ~n5616 & n5617;
  assign n5619 = ~n3422 & n5496;
  assign n5620 = ~n3291 & n5619;
  assign n5621 = ~n3317 & ~n5619;
  assign n5622 = ~n3421 & ~n5484;
  assign n5623 = ~n5501 & n5622;
  assign n5624 = ~pi216 & ~n5623;
  assign n5625 = ~n5480 & ~n5624;
  assign n5626 = ~pi221 & ~n5625;
  assign n5627 = ~n5493 & ~n5626;
  assign n5628 = ~pi215 & ~n5627;
  assign n5629 = ~n5479 & ~n5628;
  assign n5630 = n2538 & ~n5629;
  assign n5631 = ~pi56 & n5630;
  assign n5632 = ~n5621 & ~n5631;
  assign n5633 = pi62 & ~n5632;
  assign n5634 = ~n2538 & ~n5619;
  assign n5635 = pi56 & ~n5634;
  assign n5636 = ~n5630 & n5635;
  assign n5637 = ~n2577 & n5619;
  assign n5638 = n2577 & n5629;
  assign n5639 = pi55 & ~n5637;
  assign n5640 = ~n5638 & n5639;
  assign n5641 = pi299 & ~n5619;
  assign n5642 = ~n5533 & ~n5641;
  assign n5643 = ~n2533 & n5642;
  assign n5644 = ~n2628 & n5642;
  assign n5645 = pi299 & ~n5629;
  assign n5646 = ~n5533 & ~n5645;
  assign n5647 = n2628 & n5646;
  assign n5648 = ~n5644 & ~n5647;
  assign n5649 = n2534 & ~n5648;
  assign n5650 = ~n2534 & n5642;
  assign n5651 = pi92 & ~n5650;
  assign n5652 = ~n5649 & n5651;
  assign n5653 = pi75 & n5642;
  assign n5654 = pi87 & n5648;
  assign n5655 = pi38 & n5642;
  assign n5656 = pi39 & ~n5646;
  assign n5657 = ~n5318 & n5530;
  assign n5658 = ~pi223 & ~n5657;
  assign n5659 = n5551 & ~n5658;
  assign n5660 = ~pi161 & ~n3177;
  assign n5661 = pi161 & n3466;
  assign n5662 = ~pi879 & ~n5660;
  assign n5663 = ~n5661 & n5662;
  assign n5664 = ~pi161 & ~n3392;
  assign n5665 = pi879 & ~n5664;
  assign n5666 = ~pi228 & ~n5663;
  assign n5667 = ~n5665 & n5666;
  assign n5668 = n5556 & ~n5667;
  assign n5669 = ~n5480 & ~n5668;
  assign n5670 = ~pi221 & ~n5669;
  assign n5671 = ~n5493 & ~n5670;
  assign n5672 = ~pi215 & ~n5671;
  assign n5673 = n5571 & ~n5672;
  assign n5674 = ~pi39 & ~n5659;
  assign n5675 = ~n5673 & n5674;
  assign n5676 = ~pi38 & ~n5656;
  assign n5677 = ~n5675 & n5676;
  assign n5678 = ~pi100 & ~n5655;
  assign n5679 = ~n5677 & n5678;
  assign n5680 = ~n2531 & n5642;
  assign n5681 = ~n5588 & n5622;
  assign n5682 = ~pi216 & ~n5681;
  assign n5683 = ~n5480 & ~n5682;
  assign n5684 = ~pi221 & ~n5683;
  assign n5685 = ~n5493 & ~n5684;
  assign n5686 = ~pi215 & ~n5685;
  assign n5687 = ~n5479 & ~n5686;
  assign n5688 = pi299 & ~n5687;
  assign n5689 = n2531 & ~n5533;
  assign n5690 = ~n5688 & n5689;
  assign n5691 = pi100 & ~n5680;
  assign n5692 = ~n5690 & n5691;
  assign n5693 = ~n5679 & ~n5692;
  assign n5694 = ~pi87 & ~n5693;
  assign n5695 = ~pi75 & ~n5654;
  assign n5696 = ~n5694 & n5695;
  assign n5697 = ~pi92 & ~n5653;
  assign n5698 = ~n5696 & n5697;
  assign n5699 = n2533 & ~n5652;
  assign n5700 = ~n5698 & n5699;
  assign n5701 = ~pi55 & ~n5643;
  assign n5702 = ~n5700 & n5701;
  assign n5703 = ~pi56 & ~n5640;
  assign n5704 = ~n5702 & n5703;
  assign n5705 = ~pi62 & ~n5636;
  assign n5706 = ~n5704 & n5705;
  assign n5707 = n3291 & ~n5633;
  assign n5708 = ~n5706 & n5707;
  assign n5709 = pi244 & ~n5620;
  assign n5710 = ~n5708 & n5709;
  assign po164 = n5618 | n5710;
  assign n5712 = pi216 & pi278;
  assign n5713 = ~pi221 & ~n5712;
  assign n5714 = ~pi105 & pi152;
  assign n5715 = pi846 & ~n2442;
  assign n5716 = pi105 & n5715;
  assign n5717 = ~n5714 & ~n5716;
  assign n5718 = pi228 & ~n5717;
  assign n5719 = pi152 & ~pi228;
  assign n5720 = ~n5718 & ~n5719;
  assign n5721 = ~pi216 & ~n5720;
  assign n5722 = n5713 & ~n5721;
  assign n5723 = pi833 & ~pi930;
  assign n5724 = ~pi216 & pi221;
  assign n5725 = n5723 & n5724;
  assign n5726 = ~pi215 & pi221;
  assign n5727 = ~pi216 & n5726;
  assign n5728 = pi833 & n5727;
  assign n5729 = ~n2461 & ~n5728;
  assign n5730 = ~n5725 & ~n5729;
  assign n5731 = ~n5722 & n5730;
  assign n5732 = ~n3422 & ~n5731;
  assign n5733 = ~n3291 & ~n5732;
  assign n5734 = ~n3421 & ~n5718;
  assign n5735 = ~pi846 & n2523;
  assign n5736 = ~n3524 & ~n5719;
  assign n5737 = ~n5735 & ~n5736;
  assign n5738 = n5734 & ~n5737;
  assign n5739 = ~pi216 & ~n5738;
  assign n5740 = n5713 & ~n5739;
  assign n5741 = n5730 & ~n5740;
  assign n5742 = n2538 & ~n5741;
  assign n5743 = ~pi56 & n5742;
  assign n5744 = ~n3317 & n5732;
  assign n5745 = ~n5743 & ~n5744;
  assign n5746 = pi62 & ~n5745;
  assign n5747 = ~n2538 & n5732;
  assign n5748 = pi56 & ~n5747;
  assign n5749 = ~n5742 & n5748;
  assign n5750 = ~n2577 & ~n5732;
  assign n5751 = n2577 & n5741;
  assign n5752 = pi55 & ~n5750;
  assign n5753 = ~n5751 & n5752;
  assign n5754 = pi222 & ~pi224;
  assign n5755 = n5723 & n5754;
  assign n5756 = pi224 & pi278;
  assign n5757 = ~pi222 & ~n5756;
  assign n5758 = ~pi224 & n5715;
  assign n5759 = n5757 & ~n5758;
  assign n5760 = n2598 & ~n5755;
  assign n5761 = ~n5759 & n5760;
  assign n5762 = ~pi299 & ~n5761;
  assign n5763 = ~n3440 & n5762;
  assign n5764 = pi299 & n5732;
  assign n5765 = ~n5763 & ~n5764;
  assign n5766 = ~n2533 & n5765;
  assign n5767 = ~n2628 & n5765;
  assign n5768 = pi299 & ~n5741;
  assign n5769 = ~n5763 & ~n5768;
  assign n5770 = n2628 & n5769;
  assign n5771 = ~n5767 & ~n5770;
  assign n5772 = n2534 & ~n5771;
  assign n5773 = ~n2534 & n5765;
  assign n5774 = pi92 & ~n5773;
  assign n5775 = ~n5772 & n5774;
  assign n5776 = pi75 & n5765;
  assign n5777 = pi87 & n5771;
  assign n5778 = pi38 & n5765;
  assign n5779 = pi39 & ~n5769;
  assign n5780 = ~pi846 & n3176;
  assign n5781 = ~pi224 & ~n5780;
  assign n5782 = n5757 & ~n5781;
  assign n5783 = ~pi223 & ~pi299;
  assign n5784 = ~n2597 & n5783;
  assign n5785 = ~n5755 & n5784;
  assign n5786 = ~n5782 & n5785;
  assign n5787 = pi228 & ~n5714;
  assign n5788 = pi105 & ~n5780;
  assign n5789 = n5787 & ~n5788;
  assign n5790 = ~pi216 & ~n5789;
  assign n5791 = ~pi152 & n3177;
  assign n5792 = pi152 & ~n3466;
  assign n5793 = ~pi846 & ~n5791;
  assign n5794 = ~n5792 & n5793;
  assign n5795 = ~pi152 & pi846;
  assign n5796 = ~n3392 & n5795;
  assign n5797 = ~n5794 & ~n5796;
  assign n5798 = ~pi228 & ~n5797;
  assign n5799 = n5790 & ~n5798;
  assign n5800 = n5713 & ~n5799;
  assign n5801 = ~n5725 & ~n5800;
  assign n5802 = pi299 & ~n5729;
  assign n5803 = n5801 & n5802;
  assign n5804 = ~pi39 & ~n5786;
  assign n5805 = ~n5803 & n5804;
  assign n5806 = ~pi38 & ~n5779;
  assign n5807 = ~n5805 & n5806;
  assign n5808 = ~pi100 & ~n5778;
  assign n5809 = ~n5807 & n5808;
  assign n5810 = ~n2531 & n5765;
  assign n5811 = pi846 & ~n3370;
  assign n5812 = ~n3364 & ~n5811;
  assign n5813 = ~pi228 & ~n5812;
  assign n5814 = n5734 & ~n5813;
  assign n5815 = ~pi216 & ~n5814;
  assign n5816 = n5713 & ~n5815;
  assign n5817 = n5730 & ~n5816;
  assign n5818 = pi299 & ~n5817;
  assign n5819 = n2531 & ~n5763;
  assign n5820 = ~n5818 & n5819;
  assign n5821 = pi100 & ~n5810;
  assign n5822 = ~n5820 & n5821;
  assign n5823 = ~n5809 & ~n5822;
  assign n5824 = ~pi87 & ~n5823;
  assign n5825 = ~pi75 & ~n5777;
  assign n5826 = ~n5824 & n5825;
  assign n5827 = ~pi92 & ~n5776;
  assign n5828 = ~n5826 & n5827;
  assign n5829 = n2533 & ~n5775;
  assign n5830 = ~n5828 & n5829;
  assign n5831 = ~pi55 & ~n5766;
  assign n5832 = ~n5830 & n5831;
  assign n5833 = ~pi56 & ~n5753;
  assign n5834 = ~n5832 & n5833;
  assign n5835 = ~pi62 & ~n5749;
  assign n5836 = ~n5834 & n5835;
  assign n5837 = n3291 & ~n5746;
  assign n5838 = ~n5836 & n5837;
  assign n5839 = pi242 & ~n5733;
  assign n5840 = ~n5838 & n5839;
  assign n5841 = ~n3291 & n5731;
  assign n5842 = ~n3317 & ~n5731;
  assign n5843 = ~n5718 & ~n5737;
  assign n5844 = ~pi216 & ~n5843;
  assign n5845 = n5713 & ~n5844;
  assign n5846 = n5730 & ~n5845;
  assign n5847 = n2538 & ~n5846;
  assign n5848 = ~pi56 & n5847;
  assign n5849 = ~n5842 & ~n5848;
  assign n5850 = pi62 & ~n5849;
  assign n5851 = ~n2538 & ~n5731;
  assign n5852 = pi56 & ~n5851;
  assign n5853 = ~n5847 & n5852;
  assign n5854 = ~n2577 & n5731;
  assign n5855 = n2577 & n5846;
  assign n5856 = pi55 & ~n5854;
  assign n5857 = ~n5855 & n5856;
  assign n5858 = pi299 & ~n5731;
  assign n5859 = ~n5762 & ~n5858;
  assign n5860 = ~n2533 & n5859;
  assign n5861 = ~n2628 & n5859;
  assign n5862 = pi299 & ~n5846;
  assign n5863 = ~n5762 & ~n5862;
  assign n5864 = n2628 & n5863;
  assign n5865 = ~n5861 & ~n5864;
  assign n5866 = n2534 & ~n5865;
  assign n5867 = ~n2534 & n5859;
  assign n5868 = pi92 & ~n5867;
  assign n5869 = ~n5866 & n5868;
  assign n5870 = pi75 & n5859;
  assign n5871 = pi87 & n5865;
  assign n5872 = pi38 & n5859;
  assign n5873 = pi39 & ~n5863;
  assign n5874 = ~n3175 & n5758;
  assign n5875 = n5757 & ~n5874;
  assign n5876 = n5785 & ~n5875;
  assign n5877 = ~n3176 & n5787;
  assign n5878 = pi152 & ~pi846;
  assign n5879 = ~n3392 & n5878;
  assign n5880 = pi152 & n3177;
  assign n5881 = ~pi152 & ~n3466;
  assign n5882 = pi846 & ~n5880;
  assign n5883 = ~n5881 & n5882;
  assign n5884 = ~pi228 & ~n5879;
  assign n5885 = ~n5883 & n5884;
  assign n5886 = n5790 & ~n5877;
  assign n5887 = ~n5885 & n5886;
  assign n5888 = n5713 & ~n5887;
  assign n5889 = ~n5725 & ~n5888;
  assign n5890 = n5802 & n5889;
  assign n5891 = ~pi39 & ~n5876;
  assign n5892 = ~n5890 & n5891;
  assign n5893 = ~pi38 & ~n5873;
  assign n5894 = ~n5892 & n5893;
  assign n5895 = ~pi100 & ~n5872;
  assign n5896 = ~n5894 & n5895;
  assign n5897 = ~n2531 & n5859;
  assign n5898 = ~n5718 & ~n5813;
  assign n5899 = ~pi216 & ~n5898;
  assign n5900 = n5713 & ~n5899;
  assign n5901 = n5730 & ~n5900;
  assign n5902 = pi299 & ~n5901;
  assign n5903 = n2531 & ~n5762;
  assign n5904 = ~n5902 & n5903;
  assign n5905 = pi100 & ~n5897;
  assign n5906 = ~n5904 & n5905;
  assign n5907 = ~n5896 & ~n5906;
  assign n5908 = ~pi87 & ~n5907;
  assign n5909 = ~pi75 & ~n5871;
  assign n5910 = ~n5908 & n5909;
  assign n5911 = ~pi92 & ~n5870;
  assign n5912 = ~n5910 & n5911;
  assign n5913 = n2533 & ~n5869;
  assign n5914 = ~n5912 & n5913;
  assign n5915 = ~pi55 & ~n5860;
  assign n5916 = ~n5914 & n5915;
  assign n5917 = ~pi56 & ~n5857;
  assign n5918 = ~n5916 & n5917;
  assign n5919 = ~pi62 & ~n5853;
  assign n5920 = ~n5918 & n5919;
  assign n5921 = n3291 & ~n5850;
  assign n5922 = ~n5920 & n5921;
  assign n5923 = ~pi242 & ~n5841;
  assign n5924 = ~n5922 & n5923;
  assign n5925 = ~n5840 & ~n5924;
  assign n5926 = ~pi1134 & ~n5925;
  assign n5927 = ~n5722 & ~n5725;
  assign n5928 = ~pi215 & ~n5927;
  assign n5929 = ~n3422 & n5928;
  assign n5930 = ~n3291 & n5929;
  assign n5931 = ~n3317 & ~n5929;
  assign n5932 = ~n5725 & ~n5740;
  assign n5933 = ~pi215 & ~n5932;
  assign n5934 = n2538 & ~n5933;
  assign n5935 = ~pi56 & n5934;
  assign n5936 = ~n5931 & ~n5935;
  assign n5937 = pi62 & ~n5936;
  assign n5938 = ~n2538 & ~n5929;
  assign n5939 = pi56 & ~n5938;
  assign n5940 = ~n5934 & n5939;
  assign n5941 = ~n2577 & n5929;
  assign n5942 = n2577 & n5933;
  assign n5943 = pi55 & ~n5941;
  assign n5944 = ~n5942 & n5943;
  assign n5945 = n2598 & n5763;
  assign n5946 = ~pi299 & ~n5945;
  assign n5947 = pi299 & ~n5929;
  assign n5948 = ~n5946 & ~n5947;
  assign n5949 = ~n2533 & n5948;
  assign n5950 = ~n2628 & n5948;
  assign n5951 = pi299 & ~n5933;
  assign n5952 = ~n5946 & ~n5951;
  assign n5953 = n2628 & n5952;
  assign n5954 = ~n5950 & ~n5953;
  assign n5955 = n2534 & ~n5954;
  assign n5956 = ~n2534 & n5948;
  assign n5957 = pi92 & ~n5956;
  assign n5958 = ~n5955 & n5957;
  assign n5959 = pi75 & n5948;
  assign n5960 = pi87 & n5954;
  assign n5961 = pi38 & n5948;
  assign n5962 = pi39 & ~n5952;
  assign n5963 = ~n5755 & ~n5782;
  assign n5964 = n5783 & ~n5963;
  assign n5965 = ~pi39 & ~n5964;
  assign n5966 = ~pi215 & pi299;
  assign n5967 = ~n5801 & n5966;
  assign n5968 = n5965 & ~n5967;
  assign n5969 = ~pi38 & ~n5962;
  assign n5970 = ~n5968 & n5969;
  assign n5971 = ~pi100 & ~n5961;
  assign n5972 = ~n5970 & n5971;
  assign n5973 = ~n2531 & n5948;
  assign n5974 = ~n5725 & ~n5816;
  assign n5975 = ~pi215 & ~n5974;
  assign n5976 = pi299 & ~n5975;
  assign n5977 = n2531 & ~n5946;
  assign n5978 = ~n5976 & n5977;
  assign n5979 = pi100 & ~n5973;
  assign n5980 = ~n5978 & n5979;
  assign n5981 = ~n5972 & ~n5980;
  assign n5982 = ~pi87 & ~n5981;
  assign n5983 = ~pi75 & ~n5960;
  assign n5984 = ~n5982 & n5983;
  assign n5985 = ~pi92 & ~n5959;
  assign n5986 = ~n5984 & n5985;
  assign n5987 = n2533 & ~n5958;
  assign n5988 = ~n5986 & n5987;
  assign n5989 = ~pi55 & ~n5949;
  assign n5990 = ~n5988 & n5989;
  assign n5991 = ~pi56 & ~n5944;
  assign n5992 = ~n5990 & n5991;
  assign n5993 = ~pi62 & ~n5940;
  assign n5994 = ~n5992 & n5993;
  assign n5995 = n3291 & ~n5937;
  assign n5996 = ~n5994 & n5995;
  assign n5997 = pi242 & ~n5930;
  assign n5998 = ~n5996 & n5997;
  assign n5999 = ~n3291 & n5928;
  assign n6000 = ~n3317 & ~n5928;
  assign n6001 = ~n5725 & ~n5845;
  assign n6002 = ~pi215 & ~n6001;
  assign n6003 = n2538 & ~n6002;
  assign n6004 = ~pi56 & n6003;
  assign n6005 = ~n6000 & ~n6004;
  assign n6006 = pi62 & ~n6005;
  assign n6007 = ~n2538 & ~n5928;
  assign n6008 = pi56 & ~n6007;
  assign n6009 = ~n6003 & n6008;
  assign n6010 = ~n2577 & n5928;
  assign n6011 = n2577 & n6002;
  assign n6012 = pi55 & ~n6010;
  assign n6013 = ~n6011 & n6012;
  assign n6014 = pi299 & ~n5928;
  assign n6015 = ~n3440 & n5946;
  assign n6016 = ~n6014 & ~n6015;
  assign n6017 = ~n2533 & n6016;
  assign n6018 = ~n2628 & n6016;
  assign n6019 = pi299 & ~n6002;
  assign n6020 = ~n6015 & ~n6019;
  assign n6021 = n2628 & n6020;
  assign n6022 = ~n6018 & ~n6021;
  assign n6023 = n2534 & ~n6022;
  assign n6024 = ~n2534 & n6016;
  assign n6025 = pi92 & ~n6024;
  assign n6026 = ~n6023 & n6025;
  assign n6027 = pi75 & n6016;
  assign n6028 = pi87 & n6022;
  assign n6029 = pi38 & n6016;
  assign n6030 = pi39 & ~n6020;
  assign n6031 = n5783 & n5875;
  assign n6032 = ~n5889 & n5966;
  assign n6033 = n5965 & ~n6031;
  assign n6034 = ~n6032 & n6033;
  assign n6035 = ~pi38 & ~n6030;
  assign n6036 = ~n6034 & n6035;
  assign n6037 = ~pi100 & ~n6029;
  assign n6038 = ~n6036 & n6037;
  assign n6039 = ~n2531 & n6016;
  assign n6040 = ~n5725 & ~n5900;
  assign n6041 = ~pi215 & ~n6040;
  assign n6042 = pi299 & ~n6041;
  assign n6043 = n2531 & ~n6015;
  assign n6044 = ~n6042 & n6043;
  assign n6045 = pi100 & ~n6039;
  assign n6046 = ~n6044 & n6045;
  assign n6047 = ~n6038 & ~n6046;
  assign n6048 = ~pi87 & ~n6047;
  assign n6049 = ~pi75 & ~n6028;
  assign n6050 = ~n6048 & n6049;
  assign n6051 = ~pi92 & ~n6027;
  assign n6052 = ~n6050 & n6051;
  assign n6053 = n2533 & ~n6026;
  assign n6054 = ~n6052 & n6053;
  assign n6055 = ~pi55 & ~n6017;
  assign n6056 = ~n6054 & n6055;
  assign n6057 = ~pi56 & ~n6013;
  assign n6058 = ~n6056 & n6057;
  assign n6059 = ~pi62 & ~n6009;
  assign n6060 = ~n6058 & n6059;
  assign n6061 = n3291 & ~n6006;
  assign n6062 = ~n6060 & n6061;
  assign n6063 = ~pi242 & ~n5999;
  assign n6064 = ~n6062 & n6063;
  assign n6065 = pi1134 & ~n6064;
  assign n6066 = ~n5998 & n6065;
  assign po165 = ~n5926 & ~n6066;
  assign n6068 = pi57 & pi59;
  assign n6069 = n2523 & n2539;
  assign n6070 = ~n3291 & ~n6069;
  assign n6071 = ~n6068 & ~n6070;
  assign n6072 = pi57 & ~n6071;
  assign n6073 = n2513 & n2628;
  assign n6074 = ~pi54 & n2535;
  assign n6075 = n6073 & n6074;
  assign n6076 = pi74 & ~n6075;
  assign n6077 = ~pi55 & ~n6076;
  assign n6078 = ~pi54 & ~pi92;
  assign n6079 = pi87 & ~n6073;
  assign n6080 = ~pi75 & ~n6079;
  assign n6081 = ~pi39 & n2523;
  assign n6082 = ~pi38 & pi100;
  assign n6083 = n6081 & n6082;
  assign n6084 = ~pi299 & ~n2641;
  assign n6085 = pi299 & ~n2665;
  assign n6086 = ~n6084 & ~n6085;
  assign n6087 = pi146 & n6085;
  assign n6088 = pi142 & n6084;
  assign n6089 = ~n6087 & ~n6088;
  assign n6090 = ~n6086 & n6089;
  assign n6091 = ~pi41 & ~pi99;
  assign n6092 = ~pi101 & n6091;
  assign n6093 = ~pi42 & ~pi43;
  assign n6094 = ~pi52 & n6093;
  assign n6095 = ~pi113 & ~pi116;
  assign n6096 = ~pi114 & ~pi115;
  assign n6097 = n6095 & n6096;
  assign n6098 = n6094 & n6097;
  assign n6099 = n6092 & n6098;
  assign po1057 = pi44 | ~n6099;
  assign n6101 = ~pi683 & po1057;
  assign n6102 = pi950 & pi1092;
  assign n6103 = ~pi824 & ~pi829;
  assign n6104 = n6102 & ~n6103;
  assign po740 = ~pi1093 & n6104;
  assign n6106 = ~pi250 & ~po740;
  assign n6107 = pi129 & pi250;
  assign n6108 = ~n6106 & ~n6107;
  assign n6109 = ~n6101 & ~n6108;
  assign n6110 = n6090 & ~n6109;
  assign n6111 = n3365 & ~n6090;
  assign n6112 = n6090 & ~po1057;
  assign n6113 = ~n6110 & ~n6112;
  assign n6114 = ~n6111 & n6113;
  assign n6115 = n6083 & ~n6114;
  assign n6116 = ~pi39 & n2513;
  assign n6117 = pi38 & ~n6116;
  assign n6118 = ~pi100 & ~n6117;
  assign n6119 = n2720 & n2767;
  assign n6120 = n2874 & n6119;
  assign n6121 = n2778 & ~n6120;
  assign n6122 = ~n2775 & ~n6121;
  assign n6123 = ~pi108 & ~n6122;
  assign n6124 = n2774 & ~n6123;
  assign n6125 = ~pi110 & n2890;
  assign n6126 = ~n6124 & n6125;
  assign n6127 = ~n2759 & ~n2766;
  assign n6128 = ~n6126 & n6127;
  assign n6129 = ~pi47 & ~n6128;
  assign n6130 = n2705 & ~n2762;
  assign n6131 = ~n6129 & n6130;
  assign n6132 = pi58 & n2504;
  assign n6133 = ~pi90 & ~n6132;
  assign n6134 = ~n6131 & n6133;
  assign n6135 = ~n2897 & ~n6134;
  assign n6136 = ~pi93 & ~n6135;
  assign n6137 = ~pi841 & n2505;
  assign n6138 = pi93 & ~n6137;
  assign n6139 = ~n6136 & ~n6138;
  assign n6140 = ~pi35 & ~n6139;
  assign n6141 = ~pi70 & ~n2728;
  assign n6142 = ~n6140 & n6141;
  assign n6143 = ~pi51 & ~n6142;
  assign n6144 = n2748 & ~n6143;
  assign n6145 = n3149 & ~n6144;
  assign n6146 = n2745 & ~n6145;
  assign n6147 = n2743 & ~n6146;
  assign n6148 = pi210 & pi299;
  assign n6149 = pi198 & ~pi299;
  assign n6150 = ~n6148 & ~n6149;
  assign n6151 = ~n3388 & ~n6150;
  assign n6152 = pi32 & ~n2917;
  assign n6153 = n6150 & ~n6152;
  assign n6154 = ~n6151 & ~n6153;
  assign n6155 = ~n6147 & ~n6154;
  assign n6156 = ~pi95 & ~n6155;
  assign n6157 = ~n2740 & ~n6156;
  assign n6158 = ~pi39 & ~n6157;
  assign n6159 = pi603 & ~pi642;
  assign n6160 = ~pi614 & ~pi616;
  assign n6161 = n6159 & n6160;
  assign n6162 = ~pi661 & ~pi681;
  assign n6163 = ~pi662 & pi680;
  assign n6164 = n6162 & n6163;
  assign po1101 = n6161 | n6164;
  assign n6166 = ~pi332 & ~pi468;
  assign n6167 = pi835 & pi984;
  assign n6168 = ~pi252 & ~pi1001;
  assign n6169 = ~pi979 & ~n6168;
  assign n6170 = ~n6167 & n6169;
  assign n6171 = ~pi287 & n6170;
  assign n6172 = pi835 & pi950;
  assign n6173 = n6171 & n6172;
  assign n6174 = pi1092 & n6173;
  assign n6175 = pi1093 & ~n2922;
  assign n6176 = pi829 & ~n6175;
  assign n6177 = ~pi824 & ~n6176;
  assign n6178 = pi1091 & pi1093;
  assign n6179 = n2921 & n6178;
  assign n6180 = ~n6177 & ~n6179;
  assign n6181 = n6174 & n6180;
  assign n6182 = ~n6166 & ~n6181;
  assign n6183 = po1101 & ~n6182;
  assign n6184 = n2523 & ~n6183;
  assign n6185 = n2513 & n6166;
  assign n6186 = po1101 & n6185;
  assign n6187 = ~n6184 & ~n6186;
  assign n6188 = ~pi587 & ~pi602;
  assign n6189 = ~pi961 & ~pi967;
  assign n6190 = ~pi969 & ~pi971;
  assign n6191 = ~pi974 & ~pi977;
  assign n6192 = n6190 & n6191;
  assign n6193 = n6188 & n6189;
  assign n6194 = n6192 & n6193;
  assign n6195 = n6187 & n6194;
  assign n6196 = ~n6161 & ~n6166;
  assign n6197 = ~n6164 & n6196;
  assign n6198 = n6181 & ~n6197;
  assign n6199 = n2523 & ~n6198;
  assign n6200 = ~n6194 & ~n6199;
  assign n6201 = pi223 & ~n6200;
  assign n6202 = ~n6195 & n6201;
  assign n6203 = n2926 & n6173;
  assign n6204 = pi222 & pi224;
  assign n6205 = po1101 & ~n6166;
  assign n6206 = n6166 & ~n6194;
  assign n6207 = ~n6205 & ~n6206;
  assign n6208 = n6204 & ~n6207;
  assign n6209 = n6203 & n6208;
  assign n6210 = ~pi223 & ~n6209;
  assign n6211 = n2523 & n6210;
  assign n6212 = ~n6202 & ~n6211;
  assign n6213 = ~pi299 & ~n6212;
  assign n6214 = pi216 & pi221;
  assign n6215 = ~pi960 & ~pi963;
  assign n6216 = ~pi970 & ~pi972;
  assign n6217 = ~pi975 & ~pi978;
  assign n6218 = n6216 & n6217;
  assign n6219 = n6215 & n6218;
  assign n6220 = ~pi907 & ~pi947;
  assign n6221 = n6219 & n6220;
  assign n6222 = n6166 & ~n6221;
  assign n6223 = ~n6205 & ~n6222;
  assign n6224 = n6203 & n6214;
  assign n6225 = ~n6223 & n6224;
  assign n6226 = n2523 & ~n6225;
  assign n6227 = ~pi215 & ~n6226;
  assign n6228 = n6199 & ~n6221;
  assign n6229 = ~n6187 & n6221;
  assign n6230 = pi215 & ~n6228;
  assign n6231 = ~n6229 & n6230;
  assign n6232 = pi299 & ~n6227;
  assign n6233 = ~n6231 & n6232;
  assign n6234 = pi39 & ~n6233;
  assign n6235 = ~n6213 & n6234;
  assign n6236 = ~n6158 & ~n6235;
  assign n6237 = ~pi38 & ~n6236;
  assign n6238 = n6118 & ~n6237;
  assign n6239 = ~pi87 & ~n6115;
  assign n6240 = ~n6238 & n6239;
  assign n6241 = n6078 & n6080;
  assign n6242 = ~n6240 & n6241;
  assign n6243 = ~pi74 & ~n6242;
  assign n6244 = n6077 & ~n6243;
  assign n6245 = ~pi56 & ~n6244;
  assign n6246 = ~pi55 & ~pi74;
  assign n6247 = n6075 & n6246;
  assign n6248 = pi56 & ~n6247;
  assign n6249 = ~n6245 & ~n6248;
  assign n6250 = ~pi62 & ~n6249;
  assign n6251 = n3316 & n6073;
  assign n6252 = pi62 & ~n6251;
  assign n6253 = ~pi59 & ~n6252;
  assign n6254 = ~n6250 & n6253;
  assign n6255 = ~pi57 & ~n6254;
  assign po167 = ~n6072 & ~n6255;
  assign n6257 = ~pi55 & n2530;
  assign n6258 = ~pi59 & n6257;
  assign n6259 = ~pi228 & ~n6258;
  assign n6260 = pi57 & ~n6259;
  assign n6261 = ~n6164 & ~n6166;
  assign n6262 = ~pi907 & n6166;
  assign n6263 = ~n6261 & ~n6262;
  assign n6264 = ~pi228 & ~n2577;
  assign n6265 = pi30 & pi228;
  assign n6266 = ~n3524 & ~n6265;
  assign n6267 = ~n6264 & ~n6266;
  assign n6268 = n6263 & n6267;
  assign n6269 = n6260 & n6268;
  assign n6270 = ~pi228 & ~n6257;
  assign n6271 = n6268 & ~n6270;
  assign n6272 = pi59 & ~n6271;
  assign n6273 = n6263 & n6265;
  assign n6274 = ~n2530 & n6273;
  assign n6275 = pi55 & ~n6268;
  assign n6276 = ~pi54 & n2572;
  assign n6277 = pi299 & n6263;
  assign n6278 = ~pi602 & n6166;
  assign n6279 = ~n6261 & ~n6278;
  assign n6280 = ~pi299 & n6279;
  assign n6281 = ~n6277 & ~n6280;
  assign n6282 = n6265 & ~n6281;
  assign n6283 = ~n6276 & ~n6282;
  assign n6284 = ~n2615 & n6282;
  assign n6285 = ~pi39 & ~n6266;
  assign n6286 = ~n6281 & n6285;
  assign n6287 = n2574 & n6286;
  assign n6288 = ~n6284 & ~n6287;
  assign n6289 = n2572 & n6288;
  assign n6290 = ~pi54 & n6289;
  assign n6291 = pi74 & ~n6283;
  assign n6292 = ~n6290 & n6291;
  assign n6293 = ~n2572 & ~n6282;
  assign n6294 = ~n6289 & ~n6293;
  assign n6295 = pi54 & ~n6294;
  assign n6296 = ~pi75 & n6288;
  assign n6297 = pi75 & ~n6282;
  assign n6298 = pi92 & ~n6297;
  assign n6299 = ~n6296 & n6298;
  assign n6300 = pi75 & n6288;
  assign n6301 = pi87 & n6282;
  assign n6302 = ~n2531 & n6282;
  assign n6303 = pi299 & ~n6273;
  assign n6304 = pi252 & n6185;
  assign n6305 = ~n6164 & ~n6304;
  assign n6306 = pi252 & n2523;
  assign n6307 = n6164 & ~n6306;
  assign n6308 = ~n6305 & ~n6307;
  assign n6309 = ~n2666 & ~n6308;
  assign n6310 = n2523 & ~n6108;
  assign n6311 = pi683 & n6310;
  assign n6312 = po1057 & n6311;
  assign n6313 = ~n6261 & n6312;
  assign n6314 = n2666 & ~n6313;
  assign n6315 = ~pi228 & ~n6262;
  assign n6316 = ~n6314 & n6315;
  assign n6317 = ~n6309 & n6316;
  assign n6318 = n6303 & ~n6317;
  assign n6319 = n6265 & n6279;
  assign n6320 = ~pi142 & ~n2641;
  assign n6321 = n6313 & n6320;
  assign n6322 = pi252 & ~n6320;
  assign n6323 = n6308 & n6322;
  assign n6324 = ~n6321 & ~n6323;
  assign n6325 = ~pi228 & ~n6278;
  assign n6326 = ~n6324 & n6325;
  assign n6327 = ~pi299 & ~n6319;
  assign n6328 = ~n6326 & n6327;
  assign n6329 = n2531 & ~n6318;
  assign n6330 = ~n6328 & n6329;
  assign n6331 = pi100 & ~n6302;
  assign n6332 = ~n6330 & n6331;
  assign n6333 = ~pi287 & n2523;
  assign n6334 = pi835 & n6170;
  assign n6335 = n6333 & n6334;
  assign n6336 = pi824 & pi1093;
  assign n6337 = n6102 & n6336;
  assign n6338 = n6335 & n6337;
  assign n6339 = ~pi829 & ~n2921;
  assign n6340 = pi1091 & ~n6339;
  assign n6341 = n6338 & ~n6340;
  assign n6342 = ~pi216 & ~n6341;
  assign n6343 = ~pi1091 & n6338;
  assign n6344 = pi1091 & n2921;
  assign n6345 = n6337 & ~n6344;
  assign n6346 = ~n2926 & ~n6345;
  assign n6347 = pi1091 & ~n6346;
  assign n6348 = n6335 & n6347;
  assign n6349 = ~n6343 & ~n6348;
  assign n6350 = pi216 & n6349;
  assign n6351 = ~n6342 & ~n6350;
  assign n6352 = ~pi228 & n6351;
  assign n6353 = ~n6265 & ~n6352;
  assign n6354 = n5726 & ~n6353;
  assign n6355 = ~n6265 & ~n6354;
  assign n6356 = n6263 & ~n6355;
  assign n6357 = pi299 & ~n6356;
  assign n6358 = pi224 & n6349;
  assign n6359 = pi222 & ~pi223;
  assign n6360 = ~pi224 & ~n6341;
  assign n6361 = n6359 & ~n6360;
  assign n6362 = ~n6358 & n6361;
  assign n6363 = ~pi228 & n6362;
  assign n6364 = ~n6265 & ~n6363;
  assign n6365 = n6279 & ~n6364;
  assign n6366 = ~pi299 & ~n6365;
  assign n6367 = pi39 & ~n6366;
  assign n6368 = ~n6357 & n6367;
  assign n6369 = pi158 & pi159;
  assign n6370 = pi160 & pi197;
  assign n6371 = n6369 & n6370;
  assign n6372 = ~pi91 & pi314;
  assign n6373 = n2765 & ~n2766;
  assign n6374 = pi85 & n2825;
  assign n6375 = n2481 & ~n6374;
  assign n6376 = n2829 & ~n6375;
  assign n6377 = n2477 & ~n6376;
  assign n6378 = ~n2809 & ~n2834;
  assign n6379 = ~n6377 & n6378;
  assign n6380 = n2478 & n6379;
  assign n6381 = ~n2806 & ~n6380;
  assign n6382 = n2803 & ~n6381;
  assign n6383 = pi67 & n2483;
  assign n6384 = n2484 & ~n6383;
  assign n6385 = ~n6382 & n6384;
  assign n6386 = n2796 & ~n6385;
  assign n6387 = ~pi71 & ~n6386;
  assign po1049 = pi64 | ~n2489;
  assign n6389 = n2789 & ~po1049;
  assign n6390 = ~n6387 & n6389;
  assign n6391 = ~pi81 & ~n6390;
  assign n6392 = ~pi102 & ~n2784;
  assign n6393 = n2465 & n6392;
  assign n6394 = ~n6391 & n6393;
  assign n6395 = n2783 & ~n6394;
  assign n6396 = n2877 & ~n6395;
  assign n6397 = n2719 & ~n6396;
  assign n6398 = ~n2722 & ~n6397;
  assign n6399 = ~pi86 & ~n6398;
  assign n6400 = n2498 & n2780;
  assign n6401 = ~n6399 & n6400;
  assign n6402 = n2890 & ~n6401;
  assign n6403 = n6373 & ~n6402;
  assign n6404 = n6372 & ~n6403;
  assign n6405 = ~pi91 & ~pi314;
  assign n6406 = n2844 & n6389;
  assign n6407 = n6391 & ~n6406;
  assign n6408 = n6393 & ~n6407;
  assign n6409 = n2783 & ~n6408;
  assign n6410 = n2877 & ~n6409;
  assign n6411 = n2719 & ~n6410;
  assign n6412 = ~n2722 & ~n6411;
  assign n6413 = ~pi86 & ~n6412;
  assign n6414 = n6400 & ~n6413;
  assign n6415 = n2890 & ~n6414;
  assign n6416 = n6373 & ~n6415;
  assign n6417 = n6405 & ~n6416;
  assign n6418 = ~pi58 & n2756;
  assign n6419 = ~n2705 & ~n6418;
  assign n6420 = ~n6404 & ~n6419;
  assign n6421 = ~n6417 & n6420;
  assign n6422 = ~pi90 & ~n6421;
  assign n6423 = ~n2897 & ~n6422;
  assign n6424 = ~pi93 & ~n6423;
  assign n6425 = pi93 & ~n2914;
  assign n6426 = ~pi35 & ~n6425;
  assign n6427 = ~n6424 & n6426;
  assign n6428 = ~pi70 & ~n6427;
  assign n6429 = n3082 & ~n6428;
  assign n6430 = ~pi72 & ~n6429;
  assign n6431 = ~pi95 & n2462;
  assign n6432 = ~n2744 & n6431;
  assign n6433 = ~n6430 & n6432;
  assign n6434 = ~n3162 & ~n6433;
  assign n6435 = ~pi841 & n2506;
  assign n6436 = n2509 & n6435;
  assign n6437 = n2735 & n6436;
  assign n6438 = pi32 & n6437;
  assign n6439 = ~pi95 & n6438;
  assign n6440 = ~pi210 & n6439;
  assign n6441 = n6434 & ~n6440;
  assign n6442 = ~n6166 & ~n6441;
  assign n6443 = ~pi47 & n2496;
  assign n6444 = ~n2889 & ~n6414;
  assign n6445 = n6443 & ~n6444;
  assign n6446 = n6405 & ~n6445;
  assign n6447 = ~n2889 & ~n6401;
  assign n6448 = n6443 & ~n6447;
  assign n6449 = n6372 & ~n6448;
  assign n6450 = ~n6419 & ~n6449;
  assign n6451 = ~n6446 & n6450;
  assign n6452 = ~pi90 & ~n6451;
  assign n6453 = ~n2897 & ~n6452;
  assign n6454 = ~pi93 & ~n6453;
  assign n6455 = n6426 & ~n6454;
  assign n6456 = ~pi70 & ~n6455;
  assign n6457 = n3082 & ~n6456;
  assign n6458 = ~pi72 & ~n6457;
  assign n6459 = n6432 & ~n6458;
  assign n6460 = ~n3162 & ~n6459;
  assign n6461 = ~n6440 & n6460;
  assign n6462 = n6166 & ~n6461;
  assign n6463 = ~n6442 & ~n6462;
  assign n6464 = n6263 & ~n6463;
  assign n6465 = n6371 & ~n6464;
  assign n6466 = n6263 & ~n6441;
  assign n6467 = ~n6371 & ~n6466;
  assign n6468 = ~pi228 & ~n6467;
  assign n6469 = ~n6465 & n6468;
  assign n6470 = n6303 & ~n6469;
  assign n6471 = ~pi198 & n6439;
  assign n6472 = n6434 & ~n6471;
  assign n6473 = ~pi228 & ~n6472;
  assign n6474 = ~n6265 & ~n6473;
  assign n6475 = n6279 & ~n6474;
  assign n6476 = ~pi299 & ~n6475;
  assign n6477 = pi145 & pi180;
  assign n6478 = pi181 & pi182;
  assign n6479 = n6477 & n6478;
  assign n6480 = ~pi299 & n6479;
  assign n6481 = ~n6476 & ~n6480;
  assign n6482 = ~n6166 & ~n6472;
  assign n6483 = n6460 & ~n6471;
  assign n6484 = n6166 & ~n6483;
  assign n6485 = ~n6482 & ~n6484;
  assign n6486 = ~pi228 & n6279;
  assign n6487 = ~n6485 & n6486;
  assign n6488 = ~n6319 & ~n6487;
  assign n6489 = n6479 & ~n6488;
  assign n6490 = ~n6481 & ~n6489;
  assign n6491 = pi232 & ~n6470;
  assign n6492 = ~n6490 & n6491;
  assign n6493 = ~pi228 & n6466;
  assign n6494 = n6303 & ~n6493;
  assign n6495 = ~pi232 & ~n6494;
  assign n6496 = ~n6476 & n6495;
  assign n6497 = ~n6492 & ~n6496;
  assign n6498 = ~pi39 & ~n6497;
  assign n6499 = ~pi38 & ~n6368;
  assign n6500 = ~n6498 & n6499;
  assign n6501 = pi38 & ~n6282;
  assign n6502 = ~n6286 & n6501;
  assign n6503 = ~n6500 & ~n6502;
  assign n6504 = ~pi100 & ~n6503;
  assign n6505 = ~pi87 & ~n6332;
  assign n6506 = ~n6504 & n6505;
  assign n6507 = ~pi75 & ~n6301;
  assign n6508 = ~n6506 & n6507;
  assign n6509 = ~pi92 & ~n6300;
  assign n6510 = ~n6508 & n6509;
  assign n6511 = ~pi54 & ~n6299;
  assign n6512 = ~n6510 & n6511;
  assign n6513 = ~pi74 & ~n6295;
  assign n6514 = ~n6512 & n6513;
  assign n6515 = ~pi55 & ~n6292;
  assign n6516 = ~n6514 & n6515;
  assign n6517 = n2530 & ~n6275;
  assign n6518 = ~n6516 & n6517;
  assign n6519 = ~pi59 & ~n6274;
  assign n6520 = ~n6518 & n6519;
  assign n6521 = ~pi57 & ~n6272;
  assign n6522 = ~n6520 & n6521;
  assign po171 = ~n6269 & ~n6522;
  assign n6524 = ~pi947 & n6166;
  assign n6525 = ~n6196 & ~n6524;
  assign n6526 = n6267 & n6525;
  assign n6527 = n6260 & n6526;
  assign n6528 = ~n6270 & n6526;
  assign n6529 = pi59 & ~n6528;
  assign n6530 = n6265 & n6525;
  assign n6531 = ~n2530 & n6530;
  assign n6532 = pi55 & ~n6526;
  assign n6533 = pi299 & ~n6525;
  assign n6534 = ~pi587 & n6166;
  assign n6535 = ~n6196 & ~n6534;
  assign n6536 = ~pi299 & ~n6535;
  assign n6537 = ~n6533 & ~n6536;
  assign n6538 = n6265 & n6537;
  assign n6539 = ~n6276 & ~n6538;
  assign n6540 = ~n2615 & n6538;
  assign n6541 = n6285 & n6537;
  assign n6542 = n2574 & n6541;
  assign n6543 = ~n6540 & ~n6542;
  assign n6544 = n2572 & n6543;
  assign n6545 = ~pi54 & n6544;
  assign n6546 = pi74 & ~n6539;
  assign n6547 = ~n6545 & n6546;
  assign n6548 = ~n2572 & ~n6538;
  assign n6549 = ~n6544 & ~n6548;
  assign n6550 = pi54 & ~n6549;
  assign n6551 = ~pi75 & n6543;
  assign n6552 = pi75 & ~n6538;
  assign n6553 = pi92 & ~n6552;
  assign n6554 = ~n6551 & n6553;
  assign n6555 = pi75 & n6543;
  assign n6556 = pi87 & n6538;
  assign n6557 = ~n2531 & n6538;
  assign n6558 = pi299 & ~n6530;
  assign n6559 = ~n6196 & n6312;
  assign n6560 = n2666 & ~n6524;
  assign n6561 = n6559 & n6560;
  assign n6562 = ~n6161 & n6304;
  assign n6563 = n6161 & n6306;
  assign n6564 = ~n6562 & ~n6563;
  assign n6565 = n6161 & ~n6166;
  assign n6566 = ~pi947 & ~n6565;
  assign n6567 = ~n2666 & ~n6566;
  assign n6568 = ~n6564 & n6567;
  assign n6569 = ~n6561 & ~n6568;
  assign n6570 = ~pi228 & ~n6569;
  assign n6571 = n6558 & ~n6570;
  assign n6572 = ~pi228 & n2641;
  assign n6573 = ~n6534 & ~n6564;
  assign n6574 = n6572 & ~n6573;
  assign n6575 = pi142 & n6564;
  assign n6576 = ~pi142 & ~n6559;
  assign n6577 = ~pi587 & ~n6565;
  assign n6578 = ~pi228 & ~n6577;
  assign n6579 = ~n6576 & n6578;
  assign n6580 = ~n6575 & n6579;
  assign n6581 = n6265 & n6535;
  assign n6582 = ~n6572 & ~n6581;
  assign n6583 = ~n6580 & n6582;
  assign n6584 = ~n6574 & ~n6583;
  assign n6585 = ~pi299 & ~n6584;
  assign n6586 = n2531 & ~n6571;
  assign n6587 = ~n6585 & n6586;
  assign n6588 = pi100 & ~n6557;
  assign n6589 = ~n6587 & n6588;
  assign n6590 = pi299 & n5726;
  assign n6591 = ~n6558 & ~n6590;
  assign n6592 = n6354 & n6525;
  assign n6593 = ~n6591 & ~n6592;
  assign n6594 = ~n6364 & n6535;
  assign n6595 = ~pi299 & ~n6594;
  assign n6596 = pi39 & ~n6595;
  assign n6597 = ~n6593 & n6596;
  assign n6598 = ~n6463 & n6525;
  assign n6599 = n6371 & ~n6598;
  assign n6600 = ~n6441 & n6525;
  assign n6601 = ~n6371 & ~n6600;
  assign n6602 = ~pi228 & ~n6601;
  assign n6603 = ~n6599 & n6602;
  assign n6604 = n6558 & ~n6603;
  assign n6605 = ~n6474 & n6535;
  assign n6606 = ~n6479 & n6605;
  assign n6607 = ~pi228 & n6535;
  assign n6608 = ~n6485 & n6607;
  assign n6609 = ~n6581 & ~n6608;
  assign n6610 = n6479 & ~n6609;
  assign n6611 = ~pi299 & ~n6606;
  assign n6612 = ~n6610 & n6611;
  assign n6613 = pi232 & ~n6604;
  assign n6614 = ~n6612 & n6613;
  assign n6615 = ~pi228 & n6600;
  assign n6616 = n6558 & ~n6615;
  assign n6617 = ~pi299 & ~n6605;
  assign n6618 = ~pi232 & ~n6616;
  assign n6619 = ~n6617 & n6618;
  assign n6620 = ~n6614 & ~n6619;
  assign n6621 = ~pi39 & ~n6620;
  assign n6622 = ~pi38 & ~n6597;
  assign n6623 = ~n6621 & n6622;
  assign n6624 = pi38 & ~n6538;
  assign n6625 = ~n6541 & n6624;
  assign n6626 = ~n6623 & ~n6625;
  assign n6627 = ~pi100 & ~n6626;
  assign n6628 = ~pi87 & ~n6589;
  assign n6629 = ~n6627 & n6628;
  assign n6630 = ~pi75 & ~n6556;
  assign n6631 = ~n6629 & n6630;
  assign n6632 = ~pi92 & ~n6555;
  assign n6633 = ~n6631 & n6632;
  assign n6634 = ~pi54 & ~n6554;
  assign n6635 = ~n6633 & n6634;
  assign n6636 = ~pi74 & ~n6550;
  assign n6637 = ~n6635 & n6636;
  assign n6638 = ~pi55 & ~n6547;
  assign n6639 = ~n6637 & n6638;
  assign n6640 = n2530 & ~n6532;
  assign n6641 = ~n6639 & n6640;
  assign n6642 = ~pi59 & ~n6531;
  assign n6643 = ~n6641 & n6642;
  assign n6644 = ~pi57 & ~n6529;
  assign n6645 = ~n6643 & n6644;
  assign po172 = ~n6527 & ~n6645;
  assign n6647 = n6166 & n6265;
  assign n6648 = pi970 & n6647;
  assign n6649 = ~pi228 & pi970;
  assign n6650 = n2577 & n6185;
  assign n6651 = n6649 & n6650;
  assign n6652 = n6258 & n6651;
  assign n6653 = ~n6648 & ~n6652;
  assign n6654 = pi57 & ~n6653;
  assign n6655 = n6257 & n6651;
  assign n6656 = pi59 & ~n6648;
  assign n6657 = ~n6655 & n6656;
  assign n6658 = ~n2530 & n6648;
  assign n6659 = pi55 & ~n6648;
  assign n6660 = ~n6651 & n6659;
  assign n6661 = pi299 & pi970;
  assign n6662 = ~pi299 & pi967;
  assign n6663 = ~n6661 & ~n6662;
  assign n6664 = n6647 & ~n6663;
  assign n6665 = ~n6276 & ~n6664;
  assign n6666 = ~n2615 & n6664;
  assign n6667 = pi228 & ~n6647;
  assign n6668 = ~pi228 & ~n6185;
  assign n6669 = ~n6667 & ~n6668;
  assign n6670 = ~pi39 & n6669;
  assign n6671 = ~n6663 & n6670;
  assign n6672 = n2574 & n6671;
  assign n6673 = ~n6666 & ~n6672;
  assign n6674 = n2572 & n6673;
  assign n6675 = ~pi54 & n6674;
  assign n6676 = pi74 & ~n6665;
  assign n6677 = ~n6675 & n6676;
  assign n6678 = ~n2572 & ~n6664;
  assign n6679 = ~n6674 & ~n6678;
  assign n6680 = pi54 & ~n6679;
  assign n6681 = ~pi75 & n6673;
  assign n6682 = pi75 & ~n6664;
  assign n6683 = pi92 & ~n6682;
  assign n6684 = ~n6681 & n6683;
  assign n6685 = pi75 & n6673;
  assign n6686 = pi87 & n6664;
  assign n6687 = ~n2531 & n6664;
  assign n6688 = pi299 & ~n6648;
  assign n6689 = ~n2666 & ~n6304;
  assign n6690 = n6166 & n6312;
  assign n6691 = n2666 & ~n6690;
  assign n6692 = ~pi228 & ~n6689;
  assign n6693 = ~n6691 & n6692;
  assign n6694 = pi970 & n6693;
  assign n6695 = n6688 & ~n6694;
  assign n6696 = n6320 & n6690;
  assign n6697 = n6304 & ~n6320;
  assign n6698 = ~pi228 & ~n6696;
  assign n6699 = ~n6697 & n6698;
  assign n6700 = ~n6667 & ~n6699;
  assign n6701 = pi967 & n6700;
  assign n6702 = ~pi299 & ~n6701;
  assign n6703 = n2531 & ~n6695;
  assign n6704 = ~n6702 & n6703;
  assign n6705 = pi100 & ~n6687;
  assign n6706 = ~n6704 & n6705;
  assign n6707 = n5726 & n6351;
  assign n6708 = n6166 & n6707;
  assign n6709 = ~pi228 & ~n6708;
  assign n6710 = n6661 & ~n6709;
  assign n6711 = n6166 & n6362;
  assign n6712 = ~pi228 & ~n6711;
  assign n6713 = n6662 & ~n6712;
  assign n6714 = ~n6710 & ~n6713;
  assign n6715 = pi39 & ~n6667;
  assign n6716 = ~n6714 & n6715;
  assign n6717 = n6166 & ~n6474;
  assign n6718 = ~n6479 & ~n6717;
  assign n6719 = ~n6472 & ~n6479;
  assign n6720 = ~pi228 & n6484;
  assign n6721 = ~n6647 & ~n6719;
  assign n6722 = ~n6720 & n6721;
  assign n6723 = ~n6718 & ~n6722;
  assign n6724 = pi967 & n6723;
  assign n6725 = ~pi299 & ~n6724;
  assign n6726 = n6166 & ~n6441;
  assign n6727 = n6649 & n6726;
  assign n6728 = n6688 & ~n6727;
  assign n6729 = pi299 & n6369;
  assign n6730 = ~n6728 & ~n6729;
  assign n6731 = n6370 & ~n6462;
  assign n6732 = ~n6370 & n6441;
  assign n6733 = ~n6731 & ~n6732;
  assign n6734 = n6166 & n6733;
  assign n6735 = n6649 & n6734;
  assign n6736 = ~n6648 & ~n6735;
  assign n6737 = n6369 & ~n6736;
  assign n6738 = ~n6730 & ~n6737;
  assign n6739 = pi232 & ~n6725;
  assign n6740 = ~n6738 & n6739;
  assign n6741 = pi967 & n6717;
  assign n6742 = ~pi299 & ~n6741;
  assign n6743 = ~pi232 & ~n6728;
  assign n6744 = ~n6742 & n6743;
  assign n6745 = ~n6740 & ~n6744;
  assign n6746 = ~pi39 & ~n6745;
  assign n6747 = ~pi38 & ~n6716;
  assign n6748 = ~n6746 & n6747;
  assign n6749 = pi39 & n6664;
  assign n6750 = pi38 & ~n6749;
  assign n6751 = ~n6671 & n6750;
  assign n6752 = ~n6748 & ~n6751;
  assign n6753 = ~pi100 & ~n6752;
  assign n6754 = ~pi87 & ~n6706;
  assign n6755 = ~n6753 & n6754;
  assign n6756 = ~pi75 & ~n6686;
  assign n6757 = ~n6755 & n6756;
  assign n6758 = ~pi92 & ~n6685;
  assign n6759 = ~n6757 & n6758;
  assign n6760 = ~pi54 & ~n6684;
  assign n6761 = ~n6759 & n6760;
  assign n6762 = ~pi74 & ~n6680;
  assign n6763 = ~n6761 & n6762;
  assign n6764 = ~pi55 & ~n6677;
  assign n6765 = ~n6763 & n6764;
  assign n6766 = n2530 & ~n6660;
  assign n6767 = ~n6765 & n6766;
  assign n6768 = ~pi59 & ~n6658;
  assign n6769 = ~n6767 & n6768;
  assign n6770 = ~pi57 & ~n6657;
  assign n6771 = ~n6769 & n6770;
  assign po173 = ~n6654 & ~n6771;
  assign n6773 = pi972 & n6647;
  assign n6774 = ~pi228 & pi972;
  assign n6775 = n6650 & n6774;
  assign n6776 = n6258 & n6775;
  assign n6777 = ~n6773 & ~n6776;
  assign n6778 = pi57 & ~n6777;
  assign n6779 = n6257 & n6775;
  assign n6780 = pi59 & ~n6773;
  assign n6781 = ~n6779 & n6780;
  assign n6782 = ~n2530 & n6773;
  assign n6783 = pi55 & ~n6773;
  assign n6784 = ~n6775 & n6783;
  assign n6785 = ~pi299 & pi961;
  assign n6786 = pi299 & pi972;
  assign n6787 = ~n6785 & ~n6786;
  assign n6788 = n6647 & ~n6787;
  assign n6789 = ~n6276 & ~n6788;
  assign n6790 = ~n2615 & n6788;
  assign n6791 = n6670 & ~n6787;
  assign n6792 = n2574 & n6791;
  assign n6793 = ~n6790 & ~n6792;
  assign n6794 = n2572 & n6793;
  assign n6795 = ~pi54 & n6794;
  assign n6796 = pi74 & ~n6789;
  assign n6797 = ~n6795 & n6796;
  assign n6798 = ~n2572 & ~n6788;
  assign n6799 = ~n6794 & ~n6798;
  assign n6800 = pi54 & ~n6799;
  assign n6801 = ~pi75 & n6793;
  assign n6802 = pi75 & ~n6788;
  assign n6803 = pi92 & ~n6802;
  assign n6804 = ~n6801 & n6803;
  assign n6805 = pi75 & n6793;
  assign n6806 = pi87 & n6788;
  assign n6807 = ~n2531 & n6788;
  assign n6808 = pi299 & ~n6773;
  assign n6809 = pi972 & n6693;
  assign n6810 = n6808 & ~n6809;
  assign n6811 = pi961 & n6700;
  assign n6812 = ~pi299 & ~n6811;
  assign n6813 = n2531 & ~n6810;
  assign n6814 = ~n6812 & n6813;
  assign n6815 = pi100 & ~n6807;
  assign n6816 = ~n6814 & n6815;
  assign n6817 = ~n6712 & n6785;
  assign n6818 = ~n6709 & n6786;
  assign n6819 = ~n6817 & ~n6818;
  assign n6820 = n6715 & ~n6819;
  assign n6821 = pi961 & n6723;
  assign n6822 = ~pi299 & ~n6821;
  assign n6823 = n6726 & n6774;
  assign n6824 = n6808 & ~n6823;
  assign n6825 = ~n6729 & ~n6824;
  assign n6826 = n6734 & n6774;
  assign n6827 = ~n6773 & ~n6826;
  assign n6828 = n6369 & ~n6827;
  assign n6829 = ~n6825 & ~n6828;
  assign n6830 = pi232 & ~n6822;
  assign n6831 = ~n6829 & n6830;
  assign n6832 = pi961 & n6717;
  assign n6833 = ~pi299 & ~n6832;
  assign n6834 = ~pi232 & ~n6824;
  assign n6835 = ~n6833 & n6834;
  assign n6836 = ~n6831 & ~n6835;
  assign n6837 = ~pi39 & ~n6836;
  assign n6838 = ~pi38 & ~n6820;
  assign n6839 = ~n6837 & n6838;
  assign n6840 = pi39 & n6788;
  assign n6841 = pi38 & ~n6840;
  assign n6842 = ~n6791 & n6841;
  assign n6843 = ~n6839 & ~n6842;
  assign n6844 = ~pi100 & ~n6843;
  assign n6845 = ~pi87 & ~n6816;
  assign n6846 = ~n6844 & n6845;
  assign n6847 = ~pi75 & ~n6806;
  assign n6848 = ~n6846 & n6847;
  assign n6849 = ~pi92 & ~n6805;
  assign n6850 = ~n6848 & n6849;
  assign n6851 = ~pi54 & ~n6804;
  assign n6852 = ~n6850 & n6851;
  assign n6853 = ~pi74 & ~n6800;
  assign n6854 = ~n6852 & n6853;
  assign n6855 = ~pi55 & ~n6797;
  assign n6856 = ~n6854 & n6855;
  assign n6857 = n2530 & ~n6784;
  assign n6858 = ~n6856 & n6857;
  assign n6859 = ~pi59 & ~n6782;
  assign n6860 = ~n6858 & n6859;
  assign n6861 = ~pi57 & ~n6781;
  assign n6862 = ~n6860 & n6861;
  assign po174 = ~n6778 & ~n6862;
  assign n6864 = pi960 & n6647;
  assign n6865 = ~pi228 & pi960;
  assign n6866 = n6650 & n6865;
  assign n6867 = n6258 & n6866;
  assign n6868 = ~n6864 & ~n6867;
  assign n6869 = pi57 & ~n6868;
  assign n6870 = n6257 & n6866;
  assign n6871 = pi59 & ~n6864;
  assign n6872 = ~n6870 & n6871;
  assign n6873 = ~n2530 & n6864;
  assign n6874 = pi55 & ~n6864;
  assign n6875 = ~n6866 & n6874;
  assign n6876 = ~pi299 & pi977;
  assign n6877 = pi299 & pi960;
  assign n6878 = ~n6876 & ~n6877;
  assign n6879 = n6647 & ~n6878;
  assign n6880 = ~n6276 & ~n6879;
  assign n6881 = ~n2615 & n6879;
  assign n6882 = n6670 & ~n6878;
  assign n6883 = n2574 & n6882;
  assign n6884 = ~n6881 & ~n6883;
  assign n6885 = n2572 & n6884;
  assign n6886 = ~pi54 & n6885;
  assign n6887 = pi74 & ~n6880;
  assign n6888 = ~n6886 & n6887;
  assign n6889 = ~n2572 & ~n6879;
  assign n6890 = ~n6885 & ~n6889;
  assign n6891 = pi54 & ~n6890;
  assign n6892 = ~pi75 & n6884;
  assign n6893 = pi75 & ~n6879;
  assign n6894 = pi92 & ~n6893;
  assign n6895 = ~n6892 & n6894;
  assign n6896 = pi75 & n6884;
  assign n6897 = pi87 & n6879;
  assign n6898 = ~n2531 & n6879;
  assign n6899 = pi299 & ~n6864;
  assign n6900 = pi960 & n6693;
  assign n6901 = n6899 & ~n6900;
  assign n6902 = pi977 & n6700;
  assign n6903 = ~pi299 & ~n6902;
  assign n6904 = n2531 & ~n6901;
  assign n6905 = ~n6903 & n6904;
  assign n6906 = pi100 & ~n6898;
  assign n6907 = ~n6905 & n6906;
  assign n6908 = ~n6712 & n6876;
  assign n6909 = ~n6709 & n6877;
  assign n6910 = ~n6908 & ~n6909;
  assign n6911 = n6715 & ~n6910;
  assign n6912 = pi977 & n6723;
  assign n6913 = ~pi299 & ~n6912;
  assign n6914 = n6726 & n6865;
  assign n6915 = n6899 & ~n6914;
  assign n6916 = ~n6729 & ~n6915;
  assign n6917 = n6734 & n6865;
  assign n6918 = ~n6864 & ~n6917;
  assign n6919 = n6369 & ~n6918;
  assign n6920 = ~n6916 & ~n6919;
  assign n6921 = pi232 & ~n6913;
  assign n6922 = ~n6920 & n6921;
  assign n6923 = pi977 & n6717;
  assign n6924 = ~pi299 & ~n6923;
  assign n6925 = ~pi232 & ~n6915;
  assign n6926 = ~n6924 & n6925;
  assign n6927 = ~n6922 & ~n6926;
  assign n6928 = ~pi39 & ~n6927;
  assign n6929 = ~pi38 & ~n6911;
  assign n6930 = ~n6928 & n6929;
  assign n6931 = pi39 & n6879;
  assign n6932 = pi38 & ~n6931;
  assign n6933 = ~n6882 & n6932;
  assign n6934 = ~n6930 & ~n6933;
  assign n6935 = ~pi100 & ~n6934;
  assign n6936 = ~pi87 & ~n6907;
  assign n6937 = ~n6935 & n6936;
  assign n6938 = ~pi75 & ~n6897;
  assign n6939 = ~n6937 & n6938;
  assign n6940 = ~pi92 & ~n6896;
  assign n6941 = ~n6939 & n6940;
  assign n6942 = ~pi54 & ~n6895;
  assign n6943 = ~n6941 & n6942;
  assign n6944 = ~pi74 & ~n6891;
  assign n6945 = ~n6943 & n6944;
  assign n6946 = ~pi55 & ~n6888;
  assign n6947 = ~n6945 & n6946;
  assign n6948 = n2530 & ~n6875;
  assign n6949 = ~n6947 & n6948;
  assign n6950 = ~pi59 & ~n6873;
  assign n6951 = ~n6949 & n6950;
  assign n6952 = ~pi57 & ~n6872;
  assign n6953 = ~n6951 & n6952;
  assign po175 = ~n6869 & ~n6953;
  assign n6955 = pi963 & n6647;
  assign n6956 = ~pi228 & pi963;
  assign n6957 = n6650 & n6956;
  assign n6958 = n6258 & n6957;
  assign n6959 = ~n6955 & ~n6958;
  assign n6960 = pi57 & ~n6959;
  assign n6961 = n6257 & n6957;
  assign n6962 = pi59 & ~n6955;
  assign n6963 = ~n6961 & n6962;
  assign n6964 = ~n2530 & n6955;
  assign n6965 = pi55 & ~n6955;
  assign n6966 = ~n6957 & n6965;
  assign n6967 = ~pi299 & pi969;
  assign n6968 = pi299 & pi963;
  assign n6969 = ~n6967 & ~n6968;
  assign n6970 = n6647 & ~n6969;
  assign n6971 = ~n6276 & ~n6970;
  assign n6972 = ~n2615 & n6970;
  assign n6973 = n6670 & ~n6969;
  assign n6974 = n2574 & n6973;
  assign n6975 = ~n6972 & ~n6974;
  assign n6976 = n2572 & n6975;
  assign n6977 = ~pi54 & n6976;
  assign n6978 = pi74 & ~n6971;
  assign n6979 = ~n6977 & n6978;
  assign n6980 = ~n2572 & ~n6970;
  assign n6981 = ~n6976 & ~n6980;
  assign n6982 = pi54 & ~n6981;
  assign n6983 = ~pi75 & n6975;
  assign n6984 = pi75 & ~n6970;
  assign n6985 = pi92 & ~n6984;
  assign n6986 = ~n6983 & n6985;
  assign n6987 = pi75 & n6975;
  assign n6988 = pi87 & n6970;
  assign n6989 = ~n2531 & n6970;
  assign n6990 = pi299 & ~n6955;
  assign n6991 = pi963 & n6693;
  assign n6992 = n6990 & ~n6991;
  assign n6993 = pi969 & n6700;
  assign n6994 = ~pi299 & ~n6993;
  assign n6995 = n2531 & ~n6992;
  assign n6996 = ~n6994 & n6995;
  assign n6997 = pi100 & ~n6989;
  assign n6998 = ~n6996 & n6997;
  assign n6999 = ~n6712 & n6967;
  assign n7000 = ~n6709 & n6968;
  assign n7001 = ~n6999 & ~n7000;
  assign n7002 = n6715 & ~n7001;
  assign n7003 = pi969 & n6723;
  assign n7004 = ~pi299 & ~n7003;
  assign n7005 = n6726 & n6956;
  assign n7006 = n6990 & ~n7005;
  assign n7007 = ~n6729 & ~n7006;
  assign n7008 = n6734 & n6956;
  assign n7009 = ~n6955 & ~n7008;
  assign n7010 = n6369 & ~n7009;
  assign n7011 = ~n7007 & ~n7010;
  assign n7012 = pi232 & ~n7004;
  assign n7013 = ~n7011 & n7012;
  assign n7014 = pi969 & n6717;
  assign n7015 = ~pi299 & ~n7014;
  assign n7016 = ~pi232 & ~n7006;
  assign n7017 = ~n7015 & n7016;
  assign n7018 = ~n7013 & ~n7017;
  assign n7019 = ~pi39 & ~n7018;
  assign n7020 = ~pi38 & ~n7002;
  assign n7021 = ~n7019 & n7020;
  assign n7022 = pi39 & n6970;
  assign n7023 = pi38 & ~n7022;
  assign n7024 = ~n6973 & n7023;
  assign n7025 = ~n7021 & ~n7024;
  assign n7026 = ~pi100 & ~n7025;
  assign n7027 = ~pi87 & ~n6998;
  assign n7028 = ~n7026 & n7027;
  assign n7029 = ~pi75 & ~n6988;
  assign n7030 = ~n7028 & n7029;
  assign n7031 = ~pi92 & ~n6987;
  assign n7032 = ~n7030 & n7031;
  assign n7033 = ~pi54 & ~n6986;
  assign n7034 = ~n7032 & n7033;
  assign n7035 = ~pi74 & ~n6982;
  assign n7036 = ~n7034 & n7035;
  assign n7037 = ~pi55 & ~n6979;
  assign n7038 = ~n7036 & n7037;
  assign n7039 = n2530 & ~n6966;
  assign n7040 = ~n7038 & n7039;
  assign n7041 = ~pi59 & ~n6964;
  assign n7042 = ~n7040 & n7041;
  assign n7043 = ~pi57 & ~n6963;
  assign n7044 = ~n7042 & n7043;
  assign po176 = ~n6960 & ~n7044;
  assign n7046 = pi975 & n6647;
  assign n7047 = ~pi228 & pi975;
  assign n7048 = n6650 & n7047;
  assign n7049 = n6258 & n7048;
  assign n7050 = ~n7046 & ~n7049;
  assign n7051 = pi57 & ~n7050;
  assign n7052 = n6257 & n7048;
  assign n7053 = pi59 & ~n7046;
  assign n7054 = ~n7052 & n7053;
  assign n7055 = ~n2530 & n7046;
  assign n7056 = pi55 & ~n7046;
  assign n7057 = ~n7048 & n7056;
  assign n7058 = ~pi299 & pi971;
  assign n7059 = pi299 & pi975;
  assign n7060 = ~n7058 & ~n7059;
  assign n7061 = n6647 & ~n7060;
  assign n7062 = ~n6276 & ~n7061;
  assign n7063 = ~n2615 & n7061;
  assign n7064 = n6670 & ~n7060;
  assign n7065 = n2574 & n7064;
  assign n7066 = ~n7063 & ~n7065;
  assign n7067 = n2572 & n7066;
  assign n7068 = ~pi54 & n7067;
  assign n7069 = pi74 & ~n7062;
  assign n7070 = ~n7068 & n7069;
  assign n7071 = ~n2572 & ~n7061;
  assign n7072 = ~n7067 & ~n7071;
  assign n7073 = pi54 & ~n7072;
  assign n7074 = ~pi75 & n7066;
  assign n7075 = pi75 & ~n7061;
  assign n7076 = pi92 & ~n7075;
  assign n7077 = ~n7074 & n7076;
  assign n7078 = pi75 & n7066;
  assign n7079 = pi87 & n7061;
  assign n7080 = ~n2531 & n7061;
  assign n7081 = pi299 & ~n7046;
  assign n7082 = pi975 & n6693;
  assign n7083 = n7081 & ~n7082;
  assign n7084 = pi971 & n6700;
  assign n7085 = ~pi299 & ~n7084;
  assign n7086 = n2531 & ~n7083;
  assign n7087 = ~n7085 & n7086;
  assign n7088 = pi100 & ~n7080;
  assign n7089 = ~n7087 & n7088;
  assign n7090 = ~n6712 & n7058;
  assign n7091 = ~n6709 & n7059;
  assign n7092 = ~n7090 & ~n7091;
  assign n7093 = n6715 & ~n7092;
  assign n7094 = pi971 & n6723;
  assign n7095 = ~pi299 & ~n7094;
  assign n7096 = n6726 & n7047;
  assign n7097 = n7081 & ~n7096;
  assign n7098 = ~n6729 & ~n7097;
  assign n7099 = n6734 & n7047;
  assign n7100 = ~n7046 & ~n7099;
  assign n7101 = n6369 & ~n7100;
  assign n7102 = ~n7098 & ~n7101;
  assign n7103 = pi232 & ~n7095;
  assign n7104 = ~n7102 & n7103;
  assign n7105 = pi971 & n6717;
  assign n7106 = ~pi299 & ~n7105;
  assign n7107 = ~pi232 & ~n7097;
  assign n7108 = ~n7106 & n7107;
  assign n7109 = ~n7104 & ~n7108;
  assign n7110 = ~pi39 & ~n7109;
  assign n7111 = ~pi38 & ~n7093;
  assign n7112 = ~n7110 & n7111;
  assign n7113 = pi39 & n7061;
  assign n7114 = pi38 & ~n7113;
  assign n7115 = ~n7064 & n7114;
  assign n7116 = ~n7112 & ~n7115;
  assign n7117 = ~pi100 & ~n7116;
  assign n7118 = ~pi87 & ~n7089;
  assign n7119 = ~n7117 & n7118;
  assign n7120 = ~pi75 & ~n7079;
  assign n7121 = ~n7119 & n7120;
  assign n7122 = ~pi92 & ~n7078;
  assign n7123 = ~n7121 & n7122;
  assign n7124 = ~pi54 & ~n7077;
  assign n7125 = ~n7123 & n7124;
  assign n7126 = ~pi74 & ~n7073;
  assign n7127 = ~n7125 & n7126;
  assign n7128 = ~pi55 & ~n7070;
  assign n7129 = ~n7127 & n7128;
  assign n7130 = n2530 & ~n7057;
  assign n7131 = ~n7129 & n7130;
  assign n7132 = ~pi59 & ~n7055;
  assign n7133 = ~n7131 & n7132;
  assign n7134 = ~pi57 & ~n7054;
  assign n7135 = ~n7133 & n7134;
  assign po177 = ~n7051 & ~n7135;
  assign n7137 = pi978 & n6647;
  assign n7138 = ~pi228 & pi978;
  assign n7139 = n6650 & n7138;
  assign n7140 = n6258 & n7139;
  assign n7141 = ~n7137 & ~n7140;
  assign n7142 = pi57 & ~n7141;
  assign n7143 = n6257 & n7139;
  assign n7144 = pi59 & ~n7137;
  assign n7145 = ~n7143 & n7144;
  assign n7146 = ~n2530 & n7137;
  assign n7147 = pi55 & ~n7137;
  assign n7148 = ~n7139 & n7147;
  assign n7149 = ~pi299 & pi974;
  assign n7150 = pi299 & pi978;
  assign n7151 = ~n7149 & ~n7150;
  assign n7152 = n6647 & ~n7151;
  assign n7153 = ~n6276 & ~n7152;
  assign n7154 = n6669 & ~n7151;
  assign n7155 = ~pi228 & ~n2615;
  assign n7156 = n7154 & ~n7155;
  assign n7157 = n2572 & ~n7156;
  assign n7158 = ~pi54 & n7157;
  assign n7159 = pi74 & ~n7153;
  assign n7160 = ~n7158 & n7159;
  assign n7161 = ~n2572 & ~n7152;
  assign n7162 = ~n7157 & ~n7161;
  assign n7163 = pi54 & ~n7162;
  assign n7164 = ~pi75 & ~n7156;
  assign n7165 = pi75 & ~n7152;
  assign n7166 = pi92 & ~n7165;
  assign n7167 = ~n7164 & n7166;
  assign n7168 = pi75 & ~n7156;
  assign n7169 = pi87 & n7152;
  assign n7170 = ~n2531 & n7152;
  assign n7171 = pi299 & ~n7137;
  assign n7172 = pi978 & n6693;
  assign n7173 = n7171 & ~n7172;
  assign n7174 = pi974 & n6700;
  assign n7175 = ~pi299 & ~n7174;
  assign n7176 = n2531 & ~n7173;
  assign n7177 = ~n7175 & n7176;
  assign n7178 = pi100 & ~n7170;
  assign n7179 = ~n7177 & n7178;
  assign n7180 = pi39 & n7152;
  assign n7181 = ~pi39 & n7154;
  assign n7182 = pi38 & ~n7180;
  assign n7183 = ~n7181 & n7182;
  assign n7184 = ~n6712 & n7149;
  assign n7185 = ~n6709 & n7150;
  assign n7186 = ~n7184 & ~n7185;
  assign n7187 = n6715 & ~n7186;
  assign n7188 = pi974 & n6723;
  assign n7189 = ~pi299 & ~n7188;
  assign n7190 = n6726 & n7138;
  assign n7191 = n7171 & ~n7190;
  assign n7192 = ~n6729 & ~n7191;
  assign n7193 = n6734 & n7138;
  assign n7194 = ~n7137 & ~n7193;
  assign n7195 = n6369 & ~n7194;
  assign n7196 = ~n7192 & ~n7195;
  assign n7197 = pi232 & ~n7189;
  assign n7198 = ~n7196 & n7197;
  assign n7199 = pi974 & n6717;
  assign n7200 = ~pi299 & ~n7199;
  assign n7201 = ~pi232 & ~n7191;
  assign n7202 = ~n7200 & n7201;
  assign n7203 = ~n7198 & ~n7202;
  assign n7204 = ~pi39 & ~n7203;
  assign n7205 = ~pi38 & ~n7187;
  assign n7206 = ~n7204 & n7205;
  assign n7207 = ~n7183 & ~n7206;
  assign n7208 = ~pi100 & ~n7207;
  assign n7209 = ~pi87 & ~n7179;
  assign n7210 = ~n7208 & n7209;
  assign n7211 = ~pi75 & ~n7169;
  assign n7212 = ~n7210 & n7211;
  assign n7213 = ~pi92 & ~n7168;
  assign n7214 = ~n7212 & n7213;
  assign n7215 = ~pi54 & ~n7167;
  assign n7216 = ~n7214 & n7215;
  assign n7217 = ~pi74 & ~n7163;
  assign n7218 = ~n7216 & n7217;
  assign n7219 = ~pi55 & ~n7160;
  assign n7220 = ~n7218 & n7219;
  assign n7221 = n2530 & ~n7148;
  assign n7222 = ~n7220 & n7221;
  assign n7223 = ~pi59 & ~n7146;
  assign n7224 = ~n7222 & n7223;
  assign n7225 = ~pi57 & ~n7145;
  assign n7226 = ~n7224 & n7225;
  assign po178 = ~n7142 & ~n7226;
  assign n7228 = n2574 & n6081;
  assign n7229 = pi75 & ~n7228;
  assign n7230 = ~pi38 & ~pi87;
  assign n7231 = ~pi75 & ~pi100;
  assign n7232 = n7230 & n7231;
  assign n7233 = n6081 & n7232;
  assign n7234 = pi92 & ~n7233;
  assign n7235 = ~n7229 & ~n7234;
  assign n7236 = ~pi38 & n6081;
  assign n7237 = pi100 & ~n7236;
  assign n7238 = ~pi87 & ~n7237;
  assign n7239 = ~n6442 & n6729;
  assign n7240 = ~n6733 & n7239;
  assign n7241 = n6479 & n6484;
  assign n7242 = ~pi299 & ~n6482;
  assign n7243 = ~n6719 & n7242;
  assign n7244 = ~n7241 & n7243;
  assign n7245 = ~n7240 & ~n7244;
  assign n7246 = pi232 & ~n7245;
  assign n7247 = pi299 & n6441;
  assign n7248 = ~pi299 & n6472;
  assign n7249 = ~n7247 & ~n7248;
  assign n7250 = ~n6369 & n7247;
  assign n7251 = pi232 & ~n7250;
  assign n7252 = ~n7249 & ~n7251;
  assign n7253 = ~n7246 & ~n7252;
  assign n7254 = ~pi39 & ~n7253;
  assign n7255 = ~pi299 & ~n6207;
  assign n7256 = n6362 & n7255;
  assign n7257 = pi299 & ~n6223;
  assign n7258 = n6707 & n7257;
  assign n7259 = pi39 & ~n7256;
  assign n7260 = ~n7258 & n7259;
  assign n7261 = ~n7254 & ~n7260;
  assign n7262 = ~pi38 & ~n7261;
  assign n7263 = ~n6117 & ~n7262;
  assign n7264 = ~pi100 & ~n7263;
  assign n7265 = ~n6115 & n7238;
  assign n7266 = ~n7264 & n7265;
  assign n7267 = n2572 & ~n7266;
  assign n7268 = n7235 & ~n7267;
  assign n7269 = ~pi54 & ~n7268;
  assign n7270 = ~pi92 & n7233;
  assign n7271 = pi54 & ~n7270;
  assign n7272 = ~n7269 & ~n7271;
  assign n7273 = ~pi74 & ~n7272;
  assign n7274 = ~n6076 & ~n7273;
  assign n7275 = ~pi55 & ~n7274;
  assign n7276 = ~pi74 & n6075;
  assign n7277 = pi55 & ~n7276;
  assign n7278 = ~pi56 & ~n7277;
  assign n7279 = ~pi62 & n7278;
  assign n7280 = ~n7275 & n7279;
  assign n7281 = n3291 & ~n7280;
  assign po195 = n6071 & ~n7281;
  assign n7283 = ~pi954 & ~po195;
  assign n7284 = pi24 & pi954;
  assign po182 = ~n7283 & ~n7284;
  assign n7286 = n3317 & n3524;
  assign n7287 = ~n2441 & ~n7286;
  assign n7288 = pi62 & ~n7287;
  assign n7289 = n2532 & n3524;
  assign n7290 = n2537 & n7289;
  assign n7291 = pi56 & ~n2441;
  assign n7292 = ~n7290 & n7291;
  assign n7293 = n2533 & n2572;
  assign n7294 = n2531 & n3524;
  assign n7295 = n2573 & n7294;
  assign n7296 = n7293 & n7295;
  assign n7297 = ~n2441 & ~n7296;
  assign n7298 = pi55 & ~n7297;
  assign n7299 = ~n2441 & ~n2533;
  assign n7300 = ~pi75 & n7295;
  assign n7301 = ~n2441 & ~n7300;
  assign n7302 = pi92 & ~n7301;
  assign n7303 = pi75 & ~n2441;
  assign n7304 = ~n2441 & ~n7289;
  assign n7305 = pi87 & ~n7304;
  assign n7306 = ~pi100 & n4685;
  assign n7307 = n2523 & ~n6322;
  assign n7308 = ~pi299 & ~n7307;
  assign n7309 = pi299 & ~n3371;
  assign n7310 = ~n7308 & ~n7309;
  assign n7311 = pi100 & n3524;
  assign n7312 = n7310 & n7311;
  assign n7313 = ~pi39 & ~n7312;
  assign n7314 = ~n7306 & n7313;
  assign n7315 = ~pi100 & n3524;
  assign n7316 = pi39 & ~n7315;
  assign n7317 = ~pi38 & ~n7316;
  assign n7318 = ~n7314 & n7317;
  assign n7319 = ~n2441 & ~n7318;
  assign n7320 = ~pi87 & ~n7319;
  assign n7321 = ~pi75 & ~n7305;
  assign n7322 = ~n7320 & n7321;
  assign n7323 = ~pi92 & ~n7303;
  assign n7324 = ~n7322 & n7323;
  assign n7325 = n2533 & ~n7302;
  assign n7326 = ~n7324 & n7325;
  assign n7327 = ~pi55 & ~n7299;
  assign n7328 = ~n7326 & n7327;
  assign n7329 = ~pi56 & ~n7298;
  assign n7330 = ~n7328 & n7329;
  assign n7331 = ~pi62 & ~n7292;
  assign n7332 = ~n7330 & n7331;
  assign n7333 = ~n7288 & ~n7332;
  assign n7334 = n3291 & ~n7333;
  assign n7335 = n2441 & ~n3291;
  assign po183 = n7334 | n7335;
  assign n7337 = pi119 & pi1056;
  assign n7338 = ~pi228 & pi252;
  assign n7339 = ~pi119 & ~n7338;
  assign n7340 = ~pi468 & ~n7339;
  assign po184 = n7337 | ~n7340;
  assign n7342 = pi119 & pi1077;
  assign po185 = ~n7340 | n7342;
  assign n7344 = pi119 & pi1073;
  assign po186 = ~n7340 | n7344;
  assign n7346 = pi119 & pi1041;
  assign po187 = ~n7340 | n7346;
  assign n7348 = pi824 & n6102;
  assign n7349 = ~pi122 & pi1093;
  assign n7350 = n7348 & n7349;
  assign n7351 = ~pi1091 & n7350;
  assign n7352 = ~pi98 & n7351;
  assign n7353 = pi567 & n7352;
  assign n7354 = ~pi285 & ~pi286;
  assign n7355 = ~pi289 & n7354;
  assign n7356 = ~pi288 & n7355;
  assign po1038 = pi57 | ~n6258;
  assign n7358 = ~n7356 & po1038;
  assign n7359 = n7353 & n7358;
  assign n7360 = ~pi74 & n6078;
  assign n7361 = n2531 & n7231;
  assign n7362 = n2508 & ~n6138;
  assign n7363 = ~pi841 & n2708;
  assign n7364 = pi90 & n7363;
  assign n7365 = ~pi93 & ~n7364;
  assign n7366 = n7362 & ~n7365;
  assign n7367 = ~pi51 & ~n7366;
  assign n7368 = ~pi88 & pi98;
  assign n7369 = ~pi50 & ~pi77;
  assign n7370 = ~pi94 & n7369;
  assign n7371 = n2768 & n7370;
  assign n7372 = n2495 & n7368;
  assign n7373 = n7371 & n7372;
  assign n7374 = ~pi97 & ~n7373;
  assign n7375 = n2717 & ~n7374;
  assign n7376 = ~pi35 & n2709;
  assign n7377 = ~pi70 & n7376;
  assign n7378 = n7375 & n7377;
  assign n7379 = n7367 & ~n7378;
  assign n7380 = n2748 & n3174;
  assign n7381 = ~n7379 & n7380;
  assign n7382 = ~pi122 & pi829;
  assign n7383 = n6102 & n7382;
  assign n7384 = n7381 & ~n7383;
  assign n7385 = ~n2747 & ~n7379;
  assign n7386 = ~pi96 & ~n7385;
  assign n7387 = pi96 & ~n6436;
  assign n7388 = ~pi72 & n6431;
  assign n7389 = ~n7387 & n7388;
  assign n7390 = n7383 & n7389;
  assign n7391 = ~n7386 & n7390;
  assign n7392 = ~pi1093 & ~n7391;
  assign n7393 = ~n7384 & n7392;
  assign n7394 = ~pi72 & n7393;
  assign n7395 = ~pi1093 & ~n7394;
  assign n7396 = n6104 & n7381;
  assign n7397 = n7392 & ~n7396;
  assign n7398 = n7395 & ~n7397;
  assign n7399 = ~pi87 & ~n7398;
  assign n7400 = n2523 & po740;
  assign n7401 = pi87 & ~n7400;
  assign n7402 = n7361 & ~n7401;
  assign n7403 = ~n7399 & n7402;
  assign n7404 = ~pi567 & ~n7403;
  assign n7405 = n7360 & ~n7404;
  assign n7406 = pi232 & n6166;
  assign n7407 = n6086 & n7406;
  assign n7408 = n2615 & ~n7407;
  assign n7409 = n7352 & ~n7408;
  assign n7410 = ~n2921 & po1057;
  assign n7411 = pi1093 & n7383;
  assign n7412 = n7410 & n7411;
  assign n7413 = ~pi24 & n2523;
  assign n7414 = pi252 & n7413;
  assign n7415 = n7412 & n7414;
  assign n7416 = pi1091 & ~n7415;
  assign n7417 = n7408 & ~n7416;
  assign n7418 = ~pi122 & n7348;
  assign n7419 = ~pi98 & n7418;
  assign n7420 = pi1093 & n7419;
  assign n7421 = ~pi1091 & ~n7420;
  assign n7422 = n7417 & ~n7421;
  assign n7423 = pi75 & ~n7409;
  assign n7424 = ~n7422 & n7423;
  assign n7425 = pi1093 & n2921;
  assign n7426 = n6104 & ~n7425;
  assign n7427 = n2523 & n7426;
  assign n7428 = pi1091 & ~n7427;
  assign n7429 = ~pi1091 & ~n7400;
  assign n7430 = n2523 & n7348;
  assign n7431 = pi122 & n7430;
  assign n7432 = ~n7419 & ~n7431;
  assign n7433 = pi1093 & ~n7432;
  assign n7434 = n7429 & ~n7433;
  assign n7435 = n2628 & ~n7428;
  assign n7436 = ~n7434 & n7435;
  assign n7437 = ~n7352 & ~n7436;
  assign n7438 = pi87 & ~n7437;
  assign n7439 = ~n2531 & n7352;
  assign n7440 = pi228 & ~n7407;
  assign n7441 = ~n7352 & ~n7440;
  assign n7442 = pi1091 & n7412;
  assign n7443 = n2523 & n7442;
  assign n7444 = ~pi1091 & n7420;
  assign n7445 = n7440 & ~n7444;
  assign n7446 = ~n7443 & n7445;
  assign n7447 = n2531 & ~n7441;
  assign n7448 = ~n7446 & n7447;
  assign n7449 = pi100 & ~n7439;
  assign n7450 = ~n7448 & n7449;
  assign n7451 = pi38 & n7351;
  assign n7452 = ~pi98 & n7451;
  assign n7453 = pi1093 & ~n2921;
  assign n7454 = ~n7367 & n7380;
  assign n7455 = n7348 & n7454;
  assign n7456 = ~pi829 & n7455;
  assign n7457 = ~pi24 & n2756;
  assign n7458 = ~pi46 & n2496;
  assign n7459 = ~pi47 & pi97;
  assign n7460 = n7458 & n7459;
  assign n7461 = n2887 & n7460;
  assign n7462 = ~pi91 & n7461;
  assign n7463 = ~n7457 & ~n7462;
  assign n7464 = n2463 & n7362;
  assign n7465 = ~n7463 & n7464;
  assign n7466 = n7367 & ~n7465;
  assign n7467 = ~n2747 & ~n7466;
  assign n7468 = ~pi96 & ~n7467;
  assign n7469 = pi950 & n7389;
  assign n7470 = pi829 & pi1092;
  assign n7471 = n7469 & n7470;
  assign n7472 = ~n7468 & n7471;
  assign n7473 = ~n7456 & ~n7472;
  assign n7474 = ~pi122 & ~n7473;
  assign n7475 = pi122 & n6104;
  assign n7476 = n7454 & n7475;
  assign n7477 = ~n7474 & ~n7476;
  assign n7478 = n7453 & ~n7477;
  assign n7479 = pi1091 & ~n7478;
  assign n7480 = ~n7398 & n7479;
  assign n7481 = ~pi39 & ~n7480;
  assign n7482 = ~pi1091 & ~n7398;
  assign n7483 = pi122 & n7455;
  assign n7484 = ~n7419 & ~n7483;
  assign n7485 = pi1093 & ~n7484;
  assign n7486 = n7482 & ~n7485;
  assign n7487 = n7481 & ~n7486;
  assign n7488 = ~n5727 & n7352;
  assign n7489 = ~n6205 & ~n7352;
  assign n7490 = n2924 & n6335;
  assign n7491 = pi1092 & n7490;
  assign n7492 = n7453 & n7491;
  assign n7493 = pi1091 & ~n7492;
  assign n7494 = ~n7421 & ~n7493;
  assign n7495 = n6205 & ~n7494;
  assign n7496 = ~n7489 & ~n7495;
  assign n7497 = n6221 & ~n7496;
  assign n7498 = ~n6197 & n7494;
  assign n7499 = n6197 & n7352;
  assign n7500 = ~n7498 & ~n7499;
  assign n7501 = ~n6221 & n7500;
  assign n7502 = n5727 & ~n7497;
  assign n7503 = ~n7501 & n7502;
  assign n7504 = pi299 & ~n7488;
  assign n7505 = ~n7503 & n7504;
  assign n7506 = ~pi223 & n5754;
  assign n7507 = n7352 & ~n7506;
  assign n7508 = n6194 & ~n7496;
  assign n7509 = ~n6194 & n7500;
  assign n7510 = n7506 & ~n7508;
  assign n7511 = ~n7509 & n7510;
  assign n7512 = ~pi299 & ~n7507;
  assign n7513 = ~n7511 & n7512;
  assign n7514 = pi39 & ~n7505;
  assign n7515 = ~n7513 & n7514;
  assign n7516 = ~n7487 & ~n7515;
  assign n7517 = ~pi38 & ~n7516;
  assign n7518 = ~pi100 & ~n7452;
  assign n7519 = ~n7517 & n7518;
  assign n7520 = ~pi87 & ~n7450;
  assign n7521 = ~n7519 & n7520;
  assign n7522 = ~pi75 & ~n7438;
  assign n7523 = ~n7521 & n7522;
  assign n7524 = ~n7424 & ~n7523;
  assign n7525 = pi567 & ~n7524;
  assign n7526 = n7405 & ~n7525;
  assign n7527 = n7353 & ~n7360;
  assign n7528 = ~n7526 & ~n7527;
  assign n7529 = ~n7356 & n7528;
  assign n7530 = pi1091 & n7410;
  assign n7531 = n7383 & n7530;
  assign n7532 = n7414 & n7531;
  assign n7533 = pi1093 & n7532;
  assign n7534 = n7408 & n7533;
  assign n7535 = pi75 & ~n7534;
  assign n7536 = n2531 & n7440;
  assign n7537 = n7443 & n7536;
  assign n7538 = pi100 & ~n7537;
  assign n7539 = ~n7480 & ~n7482;
  assign n7540 = ~pi39 & ~n7539;
  assign n7541 = pi1093 & n2922;
  assign n7542 = n7491 & n7541;
  assign n7543 = ~n6223 & n7542;
  assign n7544 = ~pi216 & n6590;
  assign n7545 = n7543 & n7544;
  assign n7546 = ~n6207 & n7542;
  assign n7547 = ~pi299 & n6359;
  assign n7548 = ~pi224 & n7547;
  assign n7549 = n7546 & n7548;
  assign n7550 = pi39 & ~n7545;
  assign n7551 = ~n7549 & n7550;
  assign n7552 = ~pi38 & ~n7551;
  assign n7553 = ~n7540 & n7552;
  assign n7554 = ~pi100 & ~n7553;
  assign n7555 = pi1093 & n7455;
  assign n7556 = n7552 & n7555;
  assign n7557 = ~n7479 & n7556;
  assign n7558 = n7554 & ~n7557;
  assign n7559 = ~n7538 & ~n7558;
  assign n7560 = ~pi87 & ~n7559;
  assign n7561 = ~pi1091 & pi1093;
  assign n7562 = ~n7430 & n7561;
  assign n7563 = ~n7427 & ~n7561;
  assign n7564 = n2628 & ~n7563;
  assign n7565 = ~n7562 & n7564;
  assign n7566 = pi87 & ~n7565;
  assign n7567 = ~n7560 & ~n7566;
  assign n7568 = ~pi75 & ~n7567;
  assign n7569 = ~n7535 & ~n7568;
  assign n7570 = pi567 & ~n7569;
  assign n7571 = n7405 & ~n7570;
  assign n7572 = n7356 & ~n7571;
  assign n7573 = ~po1038 & ~n7529;
  assign n7574 = ~n7572 & n7573;
  assign n7575 = pi217 & ~n7359;
  assign n7576 = ~n7574 & n7575;
  assign n7577 = ~pi1161 & ~pi1162;
  assign n7578 = ~pi1163 & n7577;
  assign n7579 = ~pi590 & ~pi591;
  assign n7580 = ~pi592 & n7579;
  assign n7581 = pi437 & ~pi453;
  assign n7582 = ~pi437 & pi453;
  assign n7583 = ~n7581 & ~n7582;
  assign n7584 = pi417 & ~pi418;
  assign n7585 = ~pi417 & pi418;
  assign n7586 = ~n7584 & ~n7585;
  assign n7587 = pi464 & ~n7586;
  assign n7588 = ~pi464 & n7586;
  assign n7589 = ~n7587 & ~n7588;
  assign n7590 = n7583 & n7589;
  assign n7591 = ~n7583 & ~n7589;
  assign n7592 = ~n7590 & ~n7591;
  assign n7593 = ~pi415 & ~pi431;
  assign n7594 = pi415 & pi431;
  assign n7595 = ~n7593 & ~n7594;
  assign n7596 = pi416 & ~pi438;
  assign n7597 = ~pi416 & pi438;
  assign n7598 = ~n7596 & ~n7597;
  assign n7599 = n7595 & n7598;
  assign n7600 = ~n7595 & ~n7598;
  assign n7601 = ~n7599 & ~n7600;
  assign n7602 = n7592 & n7601;
  assign n7603 = ~n7592 & ~n7601;
  assign n7604 = pi1197 & ~n7602;
  assign n7605 = ~n7603 & n7604;
  assign n7606 = ~pi421 & ~pi454;
  assign n7607 = pi421 & pi454;
  assign n7608 = ~n7606 & ~n7607;
  assign n7609 = pi419 & ~pi420;
  assign n7610 = ~pi419 & pi420;
  assign n7611 = ~n7609 & ~n7610;
  assign n7612 = n7608 & ~n7611;
  assign n7613 = ~n7608 & n7611;
  assign n7614 = ~n7612 & ~n7613;
  assign n7615 = ~pi423 & ~pi424;
  assign n7616 = pi423 & pi424;
  assign n7617 = ~n7615 & ~n7616;
  assign n7618 = pi432 & ~pi459;
  assign n7619 = ~pi432 & pi459;
  assign n7620 = ~n7618 & ~n7619;
  assign n7621 = n7617 & ~n7620;
  assign n7622 = ~n7617 & n7620;
  assign n7623 = ~n7621 & ~n7622;
  assign n7624 = n7614 & n7623;
  assign n7625 = ~n7614 & ~n7623;
  assign n7626 = ~n7624 & ~n7625;
  assign n7627 = pi425 & n7626;
  assign n7628 = ~pi425 & ~n7626;
  assign n7629 = pi1198 & ~n7627;
  assign n7630 = ~n7628 & n7629;
  assign n7631 = ~n7605 & ~n7630;
  assign n7632 = ~pi436 & ~pi443;
  assign n7633 = pi436 & pi443;
  assign n7634 = ~n7632 & ~n7633;
  assign n7635 = ~pi444 & ~n7634;
  assign n7636 = pi444 & n7634;
  assign n7637 = ~n7635 & ~n7636;
  assign n7638 = ~pi429 & ~pi435;
  assign n7639 = pi429 & pi435;
  assign n7640 = ~n7638 & ~n7639;
  assign n7641 = ~pi434 & ~pi446;
  assign n7642 = pi434 & pi446;
  assign n7643 = ~n7641 & ~n7642;
  assign n7644 = pi414 & n7643;
  assign n7645 = ~pi414 & ~n7643;
  assign n7646 = ~n7644 & ~n7645;
  assign n7647 = pi422 & ~n7646;
  assign n7648 = ~pi422 & n7646;
  assign n7649 = ~n7647 & ~n7648;
  assign n7650 = n7640 & n7649;
  assign n7651 = ~n7640 & ~n7649;
  assign n7652 = ~n7650 & ~n7651;
  assign n7653 = ~n7637 & n7652;
  assign n7654 = ~pi592 & pi1196;
  assign n7655 = n7637 & ~n7652;
  assign n7656 = ~n7653 & n7654;
  assign n7657 = ~n7655 & n7656;
  assign n7658 = n7631 & ~n7657;
  assign n7659 = ~pi433 & ~pi451;
  assign n7660 = pi433 & pi451;
  assign n7661 = ~n7659 & ~n7660;
  assign n7662 = pi448 & ~pi449;
  assign n7663 = ~pi448 & pi449;
  assign n7664 = ~n7662 & ~n7663;
  assign n7665 = n7661 & n7664;
  assign n7666 = ~n7661 & ~n7664;
  assign n7667 = ~n7665 & ~n7666;
  assign n7668 = pi427 & ~pi428;
  assign n7669 = ~pi427 & pi428;
  assign n7670 = ~n7668 & ~n7669;
  assign n7671 = ~pi426 & ~pi430;
  assign n7672 = pi426 & pi430;
  assign n7673 = ~n7671 & ~n7672;
  assign n7674 = pi445 & ~n7673;
  assign n7675 = ~pi445 & n7673;
  assign n7676 = ~n7674 & ~n7675;
  assign n7677 = ~n7670 & n7676;
  assign n7678 = n7670 & ~n7676;
  assign n7679 = ~n7677 & ~n7678;
  assign n7680 = ~n7667 & ~n7679;
  assign n7681 = n7667 & n7679;
  assign n7682 = pi1199 & ~n7680;
  assign n7683 = ~n7681 & n7682;
  assign n7684 = n7658 & ~n7683;
  assign n7685 = n7580 & ~n7684;
  assign n7686 = n7353 & ~n7685;
  assign n7687 = pi588 & ~n7686;
  assign n7688 = ~pi592 & n7353;
  assign n7689 = ~pi379 & ~pi382;
  assign n7690 = pi379 & pi382;
  assign n7691 = ~n7689 & ~n7690;
  assign n7692 = ~pi376 & ~pi439;
  assign n7693 = pi376 & pi439;
  assign n7694 = ~n7692 & ~n7693;
  assign n7695 = pi378 & ~pi381;
  assign n7696 = ~pi378 & pi381;
  assign n7697 = ~n7695 & ~n7696;
  assign n7698 = n7694 & n7697;
  assign n7699 = ~n7694 & ~n7697;
  assign n7700 = ~n7698 & ~n7699;
  assign n7701 = n7691 & ~n7700;
  assign n7702 = ~n7691 & n7700;
  assign n7703 = ~n7701 & ~n7702;
  assign n7704 = pi317 & ~pi385;
  assign n7705 = ~pi317 & pi385;
  assign n7706 = ~n7704 & ~n7705;
  assign n7707 = pi377 & ~n7706;
  assign n7708 = ~pi377 & n7706;
  assign n7709 = ~n7707 & ~n7708;
  assign n7710 = n7703 & n7709;
  assign n7711 = ~n7703 & ~n7709;
  assign n7712 = ~n7710 & ~n7711;
  assign n7713 = pi1199 & n7712;
  assign n7714 = ~pi380 & ~pi387;
  assign n7715 = pi380 & pi387;
  assign n7716 = ~n7714 & ~n7715;
  assign n7717 = pi337 & ~pi339;
  assign n7718 = ~pi337 & pi339;
  assign n7719 = ~n7717 & ~n7718;
  assign n7720 = pi363 & ~pi372;
  assign n7721 = ~pi363 & pi372;
  assign n7722 = ~n7720 & ~n7721;
  assign n7723 = pi386 & n7722;
  assign n7724 = ~pi386 & ~n7722;
  assign n7725 = ~n7723 & ~n7724;
  assign n7726 = ~pi338 & ~pi388;
  assign n7727 = pi338 & pi388;
  assign n7728 = ~n7726 & ~n7727;
  assign n7729 = n7725 & ~n7728;
  assign n7730 = ~n7725 & n7728;
  assign n7731 = ~n7729 & ~n7730;
  assign n7732 = n7719 & n7731;
  assign n7733 = ~n7719 & ~n7731;
  assign n7734 = ~n7732 & ~n7733;
  assign n7735 = n7716 & ~n7734;
  assign n7736 = ~n7716 & n7734;
  assign n7737 = pi1196 & ~n7735;
  assign n7738 = ~n7736 & n7737;
  assign n7739 = ~pi336 & ~pi383;
  assign n7740 = pi336 & pi383;
  assign n7741 = ~n7739 & ~n7740;
  assign n7742 = pi364 & n7741;
  assign n7743 = ~pi364 & ~n7741;
  assign n7744 = ~n7742 & ~n7743;
  assign n7745 = pi366 & ~n7744;
  assign n7746 = ~pi366 & n7744;
  assign n7747 = ~n7745 & ~n7746;
  assign n7748 = ~pi365 & ~pi447;
  assign n7749 = pi365 & pi447;
  assign n7750 = ~n7748 & ~n7749;
  assign n7751 = pi368 & ~pi389;
  assign n7752 = ~pi368 & pi389;
  assign n7753 = ~n7751 & ~n7752;
  assign n7754 = n7750 & ~n7753;
  assign n7755 = ~n7750 & n7753;
  assign n7756 = ~n7754 & ~n7755;
  assign n7757 = n7747 & n7756;
  assign n7758 = ~n7747 & ~n7756;
  assign n7759 = ~n7757 & ~n7758;
  assign n7760 = pi367 & ~n7759;
  assign n7761 = ~pi367 & n7759;
  assign n7762 = pi1197 & ~n7760;
  assign n7763 = ~n7761 & n7762;
  assign n7764 = ~n7738 & ~n7763;
  assign n7765 = ~n7713 & n7764;
  assign n7766 = pi592 & n7353;
  assign n7767 = ~pi370 & ~pi371;
  assign n7768 = pi370 & pi371;
  assign n7769 = ~n7767 & ~n7768;
  assign n7770 = ~pi384 & ~pi442;
  assign n7771 = pi384 & pi442;
  assign n7772 = ~n7770 & ~n7771;
  assign n7773 = pi440 & n7772;
  assign n7774 = ~pi440 & ~n7772;
  assign n7775 = ~n7773 & ~n7774;
  assign n7776 = pi373 & ~pi375;
  assign n7777 = ~pi373 & pi375;
  assign n7778 = ~n7776 & ~n7777;
  assign n7779 = n7775 & n7778;
  assign n7780 = ~n7775 & ~n7778;
  assign n7781 = ~n7779 & ~n7780;
  assign n7782 = n7769 & n7781;
  assign n7783 = ~n7769 & ~n7781;
  assign n7784 = ~n7782 & ~n7783;
  assign n7785 = ~pi369 & n7784;
  assign n7786 = pi369 & ~n7784;
  assign n7787 = ~n7785 & ~n7786;
  assign n7788 = pi374 & n7787;
  assign n7789 = ~pi374 & ~n7787;
  assign n7790 = pi1198 & ~n7788;
  assign n7791 = ~n7789 & n7790;
  assign n7792 = n7765 & n7766;
  assign n7793 = ~n7791 & n7792;
  assign n7794 = ~pi590 & ~n7688;
  assign n7795 = ~n7793 & n7794;
  assign n7796 = pi1199 & ~n7766;
  assign n7797 = pi351 & n7796;
  assign n7798 = pi351 & pi1199;
  assign n7799 = ~pi452 & ~pi455;
  assign n7800 = pi452 & pi455;
  assign n7801 = ~n7799 & ~n7800;
  assign n7802 = ~pi361 & ~pi458;
  assign n7803 = pi361 & pi458;
  assign n7804 = ~n7802 & ~n7803;
  assign n7805 = ~pi342 & ~pi441;
  assign n7806 = pi342 & pi441;
  assign n7807 = ~n7805 & ~n7806;
  assign n7808 = n7804 & ~n7807;
  assign n7809 = ~n7804 & n7807;
  assign n7810 = ~n7808 & ~n7809;
  assign n7811 = pi320 & ~pi460;
  assign n7812 = ~pi320 & pi460;
  assign n7813 = ~n7811 & ~n7812;
  assign n7814 = pi355 & ~n7813;
  assign n7815 = ~pi355 & n7813;
  assign n7816 = ~n7814 & ~n7815;
  assign n7817 = n7810 & n7816;
  assign n7818 = ~n7810 & ~n7816;
  assign n7819 = ~n7817 & ~n7818;
  assign n7820 = n7801 & n7819;
  assign n7821 = ~n7801 & ~n7819;
  assign n7822 = ~n7820 & ~n7821;
  assign n7823 = ~pi592 & ~pi1198;
  assign n7824 = ~n7822 & n7823;
  assign n7825 = n7353 & ~n7824;
  assign n7826 = pi1196 & ~n7825;
  assign n7827 = pi315 & ~pi359;
  assign n7828 = ~pi315 & pi359;
  assign n7829 = ~n7827 & ~n7828;
  assign n7830 = ~pi321 & ~pi347;
  assign n7831 = pi321 & pi347;
  assign n7832 = ~n7830 & ~n7831;
  assign n7833 = ~pi316 & ~pi349;
  assign n7834 = pi316 & pi349;
  assign n7835 = ~n7833 & ~n7834;
  assign n7836 = pi322 & ~pi348;
  assign n7837 = ~pi322 & pi348;
  assign n7838 = ~n7836 & ~n7837;
  assign n7839 = n7835 & n7838;
  assign n7840 = ~n7835 & ~n7838;
  assign n7841 = ~n7839 & ~n7840;
  assign n7842 = n7832 & ~n7841;
  assign n7843 = ~n7832 & n7841;
  assign n7844 = ~n7842 & ~n7843;
  assign n7845 = n7829 & n7844;
  assign n7846 = ~n7829 & ~n7844;
  assign n7847 = ~n7845 & ~n7846;
  assign n7848 = ~pi350 & ~n7847;
  assign n7849 = pi1196 & ~n7822;
  assign n7850 = pi350 & n7847;
  assign n7851 = ~n7848 & ~n7849;
  assign n7852 = ~n7850 & n7851;
  assign n7853 = n7688 & n7852;
  assign n7854 = pi1198 & ~n7853;
  assign n7855 = ~pi345 & ~pi346;
  assign n7856 = pi345 & pi346;
  assign n7857 = ~n7855 & ~n7856;
  assign n7858 = pi323 & n7857;
  assign n7859 = ~pi323 & ~n7857;
  assign n7860 = ~n7858 & ~n7859;
  assign n7861 = pi358 & ~pi450;
  assign n7862 = ~pi358 & pi450;
  assign n7863 = ~n7861 & ~n7862;
  assign n7864 = n7860 & n7863;
  assign n7865 = ~n7860 & ~n7863;
  assign n7866 = ~n7864 & ~n7865;
  assign n7867 = pi327 & ~pi362;
  assign n7868 = ~pi327 & pi362;
  assign n7869 = ~n7867 & ~n7868;
  assign n7870 = pi343 & ~pi344;
  assign n7871 = ~pi343 & pi344;
  assign n7872 = ~n7870 & ~n7871;
  assign n7873 = n7869 & n7872;
  assign n7874 = ~n7869 & ~n7872;
  assign n7875 = ~n7873 & ~n7874;
  assign n7876 = ~n7866 & n7875;
  assign n7877 = n7866 & ~n7875;
  assign n7878 = pi1197 & ~n7876;
  assign n7879 = ~n7877 & n7878;
  assign n7880 = ~n7826 & ~n7879;
  assign n7881 = ~n7854 & n7880;
  assign n7882 = ~pi592 & ~n7881;
  assign n7883 = n7353 & ~n7882;
  assign n7884 = ~n7798 & ~n7883;
  assign n7885 = ~pi356 & ~pi357;
  assign n7886 = pi356 & pi357;
  assign n7887 = ~n7885 & ~n7886;
  assign n7888 = pi352 & ~pi353;
  assign n7889 = ~pi352 & pi353;
  assign n7890 = ~n7888 & ~n7889;
  assign n7891 = ~pi360 & ~pi462;
  assign n7892 = pi360 & pi462;
  assign n7893 = ~n7891 & ~n7892;
  assign n7894 = pi354 & ~n7893;
  assign n7895 = ~pi354 & n7893;
  assign n7896 = ~n7894 & ~n7895;
  assign n7897 = n7890 & n7896;
  assign n7898 = ~n7890 & ~n7896;
  assign n7899 = ~n7897 & ~n7898;
  assign n7900 = ~n7887 & ~n7899;
  assign n7901 = n7887 & n7899;
  assign n7902 = ~n7900 & ~n7901;
  assign n7903 = pi461 & ~n7902;
  assign n7904 = ~pi461 & n7902;
  assign n7905 = ~n7903 & ~n7904;
  assign n7906 = ~n7797 & n7905;
  assign n7907 = ~n7884 & n7906;
  assign n7908 = ~pi351 & n7796;
  assign n7909 = ~pi351 & pi1199;
  assign n7910 = ~n7883 & ~n7909;
  assign n7911 = ~n7905 & ~n7908;
  assign n7912 = ~n7910 & n7911;
  assign n7913 = pi590 & ~n7907;
  assign n7914 = ~n7912 & n7913;
  assign n7915 = ~pi591 & ~n7795;
  assign n7916 = ~n7914 & n7915;
  assign n7917 = pi590 & n7353;
  assign n7918 = pi318 & ~pi409;
  assign n7919 = ~pi318 & pi409;
  assign n7920 = ~n7918 & ~n7919;
  assign n7921 = pi403 & ~pi405;
  assign n7922 = ~pi403 & pi405;
  assign n7923 = ~n7921 & ~n7922;
  assign n7924 = pi325 & n7923;
  assign n7925 = ~pi325 & ~n7923;
  assign n7926 = ~n7924 & ~n7925;
  assign n7927 = ~pi401 & ~pi402;
  assign n7928 = pi401 & pi402;
  assign n7929 = ~n7927 & ~n7928;
  assign n7930 = pi326 & ~pi406;
  assign n7931 = ~pi326 & pi406;
  assign n7932 = ~n7930 & ~n7931;
  assign n7933 = n7929 & n7932;
  assign n7934 = ~n7929 & ~n7932;
  assign n7935 = ~n7933 & ~n7934;
  assign n7936 = n7926 & ~n7935;
  assign n7937 = ~n7926 & n7935;
  assign n7938 = ~n7936 & ~n7937;
  assign n7939 = n7920 & n7938;
  assign n7940 = ~n7920 & ~n7938;
  assign n7941 = ~n7939 & ~n7940;
  assign n7942 = n7444 & ~n7941;
  assign n7943 = pi567 & n7942;
  assign n7944 = ~pi390 & ~pi410;
  assign n7945 = pi390 & pi410;
  assign n7946 = ~n7944 & ~n7945;
  assign n7947 = pi411 & ~n7946;
  assign n7948 = ~pi411 & n7946;
  assign n7949 = ~n7947 & ~n7948;
  assign n7950 = ~pi397 & ~pi404;
  assign n7951 = pi397 & pi404;
  assign n7952 = ~n7950 & ~n7951;
  assign n7953 = pi412 & ~n7952;
  assign n7954 = ~pi412 & n7952;
  assign n7955 = ~n7953 & ~n7954;
  assign n7956 = ~pi319 & ~pi324;
  assign n7957 = pi319 & pi324;
  assign n7958 = ~n7956 & ~n7957;
  assign n7959 = pi456 & n7958;
  assign n7960 = ~pi456 & ~n7958;
  assign n7961 = ~n7959 & ~n7960;
  assign n7962 = n7955 & ~n7961;
  assign n7963 = ~n7955 & n7961;
  assign n7964 = ~n7962 & ~n7963;
  assign n7965 = n7949 & n7964;
  assign n7966 = ~n7949 & ~n7964;
  assign n7967 = ~n7965 & ~n7966;
  assign n7968 = pi1196 & ~n7967;
  assign n7969 = ~pi592 & ~n7968;
  assign n7970 = n7943 & n7969;
  assign n7971 = n7796 & ~n7970;
  assign n7972 = n7353 & ~n7654;
  assign n7973 = n7444 & n7967;
  assign n7974 = pi567 & n7973;
  assign n7975 = n7654 & n7974;
  assign n7976 = ~pi1199 & ~n7972;
  assign n7977 = ~n7975 & n7976;
  assign n7978 = ~n7971 & ~n7977;
  assign n7979 = pi1198 & ~n7766;
  assign n7980 = n7978 & ~n7979;
  assign n7981 = ~pi328 & ~pi408;
  assign n7982 = pi328 & pi408;
  assign n7983 = ~n7981 & ~n7982;
  assign n7984 = ~pi329 & ~pi395;
  assign n7985 = pi329 & pi395;
  assign n7986 = ~n7984 & ~n7985;
  assign n7987 = n7983 & ~n7986;
  assign n7988 = ~n7983 & n7986;
  assign n7989 = ~n7987 & ~n7988;
  assign n7990 = ~pi398 & ~pi399;
  assign n7991 = pi398 & pi399;
  assign n7992 = ~n7990 & ~n7991;
  assign n7993 = pi400 & n7992;
  assign n7994 = ~pi400 & ~n7992;
  assign n7995 = ~n7993 & ~n7994;
  assign n7996 = pi394 & ~pi396;
  assign n7997 = ~pi394 & pi396;
  assign n7998 = ~n7996 & ~n7997;
  assign n7999 = n7995 & ~n7998;
  assign n8000 = ~n7995 & n7998;
  assign n8001 = ~n7999 & ~n8000;
  assign n8002 = n7989 & n8001;
  assign n8003 = ~n7989 & ~n8001;
  assign n8004 = ~n8002 & ~n8003;
  assign n8005 = ~n7980 & ~n8004;
  assign n8006 = ~pi407 & ~pi463;
  assign n8007 = pi407 & pi463;
  assign n8008 = ~n8006 & ~n8007;
  assign n8009 = pi335 & ~pi413;
  assign n8010 = ~pi335 & pi413;
  assign n8011 = ~n8009 & ~n8010;
  assign n8012 = n8008 & n8011;
  assign n8013 = ~n8008 & ~n8011;
  assign n8014 = ~n8012 & ~n8013;
  assign n8015 = pi334 & n8014;
  assign n8016 = ~pi334 & ~n8014;
  assign n8017 = ~n8015 & ~n8016;
  assign n8018 = ~pi393 & ~n8017;
  assign n8019 = pi393 & n8017;
  assign n8020 = ~n8018 & ~n8019;
  assign n8021 = pi392 & ~n8020;
  assign n8022 = ~pi392 & n8020;
  assign n8023 = ~n8021 & ~n8022;
  assign n8024 = pi391 & n8023;
  assign n8025 = ~pi391 & ~n8023;
  assign n8026 = ~n8024 & ~n8025;
  assign n8027 = ~pi333 & pi1197;
  assign n8028 = ~n7766 & n8027;
  assign n8029 = n7978 & ~n8028;
  assign n8030 = n8026 & ~n8029;
  assign n8031 = pi333 & pi1197;
  assign n8032 = ~n7766 & n8031;
  assign n8033 = ~n8026 & n8032;
  assign n8034 = ~n7978 & ~n8031;
  assign n8035 = ~pi590 & ~n8033;
  assign n8036 = ~n8034 & n8035;
  assign n8037 = ~n8005 & n8036;
  assign n8038 = ~n8030 & n8037;
  assign n8039 = ~n7917 & ~n8038;
  assign n8040 = pi591 & ~n8039;
  assign n8041 = ~pi588 & ~n8040;
  assign n8042 = ~n7916 & n8041;
  assign n8043 = n7358 & ~n7687;
  assign n8044 = ~n8042 & n8043;
  assign n8045 = ~pi1196 & n7528;
  assign n8046 = ~pi443 & ~pi592;
  assign n8047 = ~pi87 & ~n7538;
  assign n8048 = ~n7554 & n8047;
  assign n8049 = pi87 & n2628;
  assign n8050 = ~n7428 & n8049;
  assign n8051 = ~n7429 & n8050;
  assign n8052 = ~pi75 & ~n8051;
  assign n8053 = ~n8048 & n8052;
  assign n8054 = ~n7535 & ~n8053;
  assign n8055 = pi567 & ~n8054;
  assign n8056 = n7405 & ~n8055;
  assign n8057 = n8046 & ~n8056;
  assign n8058 = n7528 & ~n8046;
  assign n8059 = ~pi436 & ~pi444;
  assign n8060 = pi436 & pi444;
  assign n8061 = ~n8059 & ~n8060;
  assign n8062 = ~n7652 & ~n8061;
  assign n8063 = n7652 & n8061;
  assign n8064 = ~n8062 & ~n8063;
  assign n8065 = ~n8057 & ~n8064;
  assign n8066 = ~n8058 & n8065;
  assign n8067 = pi443 & ~pi592;
  assign n8068 = n7528 & ~n8067;
  assign n8069 = ~n8056 & n8067;
  assign n8070 = n8064 & ~n8069;
  assign n8071 = ~n8068 & n8070;
  assign n8072 = pi1196 & ~n8066;
  assign n8073 = ~n8071 & n8072;
  assign n8074 = ~n8045 & ~n8073;
  assign n8075 = n7631 & ~n8074;
  assign n8076 = ~pi592 & ~n8056;
  assign n8077 = pi592 & n7528;
  assign n8078 = ~n8076 & ~n8077;
  assign n8079 = ~n7631 & ~n8078;
  assign n8080 = ~n8075 & ~n8079;
  assign n8081 = ~pi1199 & ~n8080;
  assign n8082 = ~pi428 & n8080;
  assign n8083 = pi428 & n8078;
  assign n8084 = ~pi427 & ~n8083;
  assign n8085 = ~n8082 & n8084;
  assign n8086 = ~pi428 & n8078;
  assign n8087 = pi428 & n8080;
  assign n8088 = pi427 & ~n8086;
  assign n8089 = ~n8087 & n8088;
  assign n8090 = ~n8085 & ~n8089;
  assign n8091 = pi445 & n7667;
  assign n8092 = ~pi445 & ~n7667;
  assign n8093 = ~n8091 & ~n8092;
  assign n8094 = ~n8090 & n8093;
  assign n8095 = ~n7670 & n8080;
  assign n8096 = n7670 & n8078;
  assign n8097 = ~n8093 & ~n8096;
  assign n8098 = ~n8095 & n8097;
  assign n8099 = ~n7673 & ~n8098;
  assign n8100 = ~n8094 & n8099;
  assign n8101 = ~n8090 & ~n8093;
  assign n8102 = n8093 & ~n8096;
  assign n8103 = ~n8095 & n8102;
  assign n8104 = n7673 & ~n8103;
  assign n8105 = ~n8101 & n8104;
  assign n8106 = pi1199 & ~n8100;
  assign n8107 = ~n8105 & n8106;
  assign n8108 = n7579 & ~n8081;
  assign n8109 = ~n8107 & n8108;
  assign n8110 = ~n7528 & ~n7579;
  assign n8111 = ~n7356 & ~n8110;
  assign n8112 = ~n8109 & n8111;
  assign n8113 = n7571 & ~n7579;
  assign n8114 = pi592 & ~n7571;
  assign n8115 = ~n8076 & ~n8114;
  assign n8116 = ~n7631 & n8115;
  assign n8117 = ~pi1196 & ~n7571;
  assign n8118 = pi443 & ~n7571;
  assign n8119 = ~n8057 & ~n8118;
  assign n8120 = ~n8064 & ~n8119;
  assign n8121 = ~pi443 & ~n7571;
  assign n8122 = ~n8069 & ~n8121;
  assign n8123 = n8064 & ~n8122;
  assign n8124 = ~n8114 & ~n8120;
  assign n8125 = ~n8123 & n8124;
  assign n8126 = pi1196 & ~n8125;
  assign n8127 = n7631 & ~n8117;
  assign n8128 = ~n8126 & n8127;
  assign n8129 = ~n8116 & ~n8128;
  assign n8130 = ~pi1199 & n8129;
  assign n8131 = pi428 & ~n8129;
  assign n8132 = ~pi428 & n8115;
  assign n8133 = ~n8131 & ~n8132;
  assign n8134 = ~pi427 & ~n8133;
  assign n8135 = pi428 & ~n8115;
  assign n8136 = ~pi428 & n8129;
  assign n8137 = ~n8135 & ~n8136;
  assign n8138 = pi427 & n8137;
  assign n8139 = ~n8134 & ~n8138;
  assign n8140 = pi430 & ~n8139;
  assign n8141 = pi427 & ~n8133;
  assign n8142 = ~pi427 & n8137;
  assign n8143 = ~n8141 & ~n8142;
  assign n8144 = ~pi430 & ~n8143;
  assign n8145 = ~n8140 & ~n8144;
  assign n8146 = ~pi426 & n8145;
  assign n8147 = pi430 & ~n8143;
  assign n8148 = ~pi430 & ~n8139;
  assign n8149 = ~n8147 & ~n8148;
  assign n8150 = pi426 & n8149;
  assign n8151 = n8093 & ~n8146;
  assign n8152 = ~n8150 & n8151;
  assign n8153 = ~pi426 & n8149;
  assign n8154 = pi426 & n8145;
  assign n8155 = ~n8093 & ~n8153;
  assign n8156 = ~n8154 & n8155;
  assign n8157 = pi1199 & ~n8152;
  assign n8158 = ~n8156 & n8157;
  assign n8159 = n7579 & ~n8130;
  assign n8160 = ~n8158 & n8159;
  assign n8161 = n7356 & ~n8113;
  assign n8162 = ~n8160 & n8161;
  assign n8163 = ~n8112 & ~n8162;
  assign n8164 = pi588 & ~n8163;
  assign n8165 = pi591 & n7571;
  assign n8166 = n7849 & ~n8115;
  assign n8167 = pi350 & ~pi592;
  assign n8168 = ~n7571 & ~n8167;
  assign n8169 = ~n8056 & n8167;
  assign n8170 = n7847 & ~n8169;
  assign n8171 = ~n8168 & n8170;
  assign n8172 = ~pi350 & ~pi592;
  assign n8173 = ~n7571 & ~n8172;
  assign n8174 = ~n8056 & n8172;
  assign n8175 = ~n7847 & ~n8174;
  assign n8176 = ~n8173 & n8175;
  assign n8177 = ~n7849 & ~n8171;
  assign n8178 = ~n8176 & n8177;
  assign n8179 = pi1198 & ~n8166;
  assign n8180 = ~n8178 & n8179;
  assign n8181 = ~pi455 & n8115;
  assign n8182 = pi455 & n7571;
  assign n8183 = ~pi452 & ~n8182;
  assign n8184 = ~n8181 & n8183;
  assign n8185 = ~pi455 & n7571;
  assign n8186 = pi455 & n8115;
  assign n8187 = pi452 & ~n8185;
  assign n8188 = ~n8186 & n8187;
  assign n8189 = ~n8184 & ~n8188;
  assign n8190 = ~n7819 & ~n8189;
  assign n8191 = n7801 & n8115;
  assign n8192 = n7571 & ~n7801;
  assign n8193 = n7819 & ~n8192;
  assign n8194 = ~n8191 & n8193;
  assign n8195 = ~n8190 & ~n8194;
  assign n8196 = pi1196 & ~n8195;
  assign n8197 = ~pi1198 & ~n8117;
  assign n8198 = ~n8196 & n8197;
  assign n8199 = ~n8180 & ~n8198;
  assign n8200 = ~n7879 & ~n8199;
  assign n8201 = n7879 & n8115;
  assign n8202 = ~n8200 & ~n8201;
  assign n8203 = ~n7798 & n8202;
  assign n8204 = pi1199 & ~n8115;
  assign n8205 = pi351 & n8204;
  assign n8206 = ~n8203 & ~n8205;
  assign n8207 = ~pi461 & ~n8206;
  assign n8208 = ~n7909 & n8202;
  assign n8209 = ~pi351 & n8204;
  assign n8210 = ~n8208 & ~n8209;
  assign n8211 = pi461 & ~n8210;
  assign n8212 = ~n8207 & ~n8211;
  assign n8213 = ~n7887 & n8212;
  assign n8214 = ~pi461 & ~n8210;
  assign n8215 = pi461 & ~n8206;
  assign n8216 = ~n8214 & ~n8215;
  assign n8217 = n7887 & n8216;
  assign n8218 = ~n7899 & ~n8213;
  assign n8219 = ~n8217 & n8218;
  assign n8220 = pi356 & ~pi357;
  assign n8221 = ~pi356 & pi357;
  assign n8222 = ~n8220 & ~n8221;
  assign n8223 = n8212 & ~n8222;
  assign n8224 = n8216 & n8222;
  assign n8225 = n7899 & ~n8223;
  assign n8226 = ~n8224 & n8225;
  assign n8227 = ~pi591 & ~n8219;
  assign n8228 = ~n8226 & n8227;
  assign n8229 = pi590 & ~n8165;
  assign n8230 = ~n8228 & n8229;
  assign n8231 = pi1198 & ~n8004;
  assign n8232 = ~pi1196 & ~n7568;
  assign n8233 = n7430 & n7967;
  assign n8234 = n7561 & ~n8233;
  assign n8235 = pi87 & n7564;
  assign n8236 = ~n8234 & n8235;
  assign n8237 = n7557 & n7967;
  assign n8238 = n7554 & ~n8237;
  assign n8239 = n8047 & ~n8238;
  assign n8240 = ~pi75 & ~pi592;
  assign n8241 = ~n8236 & n8240;
  assign n8242 = ~n8239 & n8241;
  assign n8243 = pi1196 & ~n8242;
  assign n8244 = ~pi1199 & ~n8243;
  assign n8245 = ~n8232 & n8244;
  assign n8246 = ~n7569 & ~n8240;
  assign n8247 = ~pi75 & n7968;
  assign n8248 = ~n7941 & ~n8247;
  assign n8249 = n7557 & n8248;
  assign n8250 = n7554 & ~n8249;
  assign n8251 = n8047 & ~n8250;
  assign n8252 = ~n7941 & ~n7968;
  assign n8253 = n7430 & n8252;
  assign n8254 = n7561 & ~n8253;
  assign n8255 = n8235 & ~n8254;
  assign n8256 = pi1199 & n8240;
  assign n8257 = ~n8255 & n8256;
  assign n8258 = ~n8251 & n8257;
  assign n8259 = ~n8245 & ~n8258;
  assign n8260 = ~n8246 & n8259;
  assign n8261 = pi567 & ~n8260;
  assign n8262 = n7405 & ~n8231;
  assign n8263 = ~n8261 & n8262;
  assign n8264 = n8115 & n8231;
  assign n8265 = ~n8263 & ~n8264;
  assign n8266 = pi333 & ~n8265;
  assign n8267 = ~pi1197 & ~n8265;
  assign n8268 = pi1197 & n8115;
  assign n8269 = ~n8267 & ~n8268;
  assign n8270 = ~pi333 & ~n8269;
  assign n8271 = ~n8266 & ~n8270;
  assign n8272 = ~pi391 & ~n8271;
  assign n8273 = ~n8031 & ~n8265;
  assign n8274 = pi333 & n8268;
  assign n8275 = ~n8273 & ~n8274;
  assign n8276 = pi391 & ~n8275;
  assign n8277 = ~n8272 & ~n8276;
  assign n8278 = pi392 & ~n8277;
  assign n8279 = pi391 & ~n8271;
  assign n8280 = ~pi391 & ~n8275;
  assign n8281 = ~n8279 & ~n8280;
  assign n8282 = ~pi392 & ~n8281;
  assign n8283 = ~n8278 & ~n8282;
  assign n8284 = pi393 & ~n8283;
  assign n8285 = pi392 & ~n8281;
  assign n8286 = ~pi392 & ~n8277;
  assign n8287 = ~n8285 & ~n8286;
  assign n8288 = ~pi393 & ~n8287;
  assign n8289 = ~n8284 & ~n8288;
  assign n8290 = ~pi334 & ~n8289;
  assign n8291 = pi393 & ~n8287;
  assign n8292 = ~pi393 & ~n8283;
  assign n8293 = ~n8291 & ~n8292;
  assign n8294 = pi334 & ~n8293;
  assign n8295 = ~n8014 & ~n8290;
  assign n8296 = ~n8294 & n8295;
  assign n8297 = ~pi334 & ~n8293;
  assign n8298 = pi334 & ~n8289;
  assign n8299 = n8014 & ~n8297;
  assign n8300 = ~n8298 & n8299;
  assign n8301 = pi591 & ~n8296;
  assign n8302 = ~n8300 & n8301;
  assign n8303 = pi592 & ~n7765;
  assign n8304 = n7571 & ~n8303;
  assign n8305 = n8056 & n8303;
  assign n8306 = ~n8304 & ~n8305;
  assign n8307 = pi374 & ~n8306;
  assign n8308 = ~pi1198 & n8306;
  assign n8309 = pi592 & ~n8056;
  assign n8310 = ~pi592 & ~n7571;
  assign n8311 = ~n8309 & ~n8310;
  assign n8312 = pi1198 & ~n8311;
  assign n8313 = ~n8308 & ~n8312;
  assign n8314 = ~pi374 & n8313;
  assign n8315 = ~n8307 & ~n8314;
  assign n8316 = pi369 & ~n8315;
  assign n8317 = ~pi374 & n8306;
  assign n8318 = pi374 & ~n8313;
  assign n8319 = ~n8317 & ~n8318;
  assign n8320 = ~pi369 & n8319;
  assign n8321 = ~n8316 & ~n8320;
  assign n8322 = pi370 & ~n8321;
  assign n8323 = ~pi369 & ~n8315;
  assign n8324 = pi369 & n8319;
  assign n8325 = ~n8323 & ~n8324;
  assign n8326 = ~pi370 & ~n8325;
  assign n8327 = ~n8322 & ~n8326;
  assign n8328 = pi371 & ~n8327;
  assign n8329 = pi370 & ~n8325;
  assign n8330 = ~pi370 & ~n8321;
  assign n8331 = ~n8329 & ~n8330;
  assign n8332 = ~pi371 & ~n8331;
  assign n8333 = ~n8328 & ~n8332;
  assign n8334 = pi373 & ~n8333;
  assign n8335 = pi371 & ~n8331;
  assign n8336 = ~pi371 & ~n8327;
  assign n8337 = ~n8335 & ~n8336;
  assign n8338 = ~pi373 & ~n8337;
  assign n8339 = ~n8334 & ~n8338;
  assign n8340 = ~pi375 & ~n8339;
  assign n8341 = pi373 & ~n8337;
  assign n8342 = ~pi373 & ~n8333;
  assign n8343 = ~n8341 & ~n8342;
  assign n8344 = pi375 & ~n8343;
  assign n8345 = n7775 & ~n8340;
  assign n8346 = ~n8344 & n8345;
  assign n8347 = ~pi375 & ~n8343;
  assign n8348 = pi375 & ~n8339;
  assign n8349 = ~n7775 & ~n8347;
  assign n8350 = ~n8348 & n8349;
  assign n8351 = ~pi591 & ~n8346;
  assign n8352 = ~n8350 & n8351;
  assign n8353 = ~pi590 & ~n8302;
  assign n8354 = ~n8352 & n8353;
  assign n8355 = n7356 & ~n8354;
  assign n8356 = ~n8230 & n8355;
  assign n8357 = pi591 & ~n7528;
  assign n8358 = n7849 & ~n8078;
  assign n8359 = n7528 & ~n8167;
  assign n8360 = n8170 & ~n8359;
  assign n8361 = n7528 & ~n8172;
  assign n8362 = n8175 & ~n8361;
  assign n8363 = ~n7849 & ~n8360;
  assign n8364 = ~n8362 & n8363;
  assign n8365 = pi1198 & ~n8358;
  assign n8366 = ~n8364 & n8365;
  assign n8367 = pi452 & n7819;
  assign n8368 = ~pi452 & ~n7819;
  assign n8369 = ~n8367 & ~n8368;
  assign n8370 = pi455 & ~n8369;
  assign n8371 = ~pi455 & n8369;
  assign n8372 = ~n8370 & ~n8371;
  assign n8373 = ~n7528 & ~n8372;
  assign n8374 = n8078 & n8372;
  assign n8375 = pi1196 & ~n8373;
  assign n8376 = ~n8374 & n8375;
  assign n8377 = ~pi1198 & ~n8045;
  assign n8378 = ~n8376 & n8377;
  assign n8379 = ~n8366 & ~n8378;
  assign n8380 = ~n7879 & ~n8379;
  assign n8381 = n7879 & n8078;
  assign n8382 = ~n8380 & ~n8381;
  assign n8383 = ~n7798 & n8382;
  assign n8384 = pi1199 & ~n8078;
  assign n8385 = pi351 & n8384;
  assign n8386 = ~n8383 & ~n8385;
  assign n8387 = ~pi461 & ~n8386;
  assign n8388 = ~n7909 & n8382;
  assign n8389 = ~pi351 & n8384;
  assign n8390 = ~n8388 & ~n8389;
  assign n8391 = pi461 & ~n8390;
  assign n8392 = ~n8387 & ~n8391;
  assign n8393 = ~n7887 & n8392;
  assign n8394 = ~pi461 & ~n8390;
  assign n8395 = pi461 & ~n8386;
  assign n8396 = ~n8394 & ~n8395;
  assign n8397 = n7887 & n8396;
  assign n8398 = ~n7899 & ~n8393;
  assign n8399 = ~n8397 & n8398;
  assign n8400 = ~n8222 & n8392;
  assign n8401 = n8222 & n8396;
  assign n8402 = n7899 & ~n8400;
  assign n8403 = ~n8401 & n8402;
  assign n8404 = ~pi591 & ~n8399;
  assign n8405 = ~n8403 & n8404;
  assign n8406 = pi590 & ~n8357;
  assign n8407 = ~n8405 & n8406;
  assign n8408 = ~n7528 & ~n8303;
  assign n8409 = ~n8305 & ~n8408;
  assign n8410 = pi374 & ~n8409;
  assign n8411 = ~pi1198 & n8409;
  assign n8412 = ~pi592 & n7528;
  assign n8413 = ~n8309 & ~n8412;
  assign n8414 = pi1198 & ~n8413;
  assign n8415 = ~n8411 & ~n8414;
  assign n8416 = ~pi374 & n8415;
  assign n8417 = ~n8410 & ~n8416;
  assign n8418 = ~pi369 & ~n8417;
  assign n8419 = ~pi374 & n8409;
  assign n8420 = pi374 & ~n8415;
  assign n8421 = ~n8419 & ~n8420;
  assign n8422 = pi369 & n8421;
  assign n8423 = ~n8418 & ~n8422;
  assign n8424 = pi370 & ~n8423;
  assign n8425 = pi369 & ~n8417;
  assign n8426 = ~pi369 & n8421;
  assign n8427 = ~n8425 & ~n8426;
  assign n8428 = ~pi370 & ~n8427;
  assign n8429 = pi371 & ~n7781;
  assign n8430 = ~pi371 & n7781;
  assign n8431 = ~n8429 & ~n8430;
  assign n8432 = ~n8424 & ~n8431;
  assign n8433 = ~n8428 & n8432;
  assign n8434 = pi370 & ~n8427;
  assign n8435 = ~pi370 & ~n8423;
  assign n8436 = n8431 & ~n8434;
  assign n8437 = ~n8435 & n8436;
  assign n8438 = ~pi591 & ~n8433;
  assign n8439 = ~n8437 & n8438;
  assign n8440 = n8076 & n8231;
  assign n8441 = n7420 & n7967;
  assign n8442 = ~n7360 & n7943;
  assign n8443 = n8441 & n8442;
  assign n8444 = n7654 & ~n8443;
  assign n8445 = ~pi592 & ~pi1196;
  assign n8446 = ~n8442 & n8445;
  assign n8447 = ~n8444 & ~n8446;
  assign n8448 = ~n7405 & ~n8447;
  assign n8449 = n7482 & ~n7967;
  assign n8450 = n7487 & ~n8449;
  assign n8451 = n7485 & ~n7941;
  assign n8452 = n7482 & ~n8451;
  assign n8453 = n8450 & ~n8452;
  assign n8454 = n7942 & n7967;
  assign n8455 = n6197 & ~n6221;
  assign n8456 = pi1093 & ~n6205;
  assign n8457 = n6221 & n8456;
  assign n8458 = n5727 & ~n8455;
  assign n8459 = ~n8457 & n8458;
  assign n8460 = n7542 & n8459;
  assign n8461 = pi299 & ~n8454;
  assign n8462 = ~n8460 & n8461;
  assign n8463 = ~n6194 & n6197;
  assign n8464 = n6194 & ~n6205;
  assign n8465 = n7506 & ~n8463;
  assign n8466 = ~n8464 & n8465;
  assign n8467 = n7542 & n8466;
  assign n8468 = ~pi299 & ~n8454;
  assign n8469 = ~n8467 & n8468;
  assign n8470 = pi39 & ~n8462;
  assign n8471 = ~n8469 & n8470;
  assign n8472 = ~n8453 & ~n8471;
  assign n8473 = ~pi38 & ~n8472;
  assign n8474 = pi38 & n7973;
  assign n8475 = ~pi100 & ~n8474;
  assign n8476 = pi38 & n7942;
  assign n8477 = ~pi100 & ~n8476;
  assign n8478 = ~n8475 & ~n8477;
  assign n8479 = ~n8473 & ~n8478;
  assign n8480 = n7538 & ~n8454;
  assign n8481 = ~n8479 & ~n8480;
  assign n8482 = ~pi87 & ~n8481;
  assign n8483 = ~n2628 & n7973;
  assign n8484 = pi87 & ~n8483;
  assign n8485 = ~n2628 & n7942;
  assign n8486 = pi87 & ~n8485;
  assign n8487 = ~n8484 & ~n8486;
  assign n8488 = n7429 & ~n7967;
  assign n8489 = n7429 & n7941;
  assign n8490 = n7436 & ~n8489;
  assign n8491 = ~n8488 & n8490;
  assign n8492 = ~n8487 & ~n8491;
  assign n8493 = ~n8482 & ~n8492;
  assign n8494 = ~pi75 & ~n8493;
  assign n8495 = ~n7408 & n7973;
  assign n8496 = pi75 & ~n8495;
  assign n8497 = ~n7408 & n7942;
  assign n8498 = pi75 & ~n8497;
  assign n8499 = ~n8496 & ~n8498;
  assign n8500 = ~pi1091 & ~n8454;
  assign n8501 = n7417 & ~n8500;
  assign n8502 = ~n8499 & ~n8501;
  assign n8503 = ~n8494 & ~n8502;
  assign n8504 = n8444 & ~n8503;
  assign n8505 = n8486 & ~n8490;
  assign n8506 = n7538 & ~n7942;
  assign n8507 = n7481 & ~n8452;
  assign n8508 = ~pi299 & n8467;
  assign n8509 = pi299 & n8460;
  assign n8510 = ~n8508 & ~n8509;
  assign n8511 = ~n7942 & n8510;
  assign n8512 = pi39 & ~n8511;
  assign n8513 = ~n8507 & ~n8512;
  assign n8514 = ~pi38 & ~n8513;
  assign n8515 = n8477 & ~n8514;
  assign n8516 = ~n8506 & ~n8515;
  assign n8517 = ~pi87 & ~n8516;
  assign n8518 = ~n8505 & ~n8517;
  assign n8519 = ~pi75 & ~n8518;
  assign n8520 = n7420 & ~n7941;
  assign n8521 = ~pi1091 & ~n8520;
  assign n8522 = n7417 & ~n8521;
  assign n8523 = n8498 & ~n8522;
  assign n8524 = ~n8519 & ~n8523;
  assign n8525 = n8446 & ~n8524;
  assign n8526 = ~n8504 & ~n8525;
  assign n8527 = pi567 & ~n8526;
  assign n8528 = pi1199 & ~n8448;
  assign n8529 = ~n8527 & n8528;
  assign n8530 = ~n7973 & n8510;
  assign n8531 = pi39 & ~n8530;
  assign n8532 = ~n8450 & ~n8531;
  assign n8533 = ~pi38 & ~n8532;
  assign n8534 = n8475 & ~n8533;
  assign n8535 = n7538 & ~n7973;
  assign n8536 = ~n8534 & ~n8535;
  assign n8537 = ~pi87 & ~n8536;
  assign n8538 = n7436 & ~n8488;
  assign n8539 = n8484 & ~n8538;
  assign n8540 = ~n8537 & ~n8539;
  assign n8541 = ~pi75 & ~n8540;
  assign n8542 = ~pi1091 & ~n8441;
  assign n8543 = n7417 & ~n8542;
  assign n8544 = n8496 & ~n8543;
  assign n8545 = ~n8541 & ~n8544;
  assign n8546 = pi567 & ~n8545;
  assign n8547 = n7405 & ~n8546;
  assign n8548 = ~n7360 & n7974;
  assign n8549 = n7654 & ~n8548;
  assign n8550 = ~n8547 & n8549;
  assign n8551 = ~pi1199 & ~n8045;
  assign n8552 = ~n8550 & n8551;
  assign n8553 = ~n8231 & ~n8552;
  assign n8554 = ~n8529 & n8553;
  assign n8555 = ~n8077 & ~n8440;
  assign n8556 = ~n8554 & n8555;
  assign n8557 = ~n8031 & ~n8556;
  assign n8558 = pi1197 & ~n8078;
  assign n8559 = pi333 & n8558;
  assign n8560 = ~n8557 & ~n8559;
  assign n8561 = ~pi391 & ~n8560;
  assign n8562 = ~n8027 & ~n8556;
  assign n8563 = ~pi333 & n8558;
  assign n8564 = ~n8562 & ~n8563;
  assign n8565 = pi391 & ~n8564;
  assign n8566 = ~n8561 & ~n8565;
  assign n8567 = pi392 & n8566;
  assign n8568 = ~pi391 & ~n8564;
  assign n8569 = pi391 & ~n8560;
  assign n8570 = ~n8568 & ~n8569;
  assign n8571 = ~pi392 & n8570;
  assign n8572 = ~n8020 & ~n8567;
  assign n8573 = ~n8571 & n8572;
  assign n8574 = ~pi392 & n8566;
  assign n8575 = pi392 & n8570;
  assign n8576 = n8020 & ~n8574;
  assign n8577 = ~n8575 & n8576;
  assign n8578 = pi591 & ~n8573;
  assign n8579 = ~n8577 & n8578;
  assign n8580 = ~pi590 & ~n8439;
  assign n8581 = ~n8579 & n8580;
  assign n8582 = ~n7356 & ~n8581;
  assign n8583 = ~n8407 & n8582;
  assign n8584 = ~pi588 & ~n8583;
  assign n8585 = ~n8356 & n8584;
  assign n8586 = ~po1038 & ~n8164;
  assign n8587 = ~n8585 & n8586;
  assign n8588 = ~pi217 & ~n8044;
  assign n8589 = ~n8587 & n8588;
  assign n8590 = ~n7576 & n7578;
  assign n8591 = ~n8589 & n8590;
  assign n8592 = pi1161 & ~pi1163;
  assign n8593 = n2923 & n8592;
  assign n8594 = ~pi31 & pi1162;
  assign n8595 = n8593 & n8594;
  assign po189 = n8591 | n8595;
  assign n8597 = ~pi74 & ~po1038;
  assign n8598 = n6078 & n8597;
  assign n8599 = n6112 & n6310;
  assign n8600 = po1057 & ~n7407;
  assign n8601 = pi252 & ~n8600;
  assign n8602 = pi129 & n2523;
  assign n8603 = ~n6090 & n8602;
  assign n8604 = n8601 & n8603;
  assign n8605 = ~n8599 & ~n8604;
  assign n8606 = pi100 & n2531;
  assign n8607 = ~pi137 & n8606;
  assign n8608 = ~n8605 & n8607;
  assign n8609 = ~pi24 & ~pi90;
  assign n8610 = n2916 & n8609;
  assign n8611 = n2702 & n2707;
  assign n8612 = pi50 & n2769;
  assign n8613 = n2495 & n8612;
  assign n8614 = ~pi93 & n8611;
  assign n8615 = n8613 & n8614;
  assign n8616 = n8610 & n8615;
  assign n8617 = pi829 & ~pi1093;
  assign n8618 = n6102 & n8617;
  assign po840 = n2926 | n8618;
  assign n8620 = ~n7356 & ~po840;
  assign n8621 = ~pi137 & ~n8620;
  assign n8622 = n8616 & ~n8621;
  assign n8623 = n2520 & n7376;
  assign n8624 = ~pi24 & n8612;
  assign n8625 = ~pi64 & ~pi81;
  assign n8626 = n2489 & n8625;
  assign n8627 = n2464 & n2803;
  assign n8628 = ~pi103 & n2470;
  assign n8629 = n8627 & n8628;
  assign n8630 = ~pi66 & ~pi84;
  assign n8631 = ~pi89 & ~pi102;
  assign n8632 = n7369 & n8631;
  assign n8633 = ~pi68 & ~pi73;
  assign n8634 = ~pi45 & ~pi48;
  assign n8635 = n2468 & n2484;
  assign n8636 = ~pi61 & ~pi104;
  assign n8637 = n8634 & n8636;
  assign n8638 = n8635 & n8637;
  assign n8639 = ~pi49 & pi76;
  assign n8640 = n2478 & n8639;
  assign n8641 = n8630 & n8633;
  assign n8642 = n8640 & n8641;
  assign n8643 = n8626 & n8632;
  assign n8644 = n8642 & n8643;
  assign n8645 = n8629 & n8638;
  assign n8646 = n8644 & n8645;
  assign n8647 = ~n8624 & ~n8646;
  assign n8648 = n2703 & n2707;
  assign n8649 = ~pi40 & n8623;
  assign n8650 = n8648 & n8649;
  assign n8651 = n8621 & n8650;
  assign n8652 = ~n8647 & n8651;
  assign n8653 = ~n8622 & ~n8652;
  assign n8654 = ~pi32 & ~n8653;
  assign n8655 = ~pi24 & ~pi841;
  assign n8656 = pi32 & ~n8655;
  assign n8657 = n2713 & n8656;
  assign n8658 = ~n8654 & ~n8657;
  assign n8659 = n6150 & ~n8658;
  assign n8660 = ~pi32 & ~n8616;
  assign n8661 = ~n6150 & ~n6152;
  assign n8662 = ~n8660 & n8661;
  assign n8663 = ~n8659 & ~n8662;
  assign n8664 = ~pi95 & n2532;
  assign n8665 = ~n8663 & n8664;
  assign n8666 = ~n8608 & ~n8665;
  assign n8667 = n2534 & ~n8666;
  assign n8668 = n7413 & ~po840;
  assign n8669 = ~pi87 & n2531;
  assign n8670 = pi75 & ~pi100;
  assign n8671 = n8669 & n8670;
  assign n8672 = n6090 & po1057;
  assign n8673 = ~pi137 & n8671;
  assign n8674 = ~n8601 & n8673;
  assign n8675 = ~n8672 & n8674;
  assign n8676 = n8668 & n8675;
  assign n8677 = ~n8667 & ~n8676;
  assign po190 = n8598 & ~n8677;
  assign n8679 = ~pi195 & ~pi196;
  assign n8680 = ~pi138 & n8679;
  assign n8681 = ~pi139 & n8680;
  assign n8682 = ~pi118 & n8681;
  assign n8683 = ~pi79 & n8682;
  assign n8684 = ~pi34 & n8683;
  assign n8685 = ~pi33 & ~n8684;
  assign n8686 = pi149 & pi157;
  assign n8687 = ~pi149 & ~pi157;
  assign n8688 = n6166 & ~n8687;
  assign n8689 = ~n8686 & n8688;
  assign n8690 = pi232 & n8689;
  assign n8691 = pi75 & ~n8690;
  assign n8692 = pi100 & ~n8690;
  assign n8693 = ~n8691 & ~n8692;
  assign n8694 = pi164 & n7406;
  assign n8695 = n7231 & n8694;
  assign n8696 = n8693 & ~n8695;
  assign n8697 = ~pi74 & ~n8696;
  assign n8698 = pi169 & n7406;
  assign n8699 = n7231 & n8698;
  assign n8700 = n8693 & ~n8699;
  assign n8701 = pi74 & ~n8700;
  assign n8702 = ~n3291 & ~n8697;
  assign n8703 = ~n8701 & n8702;
  assign n8704 = ~pi38 & ~pi54;
  assign n8705 = n8693 & n8704;
  assign n8706 = n8697 & ~n8705;
  assign n8707 = ~n8701 & ~n8706;
  assign n8708 = ~n2530 & ~n8707;
  assign n8709 = n3291 & ~n8708;
  assign n8710 = pi299 & ~n8689;
  assign n8711 = pi178 & pi183;
  assign n8712 = ~pi178 & ~pi183;
  assign n8713 = n6166 & ~n8712;
  assign n8714 = ~n8711 & n8713;
  assign n8715 = ~pi299 & ~n8714;
  assign n8716 = pi232 & ~n8710;
  assign n8717 = ~n8715 & n8716;
  assign n8718 = pi100 & ~n8717;
  assign n8719 = pi75 & ~n8717;
  assign n8720 = ~n8718 & ~n8719;
  assign n8721 = n7231 & n7406;
  assign n8722 = pi191 & ~pi299;
  assign n8723 = pi169 & pi299;
  assign n8724 = ~n8722 & ~n8723;
  assign n8725 = n8721 & ~n8724;
  assign n8726 = n8720 & ~n8725;
  assign n8727 = pi74 & ~n8726;
  assign n8728 = ~pi55 & ~n8727;
  assign n8729 = ~pi186 & ~pi299;
  assign n8730 = ~pi164 & pi299;
  assign n8731 = ~n8729 & ~n8730;
  assign n8732 = n7406 & n8731;
  assign n8733 = n7231 & n8732;
  assign n8734 = n8720 & ~n8733;
  assign n8735 = pi54 & ~n8734;
  assign n8736 = pi38 & n8732;
  assign n8737 = pi87 & ~n8736;
  assign n8738 = pi39 & pi232;
  assign n8739 = pi216 & n5726;
  assign n8740 = n6222 & n6341;
  assign n8741 = ~pi154 & ~n8740;
  assign n8742 = n6222 & ~n6349;
  assign n8743 = pi154 & ~n8742;
  assign n8744 = ~pi152 & ~n8741;
  assign n8745 = ~n8743 & n8744;
  assign n8746 = n6222 & n7542;
  assign n8747 = pi152 & pi154;
  assign n8748 = n8746 & n8747;
  assign n8749 = ~n8745 & ~n8748;
  assign n8750 = n8739 & ~n8749;
  assign n8751 = pi299 & ~n8750;
  assign n8752 = pi224 & n6359;
  assign n8753 = ~n6194 & n8752;
  assign n8754 = n6166 & n8753;
  assign n8755 = ~n6349 & n8754;
  assign n8756 = ~pi174 & n8755;
  assign n8757 = n7542 & n8754;
  assign n8758 = pi174 & n8757;
  assign n8759 = ~pi299 & ~n8756;
  assign n8760 = ~n8758 & n8759;
  assign n8761 = pi176 & ~n8760;
  assign n8762 = n6341 & n8754;
  assign n8763 = ~pi174 & n8762;
  assign n8764 = ~pi299 & ~n8763;
  assign n8765 = ~pi176 & ~n8764;
  assign n8766 = ~n8761 & ~n8765;
  assign n8767 = n8738 & ~n8751;
  assign n8768 = ~n8766 & n8767;
  assign n8769 = ~pi39 & pi232;
  assign n8770 = n3162 & n6166;
  assign n8771 = pi158 & n8770;
  assign n8772 = ~pi40 & n6166;
  assign n8773 = ~pi102 & n8625;
  assign n8774 = n2468 & n8773;
  assign n8775 = n2466 & n8774;
  assign n8776 = n2480 & n2486;
  assign n8777 = ~pi66 & pi73;
  assign n8778 = n8775 & n8777;
  assign n8779 = n8776 & n8778;
  assign n8780 = n2476 & n8779;
  assign n8781 = n8648 & n8780;
  assign n8782 = n2489 & n8781;
  assign n8783 = n8623 & n8782;
  assign n8784 = n2518 & n8783;
  assign n8785 = n8772 & n8784;
  assign n8786 = ~pi152 & n8785;
  assign n8787 = n2518 & n6166;
  assign n8788 = ~pi40 & n8787;
  assign n8789 = ~pi90 & n6132;
  assign n8790 = ~n7364 & ~n8789;
  assign n8791 = ~pi72 & n3080;
  assign n8792 = n7362 & n8791;
  assign n8793 = ~n8790 & n8792;
  assign n8794 = n8788 & n8793;
  assign n8795 = pi172 & n8794;
  assign n8796 = ~n8786 & ~n8795;
  assign n8797 = ~pi149 & ~n8796;
  assign n8798 = n3082 & n3174;
  assign n8799 = ~pi60 & n8612;
  assign n8800 = n2719 & ~n8799;
  assign n8801 = ~pi90 & n2717;
  assign n8802 = n2516 & n8801;
  assign n8803 = n2723 & n8802;
  assign n8804 = ~n8800 & n8803;
  assign n8805 = ~pi70 & ~n8804;
  assign n8806 = n2516 & ~n8790;
  assign n8807 = n8805 & ~n8806;
  assign n8808 = n8798 & ~n8807;
  assign n8809 = pi172 & n8808;
  assign n8810 = n8798 & ~n8805;
  assign n8811 = ~n6440 & ~n8810;
  assign n8812 = ~n8809 & n8811;
  assign n8813 = pi152 & ~n8812;
  assign n8814 = n2487 & n8775;
  assign n8815 = ~pi60 & n8814;
  assign n8816 = pi53 & ~n8815;
  assign n8817 = ~n8800 & ~n8816;
  assign n8818 = n2494 & n8780;
  assign n8819 = n2489 & ~n8818;
  assign n8820 = ~n8817 & n8819;
  assign n8821 = n2720 & ~n8820;
  assign n8822 = n2489 & n8803;
  assign n8823 = n8821 & n8822;
  assign n8824 = ~pi70 & ~n8823;
  assign n8825 = ~n8806 & n8824;
  assign n8826 = n8798 & ~n8825;
  assign n8827 = pi172 & n8826;
  assign n8828 = n8798 & ~n8824;
  assign n8829 = ~n6440 & ~n8828;
  assign n8830 = ~n8827 & n8829;
  assign n8831 = ~pi152 & ~n8830;
  assign n8832 = ~n8813 & ~n8831;
  assign n8833 = pi149 & n6166;
  assign n8834 = ~n8832 & n8833;
  assign n8835 = pi299 & ~n8771;
  assign n8836 = ~n8797 & n8835;
  assign n8837 = ~n8834 & n8836;
  assign n8838 = pi180 & n8770;
  assign n8839 = pi183 & n6166;
  assign n8840 = ~n6471 & ~n8828;
  assign n8841 = n8839 & ~n8840;
  assign n8842 = ~pi183 & n8785;
  assign n8843 = ~pi193 & ~n8842;
  assign n8844 = ~n8841 & n8843;
  assign n8845 = ~n6471 & ~n8826;
  assign n8846 = n8839 & ~n8845;
  assign n8847 = ~n8785 & ~n8794;
  assign n8848 = ~pi183 & ~n8847;
  assign n8849 = pi193 & ~n8848;
  assign n8850 = ~n8846 & n8849;
  assign n8851 = ~pi174 & ~n8844;
  assign n8852 = ~n8850 & n8851;
  assign n8853 = ~n6471 & ~n8808;
  assign n8854 = n6166 & ~n8853;
  assign n8855 = pi183 & ~n8854;
  assign n8856 = ~pi183 & ~n8794;
  assign n8857 = pi193 & ~n8856;
  assign n8858 = ~n8855 & n8857;
  assign n8859 = ~n6471 & ~n8810;
  assign n8860 = ~pi193 & n8839;
  assign n8861 = ~n8859 & n8860;
  assign n8862 = ~n8858 & ~n8861;
  assign n8863 = pi174 & ~n8862;
  assign n8864 = ~pi299 & ~n8838;
  assign n8865 = ~n8852 & n8864;
  assign n8866 = ~n8863 & n8865;
  assign n8867 = n8769 & ~n8837;
  assign n8868 = ~n8866 & n8867;
  assign n8869 = ~n8768 & ~n8868;
  assign n8870 = ~pi38 & ~n8869;
  assign n8871 = pi299 & n7406;
  assign n8872 = ~n6116 & n8871;
  assign n8873 = ~pi186 & ~n8872;
  assign n8874 = ~n6081 & n7406;
  assign n8875 = pi186 & ~n8874;
  assign n8876 = pi164 & ~n8875;
  assign n8877 = ~n8873 & n8876;
  assign n8878 = ~pi299 & n7406;
  assign n8879 = ~n6116 & n8878;
  assign n8880 = ~pi164 & pi186;
  assign n8881 = n8879 & n8880;
  assign n8882 = ~n8877 & ~n8881;
  assign n8883 = pi38 & ~n8882;
  assign n8884 = ~pi87 & ~n8883;
  assign n8885 = ~n8870 & n8884;
  assign n8886 = ~pi100 & ~n8737;
  assign n8887 = ~n8885 & n8886;
  assign n8888 = ~n8718 & ~n8887;
  assign n8889 = n2572 & ~n8888;
  assign n8890 = ~pi75 & pi92;
  assign n8891 = ~pi100 & n8736;
  assign n8892 = ~n8718 & ~n8891;
  assign n8893 = ~pi176 & ~pi299;
  assign n8894 = pi232 & ~n3361;
  assign n8895 = n6166 & ~n8893;
  assign n8896 = n8894 & n8895;
  assign n8897 = n2574 & n8896;
  assign n8898 = n6116 & n8897;
  assign n8899 = n8892 & ~n8898;
  assign n8900 = n8890 & ~n8899;
  assign n8901 = ~n8719 & ~n8900;
  assign n8902 = ~n8889 & n8901;
  assign n8903 = ~pi54 & ~n8902;
  assign n8904 = ~n8735 & ~n8903;
  assign n8905 = ~pi74 & ~n8904;
  assign n8906 = n8728 & ~n8905;
  assign n8907 = pi55 & ~n8701;
  assign n8908 = pi54 & ~n8696;
  assign n8909 = pi92 & n8693;
  assign n8910 = pi38 & n8695;
  assign n8911 = n8909 & ~n8910;
  assign n8912 = ~pi92 & ~n8691;
  assign n8913 = pi149 & n7406;
  assign n8914 = n6116 & n8913;
  assign n8915 = ~pi38 & ~n8914;
  assign n8916 = pi38 & ~n8694;
  assign n8917 = ~pi100 & ~n8916;
  assign n8918 = ~pi87 & n8917;
  assign n8919 = ~n8915 & n8918;
  assign n8920 = pi87 & n8694;
  assign n8921 = pi38 & ~pi100;
  assign n8922 = n8920 & n8921;
  assign n8923 = ~n8692 & ~n8922;
  assign n8924 = ~n8919 & n8923;
  assign n8925 = ~pi75 & ~n8924;
  assign n8926 = n8912 & ~n8925;
  assign n8927 = ~pi54 & ~n8911;
  assign n8928 = ~n8926 & n8927;
  assign n8929 = ~n8908 & ~n8928;
  assign n8930 = ~pi74 & ~n8929;
  assign n8931 = n8907 & ~n8930;
  assign n8932 = n2530 & ~n8931;
  assign n8933 = ~n8906 & n8932;
  assign n8934 = n8709 & ~n8933;
  assign n8935 = ~n8703 & ~n8934;
  assign n8936 = n8685 & ~n8935;
  assign n8937 = ~pi40 & n2489;
  assign n8938 = ~pi38 & n8937;
  assign n8939 = n7231 & n8938;
  assign n8940 = n2533 & n8939;
  assign n8941 = ~n2530 & n8940;
  assign n8942 = n2499 & n2502;
  assign n8943 = n2720 & n8942;
  assign n8944 = ~pi53 & n8943;
  assign n8945 = n8815 & n8944;
  assign n8946 = ~pi58 & n8945;
  assign n8947 = n7376 & n8946;
  assign n8948 = ~pi32 & n2520;
  assign n8949 = n8947 & n8948;
  assign n8950 = ~pi95 & n8949;
  assign n8951 = ~pi39 & ~n8913;
  assign n8952 = n8950 & n8951;
  assign n8953 = n8937 & ~n8952;
  assign n8954 = ~pi38 & ~n8953;
  assign n8955 = n8918 & ~n8954;
  assign n8956 = ~pi38 & ~n8937;
  assign n8957 = n8917 & ~n8956;
  assign n8958 = pi87 & n8957;
  assign n8959 = ~n8692 & ~n8958;
  assign n8960 = ~n8955 & n8959;
  assign n8961 = ~pi75 & ~n8960;
  assign n8962 = n8912 & ~n8961;
  assign n8963 = ~pi75 & n8957;
  assign n8964 = n8909 & ~n8963;
  assign n8965 = ~pi54 & ~n8964;
  assign n8966 = ~n8962 & n8965;
  assign n8967 = ~n8908 & ~n8966;
  assign n8968 = ~pi74 & ~n8967;
  assign n8969 = n8907 & ~n8968;
  assign n8970 = n2614 & n8950;
  assign n8971 = ~n8896 & n8970;
  assign n8972 = n2613 & n8937;
  assign n8973 = ~n8971 & n8972;
  assign n8974 = n8892 & ~n8973;
  assign n8975 = n8890 & ~n8974;
  assign n8976 = pi87 & ~n8972;
  assign n8977 = n8892 & n8976;
  assign n8978 = ~n8739 & n8937;
  assign n8979 = pi299 & ~n8978;
  assign n8980 = n6336 & ~n6340;
  assign n8981 = n6174 & n8980;
  assign n8982 = ~n6203 & ~n8981;
  assign n8983 = n8950 & ~n8982;
  assign n8984 = n6205 & n8983;
  assign n8985 = n8937 & ~n8984;
  assign n8986 = n6166 & n8983;
  assign n8987 = n8937 & ~n8986;
  assign n8988 = ~n6221 & ~n8987;
  assign n8989 = n8985 & ~n8988;
  assign n8990 = n8979 & ~n8989;
  assign n8991 = ~n8752 & n8937;
  assign n8992 = ~n8985 & ~n8991;
  assign n8993 = ~n6194 & ~n8987;
  assign n8994 = ~n8991 & n8993;
  assign n8995 = ~n8992 & ~n8994;
  assign n8996 = ~pi299 & ~n8995;
  assign n8997 = ~n8990 & ~n8996;
  assign n8998 = ~pi232 & n8997;
  assign n8999 = n8950 & n8981;
  assign n9000 = n2489 & ~n8999;
  assign n9001 = ~pi40 & n9000;
  assign n9002 = n6222 & ~n9001;
  assign n9003 = pi152 & n9002;
  assign n9004 = n8985 & ~n9003;
  assign n9005 = pi154 & ~n9004;
  assign n9006 = n6203 & n8950;
  assign n9007 = ~n6197 & n9006;
  assign n9008 = n8937 & ~n9007;
  assign n9009 = n6166 & n9008;
  assign n9010 = ~pi152 & n9009;
  assign n9011 = ~pi154 & ~n8989;
  assign n9012 = ~n9010 & n9011;
  assign n9013 = n8739 & ~n9005;
  assign n9014 = ~n9012 & n9013;
  assign n9015 = n8979 & ~n9014;
  assign n9016 = n6206 & n9006;
  assign n9017 = n8752 & n8937;
  assign n9018 = ~n9016 & n9017;
  assign n9019 = ~n8991 & ~n9018;
  assign n9020 = n8893 & n9019;
  assign n9021 = n6166 & n9001;
  assign n9022 = ~pi174 & ~n8992;
  assign n9023 = ~n9021 & ~n9022;
  assign n9024 = n8996 & n9023;
  assign n9025 = pi232 & ~n9020;
  assign n9026 = ~n9024 & n9025;
  assign n9027 = ~n9015 & n9026;
  assign n9028 = ~n8998 & ~n9027;
  assign n9029 = pi39 & ~n9028;
  assign n9030 = ~pi158 & pi299;
  assign n9031 = pi95 & ~n8937;
  assign n9032 = ~n2442 & ~n9031;
  assign n9033 = ~pi40 & ~pi479;
  assign n9034 = n2489 & ~n8949;
  assign n9035 = n9033 & n9034;
  assign n9036 = ~n9032 & ~n9035;
  assign n9037 = pi32 & ~n8937;
  assign n9038 = n2489 & ~n2507;
  assign n9039 = n2489 & ~n8947;
  assign n9040 = pi70 & ~n9039;
  assign n9041 = n2489 & ~n8945;
  assign n9042 = pi58 & ~n9041;
  assign n9043 = n8821 & n8942;
  assign n9044 = n2489 & ~n9043;
  assign n9045 = ~pi58 & ~n9044;
  assign n9046 = ~n9042 & ~n9045;
  assign n9047 = ~pi90 & ~n9046;
  assign n9048 = ~pi841 & n8946;
  assign n9049 = n2489 & ~n9048;
  assign n9050 = pi90 & ~n9049;
  assign n9051 = n2516 & ~n9050;
  assign n9052 = ~n9047 & n9051;
  assign n9053 = n2489 & ~n2516;
  assign n9054 = ~pi70 & ~n9053;
  assign n9055 = ~n9052 & n9054;
  assign n9056 = ~n9040 & ~n9055;
  assign n9057 = ~pi51 & ~n9056;
  assign n9058 = pi51 & ~n2489;
  assign n9059 = n2507 & ~n9058;
  assign n9060 = ~n9057 & n9059;
  assign n9061 = ~n9038 & ~n9060;
  assign n9062 = ~pi40 & ~n9061;
  assign n9063 = ~pi32 & ~n9062;
  assign n9064 = ~n9037 & ~n9063;
  assign n9065 = ~pi95 & ~n9064;
  assign n9066 = ~n9036 & ~n9065;
  assign n9067 = n8623 & n9048;
  assign n9068 = n8937 & ~n9067;
  assign n9069 = pi32 & ~n9068;
  assign n9070 = ~n9063 & ~n9069;
  assign n9071 = ~pi95 & ~n9070;
  assign n9072 = ~pi210 & n9071;
  assign n9073 = n9066 & ~n9072;
  assign n9074 = ~n6166 & n9073;
  assign n9075 = n6166 & ~n9031;
  assign n9076 = ~pi40 & ~n9037;
  assign n9077 = n2489 & ~n2510;
  assign n9078 = ~pi32 & ~n9077;
  assign n9079 = pi93 & ~n2489;
  assign n9080 = n2510 & ~n9079;
  assign n9081 = n2489 & ~n9042;
  assign n9082 = ~pi90 & ~n9081;
  assign n9083 = ~n9050 & ~n9082;
  assign n9084 = ~pi90 & n8781;
  assign n9085 = n9083 & ~n9084;
  assign n9086 = ~pi93 & ~n9085;
  assign n9087 = n9080 & ~n9086;
  assign n9088 = n9078 & ~n9087;
  assign n9089 = n9076 & ~n9088;
  assign n9090 = ~pi95 & ~n9089;
  assign n9091 = n9075 & ~n9090;
  assign n9092 = ~n9074 & ~n9091;
  assign n9093 = pi152 & ~n9092;
  assign n9094 = ~pi93 & ~n9083;
  assign n9095 = n9080 & ~n9094;
  assign n9096 = n9078 & ~n9095;
  assign n9097 = n9076 & ~n9096;
  assign n9098 = ~pi95 & ~n9097;
  assign n9099 = n9075 & ~n9098;
  assign n9100 = ~n9074 & ~n9099;
  assign n9101 = ~pi152 & ~n9100;
  assign n9102 = ~pi172 & ~n9093;
  assign n9103 = ~n9101 & n9102;
  assign n9104 = ~pi32 & n8623;
  assign n9105 = n8781 & n9104;
  assign n9106 = n8937 & ~n9105;
  assign n9107 = ~pi95 & ~n9106;
  assign n9108 = n9075 & ~n9107;
  assign n9109 = ~n9074 & ~n9108;
  assign n9110 = pi152 & ~n9109;
  assign n9111 = ~n6166 & ~n9073;
  assign n9112 = n6166 & ~n8937;
  assign n9113 = ~n9111 & ~n9112;
  assign n9114 = ~pi152 & n9113;
  assign n9115 = pi172 & ~n9110;
  assign n9116 = ~n9114 & n9115;
  assign n9117 = ~n9103 & ~n9116;
  assign n9118 = ~pi95 & ~n9117;
  assign n9119 = ~n9036 & ~n9118;
  assign n9120 = n9030 & ~n9119;
  assign n9121 = pi158 & pi299;
  assign n9122 = ~n9117 & n9121;
  assign n9123 = ~n9120 & ~n9122;
  assign n9124 = pi149 & ~n9123;
  assign n9125 = n2463 & n2516;
  assign n9126 = ~n2489 & ~n9125;
  assign n9127 = n8817 & n8943;
  assign n9128 = n2489 & ~n9127;
  assign n9129 = ~pi58 & ~n9128;
  assign n9130 = n7376 & n9129;
  assign n9131 = ~n9126 & ~n9130;
  assign n9132 = ~pi70 & ~n9131;
  assign n9133 = ~n9040 & ~n9132;
  assign n9134 = ~pi51 & ~n9133;
  assign n9135 = n9059 & ~n9134;
  assign n9136 = ~n9038 & ~n9135;
  assign n9137 = ~pi40 & ~n9136;
  assign n9138 = ~pi32 & ~n9137;
  assign n9139 = ~n9069 & ~n9138;
  assign n9140 = ~pi95 & ~n9139;
  assign n9141 = ~n9031 & ~n9140;
  assign n9142 = ~pi210 & ~n9141;
  assign n9143 = n6166 & ~n9142;
  assign n9144 = ~n9037 & ~n9138;
  assign n9145 = ~pi95 & ~n9144;
  assign n9146 = ~n9031 & ~n9145;
  assign n9147 = n9143 & n9146;
  assign n9148 = ~n9074 & ~n9147;
  assign n9149 = ~pi152 & ~n9148;
  assign n9150 = ~pi40 & ~n2489;
  assign n9151 = pi32 & ~n9150;
  assign n9152 = n7376 & n9045;
  assign n9153 = ~n9126 & ~n9152;
  assign n9154 = ~pi70 & ~n9153;
  assign n9155 = ~n9040 & ~n9154;
  assign n9156 = ~pi51 & ~n9155;
  assign n9157 = n9059 & ~n9156;
  assign n9158 = ~pi40 & ~n9038;
  assign n9159 = ~n9157 & n9158;
  assign n9160 = ~pi32 & ~n9159;
  assign n9161 = ~n9151 & ~n9160;
  assign n9162 = ~n2735 & ~n8937;
  assign n9163 = ~n9161 & ~n9162;
  assign n9164 = ~pi95 & ~n9163;
  assign n9165 = ~n9031 & ~n9164;
  assign n9166 = pi95 & ~n9150;
  assign n9167 = ~pi40 & ~n9068;
  assign n9168 = pi32 & ~n9167;
  assign n9169 = ~n9160 & ~n9168;
  assign n9170 = ~pi95 & ~n9169;
  assign n9171 = ~n9166 & ~n9170;
  assign n9172 = n9165 & ~n9171;
  assign n9173 = ~pi210 & ~n9172;
  assign n9174 = n6166 & ~n9173;
  assign n9175 = n9165 & n9174;
  assign n9176 = ~n9074 & ~n9175;
  assign n9177 = pi152 & ~n9176;
  assign n9178 = pi172 & ~n9149;
  assign n9179 = ~n9177 & n9178;
  assign n9180 = ~n9042 & ~n9129;
  assign n9181 = ~pi90 & ~n9180;
  assign n9182 = n9051 & ~n9181;
  assign n9183 = n9054 & ~n9182;
  assign n9184 = ~n9040 & ~n9183;
  assign n9185 = ~pi51 & ~n9184;
  assign n9186 = n9059 & ~n9185;
  assign n9187 = ~n9038 & ~n9186;
  assign n9188 = ~pi40 & ~n9187;
  assign n9189 = ~pi32 & ~n9188;
  assign n9190 = ~n9037 & ~n9189;
  assign n9191 = ~pi95 & ~n9190;
  assign n9192 = n9075 & ~n9191;
  assign n9193 = ~n9069 & ~n9189;
  assign n9194 = ~pi95 & ~n9193;
  assign n9195 = ~pi210 & n9194;
  assign n9196 = n9192 & ~n9195;
  assign n9197 = ~n9074 & ~n9196;
  assign n9198 = ~pi152 & ~n9197;
  assign n9199 = ~n9031 & ~n9065;
  assign n9200 = ~n9072 & n9199;
  assign n9201 = n6166 & ~n9200;
  assign n9202 = ~n9111 & ~n9201;
  assign n9203 = pi152 & n9202;
  assign n9204 = ~pi172 & ~n9198;
  assign n9205 = ~n9203 & n9204;
  assign n9206 = ~n9179 & ~n9205;
  assign n9207 = n9121 & ~n9206;
  assign n9208 = ~n9036 & ~n9145;
  assign n9209 = ~n9112 & ~n9143;
  assign n9210 = n9208 & ~n9209;
  assign n9211 = ~pi152 & ~n9210;
  assign n9212 = ~n9036 & ~n9164;
  assign n9213 = ~n9112 & ~n9174;
  assign n9214 = n9212 & ~n9213;
  assign n9215 = pi152 & ~n9214;
  assign n9216 = pi172 & ~n9211;
  assign n9217 = ~n9215 & n9216;
  assign n9218 = ~n9036 & ~n9191;
  assign n9219 = ~n9195 & n9218;
  assign n9220 = n6166 & n9219;
  assign n9221 = ~pi152 & ~n9220;
  assign n9222 = pi152 & ~n9073;
  assign n9223 = ~pi172 & ~n9221;
  assign n9224 = ~n9222 & n9223;
  assign n9225 = n9030 & ~n9074;
  assign n9226 = ~n9224 & n9225;
  assign n9227 = ~n9217 & n9226;
  assign n9228 = ~n9207 & ~n9227;
  assign n9229 = ~pi149 & ~n9228;
  assign n9230 = ~pi198 & n9071;
  assign n9231 = n9066 & ~n9230;
  assign n9232 = ~n6166 & n9231;
  assign n9233 = n6166 & ~n9107;
  assign n9234 = ~n9036 & n9233;
  assign n9235 = ~n9232 & ~n9234;
  assign n9236 = pi183 & ~n9235;
  assign n9237 = ~pi198 & ~n9172;
  assign n9238 = n6166 & ~n9237;
  assign n9239 = ~n9112 & ~n9238;
  assign n9240 = n9212 & ~n9239;
  assign n9241 = ~n9232 & ~n9240;
  assign n9242 = ~pi183 & ~n9241;
  assign n9243 = pi174 & ~n9236;
  assign n9244 = ~n9242 & n9243;
  assign n9245 = ~pi198 & n9140;
  assign n9246 = n9208 & ~n9245;
  assign n9247 = ~pi183 & n9246;
  assign n9248 = ~pi95 & ~n8937;
  assign n9249 = ~n9036 & ~n9248;
  assign n9250 = pi183 & n9249;
  assign n9251 = ~n9247 & ~n9250;
  assign n9252 = n6166 & ~n9251;
  assign n9253 = ~pi174 & ~n9252;
  assign n9254 = ~n9232 & n9253;
  assign n9255 = ~pi180 & ~n9254;
  assign n9256 = ~n9244 & n9255;
  assign n9257 = n9165 & n9238;
  assign n9258 = ~n9232 & ~n9257;
  assign n9259 = ~pi183 & ~n9258;
  assign n9260 = ~n9108 & ~n9232;
  assign n9261 = pi183 & ~n9260;
  assign n9262 = pi174 & ~n9261;
  assign n9263 = ~n9259 & n9262;
  assign n9264 = ~n6166 & ~n9231;
  assign n9265 = ~n9112 & ~n9264;
  assign n9266 = pi183 & n9265;
  assign n9267 = ~pi40 & n9136;
  assign n9268 = ~pi32 & ~n9267;
  assign n9269 = ~n9168 & ~n9268;
  assign n9270 = ~pi95 & ~n9269;
  assign n9271 = ~pi198 & n9270;
  assign n9272 = ~n9151 & ~n9268;
  assign n9273 = ~pi95 & ~n9272;
  assign n9274 = pi198 & n9273;
  assign n9275 = ~n9166 & ~n9271;
  assign n9276 = ~n9274 & n9275;
  assign n9277 = n8772 & ~n9276;
  assign n9278 = ~n9232 & ~n9277;
  assign n9279 = ~pi183 & ~n9278;
  assign n9280 = ~pi174 & ~n9266;
  assign n9281 = ~n9279 & n9280;
  assign n9282 = pi180 & ~n9263;
  assign n9283 = ~n9281 & n9282;
  assign n9284 = ~n9256 & ~n9283;
  assign n9285 = pi193 & ~n9284;
  assign n9286 = ~n8839 & ~n9231;
  assign n9287 = ~n9036 & ~n9090;
  assign n9288 = n6166 & ~n9287;
  assign n9289 = pi183 & n9288;
  assign n9290 = pi174 & ~n9289;
  assign n9291 = ~n9286 & n9290;
  assign n9292 = ~pi198 & n9194;
  assign n9293 = n9192 & ~n9292;
  assign n9294 = ~n9232 & ~n9293;
  assign n9295 = ~pi183 & ~n9294;
  assign n9296 = ~n9099 & ~n9232;
  assign n9297 = pi183 & ~n9296;
  assign n9298 = ~n9295 & ~n9297;
  assign n9299 = ~pi95 & n9298;
  assign n9300 = ~pi174 & ~n9036;
  assign n9301 = ~n9299 & n9300;
  assign n9302 = ~pi180 & ~n9291;
  assign n9303 = ~n9301 & n9302;
  assign n9304 = ~pi174 & ~n9298;
  assign n9305 = n9199 & ~n9230;
  assign n9306 = n8772 & n9305;
  assign n9307 = ~n9232 & ~n9306;
  assign n9308 = ~pi183 & n9307;
  assign n9309 = ~n9091 & ~n9232;
  assign n9310 = pi183 & n9309;
  assign n9311 = pi174 & ~n9308;
  assign n9312 = ~n9310 & n9311;
  assign n9313 = pi180 & ~n9304;
  assign n9314 = ~n9312 & n9313;
  assign n9315 = ~pi193 & ~n9303;
  assign n9316 = ~n9314 & n9315;
  assign n9317 = ~pi299 & ~n9285;
  assign n9318 = ~n9316 & n9317;
  assign n9319 = ~n9124 & ~n9229;
  assign n9320 = ~n9318 & n9319;
  assign n9321 = pi232 & ~n9320;
  assign n9322 = n6150 & n9071;
  assign n9323 = n9066 & ~n9322;
  assign n9324 = ~pi232 & ~n9323;
  assign n9325 = ~pi39 & ~n9324;
  assign n9326 = ~n9321 & n9325;
  assign n9327 = ~n9029 & ~n9326;
  assign n9328 = ~pi38 & ~n9327;
  assign n9329 = ~n8883 & ~n9328;
  assign n9330 = ~pi100 & ~n9329;
  assign n9331 = ~pi87 & ~n8718;
  assign n9332 = ~n9330 & n9331;
  assign n9333 = n2572 & ~n8977;
  assign n9334 = ~n9332 & n9333;
  assign n9335 = ~n8719 & ~n8975;
  assign n9336 = ~n9334 & n9335;
  assign n9337 = ~pi54 & ~n9336;
  assign n9338 = ~n8735 & ~n9337;
  assign n9339 = ~pi74 & ~n9338;
  assign n9340 = n8728 & ~n9339;
  assign n9341 = n2530 & ~n8969;
  assign n9342 = ~n9340 & n9341;
  assign n9343 = n8709 & ~n8941;
  assign n9344 = ~n9342 & n9343;
  assign n9345 = ~n8703 & ~n9344;
  assign n9346 = ~n8685 & ~n9345;
  assign n9347 = ~pi954 & ~n8936;
  assign n9348 = ~n9346 & n9347;
  assign n9349 = pi33 & ~n8935;
  assign n9350 = ~pi33 & ~n9345;
  assign n9351 = pi954 & ~n9349;
  assign n9352 = ~n9350 & n9351;
  assign po191 = ~n9348 & ~n9352;
  assign n9354 = pi197 & n8687;
  assign n9355 = ~pi197 & ~n8687;
  assign n9356 = ~n9354 & ~n9355;
  assign n9357 = pi162 & n6166;
  assign n9358 = n9356 & ~n9357;
  assign n9359 = n9354 & n9357;
  assign n9360 = ~pi162 & ~pi197;
  assign n9361 = n8688 & ~n9360;
  assign n9362 = n6166 & ~n9361;
  assign n9363 = ~n9359 & n9362;
  assign n9364 = ~n9356 & ~n9363;
  assign n9365 = ~n9358 & ~n9364;
  assign n9366 = pi232 & ~n7231;
  assign n9367 = n9365 & n9366;
  assign n9368 = pi167 & n8721;
  assign n9369 = ~n9367 & ~n9368;
  assign n9370 = ~pi74 & n9369;
  assign n9371 = pi148 & n8721;
  assign n9372 = pi74 & ~n9371;
  assign n9373 = ~n9367 & n9372;
  assign n9374 = ~n9370 & ~n9373;
  assign n9375 = ~n3291 & n9374;
  assign n9376 = ~pi54 & ~n9367;
  assign n9377 = pi38 & n9368;
  assign n9378 = n9376 & ~n9377;
  assign n9379 = ~pi74 & n9378;
  assign n9380 = n9374 & ~n9379;
  assign n9381 = ~n2530 & ~n9380;
  assign n9382 = n3291 & ~n9381;
  assign n9383 = pi140 & pi145;
  assign n9384 = n8712 & ~n9383;
  assign n9385 = ~pi140 & ~pi145;
  assign n9386 = n6166 & ~n9385;
  assign n9387 = n9384 & n9386;
  assign n9388 = ~n9383 & ~n9385;
  assign n9389 = n8713 & ~n9388;
  assign n9390 = ~pi299 & ~n9387;
  assign n9391 = ~n9389 & n9390;
  assign n9392 = pi299 & ~n9365;
  assign n9393 = pi232 & ~n9391;
  assign n9394 = ~n9392 & n9393;
  assign n9395 = pi100 & ~n9394;
  assign n9396 = pi75 & ~n9394;
  assign n9397 = ~n9395 & ~n9396;
  assign n9398 = pi141 & ~pi299;
  assign n9399 = pi148 & pi299;
  assign n9400 = ~n9398 & ~n9399;
  assign n9401 = n7406 & ~n9400;
  assign n9402 = n7231 & ~n9401;
  assign n9403 = n9397 & ~n9402;
  assign n9404 = pi74 & ~n9403;
  assign n9405 = ~pi55 & ~n9404;
  assign n9406 = ~pi167 & pi299;
  assign n9407 = ~pi188 & ~pi299;
  assign n9408 = ~n9406 & ~n9407;
  assign n9409 = n7406 & n9408;
  assign n9410 = ~pi100 & ~n9409;
  assign n9411 = ~pi75 & n9410;
  assign n9412 = n9397 & ~n9411;
  assign n9413 = pi54 & ~n9412;
  assign n9414 = ~pi38 & pi155;
  assign n9415 = ~pi161 & ~n8742;
  assign n9416 = pi161 & ~n8746;
  assign n9417 = n8739 & ~n9415;
  assign n9418 = ~n9416 & n9417;
  assign n9419 = n9414 & ~n9418;
  assign n9420 = ~pi38 & ~pi155;
  assign n9421 = ~pi161 & n8739;
  assign n9422 = n8740 & n9421;
  assign n9423 = n9420 & ~n9422;
  assign n9424 = ~n9419 & ~n9423;
  assign n9425 = pi299 & ~n9424;
  assign n9426 = ~pi177 & ~pi299;
  assign n9427 = ~pi144 & n8762;
  assign n9428 = n9426 & ~n9427;
  assign n9429 = ~pi144 & n8755;
  assign n9430 = pi177 & ~pi299;
  assign n9431 = pi144 & n8757;
  assign n9432 = ~n9429 & n9430;
  assign n9433 = ~n9431 & n9432;
  assign n9434 = pi232 & ~n9428;
  assign n9435 = ~n9433 & n9434;
  assign n9436 = ~pi38 & ~n9435;
  assign n9437 = ~n9425 & ~n9436;
  assign n9438 = pi39 & ~n9437;
  assign n9439 = ~pi167 & pi188;
  assign n9440 = n8879 & n9439;
  assign n9441 = ~pi188 & ~n8872;
  assign n9442 = pi188 & ~n8874;
  assign n9443 = pi167 & ~n9442;
  assign n9444 = ~n9441 & n9443;
  assign n9445 = pi38 & ~n9440;
  assign n9446 = ~n9444 & n9445;
  assign n9447 = pi159 & n3162;
  assign n9448 = ~pi146 & n8826;
  assign n9449 = ~pi161 & n8829;
  assign n9450 = ~n9448 & n9449;
  assign n9451 = ~pi146 & n8808;
  assign n9452 = pi161 & ~n9451;
  assign n9453 = n8811 & n9452;
  assign n9454 = pi162 & ~n9453;
  assign n9455 = ~n9450 & n9454;
  assign n9456 = ~n9447 & ~n9455;
  assign n9457 = n6166 & ~n9456;
  assign n9458 = ~pi146 & n8794;
  assign n9459 = ~pi161 & n8785;
  assign n9460 = ~n9458 & ~n9459;
  assign n9461 = ~pi162 & ~n9460;
  assign n9462 = pi299 & ~n9461;
  assign n9463 = ~n9457 & n9462;
  assign n9464 = pi181 & n8770;
  assign n9465 = ~pi142 & n8808;
  assign n9466 = pi144 & ~n9465;
  assign n9467 = n8859 & n9466;
  assign n9468 = ~pi142 & n8826;
  assign n9469 = ~pi144 & n8840;
  assign n9470 = ~n9468 & n9469;
  assign n9471 = pi140 & n6166;
  assign n9472 = ~n9467 & n9471;
  assign n9473 = ~n9470 & n9472;
  assign n9474 = ~pi142 & n8794;
  assign n9475 = ~pi144 & n8785;
  assign n9476 = ~n9474 & ~n9475;
  assign n9477 = ~pi140 & ~n9476;
  assign n9478 = ~pi299 & ~n9464;
  assign n9479 = ~n9477 & n9478;
  assign n9480 = ~n9473 & n9479;
  assign n9481 = pi232 & ~n9480;
  assign n9482 = ~n9463 & n9481;
  assign n9483 = n2531 & ~n9482;
  assign n9484 = ~n9438 & ~n9446;
  assign n9485 = ~n9483 & n9484;
  assign n9486 = ~pi100 & ~n9485;
  assign n9487 = ~n9395 & ~n9486;
  assign n9488 = ~pi87 & ~n9487;
  assign n9489 = ~n2613 & ~n9410;
  assign n9490 = ~n9395 & n9489;
  assign n9491 = pi87 & ~n9490;
  assign n9492 = ~n9488 & ~n9491;
  assign n9493 = n2572 & ~n9492;
  assign n9494 = pi38 & n9408;
  assign n9495 = ~pi155 & pi299;
  assign n9496 = ~n9426 & ~n9495;
  assign n9497 = n2531 & n9496;
  assign n9498 = n2513 & n9497;
  assign n9499 = ~n9494 & ~n9498;
  assign n9500 = n7406 & ~n9499;
  assign n9501 = ~pi100 & ~n9500;
  assign n9502 = ~n9395 & ~n9501;
  assign n9503 = ~pi87 & ~n9502;
  assign n9504 = ~n9491 & ~n9503;
  assign n9505 = n8890 & ~n9504;
  assign n9506 = ~n9396 & ~n9505;
  assign n9507 = ~n9493 & n9506;
  assign n9508 = ~pi54 & ~n9507;
  assign n9509 = ~n9413 & ~n9508;
  assign n9510 = ~pi74 & ~n9509;
  assign n9511 = n9405 & ~n9510;
  assign n9512 = pi55 & ~n9373;
  assign n9513 = pi54 & n9369;
  assign n9514 = pi167 & n7406;
  assign n9515 = pi38 & n9514;
  assign n9516 = ~pi92 & pi162;
  assign n9517 = n7230 & n9516;
  assign n9518 = n8769 & n9517;
  assign n9519 = n6185 & n9518;
  assign n9520 = ~n9515 & ~n9519;
  assign n9521 = n7231 & ~n9520;
  assign n9522 = n9376 & ~n9521;
  assign n9523 = ~n9513 & ~n9522;
  assign n9524 = ~pi74 & ~n9523;
  assign n9525 = n9512 & ~n9524;
  assign n9526 = n2530 & ~n9525;
  assign n9527 = ~n9511 & n9526;
  assign n9528 = n9382 & ~n9527;
  assign n9529 = ~n9375 & ~n9528;
  assign n9530 = pi34 & n9529;
  assign n9531 = ~n2530 & ~n8940;
  assign n9532 = n3291 & ~n9531;
  assign n9533 = ~n9382 & ~n9532;
  assign n9534 = ~n8939 & n9378;
  assign n9535 = ~n6078 & ~n9534;
  assign n9536 = pi162 & n7406;
  assign n9537 = n8970 & ~n9536;
  assign n9538 = n8938 & ~n9537;
  assign n9539 = ~n9515 & ~n9538;
  assign n9540 = n7231 & ~n9539;
  assign n9541 = ~n9367 & ~n9540;
  assign n9542 = ~pi92 & ~n9541;
  assign n9543 = ~n9535 & ~n9542;
  assign n9544 = ~n9513 & ~n9543;
  assign n9545 = ~pi74 & ~n9544;
  assign n9546 = n9512 & ~n9545;
  assign n9547 = ~pi38 & ~n8997;
  assign n9548 = ~pi232 & ~n9547;
  assign n9549 = ~pi161 & n9009;
  assign n9550 = ~n8989 & ~n9549;
  assign n9551 = n8739 & ~n9550;
  assign n9552 = n9420 & ~n9551;
  assign n9553 = pi161 & n9002;
  assign n9554 = n8739 & n8985;
  assign n9555 = ~n9553 & n9554;
  assign n9556 = n9414 & ~n9555;
  assign n9557 = ~n9552 & ~n9556;
  assign n9558 = n8979 & ~n9557;
  assign n9559 = pi144 & n8995;
  assign n9560 = ~pi144 & ~n8992;
  assign n9561 = ~n9019 & n9560;
  assign n9562 = n9426 & ~n9561;
  assign n9563 = ~n9559 & n9562;
  assign n9564 = ~n9021 & n9430;
  assign n9565 = ~n9560 & n9564;
  assign n9566 = ~n8995 & n9565;
  assign n9567 = ~n9563 & ~n9566;
  assign n9568 = ~pi38 & ~n9567;
  assign n9569 = pi232 & ~n9558;
  assign n9570 = ~n9568 & n9569;
  assign n9571 = pi39 & ~n9548;
  assign n9572 = ~n9570 & n9571;
  assign n9573 = ~pi159 & pi299;
  assign n9574 = ~pi146 & n9113;
  assign n9575 = pi146 & ~n9100;
  assign n9576 = ~pi161 & ~n9574;
  assign n9577 = ~n9575 & n9576;
  assign n9578 = pi146 & ~n9092;
  assign n9579 = ~pi146 & ~n9109;
  assign n9580 = pi161 & ~n9578;
  assign n9581 = ~n9579 & n9580;
  assign n9582 = ~n9577 & ~n9581;
  assign n9583 = ~pi95 & ~n9582;
  assign n9584 = ~n9036 & ~n9583;
  assign n9585 = pi162 & ~n9584;
  assign n9586 = ~pi161 & n9220;
  assign n9587 = pi161 & n9073;
  assign n9588 = pi146 & ~n9586;
  assign n9589 = ~n9587 & n9588;
  assign n9590 = ~pi161 & n9210;
  assign n9591 = pi161 & n9214;
  assign n9592 = ~pi146 & ~n9590;
  assign n9593 = ~n9591 & n9592;
  assign n9594 = ~n9589 & ~n9593;
  assign n9595 = ~pi162 & ~n9074;
  assign n9596 = ~n9594 & n9595;
  assign n9597 = ~n9585 & ~n9596;
  assign n9598 = n9573 & ~n9597;
  assign n9599 = pi159 & pi299;
  assign n9600 = pi146 & n9202;
  assign n9601 = ~pi146 & ~n9176;
  assign n9602 = pi161 & ~n9600;
  assign n9603 = ~n9601 & n9602;
  assign n9604 = pi146 & ~n9197;
  assign n9605 = ~pi146 & ~n9148;
  assign n9606 = ~pi161 & ~n9604;
  assign n9607 = ~n9605 & n9606;
  assign n9608 = ~pi162 & ~n9603;
  assign n9609 = ~n9607 & n9608;
  assign n9610 = pi162 & n9582;
  assign n9611 = n9599 & ~n9609;
  assign n9612 = ~n9610 & n9611;
  assign n9613 = ~pi142 & ~n9260;
  assign n9614 = pi142 & ~n9309;
  assign n9615 = ~n9613 & ~n9614;
  assign n9616 = ~pi95 & n9615;
  assign n9617 = ~n9036 & ~n9616;
  assign n9618 = pi140 & ~n9617;
  assign n9619 = pi142 & n9231;
  assign n9620 = ~pi142 & ~n9241;
  assign n9621 = ~pi140 & ~n9619;
  assign n9622 = ~n9620 & n9621;
  assign n9623 = ~pi181 & ~n9622;
  assign n9624 = ~n9618 & n9623;
  assign n9625 = ~pi142 & ~n9258;
  assign n9626 = pi142 & ~n9307;
  assign n9627 = ~pi140 & ~n9626;
  assign n9628 = ~n9625 & n9627;
  assign n9629 = pi140 & n9615;
  assign n9630 = pi181 & ~n9628;
  assign n9631 = ~n9629 & n9630;
  assign n9632 = pi144 & ~n9631;
  assign n9633 = ~n9624 & n9632;
  assign n9634 = n9218 & ~n9292;
  assign n9635 = ~pi140 & n9634;
  assign n9636 = ~n9036 & ~n9098;
  assign n9637 = pi140 & n9636;
  assign n9638 = pi142 & ~n9637;
  assign n9639 = ~n9635 & n9638;
  assign n9640 = ~pi140 & n9246;
  assign n9641 = pi140 & n9249;
  assign n9642 = ~pi142 & ~n9641;
  assign n9643 = ~n9640 & n9642;
  assign n9644 = ~n9639 & ~n9643;
  assign n9645 = n6166 & ~n9644;
  assign n9646 = ~pi181 & ~n9264;
  assign n9647 = ~n9645 & n9646;
  assign n9648 = pi142 & ~n9294;
  assign n9649 = ~pi142 & ~n9278;
  assign n9650 = ~pi140 & ~n9648;
  assign n9651 = ~n9649 & n9650;
  assign n9652 = ~pi142 & n9265;
  assign n9653 = pi142 & ~n9296;
  assign n9654 = pi140 & ~n9652;
  assign n9655 = ~n9653 & n9654;
  assign n9656 = pi181 & ~n9651;
  assign n9657 = ~n9655 & n9656;
  assign n9658 = ~pi144 & ~n9647;
  assign n9659 = ~n9657 & n9658;
  assign n9660 = ~n9633 & ~n9659;
  assign n9661 = ~pi299 & ~n9660;
  assign n9662 = ~n9598 & ~n9612;
  assign n9663 = ~n9661 & n9662;
  assign n9664 = pi232 & ~n9663;
  assign n9665 = ~n9324 & ~n9664;
  assign n9666 = n2531 & ~n9665;
  assign n9667 = ~pi87 & ~n9446;
  assign n9668 = ~n9572 & n9667;
  assign n9669 = ~n9666 & n9668;
  assign n9670 = pi38 & ~n9409;
  assign n9671 = ~n8956 & ~n9670;
  assign n9672 = pi87 & n9671;
  assign n9673 = ~pi100 & ~n9672;
  assign n9674 = ~n9669 & n9673;
  assign n9675 = ~n9395 & ~n9674;
  assign n9676 = n2572 & ~n9675;
  assign n9677 = ~pi38 & ~n9496;
  assign n9678 = n7406 & ~n9677;
  assign n9679 = n8970 & ~n9678;
  assign n9680 = n9671 & ~n9679;
  assign n9681 = ~pi100 & ~n9680;
  assign n9682 = ~n9395 & ~n9681;
  assign n9683 = n8890 & ~n9682;
  assign n9684 = ~n9396 & ~n9683;
  assign n9685 = ~n9676 & n9684;
  assign n9686 = ~pi54 & ~n9685;
  assign n9687 = ~n9413 & ~n9686;
  assign n9688 = ~pi74 & ~n9687;
  assign n9689 = n9405 & ~n9688;
  assign n9690 = n2530 & ~n9546;
  assign n9691 = ~n9689 & n9690;
  assign n9692 = ~n9533 & ~n9691;
  assign n9693 = ~n9375 & ~n9692;
  assign n9694 = ~pi34 & n9693;
  assign n9695 = ~pi33 & ~pi954;
  assign n9696 = ~n9530 & ~n9695;
  assign n9697 = ~n9694 & n9696;
  assign n9698 = ~pi34 & ~n8683;
  assign n9699 = n9529 & n9698;
  assign n9700 = n9693 & ~n9698;
  assign n9701 = n9695 & ~n9699;
  assign n9702 = ~n9700 & n9701;
  assign po192 = ~n9697 & ~n9702;
  assign n9704 = n2530 & n2577;
  assign n9705 = n7413 & n9704;
  assign n9706 = ~pi55 & n9705;
  assign n9707 = pi59 & ~n9706;
  assign n9708 = pi137 & n8599;
  assign n9709 = ~pi137 & n8601;
  assign n9710 = ~n6179 & n7348;
  assign n9711 = pi683 & n9710;
  assign n9712 = n6089 & n7406;
  assign n9713 = pi252 & ~n9711;
  assign n9714 = po1057 & n9713;
  assign n9715 = ~n9712 & n9714;
  assign n9716 = ~n9709 & ~n9715;
  assign n9717 = n8603 & n9716;
  assign n9718 = ~n9708 & ~n9717;
  assign n9719 = n8606 & ~n9718;
  assign n9720 = ~pi93 & ~n8789;
  assign n9721 = ~n6138 & ~n9720;
  assign n9722 = ~pi35 & ~n9721;
  assign n9723 = pi35 & ~n2915;
  assign n9724 = ~pi32 & n2521;
  assign n9725 = ~n9723 & n9724;
  assign n9726 = ~n9722 & n9725;
  assign n9727 = pi32 & ~pi93;
  assign n9728 = n8610 & n9727;
  assign n9729 = n7363 & n9728;
  assign n9730 = ~n9726 & ~n9729;
  assign n9731 = ~pi95 & n6150;
  assign n9732 = ~n9730 & n9731;
  assign n9733 = pi1082 & n2742;
  assign n9734 = ~pi1082 & n6150;
  assign n9735 = ~n9722 & ~n9734;
  assign n9736 = ~pi137 & n6150;
  assign n9737 = ~pi122 & n2926;
  assign n9738 = ~n7356 & ~n9737;
  assign n9739 = ~pi122 & ~po740;
  assign n9740 = n7356 & ~n9739;
  assign n9741 = n2495 & n8646;
  assign n9742 = n2709 & n8611;
  assign n9743 = n9741 & n9742;
  assign n9744 = n9722 & ~n9743;
  assign n9745 = ~n9736 & ~n9738;
  assign n9746 = ~n9740 & n9745;
  assign n9747 = ~n9744 & n9746;
  assign n9748 = ~n9735 & ~n9747;
  assign n9749 = n2521 & ~n9723;
  assign n9750 = ~n9748 & n9749;
  assign n9751 = ~n9733 & ~n9750;
  assign n9752 = n2518 & ~n9751;
  assign n9753 = ~pi38 & ~n9732;
  assign n9754 = ~n9752 & n9753;
  assign n9755 = pi38 & ~n7413;
  assign n9756 = ~pi39 & ~pi100;
  assign n9757 = ~n9755 & n9756;
  assign n9758 = ~n9754 & n9757;
  assign n9759 = ~n9719 & ~n9758;
  assign n9760 = n2534 & ~n9759;
  assign n9761 = ~pi24 & n8671;
  assign n9762 = pi137 & ~po840;
  assign n9763 = ~n8672 & n9762;
  assign n9764 = ~n8601 & ~n9763;
  assign n9765 = n9761 & ~n9764;
  assign n9766 = n2523 & n9765;
  assign n9767 = ~n9760 & ~n9766;
  assign n9768 = ~pi92 & ~n9767;
  assign n9769 = ~pi54 & ~n9768;
  assign n9770 = ~pi24 & n7270;
  assign n9771 = pi54 & ~n9770;
  assign n9772 = n2530 & n6246;
  assign n9773 = ~n9771 & n9772;
  assign n9774 = ~n9769 & n9773;
  assign n9775 = ~pi59 & ~n9774;
  assign n9776 = ~pi57 & ~n9707;
  assign po193 = ~n9775 & n9776;
  assign n9778 = n6431 & n8623;
  assign n9779 = n2532 & n6074;
  assign n9780 = ~po1038 & n9779;
  assign n9781 = ~pi74 & n9780;
  assign n9782 = n9778 & n9781;
  assign n9783 = ~pi77 & n2767;
  assign n9784 = n2720 & n9783;
  assign n9785 = n2717 & n9784;
  assign n9786 = ~pi65 & n2464;
  assign n9787 = n2489 & n9786;
  assign n9788 = n8773 & n9787;
  assign n9789 = ~pi69 & n9788;
  assign n9790 = ~pi67 & ~pi71;
  assign n9791 = ~pi83 & n2801;
  assign n9792 = pi36 & ~pi103;
  assign n9793 = n9790 & n9792;
  assign n9794 = n9789 & n9793;
  assign n9795 = n9791 & n9794;
  assign n9796 = n9785 & n9795;
  assign n9797 = ~pi58 & n7457;
  assign n9798 = ~n9796 & ~n9797;
  assign n9799 = po740 & n9782;
  assign po194 = ~n9798 & n9799;
  assign n9801 = ~pi45 & ~pi49;
  assign n9802 = n2481 & n9801;
  assign n9803 = ~pi71 & n2489;
  assign n9804 = ~pi104 & n2471;
  assign n9805 = n9803 & n9804;
  assign n9806 = ~pi48 & ~pi65;
  assign n9807 = pi89 & n9806;
  assign n9808 = n9802 & n9807;
  assign n9809 = n8776 & n9808;
  assign n9810 = n9805 & n9809;
  assign n9811 = pi332 & n9810;
  assign n9812 = ~pi64 & ~n9811;
  assign n9813 = ~pi81 & ~n2787;
  assign n9814 = n6431 & n9125;
  assign n9815 = n2503 & n9814;
  assign n9816 = n2520 & n9815;
  assign n9817 = ~pi39 & ~pi841;
  assign n9818 = n2467 & n9817;
  assign n9819 = ~n9812 & n9818;
  assign n9820 = n9816 & n9819;
  assign n9821 = n9813 & n9820;
  assign n9822 = ~pi38 & ~n9821;
  assign n9823 = ~pi39 & ~pi95;
  assign n9824 = ~pi32 & n9823;
  assign n9825 = pi24 & n2712;
  assign n9826 = n2701 & n9825;
  assign n9827 = n9824 & n9826;
  assign n9828 = pi38 & ~n9827;
  assign n9829 = n2573 & n7293;
  assign n9830 = ~po1038 & n9829;
  assign n9831 = ~n9822 & n9830;
  assign po196 = ~n9828 & n9831;
  assign n9833 = ~pi38 & n9830;
  assign n9834 = ~pi984 & ~n6102;
  assign n9835 = pi835 & ~n9834;
  assign n9836 = n6169 & ~n9835;
  assign n9837 = n6180 & ~n9836;
  assign n9838 = pi1093 & n9837;
  assign n9839 = n6170 & n6333;
  assign n9840 = ~n9838 & n9839;
  assign n9841 = ~pi215 & n9840;
  assign n9842 = n6205 & n9837;
  assign n9843 = n9839 & ~n9842;
  assign n9844 = n6221 & n9843;
  assign n9845 = ~n6197 & n9837;
  assign n9846 = n9839 & ~n9845;
  assign n9847 = ~n6221 & n9846;
  assign n9848 = pi299 & ~n9844;
  assign n9849 = ~n9847 & n9848;
  assign n9850 = ~n9841 & n9849;
  assign n9851 = ~pi223 & n9840;
  assign n9852 = n6194 & n9843;
  assign n9853 = ~n6194 & n9846;
  assign n9854 = ~pi299 & ~n9852;
  assign n9855 = ~n9853 & n9854;
  assign n9856 = ~n9851 & n9855;
  assign n9857 = pi786 & ~pi1082;
  assign n9858 = ~n9850 & ~n9857;
  assign n9859 = ~n9856 & n9858;
  assign n9860 = n5966 & ~n6223;
  assign n9861 = n5783 & ~n6207;
  assign n9862 = ~n9860 & ~n9861;
  assign n9863 = po740 & n9857;
  assign n9864 = ~n9862 & n9863;
  assign n9865 = n6335 & n9864;
  assign n9866 = ~n9859 & ~n9865;
  assign n9867 = pi39 & ~n9866;
  assign n9868 = ~n6150 & n6438;
  assign n9869 = pi35 & ~n6435;
  assign n9870 = n2520 & ~n9869;
  assign n9871 = ~pi986 & ~po740;
  assign n9872 = pi252 & ~n9871;
  assign n9873 = pi314 & ~n9872;
  assign n9874 = ~pi49 & n8633;
  assign n9875 = n8625 & n8630;
  assign n9876 = ~pi65 & ~pi69;
  assign n9877 = n9875 & n9876;
  assign n9878 = ~pi83 & ~pi103;
  assign n9879 = ~pi45 & pi48;
  assign n9880 = n2478 & n9879;
  assign n9881 = n9878 & n9880;
  assign n9882 = n8627 & n8632;
  assign n9883 = n9874 & n9882;
  assign n9884 = n9877 & n9881;
  assign n9885 = n9883 & n9884;
  assign n9886 = n9805 & n9885;
  assign n9887 = ~pi47 & ~pi841;
  assign n9888 = n9886 & n9887;
  assign n9889 = ~n2760 & ~n9888;
  assign n9890 = n2501 & n2705;
  assign n9891 = ~n9873 & n9890;
  assign n9892 = ~n9889 & n9891;
  assign n9893 = pi108 & n7458;
  assign n9894 = n2772 & n9893;
  assign n9895 = ~n2773 & n7458;
  assign n9896 = ~pi841 & n2494;
  assign n9897 = n2720 & n9896;
  assign n9898 = ~pi97 & n9897;
  assign n9899 = n9886 & n9898;
  assign n9900 = n9895 & n9899;
  assign n9901 = ~pi47 & ~n9894;
  assign n9902 = ~n9900 & n9901;
  assign n9903 = n6130 & n9873;
  assign n9904 = ~n9902 & n9903;
  assign n9905 = ~n9892 & ~n9904;
  assign n9906 = n2709 & ~n9905;
  assign n9907 = ~pi35 & ~n9906;
  assign n9908 = n2462 & n9870;
  assign n9909 = ~n9907 & n9908;
  assign n9910 = ~n9868 & ~n9909;
  assign n9911 = n9823 & ~n9910;
  assign n9912 = ~n9867 & ~n9911;
  assign po197 = n9833 & ~n9912;
  assign n9914 = n2518 & ~n3387;
  assign n9915 = pi102 & n2931;
  assign n9916 = n2466 & n9915;
  assign n9917 = n2510 & n9916;
  assign n9918 = n2503 & n9917;
  assign n9919 = n2492 & n9918;
  assign n9920 = ~pi40 & ~n9919;
  assign n9921 = n9914 & ~n9920;
  assign n9922 = ~pi1082 & ~n9921;
  assign n9923 = n6431 & n9919;
  assign n9924 = pi1082 & ~n9923;
  assign n9925 = n9781 & ~n9924;
  assign po198 = ~n9922 & n9925;
  assign n9927 = ~pi189 & n6166;
  assign n9928 = pi144 & n9927;
  assign n9929 = ~pi174 & n9928;
  assign n9930 = ~pi299 & ~n9929;
  assign n9931 = ~pi166 & n6166;
  assign n9932 = pi161 & n9931;
  assign n9933 = ~pi152 & n9932;
  assign n9934 = ~n6084 & ~n9933;
  assign n9935 = pi232 & ~n9930;
  assign n9936 = ~n9934 & n9935;
  assign n9937 = ~pi72 & ~n9936;
  assign n9938 = pi39 & ~n9937;
  assign n9939 = ~pi41 & ~pi72;
  assign n9940 = ~pi39 & ~n9939;
  assign n9941 = ~n9938 & ~n9940;
  assign n9942 = ~n7360 & ~n9941;
  assign n9943 = ~n2574 & n9941;
  assign n9944 = ~n7440 & ~n9939;
  assign n9945 = ~n2922 & n9939;
  assign n9946 = n7440 & ~n9945;
  assign n9947 = ~pi41 & pi72;
  assign n9948 = n2922 & ~n9947;
  assign n9949 = ~pi44 & n2523;
  assign n9950 = ~pi101 & n9949;
  assign n9951 = n7411 & n9950;
  assign n9952 = n7414 & n9951;
  assign n9953 = pi41 & ~n9952;
  assign n9954 = ~pi99 & n6098;
  assign n9955 = ~pi72 & pi101;
  assign n9956 = ~pi41 & ~n9955;
  assign n9957 = pi252 & n6431;
  assign n9958 = ~pi24 & n2712;
  assign n9959 = n7411 & n9957;
  assign n9960 = n9958 & n9959;
  assign n9961 = ~pi44 & n9960;
  assign n9962 = n9956 & n9961;
  assign n9963 = ~n9954 & n9962;
  assign n9964 = n9948 & ~n9963;
  assign n9965 = ~n9953 & n9964;
  assign n9966 = n9946 & ~n9965;
  assign n9967 = ~n9944 & ~n9966;
  assign n9968 = ~pi39 & ~n9967;
  assign n9969 = n2574 & ~n9938;
  assign n9970 = ~n9968 & n9969;
  assign n9971 = pi75 & ~n9943;
  assign n9972 = ~n9970 & n9971;
  assign n9973 = ~n2613 & n9940;
  assign n9974 = ~pi228 & n9939;
  assign n9975 = n2712 & n6431;
  assign n9976 = ~pi44 & n9975;
  assign n9977 = n9956 & n9976;
  assign n9978 = ~n9947 & ~n9977;
  assign n9979 = pi41 & ~n9950;
  assign n9980 = pi228 & n9978;
  assign n9981 = ~n9979 & n9980;
  assign n9982 = n2628 & ~n9974;
  assign n9983 = ~n9981 & n9982;
  assign n9984 = pi87 & ~n9973;
  assign n9985 = ~n9938 & n9984;
  assign n9986 = ~n9983 & n9985;
  assign n9987 = pi38 & ~n9941;
  assign n9988 = ~pi72 & ~n7411;
  assign n9989 = ~n9978 & ~n9988;
  assign n9990 = ~n9954 & n9989;
  assign n9991 = pi41 & ~n9951;
  assign n9992 = n2922 & ~n9954;
  assign n9993 = ~n9948 & ~n9992;
  assign n9994 = ~n9991 & ~n9993;
  assign n9995 = ~n9990 & n9994;
  assign n9996 = n9946 & ~n9995;
  assign n9997 = ~n9944 & ~n9996;
  assign n9998 = ~pi39 & ~n9997;
  assign n9999 = ~n9938 & ~n9998;
  assign n10000 = n6082 & ~n9999;
  assign n10001 = pi287 & n2523;
  assign n10002 = n9936 & n10001;
  assign n10003 = ~n9937 & ~n10002;
  assign n10004 = pi39 & ~n10003;
  assign n10005 = ~pi250 & pi252;
  assign n10006 = pi901 & ~pi959;
  assign n10007 = ~pi480 & pi949;
  assign n10008 = n2711 & n10007;
  assign n10009 = n2706 & n2758;
  assign n10010 = pi110 & n10009;
  assign n10011 = n10008 & n10010;
  assign n10012 = ~n10006 & ~n10011;
  assign n10013 = n2717 & n2777;
  assign n10014 = n2711 & n10013;
  assign n10015 = ~n10007 & n10014;
  assign n10016 = ~pi109 & n2498;
  assign n10017 = n2777 & n10016;
  assign n10018 = ~pi110 & ~n10017;
  assign n10019 = n2706 & n10008;
  assign n10020 = ~n2759 & n10019;
  assign n10021 = ~n10018 & n10020;
  assign n10022 = n10006 & ~n10015;
  assign n10023 = ~n10021 & n10022;
  assign n10024 = n6431 & n10005;
  assign n10025 = ~n10012 & n10024;
  assign n10026 = ~n10023 & n10025;
  assign n10027 = ~pi72 & n10026;
  assign n10028 = n9778 & n10010;
  assign n10029 = ~n10005 & n10007;
  assign n10030 = n10028 & n10029;
  assign n10031 = ~n10027 & ~n10030;
  assign n10032 = ~pi44 & ~n10031;
  assign n10033 = ~pi101 & n10032;
  assign n10034 = pi41 & ~n10033;
  assign n10035 = pi44 & ~pi72;
  assign n10036 = n6431 & ~n10005;
  assign n10037 = n10011 & n10036;
  assign n10038 = ~pi72 & ~n10037;
  assign n10039 = ~n10026 & n10038;
  assign n10040 = ~n10035 & ~n10039;
  assign n10041 = ~pi101 & ~n10040;
  assign n10042 = n9956 & ~n10041;
  assign n10043 = ~n10034 & ~n10042;
  assign n10044 = ~pi228 & ~n10043;
  assign n10045 = pi1093 & ~n7381;
  assign n10046 = ~pi44 & ~n10045;
  assign n10047 = ~n7393 & n10046;
  assign n10048 = ~pi101 & n10047;
  assign n10049 = pi41 & ~n10048;
  assign n10050 = ~pi72 & ~n7381;
  assign n10051 = ~n7395 & n10050;
  assign n10052 = ~n10035 & ~n10051;
  assign n10053 = ~pi101 & ~n10052;
  assign n10054 = n9956 & ~n10053;
  assign n10055 = ~n2922 & ~n10054;
  assign n10056 = ~n10049 & n10055;
  assign n10057 = n2928 & ~n7374;
  assign n10058 = n2930 & n10057;
  assign n10059 = ~n7457 & ~n10058;
  assign n10060 = n2463 & ~n10059;
  assign n10061 = n7365 & ~n10060;
  assign n10062 = n7362 & ~n10061;
  assign n10063 = ~pi51 & ~n10062;
  assign n10064 = ~n2747 & ~n10063;
  assign n10065 = ~pi96 & ~n10064;
  assign n10066 = ~pi122 & n7471;
  assign n10067 = ~n10065 & n10066;
  assign n10068 = pi1093 & ~n7384;
  assign n10069 = ~n10067 & n10068;
  assign n10070 = ~n7393 & ~n10069;
  assign n10071 = ~pi44 & n10070;
  assign n10072 = ~pi101 & n10071;
  assign n10073 = pi41 & ~n10072;
  assign n10074 = ~pi72 & ~n10072;
  assign n10075 = ~pi41 & ~n10074;
  assign n10076 = n2922 & ~n10075;
  assign n10077 = ~n10073 & n10076;
  assign n10078 = pi228 & ~n10056;
  assign n10079 = ~n10077 & n10078;
  assign n10080 = ~pi39 & ~n10044;
  assign n10081 = ~n10079 & n10080;
  assign n10082 = n2613 & ~n10004;
  assign n10083 = ~n10081 & n10082;
  assign n10084 = ~pi87 & ~n9987;
  assign n10085 = ~n10000 & n10084;
  assign n10086 = ~n10083 & n10085;
  assign n10087 = ~pi75 & ~n9986;
  assign n10088 = ~n10086 & n10087;
  assign n10089 = ~n9972 & ~n10088;
  assign n10090 = n7360 & ~n10089;
  assign n10091 = ~po1038 & ~n9942;
  assign n10092 = ~n10090 & n10091;
  assign n10093 = n8738 & n9933;
  assign n10094 = ~pi72 & ~n9940;
  assign n10095 = po1038 & n10094;
  assign n10096 = ~n10093 & n10095;
  assign po199 = ~n10092 & ~n10096;
  assign n10098 = pi211 & pi214;
  assign n10099 = pi212 & n10098;
  assign n10100 = ~pi219 & ~n10099;
  assign n10101 = pi207 & pi208;
  assign n10102 = ~pi72 & pi199;
  assign n10103 = ~pi232 & ~n10102;
  assign n10104 = ~pi299 & ~n10103;
  assign n10105 = ~pi72 & ~n9927;
  assign n10106 = pi199 & n10105;
  assign n10107 = pi232 & ~n10106;
  assign n10108 = n10104 & ~n10107;
  assign n10109 = pi39 & ~n10108;
  assign n10110 = pi42 & ~pi72;
  assign n10111 = ~n2574 & n10110;
  assign n10112 = ~n7440 & ~n10110;
  assign n10113 = ~pi115 & n2922;
  assign n10114 = n10110 & ~n10113;
  assign n10115 = n7440 & ~n10114;
  assign n10116 = pi114 & ~n10110;
  assign n10117 = n10113 & ~n10116;
  assign n10118 = n6092 & n9961;
  assign n10119 = ~pi113 & n10118;
  assign n10120 = ~pi116 & n10119;
  assign n10121 = n10110 & ~n10120;
  assign n10122 = n6091 & n9950;
  assign n10123 = n6095 & n10122;
  assign n10124 = n7411 & n10123;
  assign n10125 = ~pi114 & ~n6094;
  assign n10126 = n10124 & n10125;
  assign n10127 = ~pi42 & n10126;
  assign n10128 = n7414 & n10127;
  assign n10129 = ~pi114 & ~n10121;
  assign n10130 = ~n10128 & n10129;
  assign n10131 = n10117 & ~n10130;
  assign n10132 = n10115 & ~n10131;
  assign n10133 = n2574 & ~n10112;
  assign n10134 = ~n10132 & n10133;
  assign n10135 = ~pi39 & ~n10111;
  assign n10136 = ~n10134 & n10135;
  assign n10137 = ~n10109 & ~n10136;
  assign n10138 = pi75 & ~n10137;
  assign n10139 = ~pi39 & ~n10110;
  assign n10140 = ~n2613 & n10139;
  assign n10141 = n6092 & n9976;
  assign n10142 = pi228 & n10141;
  assign n10143 = n6097 & n10142;
  assign n10144 = n10110 & ~n10143;
  assign n10145 = ~pi42 & n6096;
  assign n10146 = pi228 & n10145;
  assign n10147 = n10123 & n10146;
  assign n10148 = n2628 & ~n10144;
  assign n10149 = ~n10147 & n10148;
  assign n10150 = pi87 & ~n10140;
  assign n10151 = ~n10149 & n10150;
  assign n10152 = ~n10109 & n10151;
  assign n10153 = ~n10109 & ~n10139;
  assign n10154 = pi38 & ~n10153;
  assign n10155 = n6095 & n10141;
  assign n10156 = ~pi72 & ~n10155;
  assign n10157 = ~n9988 & ~n10156;
  assign n10158 = pi42 & ~n10157;
  assign n10159 = ~pi114 & ~n10158;
  assign n10160 = ~n10127 & n10159;
  assign n10161 = n10117 & ~n10160;
  assign n10162 = n10115 & ~n10161;
  assign n10163 = ~n10112 & ~n10162;
  assign n10164 = ~pi39 & ~n10163;
  assign n10165 = ~n10109 & ~n10164;
  assign n10166 = n6082 & ~n10165;
  assign n10167 = n6166 & n10001;
  assign n10168 = ~pi189 & n10167;
  assign n10169 = ~n10105 & ~n10168;
  assign n10170 = pi199 & ~n10169;
  assign n10171 = pi232 & ~n10170;
  assign n10172 = n10104 & ~n10171;
  assign n10173 = pi39 & ~n10172;
  assign n10174 = pi115 & ~n10110;
  assign n10175 = n6091 & n10033;
  assign n10176 = n6095 & n10175;
  assign n10177 = ~pi42 & ~n10176;
  assign n10178 = ~pi72 & pi116;
  assign n10179 = pi72 & ~n6091;
  assign n10180 = ~pi99 & n10042;
  assign n10181 = ~n10179 & ~n10180;
  assign n10182 = ~pi72 & pi113;
  assign n10183 = ~n10181 & ~n10182;
  assign n10184 = ~n10178 & n10183;
  assign n10185 = pi42 & ~pi114;
  assign n10186 = n10184 & n10185;
  assign n10187 = ~n10116 & ~n10177;
  assign n10188 = ~n10186 & n10187;
  assign n10189 = ~pi115 & ~n10188;
  assign n10190 = ~pi228 & ~n10174;
  assign n10191 = ~n10189 & n10190;
  assign n10192 = ~pi113 & n6091;
  assign n10193 = n10072 & n10192;
  assign n10194 = ~pi116 & n10193;
  assign n10195 = ~pi114 & n10194;
  assign n10196 = ~pi42 & n10195;
  assign n10197 = n10110 & ~n10195;
  assign n10198 = n10113 & ~n10196;
  assign n10199 = ~n10197 & n10198;
  assign n10200 = pi72 & ~n10192;
  assign n10201 = ~pi99 & ~pi113;
  assign n10202 = n10054 & n10201;
  assign n10203 = ~n10200 & ~n10202;
  assign n10204 = ~n10178 & ~n10203;
  assign n10205 = pi42 & ~n10204;
  assign n10206 = n6091 & n10048;
  assign n10207 = n6095 & n10206;
  assign n10208 = ~pi42 & n10207;
  assign n10209 = ~pi114 & ~n10208;
  assign n10210 = ~n10205 & n10209;
  assign n10211 = ~n10116 & ~n10210;
  assign n10212 = ~pi115 & ~n2922;
  assign n10213 = ~n10211 & n10212;
  assign n10214 = pi228 & ~n10174;
  assign n10215 = ~n10199 & n10214;
  assign n10216 = ~n10213 & n10215;
  assign n10217 = ~pi39 & ~n10191;
  assign n10218 = ~n10216 & n10217;
  assign n10219 = ~n10173 & ~n10218;
  assign n10220 = n2613 & ~n10219;
  assign n10221 = ~pi87 & ~n10154;
  assign n10222 = ~n10166 & n10221;
  assign n10223 = ~n10220 & n10222;
  assign n10224 = ~pi75 & ~n10152;
  assign n10225 = ~n10223 & n10224;
  assign n10226 = n7360 & ~n10138;
  assign n10227 = ~n10225 & n10226;
  assign n10228 = ~n7360 & n10153;
  assign n10229 = ~n10101 & ~n10228;
  assign n10230 = ~n10227 & n10229;
  assign n10231 = ~pi72 & pi200;
  assign n10232 = ~pi232 & ~n10231;
  assign n10233 = ~pi299 & ~n10232;
  assign n10234 = pi200 & n10105;
  assign n10235 = pi232 & ~n10234;
  assign n10236 = n10233 & ~n10235;
  assign n10237 = pi39 & ~n10236;
  assign n10238 = ~n10108 & n10237;
  assign n10239 = ~n10139 & ~n10238;
  assign n10240 = ~n7360 & n10239;
  assign n10241 = n10101 & ~n10240;
  assign n10242 = ~n10136 & ~n10238;
  assign n10243 = pi75 & ~n10242;
  assign n10244 = n10151 & ~n10238;
  assign n10245 = ~n10164 & ~n10238;
  assign n10246 = n6082 & ~n10245;
  assign n10247 = pi38 & ~n10239;
  assign n10248 = ~pi87 & ~n10247;
  assign n10249 = ~n10104 & ~n10233;
  assign n10250 = pi200 & ~n10169;
  assign n10251 = pi232 & ~n10250;
  assign n10252 = ~n10170 & n10251;
  assign n10253 = ~n10249 & ~n10252;
  assign n10254 = pi39 & ~n10253;
  assign n10255 = ~n10218 & ~n10254;
  assign n10256 = n2613 & ~n10255;
  assign n10257 = ~n10246 & n10248;
  assign n10258 = ~n10256 & n10257;
  assign n10259 = ~pi75 & ~n10244;
  assign n10260 = ~n10258 & n10259;
  assign n10261 = n7360 & ~n10243;
  assign n10262 = ~n10260 & n10261;
  assign n10263 = n10241 & ~n10262;
  assign n10264 = ~n10230 & ~n10263;
  assign n10265 = n10100 & ~n10264;
  assign n10266 = pi232 & n9931;
  assign n10267 = ~pi72 & ~n10266;
  assign n10268 = pi299 & n10267;
  assign n10269 = pi39 & ~n10268;
  assign n10270 = ~n10108 & n10269;
  assign n10271 = ~n10139 & ~n10270;
  assign n10272 = ~n7360 & n10271;
  assign n10273 = ~n10136 & ~n10270;
  assign n10274 = pi75 & ~n10273;
  assign n10275 = n10151 & ~n10270;
  assign n10276 = n9931 & n10001;
  assign n10277 = pi232 & pi299;
  assign n10278 = ~n10267 & n10277;
  assign n10279 = ~n10276 & n10278;
  assign n10280 = ~pi299 & n10171;
  assign n10281 = pi72 & ~pi232;
  assign n10282 = pi299 & ~n10281;
  assign n10283 = n10103 & ~n10282;
  assign n10284 = ~n10279 & ~n10283;
  assign n10285 = ~n10280 & n10284;
  assign n10286 = pi39 & ~n10285;
  assign n10287 = ~n10218 & ~n10286;
  assign n10288 = n2613 & ~n10287;
  assign n10289 = ~n10164 & ~n10270;
  assign n10290 = n6082 & ~n10289;
  assign n10291 = pi38 & ~n10271;
  assign n10292 = ~pi87 & ~n10291;
  assign n10293 = ~n10290 & n10292;
  assign n10294 = ~n10288 & n10293;
  assign n10295 = ~pi75 & ~n10275;
  assign n10296 = ~n10294 & n10295;
  assign n10297 = n7360 & ~n10274;
  assign n10298 = ~n10296 & n10297;
  assign n10299 = ~n10101 & ~n10298;
  assign n10300 = n10237 & n10270;
  assign n10301 = ~n10136 & ~n10300;
  assign n10302 = pi75 & ~n10301;
  assign n10303 = n10151 & ~n10300;
  assign n10304 = ~n10231 & n10283;
  assign n10305 = ~pi299 & n10251;
  assign n10306 = ~n10170 & n10305;
  assign n10307 = ~n10279 & ~n10304;
  assign n10308 = ~n10306 & n10307;
  assign n10309 = pi39 & ~n10308;
  assign n10310 = ~n10218 & ~n10309;
  assign n10311 = n2613 & ~n10310;
  assign n10312 = ~n10248 & ~n10292;
  assign n10313 = ~n10164 & ~n10300;
  assign n10314 = n6082 & ~n10313;
  assign n10315 = ~n10312 & ~n10314;
  assign n10316 = ~n10311 & n10315;
  assign n10317 = ~pi75 & ~n10303;
  assign n10318 = ~n10316 & n10317;
  assign n10319 = n7360 & ~n10302;
  assign n10320 = ~n10318 & n10319;
  assign n10321 = n10241 & ~n10320;
  assign n10322 = ~n10299 & ~n10321;
  assign n10323 = ~n10100 & ~n10272;
  assign n10324 = ~n10322 & n10323;
  assign n10325 = ~po1038 & ~n10265;
  assign n10326 = ~n10324 & n10325;
  assign n10327 = ~n10100 & n10267;
  assign n10328 = pi39 & ~n10327;
  assign n10329 = po1038 & ~n10139;
  assign n10330 = ~n10328 & n10329;
  assign po200 = n10326 | n10330;
  assign n10332 = pi212 & pi214;
  assign n10333 = ~pi211 & ~pi219;
  assign n10334 = n10332 & ~n10333;
  assign n10335 = ~pi211 & ~n10332;
  assign n10336 = ~n10334 & ~n10335;
  assign n10337 = ~n10236 & n10269;
  assign n10338 = pi43 & ~pi72;
  assign n10339 = ~n2574 & n10338;
  assign n10340 = ~n7440 & ~n10338;
  assign n10341 = n2922 & n10145;
  assign n10342 = n10338 & ~n10341;
  assign n10343 = n7440 & ~n10342;
  assign n10344 = ~pi72 & ~n10120;
  assign n10345 = pi43 & n10344;
  assign n10346 = ~pi43 & pi52;
  assign n10347 = n7414 & n10124;
  assign n10348 = n10346 & n10347;
  assign n10349 = ~n10345 & ~n10348;
  assign n10350 = n10341 & ~n10349;
  assign n10351 = n10343 & ~n10350;
  assign n10352 = n2574 & ~n10340;
  assign n10353 = ~n10351 & n10352;
  assign n10354 = ~pi39 & ~n10339;
  assign n10355 = ~n10353 & n10354;
  assign n10356 = ~n10337 & ~n10355;
  assign n10357 = pi75 & ~n10356;
  assign n10358 = ~pi39 & ~n10338;
  assign n10359 = ~n2613 & n10358;
  assign n10360 = ~pi43 & n10145;
  assign n10361 = pi228 & n10360;
  assign n10362 = n10123 & n10361;
  assign n10363 = pi228 & n10155;
  assign n10364 = n10145 & n10363;
  assign n10365 = n10338 & ~n10364;
  assign n10366 = n2532 & ~n10362;
  assign n10367 = ~n10365 & n10366;
  assign n10368 = pi87 & ~n10359;
  assign n10369 = ~n10367 & n10368;
  assign n10370 = ~n10337 & n10369;
  assign n10371 = ~n10337 & ~n10358;
  assign n10372 = pi38 & ~n10371;
  assign n10373 = n10124 & n10346;
  assign n10374 = pi43 & ~n10157;
  assign n10375 = ~n10373 & ~n10374;
  assign n10376 = n10341 & ~n10375;
  assign n10377 = n10343 & ~n10376;
  assign n10378 = ~n10340 & ~n10377;
  assign n10379 = ~pi39 & ~n10378;
  assign n10380 = ~n10337 & ~n10379;
  assign n10381 = n6082 & ~n10380;
  assign n10382 = ~pi228 & ~n10176;
  assign n10383 = ~n2922 & ~n10206;
  assign n10384 = n6091 & n10072;
  assign n10385 = n2922 & ~n10384;
  assign n10386 = ~pi113 & ~n10383;
  assign n10387 = ~n10385 & n10386;
  assign n10388 = ~pi116 & n10387;
  assign n10389 = pi228 & ~n10388;
  assign n10390 = ~n10382 & ~n10389;
  assign n10391 = ~pi43 & ~n10390;
  assign n10392 = n10145 & ~n10391;
  assign n10393 = ~n10338 & ~n10392;
  assign n10394 = ~pi99 & ~n10055;
  assign n10395 = ~n10076 & n10394;
  assign n10396 = n6095 & n10395;
  assign n10397 = ~pi72 & ~n10396;
  assign n10398 = pi228 & ~n10397;
  assign n10399 = ~pi228 & n10184;
  assign n10400 = ~n10398 & ~n10399;
  assign n10401 = pi43 & n10145;
  assign n10402 = ~n10400 & n10401;
  assign n10403 = ~n10393 & ~n10402;
  assign n10404 = ~pi39 & ~n10403;
  assign n10405 = n10232 & ~n10282;
  assign n10406 = ~n10279 & ~n10405;
  assign n10407 = ~n10305 & n10406;
  assign n10408 = pi39 & ~n10407;
  assign n10409 = ~n10404 & ~n10408;
  assign n10410 = n2613 & ~n10409;
  assign n10411 = ~pi87 & ~n10372;
  assign n10412 = ~n10381 & n10411;
  assign n10413 = ~n10410 & n10412;
  assign n10414 = ~pi75 & ~n10370;
  assign n10415 = ~n10413 & n10414;
  assign n10416 = n7360 & ~n10357;
  assign n10417 = ~n10415 & n10416;
  assign n10418 = ~n7360 & n10371;
  assign n10419 = ~n10101 & ~n10418;
  assign n10420 = ~n10417 & n10419;
  assign n10421 = ~pi199 & ~pi200;
  assign n10422 = ~pi299 & ~n10421;
  assign n10423 = ~pi72 & ~n10422;
  assign n10424 = ~pi232 & ~n10423;
  assign n10425 = ~pi299 & ~n10424;
  assign n10426 = n10105 & n10421;
  assign n10427 = pi232 & ~n10426;
  assign n10428 = n10425 & ~n10427;
  assign n10429 = pi39 & ~n10428;
  assign n10430 = ~n10268 & n10429;
  assign n10431 = ~n10358 & ~n10430;
  assign n10432 = ~n7360 & n10431;
  assign n10433 = ~n10355 & ~n10430;
  assign n10434 = pi75 & ~n10433;
  assign n10435 = n10369 & ~n10430;
  assign n10436 = pi38 & ~n10431;
  assign n10437 = ~n10379 & ~n10430;
  assign n10438 = n6082 & ~n10437;
  assign n10439 = pi232 & ~pi299;
  assign n10440 = ~n10169 & n10421;
  assign n10441 = n10439 & ~n10440;
  assign n10442 = ~n10279 & ~n10424;
  assign n10443 = ~n10441 & n10442;
  assign n10444 = pi39 & ~n10443;
  assign n10445 = ~n10404 & ~n10444;
  assign n10446 = n2613 & ~n10445;
  assign n10447 = ~pi87 & ~n10436;
  assign n10448 = ~n10438 & n10447;
  assign n10449 = ~n10446 & n10448;
  assign n10450 = ~pi75 & ~n10435;
  assign n10451 = ~n10449 & n10450;
  assign n10452 = n7360 & ~n10434;
  assign n10453 = ~n10451 & n10452;
  assign n10454 = n10101 & ~n10432;
  assign n10455 = ~n10453 & n10454;
  assign n10456 = ~n10420 & ~n10455;
  assign n10457 = n10336 & ~n10456;
  assign n10458 = ~n10237 & ~n10355;
  assign n10459 = pi75 & ~n10458;
  assign n10460 = ~n10237 & n10369;
  assign n10461 = ~n10237 & ~n10358;
  assign n10462 = pi38 & ~n10461;
  assign n10463 = ~n10237 & ~n10379;
  assign n10464 = n6082 & ~n10463;
  assign n10465 = n10233 & ~n10251;
  assign n10466 = pi39 & ~n10465;
  assign n10467 = ~n10404 & ~n10466;
  assign n10468 = n2613 & ~n10467;
  assign n10469 = ~pi87 & ~n10462;
  assign n10470 = ~n10464 & n10469;
  assign n10471 = ~n10468 & n10470;
  assign n10472 = ~pi75 & ~n10460;
  assign n10473 = ~n10471 & n10472;
  assign n10474 = n7360 & ~n10459;
  assign n10475 = ~n10473 & n10474;
  assign n10476 = ~n7360 & n10461;
  assign n10477 = ~n10101 & ~n10476;
  assign n10478 = ~n10475 & n10477;
  assign n10479 = ~n10358 & ~n10429;
  assign n10480 = ~n7360 & n10479;
  assign n10481 = ~n10355 & ~n10429;
  assign n10482 = pi75 & ~n10481;
  assign n10483 = ~n2532 & ~n10479;
  assign n10484 = n10369 & ~n10483;
  assign n10485 = pi38 & ~n10479;
  assign n10486 = ~n10379 & ~n10429;
  assign n10487 = n6082 & ~n10486;
  assign n10488 = pi232 & ~n10440;
  assign n10489 = n10425 & ~n10488;
  assign n10490 = pi39 & ~n10489;
  assign n10491 = ~n10404 & ~n10490;
  assign n10492 = n2613 & ~n10491;
  assign n10493 = ~pi87 & ~n10485;
  assign n10494 = ~n10487 & n10493;
  assign n10495 = ~n10492 & n10494;
  assign n10496 = ~pi75 & ~n10484;
  assign n10497 = ~n10495 & n10496;
  assign n10498 = n7360 & ~n10482;
  assign n10499 = ~n10497 & n10498;
  assign n10500 = n10101 & ~n10480;
  assign n10501 = ~n10499 & n10500;
  assign n10502 = ~n10478 & ~n10501;
  assign n10503 = ~n10336 & ~n10502;
  assign n10504 = ~po1038 & ~n10457;
  assign n10505 = ~n10503 & n10504;
  assign n10506 = n10267 & n10336;
  assign n10507 = pi39 & ~n10506;
  assign n10508 = po1038 & ~n10358;
  assign n10509 = ~n10507 & n10508;
  assign po201 = n10505 | n10509;
  assign n10511 = ~pi39 & ~n10035;
  assign n10512 = pi39 & ~pi72;
  assign n10513 = n7407 & n10512;
  assign n10514 = pi39 & ~n10513;
  assign n10515 = ~n10511 & ~n10514;
  assign n10516 = ~n2574 & n10515;
  assign n10517 = ~n7440 & ~n10035;
  assign n10518 = ~pi39 & ~n10517;
  assign n10519 = ~n2922 & n10035;
  assign n10520 = n7440 & ~n10519;
  assign n10521 = pi44 & pi72;
  assign n10522 = n7530 & ~n10521;
  assign n10523 = n7411 & n9949;
  assign n10524 = n7414 & n10523;
  assign n10525 = pi44 & ~n9960;
  assign n10526 = ~n10524 & ~n10525;
  assign n10527 = n10522 & ~n10526;
  assign n10528 = n10520 & ~n10527;
  assign n10529 = n10518 & ~n10528;
  assign n10530 = ~n10513 & ~n10529;
  assign n10531 = n2574 & ~n10530;
  assign n10532 = pi75 & ~n10516;
  assign n10533 = ~n10531 & n10532;
  assign n10534 = pi228 & n2613;
  assign n10535 = n9949 & n10534;
  assign n10536 = n9975 & n10534;
  assign n10537 = n10035 & ~n10536;
  assign n10538 = ~pi39 & ~n10535;
  assign n10539 = ~n10537 & n10538;
  assign n10540 = pi87 & ~n10514;
  assign n10541 = ~n10539 & n10540;
  assign n10542 = pi287 & n9975;
  assign n10543 = n10513 & ~n10542;
  assign n10544 = pi44 & n10039;
  assign n10545 = ~pi228 & ~n10544;
  assign n10546 = ~n10032 & n10545;
  assign n10547 = n2922 & ~n10071;
  assign n10548 = n10035 & ~n10070;
  assign n10549 = n10547 & ~n10548;
  assign n10550 = pi44 & n10051;
  assign n10551 = ~n2922 & ~n10047;
  assign n10552 = ~n10550 & n10551;
  assign n10553 = ~n10549 & ~n10552;
  assign n10554 = pi228 & ~n10553;
  assign n10555 = ~pi39 & ~n10546;
  assign n10556 = ~n10554 & n10555;
  assign n10557 = n2613 & ~n10543;
  assign n10558 = ~n10556 & n10557;
  assign n10559 = pi38 & ~n10515;
  assign n10560 = n7411 & n9975;
  assign n10561 = pi44 & ~n10560;
  assign n10562 = ~n10523 & ~n10561;
  assign n10563 = n10522 & ~n10562;
  assign n10564 = n10520 & ~n10563;
  assign n10565 = n10518 & ~n10564;
  assign n10566 = n6082 & ~n10513;
  assign n10567 = ~n10565 & n10566;
  assign n10568 = ~pi87 & ~n10559;
  assign n10569 = ~n10567 & n10568;
  assign n10570 = ~n10558 & n10569;
  assign n10571 = ~pi75 & ~n10541;
  assign n10572 = ~n10570 & n10571;
  assign n10573 = ~n10533 & ~n10572;
  assign n10574 = n7360 & ~n10573;
  assign n10575 = ~n7360 & ~n10515;
  assign n10576 = ~po1038 & ~n10575;
  assign n10577 = ~n10574 & n10576;
  assign n10578 = n2665 & n7406;
  assign n10579 = ~pi72 & n10578;
  assign n10580 = pi39 & ~n10579;
  assign n10581 = po1038 & ~n10511;
  assign n10582 = ~n10580 & n10581;
  assign po202 = n10577 | n10582;
  assign n10584 = ~pi38 & pi39;
  assign n10585 = n9830 & n10584;
  assign n10586 = pi979 & n10585;
  assign po203 = n6333 & n10586;
  assign n10588 = ~pi76 & n9874;
  assign n10589 = ~pi102 & ~pi104;
  assign n10590 = ~pi111 & n10589;
  assign n10591 = pi61 & ~pi82;
  assign n10592 = ~pi83 & ~pi89;
  assign n10593 = n10591 & n10592;
  assign n10594 = n7369 & n8634;
  assign n10595 = n10593 & n10594;
  assign n10596 = n9803 & n10590;
  assign n10597 = n10595 & n10596;
  assign n10598 = n8629 & n9877;
  assign n10599 = n10588 & n10598;
  assign n10600 = n10597 & n10599;
  assign n10601 = n8648 & n10600;
  assign n10602 = ~pi841 & n10601;
  assign n10603 = n2707 & n2889;
  assign n10604 = pi24 & n10603;
  assign n10605 = ~n10602 & ~n10604;
  assign po204 = n9782 & ~n10605;
  assign n10607 = ~pi82 & n2473;
  assign n10608 = ~pi84 & pi104;
  assign n10609 = n2804 & n10608;
  assign n10610 = n9802 & n10609;
  assign n10611 = n10607 & n10610;
  assign n10612 = ~pi36 & ~n10611;
  assign n10613 = n8635 & n8773;
  assign n10614 = n2485 & n2489;
  assign n10615 = ~pi98 & n10614;
  assign n10616 = n10613 & n10615;
  assign n10617 = ~n10612 & n10616;
  assign n10618 = ~n2802 & n10617;
  assign n10619 = ~pi88 & ~n10618;
  assign n10620 = ~n2871 & n7369;
  assign n10621 = n2754 & ~n10619;
  assign n10622 = n10620 & n10621;
  assign n10623 = n2705 & n10622;
  assign n10624 = ~n9797 & ~n10623;
  assign n10625 = n9778 & ~n10624;
  assign n10626 = n7425 & ~n10625;
  assign n10627 = ~pi36 & n10617;
  assign n10628 = ~pi88 & ~n10627;
  assign n10629 = n10620 & ~n10628;
  assign n10630 = n9816 & n10629;
  assign n10631 = ~pi824 & n6102;
  assign n10632 = n10630 & n10631;
  assign n10633 = ~n6102 & n10625;
  assign n10634 = pi829 & ~n10632;
  assign n10635 = ~n10633 & n10634;
  assign n10636 = ~n2921 & n10635;
  assign n10637 = ~n10626 & ~n10636;
  assign n10638 = pi1091 & ~n10637;
  assign n10639 = ~n7348 & n10625;
  assign n10640 = ~pi829 & ~n10639;
  assign n10641 = ~n10635 & ~n10640;
  assign n10642 = ~pi1093 & ~n10641;
  assign n10643 = n2711 & n7348;
  assign n10644 = n3174 & n10643;
  assign n10645 = ~n9798 & n10644;
  assign n10646 = ~n6339 & ~n7561;
  assign n10647 = ~n10645 & ~n10646;
  assign n10648 = ~n10639 & n10647;
  assign n10649 = n9781 & ~n10648;
  assign n10650 = ~n10642 & n10649;
  assign po205 = ~n10638 & n10650;
  assign n10652 = pi841 & n2520;
  assign n10653 = n9781 & n10652;
  assign n10654 = n9886 & n10653;
  assign po206 = n9815 & n10654;
  assign n10656 = n2518 & n2735;
  assign n10657 = ~pi70 & n10656;
  assign n10658 = ~pi35 & ~pi51;
  assign n10659 = ~pi103 & n2803;
  assign n10660 = n9875 & n10659;
  assign n10661 = n8633 & n8635;
  assign n10662 = n10660 & n10661;
  assign n10663 = n2466 & n2489;
  assign n10664 = ~pi45 & pi49;
  assign n10665 = n10590 & n10664;
  assign n10666 = n10662 & n10665;
  assign n10667 = n10663 & n10666;
  assign n10668 = n10607 & n10667;
  assign n10669 = n8648 & n10658;
  assign n10670 = n10668 & n10669;
  assign n10671 = pi841 & n2709;
  assign n10672 = n10657 & n10671;
  assign n10673 = n10670 & n10672;
  assign n10674 = ~pi74 & ~n10673;
  assign n10675 = pi74 & ~n7413;
  assign n10676 = n9780 & ~n10674;
  assign po207 = ~n10675 & n10676;
  assign n10678 = pi24 & ~pi94;
  assign n10679 = ~n8613 & n10678;
  assign n10680 = pi24 & n8611;
  assign n10681 = ~n10013 & ~n10680;
  assign n10682 = pi252 & ~po840;
  assign n10683 = ~pi252 & ~n8600;
  assign n10684 = ~n10682 & ~n10683;
  assign n10685 = n9778 & n10684;
  assign n10686 = ~n10679 & n10685;
  assign n10687 = ~n10681 & n10686;
  assign n10688 = n2509 & n10656;
  assign n10689 = pi24 & ~pi90;
  assign n10690 = n10688 & n10689;
  assign n10691 = ~n10684 & n10690;
  assign n10692 = n8615 & n10691;
  assign n10693 = ~n10687 & ~n10692;
  assign n10694 = ~pi100 & ~n10693;
  assign n10695 = pi100 & n8672;
  assign n10696 = n6311 & n10695;
  assign n10697 = ~n10694 & ~n10696;
  assign n10698 = n2531 & n2534;
  assign n10699 = ~n10697 & n10698;
  assign n10700 = n8671 & n8672;
  assign n10701 = n8668 & n10700;
  assign n10702 = ~n10699 & ~n10701;
  assign po208 = n8598 & ~n10702;
  assign n10704 = n2705 & n9782;
  assign n10705 = n2754 & n10704;
  assign n10706 = n2489 & n8775;
  assign n10707 = n9878 & n10706;
  assign n10708 = ~pi69 & n10707;
  assign n10709 = n2803 & n10708;
  assign n10710 = n10705 & n10709;
  assign po209 = n2806 & n10710;
  assign n10712 = pi52 & ~pi72;
  assign n10713 = ~pi39 & ~n10712;
  assign n10714 = ~n10429 & ~n10713;
  assign n10715 = ~n7360 & ~n10101;
  assign n10716 = n10714 & n10715;
  assign n10717 = ~n10269 & ~n10713;
  assign n10718 = ~n7360 & n10717;
  assign n10719 = ~pi219 & n10335;
  assign n10720 = ~n2613 & n10717;
  assign n10721 = pi87 & ~n10720;
  assign n10722 = ~pi52 & n10123;
  assign n10723 = pi52 & n10156;
  assign n10724 = ~n10722 & ~n10723;
  assign n10725 = n10361 & ~n10724;
  assign n10726 = ~n10361 & n10712;
  assign n10727 = ~n10725 & ~n10726;
  assign n10728 = ~pi39 & n10727;
  assign n10729 = n2613 & ~n10269;
  assign n10730 = ~n10728 & n10729;
  assign n10731 = n10721 & ~n10730;
  assign n10732 = pi38 & ~n10717;
  assign n10733 = n2922 & n7440;
  assign n10734 = n10360 & n10733;
  assign n10735 = n7411 & n10155;
  assign n10736 = n10734 & n10735;
  assign n10737 = n10712 & ~n10736;
  assign n10738 = ~pi39 & ~n10737;
  assign n10739 = ~n10269 & ~n10738;
  assign n10740 = n6082 & ~n10739;
  assign n10741 = ~n10279 & n10282;
  assign n10742 = pi39 & ~n10741;
  assign n10743 = ~n10360 & ~n10712;
  assign n10744 = ~pi52 & n10176;
  assign n10745 = pi52 & ~n10184;
  assign n10746 = n10360 & ~n10744;
  assign n10747 = ~n10745 & n10746;
  assign n10748 = ~pi228 & ~n10743;
  assign n10749 = ~n10747 & n10748;
  assign n10750 = ~pi52 & n10388;
  assign n10751 = pi52 & n10397;
  assign n10752 = n10360 & ~n10750;
  assign n10753 = ~n10751 & n10752;
  assign n10754 = pi228 & ~n10743;
  assign n10755 = ~n10753 & n10754;
  assign n10756 = ~pi39 & ~n10749;
  assign n10757 = ~n10755 & n10756;
  assign n10758 = ~n10742 & ~n10757;
  assign n10759 = n2613 & ~n10758;
  assign n10760 = ~n10732 & ~n10740;
  assign n10761 = ~n10759 & n10760;
  assign n10762 = ~pi87 & ~n10761;
  assign n10763 = n10101 & ~n10731;
  assign n10764 = ~n10762 & n10763;
  assign n10765 = ~n2613 & n10714;
  assign n10766 = n2613 & ~n10430;
  assign n10767 = ~n10728 & n10766;
  assign n10768 = n10721 & ~n10765;
  assign n10769 = ~n10767 & n10768;
  assign n10770 = pi38 & ~n10714;
  assign n10771 = ~n10717 & n10770;
  assign n10772 = ~n10444 & ~n10757;
  assign n10773 = n2613 & ~n10772;
  assign n10774 = ~n10430 & ~n10738;
  assign n10775 = n6082 & ~n10774;
  assign n10776 = ~n10771 & ~n10775;
  assign n10777 = ~n10773 & n10776;
  assign n10778 = ~pi87 & ~n10777;
  assign n10779 = ~n10101 & ~n10769;
  assign n10780 = ~n10778 & n10779;
  assign n10781 = ~n10764 & ~n10780;
  assign n10782 = ~pi75 & ~n10781;
  assign n10783 = ~pi39 & n10712;
  assign n10784 = n2574 & n10734;
  assign n10785 = n10120 & n10784;
  assign n10786 = n10783 & ~n10785;
  assign n10787 = ~pi39 & ~n10786;
  assign n10788 = ~n10101 & n10428;
  assign n10789 = n10269 & ~n10788;
  assign n10790 = pi75 & ~n10789;
  assign n10791 = ~n10787 & n10790;
  assign n10792 = ~n10782 & ~n10791;
  assign n10793 = n7360 & ~n10792;
  assign n10794 = ~n10718 & n10719;
  assign n10795 = ~n10793 & n10794;
  assign n10796 = n2613 & ~n10429;
  assign n10797 = ~n10728 & n10796;
  assign n10798 = ~n10765 & ~n10797;
  assign n10799 = pi87 & ~n10798;
  assign n10800 = ~n10429 & ~n10738;
  assign n10801 = n6082 & ~n10800;
  assign n10802 = ~n10490 & ~n10757;
  assign n10803 = n2613 & ~n10802;
  assign n10804 = ~pi87 & ~n10770;
  assign n10805 = ~n10801 & n10804;
  assign n10806 = ~n10803 & n10805;
  assign n10807 = ~pi75 & ~n10799;
  assign n10808 = ~n10806 & n10807;
  assign n10809 = ~n10429 & ~n10787;
  assign n10810 = pi75 & ~n10809;
  assign n10811 = n7360 & ~n10101;
  assign n10812 = ~n10810 & n10811;
  assign n10813 = ~n10808 & n10812;
  assign n10814 = ~n7360 & ~n10783;
  assign n10815 = pi75 & n10786;
  assign n10816 = pi100 & ~n10783;
  assign n10817 = pi38 & ~n10783;
  assign n10818 = ~pi38 & n10727;
  assign n10819 = ~n10817 & ~n10818;
  assign n10820 = ~pi100 & ~n10819;
  assign n10821 = ~pi100 & n10584;
  assign n10822 = pi87 & ~n10821;
  assign n10823 = ~n10816 & n10822;
  assign n10824 = ~n10820 & n10823;
  assign n10825 = pi100 & ~n10737;
  assign n10826 = ~pi100 & n10757;
  assign n10827 = ~pi39 & ~n10825;
  assign n10828 = ~n10826 & n10827;
  assign n10829 = ~pi38 & ~n10828;
  assign n10830 = ~pi87 & ~n10817;
  assign n10831 = ~n10829 & n10830;
  assign n10832 = ~n10824 & ~n10831;
  assign n10833 = ~pi75 & ~n10832;
  assign n10834 = n7360 & ~n10815;
  assign n10835 = ~n10833 & n10834;
  assign n10836 = n10101 & ~n10814;
  assign n10837 = ~n10835 & n10836;
  assign n10838 = ~n10719 & ~n10813;
  assign n10839 = ~n10837 & n10838;
  assign n10840 = ~n10795 & ~n10839;
  assign n10841 = ~po1038 & ~n10716;
  assign n10842 = ~n10840 & n10841;
  assign n10843 = pi39 & n10719;
  assign n10844 = n10267 & n10843;
  assign n10845 = po1038 & ~n10783;
  assign n10846 = ~n10844 & n10845;
  assign po210 = ~n10842 & ~n10846;
  assign n10848 = ~pi287 & ~pi979;
  assign n10849 = n6167 & n10848;
  assign n10850 = pi39 & ~n10849;
  assign n10851 = pi24 & n9778;
  assign n10852 = pi53 & n2720;
  assign n10853 = n2717 & n10852;
  assign n10854 = n2721 & n10853;
  assign n10855 = n10851 & n10854;
  assign n10856 = ~pi39 & ~n10855;
  assign n10857 = n9833 & ~n10850;
  assign n10858 = ~n10856 & n10857;
  assign po211 = ~n3378 & n10858;
  assign n10860 = n8611 & n8944;
  assign n10861 = ~pi60 & ~pi85;
  assign n10862 = pi106 & n10861;
  assign n10863 = n2478 & n8631;
  assign n10864 = n10862 & n10863;
  assign n10865 = n8638 & n10864;
  assign n10866 = n10588 & n10660;
  assign n10867 = n10865 & n10866;
  assign n10868 = n10663 & n10867;
  assign n10869 = n10860 & n10868;
  assign n10870 = ~pi841 & n2709;
  assign n10871 = n10657 & n10870;
  assign n10872 = n2616 & n10658;
  assign n10873 = n10871 & n10872;
  assign n10874 = n10869 & n10873;
  assign n10875 = ~pi54 & ~n10874;
  assign n10876 = n2575 & n9827;
  assign n10877 = pi54 & ~n10876;
  assign n10878 = n8597 & ~n10875;
  assign po212 = ~n10877 & n10878;
  assign n10880 = n2577 & n9778;
  assign n10881 = n2467 & n8648;
  assign n10882 = n10880 & n10881;
  assign n10883 = pi45 & n2478;
  assign n10884 = n2489 & n10883;
  assign n10885 = n10662 & n10884;
  assign n10886 = n2475 & n10885;
  assign n10887 = n10882 & n10886;
  assign n10888 = ~pi55 & ~n10887;
  assign n10889 = n2576 & n9827;
  assign n10890 = pi55 & ~n10889;
  assign n10891 = n2530 & n3291;
  assign n10892 = ~n10888 & n10891;
  assign po213 = ~n10890 & n10892;
  assign n10894 = n2518 & n2538;
  assign n10895 = n2917 & n10894;
  assign n10896 = pi56 & ~n10895;
  assign n10897 = pi56 & ~pi62;
  assign n10898 = pi55 & n9705;
  assign n10899 = ~n10897 & ~n10898;
  assign n10900 = n3291 & ~n10896;
  assign po214 = ~n10899 & n10900;
  assign n10902 = n6257 & n10889;
  assign n10903 = pi57 & ~n10902;
  assign n10904 = n6437 & n10894;
  assign n10905 = ~pi56 & pi62;
  assign n10906 = ~pi924 & n10905;
  assign n10907 = ~n10897 & ~n10906;
  assign n10908 = n10904 & ~n10907;
  assign n10909 = ~pi57 & ~n10908;
  assign n10910 = ~pi59 & ~n10903;
  assign po215 = ~n10909 & n10910;
  assign n10912 = n9781 & n10688;
  assign n10913 = ~pi93 & n10912;
  assign po216 = n7364 & n10913;
  assign n10915 = pi59 & ~n10902;
  assign n10916 = pi924 & n10905;
  assign n10917 = n10904 & n10916;
  assign n10918 = ~pi59 & ~n10917;
  assign n10919 = ~pi57 & ~n10915;
  assign po217 = ~n10918 & n10919;
  assign n10921 = pi39 & ~pi979;
  assign n10922 = ~n6167 & n10921;
  assign n10923 = n6168 & n10922;
  assign n10924 = n6333 & n10923;
  assign n10925 = ~pi39 & n10851;
  assign n10926 = n10860 & n10925;
  assign n10927 = n2718 & n10926;
  assign n10928 = ~n10924 & ~n10927;
  assign po218 = n9833 & ~n10928;
  assign n10930 = pi841 & n10601;
  assign n10931 = ~pi24 & n10860;
  assign n10932 = n2718 & n10931;
  assign n10933 = ~n10930 & ~n10932;
  assign po219 = n9782 & ~n10933;
  assign n10935 = n10895 & n10905;
  assign n10936 = ~pi57 & ~n10935;
  assign n10937 = pi57 & ~n9706;
  assign n10938 = ~pi59 & ~n10936;
  assign po220 = ~n10937 & n10938;
  assign n10940 = n8625 & n10881;
  assign n10941 = n2862 & n10940;
  assign n10942 = pi999 & n10941;
  assign n10943 = ~pi24 & n10603;
  assign n10944 = ~n10942 & ~n10943;
  assign po221 = n9782 & ~n10944;
  assign n10946 = n2849 & n8814;
  assign n10947 = ~pi841 & ~n10946;
  assign n10948 = ~pi64 & ~n2850;
  assign n10949 = n2467 & ~n10948;
  assign n10950 = n9813 & n10949;
  assign n10951 = pi841 & ~n10950;
  assign n10952 = n10705 & ~n10947;
  assign po222 = ~n10951 & n10952;
  assign n10954 = n9857 & n10585;
  assign n10955 = ~n9849 & n10954;
  assign po223 = ~n9855 & n10955;
  assign n10957 = pi199 & ~pi299;
  assign n10958 = n2613 & n7293;
  assign n10959 = n8623 & n8648;
  assign n10960 = n6431 & n10959;
  assign n10961 = pi314 & n2466;
  assign n10962 = n10960 & n10961;
  assign n10963 = pi81 & ~pi102;
  assign n10964 = n10962 & n10963;
  assign n10965 = n2491 & n10964;
  assign n10966 = n2614 & n10957;
  assign n10967 = n10958 & n10966;
  assign n10968 = n10965 & n10967;
  assign n10969 = ~pi219 & ~n10968;
  assign n10970 = ~pi199 & ~pi299;
  assign n10971 = n2577 & n10965;
  assign n10972 = ~n10970 & n10971;
  assign n10973 = pi219 & ~n10972;
  assign n10974 = ~po1038 & ~n10969;
  assign po224 = ~n10973 & n10974;
  assign n10976 = pi83 & ~pi103;
  assign n10977 = n10706 & n10976;
  assign n10978 = n9781 & n10977;
  assign n10979 = n10962 & n10978;
  assign po225 = n2793 & n10979;
  assign n10981 = ~n6223 & n6341;
  assign n10982 = n3293 & n5966;
  assign n10983 = n10981 & n10982;
  assign n10984 = ~n6207 & n6341;
  assign n10985 = n3328 & n5783;
  assign n10986 = n10984 & n10985;
  assign n10987 = ~n10983 & ~n10986;
  assign po226 = n10585 & ~n10987;
  assign n10989 = pi69 & n10659;
  assign n10990 = n9791 & n10989;
  assign n10991 = ~pi71 & ~n10990;
  assign n10992 = ~pi81 & ~pi314;
  assign n10993 = n2467 & n10992;
  assign n10994 = n6389 & n10993;
  assign n10995 = ~n10991 & n10994;
  assign n10996 = pi71 & pi314;
  assign n10997 = n7369 & n10996;
  assign n10998 = n9788 & n10997;
  assign n10999 = n2487 & n10998;
  assign n11000 = ~n10995 & ~n10999;
  assign po227 = n10705 & ~n11000;
  assign n11002 = n2517 & n2749;
  assign n11003 = ~pi96 & n11002;
  assign n11004 = n2701 & n11003;
  assign n11005 = pi24 & n9824;
  assign n11006 = n11004 & n11005;
  assign n11007 = ~n7255 & ~n7257;
  assign n11008 = n2608 & n5783;
  assign n11009 = pi299 & n3303;
  assign n11010 = ~n11008 & ~n11009;
  assign n11011 = ~n11007 & ~n11010;
  assign n11012 = pi210 & pi589;
  assign n11013 = n3303 & ~n11012;
  assign n11014 = n7257 & n11013;
  assign n11015 = pi198 & pi589;
  assign n11016 = n2608 & ~n11015;
  assign n11017 = n9861 & n11016;
  assign n11018 = ~n11014 & ~n11017;
  assign n11019 = ~pi593 & n6334;
  assign n11020 = ~n6346 & n11019;
  assign n11021 = n11011 & n11020;
  assign n11022 = n11018 & n11021;
  assign n11023 = ~pi287 & ~n11022;
  assign n11024 = pi39 & ~n11023;
  assign n11025 = n2523 & n11024;
  assign n11026 = ~n11006 & ~n11025;
  assign po228 = n9833 & ~n11026;
  assign n11028 = n2482 & n6374;
  assign n11029 = n10614 & n11028;
  assign n11030 = ~pi64 & n8635;
  assign n11031 = n11029 & n11030;
  assign n11032 = ~pi81 & ~n11031;
  assign n11033 = ~pi50 & n8648;
  assign n11034 = n6393 & n11033;
  assign n11035 = ~pi199 & pi200;
  assign n11036 = ~pi299 & n11035;
  assign n11037 = pi211 & ~pi219;
  assign n11038 = pi299 & n11037;
  assign n11039 = ~n11036 & ~n11038;
  assign n11040 = pi314 & ~n11039;
  assign n11041 = n9778 & n11040;
  assign n11042 = ~n11032 & n11041;
  assign n11043 = n11034 & n11042;
  assign n11044 = n10613 & n11039;
  assign n11045 = n10962 & n11044;
  assign n11046 = n11029 & n11045;
  assign n11047 = ~n11043 & ~n11046;
  assign po229 = n9781 & ~n11047;
  assign n11049 = pi72 & n9825;
  assign n11050 = pi88 & n9785;
  assign n11051 = n2870 & n11050;
  assign n11052 = n6345 & n8623;
  assign n11053 = n11051 & n11052;
  assign n11054 = ~n11049 & ~n11053;
  assign n11055 = n6431 & ~n11054;
  assign n11056 = ~pi39 & ~n11055;
  assign n11057 = n7544 & n10981;
  assign n11058 = n7548 & n10984;
  assign n11059 = pi39 & ~n11057;
  assign n11060 = ~n11058 & n11059;
  assign n11061 = n9833 & ~n11060;
  assign po230 = ~n11056 & n11061;
  assign n11063 = n8752 & n10984;
  assign n11064 = ~pi299 & ~n11063;
  assign n11065 = n8739 & n10981;
  assign n11066 = pi299 & ~n11065;
  assign n11067 = ~n11064 & ~n11066;
  assign n11068 = pi39 & n11067;
  assign n11069 = ~pi314 & pi1050;
  assign n11070 = n6431 & n8783;
  assign n11071 = ~pi39 & n11069;
  assign n11072 = n11070 & n11071;
  assign n11073 = ~n11068 & ~n11072;
  assign po231 = n9833 & ~n11073;
  assign n11075 = n2955 & n7461;
  assign n11076 = ~pi96 & ~n11075;
  assign n11077 = ~pi96 & n6150;
  assign n11078 = pi479 & ~n11077;
  assign n11079 = ~pi96 & ~pi1093;
  assign n11080 = n7348 & n11079;
  assign n11081 = n3353 & n7360;
  assign n11082 = ~n11080 & n11081;
  assign n11083 = ~po840 & ~n11078;
  assign n11084 = n11082 & n11083;
  assign n11085 = n7389 & n11084;
  assign n11086 = ~n11076 & n11085;
  assign n11087 = n2574 & n9827;
  assign n11088 = pi74 & n6276;
  assign n11089 = n11087 & n11088;
  assign n11090 = ~n11086 & ~n11089;
  assign po232 = ~po1038 & ~n11090;
  assign n11092 = pi75 & ~n11087;
  assign n11093 = n2615 & ~n11079;
  assign n11094 = ~n6175 & n11093;
  assign n11095 = ~n11076 & n11094;
  assign n11096 = n7471 & n11095;
  assign n11097 = ~pi75 & ~n11096;
  assign n11098 = n8598 & ~n11092;
  assign po233 = ~n11097 & n11098;
  assign n11100 = n8646 & n9816;
  assign n11101 = ~n9739 & n11100;
  assign n11102 = po1057 & ~n11101;
  assign n11103 = n3174 & n10014;
  assign n11104 = pi829 & n6102;
  assign n11105 = pi252 & n11104;
  assign n11106 = n11103 & ~n11105;
  assign n11107 = ~pi137 & n11106;
  assign n11108 = ~pi137 & n2922;
  assign n11109 = ~n8611 & ~n10013;
  assign n11110 = ~pi94 & ~n9741;
  assign n11111 = n9778 & ~n11110;
  assign n11112 = ~n11109 & n11111;
  assign n11113 = ~n11104 & ~n11112;
  assign n11114 = ~pi252 & n11112;
  assign n11115 = pi252 & n11100;
  assign n11116 = n11104 & ~n11115;
  assign n11117 = ~n11114 & n11116;
  assign n11118 = ~n11113 & ~n11117;
  assign n11119 = pi122 & ~n11118;
  assign n11120 = n7348 & n11113;
  assign n11121 = ~n6104 & ~n11103;
  assign n11122 = ~n11117 & ~n11121;
  assign n11123 = ~n11120 & n11122;
  assign n11124 = ~pi122 & ~n11123;
  assign n11125 = ~n11119 & ~n11124;
  assign n11126 = ~pi1093 & ~n11125;
  assign n11127 = ~pi122 & ~n11106;
  assign n11128 = ~n11119 & ~n11127;
  assign n11129 = pi1093 & ~n11128;
  assign n11130 = ~n11126 & ~n11129;
  assign n11131 = n2922 & ~n11130;
  assign n11132 = ~n11108 & ~n11131;
  assign n11133 = ~n11107 & ~n11132;
  assign n11134 = ~pi122 & n11103;
  assign n11135 = pi1093 & ~n11112;
  assign n11136 = ~n7349 & ~n11135;
  assign n11137 = ~n11134 & ~n11136;
  assign n11138 = ~n11126 & ~n11137;
  assign n11139 = ~n2922 & ~n11138;
  assign n11140 = ~pi137 & ~n2922;
  assign n11141 = ~n11139 & ~n11140;
  assign n11142 = pi252 & pi1092;
  assign n11143 = ~pi1093 & n11142;
  assign n11144 = n2924 & n11143;
  assign n11145 = ~pi137 & ~n11144;
  assign n11146 = n11103 & n11145;
  assign n11147 = ~n11141 & ~n11146;
  assign n11148 = ~n11133 & ~n11147;
  assign n11149 = ~po1057 & ~n11148;
  assign n11150 = ~pi137 & po1057;
  assign n11151 = ~n11102 & ~n11150;
  assign n11152 = ~n11149 & n11151;
  assign n11153 = ~pi210 & ~n11152;
  assign n11154 = ~n11131 & ~n11139;
  assign n11155 = ~po1057 & ~n11154;
  assign n11156 = ~n11102 & ~n11155;
  assign n11157 = pi210 & ~n11156;
  assign n11158 = ~n11153 & ~n11157;
  assign n11159 = n2664 & n9931;
  assign n11160 = ~n11158 & ~n11159;
  assign n11161 = pi210 & ~n11154;
  assign n11162 = ~pi210 & ~n11148;
  assign n11163 = ~n11161 & ~n11162;
  assign n11164 = n11159 & ~n11163;
  assign n11165 = pi299 & ~n11164;
  assign n11166 = ~n11160 & n11165;
  assign n11167 = ~pi198 & ~n11152;
  assign n11168 = pi198 & ~n11156;
  assign n11169 = ~n11167 & ~n11168;
  assign n11170 = n2641 & n6166;
  assign n11171 = ~n11169 & ~n11170;
  assign n11172 = pi198 & ~n11154;
  assign n11173 = ~pi198 & ~n11148;
  assign n11174 = ~n11172 & ~n11173;
  assign n11175 = n11170 & ~n11174;
  assign n11176 = ~pi299 & ~n11175;
  assign n11177 = ~n11171 & n11176;
  assign n11178 = ~n11166 & ~n11177;
  assign n11179 = pi232 & ~n11178;
  assign n11180 = pi299 & ~n11158;
  assign n11181 = ~pi299 & ~n11169;
  assign n11182 = ~pi232 & ~n11180;
  assign n11183 = ~n11181 & n11182;
  assign n11184 = ~n11179 & ~n11183;
  assign n11185 = n7356 & ~n11184;
  assign n11186 = ~n2922 & n11135;
  assign n11187 = ~n11103 & n11104;
  assign n11188 = ~n11105 & ~n11113;
  assign n11189 = ~n11187 & n11188;
  assign n11190 = n7349 & ~n11189;
  assign n11191 = ~n11119 & ~n11190;
  assign n11192 = n2922 & ~n11191;
  assign n11193 = ~pi1093 & ~n11118;
  assign n11194 = ~n11186 & ~n11193;
  assign n11195 = ~n11192 & n11194;
  assign n11196 = ~po1057 & n11195;
  assign n11197 = po1057 & n11100;
  assign n11198 = ~n9737 & n11197;
  assign n11199 = ~n11196 & ~n11198;
  assign n11200 = pi210 & ~n11199;
  assign n11201 = n8618 & n11150;
  assign n11202 = ~pi137 & ~n11189;
  assign n11203 = pi137 & n11193;
  assign n11204 = ~n11202 & ~n11203;
  assign n11205 = ~pi1093 & ~n11204;
  assign n11206 = ~po1057 & ~n11135;
  assign n11207 = ~n11205 & n11206;
  assign n11208 = ~n11197 & ~n11207;
  assign n11209 = ~n2922 & ~n11201;
  assign n11210 = ~n11208 & n11209;
  assign n11211 = pi137 & ~n7349;
  assign n11212 = n11104 & ~n11211;
  assign n11213 = n11100 & ~n11212;
  assign n11214 = po1057 & ~n11213;
  assign n11215 = pi137 & ~n11191;
  assign n11216 = n11204 & ~n11215;
  assign n11217 = ~po1057 & ~n11216;
  assign n11218 = n2922 & ~n11214;
  assign n11219 = ~n11217 & n11218;
  assign n11220 = ~n11210 & ~n11219;
  assign n11221 = ~pi210 & ~n11220;
  assign n11222 = ~n11200 & ~n11221;
  assign n11223 = ~n11159 & ~n11222;
  assign n11224 = ~n6175 & ~n11216;
  assign n11225 = ~n11186 & ~n11224;
  assign n11226 = ~pi210 & n11225;
  assign n11227 = pi210 & n11195;
  assign n11228 = ~n11226 & ~n11227;
  assign n11229 = n11159 & ~n11228;
  assign n11230 = pi299 & ~n11229;
  assign n11231 = ~n11223 & n11230;
  assign n11232 = pi198 & ~n11199;
  assign n11233 = ~pi198 & ~n11220;
  assign n11234 = ~n11232 & ~n11233;
  assign n11235 = ~n11170 & ~n11234;
  assign n11236 = ~pi198 & ~n11225;
  assign n11237 = pi198 & ~n11195;
  assign n11238 = n11170 & ~n11237;
  assign n11239 = ~n11236 & n11238;
  assign n11240 = ~pi299 & ~n11239;
  assign n11241 = ~n11235 & n11240;
  assign n11242 = ~n11231 & ~n11241;
  assign n11243 = pi232 & ~n11242;
  assign n11244 = pi299 & ~n11222;
  assign n11245 = ~pi299 & ~n11234;
  assign n11246 = ~pi232 & ~n11244;
  assign n11247 = ~n11245 & n11246;
  assign n11248 = ~n7356 & ~n11247;
  assign n11249 = ~n11243 & n11248;
  assign n11250 = ~n11185 & ~n11249;
  assign po234 = n9781 & ~n11250;
  assign n11252 = n2767 & n2782;
  assign n11253 = ~pi86 & ~n11252;
  assign n11254 = n6400 & ~n11253;
  assign n11255 = n2707 & n11254;
  assign n11256 = ~pi314 & n11255;
  assign n11257 = pi86 & n8611;
  assign n11258 = pi314 & n11257;
  assign n11259 = n2770 & n11258;
  assign n11260 = ~n11256 & ~n11259;
  assign po235 = n9782 & ~n11260;
  assign n11262 = pi119 & pi232;
  assign po236 = ~pi468 & n11262;
  assign n11264 = pi163 & ~n9363;
  assign n11265 = ~pi163 & ~n9359;
  assign n11266 = ~n9361 & n11265;
  assign n11267 = ~n11264 & ~n11266;
  assign n11268 = pi232 & n11267;
  assign n11269 = ~n7231 & n11268;
  assign n11270 = pi74 & ~n11269;
  assign n11271 = pi75 & ~n11268;
  assign n11272 = pi100 & ~n11268;
  assign n11273 = ~n11271 & ~n11272;
  assign n11274 = pi147 & n7406;
  assign n11275 = n7231 & n11274;
  assign n11276 = n11273 & ~n11275;
  assign n11277 = ~n3291 & ~n11270;
  assign n11278 = n11276 & n11277;
  assign n11279 = pi54 & ~n11276;
  assign n11280 = ~pi38 & ~pi40;
  assign n11281 = pi38 & ~n11274;
  assign n11282 = ~pi100 & ~n11281;
  assign n11283 = ~n11280 & n11282;
  assign n11284 = ~n11272 & ~n11283;
  assign n11285 = ~pi75 & ~n11284;
  assign n11286 = ~n11271 & ~n11285;
  assign n11287 = ~pi54 & ~n11286;
  assign n11288 = ~n11279 & ~n11287;
  assign n11289 = ~pi74 & ~n11288;
  assign n11290 = ~n11270 & ~n11289;
  assign n11291 = ~n2530 & ~n11290;
  assign n11292 = n3291 & ~n11291;
  assign n11293 = ~n9384 & n9386;
  assign n11294 = ~pi184 & n11293;
  assign n11295 = pi184 & n6166;
  assign n11296 = ~n11293 & n11295;
  assign n11297 = ~pi299 & ~n11294;
  assign n11298 = ~n11296 & n11297;
  assign n11299 = pi299 & ~n11267;
  assign n11300 = pi232 & ~n11298;
  assign n11301 = ~n11299 & n11300;
  assign n11302 = ~n7231 & n11301;
  assign n11303 = pi74 & ~n11302;
  assign n11304 = ~pi55 & ~n11303;
  assign n11305 = ~pi187 & ~pi299;
  assign n11306 = ~pi147 & pi299;
  assign n11307 = ~n11305 & ~n11306;
  assign n11308 = n7406 & n11307;
  assign n11309 = n7231 & ~n11308;
  assign n11310 = pi54 & ~n11309;
  assign n11311 = ~n11302 & n11310;
  assign n11312 = pi75 & ~n11301;
  assign n11313 = pi100 & ~n11301;
  assign n11314 = pi38 & ~n11308;
  assign n11315 = ~pi100 & ~n11314;
  assign n11316 = ~pi179 & ~pi299;
  assign n11317 = ~pi156 & pi299;
  assign n11318 = ~n11316 & ~n11317;
  assign n11319 = n7406 & n11318;
  assign n11320 = n2518 & n2614;
  assign n11321 = n11319 & n11320;
  assign n11322 = n2511 & n11321;
  assign n11323 = n11280 & ~n11322;
  assign n11324 = n11315 & ~n11323;
  assign n11325 = ~n11313 & ~n11324;
  assign n11326 = n8890 & ~n11325;
  assign n11327 = ~pi187 & ~n8872;
  assign n11328 = pi187 & ~n8874;
  assign n11329 = pi147 & ~n11328;
  assign n11330 = ~n11327 & n11329;
  assign n11331 = ~pi147 & pi187;
  assign n11332 = n8879 & n11331;
  assign n11333 = ~n11330 & ~n11332;
  assign n11334 = pi38 & ~n11333;
  assign n11335 = n2511 & n8787;
  assign n11336 = pi156 & n6203;
  assign n11337 = ~pi166 & n8981;
  assign n11338 = ~n11336 & ~n11337;
  assign n11339 = ~n6221 & n8739;
  assign n11340 = ~n11338 & n11339;
  assign n11341 = n11335 & n11340;
  assign n11342 = ~pi40 & pi299;
  assign n11343 = ~n11341 & n11342;
  assign n11344 = ~pi189 & n8981;
  assign n11345 = pi179 & n6203;
  assign n11346 = ~n11344 & ~n11345;
  assign n11347 = n8753 & ~n11346;
  assign n11348 = n11335 & n11347;
  assign n11349 = ~pi40 & ~pi299;
  assign n11350 = ~n11348 & n11349;
  assign n11351 = pi39 & ~n11343;
  assign n11352 = ~n11350 & n11351;
  assign n11353 = pi40 & ~pi299;
  assign n11354 = ~pi182 & pi184;
  assign n11355 = ~pi32 & pi95;
  assign n11356 = ~pi479 & n11355;
  assign n11357 = n2511 & n11356;
  assign n11358 = pi182 & n11357;
  assign n11359 = ~pi189 & n8783;
  assign n11360 = ~n8793 & ~n11359;
  assign n11361 = n2518 & ~n11360;
  assign n11362 = ~pi184 & ~n11358;
  assign n11363 = ~n11361 & n11362;
  assign n11364 = ~pi189 & n8826;
  assign n11365 = pi189 & n8808;
  assign n11366 = ~n6471 & ~n11365;
  assign n11367 = ~n11364 & n11366;
  assign n11368 = pi184 & ~n11357;
  assign n11369 = n11367 & n11368;
  assign n11370 = n6166 & ~n11363;
  assign n11371 = ~n11369 & n11370;
  assign n11372 = ~n11354 & ~n11371;
  assign n11373 = pi175 & ~pi299;
  assign n11374 = n6166 & ~n11367;
  assign n11375 = n11354 & ~n11374;
  assign n11376 = n11373 & ~n11375;
  assign n11377 = ~n11372 & n11376;
  assign n11378 = n6166 & n11357;
  assign n11379 = pi153 & n8787;
  assign n11380 = n8793 & n11379;
  assign n11381 = n8784 & n9931;
  assign n11382 = ~pi40 & ~pi163;
  assign n11383 = ~n11381 & n11382;
  assign n11384 = ~n11380 & n11383;
  assign n11385 = ~n11378 & n11384;
  assign n11386 = pi166 & n6166;
  assign n11387 = pi153 & n8808;
  assign n11388 = n8811 & ~n11387;
  assign n11389 = n11386 & ~n11388;
  assign n11390 = pi153 & n8826;
  assign n11391 = n8829 & ~n11390;
  assign n11392 = n9931 & ~n11391;
  assign n11393 = ~pi40 & pi163;
  assign n11394 = ~n11389 & n11393;
  assign n11395 = ~n11392 & n11394;
  assign n11396 = ~n11378 & n11395;
  assign n11397 = pi160 & ~n11396;
  assign n11398 = ~n11384 & ~n11395;
  assign n11399 = ~n11397 & ~n11398;
  assign n11400 = pi299 & ~n11385;
  assign n11401 = ~n11399 & n11400;
  assign n11402 = ~pi175 & ~pi299;
  assign n11403 = pi184 & n8840;
  assign n11404 = ~pi184 & ~n8784;
  assign n11405 = ~pi189 & ~n11404;
  assign n11406 = ~n11403 & n11405;
  assign n11407 = pi184 & pi189;
  assign n11408 = ~n8859 & n11407;
  assign n11409 = ~n11358 & ~n11408;
  assign n11410 = ~n11406 & n11409;
  assign n11411 = n6166 & n11402;
  assign n11412 = ~n11410 & n11411;
  assign n11413 = ~n11353 & ~n11412;
  assign n11414 = ~n11377 & n11413;
  assign n11415 = ~n11401 & n11414;
  assign n11416 = ~pi39 & ~n11415;
  assign n11417 = pi232 & ~n11352;
  assign n11418 = ~n11416 & n11417;
  assign n11419 = ~pi40 & ~pi232;
  assign n11420 = ~pi38 & ~n11419;
  assign n11421 = ~n11418 & n11420;
  assign n11422 = ~n11334 & ~n11421;
  assign n11423 = n2573 & ~n11422;
  assign n11424 = pi87 & ~n11280;
  assign n11425 = n11315 & n11424;
  assign n11426 = ~n11313 & ~n11425;
  assign n11427 = ~n11423 & n11426;
  assign n11428 = n2572 & ~n11427;
  assign n11429 = ~n11312 & ~n11326;
  assign n11430 = ~n11428 & n11429;
  assign n11431 = ~pi54 & ~n11430;
  assign n11432 = ~n11311 & ~n11431;
  assign n11433 = ~pi74 & ~n11432;
  assign n11434 = n11304 & ~n11433;
  assign n11435 = pi55 & ~n11270;
  assign n11436 = pi163 & pi232;
  assign n11437 = ~pi92 & n2614;
  assign n11438 = n11436 & n11437;
  assign n11439 = n11335 & n11438;
  assign n11440 = n11280 & ~n11439;
  assign n11441 = ~pi75 & n11282;
  assign n11442 = ~n11440 & n11441;
  assign n11443 = n11273 & ~n11442;
  assign n11444 = ~pi54 & ~n11443;
  assign n11445 = ~n11279 & ~n11444;
  assign n11446 = ~pi74 & ~n11445;
  assign n11447 = n11435 & ~n11446;
  assign n11448 = n2530 & ~n11447;
  assign n11449 = ~n11434 & n11448;
  assign n11450 = n11292 & ~n11449;
  assign n11451 = ~n11278 & ~n11450;
  assign n11452 = pi79 & n11451;
  assign n11453 = pi39 & ~n9150;
  assign n11454 = n7230 & ~n11453;
  assign n11455 = n2489 & ~n8950;
  assign n11456 = ~pi40 & ~n11455;
  assign n11457 = ~n6166 & n8950;
  assign n11458 = n8937 & ~n11457;
  assign n11459 = n11436 & n11458;
  assign n11460 = n11456 & ~n11459;
  assign n11461 = ~pi39 & ~n11460;
  assign n11462 = n11454 & ~n11461;
  assign n11463 = pi87 & ~n2489;
  assign n11464 = n11280 & n11463;
  assign n11465 = n11282 & ~n11464;
  assign n11466 = ~n11462 & n11465;
  assign n11467 = ~n11272 & ~n11466;
  assign n11468 = n2572 & ~n11467;
  assign n11469 = ~n8972 & n11284;
  assign n11470 = n8890 & ~n11469;
  assign n11471 = ~n11271 & ~n11470;
  assign n11472 = ~n11468 & n11471;
  assign n11473 = ~pi54 & ~n11472;
  assign n11474 = ~n11279 & ~n11473;
  assign n11475 = ~pi74 & ~n11474;
  assign n11476 = n11435 & ~n11475;
  assign n11477 = n11315 & ~n11464;
  assign n11478 = n2489 & n11319;
  assign n11479 = n11456 & ~n11478;
  assign n11480 = ~pi39 & ~n11479;
  assign n11481 = n11454 & ~n11480;
  assign n11482 = n11477 & ~n11481;
  assign n11483 = ~n11313 & ~n11482;
  assign n11484 = n8890 & ~n11483;
  assign n11485 = n6197 & n9150;
  assign n11486 = n2489 & ~n8983;
  assign n11487 = ~pi40 & ~n11486;
  assign n11488 = ~n6197 & n11487;
  assign n11489 = ~n11485 & ~n11488;
  assign n11490 = ~n6221 & ~n11489;
  assign n11491 = ~pi40 & ~n8985;
  assign n11492 = n6221 & n11491;
  assign n11493 = ~n11490 & ~n11492;
  assign n11494 = n8979 & ~n11493;
  assign n11495 = n6194 & ~n11491;
  assign n11496 = ~n6194 & n11489;
  assign n11497 = ~n11495 & ~n11496;
  assign n11498 = n8752 & ~n11497;
  assign n11499 = ~n8752 & ~n9150;
  assign n11500 = ~pi299 & ~n11499;
  assign n11501 = ~n11498 & n11500;
  assign n11502 = ~pi232 & ~n11494;
  assign n11503 = ~n11501 & n11502;
  assign n11504 = ~pi189 & ~n11491;
  assign n11505 = n8772 & ~n9000;
  assign n11506 = n6205 & n11487;
  assign n11507 = ~n11485 & ~n11506;
  assign n11508 = ~n11505 & n11507;
  assign n11509 = pi189 & ~n6194;
  assign n11510 = n11508 & n11509;
  assign n11511 = ~n11504 & ~n11510;
  assign n11512 = pi179 & ~n11511;
  assign n11513 = n2489 & ~n9006;
  assign n11514 = n8772 & ~n11513;
  assign n11515 = n11507 & ~n11514;
  assign n11516 = ~pi189 & ~n11515;
  assign n11517 = pi189 & ~n11489;
  assign n11518 = ~pi179 & ~n6194;
  assign n11519 = ~n11517 & n11518;
  assign n11520 = ~n11516 & n11519;
  assign n11521 = ~n11495 & ~n11520;
  assign n11522 = ~n11512 & n11521;
  assign n11523 = n8752 & ~n11522;
  assign n11524 = ~n11499 & ~n11523;
  assign n11525 = ~pi299 & ~n11524;
  assign n11526 = ~n8739 & n9150;
  assign n11527 = pi299 & ~n11526;
  assign n11528 = ~pi166 & ~n6221;
  assign n11529 = n11493 & ~n11528;
  assign n11530 = n11515 & n11528;
  assign n11531 = n8739 & ~n11530;
  assign n11532 = ~n11529 & n11531;
  assign n11533 = n11527 & ~n11532;
  assign n11534 = ~n11525 & ~n11533;
  assign n11535 = ~pi156 & pi232;
  assign n11536 = ~n11534 & n11535;
  assign n11537 = pi166 & ~n6221;
  assign n11538 = n11508 & n11537;
  assign n11539 = ~n11491 & ~n11537;
  assign n11540 = n8739 & ~n11539;
  assign n11541 = ~n11538 & n11540;
  assign n11542 = n11527 & ~n11541;
  assign n11543 = ~n11525 & ~n11542;
  assign n11544 = pi156 & pi232;
  assign n11545 = ~n11543 & n11544;
  assign n11546 = pi39 & ~n11503;
  assign n11547 = ~n11536 & n11546;
  assign n11548 = ~n11545 & n11547;
  assign n11549 = ~n2442 & ~n9166;
  assign n11550 = n9033 & ~n9034;
  assign n11551 = ~n11549 & ~n11550;
  assign n11552 = ~pi40 & ~n9305;
  assign n11553 = ~pi95 & ~n11552;
  assign n11554 = ~n11551 & ~n11553;
  assign n11555 = ~pi299 & n11554;
  assign n11556 = ~pi40 & ~n9200;
  assign n11557 = ~pi95 & ~n11556;
  assign n11558 = ~n11551 & ~n11557;
  assign n11559 = pi299 & n11558;
  assign n11560 = ~pi232 & ~n11555;
  assign n11561 = ~n11559 & n11560;
  assign n11562 = ~n6166 & n11554;
  assign n11563 = ~pi40 & ~n9097;
  assign n11564 = ~pi95 & ~n11563;
  assign n11565 = ~pi40 & ~n9089;
  assign n11566 = pi189 & n11565;
  assign n11567 = n11564 & ~n11566;
  assign n11568 = pi182 & n9166;
  assign n11569 = ~pi182 & n11551;
  assign n11570 = n6166 & ~n11569;
  assign n11571 = ~n11568 & n11570;
  assign n11572 = ~n11567 & n11571;
  assign n11573 = pi184 & ~n11572;
  assign n11574 = ~pi40 & n9187;
  assign n11575 = ~pi32 & ~n11574;
  assign n11576 = ~n9151 & ~n11575;
  assign n11577 = ~pi95 & ~n11576;
  assign n11578 = ~n9166 & ~n11577;
  assign n11579 = pi198 & ~n11578;
  assign n11580 = ~n9168 & ~n11575;
  assign n11581 = ~pi95 & ~n11580;
  assign n11582 = ~n9166 & ~n11581;
  assign n11583 = ~pi198 & ~n11582;
  assign n11584 = n9927 & ~n11579;
  assign n11585 = ~n11583 & n11584;
  assign n11586 = pi189 & n6166;
  assign n11587 = n11552 & n11586;
  assign n11588 = pi182 & ~pi184;
  assign n11589 = ~n11585 & n11588;
  assign n11590 = ~n11587 & n11589;
  assign n11591 = ~n11573 & ~n11590;
  assign n11592 = n11402 & ~n11591;
  assign n11593 = pi95 & ~pi182;
  assign n11594 = ~pi40 & ~n9106;
  assign n11595 = ~pi95 & pi189;
  assign n11596 = n2489 & ~n11595;
  assign n11597 = n11594 & ~n11596;
  assign n11598 = ~n11593 & ~n11597;
  assign n11599 = n11295 & ~n11598;
  assign n11600 = ~n11569 & n11599;
  assign n11601 = ~pi95 & ~n9161;
  assign n11602 = pi198 & ~n11601;
  assign n11603 = ~pi198 & ~n9170;
  assign n11604 = ~n11602 & ~n11603;
  assign n11605 = pi189 & n11571;
  assign n11606 = ~n11604 & n11605;
  assign n11607 = ~n9276 & ~n11593;
  assign n11608 = ~pi189 & n11570;
  assign n11609 = ~n11607 & n11608;
  assign n11610 = ~n11606 & ~n11609;
  assign n11611 = ~pi184 & ~n11610;
  assign n11612 = n11373 & ~n11600;
  assign n11613 = ~n11611 & n11612;
  assign n11614 = ~n11592 & ~n11613;
  assign n11615 = ~n11562 & ~n11614;
  assign n11616 = ~n6166 & n11558;
  assign n11617 = ~pi95 & ~n11594;
  assign n11618 = pi166 & ~n11617;
  assign n11619 = ~n11070 & ~n11617;
  assign n11620 = pi153 & ~n11618;
  assign n11621 = ~n11619 & n11620;
  assign n11622 = pi166 & n11565;
  assign n11623 = n11564 & ~n11622;
  assign n11624 = ~pi153 & n11623;
  assign n11625 = ~pi160 & n6166;
  assign n11626 = ~n11621 & n11625;
  assign n11627 = ~n11551 & n11626;
  assign n11628 = ~n11624 & n11627;
  assign n11629 = n6166 & ~n9166;
  assign n11630 = n11618 & n11629;
  assign n11631 = n9150 & n9931;
  assign n11632 = pi153 & ~n11631;
  assign n11633 = ~n11630 & n11632;
  assign n11634 = ~n11623 & n11629;
  assign n11635 = ~pi153 & ~n11634;
  assign n11636 = pi160 & ~n11633;
  assign n11637 = ~n11635 & n11636;
  assign n11638 = pi163 & ~n11628;
  assign n11639 = ~n11637 & n11638;
  assign n11640 = ~pi210 & n9170;
  assign n11641 = pi210 & n11601;
  assign n11642 = n11386 & ~n11640;
  assign n11643 = ~n11641 & n11642;
  assign n11644 = ~pi210 & n9270;
  assign n11645 = pi210 & n9273;
  assign n11646 = n9931 & ~n11644;
  assign n11647 = ~n11645 & n11646;
  assign n11648 = pi153 & ~n11647;
  assign n11649 = ~n11643 & n11648;
  assign n11650 = n11386 & n11556;
  assign n11651 = pi210 & ~n11578;
  assign n11652 = ~pi210 & ~n11582;
  assign n11653 = ~n11651 & ~n11652;
  assign n11654 = n9931 & n11653;
  assign n11655 = ~pi153 & ~n11654;
  assign n11656 = ~n11650 & n11655;
  assign n11657 = pi153 & n9166;
  assign n11658 = pi160 & ~n11657;
  assign n11659 = ~n11656 & n11658;
  assign n11660 = pi166 & ~n11557;
  assign n11661 = ~pi166 & n11653;
  assign n11662 = ~pi95 & ~n11661;
  assign n11663 = n6166 & ~n11662;
  assign n11664 = ~pi153 & ~n11663;
  assign n11665 = ~n11660 & n11664;
  assign n11666 = ~pi160 & ~n11551;
  assign n11667 = ~n11665 & n11666;
  assign n11668 = ~n11659 & ~n11667;
  assign n11669 = ~n11649 & ~n11668;
  assign n11670 = ~pi163 & ~n11669;
  assign n11671 = ~n11639 & ~n11670;
  assign n11672 = pi299 & ~n11616;
  assign n11673 = ~n11671 & n11672;
  assign n11674 = ~n9927 & n11554;
  assign n11675 = ~n11551 & ~n11577;
  assign n11676 = pi198 & ~n11675;
  assign n11677 = ~n11551 & ~n11581;
  assign n11678 = ~pi198 & ~n11677;
  assign n11679 = n9927 & ~n11676;
  assign n11680 = ~n11678 & n11679;
  assign n11681 = ~pi182 & ~pi184;
  assign n11682 = n11402 & n11681;
  assign n11683 = ~n11680 & n11682;
  assign n11684 = ~n11674 & n11683;
  assign n11685 = ~n11615 & ~n11684;
  assign n11686 = ~n11673 & n11685;
  assign n11687 = pi232 & ~n11686;
  assign n11688 = ~pi39 & ~n11561;
  assign n11689 = ~n11687 & n11688;
  assign n11690 = ~pi38 & ~n11548;
  assign n11691 = ~n11689 & n11690;
  assign n11692 = ~n11334 & ~n11691;
  assign n11693 = n2573 & ~n11692;
  assign n11694 = pi87 & n11477;
  assign n11695 = ~n11313 & ~n11694;
  assign n11696 = ~n11693 & n11695;
  assign n11697 = n2572 & ~n11696;
  assign n11698 = ~n11312 & ~n11484;
  assign n11699 = ~n11697 & n11698;
  assign n11700 = ~pi54 & ~n11699;
  assign n11701 = ~n11311 & ~n11700;
  assign n11702 = ~pi74 & ~n11701;
  assign n11703 = n11304 & ~n11702;
  assign n11704 = n2530 & ~n11476;
  assign n11705 = ~n11703 & n11704;
  assign n11706 = ~n8941 & n11292;
  assign n11707 = ~n11705 & n11706;
  assign n11708 = ~n11278 & ~n11707;
  assign n11709 = ~pi79 & n11708;
  assign n11710 = ~pi34 & n9695;
  assign n11711 = ~n11452 & ~n11710;
  assign n11712 = ~n11709 & n11711;
  assign n11713 = ~pi79 & ~n8682;
  assign n11714 = n11451 & n11713;
  assign n11715 = n11708 & ~n11713;
  assign n11716 = n11710 & ~n11714;
  assign n11717 = ~n11715 & n11716;
  assign po237 = n11712 | n11717;
  assign n11719 = pi98 & pi1092;
  assign n11720 = pi1093 & n11719;
  assign n11721 = ~pi567 & n2923;
  assign n11722 = ~n11720 & ~n11721;
  assign n11723 = ~pi80 & ~n11722;
  assign n11724 = pi217 & ~n11723;
  assign n11725 = n7356 & n11722;
  assign n11726 = ~n7579 & n11722;
  assign n11727 = pi588 & ~n11726;
  assign n11728 = ~n7658 & n7688;
  assign n11729 = n11722 & ~n11728;
  assign n11730 = ~pi1199 & ~n11729;
  assign n11731 = n7658 & ~n7670;
  assign n11732 = n7688 & ~n11731;
  assign n11733 = n11722 & ~n11732;
  assign n11734 = ~pi430 & n11733;
  assign n11735 = n7658 & n7670;
  assign n11736 = n7688 & ~n11735;
  assign n11737 = n11722 & ~n11736;
  assign n11738 = pi430 & n11737;
  assign n11739 = ~pi426 & ~n11734;
  assign n11740 = ~n11738 & n11739;
  assign n11741 = ~pi430 & n11737;
  assign n11742 = pi430 & n11733;
  assign n11743 = pi426 & ~n11741;
  assign n11744 = ~n11742 & n11743;
  assign n11745 = ~n11740 & ~n11744;
  assign n11746 = ~n8093 & ~n11745;
  assign n11747 = n7673 & n11733;
  assign n11748 = ~n7673 & n11737;
  assign n11749 = n8093 & ~n11747;
  assign n11750 = ~n11748 & n11749;
  assign n11751 = ~n11746 & ~n11750;
  assign n11752 = pi1199 & ~n11751;
  assign n11753 = n7579 & ~n11730;
  assign n11754 = ~n11752 & n11753;
  assign n11755 = n11727 & ~n11754;
  assign n11756 = pi591 & ~n11722;
  assign n11757 = pi590 & ~n11756;
  assign n11758 = pi461 & ~n7798;
  assign n11759 = ~pi461 & ~n7909;
  assign n11760 = ~n11758 & ~n11759;
  assign n11761 = pi1199 & ~n11760;
  assign n11762 = ~n7902 & n11761;
  assign n11763 = n7902 & n11760;
  assign n11764 = ~n7766 & n11722;
  assign n11765 = ~n11762 & n11764;
  assign n11766 = ~n11763 & n11765;
  assign n11767 = n7881 & n11766;
  assign n11768 = ~n7688 & n11722;
  assign n11769 = ~pi591 & ~n11768;
  assign n11770 = ~n11767 & n11769;
  assign n11771 = n11757 & ~n11770;
  assign n11772 = n7766 & ~n7793;
  assign n11773 = n11722 & ~n11772;
  assign n11774 = ~pi591 & ~n11773;
  assign n11775 = ~pi1197 & ~n8231;
  assign n11776 = ~n11768 & ~n11775;
  assign n11777 = pi592 & ~n11722;
  assign n11778 = ~pi1196 & ~n11722;
  assign n11779 = ~n11777 & ~n11778;
  assign n11780 = ~n7949 & ~n7952;
  assign n11781 = n7949 & n7952;
  assign n11782 = ~n11780 & ~n11781;
  assign n11783 = n7348 & n11782;
  assign n11784 = ~n11719 & ~n11783;
  assign n11785 = ~pi412 & ~n11784;
  assign n11786 = n7348 & ~n11782;
  assign n11787 = ~n11719 & ~n11786;
  assign n11788 = pi412 & ~n11787;
  assign n11789 = n7961 & ~n11785;
  assign n11790 = ~n11788 & n11789;
  assign n11791 = pi412 & ~n11784;
  assign n11792 = ~pi412 & ~n11787;
  assign n11793 = ~n7961 & ~n11791;
  assign n11794 = ~n11792 & n11793;
  assign n11795 = ~pi122 & ~n11790;
  assign n11796 = ~n11794 & n11795;
  assign n11797 = ~pi122 & ~n11796;
  assign n11798 = n7561 & ~n11797;
  assign n11799 = ~n7418 & ~n11719;
  assign n11800 = n11798 & ~n11799;
  assign n11801 = pi1091 & n11720;
  assign n11802 = ~n11800 & ~n11801;
  assign n11803 = pi567 & ~n11802;
  assign n11804 = ~n11721 & ~n11803;
  assign n11805 = n7654 & ~n11804;
  assign n11806 = n11779 & ~n11805;
  assign n11807 = ~pi1199 & ~n11806;
  assign n11808 = ~n7561 & ~n11801;
  assign n11809 = n7348 & n7941;
  assign n11810 = ~pi122 & ~n11719;
  assign n11811 = ~n11809 & n11810;
  assign n11812 = ~n11808 & ~n11811;
  assign n11813 = ~n11799 & n11812;
  assign n11814 = pi567 & n11813;
  assign n11815 = ~n11721 & ~n11814;
  assign n11816 = ~n11803 & n11815;
  assign n11817 = n7654 & ~n11816;
  assign n11818 = n8445 & ~n11815;
  assign n11819 = ~n11777 & ~n11818;
  assign n11820 = ~n11817 & n11819;
  assign n11821 = pi1199 & ~n11820;
  assign n11822 = ~n11807 & ~n11821;
  assign n11823 = n11775 & ~n11822;
  assign n11824 = ~n11776 & ~n11823;
  assign n11825 = ~pi333 & ~n11824;
  assign n11826 = n8231 & ~n11768;
  assign n11827 = ~n8231 & ~n11822;
  assign n11828 = ~n11826 & ~n11827;
  assign n11829 = pi333 & ~n11828;
  assign n11830 = ~n11825 & ~n11829;
  assign n11831 = ~pi391 & ~n11830;
  assign n11832 = pi333 & ~n11824;
  assign n11833 = ~pi333 & ~n11828;
  assign n11834 = ~n11832 & ~n11833;
  assign n11835 = pi391 & ~n11834;
  assign n11836 = n8023 & ~n11831;
  assign n11837 = ~n11835 & n11836;
  assign n11838 = ~pi391 & ~n11834;
  assign n11839 = pi391 & ~n11830;
  assign n11840 = ~n8023 & ~n11838;
  assign n11841 = ~n11839 & n11840;
  assign n11842 = pi591 & ~n11837;
  assign n11843 = ~n11841 & n11842;
  assign n11844 = ~pi590 & ~n11774;
  assign n11845 = ~n11843 & n11844;
  assign n11846 = ~pi588 & ~n11771;
  assign n11847 = ~n11845 & n11846;
  assign n11848 = ~n7356 & ~n11755;
  assign n11849 = ~n11847 & n11848;
  assign n11850 = ~pi80 & po1038;
  assign n11851 = ~n11725 & n11850;
  assign n11852 = ~n11849 & n11851;
  assign n11853 = ~n7360 & n11722;
  assign n11854 = n7360 & ~n11721;
  assign n11855 = pi824 & pi950;
  assign n11856 = ~pi51 & n10656;
  assign n11857 = ~pi88 & n2495;
  assign n11858 = n10016 & n11857;
  assign n11859 = ~pi110 & n2706;
  assign n11860 = n11858 & n11859;
  assign n11861 = n7371 & n11860;
  assign n11862 = n7377 & n11861;
  assign n11863 = n11855 & n11856;
  assign n11864 = n11862 & n11863;
  assign n11865 = ~pi98 & ~n11864;
  assign n11866 = pi1092 & ~n11865;
  assign n11867 = n8049 & ~n11808;
  assign n11868 = n11866 & n11867;
  assign n11869 = pi51 & n11862;
  assign n11870 = pi90 & pi93;
  assign n11871 = ~pi841 & ~n2709;
  assign n11872 = ~n11870 & n11871;
  assign n11873 = n2509 & n11872;
  assign n11874 = n11861 & n11873;
  assign n11875 = ~n11869 & ~n11874;
  assign n11876 = n10656 & n11855;
  assign n11877 = ~n11875 & n11876;
  assign n11878 = ~pi98 & ~n11877;
  assign n11879 = pi1092 & ~n11878;
  assign n11880 = n2615 & ~n11808;
  assign n11881 = n11879 & n11880;
  assign n11882 = ~n2628 & n11720;
  assign n11883 = ~pi75 & ~n11882;
  assign n11884 = ~n11868 & n11883;
  assign n11885 = ~n11881 & n11884;
  assign n11886 = pi75 & ~n11720;
  assign n11887 = pi567 & ~n11886;
  assign n11888 = ~n11885 & n11887;
  assign n11889 = n11854 & ~n11888;
  assign n11890 = ~n11853 & ~n11889;
  assign n11891 = ~pi592 & n11890;
  assign n11892 = ~n11777 & ~n11891;
  assign n11893 = ~n7631 & n11892;
  assign n11894 = n7631 & ~n11778;
  assign n11895 = ~pi443 & ~n11722;
  assign n11896 = pi443 & ~n11892;
  assign n11897 = ~n11895 & ~n11896;
  assign n11898 = pi436 & ~pi444;
  assign n11899 = ~pi436 & pi444;
  assign n11900 = ~n11898 & ~n11899;
  assign n11901 = ~n11897 & ~n11900;
  assign n11902 = pi443 & ~n11722;
  assign n11903 = ~pi443 & ~n11892;
  assign n11904 = ~n11902 & ~n11903;
  assign n11905 = n11900 & ~n11904;
  assign n11906 = ~n7652 & ~n11901;
  assign n11907 = ~n11905 & n11906;
  assign n11908 = ~n8061 & ~n11897;
  assign n11909 = n8061 & ~n11904;
  assign n11910 = n7652 & ~n11908;
  assign n11911 = ~n11909 & n11910;
  assign n11912 = pi1196 & ~n11907;
  assign n11913 = ~n11911 & n11912;
  assign n11914 = n11894 & ~n11913;
  assign n11915 = ~n11893 & ~n11914;
  assign n11916 = ~pi1199 & n11915;
  assign n11917 = pi426 & ~n8093;
  assign n11918 = ~pi426 & n8093;
  assign n11919 = ~n11917 & ~n11918;
  assign n11920 = pi428 & ~n11915;
  assign n11921 = ~pi428 & n11892;
  assign n11922 = ~n11920 & ~n11921;
  assign n11923 = pi427 & ~n11922;
  assign n11924 = pi428 & ~n11892;
  assign n11925 = ~pi428 & n11915;
  assign n11926 = ~n11924 & ~n11925;
  assign n11927 = ~pi427 & n11926;
  assign n11928 = ~n11923 & ~n11927;
  assign n11929 = pi430 & n11928;
  assign n11930 = ~pi427 & ~n11922;
  assign n11931 = pi427 & n11926;
  assign n11932 = ~n11930 & ~n11931;
  assign n11933 = ~pi430 & n11932;
  assign n11934 = n11919 & ~n11929;
  assign n11935 = ~n11933 & n11934;
  assign n11936 = ~pi430 & n11928;
  assign n11937 = pi430 & n11932;
  assign n11938 = ~n11919 & ~n11936;
  assign n11939 = ~n11937 & n11938;
  assign n11940 = pi1199 & ~n11935;
  assign n11941 = ~n11939 & n11940;
  assign n11942 = n7579 & ~n11916;
  assign n11943 = ~n11941 & n11942;
  assign n11944 = n11727 & ~n11943;
  assign n11945 = ~n11775 & ~n11892;
  assign n11946 = n8240 & n11854;
  assign n11947 = ~n11722 & ~n11946;
  assign n11948 = ~pi592 & ~n11853;
  assign n11949 = ~n7941 & n11719;
  assign n11950 = n7941 & n11866;
  assign n11951 = ~n11949 & ~n11950;
  assign n11952 = n11868 & ~n11951;
  assign n11953 = n7941 & n11879;
  assign n11954 = ~n11949 & ~n11953;
  assign n11955 = n11881 & ~n11954;
  assign n11956 = n7967 & n11719;
  assign n11957 = ~n7967 & n11879;
  assign n11958 = ~n11956 & ~n11957;
  assign n11959 = n11880 & ~n11958;
  assign n11960 = ~n7967 & n11866;
  assign n11961 = ~n11956 & ~n11960;
  assign n11962 = n11867 & ~n11961;
  assign n11963 = ~n11959 & ~n11962;
  assign n11964 = pi1196 & ~n11963;
  assign n11965 = ~n11882 & ~n11952;
  assign n11966 = ~n11955 & n11965;
  assign n11967 = ~n11964 & n11966;
  assign n11968 = ~pi75 & pi567;
  assign n11969 = n11948 & n11968;
  assign n11970 = ~n11967 & n11969;
  assign n11971 = pi1199 & ~n11947;
  assign n11972 = ~n11970 & n11971;
  assign n11973 = ~pi98 & n11963;
  assign n11974 = n11888 & ~n11973;
  assign n11975 = n11854 & ~n11974;
  assign n11976 = pi1196 & n11948;
  assign n11977 = ~n11975 & n11976;
  assign n11978 = ~pi1199 & n11779;
  assign n11979 = ~n11977 & n11978;
  assign n11980 = ~n8231 & ~n11972;
  assign n11981 = ~n11979 & n11980;
  assign n11982 = ~pi1197 & n11981;
  assign n11983 = ~n11945 & ~n11982;
  assign n11984 = pi333 & ~n11983;
  assign n11985 = n8231 & ~n11892;
  assign n11986 = ~n11981 & ~n11985;
  assign n11987 = ~pi333 & ~n11986;
  assign n11988 = ~n11984 & ~n11987;
  assign n11989 = ~pi391 & ~n11988;
  assign n11990 = ~pi333 & ~n11983;
  assign n11991 = pi333 & ~n11986;
  assign n11992 = ~n11990 & ~n11991;
  assign n11993 = pi391 & ~n11992;
  assign n11994 = ~n11989 & ~n11993;
  assign n11995 = ~pi392 & ~n11994;
  assign n11996 = ~pi391 & ~n11992;
  assign n11997 = pi391 & ~n11988;
  assign n11998 = ~n11996 & ~n11997;
  assign n11999 = pi392 & ~n11998;
  assign n12000 = pi393 & ~n8017;
  assign n12001 = ~pi393 & n8017;
  assign n12002 = ~n12000 & ~n12001;
  assign n12003 = ~n11995 & ~n12002;
  assign n12004 = ~n11999 & n12003;
  assign n12005 = ~pi392 & ~n11998;
  assign n12006 = pi392 & ~n11994;
  assign n12007 = n12002 & ~n12005;
  assign n12008 = ~n12006 & n12007;
  assign n12009 = pi591 & ~n12004;
  assign n12010 = ~n12008 & n12009;
  assign n12011 = n7765 & n11722;
  assign n12012 = ~pi592 & ~n11722;
  assign n12013 = pi592 & n11890;
  assign n12014 = ~n12012 & ~n12013;
  assign n12015 = ~n7765 & n12014;
  assign n12016 = ~n12011 & ~n12015;
  assign n12017 = ~pi1198 & ~n12016;
  assign n12018 = pi1198 & n12014;
  assign n12019 = ~n12017 & ~n12018;
  assign n12020 = pi374 & ~n12019;
  assign n12021 = ~pi374 & ~n12016;
  assign n12022 = ~n12020 & ~n12021;
  assign n12023 = ~n7787 & ~n12022;
  assign n12024 = pi374 & ~n12016;
  assign n12025 = ~pi374 & ~n12019;
  assign n12026 = ~n12024 & ~n12025;
  assign n12027 = n7787 & ~n12026;
  assign n12028 = ~pi591 & ~n12023;
  assign n12029 = ~n12027 & n12028;
  assign n12030 = ~pi590 & ~n12029;
  assign n12031 = ~n12010 & n12030;
  assign n12032 = n7852 & n11722;
  assign n12033 = ~n7852 & n11892;
  assign n12034 = ~n12032 & ~n12033;
  assign n12035 = pi1198 & ~n12034;
  assign n12036 = ~pi1198 & ~n11778;
  assign n12037 = ~n7801 & n11722;
  assign n12038 = n7801 & n11892;
  assign n12039 = ~n12037 & ~n12038;
  assign n12040 = n7819 & ~n12039;
  assign n12041 = pi452 & ~pi455;
  assign n12042 = ~pi452 & pi455;
  assign n12043 = ~n12041 & ~n12042;
  assign n12044 = ~n11722 & ~n12043;
  assign n12045 = ~n11892 & n12043;
  assign n12046 = ~n7819 & ~n12044;
  assign n12047 = ~n12045 & n12046;
  assign n12048 = pi1196 & ~n12047;
  assign n12049 = ~n12040 & n12048;
  assign n12050 = n12036 & ~n12049;
  assign n12051 = ~n12035 & ~n12050;
  assign n12052 = ~n7879 & ~n12051;
  assign n12053 = n7879 & n11892;
  assign n12054 = ~n12052 & ~n12053;
  assign n12055 = ~n7798 & n12054;
  assign n12056 = pi1199 & ~n11892;
  assign n12057 = pi351 & n12056;
  assign n12058 = ~n12055 & ~n12057;
  assign n12059 = ~pi461 & ~n12058;
  assign n12060 = ~n7909 & n12054;
  assign n12061 = ~pi351 & n12056;
  assign n12062 = ~n12060 & ~n12061;
  assign n12063 = pi461 & ~n12062;
  assign n12064 = ~n12059 & ~n12063;
  assign n12065 = ~pi357 & ~n12064;
  assign n12066 = ~pi461 & ~n12062;
  assign n12067 = pi461 & ~n12058;
  assign n12068 = ~n12066 & ~n12067;
  assign n12069 = pi357 & ~n12068;
  assign n12070 = ~n12065 & ~n12069;
  assign n12071 = ~pi356 & ~n12070;
  assign n12072 = ~pi357 & ~n12068;
  assign n12073 = pi357 & ~n12064;
  assign n12074 = ~n12072 & ~n12073;
  assign n12075 = pi356 & ~n12074;
  assign n12076 = ~n7899 & ~n12071;
  assign n12077 = ~n12075 & n12076;
  assign n12078 = ~pi356 & ~n12074;
  assign n12079 = pi356 & ~n12070;
  assign n12080 = n7899 & ~n12078;
  assign n12081 = ~n12079 & n12080;
  assign n12082 = ~pi591 & ~n12077;
  assign n12083 = ~n12081 & n12082;
  assign n12084 = n11757 & ~n12083;
  assign n12085 = ~pi588 & ~n12031;
  assign n12086 = ~n12084 & n12085;
  assign n12087 = n7356 & ~n11944;
  assign n12088 = ~n12086 & n12087;
  assign n12089 = pi567 & n7360;
  assign n12090 = ~n7351 & ~n11720;
  assign n12091 = ~pi122 & n12090;
  assign n12092 = n7561 & ~n12091;
  assign n12093 = n2628 & ~n11801;
  assign n12094 = ~n12092 & n12093;
  assign n12095 = n2615 & ~n11801;
  assign n12096 = ~n11879 & n12095;
  assign n12097 = pi87 & n12093;
  assign n12098 = ~n11866 & n12097;
  assign n12099 = ~n12096 & ~n12098;
  assign n12100 = pi122 & ~n12099;
  assign n12101 = ~n12094 & ~n12100;
  assign n12102 = ~pi75 & ~n12101;
  assign n12103 = ~n7361 & n12090;
  assign n12104 = n12089 & ~n12103;
  assign n12105 = ~n12102 & n12104;
  assign n12106 = ~n7360 & ~n12090;
  assign n12107 = ~n11721 & ~n12106;
  assign n12108 = ~n12105 & n12107;
  assign n12109 = ~pi592 & ~n12108;
  assign n12110 = ~n11777 & ~n12109;
  assign n12111 = ~n7631 & n12110;
  assign n12112 = pi443 & ~n12110;
  assign n12113 = n8064 & ~n11895;
  assign n12114 = ~n12112 & n12113;
  assign n12115 = ~pi443 & ~n12110;
  assign n12116 = ~n8064 & ~n11902;
  assign n12117 = ~n12115 & n12116;
  assign n12118 = pi1196 & ~n12114;
  assign n12119 = ~n12117 & n12118;
  assign n12120 = n11894 & ~n12119;
  assign n12121 = ~n12111 & ~n12120;
  assign n12122 = ~pi1199 & n12121;
  assign n12123 = pi428 & ~n12121;
  assign n12124 = ~pi428 & n12110;
  assign n12125 = ~n12123 & ~n12124;
  assign n12126 = pi427 & ~n12125;
  assign n12127 = pi428 & ~n12110;
  assign n12128 = ~pi428 & n12121;
  assign n12129 = ~n12127 & ~n12128;
  assign n12130 = ~pi427 & n12129;
  assign n12131 = ~n12126 & ~n12130;
  assign n12132 = pi430 & n12131;
  assign n12133 = ~pi427 & ~n12125;
  assign n12134 = pi427 & n12129;
  assign n12135 = ~n12133 & ~n12134;
  assign n12136 = ~pi430 & n12135;
  assign n12137 = n11919 & ~n12132;
  assign n12138 = ~n12136 & n12137;
  assign n12139 = pi430 & n12135;
  assign n12140 = ~pi430 & n12131;
  assign n12141 = ~n11919 & ~n12139;
  assign n12142 = ~n12140 & n12141;
  assign n12143 = pi1199 & ~n12138;
  assign n12144 = ~n12142 & n12143;
  assign n12145 = n7579 & ~n12122;
  assign n12146 = ~n12144 & n12145;
  assign n12147 = n11727 & ~n12146;
  assign n12148 = ~pi1197 & ~n11722;
  assign n12149 = ~n7760 & ~n7761;
  assign n12150 = n11722 & ~n12149;
  assign n12151 = pi592 & ~n12108;
  assign n12152 = ~n12012 & ~n12151;
  assign n12153 = n12149 & n12152;
  assign n12154 = pi1197 & ~n12150;
  assign n12155 = ~n12153 & n12154;
  assign n12156 = ~n7738 & ~n12148;
  assign n12157 = ~n12155 & n12156;
  assign n12158 = n7738 & n12152;
  assign n12159 = ~pi1199 & ~n12158;
  assign n12160 = ~n12157 & n12159;
  assign n12161 = ~n7712 & n7764;
  assign n12162 = n12152 & ~n12161;
  assign n12163 = pi1199 & ~n12011;
  assign n12164 = ~n12162 & n12163;
  assign n12165 = ~n12160 & ~n12164;
  assign n12166 = ~pi374 & n12165;
  assign n12167 = pi1198 & ~n12152;
  assign n12168 = pi374 & ~n12167;
  assign n12169 = ~n7787 & ~n12168;
  assign n12170 = ~n12166 & n12169;
  assign n12171 = ~pi374 & ~n12167;
  assign n12172 = n7787 & ~n12171;
  assign n12173 = ~pi374 & n12172;
  assign n12174 = n12165 & ~n12173;
  assign n12175 = pi1198 & ~n12172;
  assign n12176 = ~n12174 & ~n12175;
  assign n12177 = ~pi591 & ~n12170;
  assign n12178 = ~n12176 & n12177;
  assign n12179 = n8231 & ~n12110;
  assign n12180 = ~n11815 & ~n11854;
  assign n12181 = ~n7361 & ~n11813;
  assign n12182 = n12089 & ~n12181;
  assign n12183 = n11954 & n12095;
  assign n12184 = n11951 & n12097;
  assign n12185 = ~n12183 & ~n12184;
  assign n12186 = pi122 & ~n12185;
  assign n12187 = n2628 & ~n11812;
  assign n12188 = ~n12186 & ~n12187;
  assign n12189 = ~pi75 & ~n12188;
  assign n12190 = n12182 & ~n12189;
  assign n12191 = ~n12180 & ~n12190;
  assign n12192 = n8445 & ~n12191;
  assign n12193 = ~n11816 & ~n11854;
  assign n12194 = ~n11800 & n12187;
  assign n12195 = ~pi122 & n11809;
  assign n12196 = n11961 & n12097;
  assign n12197 = n11958 & n12095;
  assign n12198 = ~n12196 & ~n12197;
  assign n12199 = ~n11796 & ~n12198;
  assign n12200 = ~n12185 & ~n12195;
  assign n12201 = n12199 & n12200;
  assign n12202 = ~n12194 & ~n12201;
  assign n12203 = ~pi75 & ~n12202;
  assign n12204 = ~n7361 & n11802;
  assign n12205 = n12089 & ~n12204;
  assign n12206 = ~n12182 & ~n12205;
  assign n12207 = ~n12203 & ~n12206;
  assign n12208 = ~n12193 & ~n12207;
  assign n12209 = n7654 & ~n12208;
  assign n12210 = pi1199 & ~n12192;
  assign n12211 = ~n12209 & n12210;
  assign n12212 = ~n11804 & ~n11854;
  assign n12213 = ~n11798 & n12093;
  assign n12214 = ~n12199 & ~n12213;
  assign n12215 = ~pi75 & ~n12214;
  assign n12216 = n12205 & ~n12215;
  assign n12217 = ~n12212 & ~n12216;
  assign n12218 = n7654 & ~n12217;
  assign n12219 = ~pi1199 & ~n11778;
  assign n12220 = ~n12218 & n12219;
  assign n12221 = ~n12211 & ~n12220;
  assign n12222 = ~n11777 & ~n12221;
  assign n12223 = ~n8231 & ~n12222;
  assign n12224 = ~n12179 & ~n12223;
  assign n12225 = pi333 & ~n12224;
  assign n12226 = ~n11775 & n12110;
  assign n12227 = n11775 & n12222;
  assign n12228 = ~n12226 & ~n12227;
  assign n12229 = ~pi333 & n12228;
  assign n12230 = ~n12225 & ~n12229;
  assign n12231 = pi391 & ~n12230;
  assign n12232 = pi333 & ~n12228;
  assign n12233 = ~pi333 & n12224;
  assign n12234 = ~n12232 & ~n12233;
  assign n12235 = ~pi391 & n12234;
  assign n12236 = ~n12231 & ~n12235;
  assign n12237 = pi392 & ~n12236;
  assign n12238 = pi391 & ~n12234;
  assign n12239 = ~pi391 & n12230;
  assign n12240 = ~n12238 & ~n12239;
  assign n12241 = ~pi392 & n12240;
  assign n12242 = ~n12237 & ~n12241;
  assign n12243 = n12002 & ~n12242;
  assign n12244 = pi392 & ~n12240;
  assign n12245 = ~pi392 & n12236;
  assign n12246 = ~n12002 & ~n12244;
  assign n12247 = ~n12245 & n12246;
  assign n12248 = pi591 & ~n12243;
  assign n12249 = ~n12247 & n12248;
  assign n12250 = ~n12178 & ~n12249;
  assign n12251 = ~pi590 & ~n12250;
  assign n12252 = ~n7852 & n12110;
  assign n12253 = ~n12032 & ~n12252;
  assign n12254 = pi1198 & ~n12253;
  assign n12255 = n7801 & n12110;
  assign n12256 = ~n12037 & ~n12255;
  assign n12257 = n7819 & ~n12256;
  assign n12258 = n12043 & ~n12110;
  assign n12259 = n12046 & ~n12258;
  assign n12260 = pi1196 & ~n12259;
  assign n12261 = ~n12257 & n12260;
  assign n12262 = n12036 & ~n12261;
  assign n12263 = ~n12254 & ~n12262;
  assign n12264 = ~n7879 & ~n12263;
  assign n12265 = n7879 & n12110;
  assign n12266 = ~n12264 & ~n12265;
  assign n12267 = ~n7909 & n12266;
  assign n12268 = pi1199 & ~n12110;
  assign n12269 = ~pi351 & n12268;
  assign n12270 = ~n12267 & ~n12269;
  assign n12271 = ~pi461 & ~n12270;
  assign n12272 = ~n7798 & n12266;
  assign n12273 = pi351 & n12268;
  assign n12274 = ~n12272 & ~n12273;
  assign n12275 = pi461 & ~n12274;
  assign n12276 = ~n12271 & ~n12275;
  assign n12277 = ~pi357 & n12276;
  assign n12278 = ~pi461 & ~n12274;
  assign n12279 = pi461 & ~n12270;
  assign n12280 = ~n12278 & ~n12279;
  assign n12281 = pi357 & n12280;
  assign n12282 = ~pi356 & ~n12277;
  assign n12283 = ~n12281 & n12282;
  assign n12284 = ~pi357 & n12280;
  assign n12285 = pi357 & n12276;
  assign n12286 = pi356 & ~n12284;
  assign n12287 = ~n12285 & n12286;
  assign n12288 = ~n12283 & ~n12287;
  assign n12289 = n7899 & ~n12288;
  assign n12290 = ~n7887 & n12280;
  assign n12291 = n7887 & n12276;
  assign n12292 = ~n7899 & ~n12290;
  assign n12293 = ~n12291 & n12292;
  assign n12294 = ~n12289 & ~n12293;
  assign n12295 = ~pi591 & ~n12294;
  assign n12296 = n11757 & ~n12295;
  assign n12297 = ~pi588 & ~n12251;
  assign n12298 = ~n12296 & n12297;
  assign n12299 = ~n7356 & ~n12147;
  assign n12300 = ~n12298 & n12299;
  assign n12301 = ~pi80 & ~po1038;
  assign n12302 = ~n12088 & n12301;
  assign n12303 = ~n12300 & n12302;
  assign n12304 = ~pi217 & ~n11852;
  assign n12305 = ~n12303 & n12304;
  assign n12306 = n7578 & ~n11724;
  assign po238 = ~n12305 & n12306;
  assign n12308 = ~po1038 & n10882;
  assign n12309 = pi68 & ~pi81;
  assign n12310 = n2479 & n12309;
  assign n12311 = n10614 & n12310;
  assign n12312 = n11030 & n12311;
  assign n12313 = n2799 & n12312;
  assign n12314 = pi81 & ~pi314;
  assign n12315 = n2491 & n12314;
  assign n12316 = ~n12313 & ~n12315;
  assign po239 = n12308 & ~n12316;
  assign n12318 = pi69 & pi314;
  assign n12319 = n2790 & n12318;
  assign n12320 = pi66 & ~pi73;
  assign n12321 = n2792 & n12320;
  assign n12322 = n2480 & n12321;
  assign n12323 = n2476 & n12322;
  assign n12324 = ~n12319 & ~n12323;
  assign n12325 = n10705 & n10707;
  assign po240 = ~n12324 & n12325;
  assign n12327 = n8648 & n10706;
  assign n12328 = n2479 & n2798;
  assign n12329 = ~pi68 & pi84;
  assign n12330 = n2792 & n12329;
  assign n12331 = n12328 & n12330;
  assign n12332 = n9878 & n12331;
  assign n12333 = n12327 & n12332;
  assign n12334 = pi314 & ~n12333;
  assign n12335 = ~pi83 & ~n12331;
  assign n12336 = n2795 & n12327;
  assign n12337 = ~n12335 & n12336;
  assign n12338 = ~pi314 & ~n12337;
  assign n12339 = n9782 & ~n12334;
  assign po241 = ~n12338 & n12339;
  assign n12341 = ~pi299 & n10421;
  assign n12342 = ~pi211 & pi299;
  assign n12343 = ~pi219 & n12342;
  assign n12344 = ~n12341 & ~n12343;
  assign n12345 = ~po1038 & ~n12344;
  assign po242 = n10971 & n12345;
  assign n12347 = n6383 & n10708;
  assign n12348 = ~pi314 & n10709;
  assign n12349 = n11028 & n12348;
  assign n12350 = ~n12347 & ~n12349;
  assign po243 = n10705 & ~n12350;
  assign n12352 = n7543 & n10982;
  assign n12353 = n7546 & n10985;
  assign n12354 = ~n12352 & ~n12353;
  assign po244 = n10585 & ~n12354;
  assign n12356 = pi314 & n9782;
  assign n12357 = n2703 & n10706;
  assign n12358 = n2844 & n12357;
  assign n12359 = n2707 & n12356;
  assign po245 = n12358 & n12359;
  assign n12361 = ~pi1093 & n2577;
  assign n12362 = n10644 & n12361;
  assign n12363 = n11051 & n12362;
  assign n12364 = ~n7356 & ~n12363;
  assign n12365 = n7348 & n10630;
  assign n12366 = ~pi1093 & ~n12365;
  assign n12367 = n2706 & n10644;
  assign n12368 = n7370 & n11858;
  assign n12369 = n10627 & n12368;
  assign n12370 = ~pi110 & n12367;
  assign n12371 = n12369 & n12370;
  assign n12372 = pi1093 & ~n12371;
  assign n12373 = n2577 & ~n6179;
  assign n12374 = ~n12372 & n12373;
  assign n12375 = ~n12366 & n12374;
  assign n12376 = n7356 & ~n12375;
  assign n12377 = ~po1038 & ~n12364;
  assign po246 = ~n12376 & n12377;
  assign n12379 = n9810 & n10940;
  assign n12380 = pi841 & n7377;
  assign n12381 = n12379 & n12380;
  assign n12382 = ~pi24 & pi70;
  assign n12383 = n2517 & n12382;
  assign n12384 = ~n12381 & ~n12383;
  assign n12385 = n9781 & n11856;
  assign po247 = ~n12384 & n12385;
  assign n12387 = ~pi1050 & n8782;
  assign n12388 = ~pi90 & ~n12387;
  assign n12389 = n10912 & ~n12388;
  assign n12390 = n2898 & n12389;
  assign po248 = ~n7364 & n12390;
  assign n12392 = ~n6418 & ~n9796;
  assign n12393 = n2926 & n9778;
  assign n12394 = ~n12392 & n12393;
  assign n12395 = pi24 & n2931;
  assign n12396 = ~n2926 & n12395;
  assign n12397 = n10688 & n12396;
  assign n12398 = n2756 & n12397;
  assign n12399 = ~pi39 & ~n12398;
  assign n12400 = ~n12394 & n12399;
  assign n12401 = n9830 & ~n12400;
  assign po249 = n7552 & n12401;
  assign n12403 = n2533 & ~po1038;
  assign n12404 = pi92 & n2523;
  assign n12405 = n3353 & n11069;
  assign n12406 = n12404 & n12405;
  assign n12407 = n5966 & n6214;
  assign n12408 = n7543 & n12407;
  assign n12409 = n5783 & n6204;
  assign n12410 = n7546 & n12409;
  assign n12411 = ~n12408 & ~n12410;
  assign n12412 = n2535 & n10821;
  assign n12413 = ~n12411 & n12412;
  assign n12414 = ~n12406 & ~n12413;
  assign po250 = n12403 & ~n12414;
  assign n12416 = pi93 & n10688;
  assign n12417 = n2914 & n12416;
  assign n12418 = ~pi92 & ~n12417;
  assign n12419 = ~pi1050 & n2523;
  assign n12420 = pi92 & ~n12419;
  assign n12421 = n3353 & n12403;
  assign n12422 = ~n12418 & n12421;
  assign po251 = ~n12420 & n12422;
  assign n12424 = n10670 & n10871;
  assign n12425 = pi252 & n8600;
  assign n12426 = n12424 & ~n12425;
  assign n12427 = n8600 & n10682;
  assign n12428 = ~n12424 & ~n12427;
  assign n12429 = n2717 & n9778;
  assign n12430 = n9897 & n10668;
  assign n12431 = ~n2777 & ~n12430;
  assign n12432 = ~n12428 & n12429;
  assign n12433 = ~n12431 & n12432;
  assign n12434 = ~n6175 & n12424;
  assign n12435 = ~pi1093 & ~po840;
  assign n12436 = ~n12434 & ~n12435;
  assign n12437 = n8600 & n11104;
  assign n12438 = ~n12436 & n12437;
  assign n12439 = ~n12426 & ~n12438;
  assign n12440 = ~n12433 & n12439;
  assign po252 = n9781 & ~n12440;
  assign n12442 = ~n6349 & ~n11018;
  assign n12443 = pi39 & ~n12442;
  assign n12444 = n9826 & n11355;
  assign n12445 = ~pi332 & n9778;
  assign n12446 = n10870 & n12445;
  assign n12447 = n12379 & n12446;
  assign n12448 = ~pi39 & ~n12447;
  assign n12449 = ~n12444 & n12448;
  assign n12450 = n9833 & ~n12449;
  assign po253 = ~n12443 & n12450;
  assign n12452 = pi479 & ~po840;
  assign n12453 = n3164 & n12452;
  assign n12454 = pi96 & pi841;
  assign n12455 = n2508 & n12454;
  assign n12456 = n3163 & n12455;
  assign n12457 = ~n12452 & n12456;
  assign n12458 = n2965 & n12457;
  assign n12459 = ~n12453 & ~n12458;
  assign n12460 = ~pi95 & ~n12459;
  assign n12461 = n2701 & n11355;
  assign n12462 = n9958 & n12461;
  assign n12463 = ~n12460 & ~n12462;
  assign po254 = n9781 & ~n12463;
  assign n12465 = pi39 & n11011;
  assign n12466 = pi593 & n11018;
  assign n12467 = n12465 & n12466;
  assign n12468 = ~n6349 & n12467;
  assign n12469 = ~n6150 & n12452;
  assign n12470 = ~po740 & ~n12469;
  assign n12471 = n2735 & n9824;
  assign n12472 = ~n12470 & n12471;
  assign n12473 = n11075 & n12472;
  assign n12474 = ~n12468 & ~n12473;
  assign po255 = n9833 & ~n12474;
  assign n12476 = ~pi92 & n11070;
  assign n12477 = ~n12404 & ~n12476;
  assign n12478 = pi314 & pi1050;
  assign n12479 = n12421 & n12478;
  assign po256 = ~n12477 & n12479;
  assign n12481 = ~pi72 & pi152;
  assign n12482 = n9932 & n12481;
  assign n12483 = pi299 & n12482;
  assign n12484 = ~pi72 & n9928;
  assign n12485 = n9930 & n12484;
  assign n12486 = ~n12483 & ~n12485;
  assign n12487 = pi232 & ~n12486;
  assign n12488 = pi39 & ~n12487;
  assign n12489 = ~pi72 & pi99;
  assign n12490 = ~pi39 & ~n12489;
  assign n12491 = ~n12488 & ~n12490;
  assign n12492 = ~n2574 & n12491;
  assign n12493 = ~n7440 & ~n12489;
  assign n12494 = ~n2922 & n12489;
  assign n12495 = n7440 & ~n12494;
  assign n12496 = ~n9962 & n12489;
  assign n12497 = n6092 & n10524;
  assign n12498 = ~n12496 & ~n12497;
  assign n12499 = n9992 & ~n12498;
  assign n12500 = n12495 & ~n12499;
  assign n12501 = ~n12493 & ~n12500;
  assign n12502 = ~pi39 & ~n12501;
  assign n12503 = n2574 & ~n12488;
  assign n12504 = ~n12502 & n12503;
  assign n12505 = pi75 & ~n12492;
  assign n12506 = ~n12504 & n12505;
  assign n12507 = ~n2532 & ~n12491;
  assign n12508 = pi228 & n10122;
  assign n12509 = pi228 & n9977;
  assign n12510 = n12489 & ~n12509;
  assign n12511 = n2532 & ~n12508;
  assign n12512 = ~n12510 & n12511;
  assign n12513 = pi87 & ~n12507;
  assign n12514 = ~n12512 & n12513;
  assign n12515 = n8738 & ~n12486;
  assign n12516 = ~n10542 & n12515;
  assign n12517 = pi41 & pi72;
  assign n12518 = pi99 & ~n12517;
  assign n12519 = ~n10042 & n12518;
  assign n12520 = ~pi228 & ~n10175;
  assign n12521 = ~n12519 & n12520;
  assign n12522 = ~n10075 & n12518;
  assign n12523 = n10385 & ~n12522;
  assign n12524 = ~n10054 & n12518;
  assign n12525 = n10383 & ~n12524;
  assign n12526 = ~n12523 & ~n12525;
  assign n12527 = pi228 & ~n12526;
  assign n12528 = ~pi39 & ~n12521;
  assign n12529 = ~n12527 & n12528;
  assign n12530 = n2613 & ~n12516;
  assign n12531 = ~n12529 & n12530;
  assign n12532 = pi38 & ~n12491;
  assign n12533 = ~n9989 & n12489;
  assign n12534 = n6091 & n9951;
  assign n12535 = ~n12533 & ~n12534;
  assign n12536 = n9992 & ~n12535;
  assign n12537 = n12495 & ~n12536;
  assign n12538 = ~pi39 & ~n12493;
  assign n12539 = ~n12537 & n12538;
  assign n12540 = n6082 & ~n12515;
  assign n12541 = ~n12539 & n12540;
  assign n12542 = ~pi87 & ~n12532;
  assign n12543 = ~n12541 & n12542;
  assign n12544 = ~n12531 & n12543;
  assign n12545 = ~pi75 & ~n12514;
  assign n12546 = ~n12544 & n12545;
  assign n12547 = ~n12506 & ~n12546;
  assign n12548 = n7360 & ~n12547;
  assign n12549 = ~n7360 & ~n12491;
  assign n12550 = ~po1038 & ~n12549;
  assign n12551 = ~n12548 & n12550;
  assign n12552 = pi232 & n12482;
  assign n12553 = pi39 & ~n12552;
  assign n12554 = po1038 & ~n12490;
  assign n12555 = ~n12553 & n12554;
  assign po257 = n12551 | n12555;
  assign n12557 = pi129 & ~n9715;
  assign n12558 = ~n6090 & ~n12557;
  assign n12559 = ~n6110 & ~n12558;
  assign n12560 = ~pi75 & n2614;
  assign n12561 = n6082 & n12560;
  assign n12562 = ~n12559 & n12561;
  assign n12563 = po840 & n9761;
  assign n12564 = ~n8601 & n12563;
  assign n12565 = ~n12562 & ~n12564;
  assign n12566 = n8598 & ~n12565;
  assign po258 = n2523 & n12566;
  assign n12568 = ~pi72 & ~pi144;
  assign n12569 = pi174 & n12568;
  assign n12570 = n9927 & n12569;
  assign n12571 = ~pi299 & ~n12570;
  assign n12572 = n3366 & n6166;
  assign n12573 = n12481 & n12572;
  assign n12574 = pi299 & ~n12573;
  assign n12575 = pi232 & ~n12571;
  assign n12576 = ~n12574 & n12575;
  assign n12577 = pi39 & ~n12576;
  assign n12578 = ~pi39 & ~n9955;
  assign n12579 = ~n12577 & ~n12578;
  assign n12580 = ~n7360 & ~n12579;
  assign n12581 = ~n2574 & n12579;
  assign n12582 = ~n7440 & ~n9955;
  assign n12583 = ~n2922 & n9955;
  assign n12584 = n7440 & ~n12583;
  assign n12585 = n2922 & ~n6099;
  assign n12586 = n9955 & ~n9961;
  assign n12587 = ~n9952 & ~n12586;
  assign n12588 = n12585 & ~n12587;
  assign n12589 = n12584 & ~n12588;
  assign n12590 = ~n12582 & ~n12589;
  assign n12591 = ~pi39 & ~n12590;
  assign n12592 = n2574 & ~n12577;
  assign n12593 = ~n12591 & n12592;
  assign n12594 = pi75 & ~n12581;
  assign n12595 = ~n12593 & n12594;
  assign n12596 = n9976 & n10534;
  assign n12597 = n9955 & ~n12596;
  assign n12598 = ~pi101 & n10535;
  assign n12599 = ~pi39 & ~n12597;
  assign n12600 = ~n12598 & n12599;
  assign n12601 = pi87 & ~n12577;
  assign n12602 = ~n12600 & n12601;
  assign n12603 = pi38 & ~n12579;
  assign n12604 = pi39 & n12576;
  assign n12605 = n7411 & n9976;
  assign n12606 = n9955 & ~n12605;
  assign n12607 = ~n9951 & ~n12606;
  assign n12608 = n12585 & ~n12607;
  assign n12609 = n12584 & ~n12608;
  assign n12610 = ~pi39 & ~n12582;
  assign n12611 = ~n12609 & n12610;
  assign n12612 = n6082 & ~n12604;
  assign n12613 = ~n12611 & n12612;
  assign n12614 = ~n10542 & n12604;
  assign n12615 = pi101 & ~n10040;
  assign n12616 = ~pi228 & ~n12615;
  assign n12617 = ~n10033 & n12616;
  assign n12618 = ~n10547 & ~n10551;
  assign n12619 = ~pi101 & ~n12618;
  assign n12620 = ~pi72 & n2922;
  assign n12621 = ~n10071 & n12620;
  assign n12622 = ~n2922 & ~n10052;
  assign n12623 = pi101 & ~n12622;
  assign n12624 = ~n12621 & n12623;
  assign n12625 = ~n12619 & ~n12624;
  assign n12626 = pi228 & ~n12625;
  assign n12627 = ~pi39 & ~n12617;
  assign n12628 = ~n12626 & n12627;
  assign n12629 = n2613 & ~n12614;
  assign n12630 = ~n12628 & n12629;
  assign n12631 = ~pi87 & ~n12603;
  assign n12632 = ~n12613 & n12631;
  assign n12633 = ~n12630 & n12632;
  assign n12634 = ~pi75 & ~n12602;
  assign n12635 = ~n12633 & n12634;
  assign n12636 = ~n12595 & ~n12635;
  assign n12637 = n7360 & ~n12636;
  assign n12638 = ~po1038 & ~n12580;
  assign n12639 = ~n12637 & n12638;
  assign n12640 = pi232 & n12573;
  assign n12641 = pi39 & ~n12640;
  assign n12642 = po1038 & ~n12578;
  assign n12643 = ~n12641 & n12642;
  assign po259 = n12639 | n12643;
  assign n12645 = n2854 & n8626;
  assign po260 = n12308 & n12645;
  assign n12647 = pi109 & n2765;
  assign n12648 = n2704 & n12647;
  assign n12649 = pi314 & ~n12648;
  assign n12650 = ~pi109 & ~n12358;
  assign n12651 = n6373 & ~n12650;
  assign n12652 = ~pi314 & ~n12651;
  assign n12653 = n10704 & ~n12649;
  assign po261 = ~n12652 & n12653;
  assign n12655 = n7356 & ~n8600;
  assign n12656 = n9710 & ~n12655;
  assign n12657 = n10028 & ~n12656;
  assign n12658 = ~pi110 & ~n12369;
  assign n12659 = n12367 & ~n12658;
  assign n12660 = ~n2759 & n12659;
  assign n12661 = ~n8600 & ~n12660;
  assign n12662 = n8600 & ~n12371;
  assign n12663 = ~n6179 & ~n7356;
  assign n12664 = ~n12662 & n12663;
  assign n12665 = ~n12661 & n12664;
  assign n12666 = ~n12657 & ~n12665;
  assign po262 = n9781 & ~n12666;
  assign n12668 = pi24 & n10869;
  assign n12669 = ~pi53 & ~n10868;
  assign n12670 = n2723 & ~n12669;
  assign n12671 = ~pi24 & n2717;
  assign n12672 = n12670 & n12671;
  assign n12673 = ~n12668 & ~n12672;
  assign n12674 = pi841 & ~n12673;
  assign n12675 = n8655 & n10854;
  assign n12676 = ~n12674 & ~n12675;
  assign po264 = n9782 & ~n12676;
  assign n12678 = ~pi999 & n9782;
  assign po265 = n10941 & n12678;
  assign n12680 = pi314 & ~n7375;
  assign n12681 = ~pi97 & n7373;
  assign n12682 = ~pi108 & ~n12681;
  assign n12683 = n2706 & ~n12682;
  assign n12684 = n9895 & n12683;
  assign n12685 = ~pi314 & ~n12684;
  assign n12686 = n7377 & ~n9872;
  assign n12687 = ~n12680 & n12686;
  assign n12688 = ~n12685 & n12687;
  assign n12689 = n7377 & n9872;
  assign n12690 = n12684 & n12689;
  assign n12691 = ~pi51 & ~n12690;
  assign n12692 = ~n12688 & n12691;
  assign n12693 = n2532 & n7380;
  assign n12694 = ~n12692 & n12693;
  assign n12695 = ~pi87 & ~n12694;
  assign n12696 = n6080 & n8598;
  assign po266 = ~n12695 & n12696;
  assign n12698 = n2782 & n11033;
  assign po267 = n12356 & n12698;
  assign n12700 = ~pi82 & pi111;
  assign n12701 = n8648 & n12700;
  assign n12702 = n10709 & n12701;
  assign n12703 = n2800 & n12702;
  assign n12704 = pi314 & n12703;
  assign n12705 = n8600 & n9710;
  assign n12706 = n10010 & n12705;
  assign n12707 = ~n12704 & ~n12706;
  assign po268 = n9782 & ~n12707;
  assign n12709 = pi72 & n9958;
  assign n12710 = ~pi314 & n12703;
  assign n12711 = n8623 & n12710;
  assign n12712 = ~n12709 & ~n12711;
  assign n12713 = n6431 & n9781;
  assign po269 = ~n12712 & n12713;
  assign po270 = ~pi124 | pi468;
  assign n12716 = ~pi39 & n10182;
  assign n12717 = pi38 & ~n12716;
  assign n12718 = n7411 & n10141;
  assign n12719 = ~n6098 & ~n12718;
  assign n12720 = n10733 & ~n12719;
  assign n12721 = n10182 & ~n12720;
  assign n12722 = ~n6098 & n10733;
  assign n12723 = n10192 & n12722;
  assign n12724 = n9951 & n12723;
  assign n12725 = ~n12721 & ~n12724;
  assign n12726 = ~pi39 & ~n12725;
  assign n12727 = n6082 & ~n12726;
  assign n12728 = ~pi113 & n10175;
  assign n12729 = pi113 & n10181;
  assign n12730 = ~pi228 & ~n12728;
  assign n12731 = ~n12729 & n12730;
  assign n12732 = pi113 & ~n10179;
  assign n12733 = ~n10395 & n12732;
  assign n12734 = pi228 & ~n10387;
  assign n12735 = ~n12733 & n12734;
  assign n12736 = ~pi39 & ~n12731;
  assign n12737 = ~n12735 & n12736;
  assign n12738 = n2613 & ~n12737;
  assign n12739 = ~n12717 & ~n12727;
  assign n12740 = ~n12738 & n12739;
  assign n12741 = ~pi87 & ~n12740;
  assign n12742 = ~n2613 & n12716;
  assign n12743 = ~n10142 & n10182;
  assign n12744 = ~pi113 & n12508;
  assign n12745 = ~n12743 & ~n12744;
  assign n12746 = n2532 & ~n12745;
  assign n12747 = pi87 & ~n12742;
  assign n12748 = ~n12746 & n12747;
  assign n12749 = ~n12741 & ~n12748;
  assign n12750 = ~pi75 & ~n12749;
  assign n12751 = n7414 & n12724;
  assign n12752 = ~n6098 & ~n10118;
  assign n12753 = n10733 & ~n12752;
  assign n12754 = n10182 & ~n12753;
  assign n12755 = ~n12751 & ~n12754;
  assign n12756 = n2615 & ~n12755;
  assign n12757 = ~n2574 & n12716;
  assign n12758 = pi75 & ~n12757;
  assign n12759 = ~n12756 & n12758;
  assign n12760 = ~n12750 & ~n12759;
  assign n12761 = n8598 & ~n12760;
  assign n12762 = ~n8598 & ~n12716;
  assign po271 = ~n12761 & ~n12762;
  assign n12764 = ~pi72 & pi114;
  assign n12765 = ~pi39 & n12764;
  assign n12766 = ~n2574 & n12765;
  assign n12767 = n7440 & n10113;
  assign n12768 = ~n12764 & ~n12767;
  assign n12769 = n7414 & n10126;
  assign n12770 = pi114 & n10344;
  assign n12771 = n12767 & ~n12769;
  assign n12772 = ~n12770 & n12771;
  assign n12773 = n2615 & ~n12768;
  assign n12774 = ~n12772 & n12773;
  assign n12775 = pi75 & ~n12766;
  assign n12776 = ~n12774 & n12775;
  assign n12777 = ~n2613 & ~n12765;
  assign n12778 = ~pi115 & n10363;
  assign n12779 = n12764 & ~n12778;
  assign n12780 = pi228 & n10123;
  assign n12781 = ~pi115 & n12780;
  assign n12782 = ~pi114 & n12781;
  assign n12783 = n2613 & ~n12779;
  assign n12784 = ~n12782 & n12783;
  assign n12785 = n10822 & ~n12777;
  assign n12786 = ~n12784 & n12785;
  assign n12787 = pi38 & ~n12765;
  assign n12788 = ~n10735 & n12764;
  assign n12789 = n12767 & ~n12788;
  assign n12790 = ~n10126 & n12789;
  assign n12791 = ~pi39 & ~n12768;
  assign n12792 = ~n12790 & n12791;
  assign n12793 = n6082 & ~n12792;
  assign n12794 = pi114 & ~n10400;
  assign n12795 = ~pi114 & ~n10390;
  assign n12796 = ~n12794 & ~n12795;
  assign n12797 = ~pi115 & ~n12796;
  assign n12798 = pi115 & ~n12764;
  assign n12799 = ~pi39 & ~n12798;
  assign n12800 = ~n12797 & n12799;
  assign n12801 = n2613 & ~n12800;
  assign n12802 = ~pi87 & ~n12787;
  assign n12803 = ~n12793 & n12802;
  assign n12804 = ~n12801 & n12803;
  assign n12805 = ~pi75 & ~n12786;
  assign n12806 = ~n12804 & n12805;
  assign n12807 = ~n12776 & ~n12806;
  assign n12808 = n8598 & ~n12807;
  assign n12809 = ~n8598 & ~n12765;
  assign po272 = ~n12808 & ~n12809;
  assign n12811 = ~pi72 & pi115;
  assign n12812 = ~pi39 & n12811;
  assign n12813 = ~n2574 & n12812;
  assign n12814 = ~n10733 & ~n12811;
  assign n12815 = pi115 & n10344;
  assign n12816 = ~pi114 & n6094;
  assign n12817 = ~pi115 & ~n12816;
  assign n12818 = n10124 & n12817;
  assign n12819 = n7414 & n12818;
  assign n12820 = n10733 & ~n12815;
  assign n12821 = ~n12819 & n12820;
  assign n12822 = n2615 & ~n12814;
  assign n12823 = ~n12821 & n12822;
  assign n12824 = pi75 & ~n12813;
  assign n12825 = ~n12823 & n12824;
  assign n12826 = ~n2613 & ~n12812;
  assign n12827 = ~n10363 & n12811;
  assign n12828 = n2613 & ~n12827;
  assign n12829 = ~n12781 & n12828;
  assign n12830 = n10822 & ~n12826;
  assign n12831 = ~n12829 & n12830;
  assign n12832 = pi38 & ~n12812;
  assign n12833 = ~n10735 & n12811;
  assign n12834 = n10733 & ~n12833;
  assign n12835 = ~n12818 & n12834;
  assign n12836 = ~pi39 & ~n12814;
  assign n12837 = ~n12835 & n12836;
  assign n12838 = n6082 & ~n12837;
  assign n12839 = pi115 & ~n10400;
  assign n12840 = ~pi115 & ~n10390;
  assign n12841 = ~pi39 & ~n12840;
  assign n12842 = ~n12839 & n12841;
  assign n12843 = n2613 & ~n12842;
  assign n12844 = ~pi87 & ~n12832;
  assign n12845 = ~n12838 & n12844;
  assign n12846 = ~n12843 & n12845;
  assign n12847 = ~pi75 & ~n12831;
  assign n12848 = ~n12846 & n12847;
  assign n12849 = ~n12825 & ~n12848;
  assign n12850 = n8598 & ~n12849;
  assign n12851 = ~n8598 & ~n12812;
  assign po273 = ~n12850 & ~n12851;
  assign n12853 = n10178 & ~n10733;
  assign n12854 = ~n10119 & n10178;
  assign n12855 = ~n10347 & ~n12854;
  assign n12856 = n12722 & ~n12855;
  assign n12857 = ~n12853 & ~n12856;
  assign n12858 = n2615 & ~n12857;
  assign n12859 = ~pi39 & n10178;
  assign n12860 = ~n2574 & n12859;
  assign n12861 = pi75 & ~n12860;
  assign n12862 = ~n12858 & n12861;
  assign n12863 = pi38 & ~n12859;
  assign n12864 = ~pi38 & ~pi113;
  assign n12865 = n10142 & n12864;
  assign n12866 = n10178 & ~n12865;
  assign n12867 = ~n12780 & ~n12866;
  assign n12868 = ~n12863 & ~n12867;
  assign n12869 = ~pi100 & ~n12868;
  assign n12870 = pi100 & ~n12859;
  assign n12871 = n10822 & ~n12870;
  assign n12872 = ~n12869 & n12871;
  assign n12873 = ~pi113 & n12718;
  assign n12874 = n10178 & ~n12873;
  assign n12875 = ~n10124 & ~n12874;
  assign n12876 = n12722 & ~n12875;
  assign n12877 = ~n12853 & ~n12876;
  assign n12878 = ~pi39 & ~n12877;
  assign n12879 = n6082 & ~n12878;
  assign n12880 = ~n2922 & n10207;
  assign n12881 = n10178 & ~n10193;
  assign n12882 = ~n10194 & ~n12881;
  assign n12883 = n2922 & ~n12882;
  assign n12884 = pi116 & ~n2922;
  assign n12885 = n10203 & n12884;
  assign n12886 = pi228 & ~n12880;
  assign n12887 = ~n12885 & n12886;
  assign n12888 = ~n12883 & n12887;
  assign n12889 = pi116 & ~n10183;
  assign n12890 = n10382 & ~n12889;
  assign n12891 = ~pi39 & ~n12890;
  assign n12892 = ~n12888 & n12891;
  assign n12893 = n2613 & ~n12892;
  assign n12894 = ~pi87 & ~n12863;
  assign n12895 = ~n12879 & n12894;
  assign n12896 = ~n12893 & n12895;
  assign n12897 = ~pi75 & ~n12872;
  assign n12898 = ~n12896 & n12897;
  assign n12899 = ~n12862 & ~n12898;
  assign n12900 = n8598 & ~n12899;
  assign n12901 = ~n8598 & ~n12859;
  assign po274 = ~n12900 & ~n12901;
  assign n12903 = n3651 & n7310;
  assign n12904 = ~n3650 & ~n12903;
  assign n12905 = ~pi38 & ~n12904;
  assign n12906 = ~pi87 & ~n12905;
  assign n12907 = n6080 & ~n12906;
  assign n12908 = ~pi92 & ~n12907;
  assign n12909 = ~pi54 & ~n7234;
  assign n12910 = ~pi74 & n12909;
  assign n12911 = ~n12908 & n12910;
  assign n12912 = ~pi55 & ~n12911;
  assign n12913 = ~n7277 & ~n12912;
  assign n12914 = ~pi56 & ~n12913;
  assign n12915 = ~n6248 & ~n12914;
  assign n12916 = ~pi62 & ~n12915;
  assign n12917 = ~pi57 & n6253;
  assign po275 = ~n12916 & n12917;
  assign n12919 = ~pi79 & n11710;
  assign n12920 = pi163 & n6166;
  assign n12921 = ~n11267 & ~n12920;
  assign n12922 = ~pi150 & ~n12921;
  assign n12923 = pi150 & n9362;
  assign n12924 = n11265 & n12923;
  assign n12925 = ~n12922 & ~n12924;
  assign n12926 = n9366 & ~n12925;
  assign n12927 = pi74 & ~n12926;
  assign n12928 = ~pi74 & ~n12926;
  assign n12929 = pi165 & n7406;
  assign n12930 = ~n8704 & ~n12929;
  assign n12931 = n7231 & n12930;
  assign n12932 = n12928 & ~n12931;
  assign n12933 = ~n12927 & ~n12932;
  assign n12934 = ~n2530 & ~n12933;
  assign n12935 = n3291 & ~n12934;
  assign n12936 = ~n9532 & ~n12935;
  assign n12937 = pi55 & ~n12927;
  assign n12938 = pi150 & n7406;
  assign n12939 = ~pi92 & n8970;
  assign n12940 = n12938 & n12939;
  assign n12941 = n8704 & n8937;
  assign n12942 = ~n12940 & n12941;
  assign n12943 = ~n12930 & ~n12942;
  assign n12944 = n7231 & ~n12943;
  assign n12945 = n12928 & ~n12944;
  assign n12946 = n12937 & ~n12945;
  assign n12947 = ~pi184 & ~n11293;
  assign n12948 = pi185 & ~n12947;
  assign n12949 = ~pi185 & n12947;
  assign n12950 = n6166 & ~n12948;
  assign n12951 = ~n12949 & n12950;
  assign n12952 = ~pi299 & ~n12951;
  assign n12953 = pi299 & n12925;
  assign n12954 = pi232 & ~n12952;
  assign n12955 = ~n12953 & n12954;
  assign n12956 = ~n7231 & n12955;
  assign n12957 = pi74 & ~n12956;
  assign n12958 = ~pi55 & ~n12957;
  assign n12959 = ~pi143 & ~pi299;
  assign n12960 = ~pi165 & pi299;
  assign n12961 = ~n12959 & ~n12960;
  assign n12962 = n7406 & n12961;
  assign n12963 = n7231 & ~n12962;
  assign n12964 = pi54 & ~n12963;
  assign n12965 = ~n12956 & n12964;
  assign n12966 = pi75 & ~n12955;
  assign n12967 = pi100 & ~n12955;
  assign n12968 = pi38 & ~n12962;
  assign n12969 = ~pi100 & ~n12968;
  assign n12970 = ~pi157 & pi299;
  assign n12971 = ~pi178 & ~pi299;
  assign n12972 = ~n12970 & ~n12971;
  assign n12973 = n7406 & n12972;
  assign n12974 = n8970 & n12973;
  assign n12975 = n8938 & ~n12974;
  assign n12976 = n12969 & ~n12975;
  assign n12977 = ~n12967 & ~n12976;
  assign n12978 = n8890 & ~n12977;
  assign n12979 = ~pi143 & ~n8872;
  assign n12980 = pi143 & ~n8874;
  assign n12981 = pi165 & ~n12980;
  assign n12982 = ~n12979 & n12981;
  assign n12983 = pi143 & ~pi165;
  assign n12984 = n8879 & n12983;
  assign n12985 = pi38 & ~n12984;
  assign n12986 = ~n12982 & n12985;
  assign n12987 = n2573 & ~n12986;
  assign n12988 = ~pi232 & n9249;
  assign n12989 = pi168 & n6166;
  assign n12990 = n9249 & ~n12989;
  assign n12991 = pi168 & n9234;
  assign n12992 = ~pi151 & ~n12990;
  assign n12993 = ~n12991 & n12992;
  assign n12994 = ~n6166 & n9249;
  assign n12995 = n6166 & n9636;
  assign n12996 = ~n12994 & ~n12995;
  assign n12997 = ~pi168 & ~n12996;
  assign n12998 = ~n6166 & ~n9249;
  assign n12999 = ~n9288 & ~n12998;
  assign n13000 = pi168 & n12999;
  assign n13001 = pi151 & ~n12997;
  assign n13002 = ~n13000 & n13001;
  assign n13003 = ~pi150 & ~n12993;
  assign n13004 = ~n13002 & n13003;
  assign n13005 = n6166 & ~n9073;
  assign n13006 = ~n12998 & ~n13005;
  assign n13007 = pi151 & pi168;
  assign n13008 = ~n13006 & n13007;
  assign n13009 = ~pi168 & n9210;
  assign n13010 = pi168 & n9214;
  assign n13011 = ~pi151 & ~n13009;
  assign n13012 = ~n13010 & n13011;
  assign n13013 = pi151 & ~pi168;
  assign n13014 = ~n9220 & n13013;
  assign n13015 = ~n13012 & ~n13014;
  assign n13016 = ~n12994 & ~n13015;
  assign n13017 = pi150 & ~n13008;
  assign n13018 = ~n13016 & n13017;
  assign n13019 = pi299 & ~n13004;
  assign n13020 = ~n13018 & n13019;
  assign n13021 = pi173 & ~n12999;
  assign n13022 = ~pi173 & ~n9234;
  assign n13023 = ~n12994 & n13022;
  assign n13024 = ~n13021 & ~n13023;
  assign n13025 = ~pi185 & ~n13024;
  assign n13026 = n6166 & ~n9231;
  assign n13027 = pi173 & ~n12998;
  assign n13028 = ~n13026 & n13027;
  assign n13029 = ~n9240 & ~n12994;
  assign n13030 = ~pi173 & ~n13029;
  assign n13031 = pi185 & ~n13028;
  assign n13032 = ~n13030 & n13031;
  assign n13033 = pi190 & ~n13025;
  assign n13034 = ~n13032 & n13033;
  assign n13035 = pi173 & ~n12996;
  assign n13036 = ~pi173 & n9249;
  assign n13037 = ~pi185 & ~n13036;
  assign n13038 = ~n13035 & n13037;
  assign n13039 = ~pi173 & n9246;
  assign n13040 = pi173 & n9634;
  assign n13041 = ~n13039 & ~n13040;
  assign n13042 = n6166 & ~n13041;
  assign n13043 = pi185 & ~n12994;
  assign n13044 = ~n13042 & n13043;
  assign n13045 = ~pi190 & ~n13038;
  assign n13046 = ~n13044 & n13045;
  assign n13047 = ~pi299 & ~n13046;
  assign n13048 = ~n13034 & n13047;
  assign n13049 = pi232 & ~n13048;
  assign n13050 = ~n13020 & n13049;
  assign n13051 = ~pi39 & ~n12988;
  assign n13052 = ~n13050 & n13051;
  assign n13053 = ~pi232 & n8937;
  assign n13054 = pi168 & n8999;
  assign n13055 = pi157 & n9006;
  assign n13056 = ~n13054 & ~n13055;
  assign n13057 = pi299 & n8739;
  assign n13058 = n6222 & n13057;
  assign n13059 = ~n13056 & n13058;
  assign n13060 = pi178 & ~pi190;
  assign n13061 = n9016 & n13060;
  assign n13062 = ~pi178 & ~n8981;
  assign n13063 = pi190 & ~n6194;
  assign n13064 = ~n13062 & n13063;
  assign n13065 = n8986 & n13064;
  assign n13066 = ~n13061 & ~n13065;
  assign n13067 = ~pi299 & n8752;
  assign n13068 = ~n13066 & n13067;
  assign n13069 = pi232 & n8937;
  assign n13070 = ~n13059 & n13069;
  assign n13071 = ~n13068 & n13070;
  assign n13072 = pi39 & ~n13053;
  assign n13073 = ~n13071 & n13072;
  assign n13074 = ~pi38 & ~n13073;
  assign n13075 = ~n13052 & n13074;
  assign n13076 = n12987 & ~n13075;
  assign n13077 = pi87 & n12969;
  assign n13078 = ~n8938 & n13077;
  assign n13079 = ~n12967 & ~n13078;
  assign n13080 = ~n13076 & n13079;
  assign n13081 = n2572 & ~n13080;
  assign n13082 = ~n12966 & ~n12978;
  assign n13083 = ~n13081 & n13082;
  assign n13084 = ~pi54 & ~n13083;
  assign n13085 = ~n12965 & ~n13084;
  assign n13086 = ~pi74 & ~n13085;
  assign n13087 = n12958 & ~n13086;
  assign n13088 = n2530 & ~n12946;
  assign n13089 = ~n13087 & n13088;
  assign n13090 = ~n12936 & ~n13089;
  assign n13091 = ~pi74 & n7231;
  assign n13092 = ~n12929 & n13091;
  assign n13093 = ~n12926 & ~n13092;
  assign n13094 = ~n3291 & ~n13093;
  assign n13095 = ~n13090 & ~n13094;
  assign n13096 = pi118 & n13095;
  assign n13097 = n8669 & ~n12973;
  assign n13098 = n2523 & n13097;
  assign n13099 = n12969 & ~n13098;
  assign n13100 = ~n12967 & ~n13099;
  assign n13101 = n8890 & ~n13100;
  assign n13102 = n7257 & n8739;
  assign n13103 = n5783 & n6208;
  assign n13104 = ~n13102 & ~n13103;
  assign n13105 = ~n6349 & ~n13104;
  assign n13106 = ~pi232 & ~n13105;
  assign n13107 = ~pi157 & ~n8742;
  assign n13108 = pi157 & ~n8740;
  assign n13109 = ~pi168 & ~n13108;
  assign n13110 = ~n13107 & n13109;
  assign n13111 = n6205 & ~n6349;
  assign n13112 = ~pi157 & pi168;
  assign n13113 = n8746 & n13112;
  assign n13114 = ~n13111 & ~n13113;
  assign n13115 = ~n13110 & n13114;
  assign n13116 = n12407 & ~n13115;
  assign n13117 = ~pi178 & n6349;
  assign n13118 = pi178 & ~n6341;
  assign n13119 = ~pi190 & ~n13118;
  assign n13120 = ~n13117 & n13119;
  assign n13121 = ~pi178 & pi190;
  assign n13122 = n7542 & n13121;
  assign n13123 = ~n13120 & ~n13122;
  assign n13124 = n6206 & ~n13123;
  assign n13125 = ~n13111 & ~n13124;
  assign n13126 = n12409 & ~n13125;
  assign n13127 = pi232 & ~n13116;
  assign n13128 = ~n13126 & n13127;
  assign n13129 = pi39 & ~n13106;
  assign n13130 = ~n13128 & n13129;
  assign n13131 = n6150 & n6439;
  assign n13132 = ~pi232 & ~n13131;
  assign n13133 = ~n8826 & n13132;
  assign n13134 = ~pi151 & n8793;
  assign n13135 = ~pi168 & n8783;
  assign n13136 = ~n13134 & ~n13135;
  assign n13137 = n8788 & ~n13136;
  assign n13138 = pi150 & ~n13137;
  assign n13139 = ~pi151 & n8808;
  assign n13140 = n8811 & ~n13139;
  assign n13141 = n12989 & ~n13140;
  assign n13142 = ~pi151 & n8826;
  assign n13143 = n8829 & ~n13142;
  assign n13144 = ~pi168 & ~n13143;
  assign n13145 = ~pi150 & ~n13141;
  assign n13146 = ~n13144 & n13145;
  assign n13147 = ~n13138 & ~n13146;
  assign n13148 = ~n6440 & ~n8826;
  assign n13149 = ~n6166 & ~n13148;
  assign n13150 = ~n13147 & ~n13149;
  assign n13151 = pi299 & ~n13150;
  assign n13152 = ~n6166 & ~n8845;
  assign n13153 = pi173 & n8859;
  assign n13154 = pi190 & n8854;
  assign n13155 = ~n13153 & n13154;
  assign n13156 = ~pi173 & n8826;
  assign n13157 = n8840 & ~n13156;
  assign n13158 = ~pi190 & ~n13157;
  assign n13159 = ~pi185 & ~n13155;
  assign n13160 = ~n13158 & n13159;
  assign n13161 = pi173 & ~n8783;
  assign n13162 = ~pi190 & ~n13161;
  assign n13163 = ~n8847 & n13162;
  assign n13164 = ~pi173 & pi190;
  assign n13165 = n8794 & n13164;
  assign n13166 = pi185 & ~n13165;
  assign n13167 = ~n13163 & n13166;
  assign n13168 = ~n13160 & ~n13167;
  assign n13169 = ~n13152 & ~n13168;
  assign n13170 = ~pi299 & ~n13169;
  assign n13171 = pi232 & ~n13151;
  assign n13172 = ~n13170 & n13171;
  assign n13173 = ~pi39 & ~n13133;
  assign n13174 = ~n13172 & n13173;
  assign n13175 = ~n13130 & ~n13174;
  assign n13176 = ~pi38 & ~n13175;
  assign n13177 = n12987 & ~n13176;
  assign n13178 = ~n12967 & ~n13077;
  assign n13179 = ~n13177 & n13178;
  assign n13180 = n2572 & ~n13179;
  assign n13181 = ~n12966 & ~n13101;
  assign n13182 = ~n13180 & n13181;
  assign n13183 = ~pi54 & ~n13182;
  assign n13184 = ~n12965 & ~n13183;
  assign n13185 = ~pi74 & ~n13184;
  assign n13186 = n12958 & ~n13185;
  assign n13187 = pi54 & n12929;
  assign n13188 = ~pi92 & n3353;
  assign n13189 = ~n12938 & n13188;
  assign n13190 = ~n13187 & n13189;
  assign n13191 = n2523 & n13190;
  assign n13192 = n12932 & ~n13191;
  assign n13193 = n12937 & ~n13192;
  assign n13194 = n2530 & ~n13193;
  assign n13195 = ~n13186 & n13194;
  assign n13196 = n12935 & ~n13195;
  assign n13197 = ~n13094 & ~n13196;
  assign n13198 = ~pi118 & n13197;
  assign n13199 = ~n12919 & ~n13198;
  assign n13200 = ~n13096 & n13199;
  assign n13201 = ~pi118 & ~n8681;
  assign n13202 = n13197 & ~n13201;
  assign n13203 = n13095 & n13201;
  assign n13204 = n12919 & ~n13202;
  assign n13205 = ~n13203 & n13204;
  assign po276 = n13200 | n13205;
  assign n13207 = pi128 & pi228;
  assign n13208 = ~n12403 & n13207;
  assign n13209 = ~n7295 & ~n13207;
  assign n13210 = pi75 & ~n13209;
  assign n13211 = pi87 & ~n13207;
  assign n13212 = ~n7294 & ~n13207;
  assign n13213 = pi100 & ~n13212;
  assign n13214 = ~n2608 & n5783;
  assign n13215 = n7546 & n13214;
  assign n13216 = ~n3302 & n5966;
  assign n13217 = n7543 & n13216;
  assign n13218 = ~n13215 & ~n13217;
  assign n13219 = pi39 & ~n13218;
  assign n13220 = pi299 & n6371;
  assign n13221 = ~n6480 & ~n13220;
  assign n13222 = n7406 & ~n13221;
  assign n13223 = ~n6443 & n13222;
  assign n13224 = ~n6373 & ~n13222;
  assign n13225 = pi109 & ~n13222;
  assign n13226 = ~n2926 & n11254;
  assign n13227 = n9783 & n9795;
  assign n13228 = n11253 & ~n13227;
  assign n13229 = n2780 & ~n13228;
  assign n13230 = ~pi97 & ~n13229;
  assign n13231 = ~pi46 & n2926;
  assign n13232 = n2929 & n13231;
  assign n13233 = ~n13230 & n13232;
  assign n13234 = ~n13225 & ~n13226;
  assign n13235 = ~n13233 & n13234;
  assign n13236 = ~n13223 & ~n13224;
  assign n13237 = ~n13235 & n13236;
  assign n13238 = ~pi91 & ~n13237;
  assign n13239 = n2709 & ~n6419;
  assign n13240 = ~n13238 & n13239;
  assign n13241 = ~n2752 & ~n13240;
  assign n13242 = n2509 & n12471;
  assign n13243 = ~n13241 & n13242;
  assign n13244 = ~n13219 & ~n13243;
  assign n13245 = ~pi38 & ~n13244;
  assign n13246 = ~pi228 & n13245;
  assign n13247 = ~n13207 & ~n13246;
  assign n13248 = ~pi100 & ~n13247;
  assign n13249 = ~pi87 & ~n13213;
  assign n13250 = ~n13248 & n13249;
  assign n13251 = ~pi75 & ~n13211;
  assign n13252 = ~n13250 & n13251;
  assign n13253 = ~pi92 & ~n13210;
  assign n13254 = ~n13252 & n13253;
  assign n13255 = pi92 & ~n13207;
  assign n13256 = ~n7300 & n13255;
  assign n13257 = n12403 & ~n13256;
  assign n13258 = ~n13254 & n13257;
  assign po277 = n13208 | n13258;
  assign n13260 = ~pi31 & ~pi80;
  assign n13261 = pi818 & n13260;
  assign n13262 = n7351 & ~n7360;
  assign n13263 = ~n7356 & ~n13262;
  assign n13264 = ~pi120 & ~n7360;
  assign n13265 = ~pi1093 & n13264;
  assign n13266 = n13263 & ~n13265;
  assign n13267 = n2523 & n7531;
  assign n13268 = pi120 & ~n7351;
  assign n13269 = ~n7443 & n13268;
  assign n13270 = n13267 & ~n13269;
  assign n13271 = ~pi120 & pi1093;
  assign n13272 = n7443 & ~n13271;
  assign n13273 = ~n13270 & ~n13272;
  assign n13274 = n7536 & ~n13273;
  assign n13275 = ~pi120 & ~pi1093;
  assign n13276 = pi100 & ~n13275;
  assign n13277 = ~n7351 & n13276;
  assign n13278 = ~n13274 & n13277;
  assign n13279 = pi120 & n7397;
  assign n13280 = ~pi39 & ~n13279;
  assign n13281 = pi122 & n7396;
  assign n13282 = n7384 & n7418;
  assign n13283 = ~n13281 & ~n13282;
  assign n13284 = ~n10067 & n13283;
  assign n13285 = ~n2921 & ~n13284;
  assign n13286 = n6178 & ~n13285;
  assign n13287 = n7348 & n7381;
  assign n13288 = n7561 & ~n13287;
  assign n13289 = ~n7418 & n13288;
  assign n13290 = ~n13286 & ~n13289;
  assign n13291 = n13280 & n13290;
  assign n13292 = ~n7351 & ~n13275;
  assign n13293 = n6205 & n7542;
  assign n13294 = n13292 & ~n13293;
  assign n13295 = n6221 & n13294;
  assign n13296 = ~n6197 & n7542;
  assign n13297 = n13292 & ~n13296;
  assign n13298 = ~n6221 & n13297;
  assign n13299 = n5727 & ~n13295;
  assign n13300 = ~n13298 & n13299;
  assign n13301 = ~n5727 & ~n13292;
  assign n13302 = pi299 & ~n13301;
  assign n13303 = ~n13300 & n13302;
  assign n13304 = ~n7506 & ~n13292;
  assign n13305 = n6194 & n13294;
  assign n13306 = ~n6194 & n13297;
  assign n13307 = n7506 & ~n13305;
  assign n13308 = ~n13306 & n13307;
  assign n13309 = ~pi299 & ~n13304;
  assign n13310 = ~n13308 & n13309;
  assign n13311 = pi39 & ~n13303;
  assign n13312 = ~n13310 & n13311;
  assign n13313 = ~n13291 & ~n13312;
  assign n13314 = ~pi38 & ~n13313;
  assign n13315 = pi38 & n13275;
  assign n13316 = ~pi100 & ~n13315;
  assign n13317 = ~n7451 & n13316;
  assign n13318 = ~n13314 & n13317;
  assign n13319 = ~n13278 & ~n13318;
  assign n13320 = ~pi87 & ~n13319;
  assign n13321 = n7566 & ~n13275;
  assign n13322 = ~n2628 & n7351;
  assign n13323 = ~n7418 & n7561;
  assign n13324 = ~n7431 & n13323;
  assign n13325 = n7564 & ~n13324;
  assign n13326 = pi87 & ~n13322;
  assign n13327 = ~n13325 & n13326;
  assign n13328 = n13321 & n13327;
  assign n13329 = ~n13320 & ~n13328;
  assign n13330 = ~pi75 & ~n13329;
  assign n13331 = ~n7351 & n13271;
  assign n13332 = ~n7532 & n13331;
  assign n13333 = ~pi1091 & ~n7350;
  assign n13334 = ~n7416 & ~n13333;
  assign n13335 = pi120 & ~n13334;
  assign n13336 = ~n7407 & ~n13335;
  assign n13337 = ~n13332 & n13336;
  assign n13338 = n7407 & ~n13292;
  assign n13339 = ~n13337 & ~n13338;
  assign n13340 = n2615 & ~n13339;
  assign n13341 = ~n2615 & ~n13292;
  assign n13342 = pi75 & ~n13341;
  assign n13343 = ~n13340 & n13342;
  assign n13344 = n7360 & ~n13343;
  assign n13345 = ~n13330 & n13344;
  assign n13346 = n13266 & ~n13345;
  assign n13347 = n7535 & ~n13275;
  assign n13348 = ~n13286 & ~n13288;
  assign n13349 = n13280 & n13348;
  assign n13350 = pi299 & ~n13275;
  assign n13351 = ~n8460 & n13350;
  assign n13352 = ~pi299 & ~n13275;
  assign n13353 = ~n8467 & n13352;
  assign n13354 = pi39 & ~n13351;
  assign n13355 = ~n13353 & n13354;
  assign n13356 = ~n13349 & ~n13355;
  assign n13357 = ~pi38 & ~n13356;
  assign n13358 = n13316 & ~n13357;
  assign n13359 = pi120 & n7443;
  assign n13360 = ~pi120 & n13267;
  assign n13361 = ~n13359 & ~n13360;
  assign n13362 = n7536 & ~n13361;
  assign n13363 = n13276 & ~n13362;
  assign n13364 = ~n13358 & ~n13363;
  assign n13365 = ~pi87 & ~n13364;
  assign n13366 = ~n13321 & ~n13365;
  assign n13367 = ~pi75 & ~n13366;
  assign n13368 = n7360 & ~n13347;
  assign n13369 = ~n13367 & n13368;
  assign n13370 = n7356 & ~n13265;
  assign n13371 = ~n13369 & n13370;
  assign n13372 = ~n13346 & ~n13371;
  assign n13373 = n13261 & ~n13372;
  assign n13374 = ~po1038 & ~n13373;
  assign n13375 = ~n7356 & ~n13292;
  assign n13376 = pi120 & ~n13375;
  assign n13377 = n13261 & ~n13275;
  assign n13378 = ~n13375 & n13377;
  assign n13379 = po1038 & ~n13378;
  assign n13380 = ~n13376 & n13379;
  assign n13381 = ~n7578 & ~n13380;
  assign n13382 = pi951 & pi982;
  assign n13383 = pi1092 & n13382;
  assign n13384 = pi1093 & n13383;
  assign n13385 = ~pi120 & ~n13384;
  assign n13386 = ~n13375 & ~n13385;
  assign n13387 = n13379 & ~n13386;
  assign n13388 = n7578 & ~n13387;
  assign n13389 = ~n13381 & ~n13388;
  assign n13390 = ~n13374 & ~n13389;
  assign n13391 = n13264 & ~n13384;
  assign n13392 = ~n2615 & ~n13385;
  assign n13393 = pi120 & n7533;
  assign n13394 = ~pi1091 & n13384;
  assign n13395 = ~pi120 & ~n13394;
  assign n13396 = n6178 & n13383;
  assign n13397 = ~pi93 & pi950;
  assign n13398 = n7382 & n13397;
  assign n13399 = n8609 & n13398;
  assign n13400 = n2510 & n13399;
  assign n13401 = n9957 & n13400;
  assign n13402 = n7410 & n13401;
  assign n13403 = n2708 & n13402;
  assign n13404 = n13396 & ~n13403;
  assign n13405 = n13395 & ~n13404;
  assign n13406 = ~n13393 & ~n13405;
  assign n13407 = ~n7407 & ~n13406;
  assign n13408 = n7407 & n13385;
  assign n13409 = n2615 & ~n13408;
  assign n13410 = ~n13407 & n13409;
  assign n13411 = pi75 & ~n13392;
  assign n13412 = ~n13410 & n13411;
  assign n13413 = ~n2628 & n13385;
  assign n13414 = pi87 & ~n13413;
  assign n13415 = pi950 & n2523;
  assign n13416 = ~n2921 & ~n6103;
  assign n13417 = n13415 & n13416;
  assign n13418 = n13396 & ~n13417;
  assign n13419 = n2523 & n11855;
  assign n13420 = n13394 & ~n13419;
  assign n13421 = ~n13418 & ~n13420;
  assign n13422 = ~pi120 & ~n13421;
  assign n13423 = ~n7562 & ~n7563;
  assign n13424 = pi120 & ~n13423;
  assign n13425 = n2628 & ~n13424;
  assign n13426 = ~n13422 & n13425;
  assign n13427 = n13414 & ~n13426;
  assign n13428 = n7382 & n7410;
  assign n13429 = n13415 & n13428;
  assign n13430 = n13396 & ~n13429;
  assign n13431 = n13395 & ~n13430;
  assign n13432 = ~n13359 & ~n13431;
  assign n13433 = ~pi39 & n7440;
  assign n13434 = ~n13432 & n13433;
  assign n13435 = pi100 & ~n13434;
  assign n13436 = ~pi38 & ~n13435;
  assign n13437 = ~n7536 & n13385;
  assign n13438 = ~n13436 & ~n13437;
  assign n13439 = n7368 & n9784;
  assign n13440 = n2768 & n13439;
  assign n13441 = n8801 & n13440;
  assign n13442 = n7362 & n13441;
  assign n13443 = n7367 & ~n13442;
  assign n13444 = pi950 & n7380;
  assign n13445 = ~n13443 & n13444;
  assign n13446 = pi824 & n13445;
  assign n13447 = n13383 & ~n13446;
  assign n13448 = ~pi829 & n13447;
  assign n13449 = ~pi97 & ~n13440;
  assign n13450 = n2928 & ~n13449;
  assign n13451 = n2930 & n13450;
  assign n13452 = ~n7457 & ~n13451;
  assign n13453 = n2463 & ~n13452;
  assign n13454 = n7365 & ~n13453;
  assign n13455 = n7362 & ~n13454;
  assign n13456 = ~pi51 & ~n13455;
  assign n13457 = ~n2747 & ~n13456;
  assign n13458 = ~pi96 & ~n13457;
  assign n13459 = n7469 & ~n13458;
  assign n13460 = n7382 & n13383;
  assign n13461 = ~n13459 & n13460;
  assign n13462 = pi122 & n7470;
  assign n13463 = n13382 & n13462;
  assign n13464 = ~n13445 & n13463;
  assign n13465 = ~n13448 & ~n13464;
  assign n13466 = ~n13461 & n13465;
  assign n13467 = n7453 & ~n13466;
  assign n13468 = n7425 & n13383;
  assign n13469 = ~n13467 & ~n13468;
  assign n13470 = pi1091 & ~n13469;
  assign n13471 = n7561 & n13447;
  assign n13472 = ~pi120 & ~n13471;
  assign n13473 = ~n13470 & n13472;
  assign n13474 = ~n7397 & n13348;
  assign n13475 = pi120 & n13474;
  assign n13476 = ~pi39 & ~n13473;
  assign n13477 = ~n13475 & n13476;
  assign n13478 = pi39 & ~n8508;
  assign n13479 = ~n8509 & ~n13385;
  assign n13480 = n13478 & n13479;
  assign n13481 = ~n13477 & ~n13480;
  assign n13482 = n2613 & ~n13481;
  assign n13483 = ~n13438 & ~n13482;
  assign n13484 = ~pi87 & ~n13483;
  assign n13485 = ~pi75 & ~n13427;
  assign n13486 = ~n13484 & n13485;
  assign n13487 = ~n13412 & ~n13486;
  assign n13488 = n7360 & ~n13487;
  assign n13489 = n7356 & ~n13488;
  assign n13490 = n13292 & ~n13385;
  assign n13491 = ~n2531 & ~n13490;
  assign n13492 = ~n7440 & n13490;
  assign n13493 = ~n7418 & n13394;
  assign n13494 = ~n13430 & ~n13493;
  assign n13495 = ~pi120 & ~n13494;
  assign n13496 = ~n13269 & ~n13495;
  assign n13497 = n7440 & ~n13496;
  assign n13498 = n2531 & ~n13492;
  assign n13499 = ~n13497 & n13498;
  assign n13500 = pi100 & ~n13491;
  assign n13501 = ~n13499 & n13500;
  assign n13502 = pi38 & ~n13490;
  assign n13503 = ~n5727 & ~n13490;
  assign n13504 = ~n6205 & ~n13490;
  assign n13505 = ~n7542 & n13268;
  assign n13506 = ~n2921 & n7490;
  assign n13507 = n13396 & ~n13506;
  assign n13508 = ~n13493 & ~n13507;
  assign n13509 = ~pi120 & ~n13508;
  assign n13510 = ~n13505 & ~n13509;
  assign n13511 = n6205 & n13510;
  assign n13512 = ~n13504 & ~n13511;
  assign n13513 = n6221 & n13512;
  assign n13514 = ~n6197 & ~n13510;
  assign n13515 = n6197 & n13490;
  assign n13516 = ~n13514 & ~n13515;
  assign n13517 = ~n6221 & ~n13516;
  assign n13518 = n5727 & ~n13513;
  assign n13519 = ~n13517 & n13518;
  assign n13520 = pi299 & ~n13503;
  assign n13521 = ~n13519 & n13520;
  assign n13522 = ~n7506 & ~n13490;
  assign n13523 = n6194 & n13512;
  assign n13524 = ~n6194 & ~n13516;
  assign n13525 = n7506 & ~n13523;
  assign n13526 = ~n13524 & n13525;
  assign n13527 = ~pi299 & ~n13522;
  assign n13528 = ~n13526 & n13527;
  assign n13529 = ~n13521 & ~n13528;
  assign n13530 = pi39 & ~n13529;
  assign n13531 = ~n7397 & n13290;
  assign n13532 = pi120 & n13531;
  assign n13533 = n13323 & n13447;
  assign n13534 = ~pi120 & ~n13533;
  assign n13535 = ~n13470 & n13534;
  assign n13536 = ~pi39 & ~n13532;
  assign n13537 = ~n13535 & n13536;
  assign n13538 = ~pi38 & ~n13530;
  assign n13539 = ~n13537 & n13538;
  assign n13540 = ~pi100 & ~n13502;
  assign n13541 = ~n13539 & n13540;
  assign n13542 = ~n13501 & ~n13541;
  assign n13543 = ~pi87 & ~n13542;
  assign n13544 = ~n13325 & ~n13425;
  assign n13545 = ~n13418 & ~n13493;
  assign n13546 = n13422 & ~n13545;
  assign n13547 = ~n13544 & ~n13546;
  assign n13548 = ~n13322 & n13414;
  assign n13549 = ~n13547 & n13548;
  assign n13550 = ~n13543 & ~n13549;
  assign n13551 = ~pi75 & ~n13550;
  assign n13552 = n7407 & ~n13490;
  assign n13553 = ~n13404 & ~n13493;
  assign n13554 = ~pi120 & ~n13553;
  assign n13555 = n13336 & ~n13554;
  assign n13556 = ~n13552 & ~n13555;
  assign n13557 = n2615 & ~n13556;
  assign n13558 = ~n2615 & ~n13490;
  assign n13559 = pi75 & ~n13558;
  assign n13560 = ~n13557 & n13559;
  assign n13561 = n7360 & ~n13560;
  assign n13562 = ~n13551 & n13561;
  assign n13563 = n13266 & ~n13562;
  assign n13564 = ~n13489 & ~n13563;
  assign n13565 = n13388 & ~n13391;
  assign n13566 = ~n13564 & n13565;
  assign n13567 = ~n7360 & ~n13375;
  assign n13568 = ~n7351 & n7538;
  assign n13569 = ~n7351 & ~n8509;
  assign n13570 = n13478 & n13569;
  assign n13571 = ~pi39 & ~n13531;
  assign n13572 = ~pi38 & ~n13570;
  assign n13573 = ~n13571 & n13572;
  assign n13574 = ~pi100 & ~n7451;
  assign n13575 = ~n13573 & n13574;
  assign n13576 = ~n13568 & ~n13575;
  assign n13577 = ~pi87 & ~n13576;
  assign n13578 = ~n13327 & ~n13577;
  assign n13579 = ~pi75 & ~n13578;
  assign n13580 = n7351 & ~n7408;
  assign n13581 = n7408 & n13334;
  assign n13582 = pi75 & ~n13580;
  assign n13583 = ~n13581 & n13582;
  assign n13584 = ~n13579 & ~n13583;
  assign n13585 = n13263 & ~n13584;
  assign n13586 = ~pi39 & ~n13474;
  assign n13587 = n7552 & ~n13586;
  assign n13588 = ~pi100 & ~n13587;
  assign n13589 = ~n7538 & ~n13588;
  assign n13590 = ~pi87 & ~n13589;
  assign n13591 = ~n7566 & ~n13590;
  assign n13592 = ~pi75 & ~n13591;
  assign n13593 = ~n7535 & ~n13592;
  assign n13594 = n7356 & ~n13264;
  assign n13595 = ~n13593 & n13594;
  assign n13596 = ~n13567 & ~n13585;
  assign n13597 = ~n13595 & n13596;
  assign n13598 = pi120 & n13381;
  assign n13599 = ~n13597 & n13598;
  assign n13600 = ~n13566 & ~n13599;
  assign n13601 = ~n13261 & ~n13600;
  assign po278 = n13390 | n13601;
  assign n13603 = ~pi134 & ~pi135;
  assign n13604 = ~pi136 & n13603;
  assign n13605 = ~pi130 & n13604;
  assign n13606 = ~pi132 & n13605;
  assign n13607 = ~pi126 & n13606;
  assign n13608 = ~pi121 & n13607;
  assign n13609 = ~pi125 & ~pi133;
  assign n13610 = pi121 & ~n13609;
  assign n13611 = ~pi121 & n13609;
  assign n13612 = ~n13610 & ~n13611;
  assign n13613 = ~n13608 & ~n13612;
  assign n13614 = n2477 & n9790;
  assign n13615 = ~pi51 & n13614;
  assign n13616 = ~pi87 & n13615;
  assign n13617 = ~n13613 & n13616;
  assign n13618 = pi87 & ~n12920;
  assign n13619 = n6166 & ~n13615;
  assign n13620 = pi51 & n6166;
  assign n13621 = ~pi146 & n13620;
  assign n13622 = pi161 & ~n13621;
  assign n13623 = pi51 & pi146;
  assign n13624 = n13619 & ~n13623;
  assign n13625 = ~n13622 & n13624;
  assign n13626 = ~pi87 & ~n13625;
  assign n13627 = pi232 & ~n13618;
  assign n13628 = ~n13626 & n13627;
  assign n13629 = po1038 & ~n13617;
  assign n13630 = ~n13628 & n13629;
  assign n13631 = ~pi184 & ~pi299;
  assign n13632 = ~pi163 & pi299;
  assign n13633 = ~n13631 & ~n13632;
  assign n13634 = n7406 & n13633;
  assign n13635 = pi87 & ~n13634;
  assign n13636 = ~pi87 & ~n7293;
  assign n13637 = ~n13615 & n13636;
  assign n13638 = ~pi142 & n13620;
  assign n13639 = pi144 & ~n13638;
  assign n13640 = pi51 & pi142;
  assign n13641 = n13619 & ~n13640;
  assign n13642 = ~n13639 & n13641;
  assign n13643 = ~pi299 & ~n13642;
  assign n13644 = pi299 & ~n13625;
  assign n13645 = pi232 & ~n13643;
  assign n13646 = ~n13644 & n13645;
  assign n13647 = n13637 & ~n13646;
  assign n13648 = pi38 & ~n13646;
  assign n13649 = ~pi100 & ~n13648;
  assign n13650 = pi38 & ~n13615;
  assign n13651 = ~pi100 & ~n13650;
  assign n13652 = ~n13649 & ~n13651;
  assign n13653 = ~pi161 & ~n13621;
  assign n13654 = ~pi96 & n7377;
  assign n13655 = ~pi24 & pi314;
  assign n13656 = n13654 & n13655;
  assign n13657 = n2767 & n9878;
  assign n13658 = n9789 & n13657;
  assign n13659 = n12328 & n13658;
  assign n13660 = pi77 & ~pi86;
  assign n13661 = n13659 & n13660;
  assign n13662 = n8611 & n13656;
  assign n13663 = n13661 & n13662;
  assign n13664 = n3174 & n13663;
  assign n13665 = ~pi51 & ~n13614;
  assign n13666 = ~n2711 & ~n13665;
  assign n13667 = ~pi77 & n13659;
  assign n13668 = ~pi24 & n11257;
  assign n13669 = n13667 & n13668;
  assign n13670 = pi86 & n13667;
  assign n13671 = ~n13661 & ~n13670;
  assign n13672 = n10680 & ~n13671;
  assign n13673 = n13614 & ~n13669;
  assign n13674 = ~n13672 & n13673;
  assign n13675 = ~n13666 & ~n13674;
  assign n13676 = n3174 & n13675;
  assign n13677 = n13615 & ~n13676;
  assign n13678 = ~pi58 & n13654;
  assign n13679 = n8943 & n13678;
  assign n13680 = n13667 & n13679;
  assign n13681 = pi72 & n6431;
  assign n13682 = n13680 & n13681;
  assign n13683 = n13677 & ~n13682;
  assign n13684 = ~n13664 & n13683;
  assign n13685 = ~n6166 & ~n13684;
  assign n13686 = pi72 & n9975;
  assign n13687 = ~n13620 & ~n13686;
  assign n13688 = n6166 & ~n13687;
  assign n13689 = ~n13685 & ~n13688;
  assign n13690 = n13653 & ~n13689;
  assign n13691 = n13615 & ~n13664;
  assign n13692 = ~n13676 & n13691;
  assign n13693 = ~n6166 & ~n13692;
  assign n13694 = ~n13619 & ~n13693;
  assign n13695 = ~n13682 & n13694;
  assign n13696 = n13622 & ~n13695;
  assign n13697 = ~n13690 & ~n13696;
  assign n13698 = n9121 & ~n13697;
  assign n13699 = ~n13664 & n13695;
  assign n13700 = n13622 & ~n13699;
  assign n13701 = ~pi51 & n13656;
  assign n13702 = n12698 & n13701;
  assign n13703 = n2701 & n8787;
  assign n13704 = n13702 & n13703;
  assign n13705 = n13689 & ~n13704;
  assign n13706 = pi146 & n13705;
  assign n13707 = ~n6166 & n13684;
  assign n13708 = ~pi72 & ~n13702;
  assign n13709 = n6432 & ~n13708;
  assign n13710 = n6166 & ~n13709;
  assign n13711 = ~n13707 & ~n13710;
  assign n13712 = ~pi146 & ~n13711;
  assign n13713 = ~pi161 & ~n13712;
  assign n13714 = ~n13706 & n13713;
  assign n13715 = ~n13700 & ~n13714;
  assign n13716 = n9030 & ~n13715;
  assign n13717 = ~n13698 & ~n13716;
  assign n13718 = pi156 & ~n13717;
  assign n13719 = n9030 & ~n13621;
  assign n13720 = ~n13684 & n13719;
  assign n13721 = ~pi51 & n6166;
  assign n13722 = ~n13683 & n13721;
  assign n13723 = ~n13685 & ~n13722;
  assign n13724 = n6166 & n13665;
  assign n13725 = ~n13703 & ~n13724;
  assign n13726 = n3174 & ~n13675;
  assign n13727 = ~n13725 & ~n13726;
  assign n13728 = pi146 & ~n13727;
  assign n13729 = n6166 & ~n13677;
  assign n13730 = ~pi146 & ~n13729;
  assign n13731 = ~n13728 & ~n13730;
  assign n13732 = ~n13694 & ~n13731;
  assign n13733 = n13723 & ~n13732;
  assign n13734 = n9121 & ~n13733;
  assign n13735 = pi161 & ~n13720;
  assign n13736 = ~n13734 & n13735;
  assign n13737 = ~n10680 & ~n11257;
  assign n13738 = n11254 & ~n13737;
  assign n13739 = n2711 & n13738;
  assign n13740 = ~pi72 & ~n13739;
  assign n13741 = n6432 & ~n13740;
  assign n13742 = n6166 & ~n13741;
  assign n13743 = ~n13707 & ~n13742;
  assign n13744 = ~pi146 & ~n13743;
  assign n13745 = n13703 & n13739;
  assign n13746 = ~n13688 & ~n13745;
  assign n13747 = ~n13685 & n13746;
  assign n13748 = pi146 & n13747;
  assign n13749 = n9121 & ~n13748;
  assign n13750 = ~n13744 & n13749;
  assign n13751 = ~pi314 & ~n13738;
  assign n13752 = pi314 & ~n11255;
  assign n13753 = ~n13751 & ~n13752;
  assign n13754 = n2711 & n13753;
  assign n13755 = ~pi72 & ~n13754;
  assign n13756 = n6432 & ~n13755;
  assign n13757 = n6166 & ~n13756;
  assign n13758 = ~n13707 & ~n13757;
  assign n13759 = ~pi146 & ~n13758;
  assign n13760 = n7376 & n10657;
  assign n13761 = n13753 & n13760;
  assign n13762 = ~pi51 & ~n13761;
  assign n13763 = ~n13686 & n13762;
  assign n13764 = n6166 & ~n13763;
  assign n13765 = ~n13685 & ~n13764;
  assign n13766 = pi146 & n13765;
  assign n13767 = n9030 & ~n13759;
  assign n13768 = ~n13766 & n13767;
  assign n13769 = ~pi161 & ~n13750;
  assign n13770 = ~n13768 & n13769;
  assign n13771 = ~pi156 & ~n13736;
  assign n13772 = ~n13770 & n13771;
  assign n13773 = n13639 & ~n13684;
  assign n13774 = ~pi142 & ~n13758;
  assign n13775 = pi142 & n13765;
  assign n13776 = ~pi144 & ~n13774;
  assign n13777 = ~n13775 & n13776;
  assign n13778 = ~n13773 & ~n13777;
  assign n13779 = ~pi180 & ~n13778;
  assign n13780 = pi142 & ~n13727;
  assign n13781 = ~pi142 & ~n13729;
  assign n13782 = ~n13780 & ~n13781;
  assign n13783 = ~n13694 & ~n13782;
  assign n13784 = pi144 & n13723;
  assign n13785 = ~n13783 & n13784;
  assign n13786 = ~pi142 & n13743;
  assign n13787 = pi142 & ~n13747;
  assign n13788 = ~pi144 & ~n13787;
  assign n13789 = ~n13786 & n13788;
  assign n13790 = pi180 & ~n13785;
  assign n13791 = ~n13789 & n13790;
  assign n13792 = ~n13779 & ~n13791;
  assign n13793 = ~pi179 & ~n13792;
  assign n13794 = ~pi144 & n13689;
  assign n13795 = pi144 & n13695;
  assign n13796 = ~n13638 & ~n13795;
  assign n13797 = ~n13794 & n13796;
  assign n13798 = pi180 & ~n13797;
  assign n13799 = n13639 & ~n13699;
  assign n13800 = pi142 & n13705;
  assign n13801 = ~pi142 & ~n13711;
  assign n13802 = ~pi144 & ~n13801;
  assign n13803 = ~n13800 & n13802;
  assign n13804 = ~pi180 & ~n13799;
  assign n13805 = ~n13803 & n13804;
  assign n13806 = pi179 & ~n13798;
  assign n13807 = ~n13805 & n13806;
  assign n13808 = ~n13793 & ~n13807;
  assign n13809 = ~pi299 & ~n13808;
  assign n13810 = ~n13718 & ~n13772;
  assign n13811 = ~n13809 & n13810;
  assign n13812 = n8769 & ~n13811;
  assign n13813 = n3174 & n13680;
  assign n13814 = ~n6590 & ~n7547;
  assign n13815 = n13813 & ~n13814;
  assign n13816 = ~pi232 & n13615;
  assign n13817 = ~n13815 & n13816;
  assign n13818 = n13615 & ~n13813;
  assign n13819 = ~pi51 & ~n13818;
  assign n13820 = ~pi287 & ~n13819;
  assign n13821 = ~pi287 & n6166;
  assign n13822 = ~n13724 & ~n13821;
  assign n13823 = ~n13820 & ~n13822;
  assign n13824 = ~n13641 & ~n13823;
  assign n13825 = n8752 & ~n13824;
  assign n13826 = n13614 & n13825;
  assign n13827 = ~n13615 & ~n13638;
  assign n13828 = ~n6359 & ~n13827;
  assign n13829 = pi144 & ~n13828;
  assign n13830 = pi51 & ~n6166;
  assign n13831 = ~n13819 & ~n13830;
  assign n13832 = n6359 & ~n13640;
  assign n13833 = n13831 & n13832;
  assign n13834 = n13829 & ~n13833;
  assign n13835 = ~n13826 & n13834;
  assign n13836 = ~n6166 & ~n13818;
  assign n13837 = ~n6185 & ~n13836;
  assign n13838 = ~pi142 & ~n13837;
  assign n13839 = n2517 & n10657;
  assign n13840 = ~pi51 & ~n13839;
  assign n13841 = n6166 & ~n13840;
  assign n13842 = ~n13836 & ~n13841;
  assign n13843 = pi142 & ~n13842;
  assign n13844 = n6359 & ~n13843;
  assign n13845 = ~n13838 & n13844;
  assign n13846 = ~n8752 & ~n13845;
  assign n13847 = ~pi51 & n13821;
  assign n13848 = ~n13842 & ~n13847;
  assign n13849 = pi224 & ~n13638;
  assign n13850 = n13848 & n13849;
  assign n13851 = ~n13846 & ~n13850;
  assign n13852 = ~n6359 & n13724;
  assign n13853 = ~n13828 & ~n13852;
  assign n13854 = ~n13829 & n13853;
  assign n13855 = ~n13851 & n13854;
  assign n13856 = pi181 & ~n13835;
  assign n13857 = ~n13855 & n13856;
  assign n13858 = ~n13845 & n13854;
  assign n13859 = ~pi181 & ~n13834;
  assign n13860 = ~n13858 & n13859;
  assign n13861 = ~pi299 & ~n13860;
  assign n13862 = ~n13857 & n13861;
  assign n13863 = ~n13615 & ~n13625;
  assign n13864 = ~n5726 & ~n13863;
  assign n13865 = ~n13621 & ~n13818;
  assign n13866 = pi161 & ~n13865;
  assign n13867 = ~pi146 & ~n13837;
  assign n13868 = pi146 & ~n13842;
  assign n13869 = ~pi161 & ~n13868;
  assign n13870 = ~n13867 & n13869;
  assign n13871 = ~n13866 & ~n13870;
  assign n13872 = n5726 & ~n13871;
  assign n13873 = ~n8739 & ~n13872;
  assign n13874 = n13653 & n13848;
  assign n13875 = n13813 & ~n13821;
  assign n13876 = n13615 & ~n13875;
  assign n13877 = n13622 & ~n13876;
  assign n13878 = ~n13874 & ~n13877;
  assign n13879 = pi216 & ~n13878;
  assign n13880 = ~n13873 & ~n13879;
  assign n13881 = n9599 & ~n13864;
  assign n13882 = ~n13880 & n13881;
  assign n13883 = n9573 & ~n13864;
  assign n13884 = ~n13872 & n13883;
  assign n13885 = pi232 & ~n13884;
  assign n13886 = ~n13862 & n13885;
  assign n13887 = ~n13882 & n13886;
  assign n13888 = pi39 & ~n13817;
  assign n13889 = ~n13887 & n13888;
  assign n13890 = ~pi39 & ~pi232;
  assign n13891 = ~n13684 & n13890;
  assign n13892 = ~n13889 & ~n13891;
  assign n13893 = ~n13812 & n13892;
  assign n13894 = ~pi38 & ~n13893;
  assign n13895 = ~n13652 & ~n13894;
  assign n13896 = pi100 & n13646;
  assign n13897 = pi100 & n13615;
  assign n13898 = n2536 & ~n13897;
  assign n13899 = ~n13896 & n13898;
  assign n13900 = ~n13895 & n13899;
  assign n13901 = ~n13613 & ~n13635;
  assign n13902 = ~n13647 & n13901;
  assign n13903 = ~n13900 & n13902;
  assign n13904 = n13636 & ~n13646;
  assign n13905 = ~pi159 & n13644;
  assign n13906 = ~n8739 & n13625;
  assign n13907 = n13653 & ~n13823;
  assign n13908 = n6166 & n6333;
  assign n13909 = n13622 & ~n13908;
  assign n13910 = n8739 & ~n13907;
  assign n13911 = ~n13909 & n13910;
  assign n13912 = n9599 & ~n13906;
  assign n13913 = ~n13911 & n13912;
  assign n13914 = ~pi181 & n13642;
  assign n13915 = ~pi144 & ~n13641;
  assign n13916 = ~n13825 & n13915;
  assign n13917 = n8752 & n13821;
  assign n13918 = ~n13640 & n13917;
  assign n13919 = n13839 & n13918;
  assign n13920 = n13639 & ~n13919;
  assign n13921 = pi181 & ~n13916;
  assign n13922 = ~n13920 & n13921;
  assign n13923 = ~pi299 & ~n13914;
  assign n13924 = ~n13922 & n13923;
  assign n13925 = n8738 & ~n13905;
  assign n13926 = ~n13913 & n13925;
  assign n13927 = ~n13924 & n13926;
  assign n13928 = n6166 & ~n13692;
  assign n13929 = ~pi142 & n13928;
  assign n13930 = n13614 & ~n13663;
  assign n13931 = n13654 & n13930;
  assign n13932 = n13674 & n13931;
  assign n13933 = ~n13666 & ~n13932;
  assign n13934 = n3174 & ~n13933;
  assign n13935 = ~n13725 & ~n13934;
  assign n13936 = pi142 & n13935;
  assign n13937 = ~pi144 & ~n13929;
  assign n13938 = ~n13936 & n13937;
  assign n13939 = n6166 & ~n13762;
  assign n13940 = ~n13640 & n13939;
  assign n13941 = pi144 & ~n13940;
  assign n13942 = pi180 & ~n13938;
  assign n13943 = ~n13941 & n13942;
  assign n13944 = n13639 & ~n13745;
  assign n13945 = ~pi144 & ~n13782;
  assign n13946 = ~pi180 & ~n13945;
  assign n13947 = ~n13944 & n13946;
  assign n13948 = pi179 & ~n13947;
  assign n13949 = ~n13943 & n13948;
  assign n13950 = ~pi180 & n13642;
  assign n13951 = n6166 & ~n13691;
  assign n13952 = ~pi142 & n13951;
  assign n13953 = ~pi51 & ~n13930;
  assign n13954 = n3174 & ~n13953;
  assign n13955 = ~n13725 & ~n13954;
  assign n13956 = pi142 & n13955;
  assign n13957 = ~pi144 & ~n13952;
  assign n13958 = ~n13956 & n13957;
  assign n13959 = n13639 & ~n13704;
  assign n13960 = pi180 & ~n13958;
  assign n13961 = ~n13959 & n13960;
  assign n13962 = ~pi179 & ~n13950;
  assign n13963 = ~n13961 & n13962;
  assign n13964 = ~n13949 & ~n13963;
  assign n13965 = ~pi299 & ~n13964;
  assign n13966 = ~n13623 & n13939;
  assign n13967 = pi161 & ~n13966;
  assign n13968 = pi146 & n13935;
  assign n13969 = ~pi146 & n13928;
  assign n13970 = ~pi161 & ~n13968;
  assign n13971 = ~n13969 & n13970;
  assign n13972 = ~n13967 & ~n13971;
  assign n13973 = n9121 & ~n13972;
  assign n13974 = n13622 & ~n13745;
  assign n13975 = ~pi161 & ~n13731;
  assign n13976 = ~n13974 & ~n13975;
  assign n13977 = n9030 & ~n13976;
  assign n13978 = pi232 & ~n13977;
  assign n13979 = ~n13973 & n13978;
  assign n13980 = pi156 & ~n13979;
  assign n13981 = ~pi39 & ~n13965;
  assign n13982 = ~n13980 & n13981;
  assign n13983 = ~pi38 & ~n13927;
  assign n13984 = ~n13982 & n13983;
  assign n13985 = ~pi158 & n13644;
  assign n13986 = n13622 & ~n13704;
  assign n13987 = ~pi146 & n13951;
  assign n13988 = pi146 & n13955;
  assign n13989 = ~pi161 & ~n13987;
  assign n13990 = ~n13988 & n13989;
  assign n13991 = ~n13986 & ~n13990;
  assign n13992 = n9121 & ~n13991;
  assign n13993 = pi232 & ~n13985;
  assign n13994 = ~n13992 & n13993;
  assign n13995 = ~pi156 & n2531;
  assign n13996 = ~n13994 & n13995;
  assign n13997 = n13649 & ~n13996;
  assign n13998 = ~n13984 & n13997;
  assign n13999 = n2536 & ~n13896;
  assign n14000 = ~n13998 & n13999;
  assign n14001 = n13613 & ~n13635;
  assign n14002 = ~n13904 & n14001;
  assign n14003 = ~n14000 & n14002;
  assign n14004 = ~po1038 & ~n14003;
  assign n14005 = ~n13903 & n14004;
  assign po279 = n13630 | n14005;
  assign n14007 = n7351 & n7358;
  assign n14008 = n7360 & n13584;
  assign n14009 = n13263 & ~n14008;
  assign n14010 = n7360 & n13593;
  assign n14011 = n7356 & ~n14010;
  assign n14012 = ~po1038 & ~n14009;
  assign n14013 = ~n14011 & n14012;
  assign po280 = n14007 | n14013;
  assign n14015 = ~pi39 & pi110;
  assign n14016 = n9710 & n14015;
  assign n14017 = ~n10578 & n14016;
  assign n14018 = po1057 & n14017;
  assign n14019 = ~pi110 & n8981;
  assign n14020 = ~n6223 & n14019;
  assign n14021 = pi39 & n5726;
  assign n14022 = n14020 & n14021;
  assign n14023 = ~n14018 & ~n14022;
  assign n14024 = po1038 & ~n14023;
  assign n14025 = pi110 & n12705;
  assign n14026 = ~pi39 & ~n14025;
  assign n14027 = ~n6207 & n7547;
  assign n14028 = n14019 & n14027;
  assign n14029 = n6590 & n14020;
  assign n14030 = pi39 & ~n14028;
  assign n14031 = ~n14029 & n14030;
  assign n14032 = ~n14026 & ~n14031;
  assign n14033 = ~n2576 & ~n14032;
  assign n14034 = pi72 & n2711;
  assign n14035 = n10009 & n14034;
  assign n14036 = ~pi111 & ~n6379;
  assign n14037 = ~pi36 & n2808;
  assign n14038 = ~n14036 & n14037;
  assign n14039 = n2792 & ~n14038;
  assign n14040 = ~n2791 & ~n2797;
  assign n14041 = ~n14039 & n14040;
  assign n14042 = ~pi83 & ~n14041;
  assign n14043 = n2795 & ~n14042;
  assign n14044 = ~pi71 & ~n14043;
  assign n14045 = n6389 & ~n14044;
  assign n14046 = ~pi81 & ~n14045;
  assign n14047 = n11034 & ~n14046;
  assign n14048 = ~pi90 & ~n14047;
  assign n14049 = n2710 & ~n14048;
  assign n14050 = pi90 & ~n10009;
  assign n14051 = ~pi72 & ~pi93;
  assign n14052 = ~n14050 & n14051;
  assign n14053 = n14049 & n14052;
  assign n14054 = ~n14035 & ~n14053;
  assign n14055 = n6431 & ~n14054;
  assign n14056 = ~pi110 & ~n14055;
  assign n14057 = n12705 & ~n14056;
  assign n14058 = n2898 & n14049;
  assign n14059 = ~pi72 & ~n14058;
  assign n14060 = n6432 & ~n12705;
  assign n14061 = ~n14059 & n14060;
  assign n14062 = ~pi39 & ~n14061;
  assign n14063 = ~n14057 & n14062;
  assign n14064 = ~n14031 & ~n14063;
  assign n14065 = n2576 & ~n14064;
  assign n14066 = ~po1038 & ~n14033;
  assign n14067 = ~n14065 & n14066;
  assign po281 = ~n14024 & ~n14067;
  assign n14069 = ~pi125 & n13608;
  assign n14070 = pi125 & pi133;
  assign n14071 = ~n13609 & ~n14070;
  assign n14072 = ~n14069 & ~n14071;
  assign n14073 = n13615 & ~n14072;
  assign n14074 = pi172 & n13620;
  assign n14075 = ~pi152 & n13724;
  assign n14076 = ~n14074 & ~n14075;
  assign n14077 = pi232 & ~n14076;
  assign n14078 = ~n14073 & ~n14077;
  assign n14079 = ~pi87 & ~n14078;
  assign n14080 = pi87 & n9536;
  assign n14081 = po1038 & ~n14080;
  assign n14082 = ~n14079 & n14081;
  assign n14083 = pi193 & n13620;
  assign n14084 = ~pi174 & n13724;
  assign n14085 = ~pi299 & ~n14083;
  assign n14086 = ~n14084 & n14085;
  assign n14087 = pi299 & n14076;
  assign n14088 = pi232 & ~n14086;
  assign n14089 = ~n14087 & n14088;
  assign n14090 = pi100 & n14089;
  assign n14091 = pi38 & ~n14089;
  assign n14092 = ~pi100 & ~n14091;
  assign n14093 = ~n13651 & ~n14092;
  assign n14094 = ~pi193 & n13620;
  assign n14095 = ~pi145 & n13955;
  assign n14096 = ~n13724 & ~n14095;
  assign n14097 = pi174 & ~n14096;
  assign n14098 = ~pi145 & n13704;
  assign n14099 = ~pi174 & n14098;
  assign n14100 = ~n13693 & ~n14094;
  assign n14101 = ~n14097 & n14100;
  assign n14102 = ~n14099 & n14101;
  assign n14103 = n9430 & ~n14102;
  assign n14104 = ~n13693 & ~n13745;
  assign n14105 = pi145 & n14104;
  assign n14106 = n13703 & n13754;
  assign n14107 = ~n13693 & ~n14106;
  assign n14108 = ~pi145 & n14107;
  assign n14109 = ~pi174 & ~n14105;
  assign n14110 = ~n14108 & n14109;
  assign n14111 = ~n13693 & ~n13935;
  assign n14112 = ~n6166 & ~n13691;
  assign n14113 = ~n13619 & ~n14112;
  assign n14114 = ~n13676 & n14113;
  assign n14115 = ~n14095 & n14114;
  assign n14116 = n3174 & n14115;
  assign n14117 = pi174 & ~n14111;
  assign n14118 = ~n14116 & n14117;
  assign n14119 = pi193 & ~n14118;
  assign n14120 = ~n14110 & n14119;
  assign n14121 = pi174 & ~n14115;
  assign n14122 = ~pi51 & n14105;
  assign n14123 = ~pi145 & ~n13693;
  assign n14124 = ~n13939 & n14123;
  assign n14125 = ~pi174 & ~n14122;
  assign n14126 = ~n14124 & n14125;
  assign n14127 = ~pi193 & ~n14121;
  assign n14128 = ~n14126 & n14127;
  assign n14129 = n9426 & ~n14120;
  assign n14130 = ~n14128 & n14129;
  assign n14131 = ~n14103 & ~n14130;
  assign n14132 = ~pi38 & ~n14131;
  assign n14133 = ~pi172 & n13620;
  assign n14134 = ~pi172 & ~n14114;
  assign n14135 = ~n13693 & ~n13727;
  assign n14136 = pi172 & ~n14135;
  assign n14137 = ~n14134 & ~n14136;
  assign n14138 = pi152 & ~n14137;
  assign n14139 = ~pi152 & ~n14104;
  assign n14140 = pi197 & ~n14133;
  assign n14141 = ~n14138 & n14140;
  assign n14142 = ~n14139 & n14141;
  assign n14143 = pi152 & ~n14111;
  assign n14144 = ~pi152 & ~n14107;
  assign n14145 = pi172 & ~n14143;
  assign n14146 = ~n14144 & n14145;
  assign n14147 = ~pi152 & n13939;
  assign n14148 = ~pi152 & n6166;
  assign n14149 = ~n13692 & ~n14148;
  assign n14150 = ~pi172 & ~n14149;
  assign n14151 = ~n14147 & n14150;
  assign n14152 = ~n14146 & ~n14151;
  assign n14153 = ~pi197 & ~n14152;
  assign n14154 = pi299 & n9420;
  assign n14155 = ~n14142 & n14154;
  assign n14156 = ~n14153 & n14155;
  assign n14157 = ~pi172 & ~n14075;
  assign n14158 = ~n13694 & n14157;
  assign n14159 = pi152 & n13724;
  assign n14160 = ~n13693 & ~n14159;
  assign n14161 = pi172 & ~n14160;
  assign n14162 = pi197 & ~n14158;
  assign n14163 = ~n14161 & n14162;
  assign n14164 = ~n13693 & ~n13955;
  assign n14165 = pi172 & ~n14164;
  assign n14166 = ~n13693 & ~n13951;
  assign n14167 = ~pi172 & ~n14166;
  assign n14168 = pi152 & ~n14165;
  assign n14169 = ~n14167 & n14168;
  assign n14170 = ~n13693 & ~n13704;
  assign n14171 = ~pi152 & ~n14133;
  assign n14172 = n14170 & n14171;
  assign n14173 = ~n14169 & ~n14172;
  assign n14174 = ~pi197 & ~n14173;
  assign n14175 = pi299 & n9414;
  assign n14176 = ~n14163 & n14175;
  assign n14177 = ~n14174 & n14176;
  assign n14178 = ~n14156 & ~n14177;
  assign n14179 = ~n14132 & n14178;
  assign n14180 = n8769 & ~n14179;
  assign n14181 = n8752 & n13813;
  assign n14182 = n13615 & ~n14181;
  assign n14183 = ~pi299 & ~n14182;
  assign n14184 = n8739 & n13813;
  assign n14185 = n13615 & ~n14184;
  assign n14186 = pi299 & ~n14185;
  assign n14187 = ~n14183 & ~n14186;
  assign n14188 = ~pi232 & ~n14187;
  assign n14189 = pi39 & ~n14188;
  assign n14190 = ~n13615 & n14076;
  assign n14191 = ~n8739 & ~n14190;
  assign n14192 = ~pi152 & ~n13848;
  assign n14193 = pi152 & n13876;
  assign n14194 = ~n14074 & ~n14193;
  assign n14195 = ~n14192 & n14194;
  assign n14196 = n8739 & ~n14195;
  assign n14197 = n9121 & ~n14196;
  assign n14198 = ~n13818 & ~n14148;
  assign n14199 = ~pi152 & n13841;
  assign n14200 = ~n14198 & ~n14199;
  assign n14201 = ~pi172 & ~n14200;
  assign n14202 = ~pi152 & n13837;
  assign n14203 = pi152 & n13831;
  assign n14204 = pi172 & ~n14203;
  assign n14205 = ~n14202 & n14204;
  assign n14206 = n8739 & ~n14201;
  assign n14207 = ~n14205 & n14206;
  assign n14208 = n9030 & ~n14207;
  assign n14209 = ~n14197 & ~n14208;
  assign n14210 = ~n14191 & ~n14209;
  assign n14211 = pi180 & n13847;
  assign n14212 = ~n6166 & ~n13614;
  assign n14213 = ~n8752 & ~n14212;
  assign n14214 = ~pi51 & n14213;
  assign n14215 = ~n13842 & ~n14214;
  assign n14216 = ~pi174 & ~n14211;
  assign n14217 = n14215 & n14216;
  assign n14218 = pi180 & n13876;
  assign n14219 = pi174 & ~n14182;
  assign n14220 = ~n14218 & n14219;
  assign n14221 = ~pi193 & ~n14220;
  assign n14222 = ~n14217 & n14221;
  assign n14223 = ~n13830 & n14213;
  assign n14224 = n8752 & n13837;
  assign n14225 = ~n14223 & ~n14224;
  assign n14226 = ~pi174 & ~n14225;
  assign n14227 = ~n13620 & ~n14182;
  assign n14228 = pi174 & ~n14227;
  assign n14229 = ~pi180 & ~n14228;
  assign n14230 = ~n14226 & n14229;
  assign n14231 = ~n10167 & ~n13836;
  assign n14232 = n8752 & n14231;
  assign n14233 = ~n14223 & ~n14232;
  assign n14234 = ~pi174 & ~n14233;
  assign n14235 = ~pi51 & ~n13876;
  assign n14236 = n6166 & ~n14235;
  assign n14237 = ~n14182 & ~n14236;
  assign n14238 = pi174 & ~n14237;
  assign n14239 = pi180 & ~n14238;
  assign n14240 = ~n14234 & n14239;
  assign n14241 = pi193 & ~n14240;
  assign n14242 = ~n14230 & n14241;
  assign n14243 = ~pi299 & ~n14222;
  assign n14244 = ~n14242 & n14243;
  assign n14245 = ~n14210 & ~n14244;
  assign n14246 = pi232 & ~n14245;
  assign n14247 = n14189 & ~n14246;
  assign n14248 = ~pi232 & ~n13692;
  assign n14249 = ~pi39 & ~n14248;
  assign n14250 = ~pi38 & ~n14249;
  assign n14251 = ~n14247 & n14250;
  assign n14252 = ~n14093 & ~n14251;
  assign n14253 = ~n14180 & n14252;
  assign n14254 = n13898 & ~n14090;
  assign n14255 = ~n14253 & n14254;
  assign n14256 = pi140 & ~pi299;
  assign n14257 = pi162 & pi299;
  assign n14258 = ~n14256 & ~n14257;
  assign n14259 = n7406 & ~n14258;
  assign n14260 = pi87 & ~n14259;
  assign n14261 = n13637 & ~n14089;
  assign n14262 = ~n14072 & ~n14260;
  assign n14263 = ~n14261 & n14262;
  assign n14264 = ~n14255 & n14263;
  assign n14265 = ~n7544 & ~n7548;
  assign n14266 = n2523 & ~n14265;
  assign n14267 = ~pi232 & ~n14266;
  assign n14268 = pi39 & ~n14267;
  assign n14269 = ~n5727 & n14076;
  assign n14270 = n2523 & ~n6166;
  assign n14271 = n6166 & ~n13818;
  assign n14272 = ~n14270 & ~n14271;
  assign n14273 = ~pi152 & n14272;
  assign n14274 = pi51 & ~pi172;
  assign n14275 = ~n13830 & ~n13840;
  assign n14276 = pi152 & ~n14275;
  assign n14277 = ~n14273 & ~n14274;
  assign n14278 = ~n14276 & n14277;
  assign n14279 = ~pi216 & ~n14278;
  assign n14280 = n5726 & n14279;
  assign n14281 = ~n14269 & ~n14280;
  assign n14282 = n9030 & ~n14281;
  assign n14283 = ~n5726 & ~n14076;
  assign n14284 = n13813 & n13821;
  assign n14285 = ~n13619 & ~n14284;
  assign n14286 = ~pi152 & ~n14285;
  assign n14287 = n13821 & n13839;
  assign n14288 = ~n13620 & ~n14287;
  assign n14289 = pi152 & ~n14288;
  assign n14290 = pi172 & ~n14286;
  assign n14291 = ~n14289 & n14290;
  assign n14292 = ~pi152 & n13823;
  assign n14293 = pi152 & n13908;
  assign n14294 = ~pi172 & ~n14292;
  assign n14295 = ~n14293 & n14294;
  assign n14296 = ~n14291 & ~n14295;
  assign n14297 = pi216 & ~n14296;
  assign n14298 = n5726 & ~n14279;
  assign n14299 = ~n14297 & n14298;
  assign n14300 = n9121 & ~n14283;
  assign n14301 = ~n14299 & n14300;
  assign n14302 = ~n7506 & ~n13619;
  assign n14303 = n6166 & n13819;
  assign n14304 = ~n14270 & ~n14303;
  assign n14305 = ~n14302 & ~n14304;
  assign n14306 = ~pi174 & n14305;
  assign n14307 = n7506 & n13839;
  assign n14308 = ~pi51 & n14307;
  assign n14309 = pi174 & n14308;
  assign n14310 = ~n14083 & ~n14309;
  assign n14311 = ~n14306 & n14310;
  assign n14312 = ~pi180 & ~n14311;
  assign n14313 = n7506 & n14272;
  assign n14314 = pi224 & ~n14284;
  assign n14315 = n6359 & ~n14314;
  assign n14316 = ~n13619 & ~n14315;
  assign n14317 = ~n14313 & ~n14316;
  assign n14318 = ~pi174 & ~n14317;
  assign n14319 = pi224 & n14288;
  assign n14320 = n6359 & ~n14319;
  assign n14321 = n7506 & ~n14275;
  assign n14322 = n14320 & ~n14321;
  assign n14323 = ~n13620 & ~n14322;
  assign n14324 = pi174 & n14323;
  assign n14325 = pi193 & ~n14318;
  assign n14326 = ~n14324 & n14325;
  assign n14327 = ~n7506 & ~n13917;
  assign n14328 = n2523 & ~n14327;
  assign n14329 = pi174 & ~n14328;
  assign n14330 = pi224 & ~n13823;
  assign n14331 = ~pi224 & n14304;
  assign n14332 = n6359 & ~n14330;
  assign n14333 = ~n14331 & n14332;
  assign n14334 = ~n13852 & ~n14333;
  assign n14335 = ~pi174 & n14334;
  assign n14336 = ~pi193 & ~n14329;
  assign n14337 = ~n14335 & n14336;
  assign n14338 = ~n14326 & ~n14337;
  assign n14339 = pi180 & ~n14338;
  assign n14340 = ~pi299 & ~n14312;
  assign n14341 = ~n14339 & n14340;
  assign n14342 = ~n14282 & ~n14301;
  assign n14343 = ~n14341 & n14342;
  assign n14344 = pi232 & ~n14343;
  assign n14345 = n14268 & ~n14344;
  assign n14346 = ~pi232 & ~n13686;
  assign n14347 = ~pi39 & ~n14346;
  assign n14348 = ~pi38 & ~n14347;
  assign n14349 = ~n14345 & n14348;
  assign n14350 = pi145 & n13955;
  assign n14351 = n13614 & ~n13682;
  assign n14352 = n13721 & ~n14351;
  assign n14353 = ~n6166 & n13686;
  assign n14354 = ~n14352 & ~n14353;
  assign n14355 = ~pi174 & ~n14350;
  assign n14356 = n14354 & n14355;
  assign n14357 = ~pi145 & n13686;
  assign n14358 = ~n6166 & ~n13686;
  assign n14359 = ~n13710 & ~n14358;
  assign n14360 = pi145 & n14359;
  assign n14361 = pi174 & ~n14357;
  assign n14362 = ~n14360 & n14361;
  assign n14363 = ~n14356 & ~n14362;
  assign n14364 = ~pi193 & ~n14363;
  assign n14365 = n13721 & n14351;
  assign n14366 = ~n13620 & ~n13664;
  assign n14367 = pi145 & ~n14366;
  assign n14368 = n14365 & ~n14367;
  assign n14369 = ~pi174 & ~n14368;
  assign n14370 = ~n14358 & n14369;
  assign n14371 = n13687 & ~n13704;
  assign n14372 = pi174 & ~n14098;
  assign n14373 = ~n14371 & n14372;
  assign n14374 = pi193 & ~n14370;
  assign n14375 = ~n14373 & n14374;
  assign n14376 = ~n14364 & ~n14375;
  assign n14377 = n9426 & ~n14376;
  assign n14378 = ~n13763 & ~n14358;
  assign n14379 = pi145 & n14378;
  assign n14380 = n13687 & ~n13745;
  assign n14381 = ~pi145 & ~n14380;
  assign n14382 = pi193 & ~n14381;
  assign n14383 = ~n14379 & n14382;
  assign n14384 = ~n13742 & ~n14358;
  assign n14385 = ~pi145 & n14384;
  assign n14386 = ~n13757 & ~n14358;
  assign n14387 = pi145 & n14386;
  assign n14388 = ~pi193 & ~n14385;
  assign n14389 = ~n14387 & n14388;
  assign n14390 = ~n14383 & ~n14389;
  assign n14391 = pi174 & ~n14390;
  assign n14392 = ~n13722 & ~n14083;
  assign n14393 = n14356 & n14392;
  assign n14394 = ~n14391 & ~n14393;
  assign n14395 = n9430 & ~n14394;
  assign n14396 = ~n14377 & ~n14395;
  assign n14397 = ~pi38 & ~n14396;
  assign n14398 = ~pi152 & n14352;
  assign n14399 = n13686 & ~n14148;
  assign n14400 = ~pi197 & ~n14398;
  assign n14401 = ~n14399 & n14400;
  assign n14402 = ~n13955 & n14354;
  assign n14403 = ~pi152 & pi197;
  assign n14404 = n14402 & n14403;
  assign n14405 = ~n14401 & ~n14404;
  assign n14406 = ~n14074 & ~n14405;
  assign n14407 = pi172 & ~n14371;
  assign n14408 = ~pi172 & n14359;
  assign n14409 = pi152 & pi197;
  assign n14410 = ~n14407 & n14409;
  assign n14411 = ~n14408 & n14410;
  assign n14412 = ~n14406 & ~n14411;
  assign n14413 = n9420 & ~n14412;
  assign n14414 = ~n13722 & n14402;
  assign n14415 = ~pi152 & ~n14074;
  assign n14416 = n14414 & n14415;
  assign n14417 = ~pi172 & n14386;
  assign n14418 = pi172 & n14378;
  assign n14419 = pi152 & ~n14418;
  assign n14420 = ~n14417 & n14419;
  assign n14421 = pi197 & ~n14416;
  assign n14422 = ~n14420 & n14421;
  assign n14423 = pi152 & ~n14380;
  assign n14424 = n13677 & n14365;
  assign n14425 = ~n14358 & ~n14424;
  assign n14426 = ~pi152 & n14425;
  assign n14427 = pi172 & ~n14426;
  assign n14428 = ~n14423 & n14427;
  assign n14429 = ~n13722 & ~n14353;
  assign n14430 = ~pi152 & ~n14429;
  assign n14431 = pi152 & n14384;
  assign n14432 = ~pi172 & ~n14430;
  assign n14433 = ~n14431 & n14432;
  assign n14434 = ~pi197 & ~n14428;
  assign n14435 = ~n14433 & n14434;
  assign n14436 = n9414 & ~n14435;
  assign n14437 = ~n14422 & n14436;
  assign n14438 = ~n14413 & ~n14437;
  assign n14439 = pi299 & ~n14438;
  assign n14440 = ~n14397 & ~n14439;
  assign n14441 = n8769 & ~n14440;
  assign n14442 = n14092 & ~n14349;
  assign n14443 = ~n14441 & n14442;
  assign n14444 = n2536 & ~n14090;
  assign n14445 = ~n14443 & n14444;
  assign n14446 = n13636 & ~n14089;
  assign n14447 = n14072 & ~n14260;
  assign n14448 = ~n14446 & n14447;
  assign n14449 = ~n14445 & n14448;
  assign n14450 = ~po1038 & ~n14264;
  assign n14451 = ~n14449 & n14450;
  assign po282 = n14082 | n14451;
  assign n14453 = pi175 & n13620;
  assign n14454 = n9927 & n13665;
  assign n14455 = ~pi299 & ~n14453;
  assign n14456 = ~n14454 & n14455;
  assign n14457 = ~pi51 & ~n13724;
  assign n14458 = pi153 & n13620;
  assign n14459 = ~n9931 & ~n13614;
  assign n14460 = ~pi51 & ~n14459;
  assign n14461 = ~n14458 & ~n14460;
  assign n14462 = ~n14457 & ~n14461;
  assign n14463 = pi299 & ~n14462;
  assign n14464 = pi232 & ~n14456;
  assign n14465 = ~n14463 & n14464;
  assign n14466 = n13636 & ~n14465;
  assign n14467 = ~pi150 & pi299;
  assign n14468 = ~pi185 & ~pi299;
  assign n14469 = ~n14467 & ~n14468;
  assign n14470 = n7406 & n14469;
  assign n14471 = pi87 & ~n14470;
  assign n14472 = ~n14466 & ~n14471;
  assign n14473 = ~pi126 & n13611;
  assign n14474 = pi126 & ~n13611;
  assign n14475 = ~n14473 & ~n14474;
  assign n14476 = ~n13607 & ~n14475;
  assign n14477 = n13616 & ~n14476;
  assign n14478 = ~n14472 & ~n14477;
  assign n14479 = ~n2613 & n14465;
  assign n14480 = ~n2613 & n13615;
  assign n14481 = ~n14476 & n14480;
  assign n14482 = ~pi160 & pi216;
  assign n14483 = n6590 & ~n14482;
  assign n14484 = ~n14463 & ~n14483;
  assign n14485 = n6333 & n11386;
  assign n14486 = ~pi166 & n13823;
  assign n14487 = ~pi153 & ~n14486;
  assign n14488 = ~n14485 & n14487;
  assign n14489 = ~pi166 & ~n14285;
  assign n14490 = pi166 & ~n14288;
  assign n14491 = pi153 & ~n14489;
  assign n14492 = ~n14490 & n14491;
  assign n14493 = pi160 & ~n14488;
  assign n14494 = ~n14492 & n14493;
  assign n14495 = pi216 & ~n14494;
  assign n14496 = ~pi166 & n14272;
  assign n14497 = pi51 & ~pi153;
  assign n14498 = pi166 & ~n14275;
  assign n14499 = ~n14496 & ~n14497;
  assign n14500 = ~n14498 & n14499;
  assign n14501 = ~pi216 & ~n14500;
  assign n14502 = n5726 & ~n14495;
  assign n14503 = ~n14501 & n14502;
  assign n14504 = ~n14484 & ~n14503;
  assign n14505 = ~pi189 & n14305;
  assign n14506 = pi189 & n14308;
  assign n14507 = ~pi182 & ~n14506;
  assign n14508 = ~n14505 & n14507;
  assign n14509 = ~pi189 & ~n14334;
  assign n14510 = pi189 & n14328;
  assign n14511 = pi182 & ~n14510;
  assign n14512 = ~n14509 & n14511;
  assign n14513 = ~n14508 & ~n14512;
  assign n14514 = n11402 & ~n14513;
  assign n14515 = ~n13620 & n14508;
  assign n14516 = ~pi189 & n14317;
  assign n14517 = pi189 & ~n14323;
  assign n14518 = pi182 & ~n14516;
  assign n14519 = ~n14517 & n14518;
  assign n14520 = ~n14515 & ~n14519;
  assign n14521 = n11373 & ~n14520;
  assign n14522 = ~n14504 & ~n14514;
  assign n14523 = ~n14521 & n14522;
  assign n14524 = pi232 & ~n14523;
  assign n14525 = n14268 & ~n14524;
  assign n14526 = ~pi153 & n14386;
  assign n14527 = pi153 & n14378;
  assign n14528 = pi157 & ~n14527;
  assign n14529 = ~n14526 & n14528;
  assign n14530 = ~pi153 & n14359;
  assign n14531 = pi153 & ~n14371;
  assign n14532 = ~pi157 & ~n14531;
  assign n14533 = ~n14530 & n14532;
  assign n14534 = ~n14529 & ~n14533;
  assign n14535 = pi166 & ~n14534;
  assign n14536 = pi157 & n13722;
  assign n14537 = ~pi166 & ~n14458;
  assign n14538 = ~n14536 & n14537;
  assign n14539 = n14402 & n14538;
  assign n14540 = ~n14535 & ~n14539;
  assign n14541 = n9599 & ~n14540;
  assign n14542 = ~pi166 & n14425;
  assign n14543 = pi166 & ~n14380;
  assign n14544 = pi153 & ~n14542;
  assign n14545 = ~n14543 & n14544;
  assign n14546 = ~pi166 & ~n14429;
  assign n14547 = pi166 & n14384;
  assign n14548 = ~pi153 & ~n14546;
  assign n14549 = ~n14547 & n14548;
  assign n14550 = ~n14545 & ~n14549;
  assign n14551 = pi157 & ~n14550;
  assign n14552 = pi166 & n13686;
  assign n14553 = ~pi166 & ~n14354;
  assign n14554 = ~pi157 & ~n14458;
  assign n14555 = ~n14552 & n14554;
  assign n14556 = ~n14553 & n14555;
  assign n14557 = ~n14551 & ~n14556;
  assign n14558 = n9573 & ~n14557;
  assign n14559 = ~pi189 & ~n14354;
  assign n14560 = pi189 & n13686;
  assign n14561 = ~pi178 & ~n14560;
  assign n14562 = ~n13620 & n14561;
  assign n14563 = ~n14559 & n14562;
  assign n14564 = ~pi181 & ~n14563;
  assign n14565 = pi189 & ~n14380;
  assign n14566 = ~pi189 & n14425;
  assign n14567 = pi178 & ~n14566;
  assign n14568 = ~n14565 & n14567;
  assign n14569 = n14564 & ~n14568;
  assign n14570 = pi189 & n14371;
  assign n14571 = ~pi189 & n14402;
  assign n14572 = ~n13620 & n14571;
  assign n14573 = ~n14570 & ~n14572;
  assign n14574 = ~pi178 & ~n14573;
  assign n14575 = ~pi189 & ~n14414;
  assign n14576 = ~n13620 & ~n13693;
  assign n14577 = ~pi189 & n14576;
  assign n14578 = n14378 & ~n14577;
  assign n14579 = pi178 & ~n14575;
  assign n14580 = ~n14578 & n14579;
  assign n14581 = pi181 & ~n14574;
  assign n14582 = ~n14580 & n14581;
  assign n14583 = n11373 & ~n14569;
  assign n14584 = ~n14582 & n14583;
  assign n14585 = n14354 & n14561;
  assign n14586 = pi189 & n14384;
  assign n14587 = ~pi189 & ~n14429;
  assign n14588 = pi178 & ~n14587;
  assign n14589 = ~n14586 & n14588;
  assign n14590 = n14564 & ~n14585;
  assign n14591 = ~n14589 & n14590;
  assign n14592 = pi189 & n14386;
  assign n14593 = ~n14575 & ~n14592;
  assign n14594 = pi178 & ~n14593;
  assign n14595 = pi189 & ~n14359;
  assign n14596 = ~pi178 & ~n14571;
  assign n14597 = ~n14595 & n14596;
  assign n14598 = ~n14594 & ~n14597;
  assign n14599 = pi181 & ~n14598;
  assign n14600 = n11402 & ~n14591;
  assign n14601 = ~n14599 & n14600;
  assign n14602 = ~n14558 & ~n14584;
  assign n14603 = ~n14541 & n14602;
  assign n14604 = ~n14601 & n14603;
  assign n14605 = pi232 & ~n14604;
  assign n14606 = n14347 & ~n14605;
  assign n14607 = n14476 & ~n14525;
  assign n14608 = ~n14606 & n14607;
  assign n14609 = pi178 & ~n13694;
  assign n14610 = ~n14577 & n14609;
  assign n14611 = pi189 & n14114;
  assign n14612 = ~pi189 & ~n13745;
  assign n14613 = n14576 & n14612;
  assign n14614 = ~pi178 & ~n14611;
  assign n14615 = ~n14613 & n14614;
  assign n14616 = pi181 & ~n14610;
  assign n14617 = ~n14615 & n14616;
  assign n14618 = ~n9927 & ~n13692;
  assign n14619 = ~pi189 & n13939;
  assign n14620 = ~n14618 & ~n14619;
  assign n14621 = ~pi178 & ~n14620;
  assign n14622 = ~pi189 & n14170;
  assign n14623 = pi189 & n14164;
  assign n14624 = pi178 & ~n14622;
  assign n14625 = ~n14623 & n14624;
  assign n14626 = ~pi181 & ~n14625;
  assign n14627 = ~n14610 & n14626;
  assign n14628 = ~n14621 & n14627;
  assign n14629 = n11402 & ~n14617;
  assign n14630 = ~n14628 & n14629;
  assign n14631 = n11386 & n13665;
  assign n14632 = ~n13693 & ~n14631;
  assign n14633 = pi153 & ~n14632;
  assign n14634 = ~pi153 & ~n14462;
  assign n14635 = ~n13694 & n14634;
  assign n14636 = pi157 & ~n14633;
  assign n14637 = ~n14635 & n14636;
  assign n14638 = pi166 & ~n14114;
  assign n14639 = pi51 & n9931;
  assign n14640 = ~n14638 & ~n14639;
  assign n14641 = ~pi153 & ~n14640;
  assign n14642 = ~pi166 & ~n14104;
  assign n14643 = pi153 & pi166;
  assign n14644 = ~n14135 & n14643;
  assign n14645 = ~pi157 & ~n14641;
  assign n14646 = ~n14644 & n14645;
  assign n14647 = ~n14642 & n14646;
  assign n14648 = n9599 & ~n14637;
  assign n14649 = ~n14647 & n14648;
  assign n14650 = ~pi189 & n14107;
  assign n14651 = pi189 & n14111;
  assign n14652 = ~pi178 & ~n14651;
  assign n14653 = ~n14650 & n14652;
  assign n14654 = n14626 & ~n14653;
  assign n14655 = pi178 & n11586;
  assign n14656 = n13665 & n14655;
  assign n14657 = pi189 & ~n13727;
  assign n14658 = ~pi178 & ~n14657;
  assign n14659 = ~n14612 & n14658;
  assign n14660 = pi181 & ~n14656;
  assign n14661 = ~n13693 & n14660;
  assign n14662 = ~n14659 & n14661;
  assign n14663 = n11373 & ~n14662;
  assign n14664 = ~n14654 & n14663;
  assign n14665 = ~n14164 & n14643;
  assign n14666 = pi166 & ~n14166;
  assign n14667 = ~n14639 & ~n14666;
  assign n14668 = ~pi153 & ~n14667;
  assign n14669 = ~pi166 & ~n14170;
  assign n14670 = pi157 & ~n14665;
  assign n14671 = ~n14669 & n14670;
  assign n14672 = ~n14668 & n14671;
  assign n14673 = pi166 & ~n14111;
  assign n14674 = ~pi166 & ~n14107;
  assign n14675 = pi153 & ~n14673;
  assign n14676 = ~n14674 & n14675;
  assign n14677 = ~pi166 & n13939;
  assign n14678 = ~n9931 & ~n13692;
  assign n14679 = ~pi153 & ~n14678;
  assign n14680 = ~n14677 & n14679;
  assign n14681 = ~n14676 & ~n14680;
  assign n14682 = ~pi157 & ~n14681;
  assign n14683 = n9573 & ~n14672;
  assign n14684 = ~n14682 & n14683;
  assign n14685 = ~n14649 & ~n14664;
  assign n14686 = ~n14630 & n14685;
  assign n14687 = ~n14684 & n14686;
  assign n14688 = pi232 & ~n14687;
  assign n14689 = n14249 & ~n14688;
  assign n14690 = pi189 & ~n14227;
  assign n14691 = ~pi189 & ~n14225;
  assign n14692 = ~pi182 & ~n14690;
  assign n14693 = ~n14691 & n14692;
  assign n14694 = pi189 & ~n14237;
  assign n14695 = ~pi189 & ~n14233;
  assign n14696 = pi182 & ~n14694;
  assign n14697 = ~n14695 & n14696;
  assign n14698 = ~n14693 & ~n14697;
  assign n14699 = n11373 & ~n14698;
  assign n14700 = pi182 & n13876;
  assign n14701 = pi189 & ~n14182;
  assign n14702 = ~n14700 & n14701;
  assign n14703 = pi182 & n13847;
  assign n14704 = ~pi189 & ~n14703;
  assign n14705 = n14215 & n14704;
  assign n14706 = ~n14702 & ~n14705;
  assign n14707 = n11402 & ~n14706;
  assign n14708 = ~n8739 & ~n14461;
  assign n14709 = ~pi166 & ~n13848;
  assign n14710 = pi166 & n13876;
  assign n14711 = pi160 & ~n14458;
  assign n14712 = ~n14710 & n14711;
  assign n14713 = ~n14709 & n14712;
  assign n14714 = ~pi166 & n13841;
  assign n14715 = ~n9931 & ~n13818;
  assign n14716 = ~pi153 & ~n14715;
  assign n14717 = ~n14714 & n14716;
  assign n14718 = ~pi166 & ~n13837;
  assign n14719 = pi166 & ~n13831;
  assign n14720 = pi153 & ~n14719;
  assign n14721 = ~n14718 & n14720;
  assign n14722 = ~pi160 & ~n14717;
  assign n14723 = ~n14721 & n14722;
  assign n14724 = n8739 & ~n14713;
  assign n14725 = ~n14723 & n14724;
  assign n14726 = pi299 & ~n14708;
  assign n14727 = ~n14725 & n14726;
  assign n14728 = ~n14707 & ~n14727;
  assign n14729 = ~n14699 & n14728;
  assign n14730 = pi232 & ~n14729;
  assign n14731 = n14189 & ~n14730;
  assign n14732 = ~n14476 & ~n14731;
  assign n14733 = ~n14689 & n14732;
  assign n14734 = n2613 & ~n14733;
  assign n14735 = ~n14608 & n14734;
  assign n14736 = n2536 & ~n14481;
  assign n14737 = ~n14479 & n14736;
  assign n14738 = ~n14735 & n14737;
  assign n14739 = ~po1038 & ~n14478;
  assign n14740 = ~n14738 & n14739;
  assign n14741 = pi87 & ~n12938;
  assign n14742 = pi232 & ~n14457;
  assign n14743 = n14476 & ~n14742;
  assign n14744 = ~pi232 & ~n13615;
  assign n14745 = ~n14461 & ~n14744;
  assign n14746 = ~n14743 & n14745;
  assign n14747 = ~pi87 & ~n14746;
  assign n14748 = po1038 & ~n14741;
  assign n14749 = ~n14747 & n14748;
  assign po283 = ~n14740 & ~n14749;
  assign n14751 = ~pi129 & ~n3291;
  assign n14752 = n2538 & n8602;
  assign n14753 = ~n2530 & ~n14752;
  assign n14754 = pi129 & n7228;
  assign n14755 = n6276 & n14754;
  assign n14756 = pi74 & ~n14755;
  assign n14757 = pi54 & n2616;
  assign n14758 = n8602 & n14757;
  assign n14759 = pi92 & ~pi129;
  assign n14760 = pi75 & n14754;
  assign n14761 = ~n2628 & ~n8669;
  assign n14762 = n8602 & ~n14761;
  assign n14763 = ~n2573 & ~n14762;
  assign n14764 = pi129 & n6116;
  assign n14765 = pi38 & ~n14764;
  assign n14766 = pi39 & n8602;
  assign n14767 = ~n2728 & ~n3088;
  assign n14768 = n2786 & ~n2860;
  assign n14769 = n2464 & ~n14768;
  assign n14770 = n2873 & ~n14769;
  assign n14771 = n2783 & ~n14770;
  assign n14772 = n2877 & ~n14771;
  assign n14773 = n2719 & ~n14772;
  assign n14774 = ~n2722 & ~n14773;
  assign n14775 = ~pi86 & ~n14774;
  assign n14776 = n2780 & ~n14775;
  assign n14777 = pi250 & n12425;
  assign n14778 = ~pi127 & ~n14777;
  assign n14779 = po740 & n14777;
  assign n14780 = ~n14778 & ~n14779;
  assign n14781 = n2777 & n14780;
  assign n14782 = ~pi97 & ~n14781;
  assign n14783 = ~n14776 & n14782;
  assign n14784 = ~n2775 & ~n14783;
  assign n14785 = ~pi108 & ~n14784;
  assign n14786 = n2774 & ~n14785;
  assign n14787 = n2890 & ~n14786;
  assign n14788 = ~n2766 & ~n14787;
  assign n14789 = n2765 & ~n14788;
  assign n14790 = n2764 & ~n14789;
  assign n14791 = n2757 & ~n14790;
  assign n14792 = n3090 & ~n14791;
  assign n14793 = n2516 & ~n14792;
  assign n14794 = n14767 & ~n14793;
  assign n14795 = ~pi70 & ~n14794;
  assign n14796 = ~n3081 & ~n14795;
  assign n14797 = ~pi51 & ~n14796;
  assign n14798 = n2748 & ~n14797;
  assign n14799 = n3149 & ~n14798;
  assign n14800 = ~n2744 & ~n14799;
  assign n14801 = n2462 & ~n14800;
  assign n14802 = n3389 & ~n14801;
  assign n14803 = ~pi95 & ~n14802;
  assign n14804 = ~pi39 & pi129;
  assign n14805 = ~n2740 & n14804;
  assign n14806 = ~n14803 & n14805;
  assign n14807 = ~pi38 & ~n14766;
  assign n14808 = ~n14806 & n14807;
  assign n14809 = ~n14765 & ~n14808;
  assign n14810 = n2573 & ~n14809;
  assign n14811 = ~pi75 & ~n14763;
  assign n14812 = ~n14810 & n14811;
  assign n14813 = ~pi92 & ~n14760;
  assign n14814 = ~n14812 & n14813;
  assign n14815 = n12909 & ~n14759;
  assign n14816 = ~n14814 & n14815;
  assign n14817 = ~pi74 & ~n14758;
  assign n14818 = ~n14816 & n14817;
  assign n14819 = ~pi55 & ~n14756;
  assign n14820 = ~n14818 & n14819;
  assign n14821 = pi55 & n7293;
  assign n14822 = n14754 & n14821;
  assign n14823 = ~n14820 & ~n14822;
  assign n14824 = ~pi56 & ~n14823;
  assign n14825 = ~n10897 & ~n10905;
  assign n14826 = ~n14824 & n14825;
  assign n14827 = ~n14753 & ~n14826;
  assign n14828 = n3291 & ~n14827;
  assign n14829 = n6071 & ~n14751;
  assign po284 = ~n14828 & n14829;
  assign n14831 = ~n6076 & ~n7277;
  assign n14832 = ~pi38 & ~n3394;
  assign n14833 = n6118 & ~n14832;
  assign n14834 = n6310 & n8606;
  assign n14835 = ~pi87 & ~n14834;
  assign n14836 = ~n14833 & n14835;
  assign n14837 = n6080 & ~n14836;
  assign n14838 = ~pi250 & n12425;
  assign n14839 = ~pi129 & ~n14838;
  assign n14840 = po740 & n14838;
  assign n14841 = n8671 & ~n14839;
  assign n14842 = ~n14840 & n14841;
  assign n14843 = n2523 & n14842;
  assign n14844 = n6078 & ~n14843;
  assign n14845 = ~n14837 & n14844;
  assign n14846 = ~n7234 & ~n7271;
  assign n14847 = ~n14845 & n14846;
  assign n14848 = n6246 & ~n14847;
  assign n14849 = n14831 & ~n14848;
  assign n14850 = ~pi56 & ~n14849;
  assign n14851 = ~n6248 & ~n14850;
  assign n14852 = ~pi62 & ~n14851;
  assign n14853 = ~n6252 & ~n14852;
  assign n14854 = n3291 & ~n14853;
  assign po286 = n6071 & ~n14854;
  assign n14856 = ~pi132 & n14473;
  assign n14857 = pi130 & ~n14856;
  assign n14858 = ~pi130 & n14856;
  assign n14859 = ~n14857 & ~n14858;
  assign n14860 = ~n13605 & ~n14859;
  assign n14861 = pi87 & ~n9409;
  assign n14862 = n7406 & ~n8724;
  assign n14863 = n13665 & ~n14862;
  assign n14864 = ~n14457 & ~n14863;
  assign n14865 = n13636 & ~n14864;
  assign n14866 = ~n14861 & ~n14865;
  assign n14867 = ~n13616 & ~n14866;
  assign n14868 = pi100 & n14864;
  assign n14869 = ~n10584 & n14863;
  assign n14870 = ~pi51 & ~n14187;
  assign n14871 = ~pi232 & ~n14870;
  assign n14872 = n10584 & ~n14871;
  assign n14873 = pi140 & n13821;
  assign n14874 = ~pi51 & ~n13842;
  assign n14875 = ~n14214 & n14874;
  assign n14876 = ~n14873 & n14875;
  assign n14877 = n8722 & ~n14876;
  assign n14878 = ~pi191 & ~pi299;
  assign n14879 = ~pi51 & ~n14182;
  assign n14880 = pi140 & n14236;
  assign n14881 = n14879 & ~n14880;
  assign n14882 = n14878 & ~n14881;
  assign n14883 = pi169 & n6166;
  assign n14884 = ~n8739 & n13665;
  assign n14885 = ~n14883 & n14884;
  assign n14886 = pi162 & n8739;
  assign n14887 = ~n13821 & n14874;
  assign n14888 = pi169 & ~n14887;
  assign n14889 = ~pi169 & ~n14235;
  assign n14890 = n14886 & ~n14889;
  assign n14891 = ~n14888 & n14890;
  assign n14892 = ~n13819 & ~n14883;
  assign n14893 = ~n2523 & n14883;
  assign n14894 = ~pi162 & n8739;
  assign n14895 = ~n14892 & n14894;
  assign n14896 = ~n14893 & n14895;
  assign n14897 = pi299 & ~n14885;
  assign n14898 = ~n14896 & n14897;
  assign n14899 = ~n14891 & n14898;
  assign n14900 = ~n14877 & ~n14882;
  assign n14901 = ~n14899 & n14900;
  assign n14902 = pi232 & ~n14901;
  assign n14903 = n14872 & ~n14902;
  assign n14904 = ~pi100 & ~n14869;
  assign n14905 = ~n14903 & n14904;
  assign n14906 = n13898 & ~n14868;
  assign n14907 = ~n14905 & n14906;
  assign n14908 = ~n14860 & ~n14867;
  assign n14909 = ~n14907 & n14908;
  assign n14910 = pi38 & ~n14864;
  assign n14911 = ~n13840 & ~n14883;
  assign n14912 = pi169 & n14271;
  assign n14913 = ~n14911 & ~n14912;
  assign n14914 = ~pi216 & ~n14913;
  assign n14915 = ~n13830 & n14285;
  assign n14916 = pi169 & n14915;
  assign n14917 = ~pi51 & ~n14287;
  assign n14918 = ~pi169 & n14917;
  assign n14919 = pi162 & pi216;
  assign n14920 = ~n14916 & n14919;
  assign n14921 = ~n14918 & n14920;
  assign n14922 = ~n14914 & ~n14921;
  assign n14923 = n5726 & ~n14922;
  assign n14924 = pi169 & n13724;
  assign n14925 = ~pi51 & ~n14924;
  assign n14926 = ~n5727 & ~n14886;
  assign n14927 = ~n14925 & n14926;
  assign n14928 = ~n14923 & ~n14927;
  assign n14929 = pi299 & ~n14928;
  assign n14930 = ~pi51 & ~n14307;
  assign n14931 = ~pi140 & n14930;
  assign n14932 = n13839 & n14320;
  assign n14933 = ~pi51 & ~n14932;
  assign n14934 = pi140 & n14933;
  assign n14935 = n14878 & ~n14931;
  assign n14936 = ~n14934 & n14935;
  assign n14937 = ~pi51 & ~n14305;
  assign n14938 = ~pi140 & n14937;
  assign n14939 = ~pi51 & n14334;
  assign n14940 = pi140 & n14939;
  assign n14941 = n8722 & ~n14938;
  assign n14942 = ~n14940 & n14941;
  assign n14943 = ~n14929 & ~n14936;
  assign n14944 = ~n14942 & n14943;
  assign n14945 = pi232 & ~n14944;
  assign n14946 = ~pi51 & ~n14266;
  assign n14947 = ~pi232 & ~n14946;
  assign n14948 = pi39 & ~n14947;
  assign n14949 = ~n14945 & n14948;
  assign n14950 = ~pi232 & ~n13763;
  assign n14951 = ~pi39 & ~n14950;
  assign n14952 = ~n6166 & n13763;
  assign n14953 = n6166 & n13684;
  assign n14954 = ~n14952 & ~n14953;
  assign n14955 = ~n8724 & ~n14954;
  assign n14956 = n8724 & n13763;
  assign n14957 = pi232 & ~n14956;
  assign n14958 = ~n14955 & n14957;
  assign n14959 = n14951 & ~n14958;
  assign n14960 = ~n14949 & ~n14959;
  assign n14961 = ~pi38 & ~n14960;
  assign n14962 = ~pi100 & ~n14910;
  assign n14963 = ~n14961 & n14962;
  assign n14964 = n2536 & ~n14868;
  assign n14965 = ~n14963 & n14964;
  assign n14966 = n14860 & n14866;
  assign n14967 = ~n14965 & n14966;
  assign n14968 = ~n14909 & ~n14967;
  assign n14969 = ~po1038 & ~n14968;
  assign n14970 = pi87 & ~n9514;
  assign n14971 = ~pi51 & ~pi87;
  assign n14972 = ~n13614 & n14971;
  assign n14973 = ~n8698 & n14972;
  assign n14974 = ~n14924 & n14971;
  assign n14975 = n14860 & n14974;
  assign n14976 = po1038 & ~n14970;
  assign n14977 = ~n14973 & n14976;
  assign n14978 = ~n14975 & n14977;
  assign po287 = ~n14969 & ~n14978;
  assign n14980 = ~pi100 & ~n13245;
  assign n14981 = n7238 & ~n14980;
  assign n14982 = ~pi75 & ~n14981;
  assign n14983 = ~n7229 & ~n14982;
  assign n14984 = ~pi92 & ~n14983;
  assign n14985 = ~n7234 & n12403;
  assign po288 = ~n14984 & n14985;
  assign n14987 = pi132 & ~n14473;
  assign n14988 = ~n14856 & ~n14987;
  assign n14989 = ~n13606 & ~n14988;
  assign n14990 = pi87 & ~n8732;
  assign n14991 = pi190 & n13724;
  assign n14992 = pi173 & n13620;
  assign n14993 = ~pi299 & ~n14992;
  assign n14994 = ~n14991 & n14993;
  assign n14995 = pi51 & ~pi151;
  assign n14996 = ~n12989 & ~n13620;
  assign n14997 = ~n14995 & ~n14996;
  assign n14998 = n13619 & n14997;
  assign n14999 = pi299 & ~n14998;
  assign n15000 = pi232 & ~n14994;
  assign n15001 = ~n14999 & n15000;
  assign n15002 = ~n2613 & n15001;
  assign n15003 = n2536 & ~n15002;
  assign n15004 = pi190 & ~pi299;
  assign n15005 = ~pi183 & n14302;
  assign n15006 = ~pi183 & ~n14304;
  assign n15007 = pi183 & ~n14334;
  assign n15008 = ~pi173 & ~n15006;
  assign n15009 = ~n15007 & n15008;
  assign n15010 = ~pi183 & ~n14313;
  assign n15011 = pi173 & ~n14317;
  assign n15012 = ~n15010 & n15011;
  assign n15013 = ~n15005 & ~n15012;
  assign n15014 = ~n15009 & n15013;
  assign n15015 = n15004 & ~n15014;
  assign n15016 = ~pi149 & pi216;
  assign n15017 = n6590 & ~n15016;
  assign n15018 = ~n14999 & ~n15017;
  assign n15019 = ~pi168 & ~n14275;
  assign n15020 = pi168 & n14272;
  assign n15021 = ~n14995 & ~n15019;
  assign n15022 = ~n15020 & n15021;
  assign n15023 = ~pi216 & ~n15022;
  assign n15024 = ~pi168 & n13908;
  assign n15025 = pi168 & n13823;
  assign n15026 = ~pi151 & ~n15025;
  assign n15027 = ~n15024 & n15026;
  assign n15028 = pi168 & ~n14285;
  assign n15029 = ~pi168 & ~n14288;
  assign n15030 = pi151 & ~n15028;
  assign n15031 = ~n15029 & n15030;
  assign n15032 = pi149 & ~n15027;
  assign n15033 = ~n15031 & n15032;
  assign n15034 = pi216 & ~n15033;
  assign n15035 = n5726 & ~n15023;
  assign n15036 = ~n15034 & n15035;
  assign n15037 = ~n15018 & ~n15036;
  assign n15038 = ~pi183 & ~n7506;
  assign n15039 = ~pi173 & ~n15038;
  assign n15040 = n14328 & n15039;
  assign n15041 = ~pi190 & ~pi299;
  assign n15042 = ~pi183 & ~n13620;
  assign n15043 = ~n14308 & n15042;
  assign n15044 = pi183 & n14323;
  assign n15045 = pi173 & ~n15043;
  assign n15046 = ~n15044 & n15045;
  assign n15047 = ~n15040 & n15041;
  assign n15048 = ~n15046 & n15047;
  assign n15049 = ~n15015 & ~n15037;
  assign n15050 = ~n15048 & n15049;
  assign n15051 = pi232 & ~n15050;
  assign n15052 = n14268 & ~n15051;
  assign n15053 = ~pi232 & ~n13741;
  assign n15054 = ~n6166 & n13741;
  assign n15055 = pi182 & n13664;
  assign n15056 = n13683 & ~n15055;
  assign n15057 = pi51 & ~pi173;
  assign n15058 = n6166 & ~n15057;
  assign n15059 = ~n15056 & n15058;
  assign n15060 = n15004 & ~n15059;
  assign n15061 = ~pi173 & ~n13741;
  assign n15062 = pi173 & n13746;
  assign n15063 = ~pi182 & ~n15061;
  assign n15064 = ~n15062 & n15063;
  assign n15065 = ~pi173 & ~n13756;
  assign n15066 = pi173 & n13763;
  assign n15067 = pi182 & n6166;
  assign n15068 = ~n15065 & n15067;
  assign n15069 = ~n15066 & n15068;
  assign n15070 = n15041 & ~n15064;
  assign n15071 = ~n15069 & n15070;
  assign n15072 = ~n15060 & ~n15071;
  assign n15073 = ~n15054 & ~n15072;
  assign n15074 = ~n6166 & ~n13741;
  assign n15075 = pi168 & ~n14995;
  assign n15076 = ~n13684 & n15075;
  assign n15077 = pi151 & n13763;
  assign n15078 = ~pi151 & ~n13756;
  assign n15079 = ~pi168 & ~n15077;
  assign n15080 = ~n15078 & n15079;
  assign n15081 = n6166 & ~n15076;
  assign n15082 = ~n15080 & n15081;
  assign n15083 = pi160 & ~n15074;
  assign n15084 = ~n15082 & n15083;
  assign n15085 = pi168 & ~n14424;
  assign n15086 = ~n15074 & n15085;
  assign n15087 = n13746 & ~n15054;
  assign n15088 = ~pi168 & ~n15087;
  assign n15089 = pi151 & ~n15086;
  assign n15090 = ~n15088 & n15089;
  assign n15091 = ~n12989 & n13741;
  assign n15092 = pi168 & n13722;
  assign n15093 = ~pi151 & ~n15092;
  assign n15094 = ~n15091 & n15093;
  assign n15095 = ~pi160 & ~n15094;
  assign n15096 = ~n15090 & n15095;
  assign n15097 = pi299 & ~n15096;
  assign n15098 = ~n15084 & n15097;
  assign n15099 = ~n15073 & ~n15098;
  assign n15100 = pi232 & ~n15099;
  assign n15101 = ~pi39 & ~n15053;
  assign n15102 = ~n15100 & n15101;
  assign n15103 = ~n15052 & ~n15102;
  assign n15104 = n2613 & ~n15103;
  assign n15105 = n15003 & ~n15104;
  assign n15106 = n13636 & ~n15001;
  assign n15107 = n14989 & ~n14990;
  assign n15108 = ~n15106 & n15107;
  assign n15109 = ~n15105 & n15108;
  assign n15110 = ~pi183 & ~n14225;
  assign n15111 = pi183 & ~n14233;
  assign n15112 = pi173 & ~n15111;
  assign n15113 = ~n15110 & n15112;
  assign n15114 = pi183 & n13847;
  assign n15115 = ~pi173 & ~n15114;
  assign n15116 = n14215 & n15115;
  assign n15117 = ~n15113 & ~n15116;
  assign n15118 = n15004 & ~n15117;
  assign n15119 = ~n13615 & n14999;
  assign n15120 = ~n12407 & ~n15119;
  assign n15121 = pi168 & n13841;
  assign n15122 = ~n12989 & ~n13818;
  assign n15123 = ~pi151 & ~n15122;
  assign n15124 = ~n15121 & n15123;
  assign n15125 = pi168 & ~n13837;
  assign n15126 = ~pi168 & ~n13831;
  assign n15127 = pi151 & ~n15126;
  assign n15128 = ~n15125 & n15127;
  assign n15129 = ~pi149 & ~n15124;
  assign n15130 = ~n15128 & n15129;
  assign n15131 = ~pi151 & n13620;
  assign n15132 = pi168 & ~n15131;
  assign n15133 = n14231 & n15132;
  assign n15134 = ~n13876 & ~n14997;
  assign n15135 = ~pi168 & ~n15134;
  assign n15136 = pi149 & ~n15135;
  assign n15137 = ~n15133 & n15136;
  assign n15138 = n8739 & ~n15137;
  assign n15139 = ~n15130 & n15138;
  assign n15140 = ~n15120 & ~n15139;
  assign n15141 = pi183 & n13876;
  assign n15142 = ~n14992 & n15041;
  assign n15143 = ~n14182 & n15142;
  assign n15144 = ~n15141 & n15143;
  assign n15145 = ~n15140 & ~n15144;
  assign n15146 = ~n15118 & n15145;
  assign n15147 = pi232 & ~n15146;
  assign n15148 = ~n14188 & ~n15147;
  assign n15149 = pi39 & ~n15148;
  assign n15150 = pi182 & n14113;
  assign n15151 = ~n13691 & n15142;
  assign n15152 = ~n15150 & n15151;
  assign n15153 = ~pi182 & n13704;
  assign n15154 = ~n14112 & ~n15057;
  assign n15155 = ~n15153 & n15154;
  assign n15156 = n15004 & ~n15155;
  assign n15157 = ~pi168 & n13724;
  assign n15158 = ~n14112 & ~n15157;
  assign n15159 = pi151 & ~n15158;
  assign n15160 = ~pi151 & ~n14998;
  assign n15161 = ~n14113 & n15160;
  assign n15162 = pi160 & ~n15159;
  assign n15163 = ~n15161 & n15162;
  assign n15164 = ~n13704 & n15132;
  assign n15165 = pi151 & n13955;
  assign n15166 = ~pi151 & ~n13691;
  assign n15167 = ~pi168 & ~n15166;
  assign n15168 = ~n15165 & n15167;
  assign n15169 = ~n15164 & ~n15168;
  assign n15170 = ~pi160 & ~n14112;
  assign n15171 = ~n15169 & n15170;
  assign n15172 = pi299 & ~n15163;
  assign n15173 = ~n15171 & n15172;
  assign n15174 = pi232 & ~n15152;
  assign n15175 = ~n15156 & n15174;
  assign n15176 = ~n15173 & n15175;
  assign n15177 = ~pi232 & n13691;
  assign n15178 = ~pi39 & ~n15177;
  assign n15179 = ~n15176 & n15178;
  assign n15180 = n2613 & ~n15179;
  assign n15181 = ~n15149 & n15180;
  assign n15182 = ~n14480 & n15003;
  assign n15183 = ~n15181 & n15182;
  assign n15184 = n13637 & ~n15001;
  assign n15185 = ~n14989 & ~n14990;
  assign n15186 = ~n15184 & n15185;
  assign n15187 = ~n15183 & n15186;
  assign n15188 = ~po1038 & ~n15187;
  assign n15189 = ~n15109 & n15188;
  assign n15190 = pi232 & n14998;
  assign n15191 = n13615 & ~n14989;
  assign n15192 = ~n15190 & ~n15191;
  assign n15193 = ~pi87 & ~n15192;
  assign n15194 = po1038 & ~n8920;
  assign n15195 = ~n15193 & n15194;
  assign po289 = n15189 | n15195;
  assign n15197 = ~pi183 & ~pi299;
  assign n15198 = ~pi149 & pi299;
  assign n15199 = ~n15197 & ~n15198;
  assign n15200 = n7406 & n15199;
  assign n15201 = pi87 & ~n15200;
  assign n15202 = ~pi133 & ~n14069;
  assign n15203 = ~n8896 & n13676;
  assign n15204 = ~pi39 & n13615;
  assign n15205 = ~n15203 & n15204;
  assign n15206 = pi145 & n13876;
  assign n15207 = n14183 & ~n15206;
  assign n15208 = pi197 & n13821;
  assign n15209 = n14184 & ~n15208;
  assign n15210 = n13615 & ~n15209;
  assign n15211 = pi299 & ~n15210;
  assign n15212 = ~n15207 & ~n15211;
  assign n15213 = pi232 & ~n15212;
  assign n15214 = n14189 & ~n15213;
  assign n15215 = ~pi38 & ~n15205;
  assign n15216 = ~n15214 & n15215;
  assign n15217 = n13651 & ~n15216;
  assign n15218 = n13898 & ~n15217;
  assign n15219 = ~n13637 & ~n15218;
  assign n15220 = ~n15202 & ~n15219;
  assign n15221 = pi299 & n8894;
  assign n15222 = n13709 & ~n15221;
  assign n15223 = n8893 & ~n15222;
  assign n15224 = ~n6166 & ~n13709;
  assign n15225 = n8894 & ~n15224;
  assign n15226 = ~n15223 & n15225;
  assign n15227 = ~n13757 & n15226;
  assign n15228 = ~n8893 & n8894;
  assign n15229 = n13709 & ~n15228;
  assign n15230 = ~n15227 & ~n15229;
  assign n15231 = ~pi39 & ~n15230;
  assign n15232 = ~n5724 & ~n15208;
  assign n15233 = n6590 & ~n15232;
  assign n15234 = ~pi145 & ~n7506;
  assign n15235 = ~pi299 & ~n15234;
  assign n15236 = ~n14327 & n15235;
  assign n15237 = ~n15233 & ~n15236;
  assign n15238 = n2523 & ~n15237;
  assign n15239 = pi232 & ~n15238;
  assign n15240 = n14268 & ~n15239;
  assign n15241 = ~n15231 & ~n15240;
  assign n15242 = n10958 & ~n15241;
  assign n15243 = ~pi87 & n15202;
  assign n15244 = ~n15242 & n15243;
  assign n15245 = ~n15201 & ~n15220;
  assign n15246 = ~n15244 & n15245;
  assign n15247 = ~po1038 & ~n15246;
  assign n15248 = pi87 & n8913;
  assign n15249 = n13616 & ~n15202;
  assign n15250 = po1038 & ~n15248;
  assign n15251 = ~n15249 & n15250;
  assign po290 = n15247 | n15251;
  assign n15253 = po1038 & n14971;
  assign n15254 = ~pi136 & n14858;
  assign n15255 = ~pi135 & n15254;
  assign n15256 = pi134 & ~n15255;
  assign n15257 = n13614 & ~n15256;
  assign n15258 = pi171 & n6166;
  assign n15259 = ~n13614 & n15258;
  assign n15260 = pi232 & n15259;
  assign n15261 = n15253 & ~n15260;
  assign n15262 = ~n15257 & n15261;
  assign n15263 = pi192 & ~pi299;
  assign n15264 = pi171 & pi299;
  assign n15265 = ~n15263 & ~n15264;
  assign n15266 = n7406 & ~n15265;
  assign n15267 = n13665 & ~n15266;
  assign n15268 = ~n14457 & ~n15267;
  assign n15269 = n13636 & ~n15268;
  assign n15270 = ~n2613 & n15268;
  assign n15271 = n2536 & ~n15270;
  assign n15272 = pi232 & ~n15265;
  assign n15273 = ~n13763 & ~n15272;
  assign n15274 = n14954 & n15272;
  assign n15275 = ~pi39 & ~n15273;
  assign n15276 = ~n15274 & n15275;
  assign n15277 = ~pi51 & ~n15259;
  assign n15278 = ~pi164 & pi216;
  assign n15279 = n5726 & ~n15278;
  assign n15280 = ~n15277 & ~n15279;
  assign n15281 = ~n13840 & ~n15258;
  assign n15282 = pi171 & n14271;
  assign n15283 = ~n15281 & ~n15282;
  assign n15284 = ~pi216 & ~n15283;
  assign n15285 = pi171 & n14915;
  assign n15286 = ~pi171 & n14917;
  assign n15287 = pi164 & pi216;
  assign n15288 = ~n15285 & n15287;
  assign n15289 = ~n15286 & n15288;
  assign n15290 = ~n15284 & ~n15289;
  assign n15291 = n5726 & ~n15290;
  assign n15292 = ~n15280 & ~n15291;
  assign n15293 = pi299 & ~n15292;
  assign n15294 = ~n14937 & n15263;
  assign n15295 = pi39 & pi186;
  assign n15296 = ~pi192 & ~pi299;
  assign n15297 = ~n14930 & n15296;
  assign n15298 = ~n15295 & ~n15297;
  assign n15299 = ~n15294 & n15298;
  assign n15300 = ~n14939 & n15263;
  assign n15301 = ~n14933 & n15296;
  assign n15302 = pi186 & ~n15300;
  assign n15303 = ~n15301 & n15302;
  assign n15304 = ~n15299 & ~n15303;
  assign n15305 = ~n15293 & ~n15304;
  assign n15306 = pi232 & ~n15305;
  assign n15307 = n14948 & ~n15306;
  assign n15308 = n2613 & ~n15276;
  assign n15309 = ~n15307 & n15308;
  assign n15310 = n15271 & ~n15309;
  assign n15311 = n15256 & ~n15269;
  assign n15312 = ~n15310 & n15311;
  assign n15313 = n13636 & n15267;
  assign n15314 = ~n14214 & n14887;
  assign n15315 = n15263 & ~n15314;
  assign n15316 = ~n14236 & n14879;
  assign n15317 = n15296 & ~n15316;
  assign n15318 = ~n15315 & ~n15317;
  assign n15319 = n14884 & ~n15258;
  assign n15320 = pi299 & ~n15319;
  assign n15321 = ~n13819 & ~n15258;
  assign n15322 = n4156 & n6166;
  assign n15323 = n8739 & ~n15321;
  assign n15324 = ~n15322 & n15323;
  assign n15325 = n15320 & ~n15324;
  assign n15326 = n15318 & ~n15325;
  assign n15327 = pi232 & ~n15326;
  assign n15328 = ~n14871 & ~n15327;
  assign n15329 = n15295 & ~n15328;
  assign n15330 = ~pi39 & ~n15267;
  assign n15331 = pi39 & ~pi186;
  assign n15332 = ~n14875 & n15263;
  assign n15333 = ~n14879 & n15296;
  assign n15334 = ~n15332 & ~n15333;
  assign n15335 = ~n15325 & n15334;
  assign n15336 = pi232 & ~n15335;
  assign n15337 = ~n14871 & ~n15336;
  assign n15338 = n15331 & ~n15337;
  assign n15339 = ~pi164 & ~n15330;
  assign n15340 = ~n15338 & n15339;
  assign n15341 = ~n15329 & n15340;
  assign n15342 = n15295 & ~n15318;
  assign n15343 = n15331 & ~n15334;
  assign n15344 = ~n15342 & ~n15343;
  assign n15345 = pi232 & ~n15344;
  assign n15346 = pi171 & ~n14887;
  assign n15347 = ~pi171 & ~n14235;
  assign n15348 = n8739 & ~n15347;
  assign n15349 = ~n15346 & n15348;
  assign n15350 = pi232 & n15320;
  assign n15351 = ~n15349 & n15350;
  assign n15352 = ~n14871 & ~n15351;
  assign n15353 = pi39 & ~n15352;
  assign n15354 = pi164 & ~n15330;
  assign n15355 = ~n15353 & n15354;
  assign n15356 = ~n15345 & n15355;
  assign n15357 = n2613 & ~n15356;
  assign n15358 = ~n15341 & n15357;
  assign n15359 = ~n14480 & n15271;
  assign n15360 = ~n15358 & n15359;
  assign n15361 = ~n15256 & ~n15313;
  assign n15362 = ~n15360 & n15361;
  assign n15363 = ~po1038 & ~n15312;
  assign n15364 = ~n15362 & n15363;
  assign po291 = n15262 | n15364;
  assign n15366 = pi135 & ~n15254;
  assign n15367 = pi134 & n15255;
  assign n15368 = ~n15366 & ~n15367;
  assign n15369 = pi170 & n6166;
  assign n15370 = n10277 & n15369;
  assign n15371 = n13665 & ~n15370;
  assign n15372 = pi194 & n8878;
  assign n15373 = n15371 & ~n15372;
  assign n15374 = n13636 & n15373;
  assign n15375 = pi185 & n14236;
  assign n15376 = n14879 & ~n15375;
  assign n15377 = ~n10584 & n15371;
  assign n15378 = ~pi194 & ~n15377;
  assign n15379 = ~n15376 & n15378;
  assign n15380 = pi170 & n7406;
  assign n15381 = ~n8878 & ~n15380;
  assign n15382 = n13665 & n15381;
  assign n15383 = ~n10584 & n15382;
  assign n15384 = pi194 & ~n15383;
  assign n15385 = ~pi185 & n14875;
  assign n15386 = ~n15314 & n15384;
  assign n15387 = ~n15385 & n15386;
  assign n15388 = ~n15379 & ~n15387;
  assign n15389 = ~pi299 & ~n15388;
  assign n15390 = n14884 & ~n15369;
  assign n15391 = pi150 & pi299;
  assign n15392 = pi170 & ~n14887;
  assign n15393 = ~pi170 & ~n14235;
  assign n15394 = n8739 & ~n15393;
  assign n15395 = ~n15392 & n15394;
  assign n15396 = n15391 & ~n15395;
  assign n15397 = ~n13819 & ~n15369;
  assign n15398 = n4378 & n6166;
  assign n15399 = n8739 & ~n15397;
  assign n15400 = ~n15398 & n15399;
  assign n15401 = n14467 & ~n15400;
  assign n15402 = ~n15396 & ~n15401;
  assign n15403 = ~n15378 & ~n15384;
  assign n15404 = ~n15390 & ~n15403;
  assign n15405 = ~n15402 & n15404;
  assign n15406 = ~n15389 & ~n15405;
  assign n15407 = pi232 & ~n15406;
  assign n15408 = ~n14872 & ~n15403;
  assign n15409 = ~n15407 & ~n15408;
  assign n15410 = ~pi100 & ~n15409;
  assign n15411 = ~n14457 & ~n15373;
  assign n15412 = pi100 & n15411;
  assign n15413 = n2536 & ~n15412;
  assign n15414 = ~n13897 & n15413;
  assign n15415 = ~n15410 & n15414;
  assign n15416 = n15368 & ~n15374;
  assign n15417 = ~n15415 & n15416;
  assign n15418 = ~n14457 & ~n15371;
  assign n15419 = pi38 & ~n15418;
  assign n15420 = ~n13614 & n15369;
  assign n15421 = ~pi51 & ~n15420;
  assign n15422 = ~n5726 & n15421;
  assign n15423 = pi170 & n14271;
  assign n15424 = ~n13840 & ~n15369;
  assign n15425 = n5727 & ~n15423;
  assign n15426 = ~n15424 & n15425;
  assign n15427 = ~n8739 & ~n15426;
  assign n15428 = ~pi170 & n14917;
  assign n15429 = pi170 & n14915;
  assign n15430 = pi216 & ~n15429;
  assign n15431 = ~n15428 & n15430;
  assign n15432 = ~n15427 & ~n15431;
  assign n15433 = n15391 & ~n15422;
  assign n15434 = ~n15432 & n15433;
  assign n15435 = ~n5727 & n15421;
  assign n15436 = n14467 & ~n15435;
  assign n15437 = ~n15426 & n15436;
  assign n15438 = ~n15434 & ~n15437;
  assign n15439 = ~pi185 & n14930;
  assign n15440 = pi185 & n14933;
  assign n15441 = ~pi299 & ~n15439;
  assign n15442 = ~n15440 & n15441;
  assign n15443 = n15438 & ~n15442;
  assign n15444 = pi232 & ~n15443;
  assign n15445 = n14948 & ~n15444;
  assign n15446 = ~pi299 & ~n13763;
  assign n15447 = pi170 & ~n14954;
  assign n15448 = ~pi170 & n13763;
  assign n15449 = n10277 & ~n15448;
  assign n15450 = ~n15447 & n15449;
  assign n15451 = n14951 & ~n15450;
  assign n15452 = ~n15446 & n15451;
  assign n15453 = ~n15445 & ~n15452;
  assign n15454 = ~pi38 & ~n15453;
  assign n15455 = ~pi194 & ~n15419;
  assign n15456 = ~n15454 & n15455;
  assign n15457 = ~n14457 & ~n15382;
  assign n15458 = pi38 & ~n15457;
  assign n15459 = ~pi185 & n14937;
  assign n15460 = pi185 & n14939;
  assign n15461 = ~pi299 & ~n15459;
  assign n15462 = ~n15460 & n15461;
  assign n15463 = n15438 & ~n15462;
  assign n15464 = pi232 & ~n15463;
  assign n15465 = n14948 & ~n15464;
  assign n15466 = n10439 & n14954;
  assign n15467 = n15451 & ~n15466;
  assign n15468 = ~n15465 & ~n15467;
  assign n15469 = ~pi38 & ~n15468;
  assign n15470 = pi194 & ~n15458;
  assign n15471 = ~n15469 & n15470;
  assign n15472 = ~n15456 & ~n15471;
  assign n15473 = ~pi100 & ~n15472;
  assign n15474 = n15413 & ~n15473;
  assign n15475 = n13636 & ~n15411;
  assign n15476 = ~n15368 & ~n15475;
  assign n15477 = ~n15474 & n15476;
  assign n15478 = ~po1038 & ~n15417;
  assign n15479 = ~n15477 & n15478;
  assign n15480 = n13614 & n15368;
  assign n15481 = ~n13614 & n15380;
  assign n15482 = n15253 & ~n15481;
  assign n15483 = ~n15480 & n15482;
  assign po292 = n15479 | n15483;
  assign n15485 = pi136 & ~n14858;
  assign n15486 = ~n15254 & ~n15485;
  assign n15487 = ~n13604 & ~n15486;
  assign n15488 = ~n13665 & n15487;
  assign n15489 = pi148 & n7406;
  assign n15490 = ~n13614 & ~n15489;
  assign n15491 = ~n15488 & ~n15490;
  assign n15492 = n15253 & ~n15491;
  assign n15493 = n9401 & ~n13614;
  assign n15494 = ~pi51 & ~n15493;
  assign n15495 = n13636 & n15494;
  assign n15496 = ~n2613 & ~n15494;
  assign n15497 = ~pi184 & n14930;
  assign n15498 = ~pi141 & ~pi299;
  assign n15499 = pi184 & n14933;
  assign n15500 = ~n15497 & n15498;
  assign n15501 = ~n15499 & n15500;
  assign n15502 = ~pi287 & n12920;
  assign n15503 = pi216 & ~n15502;
  assign n15504 = n5726 & ~n15503;
  assign n15505 = n13839 & n15504;
  assign n15506 = ~pi51 & ~pi148;
  assign n15507 = ~n15505 & n15506;
  assign n15508 = ~pi51 & n14272;
  assign n15509 = n5727 & ~n15508;
  assign n15510 = pi163 & n5726;
  assign n15511 = ~n5727 & ~n15510;
  assign n15512 = ~n14457 & n15511;
  assign n15513 = ~n14915 & n15510;
  assign n15514 = pi148 & ~n15512;
  assign n15515 = ~n15513 & n15514;
  assign n15516 = ~n15509 & n15515;
  assign n15517 = pi299 & ~n15507;
  assign n15518 = ~n15516 & n15517;
  assign n15519 = ~pi184 & n14937;
  assign n15520 = pi184 & n14939;
  assign n15521 = n9398 & ~n15519;
  assign n15522 = ~n15520 & n15521;
  assign n15523 = ~n15501 & ~n15518;
  assign n15524 = ~n15522 & n15523;
  assign n15525 = pi232 & ~n15524;
  assign n15526 = n14948 & ~n15525;
  assign n15527 = ~n9400 & ~n14954;
  assign n15528 = n9400 & n13763;
  assign n15529 = pi232 & ~n15528;
  assign n15530 = ~n15527 & n15529;
  assign n15531 = n14951 & ~n15530;
  assign n15532 = n2613 & ~n15526;
  assign n15533 = ~n15531 & n15532;
  assign n15534 = n2536 & ~n15496;
  assign n15535 = ~n15533 & n15534;
  assign n15536 = n15487 & ~n15495;
  assign n15537 = ~n15535 & n15536;
  assign n15538 = ~n13614 & n15495;
  assign n15539 = ~n10821 & ~n13614;
  assign n15540 = n15494 & n15539;
  assign n15541 = ~pi51 & n14184;
  assign n15542 = ~pi148 & ~n15541;
  assign n15543 = ~n15502 & ~n15542;
  assign n15544 = ~pi148 & n13665;
  assign n15545 = ~n15543 & ~n15544;
  assign n15546 = ~n6166 & n14884;
  assign n15547 = n8739 & n14874;
  assign n15548 = pi148 & ~n15546;
  assign n15549 = ~n15547 & n15548;
  assign n15550 = ~n15545 & ~n15549;
  assign n15551 = pi299 & ~n15550;
  assign n15552 = pi184 & n13821;
  assign n15553 = n14875 & ~n15552;
  assign n15554 = n9398 & ~n15553;
  assign n15555 = pi184 & n14236;
  assign n15556 = n14879 & ~n15555;
  assign n15557 = n15498 & ~n15556;
  assign n15558 = ~n15554 & ~n15557;
  assign n15559 = ~n15551 & n15558;
  assign n15560 = pi232 & ~n15559;
  assign n15561 = ~pi100 & n14872;
  assign n15562 = ~n15560 & n15561;
  assign n15563 = ~n15540 & ~n15562;
  assign n15564 = n2536 & ~n15563;
  assign n15565 = ~n15487 & ~n15538;
  assign n15566 = ~n15564 & n15565;
  assign n15567 = ~po1038 & ~n15566;
  assign n15568 = ~n15537 & n15567;
  assign po293 = n15492 | n15568;
  assign n15570 = ~pi39 & pi137;
  assign n15571 = n2576 & n10001;
  assign n15572 = ~pi210 & n11159;
  assign n15573 = pi299 & n15572;
  assign n15574 = ~pi299 & ~po1038;
  assign n15575 = ~pi198 & n11170;
  assign n15576 = n15574 & n15575;
  assign n15577 = ~n15573 & ~n15576;
  assign n15578 = ~n15571 & ~n15577;
  assign n15579 = po1038 & n15572;
  assign n15580 = ~n15578 & ~n15579;
  assign n15581 = n8738 & ~n15580;
  assign po294 = n15570 | n15581;
  assign n15583 = ~n9401 & n11070;
  assign n15584 = ~pi39 & ~n15583;
  assign n15585 = ~n6205 & n9399;
  assign n15586 = n6205 & n6341;
  assign n15587 = n8752 & n15586;
  assign n15588 = n9398 & ~n15587;
  assign n15589 = ~n15585 & ~n15588;
  assign n15590 = pi232 & ~n15589;
  assign n15591 = pi141 & n10439;
  assign n15592 = ~n11067 & ~n15591;
  assign n15593 = ~n15590 & ~n15592;
  assign n15594 = pi39 & ~n15593;
  assign n15595 = n9833 & ~n15584;
  assign n15596 = ~n15594 & n15595;
  assign n15597 = ~pi138 & n15596;
  assign n15598 = n8939 & ~n8970;
  assign n15599 = pi92 & ~n15598;
  assign n15600 = n2533 & ~n15599;
  assign n15601 = ~pi75 & ~n8976;
  assign n15602 = ~pi299 & ~n8991;
  assign n15603 = ~n9008 & ~n11458;
  assign n15604 = n9018 & ~n15603;
  assign n15605 = n15602 & ~n15604;
  assign n15606 = ~n6221 & ~n9008;
  assign n15607 = n8739 & ~n15603;
  assign n15608 = ~n15606 & n15607;
  assign n15609 = n8979 & ~n15608;
  assign n15610 = ~n15605 & ~n15609;
  assign n15611 = ~pi232 & ~n15610;
  assign n15612 = ~n8988 & ~n15603;
  assign n15613 = ~n8978 & ~n15612;
  assign n15614 = pi148 & ~n15613;
  assign n15615 = ~n9399 & ~n15609;
  assign n15616 = ~n15614 & ~n15615;
  assign n15617 = pi141 & n8993;
  assign n15618 = n15604 & ~n15617;
  assign n15619 = n15602 & ~n15618;
  assign n15620 = ~n15616 & ~n15619;
  assign n15621 = pi232 & ~n15620;
  assign n15622 = ~n15611 & ~n15621;
  assign n15623 = pi39 & ~n15622;
  assign n15624 = pi299 & ~n9219;
  assign n15625 = ~pi299 & ~n9634;
  assign n15626 = ~pi232 & ~n15624;
  assign n15627 = ~n15625 & n15626;
  assign n15628 = ~pi39 & ~n15627;
  assign n15629 = ~pi141 & n15625;
  assign n15630 = ~n6166 & ~n9634;
  assign n15631 = ~n13026 & ~n15630;
  assign n15632 = n9398 & ~n15631;
  assign n15633 = pi148 & n6166;
  assign n15634 = ~n9219 & ~n15633;
  assign n15635 = pi148 & n13005;
  assign n15636 = ~n15634 & ~n15635;
  assign n15637 = pi299 & ~n15636;
  assign n15638 = pi232 & ~n15629;
  assign n15639 = ~n15632 & n15638;
  assign n15640 = ~n15637 & n15639;
  assign n15641 = n15628 & ~n15640;
  assign n15642 = n2613 & ~n15623;
  assign n15643 = ~n15641 & n15642;
  assign n15644 = ~pi87 & ~n15643;
  assign n15645 = n15601 & ~n15644;
  assign n15646 = ~pi92 & ~n15645;
  assign n15647 = n15600 & ~n15646;
  assign n15648 = ~pi55 & ~n15647;
  assign n15649 = n8940 & ~n12939;
  assign n15650 = pi55 & ~n15649;
  assign n15651 = ~n15648 & ~n15650;
  assign n15652 = n2530 & ~n15651;
  assign n15653 = n9532 & ~n15652;
  assign n15654 = pi138 & n15653;
  assign n15655 = ~pi118 & n12919;
  assign n15656 = ~pi139 & n15655;
  assign n15657 = ~n15597 & ~n15656;
  assign n15658 = ~n15654 & n15657;
  assign n15659 = ~pi138 & ~n8679;
  assign n15660 = n15596 & ~n15659;
  assign n15661 = n15653 & n15659;
  assign n15662 = n15656 & ~n15660;
  assign n15663 = ~n15661 & n15662;
  assign po295 = ~n15658 & ~n15663;
  assign n15665 = n11070 & ~n14862;
  assign n15666 = ~pi39 & ~n15665;
  assign n15667 = ~pi232 & ~n11067;
  assign n15668 = ~n11063 & n14878;
  assign n15669 = ~n6205 & n8723;
  assign n15670 = n8722 & ~n15587;
  assign n15671 = ~n11066 & ~n15669;
  assign n15672 = ~n15668 & ~n15670;
  assign n15673 = n15671 & n15672;
  assign n15674 = pi232 & ~n15673;
  assign n15675 = ~n15667 & ~n15674;
  assign n15676 = pi39 & ~n15675;
  assign n15677 = n9833 & ~n15666;
  assign n15678 = ~n15676 & n15677;
  assign n15679 = ~pi139 & n15678;
  assign n15680 = ~pi191 & n15625;
  assign n15681 = n8722 & ~n15631;
  assign n15682 = ~n9219 & ~n14883;
  assign n15683 = pi169 & n13005;
  assign n15684 = ~n15682 & ~n15683;
  assign n15685 = pi299 & ~n15684;
  assign n15686 = pi232 & ~n15680;
  assign n15687 = ~n15681 & n15686;
  assign n15688 = ~n15685 & n15687;
  assign n15689 = n15628 & ~n15688;
  assign n15690 = ~pi191 & n15605;
  assign n15691 = ~pi169 & n9008;
  assign n15692 = ~n15612 & ~n15691;
  assign n15693 = n8739 & ~n15692;
  assign n15694 = n8979 & ~n15693;
  assign n15695 = ~n8993 & n15604;
  assign n15696 = n15602 & ~n15695;
  assign n15697 = pi191 & n15696;
  assign n15698 = ~n15694 & ~n15697;
  assign n15699 = pi232 & ~n15698;
  assign n15700 = ~n15611 & ~n15690;
  assign n15701 = ~n15699 & n15700;
  assign n15702 = pi39 & ~n15701;
  assign n15703 = n2613 & ~n15702;
  assign n15704 = ~n15689 & n15703;
  assign n15705 = ~pi87 & ~n15704;
  assign n15706 = n15601 & ~n15705;
  assign n15707 = ~pi92 & ~n15706;
  assign n15708 = n15600 & ~n15707;
  assign n15709 = ~pi55 & ~n15708;
  assign n15710 = ~n15650 & ~n15709;
  assign n15711 = n2530 & ~n15710;
  assign n15712 = n9532 & ~n15711;
  assign n15713 = pi139 & n15712;
  assign n15714 = ~n15655 & ~n15679;
  assign n15715 = ~n15713 & n15714;
  assign n15716 = ~pi139 & ~n8680;
  assign n15717 = n15678 & ~n15716;
  assign n15718 = n15712 & n15716;
  assign n15719 = n15655 & ~n15717;
  assign n15720 = ~n15718 & n15719;
  assign po296 = ~n15715 & ~n15720;
  assign n15722 = ~pi140 & ~n2923;
  assign n15723 = ~pi647 & n15722;
  assign n15724 = pi665 & pi1091;
  assign n15725 = pi680 & ~n15724;
  assign n15726 = n2923 & n15725;
  assign n15727 = ~pi738 & n15726;
  assign n15728 = ~n15722 & ~n15727;
  assign n15729 = ~pi778 & n15728;
  assign n15730 = ~pi625 & n15727;
  assign n15731 = ~n15728 & ~n15730;
  assign n15732 = pi1153 & ~n15731;
  assign n15733 = ~pi1153 & ~n15722;
  assign n15734 = ~n15730 & n15733;
  assign n15735 = ~n15732 & ~n15734;
  assign n15736 = pi778 & ~n15735;
  assign n15737 = ~n15729 & ~n15736;
  assign n15738 = pi660 & ~pi1155;
  assign n15739 = ~pi660 & pi1155;
  assign n15740 = ~n15738 & ~n15739;
  assign n15741 = pi785 & ~n15740;
  assign n15742 = n2923 & n15741;
  assign n15743 = n15737 & ~n15742;
  assign n15744 = pi627 & ~pi1154;
  assign n15745 = ~pi627 & pi1154;
  assign n15746 = ~n15744 & ~n15745;
  assign n15747 = pi781 & ~n15746;
  assign n15748 = n2923 & n15747;
  assign n15749 = n15743 & ~n15748;
  assign n15750 = ~pi648 & pi1159;
  assign n15751 = pi648 & ~pi1159;
  assign n15752 = ~n15750 & ~n15751;
  assign n15753 = pi789 & ~n15752;
  assign n15754 = n2923 & n15753;
  assign n15755 = n15749 & ~n15754;
  assign n15756 = ~pi641 & pi1158;
  assign n15757 = pi641 & ~pi1158;
  assign n15758 = ~n15756 & ~n15757;
  assign n15759 = pi788 & ~n15758;
  assign n15760 = n2923 & n15759;
  assign n15761 = n15755 & ~n15760;
  assign n15762 = ~pi628 & pi1156;
  assign n15763 = pi628 & ~pi1156;
  assign n15764 = ~n15762 & ~n15763;
  assign n15765 = pi792 & ~n15764;
  assign n15766 = n2923 & n15765;
  assign n15767 = n15761 & ~n15766;
  assign n15768 = pi647 & n15767;
  assign n15769 = pi1157 & ~n15723;
  assign n15770 = ~n15768 & n15769;
  assign n15771 = ~pi628 & n2923;
  assign n15772 = pi1156 & ~n15771;
  assign n15773 = n15761 & n15772;
  assign n15774 = pi608 & ~pi1153;
  assign n15775 = ~pi608 & pi1153;
  assign n15776 = ~n15774 & ~n15775;
  assign n15777 = pi778 & ~n15776;
  assign n15778 = n2923 & n15777;
  assign n15779 = pi621 & pi1091;
  assign n15780 = pi603 & ~n15779;
  assign n15781 = n2923 & n15780;
  assign n15782 = ~pi761 & n15781;
  assign n15783 = ~n15722 & ~n15782;
  assign n15784 = ~n15778 & ~n15783;
  assign n15785 = ~pi785 & ~n15784;
  assign n15786 = pi609 & ~n15777;
  assign n15787 = n2923 & ~n15786;
  assign n15788 = ~n15783 & ~n15787;
  assign n15789 = pi1155 & ~n15788;
  assign n15790 = pi609 & n2923;
  assign n15791 = n15784 & ~n15790;
  assign n15792 = ~pi1155 & ~n15791;
  assign n15793 = ~n15789 & ~n15792;
  assign n15794 = pi785 & ~n15793;
  assign n15795 = ~n15785 & ~n15794;
  assign n15796 = ~pi781 & ~n15795;
  assign n15797 = ~pi618 & n2923;
  assign n15798 = n15795 & ~n15797;
  assign n15799 = pi1154 & ~n15798;
  assign n15800 = pi618 & n2923;
  assign n15801 = n15795 & ~n15800;
  assign n15802 = ~pi1154 & ~n15801;
  assign n15803 = ~n15799 & ~n15802;
  assign n15804 = pi781 & ~n15803;
  assign n15805 = ~n15796 & ~n15804;
  assign n15806 = ~pi789 & ~n15805;
  assign n15807 = ~pi619 & n15722;
  assign n15808 = pi619 & n15805;
  assign n15809 = pi1159 & ~n15807;
  assign n15810 = ~n15808 & n15809;
  assign n15811 = ~pi619 & n15805;
  assign n15812 = pi619 & n15722;
  assign n15813 = ~pi1159 & ~n15812;
  assign n15814 = ~n15811 & n15813;
  assign n15815 = ~n15810 & ~n15814;
  assign n15816 = pi789 & ~n15815;
  assign n15817 = ~n15806 & ~n15816;
  assign n15818 = ~pi626 & pi1158;
  assign n15819 = pi626 & ~pi1158;
  assign n15820 = ~n15818 & ~n15819;
  assign n15821 = n15817 & n15820;
  assign n15822 = n15722 & ~n15820;
  assign n15823 = ~n15821 & ~n15822;
  assign n15824 = ~n15758 & ~n15823;
  assign n15825 = ~pi626 & pi641;
  assign n15826 = pi626 & ~pi641;
  assign n15827 = ~n15825 & ~n15826;
  assign n15828 = ~n15820 & ~n15827;
  assign n15829 = n15755 & n15828;
  assign n15830 = ~n15824 & ~n15829;
  assign n15831 = pi788 & ~n15830;
  assign n15832 = pi788 & ~n15820;
  assign n15833 = ~n15759 & ~n15832;
  assign n15834 = pi618 & n15743;
  assign n15835 = pi609 & n15737;
  assign n15836 = ~n15728 & ~n15780;
  assign n15837 = pi625 & n15836;
  assign n15838 = n15783 & ~n15836;
  assign n15839 = ~n15837 & ~n15838;
  assign n15840 = n15733 & ~n15839;
  assign n15841 = ~pi608 & ~n15732;
  assign n15842 = ~n15840 & n15841;
  assign n15843 = pi1153 & n15783;
  assign n15844 = ~n15837 & n15843;
  assign n15845 = pi608 & ~n15734;
  assign n15846 = ~n15844 & n15845;
  assign n15847 = ~n15842 & ~n15846;
  assign n15848 = pi778 & ~n15847;
  assign n15849 = ~pi778 & ~n15838;
  assign n15850 = ~n15848 & ~n15849;
  assign n15851 = ~pi609 & ~n15850;
  assign n15852 = ~pi1155 & ~n15835;
  assign n15853 = ~n15851 & n15852;
  assign n15854 = ~pi660 & ~n15789;
  assign n15855 = ~n15853 & n15854;
  assign n15856 = ~pi609 & n15737;
  assign n15857 = pi609 & ~n15850;
  assign n15858 = pi1155 & ~n15856;
  assign n15859 = ~n15857 & n15858;
  assign n15860 = pi660 & ~n15792;
  assign n15861 = ~n15859 & n15860;
  assign n15862 = ~n15855 & ~n15861;
  assign n15863 = pi785 & ~n15862;
  assign n15864 = ~pi785 & ~n15850;
  assign n15865 = ~n15863 & ~n15864;
  assign n15866 = ~pi618 & ~n15865;
  assign n15867 = ~pi1154 & ~n15834;
  assign n15868 = ~n15866 & n15867;
  assign n15869 = ~pi627 & ~n15799;
  assign n15870 = ~n15868 & n15869;
  assign n15871 = ~pi618 & n15743;
  assign n15872 = pi618 & ~n15865;
  assign n15873 = pi1154 & ~n15871;
  assign n15874 = ~n15872 & n15873;
  assign n15875 = pi627 & ~n15802;
  assign n15876 = ~n15874 & n15875;
  assign n15877 = ~n15870 & ~n15876;
  assign n15878 = pi781 & ~n15877;
  assign n15879 = ~pi781 & ~n15865;
  assign n15880 = ~n15878 & ~n15879;
  assign n15881 = ~pi789 & n15880;
  assign n15882 = ~pi619 & n15749;
  assign n15883 = pi619 & ~n15880;
  assign n15884 = pi1159 & ~n15882;
  assign n15885 = ~n15883 & n15884;
  assign n15886 = pi648 & ~n15814;
  assign n15887 = ~n15885 & n15886;
  assign n15888 = pi619 & n15749;
  assign n15889 = ~pi619 & ~n15880;
  assign n15890 = ~pi1159 & ~n15888;
  assign n15891 = ~n15889 & n15890;
  assign n15892 = ~pi648 & ~n15810;
  assign n15893 = ~n15891 & n15892;
  assign n15894 = pi789 & ~n15887;
  assign n15895 = ~n15893 & n15894;
  assign n15896 = n15833 & ~n15881;
  assign n15897 = ~n15895 & n15896;
  assign n15898 = ~n15831 & ~n15897;
  assign n15899 = ~pi628 & n15898;
  assign n15900 = pi788 & ~n15823;
  assign n15901 = ~pi788 & n15817;
  assign n15902 = ~n15900 & ~n15901;
  assign n15903 = pi628 & n15902;
  assign n15904 = ~pi1156 & ~n15903;
  assign n15905 = ~n15899 & n15904;
  assign n15906 = ~pi629 & ~n15773;
  assign n15907 = ~n15905 & n15906;
  assign n15908 = pi628 & n2923;
  assign n15909 = ~pi1156 & ~n15908;
  assign n15910 = n15761 & n15909;
  assign n15911 = ~pi628 & n15902;
  assign n15912 = pi628 & n15898;
  assign n15913 = pi1156 & ~n15911;
  assign n15914 = ~n15912 & n15913;
  assign n15915 = pi629 & ~n15910;
  assign n15916 = ~n15914 & n15915;
  assign n15917 = ~n15907 & ~n15916;
  assign n15918 = pi792 & ~n15917;
  assign n15919 = ~pi792 & n15898;
  assign n15920 = ~n15918 & ~n15919;
  assign n15921 = ~pi647 & n15920;
  assign n15922 = ~pi629 & pi1156;
  assign n15923 = pi629 & ~pi1156;
  assign n15924 = ~n15922 & ~n15923;
  assign n15925 = pi792 & ~n15924;
  assign n15926 = n15902 & ~n15925;
  assign n15927 = ~n15722 & n15925;
  assign n15928 = ~n15926 & ~n15927;
  assign n15929 = pi647 & n15928;
  assign n15930 = ~pi1157 & ~n15929;
  assign n15931 = ~n15921 & n15930;
  assign n15932 = ~pi630 & ~n15770;
  assign n15933 = ~n15931 & n15932;
  assign n15934 = ~pi647 & n15767;
  assign n15935 = pi647 & n15722;
  assign n15936 = ~pi1157 & ~n15935;
  assign n15937 = ~n15934 & n15936;
  assign n15938 = ~pi647 & n15928;
  assign n15939 = pi647 & n15920;
  assign n15940 = pi1157 & ~n15938;
  assign n15941 = ~n15939 & n15940;
  assign n15942 = pi630 & ~n15937;
  assign n15943 = ~n15941 & n15942;
  assign n15944 = ~n15933 & ~n15943;
  assign n15945 = pi787 & ~n15944;
  assign n15946 = ~pi787 & n15920;
  assign n15947 = ~n15945 & ~n15946;
  assign n15948 = ~pi790 & ~n15947;
  assign n15949 = ~pi787 & ~n15767;
  assign n15950 = ~n15770 & ~n15937;
  assign n15951 = pi787 & ~n15950;
  assign n15952 = ~n15949 & ~n15951;
  assign n15953 = ~pi644 & n15952;
  assign n15954 = pi644 & ~n15947;
  assign n15955 = pi715 & ~n15953;
  assign n15956 = ~n15954 & n15955;
  assign n15957 = ~pi630 & pi1157;
  assign n15958 = pi630 & ~pi1157;
  assign n15959 = ~n15957 & ~n15958;
  assign n15960 = pi787 & ~n15959;
  assign n15961 = n15928 & ~n15960;
  assign n15962 = n15722 & n15960;
  assign n15963 = ~n15961 & ~n15962;
  assign n15964 = pi644 & ~n15963;
  assign n15965 = ~pi644 & n15722;
  assign n15966 = ~pi715 & ~n15965;
  assign n15967 = ~n15964 & n15966;
  assign n15968 = pi1160 & ~n15967;
  assign n15969 = ~n15956 & n15968;
  assign n15970 = ~pi644 & ~n15963;
  assign n15971 = pi644 & n15722;
  assign n15972 = pi715 & ~n15971;
  assign n15973 = ~n15970 & n15972;
  assign n15974 = pi644 & n15952;
  assign n15975 = ~pi644 & ~n15947;
  assign n15976 = ~pi715 & ~n15974;
  assign n15977 = ~n15975 & n15976;
  assign n15978 = ~pi1160 & ~n15973;
  assign n15979 = ~n15977 & n15978;
  assign n15980 = ~n15969 & ~n15979;
  assign n15981 = pi790 & ~n15980;
  assign n15982 = pi832 & ~n15948;
  assign n15983 = ~n15981 & n15982;
  assign n15984 = ~pi140 & po1038;
  assign n15985 = ~pi102 & ~n10886;
  assign n15986 = ~pi98 & ~n2785;
  assign n15987 = ~n15985 & n15986;
  assign n15988 = n7369 & n11857;
  assign n15989 = n15987 & n15988;
  assign n15990 = n8611 & n8623;
  assign n15991 = n15989 & n15990;
  assign n15992 = ~pi40 & ~n15991;
  assign n15993 = n9914 & ~n15992;
  assign n15994 = ~pi252 & ~n15993;
  assign n15995 = n2709 & n6130;
  assign n15996 = n2500 & n15989;
  assign n15997 = ~pi47 & ~n15996;
  assign n15998 = pi314 & n9894;
  assign n15999 = n15997 & ~n15998;
  assign n16000 = n15995 & ~n15999;
  assign n16001 = ~pi35 & ~n16000;
  assign n16002 = ~pi40 & n9870;
  assign n16003 = ~n16001 & n16002;
  assign n16004 = pi252 & ~n2742;
  assign n16005 = ~n16003 & n16004;
  assign n16006 = ~n15994 & ~n16005;
  assign n16007 = n2518 & n16006;
  assign n16008 = pi1092 & n16007;
  assign n16009 = ~n11855 & n16008;
  assign n16010 = ~pi88 & ~n15987;
  assign n16011 = n10620 & ~n16010;
  assign n16012 = ~pi252 & n10959;
  assign n16013 = n16011 & n16012;
  assign n16014 = n2501 & n16011;
  assign n16015 = ~pi47 & ~n16014;
  assign n16016 = ~n15998 & n16015;
  assign n16017 = n15995 & ~n16016;
  assign n16018 = ~pi35 & ~n16017;
  assign n16019 = pi252 & n9870;
  assign n16020 = ~n16018 & n16019;
  assign n16021 = ~pi40 & ~n16013;
  assign n16022 = ~n16020 & n16021;
  assign n16023 = n7348 & n9914;
  assign n16024 = ~n16022 & n16023;
  assign n16025 = ~n16009 & ~n16024;
  assign n16026 = pi1093 & ~n16025;
  assign n16027 = ~n2921 & ~n16026;
  assign n16028 = n6179 & n16008;
  assign n16029 = ~n2922 & ~n16028;
  assign n16030 = ~n16027 & ~n16029;
  assign n16031 = ~pi1091 & n16026;
  assign n16032 = ~n16030 & ~n16031;
  assign n16033 = ~pi210 & n16032;
  assign n16034 = ~n2518 & ~n6439;
  assign n16035 = ~n3387 & ~n16022;
  assign n16036 = ~pi32 & ~n16035;
  assign n16037 = n7348 & ~n16034;
  assign n16038 = ~n16036 & n16037;
  assign n16039 = ~n16009 & ~n16038;
  assign n16040 = n7561 & ~n16039;
  assign n16041 = ~pi32 & ~n16006;
  assign n16042 = pi829 & n10631;
  assign n16043 = ~n16034 & n16042;
  assign n16044 = ~n16041 & n16043;
  assign n16045 = n16039 & ~n16044;
  assign n16046 = pi1093 & ~n16045;
  assign n16047 = ~n2921 & ~n16046;
  assign n16048 = ~n16029 & ~n16047;
  assign n16049 = ~n16040 & ~n16048;
  assign n16050 = pi210 & n16049;
  assign n16051 = ~n16033 & ~n16050;
  assign n16052 = pi299 & ~n16051;
  assign n16053 = ~pi198 & n16032;
  assign n16054 = pi198 & n16049;
  assign n16055 = ~n16053 & ~n16054;
  assign n16056 = ~pi299 & ~n16055;
  assign n16057 = ~n16052 & ~n16056;
  assign n16058 = ~pi39 & ~n16057;
  assign n16059 = ~n6170 & n6333;
  assign n16060 = ~pi120 & ~n16059;
  assign n16061 = pi120 & ~n2523;
  assign n16062 = ~n16060 & ~n16061;
  assign n16063 = n2923 & n16062;
  assign n16064 = ~n6166 & n16063;
  assign n16065 = n2523 & n2923;
  assign n16066 = n6173 & n13416;
  assign n16067 = n16065 & ~n16066;
  assign n16068 = pi120 & ~n16067;
  assign n16069 = n2923 & n16059;
  assign n16070 = ~pi120 & ~n16069;
  assign n16071 = pi1091 & ~n16068;
  assign n16072 = ~n16070 & n16071;
  assign n16073 = pi120 & ~n16065;
  assign n16074 = ~pi1091 & ~n16073;
  assign n16075 = pi120 & pi824;
  assign n16076 = n6173 & n16075;
  assign n16077 = n16074 & ~n16076;
  assign n16078 = ~n16070 & n16077;
  assign n16079 = ~n16072 & ~n16078;
  assign n16080 = n6166 & ~n16079;
  assign n16081 = ~n16064 & ~n16080;
  assign n16082 = ~n6159 & ~n16063;
  assign n16083 = ~n6166 & n16079;
  assign n16084 = n6166 & ~n16063;
  assign n16085 = ~n16083 & ~n16084;
  assign n16086 = n6159 & ~n16085;
  assign n16087 = ~n16082 & ~n16086;
  assign n16088 = n6160 & ~n16087;
  assign n16089 = ~n16081 & ~n16088;
  assign n16090 = pi681 & ~n16089;
  assign n16091 = pi661 & n16089;
  assign n16092 = pi616 & ~n16063;
  assign n16093 = pi614 & ~n16063;
  assign n16094 = ~n16092 & ~n16093;
  assign n16095 = ~n16088 & n16094;
  assign n16096 = ~n6163 & ~n16095;
  assign n16097 = n6163 & n16079;
  assign n16098 = ~n6166 & ~n16097;
  assign n16099 = ~n16096 & n16098;
  assign n16100 = ~n16080 & ~n16099;
  assign n16101 = ~pi661 & ~n16100;
  assign n16102 = ~pi681 & ~n16091;
  assign n16103 = ~n16101 & n16102;
  assign n16104 = ~n16090 & ~n16103;
  assign n16105 = ~n6194 & n16104;
  assign n16106 = pi681 & ~n16095;
  assign n16107 = pi680 & ~n16085;
  assign n16108 = ~pi662 & n6162;
  assign n16109 = ~pi680 & ~n16063;
  assign n16110 = pi616 & n16108;
  assign n16111 = ~n16109 & n16110;
  assign n16112 = ~n16107 & n16111;
  assign n16113 = pi616 & n16063;
  assign n16114 = ~n16108 & n16113;
  assign n16115 = ~n16112 & ~n16114;
  assign n16116 = n6164 & ~n16085;
  assign n16117 = ~n6164 & ~n16095;
  assign n16118 = ~pi616 & ~n16116;
  assign n16119 = ~n16117 & n16118;
  assign n16120 = ~pi681 & n16115;
  assign n16121 = ~n16119 & n16120;
  assign n16122 = ~n16106 & ~n16121;
  assign n16123 = n6194 & n16122;
  assign n16124 = ~n16105 & ~n16123;
  assign n16125 = pi223 & n16124;
  assign n16126 = n2608 & ~n16063;
  assign n16127 = ~pi824 & ~n16059;
  assign n16128 = n6333 & ~n9836;
  assign n16129 = pi1092 & n16128;
  assign n16130 = ~n10631 & ~n16129;
  assign n16131 = ~n16127 & ~n16130;
  assign n16132 = pi1093 & n16131;
  assign n16133 = ~pi120 & ~n16132;
  assign n16134 = n16074 & ~n16133;
  assign n16135 = n2921 & n16069;
  assign n16136 = pi829 & ~n16129;
  assign n16137 = ~pi829 & ~n16131;
  assign n16138 = n7453 & ~n16136;
  assign n16139 = ~n16137 & n16138;
  assign n16140 = ~n16135 & ~n16139;
  assign n16141 = pi1091 & ~n16140;
  assign n16142 = ~pi120 & ~n16141;
  assign n16143 = ~n16073 & ~n16142;
  assign n16144 = ~n16134 & ~n16143;
  assign n16145 = n6166 & ~n16144;
  assign n16146 = ~n16064 & ~n16145;
  assign n16147 = ~n6161 & ~n16146;
  assign n16148 = n6161 & ~n16144;
  assign n16149 = ~n16147 & ~n16148;
  assign n16150 = ~n6164 & n16149;
  assign n16151 = pi680 & n16144;
  assign n16152 = n16108 & n16151;
  assign n16153 = ~n16150 & ~n16152;
  assign n16154 = ~n6194 & n16153;
  assign n16155 = ~pi603 & ~n16063;
  assign n16156 = ~n6166 & n16144;
  assign n16157 = ~n16084 & ~n16156;
  assign n16158 = pi603 & ~n16157;
  assign n16159 = ~n16155 & ~n16158;
  assign n16160 = ~pi642 & ~n16159;
  assign n16161 = ~n16082 & ~n16160;
  assign n16162 = ~pi614 & ~n16161;
  assign n16163 = ~n16093 & ~n16162;
  assign n16164 = ~pi616 & ~n16163;
  assign n16165 = ~n16092 & ~n16164;
  assign n16166 = pi681 & ~n16165;
  assign n16167 = pi614 & n16063;
  assign n16168 = ~n16108 & n16167;
  assign n16169 = pi680 & ~n16157;
  assign n16170 = pi614 & n16108;
  assign n16171 = ~n16109 & n16170;
  assign n16172 = ~n16169 & n16171;
  assign n16173 = ~pi614 & ~n6164;
  assign n16174 = ~pi616 & ~n16161;
  assign n16175 = ~n16092 & n16173;
  assign n16176 = ~n16174 & n16175;
  assign n16177 = ~pi614 & pi680;
  assign n16178 = n16108 & n16177;
  assign n16179 = n16157 & n16178;
  assign n16180 = ~n16176 & ~n16179;
  assign n16181 = ~n16172 & n16180;
  assign n16182 = ~pi681 & ~n16168;
  assign n16183 = n16181 & n16182;
  assign n16184 = ~n16166 & ~n16183;
  assign n16185 = n6194 & n16184;
  assign n16186 = ~n16154 & ~n16185;
  assign n16187 = ~n2608 & n16186;
  assign n16188 = ~n16126 & ~n16187;
  assign n16189 = ~pi223 & ~n16188;
  assign n16190 = ~n16125 & ~n16189;
  assign n16191 = ~pi299 & ~n16190;
  assign n16192 = ~n6220 & n16153;
  assign n16193 = ~n3302 & n16192;
  assign n16194 = ~n6221 & n16153;
  assign n16195 = n6221 & n16184;
  assign n16196 = ~n16194 & ~n16195;
  assign n16197 = n6220 & ~n16196;
  assign n16198 = ~n3302 & n16197;
  assign n16199 = n3302 & n16063;
  assign n16200 = ~pi215 & ~n16199;
  assign n16201 = ~n16193 & n16200;
  assign n16202 = ~n16198 & n16201;
  assign n16203 = ~n6220 & n16104;
  assign n16204 = n6219 & ~n16122;
  assign n16205 = ~n6219 & ~n16104;
  assign n16206 = n6220 & ~n16204;
  assign n16207 = ~n16205 & n16206;
  assign n16208 = ~n16203 & ~n16207;
  assign n16209 = pi215 & n16208;
  assign n16210 = ~n16202 & ~n16209;
  assign n16211 = pi299 & ~n16210;
  assign n16212 = ~n16191 & ~n16211;
  assign n16213 = pi39 & ~n16212;
  assign n16214 = ~n16058 & ~n16213;
  assign n16215 = ~pi38 & ~n16214;
  assign n16216 = n2923 & n6116;
  assign n16217 = pi38 & ~n16216;
  assign n16218 = ~n16215 & ~n16217;
  assign n16219 = n9829 & n16218;
  assign n16220 = ~pi140 & ~n16219;
  assign n16221 = n15759 & ~n16220;
  assign n16222 = n15747 & ~n16220;
  assign n16223 = pi140 & ~n9829;
  assign n16224 = ~pi140 & pi738;
  assign n16225 = ~n16218 & n16224;
  assign n16226 = n6081 & n15726;
  assign n16227 = pi38 & ~n16226;
  assign n16228 = ~pi39 & n16065;
  assign n16229 = ~pi140 & ~n16228;
  assign n16230 = n16227 & ~n16229;
  assign n16231 = n2608 & n16062;
  assign n16232 = n2923 & ~n15725;
  assign n16233 = n16231 & n16232;
  assign n16234 = ~n15725 & n16153;
  assign n16235 = ~n6194 & ~n16234;
  assign n16236 = ~pi680 & ~n16165;
  assign n16237 = n15724 & n16063;
  assign n16238 = n6166 & ~n16237;
  assign n16239 = n15724 & n16143;
  assign n16240 = ~n6166 & ~n16239;
  assign n16241 = ~n16238 & ~n16240;
  assign n16242 = n6161 & n16241;
  assign n16243 = ~n6161 & n16237;
  assign n16244 = pi680 & ~n16243;
  assign n16245 = ~n16242 & n16244;
  assign n16246 = ~n16236 & ~n16245;
  assign n16247 = ~n16108 & n16246;
  assign n16248 = pi680 & ~n16241;
  assign n16249 = n16108 & ~n16248;
  assign n16250 = ~n16236 & n16249;
  assign n16251 = ~n16247 & ~n16250;
  assign n16252 = n6194 & n16251;
  assign n16253 = ~n2608 & ~n16235;
  assign n16254 = ~n16252 & n16253;
  assign n16255 = ~pi223 & ~n16233;
  assign n16256 = ~n16254 & n16255;
  assign n16257 = ~pi680 & ~n16095;
  assign n16258 = pi665 & n16072;
  assign n16259 = ~n6166 & ~n16258;
  assign n16260 = ~n16238 & ~n16259;
  assign n16261 = n6164 & ~n16260;
  assign n16262 = n16244 & ~n16260;
  assign n16263 = ~n16261 & ~n16262;
  assign n16264 = ~n16257 & n16263;
  assign n16265 = n6194 & n16264;
  assign n16266 = ~pi680 & ~n16089;
  assign n16267 = pi680 & ~n16258;
  assign n16268 = n15724 & n16064;
  assign n16269 = ~n6161 & n16268;
  assign n16270 = n16267 & ~n16269;
  assign n16271 = ~n16266 & ~n16270;
  assign n16272 = n16263 & n16271;
  assign n16273 = ~n6194 & n16272;
  assign n16274 = pi223 & ~n16265;
  assign n16275 = ~n16273 & n16274;
  assign n16276 = ~n16256 & ~n16275;
  assign n16277 = ~pi299 & ~n16276;
  assign n16278 = ~n15725 & n16199;
  assign n16279 = ~n6221 & ~n16234;
  assign n16280 = n6221 & n16251;
  assign n16281 = ~n3302 & ~n16279;
  assign n16282 = ~n16280 & n16281;
  assign n16283 = ~pi215 & ~n16278;
  assign n16284 = ~n16282 & n16283;
  assign n16285 = n6221 & n16264;
  assign n16286 = ~n6221 & n16272;
  assign n16287 = pi215 & ~n16285;
  assign n16288 = ~n16286 & n16287;
  assign n16289 = ~n16284 & ~n16288;
  assign n16290 = pi299 & ~n16289;
  assign n16291 = ~n16277 & ~n16290;
  assign n16292 = ~pi140 & n16291;
  assign n16293 = ~n6221 & n16081;
  assign n16294 = ~n15724 & n16063;
  assign n16295 = ~n16083 & n16294;
  assign n16296 = n16108 & ~n16295;
  assign n16297 = n6161 & n16083;
  assign n16298 = n15725 & n16063;
  assign n16299 = ~n16297 & n16298;
  assign n16300 = ~n16296 & n16299;
  assign n16301 = ~n16293 & n16300;
  assign n16302 = pi215 & ~n16301;
  assign n16303 = n15725 & n16153;
  assign n16304 = ~n6221 & ~n16303;
  assign n16305 = ~n6161 & n16294;
  assign n16306 = ~n15724 & n16157;
  assign n16307 = n6161 & n16306;
  assign n16308 = ~n16305 & ~n16307;
  assign n16309 = ~n16108 & n16308;
  assign n16310 = n16108 & ~n16306;
  assign n16311 = pi680 & ~n16310;
  assign n16312 = ~n16309 & n16311;
  assign n16313 = n6221 & ~n16312;
  assign n16314 = ~n3302 & ~n16304;
  assign n16315 = ~n16313 & n16314;
  assign n16316 = n3302 & n16062;
  assign n16317 = n15726 & n16316;
  assign n16318 = ~pi215 & ~n16317;
  assign n16319 = ~n16315 & n16318;
  assign n16320 = ~n16302 & ~n16319;
  assign n16321 = pi299 & ~n16320;
  assign n16322 = n15726 & n16231;
  assign n16323 = ~n6194 & ~n16303;
  assign n16324 = n6194 & ~n16312;
  assign n16325 = ~n2608 & ~n16323;
  assign n16326 = ~n16324 & n16325;
  assign n16327 = ~n16322 & ~n16326;
  assign n16328 = ~pi223 & ~n16327;
  assign n16329 = ~n6194 & n16081;
  assign n16330 = n16299 & ~n16329;
  assign n16331 = pi223 & ~n16296;
  assign n16332 = n16330 & n16331;
  assign n16333 = ~n16328 & ~n16332;
  assign n16334 = ~pi299 & n16333;
  assign n16335 = ~n16321 & ~n16334;
  assign n16336 = pi140 & ~n16335;
  assign n16337 = pi39 & ~n16336;
  assign n16338 = ~n16292 & n16337;
  assign n16339 = pi665 & ~n16031;
  assign n16340 = ~n16032 & ~n16339;
  assign n16341 = ~pi198 & ~n16340;
  assign n16342 = pi665 & ~n16040;
  assign n16343 = ~n16049 & ~n16342;
  assign n16344 = pi198 & ~n16343;
  assign n16345 = ~n16341 & ~n16344;
  assign n16346 = pi680 & n16345;
  assign n16347 = ~pi299 & ~n16346;
  assign n16348 = pi210 & ~n16343;
  assign n16349 = ~pi210 & ~n16340;
  assign n16350 = ~n16348 & ~n16349;
  assign n16351 = pi680 & n16350;
  assign n16352 = pi299 & ~n16351;
  assign n16353 = ~n16347 & ~n16352;
  assign n16354 = pi140 & ~n16353;
  assign n16355 = pi665 & n16048;
  assign n16356 = pi198 & ~n16355;
  assign n16357 = pi665 & n16030;
  assign n16358 = ~pi198 & ~n16357;
  assign n16359 = ~n16356 & ~n16358;
  assign n16360 = pi680 & ~n16359;
  assign n16361 = n16055 & ~n16360;
  assign n16362 = ~pi210 & ~n16357;
  assign n16363 = pi210 & ~n16355;
  assign n16364 = ~n16362 & ~n16363;
  assign n16365 = pi680 & ~n16364;
  assign n16366 = n16051 & ~n16365;
  assign n16367 = ~n16361 & ~n16366;
  assign n16368 = n16057 & ~n16367;
  assign n16369 = ~pi140 & n16368;
  assign n16370 = ~pi39 & ~n16354;
  assign n16371 = ~n16369 & n16370;
  assign n16372 = ~pi38 & ~n16371;
  assign n16373 = ~n16338 & n16372;
  assign n16374 = ~pi738 & ~n16230;
  assign n16375 = ~n16373 & n16374;
  assign n16376 = n9829 & ~n16375;
  assign n16377 = ~n16225 & n16376;
  assign n16378 = ~n16223 & ~n16377;
  assign n16379 = ~pi778 & ~n16378;
  assign n16380 = ~pi625 & n16220;
  assign n16381 = pi625 & n16378;
  assign n16382 = pi1153 & ~n16380;
  assign n16383 = ~n16381 & n16382;
  assign n16384 = ~pi625 & n16378;
  assign n16385 = pi625 & n16220;
  assign n16386 = ~pi1153 & ~n16385;
  assign n16387 = ~n16384 & n16386;
  assign n16388 = ~n16383 & ~n16387;
  assign n16389 = pi778 & ~n16388;
  assign n16390 = ~n16379 & ~n16389;
  assign n16391 = ~n15741 & n16390;
  assign n16392 = n15741 & n16220;
  assign n16393 = ~n16391 & ~n16392;
  assign n16394 = ~n15747 & n16393;
  assign n16395 = ~n16222 & ~n16394;
  assign n16396 = ~n15753 & n16395;
  assign n16397 = n15753 & n16220;
  assign n16398 = ~n16396 & ~n16397;
  assign n16399 = ~n15759 & n16398;
  assign n16400 = ~n16221 & ~n16399;
  assign n16401 = ~pi792 & ~n16400;
  assign n16402 = ~pi628 & ~n16220;
  assign n16403 = pi628 & ~n16400;
  assign n16404 = ~n16402 & ~n16403;
  assign n16405 = pi1156 & ~n16404;
  assign n16406 = ~pi628 & n16400;
  assign n16407 = pi628 & n16220;
  assign n16408 = ~pi1156 & ~n16407;
  assign n16409 = ~n16406 & n16408;
  assign n16410 = ~n16405 & ~n16409;
  assign n16411 = pi792 & ~n16410;
  assign n16412 = ~n16401 & ~n16411;
  assign n16413 = ~pi787 & ~n16412;
  assign n16414 = ~pi647 & n16220;
  assign n16415 = pi647 & n16412;
  assign n16416 = pi1157 & ~n16414;
  assign n16417 = ~n16415 & n16416;
  assign n16418 = ~pi647 & n16412;
  assign n16419 = pi647 & n16220;
  assign n16420 = ~pi1157 & ~n16419;
  assign n16421 = ~n16418 & n16420;
  assign n16422 = ~n16417 & ~n16421;
  assign n16423 = pi787 & ~n16422;
  assign n16424 = ~n16413 & ~n16423;
  assign n16425 = ~pi644 & n16424;
  assign n16426 = ~pi629 & n16405;
  assign n16427 = pi621 & n16030;
  assign n16428 = ~pi210 & ~n16427;
  assign n16429 = pi621 & n16048;
  assign n16430 = pi210 & ~n16429;
  assign n16431 = ~n16428 & ~n16430;
  assign n16432 = pi603 & ~n16431;
  assign n16433 = n16051 & ~n16432;
  assign n16434 = ~pi198 & ~n16427;
  assign n16435 = pi198 & ~n16429;
  assign n16436 = ~n16434 & ~n16435;
  assign n16437 = pi621 & ~n16031;
  assign n16438 = ~n16032 & ~n16437;
  assign n16439 = ~pi198 & n16438;
  assign n16440 = pi621 & ~n16040;
  assign n16441 = ~n16049 & ~n16440;
  assign n16442 = pi198 & n16441;
  assign n16443 = ~n16439 & ~n16442;
  assign n16444 = ~pi603 & ~n16443;
  assign n16445 = ~n16436 & ~n16444;
  assign n16446 = ~n16433 & n16445;
  assign n16447 = n16057 & ~n16446;
  assign n16448 = ~pi39 & ~n16447;
  assign n16449 = ~n15780 & n16063;
  assign n16450 = n3302 & n16449;
  assign n16451 = ~pi614 & ~pi642;
  assign n16452 = ~pi616 & n16451;
  assign n16453 = n16449 & ~n16452;
  assign n16454 = n15779 & n16063;
  assign n16455 = n6166 & ~n16454;
  assign n16456 = n15779 & n16143;
  assign n16457 = ~n6166 & ~n16456;
  assign n16458 = ~n16455 & ~n16457;
  assign n16459 = pi603 & ~n16458;
  assign n16460 = ~n16155 & n16452;
  assign n16461 = ~n16459 & n16460;
  assign n16462 = ~n16453 & ~n16461;
  assign n16463 = ~n6164 & ~n16462;
  assign n16464 = n15780 & n16157;
  assign n16465 = n6164 & ~n16464;
  assign n16466 = n16157 & n16465;
  assign n16467 = ~n16463 & ~n16466;
  assign n16468 = n6221 & ~n16467;
  assign n16469 = ~n15780 & n16153;
  assign n16470 = ~n6221 & n16469;
  assign n16471 = ~n16468 & ~n16470;
  assign n16472 = ~n3302 & ~n16471;
  assign n16473 = ~pi215 & ~n16450;
  assign n16474 = ~n16472 & n16473;
  assign n16475 = pi621 & n16072;
  assign n16476 = ~n6166 & ~n16475;
  assign n16477 = ~n16455 & ~n16476;
  assign n16478 = pi603 & ~n16477;
  assign n16479 = n16460 & ~n16478;
  assign n16480 = ~n16453 & ~n16479;
  assign n16481 = ~n6164 & ~n16480;
  assign n16482 = n6164 & n16085;
  assign n16483 = ~n16478 & n16482;
  assign n16484 = ~n16481 & ~n16483;
  assign n16485 = n6221 & ~n16484;
  assign n16486 = n2923 & ~n15780;
  assign n16487 = ~n16081 & n16486;
  assign n16488 = n6161 & ~n16072;
  assign n16489 = n16487 & ~n16488;
  assign n16490 = ~n6164 & ~n16489;
  assign n16491 = ~n16079 & n16486;
  assign n16492 = n6164 & ~n16491;
  assign n16493 = ~n16490 & ~n16492;
  assign n16494 = ~n6221 & n16493;
  assign n16495 = pi215 & ~n16494;
  assign n16496 = ~n16485 & n16495;
  assign n16497 = ~n16474 & ~n16496;
  assign n16498 = pi299 & ~n16497;
  assign n16499 = n2608 & n16449;
  assign n16500 = n6194 & ~n16467;
  assign n16501 = ~n6194 & n16469;
  assign n16502 = ~n16500 & ~n16501;
  assign n16503 = ~n2608 & ~n16502;
  assign n16504 = ~pi223 & ~n16499;
  assign n16505 = ~n16503 & n16504;
  assign n16506 = n6194 & ~n16484;
  assign n16507 = ~n6194 & n16493;
  assign n16508 = pi223 & ~n16507;
  assign n16509 = ~n16506 & n16508;
  assign n16510 = ~n16505 & ~n16509;
  assign n16511 = ~pi299 & ~n16510;
  assign n16512 = ~n16498 & ~n16511;
  assign n16513 = pi39 & ~n16512;
  assign n16514 = ~n16448 & ~n16513;
  assign n16515 = ~pi761 & n16514;
  assign n16516 = pi761 & n16214;
  assign n16517 = ~pi140 & ~n16515;
  assign n16518 = ~n16516 & n16517;
  assign n16519 = pi603 & ~n16443;
  assign n16520 = ~pi299 & ~n16519;
  assign n16521 = ~pi210 & ~n16438;
  assign n16522 = pi210 & ~n16441;
  assign n16523 = ~n16521 & ~n16522;
  assign n16524 = pi603 & n16523;
  assign n16525 = pi299 & ~n16524;
  assign n16526 = ~n16520 & ~n16525;
  assign n16527 = ~pi39 & ~n16526;
  assign n16528 = n15780 & n16063;
  assign n16529 = ~n16083 & n16528;
  assign n16530 = ~n16081 & n16528;
  assign n16531 = n16083 & n16452;
  assign n16532 = n16530 & ~n16531;
  assign n16533 = ~n6164 & n16532;
  assign n16534 = ~n16529 & ~n16533;
  assign n16535 = ~n16329 & ~n16534;
  assign n16536 = pi223 & ~n16535;
  assign n16537 = n2608 & n16528;
  assign n16538 = n15780 & n16153;
  assign n16539 = ~n6194 & ~n16538;
  assign n16540 = n16452 & ~n16464;
  assign n16541 = ~n16452 & ~n16528;
  assign n16542 = ~n16540 & ~n16541;
  assign n16543 = ~n6164 & ~n16542;
  assign n16544 = ~n16465 & ~n16543;
  assign n16545 = n6194 & ~n16544;
  assign n16546 = ~n2608 & ~n16539;
  assign n16547 = ~n16545 & n16546;
  assign n16548 = ~pi223 & ~n16537;
  assign n16549 = ~n16547 & n16548;
  assign n16550 = ~n16536 & ~n16549;
  assign n16551 = ~pi299 & ~n16550;
  assign n16552 = pi215 & ~n16293;
  assign n16553 = ~n16534 & n16552;
  assign n16554 = n6221 & n16544;
  assign n16555 = ~n6221 & n16538;
  assign n16556 = ~n16554 & ~n16555;
  assign n16557 = ~n3302 & ~n16556;
  assign n16558 = n3302 & n16528;
  assign n16559 = ~n16557 & ~n16558;
  assign n16560 = ~pi215 & ~n16559;
  assign n16561 = pi299 & ~n16553;
  assign n16562 = ~n16560 & n16561;
  assign n16563 = ~n16551 & ~n16562;
  assign n16564 = pi39 & ~n16563;
  assign n16565 = ~n16527 & ~n16564;
  assign n16566 = pi140 & ~pi761;
  assign n16567 = n16565 & n16566;
  assign n16568 = ~n16518 & ~n16567;
  assign n16569 = ~pi38 & ~n16568;
  assign n16570 = n6081 & n15781;
  assign n16571 = ~pi761 & n16570;
  assign n16572 = ~n16229 & ~n16571;
  assign n16573 = pi38 & ~n16572;
  assign n16574 = ~n16569 & ~n16573;
  assign n16575 = n9829 & n16574;
  assign n16576 = ~n16223 & ~n16575;
  assign n16577 = ~n15777 & ~n16576;
  assign n16578 = n15777 & ~n16220;
  assign n16579 = ~n16577 & ~n16578;
  assign n16580 = ~pi785 & ~n16579;
  assign n16581 = ~n15786 & ~n16220;
  assign n16582 = pi609 & n16577;
  assign n16583 = ~n16581 & ~n16582;
  assign n16584 = pi1155 & ~n16583;
  assign n16585 = ~pi609 & ~n15777;
  assign n16586 = ~n16220 & ~n16585;
  assign n16587 = ~pi609 & n16577;
  assign n16588 = ~n16586 & ~n16587;
  assign n16589 = ~pi1155 & ~n16588;
  assign n16590 = ~n16584 & ~n16589;
  assign n16591 = pi785 & ~n16590;
  assign n16592 = ~n16580 & ~n16591;
  assign n16593 = ~pi781 & ~n16592;
  assign n16594 = ~pi618 & n16220;
  assign n16595 = pi618 & n16592;
  assign n16596 = pi1154 & ~n16594;
  assign n16597 = ~n16595 & n16596;
  assign n16598 = ~pi618 & n16592;
  assign n16599 = pi618 & n16220;
  assign n16600 = ~pi1154 & ~n16599;
  assign n16601 = ~n16598 & n16600;
  assign n16602 = ~n16597 & ~n16601;
  assign n16603 = pi781 & ~n16602;
  assign n16604 = ~n16593 & ~n16603;
  assign n16605 = ~pi789 & ~n16604;
  assign n16606 = ~pi619 & n16220;
  assign n16607 = pi619 & n16604;
  assign n16608 = pi1159 & ~n16606;
  assign n16609 = ~n16607 & n16608;
  assign n16610 = ~pi619 & n16604;
  assign n16611 = pi619 & n16220;
  assign n16612 = ~pi1159 & ~n16611;
  assign n16613 = ~n16610 & n16612;
  assign n16614 = ~n16609 & ~n16613;
  assign n16615 = pi789 & ~n16614;
  assign n16616 = ~n16605 & ~n16615;
  assign n16617 = ~pi626 & n16616;
  assign n16618 = pi626 & n16220;
  assign n16619 = ~pi1158 & ~n16618;
  assign n16620 = ~n16617 & n16619;
  assign n16621 = ~pi626 & n16220;
  assign n16622 = pi626 & n16616;
  assign n16623 = pi1158 & ~n16621;
  assign n16624 = ~n16622 & n16623;
  assign n16625 = ~n16620 & ~n16624;
  assign n16626 = pi788 & ~n16625;
  assign n16627 = ~pi788 & ~n16616;
  assign n16628 = ~n16626 & ~n16627;
  assign n16629 = ~pi628 & pi629;
  assign n16630 = pi1156 & n16629;
  assign n16631 = pi628 & ~pi629;
  assign n16632 = ~pi1156 & n16631;
  assign n16633 = ~n16630 & ~n16632;
  assign n16634 = ~n16628 & ~n16633;
  assign n16635 = pi629 & n16409;
  assign n16636 = ~n16426 & ~n16635;
  assign n16637 = ~n16634 & n16636;
  assign n16638 = pi792 & ~n16637;
  assign n16639 = ~pi628 & ~pi629;
  assign n16640 = ~pi1156 & n16639;
  assign n16641 = pi628 & pi629;
  assign n16642 = pi1156 & n16641;
  assign n16643 = ~n16640 & ~n16642;
  assign n16644 = pi792 & n16643;
  assign n16645 = pi618 & ~n16393;
  assign n16646 = pi609 & n16390;
  assign n16647 = n16368 & ~n16446;
  assign n16648 = ~pi140 & n16647;
  assign n16649 = n16354 & ~n16526;
  assign n16650 = ~pi761 & ~n16648;
  assign n16651 = ~n16649 & n16650;
  assign n16652 = pi680 & n16526;
  assign n16653 = ~n16368 & ~n16652;
  assign n16654 = ~pi140 & ~n16653;
  assign n16655 = pi603 & pi665;
  assign n16656 = n16353 & ~n16655;
  assign n16657 = n16447 & n16656;
  assign n16658 = pi140 & ~n16657;
  assign n16659 = pi761 & ~n16654;
  assign n16660 = ~n16658 & n16659;
  assign n16661 = ~n16651 & ~n16660;
  assign n16662 = ~pi39 & ~n16661;
  assign n16663 = ~n15724 & ~n15780;
  assign n16664 = pi680 & n16663;
  assign n16665 = n16063 & ~n16664;
  assign n16666 = n2608 & n16665;
  assign n16667 = pi603 & ~pi621;
  assign n16668 = n16239 & ~n16667;
  assign n16669 = n6164 & ~n16668;
  assign n16670 = n15780 & ~n16144;
  assign n16671 = n16669 & ~n16670;
  assign n16672 = pi680 & ~n16108;
  assign n16673 = ~n16149 & ~n16663;
  assign n16674 = n16672 & ~n16673;
  assign n16675 = ~pi680 & n16149;
  assign n16676 = ~n16671 & ~n16675;
  assign n16677 = ~n16674 & n16676;
  assign n16678 = ~n6194 & n16677;
  assign n16679 = n15724 & ~n16667;
  assign n16680 = n16241 & n16679;
  assign n16681 = n16465 & ~n16680;
  assign n16682 = n16063 & ~n16663;
  assign n16683 = pi616 & ~n16682;
  assign n16684 = pi614 & ~n16682;
  assign n16685 = pi642 & ~n16682;
  assign n16686 = n16159 & ~n16663;
  assign n16687 = ~pi642 & ~n16686;
  assign n16688 = ~n16685 & ~n16687;
  assign n16689 = ~pi614 & ~n16688;
  assign n16690 = ~n16684 & ~n16689;
  assign n16691 = ~pi616 & ~n16690;
  assign n16692 = ~n16683 & ~n16691;
  assign n16693 = n16672 & ~n16692;
  assign n16694 = ~n16236 & ~n16681;
  assign n16695 = ~n16693 & n16694;
  assign n16696 = n6194 & n16695;
  assign n16697 = ~n16678 & ~n16696;
  assign n16698 = ~n2608 & ~n16697;
  assign n16699 = ~pi223 & ~n16666;
  assign n16700 = ~n16698 & n16699;
  assign n16701 = ~n16079 & n16528;
  assign n16702 = ~n16258 & ~n16701;
  assign n16703 = n6164 & n16702;
  assign n16704 = ~n16258 & ~n16268;
  assign n16705 = ~n16530 & n16704;
  assign n16706 = ~pi603 & n16268;
  assign n16707 = n16702 & ~n16706;
  assign n16708 = n16452 & n16707;
  assign n16709 = ~n16705 & ~n16708;
  assign n16710 = n16672 & ~n16709;
  assign n16711 = ~n16703 & ~n16710;
  assign n16712 = ~n16266 & n16711;
  assign n16713 = ~n6194 & n16712;
  assign n16714 = n16261 & ~n16529;
  assign n16715 = n15780 & n16167;
  assign n16716 = n16237 & ~n16667;
  assign n16717 = pi614 & ~n16716;
  assign n16718 = ~n16260 & n16451;
  assign n16719 = ~n16529 & n16718;
  assign n16720 = n16707 & n16719;
  assign n16721 = ~n16685 & ~n16717;
  assign n16722 = ~n16720 & n16721;
  assign n16723 = ~pi616 & ~n16722;
  assign n16724 = ~n16715 & n16723;
  assign n16725 = ~n16683 & ~n16724;
  assign n16726 = n16672 & ~n16725;
  assign n16727 = ~n16257 & ~n16714;
  assign n16728 = ~n16726 & n16727;
  assign n16729 = n6194 & n16728;
  assign n16730 = pi223 & ~n16713;
  assign n16731 = ~n16729 & n16730;
  assign n16732 = ~n16700 & ~n16731;
  assign n16733 = ~pi299 & ~n16732;
  assign n16734 = n3302 & ~n16665;
  assign n16735 = ~pi215 & ~n16734;
  assign n16736 = ~n6221 & n16677;
  assign n16737 = n6221 & n16695;
  assign n16738 = ~n3302 & ~n16736;
  assign n16739 = ~n16737 & n16738;
  assign n16740 = n16735 & ~n16739;
  assign n16741 = ~n6221 & ~n16712;
  assign n16742 = n6221 & ~n16728;
  assign n16743 = pi215 & ~n16741;
  assign n16744 = ~n16742 & n16743;
  assign n16745 = pi299 & ~n16744;
  assign n16746 = ~n16740 & n16745;
  assign n16747 = ~n16733 & ~n16746;
  assign n16748 = ~pi140 & ~n16747;
  assign n16749 = ~n16200 & ~n16735;
  assign n16750 = ~n15780 & n16294;
  assign n16751 = pi616 & ~n16750;
  assign n16752 = n16672 & ~n16751;
  assign n16753 = ~pi603 & ~n16294;
  assign n16754 = ~n16655 & ~n16753;
  assign n16755 = ~n16459 & n16754;
  assign n16756 = n16451 & n16755;
  assign n16757 = ~pi616 & ~n16756;
  assign n16758 = ~n16451 & n16750;
  assign n16759 = n16757 & ~n16758;
  assign n16760 = n16752 & ~n16759;
  assign n16761 = n16157 & n16681;
  assign n16762 = ~n16760 & ~n16761;
  assign n16763 = n6221 & n16762;
  assign n16764 = ~pi665 & n16456;
  assign n16765 = pi603 & ~n16764;
  assign n16766 = n16108 & n16765;
  assign n16767 = pi616 & n15780;
  assign n16768 = ~n16146 & n16663;
  assign n16769 = n16757 & ~n16768;
  assign n16770 = ~n6196 & n16239;
  assign n16771 = ~n16269 & ~n16770;
  assign n16772 = n16679 & ~n16771;
  assign n16773 = ~n16149 & ~n16772;
  assign n16774 = ~n16769 & n16773;
  assign n16775 = ~n16767 & n16774;
  assign n16776 = ~n16108 & ~n16775;
  assign n16777 = ~n15724 & ~n16144;
  assign n16778 = n16108 & ~n16777;
  assign n16779 = pi680 & ~n16778;
  assign n16780 = ~n16766 & n16779;
  assign n16781 = ~n16776 & n16780;
  assign n16782 = ~n6221 & ~n16781;
  assign n16783 = ~n3302 & ~n16763;
  assign n16784 = ~n16782 & n16783;
  assign n16785 = ~n16749 & ~n16784;
  assign n16786 = ~n15724 & ~n16480;
  assign n16787 = ~pi616 & ~n16786;
  assign n16788 = n16752 & ~n16787;
  assign n16789 = n16483 & n16754;
  assign n16790 = ~n16788 & ~n16789;
  assign n16791 = n6221 & ~n16790;
  assign n16792 = n16487 & n16754;
  assign n16793 = ~n16478 & n16754;
  assign n16794 = ~pi642 & ~n16793;
  assign n16795 = n16792 & ~n16794;
  assign n16796 = n6160 & ~n16795;
  assign n16797 = n16792 & ~n16796;
  assign n16798 = ~n16108 & ~n16797;
  assign n16799 = ~n16079 & n16664;
  assign n16800 = ~n16672 & ~n16799;
  assign n16801 = ~n16798 & ~n16800;
  assign n16802 = ~n6221 & n16801;
  assign n16803 = pi215 & ~n16791;
  assign n16804 = ~n16802 & n16803;
  assign n16805 = ~n16785 & ~n16804;
  assign n16806 = pi299 & ~n16805;
  assign n16807 = ~n15725 & ~n15780;
  assign n16808 = n16065 & n16807;
  assign n16809 = ~n16060 & n16808;
  assign n16810 = n2608 & n16809;
  assign n16811 = ~pi223 & ~n16810;
  assign n16812 = ~n16126 & n16811;
  assign n16813 = ~n6194 & n16781;
  assign n16814 = n6194 & ~n16762;
  assign n16815 = ~n2608 & ~n16814;
  assign n16816 = ~n16813 & n16815;
  assign n16817 = ~n16537 & n16812;
  assign n16818 = ~n16816 & n16817;
  assign n16819 = n6194 & n16790;
  assign n16820 = ~n6194 & ~n16801;
  assign n16821 = pi223 & ~n16819;
  assign n16822 = ~n16820 & n16821;
  assign n16823 = ~pi299 & ~n16822;
  assign n16824 = ~n16818 & n16823;
  assign n16825 = ~n16806 & ~n16824;
  assign n16826 = pi140 & n16825;
  assign n16827 = pi761 & ~n16826;
  assign n16828 = ~n16748 & n16827;
  assign n16829 = n3302 & ~n16809;
  assign n16830 = n6164 & ~n16680;
  assign n16831 = ~pi680 & n16462;
  assign n16832 = n15724 & n16461;
  assign n16833 = ~n16452 & n16716;
  assign n16834 = n16672 & ~n16833;
  assign n16835 = ~n16832 & n16834;
  assign n16836 = ~n16830 & ~n16831;
  assign n16837 = ~n16835 & n16836;
  assign n16838 = n6221 & ~n16837;
  assign n16839 = n16672 & ~n16772;
  assign n16840 = ~n15780 & ~n16149;
  assign n16841 = ~pi680 & ~n16840;
  assign n16842 = ~n16669 & ~n16839;
  assign n16843 = ~n16841 & n16842;
  assign n16844 = ~n6221 & ~n16843;
  assign n16845 = ~n16838 & ~n16844;
  assign n16846 = ~n3302 & ~n16845;
  assign n16847 = ~pi215 & ~n16829;
  assign n16848 = ~n16846 & n16847;
  assign n16849 = ~n15725 & n16481;
  assign n16850 = n6164 & ~n16667;
  assign n16851 = n16260 & n16850;
  assign n16852 = ~n16849 & ~n16851;
  assign n16853 = n6221 & n16852;
  assign n16854 = ~pi680 & ~n16489;
  assign n16855 = ~n16480 & ~n16704;
  assign n16856 = n16672 & ~n16855;
  assign n16857 = ~n16267 & ~n16667;
  assign n16858 = n6164 & ~n16857;
  assign n16859 = ~n16854 & ~n16858;
  assign n16860 = ~n16856 & n16859;
  assign n16861 = ~n6221 & ~n16860;
  assign n16862 = pi215 & ~n16853;
  assign n16863 = ~n16861 & n16862;
  assign n16864 = ~n16848 & ~n16863;
  assign n16865 = pi299 & ~n16864;
  assign n16866 = n6194 & ~n16837;
  assign n16867 = ~n6194 & ~n16843;
  assign n16868 = ~n2608 & ~n16867;
  assign n16869 = ~n16866 & n16868;
  assign n16870 = n16811 & ~n16869;
  assign n16871 = ~n6194 & n16860;
  assign n16872 = n6194 & ~n16852;
  assign n16873 = pi223 & ~n16871;
  assign n16874 = ~n16872 & n16873;
  assign n16875 = ~pi299 & ~n16874;
  assign n16876 = ~n16870 & n16875;
  assign n16877 = ~n16865 & ~n16876;
  assign n16878 = ~pi140 & n16877;
  assign n16879 = ~n16300 & n16534;
  assign n16880 = ~n16293 & ~n16879;
  assign n16881 = pi215 & ~n16880;
  assign n16882 = n16199 & ~n16807;
  assign n16883 = ~pi680 & ~n16542;
  assign n16884 = ~n16306 & n16465;
  assign n16885 = n16063 & ~n16679;
  assign n16886 = ~n16452 & n16885;
  assign n16887 = n16159 & n16452;
  assign n16888 = ~n16832 & n16887;
  assign n16889 = n16672 & ~n16886;
  assign n16890 = ~n16888 & n16889;
  assign n16891 = ~n16883 & ~n16884;
  assign n16892 = ~n16890 & n16891;
  assign n16893 = n6221 & ~n16892;
  assign n16894 = ~n16538 & ~n16779;
  assign n16895 = n16672 & ~n16773;
  assign n16896 = ~n16894 & ~n16895;
  assign n16897 = ~n6221 & ~n16896;
  assign n16898 = ~n3302 & ~n16893;
  assign n16899 = ~n16897 & n16898;
  assign n16900 = ~pi215 & ~n16882;
  assign n16901 = ~n16899 & n16900;
  assign n16902 = ~n16881 & ~n16901;
  assign n16903 = pi299 & ~n16902;
  assign n16904 = pi223 & ~n16329;
  assign n16905 = ~n16879 & n16904;
  assign n16906 = ~n6194 & n16896;
  assign n16907 = n6194 & n16892;
  assign n16908 = ~n2608 & ~n16907;
  assign n16909 = ~n16906 & n16908;
  assign n16910 = n16812 & ~n16909;
  assign n16911 = ~pi299 & ~n16905;
  assign n16912 = ~n16910 & n16911;
  assign n16913 = ~n16903 & ~n16912;
  assign n16914 = pi140 & n16913;
  assign n16915 = ~pi761 & ~n16878;
  assign n16916 = ~n16914 & n16915;
  assign n16917 = pi39 & ~n16916;
  assign n16918 = ~n16828 & n16917;
  assign n16919 = ~pi38 & ~n16662;
  assign n16920 = ~n16918 & n16919;
  assign n16921 = n15726 & ~n15780;
  assign n16922 = ~n15782 & ~n16921;
  assign n16923 = n6081 & ~n16922;
  assign n16924 = pi38 & ~n16923;
  assign n16925 = ~n16229 & n16924;
  assign n16926 = ~pi738 & ~n16925;
  assign n16927 = ~n16920 & n16926;
  assign n16928 = pi738 & ~n16574;
  assign n16929 = n9829 & ~n16927;
  assign n16930 = ~n16928 & n16929;
  assign n16931 = ~n16223 & ~n16930;
  assign n16932 = ~pi625 & n16931;
  assign n16933 = pi625 & n16576;
  assign n16934 = ~pi1153 & ~n16933;
  assign n16935 = ~n16932 & n16934;
  assign n16936 = ~pi608 & ~n16383;
  assign n16937 = ~n16935 & n16936;
  assign n16938 = ~pi625 & n16576;
  assign n16939 = pi625 & n16931;
  assign n16940 = pi1153 & ~n16938;
  assign n16941 = ~n16939 & n16940;
  assign n16942 = pi608 & ~n16387;
  assign n16943 = ~n16941 & n16942;
  assign n16944 = ~n16937 & ~n16943;
  assign n16945 = pi778 & ~n16944;
  assign n16946 = ~pi778 & n16931;
  assign n16947 = ~n16945 & ~n16946;
  assign n16948 = ~pi609 & ~n16947;
  assign n16949 = ~pi1155 & ~n16646;
  assign n16950 = ~n16948 & n16949;
  assign n16951 = ~pi660 & ~n16584;
  assign n16952 = ~n16950 & n16951;
  assign n16953 = ~pi609 & n16390;
  assign n16954 = pi609 & ~n16947;
  assign n16955 = pi1155 & ~n16953;
  assign n16956 = ~n16954 & n16955;
  assign n16957 = pi660 & ~n16589;
  assign n16958 = ~n16956 & n16957;
  assign n16959 = ~n16952 & ~n16958;
  assign n16960 = pi785 & ~n16959;
  assign n16961 = ~pi785 & ~n16947;
  assign n16962 = ~n16960 & ~n16961;
  assign n16963 = ~pi618 & ~n16962;
  assign n16964 = ~pi1154 & ~n16645;
  assign n16965 = ~n16963 & n16964;
  assign n16966 = ~pi627 & ~n16597;
  assign n16967 = ~n16965 & n16966;
  assign n16968 = ~pi618 & ~n16393;
  assign n16969 = pi618 & ~n16962;
  assign n16970 = pi1154 & ~n16968;
  assign n16971 = ~n16969 & n16970;
  assign n16972 = pi627 & ~n16601;
  assign n16973 = ~n16971 & n16972;
  assign n16974 = ~n16967 & ~n16973;
  assign n16975 = pi781 & ~n16974;
  assign n16976 = ~pi781 & ~n16962;
  assign n16977 = ~n16975 & ~n16976;
  assign n16978 = ~pi619 & ~n16977;
  assign n16979 = pi619 & n16395;
  assign n16980 = ~pi1159 & ~n16979;
  assign n16981 = ~n16978 & n16980;
  assign n16982 = ~pi648 & ~n16609;
  assign n16983 = ~n16981 & n16982;
  assign n16984 = ~pi619 & n16395;
  assign n16985 = pi619 & ~n16977;
  assign n16986 = pi1159 & ~n16984;
  assign n16987 = ~n16985 & n16986;
  assign n16988 = pi648 & ~n16613;
  assign n16989 = ~n16987 & n16988;
  assign n16990 = ~n16983 & ~n16989;
  assign n16991 = pi789 & ~n16990;
  assign n16992 = ~pi789 & ~n16977;
  assign n16993 = ~n16991 & ~n16992;
  assign n16994 = ~pi788 & ~n16993;
  assign n16995 = ~pi641 & ~pi1158;
  assign n16996 = ~n16620 & ~n16995;
  assign n16997 = ~pi626 & n16993;
  assign n16998 = pi626 & n16398;
  assign n16999 = ~pi641 & ~n16998;
  assign n17000 = ~n16997 & n16999;
  assign n17001 = ~n16996 & ~n17000;
  assign n17002 = pi641 & pi1158;
  assign n17003 = ~n16624 & ~n17002;
  assign n17004 = ~pi626 & n16398;
  assign n17005 = pi626 & n16993;
  assign n17006 = pi641 & ~n17004;
  assign n17007 = ~n17005 & n17006;
  assign n17008 = ~n17003 & ~n17007;
  assign n17009 = pi788 & ~n17001;
  assign n17010 = ~n17008 & n17009;
  assign n17011 = ~n16644 & ~n16994;
  assign n17012 = ~n17010 & n17011;
  assign n17013 = ~n16638 & ~n17012;
  assign n17014 = ~pi647 & n17013;
  assign n17015 = ~n15925 & n16628;
  assign n17016 = n15925 & n16220;
  assign n17017 = ~n17015 & ~n17016;
  assign n17018 = pi647 & ~n17017;
  assign n17019 = ~pi1157 & ~n17018;
  assign n17020 = ~n17014 & n17019;
  assign n17021 = ~pi630 & ~n16417;
  assign n17022 = ~n17020 & n17021;
  assign n17023 = pi647 & n17013;
  assign n17024 = ~pi647 & ~n17017;
  assign n17025 = pi1157 & ~n17024;
  assign n17026 = ~n17023 & n17025;
  assign n17027 = pi630 & ~n16421;
  assign n17028 = ~n17026 & n17027;
  assign n17029 = ~n17022 & ~n17028;
  assign n17030 = pi787 & ~n17029;
  assign n17031 = ~pi787 & n17013;
  assign n17032 = ~n17030 & ~n17031;
  assign n17033 = pi644 & ~n17032;
  assign n17034 = pi715 & ~n16425;
  assign n17035 = ~n17033 & n17034;
  assign n17036 = ~n15960 & ~n17017;
  assign n17037 = n15960 & n16220;
  assign n17038 = ~n17036 & ~n17037;
  assign n17039 = pi644 & ~n17038;
  assign n17040 = ~pi644 & n16220;
  assign n17041 = ~pi715 & ~n17040;
  assign n17042 = ~n17039 & n17041;
  assign n17043 = pi1160 & ~n17042;
  assign n17044 = ~n17035 & n17043;
  assign n17045 = pi644 & n16424;
  assign n17046 = ~pi715 & ~n17045;
  assign n17047 = ~pi644 & ~n17038;
  assign n17048 = pi644 & n16220;
  assign n17049 = pi715 & ~n17048;
  assign n17050 = ~n17047 & n17049;
  assign n17051 = ~pi1160 & ~n17050;
  assign n17052 = ~n17046 & n17051;
  assign n17053 = ~n17044 & ~n17052;
  assign n17054 = pi790 & ~n17053;
  assign n17055 = ~pi644 & n17051;
  assign n17056 = pi790 & ~n17055;
  assign n17057 = ~n17032 & ~n17056;
  assign n17058 = ~n17054 & ~n17057;
  assign n17059 = ~po1038 & ~n17058;
  assign n17060 = ~pi832 & ~n15984;
  assign n17061 = ~n17059 & n17060;
  assign po297 = ~n15983 & ~n17061;
  assign n17063 = ~pi141 & ~n2923;
  assign n17064 = ~pi647 & n17063;
  assign n17065 = pi706 & n15726;
  assign n17066 = ~n17063 & ~n17065;
  assign n17067 = ~pi778 & n17066;
  assign n17068 = ~pi625 & n17065;
  assign n17069 = ~n17066 & ~n17068;
  assign n17070 = pi1153 & ~n17069;
  assign n17071 = ~pi1153 & ~n17063;
  assign n17072 = ~n17068 & n17071;
  assign n17073 = ~n17070 & ~n17072;
  assign n17074 = pi778 & ~n17073;
  assign n17075 = ~n17067 & ~n17074;
  assign n17076 = ~n15742 & n17075;
  assign n17077 = ~n15748 & n17076;
  assign n17078 = ~n15754 & n17077;
  assign n17079 = ~n15760 & n17078;
  assign n17080 = ~n15766 & n17079;
  assign n17081 = pi647 & n17080;
  assign n17082 = pi1157 & ~n17064;
  assign n17083 = ~n17081 & n17082;
  assign n17084 = n15772 & n17079;
  assign n17085 = pi749 & n15781;
  assign n17086 = ~n17063 & ~n17085;
  assign n17087 = ~n15778 & ~n17086;
  assign n17088 = ~pi785 & ~n17087;
  assign n17089 = ~n15787 & ~n17086;
  assign n17090 = pi1155 & ~n17089;
  assign n17091 = ~n15790 & n17087;
  assign n17092 = ~pi1155 & ~n17091;
  assign n17093 = ~n17090 & ~n17092;
  assign n17094 = pi785 & ~n17093;
  assign n17095 = ~n17088 & ~n17094;
  assign n17096 = ~pi781 & ~n17095;
  assign n17097 = ~n15797 & n17095;
  assign n17098 = pi1154 & ~n17097;
  assign n17099 = ~n15800 & n17095;
  assign n17100 = ~pi1154 & ~n17099;
  assign n17101 = ~n17098 & ~n17100;
  assign n17102 = pi781 & ~n17101;
  assign n17103 = ~n17096 & ~n17102;
  assign n17104 = ~pi789 & ~n17103;
  assign n17105 = ~pi619 & n17063;
  assign n17106 = pi619 & n17103;
  assign n17107 = pi1159 & ~n17105;
  assign n17108 = ~n17106 & n17107;
  assign n17109 = ~pi619 & n17103;
  assign n17110 = pi619 & n17063;
  assign n17111 = ~pi1159 & ~n17110;
  assign n17112 = ~n17109 & n17111;
  assign n17113 = ~n17108 & ~n17112;
  assign n17114 = pi789 & ~n17113;
  assign n17115 = ~n17104 & ~n17114;
  assign n17116 = n15820 & n17115;
  assign n17117 = ~n15820 & n17063;
  assign n17118 = ~n17116 & ~n17117;
  assign n17119 = ~n15758 & ~n17118;
  assign n17120 = n15828 & n17078;
  assign n17121 = ~n17119 & ~n17120;
  assign n17122 = pi788 & ~n17121;
  assign n17123 = pi618 & n17076;
  assign n17124 = pi609 & n17075;
  assign n17125 = ~n15780 & ~n17066;
  assign n17126 = pi625 & n17125;
  assign n17127 = n17086 & ~n17125;
  assign n17128 = ~n17126 & ~n17127;
  assign n17129 = n17071 & ~n17128;
  assign n17130 = ~pi608 & ~n17070;
  assign n17131 = ~n17129 & n17130;
  assign n17132 = pi1153 & n17086;
  assign n17133 = ~n17126 & n17132;
  assign n17134 = pi608 & ~n17072;
  assign n17135 = ~n17133 & n17134;
  assign n17136 = ~n17131 & ~n17135;
  assign n17137 = pi778 & ~n17136;
  assign n17138 = ~pi778 & ~n17127;
  assign n17139 = ~n17137 & ~n17138;
  assign n17140 = ~pi609 & ~n17139;
  assign n17141 = ~pi1155 & ~n17124;
  assign n17142 = ~n17140 & n17141;
  assign n17143 = ~pi660 & ~n17090;
  assign n17144 = ~n17142 & n17143;
  assign n17145 = ~pi609 & n17075;
  assign n17146 = pi609 & ~n17139;
  assign n17147 = pi1155 & ~n17145;
  assign n17148 = ~n17146 & n17147;
  assign n17149 = pi660 & ~n17092;
  assign n17150 = ~n17148 & n17149;
  assign n17151 = ~n17144 & ~n17150;
  assign n17152 = pi785 & ~n17151;
  assign n17153 = ~pi785 & ~n17139;
  assign n17154 = ~n17152 & ~n17153;
  assign n17155 = ~pi618 & ~n17154;
  assign n17156 = ~pi1154 & ~n17123;
  assign n17157 = ~n17155 & n17156;
  assign n17158 = ~pi627 & ~n17098;
  assign n17159 = ~n17157 & n17158;
  assign n17160 = ~pi618 & n17076;
  assign n17161 = pi618 & ~n17154;
  assign n17162 = pi1154 & ~n17160;
  assign n17163 = ~n17161 & n17162;
  assign n17164 = pi627 & ~n17100;
  assign n17165 = ~n17163 & n17164;
  assign n17166 = ~n17159 & ~n17165;
  assign n17167 = pi781 & ~n17166;
  assign n17168 = ~pi781 & ~n17154;
  assign n17169 = ~n17167 & ~n17168;
  assign n17170 = ~pi789 & n17169;
  assign n17171 = ~pi619 & n17077;
  assign n17172 = pi619 & ~n17169;
  assign n17173 = pi1159 & ~n17171;
  assign n17174 = ~n17172 & n17173;
  assign n17175 = pi648 & ~n17112;
  assign n17176 = ~n17174 & n17175;
  assign n17177 = pi619 & n17077;
  assign n17178 = ~pi619 & ~n17169;
  assign n17179 = ~pi1159 & ~n17177;
  assign n17180 = ~n17178 & n17179;
  assign n17181 = ~pi648 & ~n17108;
  assign n17182 = ~n17180 & n17181;
  assign n17183 = pi789 & ~n17176;
  assign n17184 = ~n17182 & n17183;
  assign n17185 = n15833 & ~n17170;
  assign n17186 = ~n17184 & n17185;
  assign n17187 = ~n17122 & ~n17186;
  assign n17188 = ~pi628 & n17187;
  assign n17189 = pi788 & ~n17118;
  assign n17190 = ~pi788 & n17115;
  assign n17191 = ~n17189 & ~n17190;
  assign n17192 = pi628 & n17191;
  assign n17193 = ~pi1156 & ~n17192;
  assign n17194 = ~n17188 & n17193;
  assign n17195 = ~pi629 & ~n17084;
  assign n17196 = ~n17194 & n17195;
  assign n17197 = n15909 & n17079;
  assign n17198 = ~pi628 & n17191;
  assign n17199 = pi628 & n17187;
  assign n17200 = pi1156 & ~n17198;
  assign n17201 = ~n17199 & n17200;
  assign n17202 = pi629 & ~n17197;
  assign n17203 = ~n17201 & n17202;
  assign n17204 = ~n17196 & ~n17203;
  assign n17205 = pi792 & ~n17204;
  assign n17206 = ~pi792 & n17187;
  assign n17207 = ~n17205 & ~n17206;
  assign n17208 = ~pi647 & n17207;
  assign n17209 = n15925 & ~n17063;
  assign n17210 = ~n15925 & n17191;
  assign n17211 = ~n17209 & ~n17210;
  assign n17212 = pi647 & n17211;
  assign n17213 = ~pi1157 & ~n17212;
  assign n17214 = ~n17208 & n17213;
  assign n17215 = ~pi630 & ~n17083;
  assign n17216 = ~n17214 & n17215;
  assign n17217 = ~pi647 & n17080;
  assign n17218 = pi647 & n17063;
  assign n17219 = ~pi1157 & ~n17218;
  assign n17220 = ~n17217 & n17219;
  assign n17221 = ~pi647 & n17211;
  assign n17222 = pi647 & n17207;
  assign n17223 = pi1157 & ~n17221;
  assign n17224 = ~n17222 & n17223;
  assign n17225 = pi630 & ~n17220;
  assign n17226 = ~n17224 & n17225;
  assign n17227 = ~n17216 & ~n17226;
  assign n17228 = pi787 & ~n17227;
  assign n17229 = ~pi787 & n17207;
  assign n17230 = ~n17228 & ~n17229;
  assign n17231 = ~pi790 & ~n17230;
  assign n17232 = ~pi787 & ~n17080;
  assign n17233 = ~n17083 & ~n17220;
  assign n17234 = pi787 & ~n17233;
  assign n17235 = ~n17232 & ~n17234;
  assign n17236 = ~pi644 & n17235;
  assign n17237 = pi644 & ~n17230;
  assign n17238 = pi715 & ~n17236;
  assign n17239 = ~n17237 & n17238;
  assign n17240 = ~n15960 & n17211;
  assign n17241 = n15960 & n17063;
  assign n17242 = ~n17240 & ~n17241;
  assign n17243 = pi644 & ~n17242;
  assign n17244 = ~pi644 & n17063;
  assign n17245 = ~pi715 & ~n17244;
  assign n17246 = ~n17243 & n17245;
  assign n17247 = pi1160 & ~n17246;
  assign n17248 = ~n17239 & n17247;
  assign n17249 = ~pi644 & ~n17242;
  assign n17250 = pi644 & n17063;
  assign n17251 = pi715 & ~n17250;
  assign n17252 = ~n17249 & n17251;
  assign n17253 = pi644 & n17235;
  assign n17254 = ~pi644 & ~n17230;
  assign n17255 = ~pi715 & ~n17253;
  assign n17256 = ~n17254 & n17255;
  assign n17257 = ~pi1160 & ~n17252;
  assign n17258 = ~n17256 & n17257;
  assign n17259 = ~n17248 & ~n17258;
  assign n17260 = pi790 & ~n17259;
  assign n17261 = pi832 & ~n17231;
  assign n17262 = ~n17260 & n17261;
  assign n17263 = ~pi141 & po1038;
  assign n17264 = ~pi141 & ~n16219;
  assign n17265 = n15759 & ~n17264;
  assign n17266 = n15747 & ~n17264;
  assign n17267 = pi141 & ~n9829;
  assign n17268 = ~pi141 & ~n16228;
  assign n17269 = n16227 & ~n17268;
  assign n17270 = ~pi39 & ~n16353;
  assign n17271 = pi39 & ~n16335;
  assign n17272 = ~n17270 & ~n17271;
  assign n17273 = pi141 & n17272;
  assign n17274 = ~pi39 & ~n16368;
  assign n17275 = pi39 & ~n16291;
  assign n17276 = ~n17274 & ~n17275;
  assign n17277 = ~pi141 & ~n17276;
  assign n17278 = ~pi38 & ~n17273;
  assign n17279 = ~n17277 & n17278;
  assign n17280 = pi706 & ~n17269;
  assign n17281 = ~n17279 & n17280;
  assign n17282 = ~pi141 & ~pi706;
  assign n17283 = ~n16218 & n17282;
  assign n17284 = n9829 & ~n17281;
  assign n17285 = ~n17283 & n17284;
  assign n17286 = ~n17267 & ~n17285;
  assign n17287 = ~pi778 & ~n17286;
  assign n17288 = ~pi625 & n17264;
  assign n17289 = pi625 & n17286;
  assign n17290 = pi1153 & ~n17288;
  assign n17291 = ~n17289 & n17290;
  assign n17292 = ~pi625 & n17286;
  assign n17293 = pi625 & n17264;
  assign n17294 = ~pi1153 & ~n17293;
  assign n17295 = ~n17292 & n17294;
  assign n17296 = ~n17291 & ~n17295;
  assign n17297 = pi778 & ~n17296;
  assign n17298 = ~n17287 & ~n17297;
  assign n17299 = ~n15741 & n17298;
  assign n17300 = n15741 & n17264;
  assign n17301 = ~n17299 & ~n17300;
  assign n17302 = ~n15747 & n17301;
  assign n17303 = ~n17266 & ~n17302;
  assign n17304 = ~n15753 & n17303;
  assign n17305 = n15753 & n17264;
  assign n17306 = ~n17304 & ~n17305;
  assign n17307 = ~n15759 & n17306;
  assign n17308 = ~n17265 & ~n17307;
  assign n17309 = ~pi792 & ~n17308;
  assign n17310 = ~pi628 & ~n17264;
  assign n17311 = pi628 & ~n17308;
  assign n17312 = ~n17310 & ~n17311;
  assign n17313 = pi1156 & ~n17312;
  assign n17314 = ~pi628 & n17308;
  assign n17315 = pi628 & n17264;
  assign n17316 = ~pi1156 & ~n17315;
  assign n17317 = ~n17314 & n17316;
  assign n17318 = ~n17313 & ~n17317;
  assign n17319 = pi792 & ~n17318;
  assign n17320 = ~n17309 & ~n17319;
  assign n17321 = ~pi787 & ~n17320;
  assign n17322 = ~pi647 & n17264;
  assign n17323 = pi647 & n17320;
  assign n17324 = pi1157 & ~n17322;
  assign n17325 = ~n17323 & n17324;
  assign n17326 = ~pi647 & n17320;
  assign n17327 = pi647 & n17264;
  assign n17328 = ~pi1157 & ~n17327;
  assign n17329 = ~n17326 & n17328;
  assign n17330 = ~n17325 & ~n17329;
  assign n17331 = pi787 & ~n17330;
  assign n17332 = ~n17321 & ~n17331;
  assign n17333 = ~pi644 & n17332;
  assign n17334 = ~pi629 & n17313;
  assign n17335 = ~pi619 & n17264;
  assign n17336 = pi749 & n16570;
  assign n17337 = ~n17268 & ~n17336;
  assign n17338 = pi38 & ~n17337;
  assign n17339 = ~pi749 & n16212;
  assign n17340 = pi141 & ~n16563;
  assign n17341 = ~n17339 & ~n17340;
  assign n17342 = pi39 & ~n17341;
  assign n17343 = ~pi141 & n16514;
  assign n17344 = pi141 & n16527;
  assign n17345 = pi749 & ~n17344;
  assign n17346 = ~n17343 & n17345;
  assign n17347 = ~pi39 & n16057;
  assign n17348 = ~pi141 & ~pi749;
  assign n17349 = ~n17347 & n17348;
  assign n17350 = ~n17346 & ~n17349;
  assign n17351 = ~pi38 & ~n17350;
  assign n17352 = ~n17342 & n17351;
  assign n17353 = ~n17338 & ~n17352;
  assign n17354 = n9829 & n17353;
  assign n17355 = ~n17267 & ~n17354;
  assign n17356 = ~n15777 & ~n17355;
  assign n17357 = n15777 & ~n17264;
  assign n17358 = ~n17356 & ~n17357;
  assign n17359 = ~pi785 & ~n17358;
  assign n17360 = ~n15786 & ~n17264;
  assign n17361 = pi609 & n17356;
  assign n17362 = ~n17360 & ~n17361;
  assign n17363 = pi1155 & ~n17362;
  assign n17364 = ~n16585 & ~n17264;
  assign n17365 = ~pi609 & n17356;
  assign n17366 = ~n17364 & ~n17365;
  assign n17367 = ~pi1155 & ~n17366;
  assign n17368 = ~n17363 & ~n17367;
  assign n17369 = pi785 & ~n17368;
  assign n17370 = ~n17359 & ~n17369;
  assign n17371 = ~pi781 & ~n17370;
  assign n17372 = ~pi618 & n17264;
  assign n17373 = pi618 & n17370;
  assign n17374 = pi1154 & ~n17372;
  assign n17375 = ~n17373 & n17374;
  assign n17376 = ~pi618 & n17370;
  assign n17377 = pi618 & n17264;
  assign n17378 = ~pi1154 & ~n17377;
  assign n17379 = ~n17376 & n17378;
  assign n17380 = ~n17375 & ~n17379;
  assign n17381 = pi781 & ~n17380;
  assign n17382 = ~n17371 & ~n17381;
  assign n17383 = pi619 & n17382;
  assign n17384 = pi1159 & ~n17335;
  assign n17385 = ~n17383 & n17384;
  assign n17386 = pi618 & ~n17301;
  assign n17387 = pi609 & n17298;
  assign n17388 = ~pi706 & ~n17353;
  assign n17389 = ~n15780 & n16226;
  assign n17390 = pi38 & ~n17389;
  assign n17391 = n17337 & n17390;
  assign n17392 = ~pi141 & n16653;
  assign n17393 = pi141 & n16657;
  assign n17394 = ~pi749 & ~n17392;
  assign n17395 = ~n17393 & n17394;
  assign n17396 = ~pi141 & ~n16647;
  assign n17397 = ~n16353 & ~n16526;
  assign n17398 = pi141 & ~n17397;
  assign n17399 = pi749 & ~n17396;
  assign n17400 = ~n17398 & n17399;
  assign n17401 = ~pi39 & ~n17400;
  assign n17402 = ~n17395 & n17401;
  assign n17403 = ~pi141 & n16877;
  assign n17404 = pi141 & n16913;
  assign n17405 = pi749 & ~n17403;
  assign n17406 = ~n17404 & n17405;
  assign n17407 = pi141 & n16825;
  assign n17408 = ~pi141 & ~n16747;
  assign n17409 = ~pi749 & ~n17407;
  assign n17410 = ~n17408 & n17409;
  assign n17411 = pi39 & ~n17406;
  assign n17412 = ~n17410 & n17411;
  assign n17413 = ~pi38 & ~n17402;
  assign n17414 = ~n17412 & n17413;
  assign n17415 = pi706 & ~n17391;
  assign n17416 = ~n17414 & n17415;
  assign n17417 = n9829 & ~n17416;
  assign n17418 = ~n17388 & n17417;
  assign n17419 = ~n17267 & ~n17418;
  assign n17420 = ~pi625 & n17419;
  assign n17421 = pi625 & n17355;
  assign n17422 = ~pi1153 & ~n17421;
  assign n17423 = ~n17420 & n17422;
  assign n17424 = ~pi608 & ~n17291;
  assign n17425 = ~n17423 & n17424;
  assign n17426 = ~pi625 & n17355;
  assign n17427 = pi625 & n17419;
  assign n17428 = pi1153 & ~n17426;
  assign n17429 = ~n17427 & n17428;
  assign n17430 = pi608 & ~n17295;
  assign n17431 = ~n17429 & n17430;
  assign n17432 = ~n17425 & ~n17431;
  assign n17433 = pi778 & ~n17432;
  assign n17434 = ~pi778 & n17419;
  assign n17435 = ~n17433 & ~n17434;
  assign n17436 = ~pi609 & ~n17435;
  assign n17437 = ~pi1155 & ~n17387;
  assign n17438 = ~n17436 & n17437;
  assign n17439 = ~pi660 & ~n17363;
  assign n17440 = ~n17438 & n17439;
  assign n17441 = ~pi609 & n17298;
  assign n17442 = pi609 & ~n17435;
  assign n17443 = pi1155 & ~n17441;
  assign n17444 = ~n17442 & n17443;
  assign n17445 = pi660 & ~n17367;
  assign n17446 = ~n17444 & n17445;
  assign n17447 = ~n17440 & ~n17446;
  assign n17448 = pi785 & ~n17447;
  assign n17449 = ~pi785 & ~n17435;
  assign n17450 = ~n17448 & ~n17449;
  assign n17451 = ~pi618 & ~n17450;
  assign n17452 = ~pi1154 & ~n17386;
  assign n17453 = ~n17451 & n17452;
  assign n17454 = ~pi627 & ~n17375;
  assign n17455 = ~n17453 & n17454;
  assign n17456 = ~pi618 & ~n17301;
  assign n17457 = pi618 & ~n17450;
  assign n17458 = pi1154 & ~n17456;
  assign n17459 = ~n17457 & n17458;
  assign n17460 = pi627 & ~n17379;
  assign n17461 = ~n17459 & n17460;
  assign n17462 = ~n17455 & ~n17461;
  assign n17463 = pi781 & ~n17462;
  assign n17464 = ~pi781 & ~n17450;
  assign n17465 = ~n17463 & ~n17464;
  assign n17466 = ~pi619 & ~n17465;
  assign n17467 = pi619 & n17303;
  assign n17468 = ~pi1159 & ~n17467;
  assign n17469 = ~n17466 & n17468;
  assign n17470 = ~pi648 & ~n17385;
  assign n17471 = ~n17469 & n17470;
  assign n17472 = ~pi619 & n17382;
  assign n17473 = pi619 & n17264;
  assign n17474 = ~pi1159 & ~n17473;
  assign n17475 = ~n17472 & n17474;
  assign n17476 = ~pi619 & n17303;
  assign n17477 = pi619 & ~n17465;
  assign n17478 = pi1159 & ~n17476;
  assign n17479 = ~n17477 & n17478;
  assign n17480 = pi648 & ~n17475;
  assign n17481 = ~n17479 & n17480;
  assign n17482 = ~n17471 & ~n17481;
  assign n17483 = pi789 & ~n17482;
  assign n17484 = ~pi789 & ~n17465;
  assign n17485 = ~n17483 & ~n17484;
  assign n17486 = ~pi788 & n17485;
  assign n17487 = ~pi789 & ~n17382;
  assign n17488 = ~n17385 & ~n17475;
  assign n17489 = pi789 & ~n17488;
  assign n17490 = ~n17487 & ~n17489;
  assign n17491 = ~pi626 & n17490;
  assign n17492 = pi626 & n17264;
  assign n17493 = ~pi1158 & ~n17492;
  assign n17494 = ~n17491 & n17493;
  assign n17495 = ~n16995 & ~n17494;
  assign n17496 = ~pi626 & n17485;
  assign n17497 = pi626 & n17306;
  assign n17498 = ~pi641 & ~n17497;
  assign n17499 = ~n17496 & n17498;
  assign n17500 = ~n17495 & ~n17499;
  assign n17501 = ~pi626 & n17264;
  assign n17502 = pi626 & n17490;
  assign n17503 = pi1158 & ~n17501;
  assign n17504 = ~n17502 & n17503;
  assign n17505 = ~n17002 & ~n17504;
  assign n17506 = ~pi626 & n17306;
  assign n17507 = pi626 & n17485;
  assign n17508 = pi641 & ~n17506;
  assign n17509 = ~n17507 & n17508;
  assign n17510 = ~n17505 & ~n17509;
  assign n17511 = ~n17500 & ~n17510;
  assign n17512 = pi788 & ~n17511;
  assign n17513 = ~n17486 & ~n17512;
  assign n17514 = ~n16643 & ~n17513;
  assign n17515 = ~n17494 & ~n17504;
  assign n17516 = pi788 & ~n17515;
  assign n17517 = ~pi788 & ~n17490;
  assign n17518 = ~n17516 & ~n17517;
  assign n17519 = ~n16633 & ~n17518;
  assign n17520 = pi629 & n17317;
  assign n17521 = ~n17334 & ~n17520;
  assign n17522 = ~n17519 & n17521;
  assign n17523 = ~n17514 & n17522;
  assign n17524 = pi792 & ~n17523;
  assign n17525 = ~pi792 & ~n17513;
  assign n17526 = ~n17524 & ~n17525;
  assign n17527 = ~pi647 & n17526;
  assign n17528 = ~n15925 & n17518;
  assign n17529 = n15925 & n17264;
  assign n17530 = ~n17528 & ~n17529;
  assign n17531 = pi647 & ~n17530;
  assign n17532 = ~pi1157 & ~n17531;
  assign n17533 = ~n17527 & n17532;
  assign n17534 = ~pi630 & ~n17325;
  assign n17535 = ~n17533 & n17534;
  assign n17536 = ~pi647 & ~n17530;
  assign n17537 = pi647 & n17526;
  assign n17538 = pi1157 & ~n17536;
  assign n17539 = ~n17537 & n17538;
  assign n17540 = pi630 & ~n17329;
  assign n17541 = ~n17539 & n17540;
  assign n17542 = ~n17535 & ~n17541;
  assign n17543 = pi787 & ~n17542;
  assign n17544 = ~pi787 & n17526;
  assign n17545 = ~n17543 & ~n17544;
  assign n17546 = pi644 & ~n17545;
  assign n17547 = pi715 & ~n17333;
  assign n17548 = ~n17546 & n17547;
  assign n17549 = ~n15960 & ~n17530;
  assign n17550 = n15960 & n17264;
  assign n17551 = ~n17549 & ~n17550;
  assign n17552 = pi644 & ~n17551;
  assign n17553 = ~pi644 & n17264;
  assign n17554 = ~pi715 & ~n17553;
  assign n17555 = ~n17552 & n17554;
  assign n17556 = pi1160 & ~n17555;
  assign n17557 = ~n17548 & n17556;
  assign n17558 = pi644 & n17332;
  assign n17559 = ~pi715 & ~n17558;
  assign n17560 = ~pi644 & ~n17551;
  assign n17561 = pi644 & n17264;
  assign n17562 = pi715 & ~n17561;
  assign n17563 = ~n17560 & n17562;
  assign n17564 = ~pi1160 & ~n17563;
  assign n17565 = ~n17559 & n17564;
  assign n17566 = ~n17557 & ~n17565;
  assign n17567 = pi790 & ~n17566;
  assign n17568 = ~pi644 & n17564;
  assign n17569 = pi790 & ~n17568;
  assign n17570 = ~n17545 & ~n17569;
  assign n17571 = ~n17567 & ~n17570;
  assign n17572 = ~po1038 & ~n17571;
  assign n17573 = ~pi832 & ~n17263;
  assign n17574 = ~n17572 & n17573;
  assign po298 = ~n17262 & ~n17574;
  assign n17576 = pi142 & ~n2923;
  assign n17577 = pi735 & n15726;
  assign n17578 = ~pi625 & ~pi1153;
  assign n17579 = pi625 & pi1153;
  assign n17580 = pi778 & ~n17578;
  assign n17581 = ~n17579 & n17580;
  assign n17582 = n17577 & ~n17581;
  assign n17583 = ~n17576 & ~n17582;
  assign n17584 = ~n15741 & ~n15747;
  assign n17585 = ~n15753 & ~n15759;
  assign n17586 = n17584 & n17585;
  assign n17587 = ~n17583 & n17586;
  assign n17588 = ~n15765 & n17587;
  assign n17589 = pi647 & n17588;
  assign n17590 = ~n17576 & ~n17589;
  assign n17591 = pi1157 & ~n17590;
  assign n17592 = pi743 & n15781;
  assign n17593 = ~n15777 & n17592;
  assign n17594 = pi609 & n17593;
  assign n17595 = pi1155 & ~n17576;
  assign n17596 = ~n17594 & n17595;
  assign n17597 = ~pi609 & n17593;
  assign n17598 = ~pi1155 & ~n17576;
  assign n17599 = ~n17597 & n17598;
  assign n17600 = ~n17596 & ~n17599;
  assign n17601 = pi785 & ~n17600;
  assign n17602 = ~pi785 & ~n17576;
  assign n17603 = ~n17593 & n17602;
  assign n17604 = ~n17601 & ~n17603;
  assign n17605 = ~pi781 & ~n17604;
  assign n17606 = ~pi618 & n17576;
  assign n17607 = pi618 & n17604;
  assign n17608 = pi1154 & ~n17606;
  assign n17609 = ~n17607 & n17608;
  assign n17610 = ~pi618 & n17604;
  assign n17611 = pi618 & n17576;
  assign n17612 = ~pi1154 & ~n17611;
  assign n17613 = ~n17610 & n17612;
  assign n17614 = ~n17609 & ~n17613;
  assign n17615 = pi781 & ~n17614;
  assign n17616 = ~n17605 & ~n17615;
  assign n17617 = ~pi789 & ~n17616;
  assign n17618 = ~pi619 & n17576;
  assign n17619 = pi619 & n17616;
  assign n17620 = pi1159 & ~n17618;
  assign n17621 = ~n17619 & n17620;
  assign n17622 = ~pi619 & n17616;
  assign n17623 = pi619 & n17576;
  assign n17624 = ~pi1159 & ~n17623;
  assign n17625 = ~n17622 & n17624;
  assign n17626 = ~n17621 & ~n17625;
  assign n17627 = pi789 & ~n17626;
  assign n17628 = ~n17617 & ~n17627;
  assign n17629 = n15820 & n17628;
  assign n17630 = ~n15820 & n17576;
  assign n17631 = ~n17629 & ~n17630;
  assign n17632 = pi788 & ~n17631;
  assign n17633 = ~pi788 & n17628;
  assign n17634 = ~n17632 & ~n17633;
  assign n17635 = pi628 & ~n17634;
  assign n17636 = ~n15758 & ~n17631;
  assign n17637 = ~n15742 & ~n17583;
  assign n17638 = ~n15748 & n17637;
  assign n17639 = ~n15754 & n15828;
  assign n17640 = n17638 & n17639;
  assign n17641 = ~n17636 & ~n17640;
  assign n17642 = pi788 & ~n17641;
  assign n17643 = pi618 & n17637;
  assign n17644 = pi609 & ~n17583;
  assign n17645 = pi625 & n17577;
  assign n17646 = pi1153 & ~n17576;
  assign n17647 = ~n17645 & n17646;
  assign n17648 = pi735 & n16921;
  assign n17649 = pi625 & n17648;
  assign n17650 = ~n17576 & ~n17592;
  assign n17651 = ~n17648 & n17650;
  assign n17652 = ~n17649 & ~n17651;
  assign n17653 = ~pi1153 & ~n17652;
  assign n17654 = ~pi608 & ~n17647;
  assign n17655 = ~n17653 & n17654;
  assign n17656 = ~n17592 & ~n17649;
  assign n17657 = pi1153 & ~n17656;
  assign n17658 = n17577 & n17578;
  assign n17659 = ~n17576 & ~n17658;
  assign n17660 = ~n17657 & n17659;
  assign n17661 = pi608 & ~n17660;
  assign n17662 = ~n17655 & ~n17661;
  assign n17663 = pi778 & ~n17662;
  assign n17664 = ~pi778 & ~n17651;
  assign n17665 = ~n17663 & ~n17664;
  assign n17666 = ~pi609 & ~n17665;
  assign n17667 = ~pi1155 & ~n17644;
  assign n17668 = ~n17666 & n17667;
  assign n17669 = ~pi660 & ~n17596;
  assign n17670 = ~n17668 & n17669;
  assign n17671 = ~pi609 & ~n17583;
  assign n17672 = pi609 & ~n17665;
  assign n17673 = pi1155 & ~n17671;
  assign n17674 = ~n17672 & n17673;
  assign n17675 = pi660 & ~n17599;
  assign n17676 = ~n17674 & n17675;
  assign n17677 = ~n17670 & ~n17676;
  assign n17678 = pi785 & ~n17677;
  assign n17679 = ~pi785 & ~n17665;
  assign n17680 = ~n17678 & ~n17679;
  assign n17681 = ~pi618 & ~n17680;
  assign n17682 = ~pi1154 & ~n17643;
  assign n17683 = ~n17681 & n17682;
  assign n17684 = ~pi627 & ~n17609;
  assign n17685 = ~n17683 & n17684;
  assign n17686 = ~pi618 & n17637;
  assign n17687 = pi618 & ~n17680;
  assign n17688 = pi1154 & ~n17686;
  assign n17689 = ~n17687 & n17688;
  assign n17690 = pi627 & ~n17613;
  assign n17691 = ~n17689 & n17690;
  assign n17692 = ~n17685 & ~n17691;
  assign n17693 = pi781 & ~n17692;
  assign n17694 = ~pi781 & ~n17680;
  assign n17695 = ~n17693 & ~n17694;
  assign n17696 = ~pi789 & n17695;
  assign n17697 = pi619 & n17638;
  assign n17698 = ~pi619 & ~n17695;
  assign n17699 = ~pi1159 & ~n17697;
  assign n17700 = ~n17698 & n17699;
  assign n17701 = ~pi648 & ~n17621;
  assign n17702 = ~n17700 & n17701;
  assign n17703 = ~pi619 & n17638;
  assign n17704 = pi619 & ~n17695;
  assign n17705 = pi1159 & ~n17703;
  assign n17706 = ~n17704 & n17705;
  assign n17707 = pi648 & ~n17625;
  assign n17708 = ~n17706 & n17707;
  assign n17709 = pi789 & ~n17702;
  assign n17710 = ~n17708 & n17709;
  assign n17711 = n15833 & ~n17696;
  assign n17712 = ~n17710 & n17711;
  assign n17713 = ~n17642 & ~n17712;
  assign n17714 = ~pi628 & ~n17713;
  assign n17715 = ~pi1156 & ~n17635;
  assign n17716 = ~n17714 & n17715;
  assign n17717 = pi628 & n17587;
  assign n17718 = pi1156 & ~n17576;
  assign n17719 = ~n17717 & n17718;
  assign n17720 = ~pi629 & ~n17719;
  assign n17721 = ~n17716 & n17720;
  assign n17722 = ~pi628 & ~n17634;
  assign n17723 = pi628 & ~n17713;
  assign n17724 = pi1156 & ~n17722;
  assign n17725 = ~n17723 & n17724;
  assign n17726 = ~pi628 & n17587;
  assign n17727 = ~pi1156 & ~n17576;
  assign n17728 = ~n17726 & n17727;
  assign n17729 = pi629 & ~n17728;
  assign n17730 = ~n17725 & n17729;
  assign n17731 = ~n17721 & ~n17730;
  assign n17732 = pi792 & ~n17731;
  assign n17733 = ~pi792 & ~n17713;
  assign n17734 = ~n17732 & ~n17733;
  assign n17735 = ~pi647 & n17734;
  assign n17736 = n15925 & ~n17576;
  assign n17737 = ~n15925 & n17634;
  assign n17738 = ~n17736 & ~n17737;
  assign n17739 = pi647 & ~n17738;
  assign n17740 = ~pi1157 & ~n17739;
  assign n17741 = ~n17735 & n17740;
  assign n17742 = ~pi630 & ~n17591;
  assign n17743 = ~n17741 & n17742;
  assign n17744 = ~pi647 & n17588;
  assign n17745 = ~n17576 & ~n17744;
  assign n17746 = ~pi1157 & ~n17745;
  assign n17747 = ~pi647 & ~n17738;
  assign n17748 = pi647 & n17734;
  assign n17749 = pi1157 & ~n17747;
  assign n17750 = ~n17748 & n17749;
  assign n17751 = pi630 & ~n17746;
  assign n17752 = ~n17750 & n17751;
  assign n17753 = ~n17743 & ~n17752;
  assign n17754 = pi787 & ~n17753;
  assign n17755 = ~pi787 & n17734;
  assign n17756 = ~n17754 & ~n17755;
  assign n17757 = ~pi790 & n17756;
  assign n17758 = ~n15960 & n17738;
  assign n17759 = n15960 & n17576;
  assign n17760 = ~n17758 & ~n17759;
  assign n17761 = pi644 & ~n17760;
  assign n17762 = ~pi644 & n17576;
  assign n17763 = ~pi715 & ~n17762;
  assign n17764 = ~n17761 & n17763;
  assign n17765 = ~pi647 & ~pi1157;
  assign n17766 = pi647 & pi1157;
  assign n17767 = pi787 & ~n17765;
  assign n17768 = ~n17766 & n17767;
  assign n17769 = n17588 & ~n17768;
  assign n17770 = ~n17576 & ~n17769;
  assign n17771 = ~pi644 & ~n17770;
  assign n17772 = pi644 & n17756;
  assign n17773 = pi715 & ~n17771;
  assign n17774 = ~n17772 & n17773;
  assign n17775 = pi1160 & ~n17764;
  assign n17776 = ~n17774 & n17775;
  assign n17777 = ~pi644 & ~n17760;
  assign n17778 = pi644 & n17576;
  assign n17779 = pi715 & ~n17778;
  assign n17780 = ~n17777 & n17779;
  assign n17781 = ~pi644 & n17756;
  assign n17782 = pi644 & ~n17770;
  assign n17783 = ~pi715 & ~n17782;
  assign n17784 = ~n17781 & n17783;
  assign n17785 = ~pi1160 & ~n17780;
  assign n17786 = ~n17784 & n17785;
  assign n17787 = ~n17776 & ~n17786;
  assign n17788 = pi790 & ~n17787;
  assign n17789 = pi832 & ~n17757;
  assign n17790 = ~n17788 & n17789;
  assign n17791 = pi57 & pi142;
  assign n17792 = ~pi142 & ~n6258;
  assign n17793 = n9829 & ~n16217;
  assign n17794 = pi142 & ~n17793;
  assign n17795 = pi39 & ~n16191;
  assign n17796 = pi142 & ~n17347;
  assign n17797 = ~n17795 & n17796;
  assign n17798 = pi142 & ~n16122;
  assign n17799 = n6221 & ~n17798;
  assign n17800 = pi142 & ~n16104;
  assign n17801 = ~n6221 & ~n17800;
  assign n17802 = pi215 & ~n17799;
  assign n17803 = ~n17801 & n17802;
  assign n17804 = pi142 & n16196;
  assign n17805 = ~n3302 & ~n17804;
  assign n17806 = pi142 & ~n16063;
  assign n17807 = n3302 & ~n17806;
  assign n17808 = ~pi215 & ~n17807;
  assign n17809 = ~n17805 & n17808;
  assign n17810 = ~n17803 & ~n17809;
  assign n17811 = pi39 & pi299;
  assign n17812 = ~n17810 & n17811;
  assign n17813 = ~n17797 & ~n17812;
  assign n17814 = n2576 & ~n17813;
  assign n17815 = ~n17794 & ~n17814;
  assign n17816 = n15753 & ~n17815;
  assign n17817 = pi142 & ~n9829;
  assign n17818 = pi39 & pi142;
  assign n17819 = pi38 & ~n17818;
  assign n17820 = pi142 & ~n16065;
  assign n17821 = n2523 & n17577;
  assign n17822 = ~n17820 & ~n17821;
  assign n17823 = ~pi39 & ~n17822;
  assign n17824 = n17819 & ~n17823;
  assign n17825 = ~pi142 & ~n16353;
  assign n17826 = pi142 & n16368;
  assign n17827 = pi735 & ~n17825;
  assign n17828 = ~n17826 & n17827;
  assign n17829 = pi142 & ~pi735;
  assign n17830 = ~n16057 & n17829;
  assign n17831 = ~n17828 & ~n17830;
  assign n17832 = ~pi39 & ~n17831;
  assign n17833 = ~pi735 & ~n17800;
  assign n17834 = pi142 & ~n16272;
  assign n17835 = ~n16081 & n16294;
  assign n17836 = ~pi142 & n16300;
  assign n17837 = n17835 & n17836;
  assign n17838 = pi735 & ~n17837;
  assign n17839 = ~n17834 & n17838;
  assign n17840 = ~n17833 & ~n17839;
  assign n17841 = ~n6221 & ~n17840;
  assign n17842 = ~pi735 & ~n17798;
  assign n17843 = pi142 & ~n16264;
  assign n17844 = pi735 & ~n17836;
  assign n17845 = ~n17843 & n17844;
  assign n17846 = ~n17842 & ~n17845;
  assign n17847 = n6221 & ~n17846;
  assign n17848 = pi215 & ~n17847;
  assign n17849 = ~n17841 & n17848;
  assign n17850 = pi735 & n16298;
  assign n17851 = n17807 & ~n17850;
  assign n17852 = pi142 & ~n16153;
  assign n17853 = pi735 & n16303;
  assign n17854 = ~n17852 & ~n17853;
  assign n17855 = ~n6221 & ~n17854;
  assign n17856 = pi142 & ~n16251;
  assign n17857 = ~pi142 & ~n16312;
  assign n17858 = ~n17856 & ~n17857;
  assign n17859 = pi735 & ~n17858;
  assign n17860 = pi142 & ~n16184;
  assign n17861 = ~pi735 & ~n17860;
  assign n17862 = ~n17859 & ~n17861;
  assign n17863 = n6221 & n17862;
  assign n17864 = ~n3302 & ~n17855;
  assign n17865 = ~n17863 & n17864;
  assign n17866 = ~pi215 & ~n17851;
  assign n17867 = ~n17865 & n17866;
  assign n17868 = pi299 & ~n17849;
  assign n17869 = ~n17867 & n17868;
  assign n17870 = ~n6194 & ~n17840;
  assign n17871 = n6194 & ~n17846;
  assign n17872 = pi223 & ~n17871;
  assign n17873 = ~n17870 & n17872;
  assign n17874 = n2608 & ~n17806;
  assign n17875 = ~n17850 & n17874;
  assign n17876 = ~n6194 & ~n17854;
  assign n17877 = n6194 & n17862;
  assign n17878 = ~n2608 & ~n17876;
  assign n17879 = ~n17877 & n17878;
  assign n17880 = ~pi223 & ~n17875;
  assign n17881 = ~n17879 & n17880;
  assign n17882 = ~pi299 & ~n17873;
  assign n17883 = ~n17881 & n17882;
  assign n17884 = pi39 & ~n17869;
  assign n17885 = ~n17883 & n17884;
  assign n17886 = ~pi38 & ~n17832;
  assign n17887 = ~n17885 & n17886;
  assign n17888 = n9829 & ~n17824;
  assign n17889 = ~n17887 & n17888;
  assign n17890 = ~n17817 & ~n17889;
  assign n17891 = ~pi778 & ~n17890;
  assign n17892 = ~pi625 & n17890;
  assign n17893 = pi625 & n17815;
  assign n17894 = ~pi1153 & ~n17893;
  assign n17895 = ~n17892 & n17894;
  assign n17896 = ~pi625 & n17815;
  assign n17897 = pi625 & n17890;
  assign n17898 = pi1153 & ~n17896;
  assign n17899 = ~n17897 & n17898;
  assign n17900 = ~n17895 & ~n17899;
  assign n17901 = pi778 & ~n17900;
  assign n17902 = ~n17891 & ~n17901;
  assign n17903 = ~n15741 & ~n17902;
  assign n17904 = n15741 & ~n17815;
  assign n17905 = ~n17903 & ~n17904;
  assign n17906 = ~n15747 & n17905;
  assign n17907 = n15747 & n17815;
  assign n17908 = ~n17906 & ~n17907;
  assign n17909 = ~n15753 & n17908;
  assign n17910 = ~n17816 & ~n17909;
  assign n17911 = ~n15759 & ~n17910;
  assign n17912 = n15759 & ~n17815;
  assign n17913 = ~n17911 & ~n17912;
  assign n17914 = ~pi792 & ~n17913;
  assign n17915 = ~pi628 & ~n17815;
  assign n17916 = pi628 & ~n17913;
  assign n17917 = ~n17915 & ~n17916;
  assign n17918 = pi1156 & ~n17917;
  assign n17919 = ~pi628 & n17913;
  assign n17920 = pi628 & n17815;
  assign n17921 = ~pi1156 & ~n17920;
  assign n17922 = ~n17919 & n17921;
  assign n17923 = ~n17918 & ~n17922;
  assign n17924 = pi792 & ~n17923;
  assign n17925 = ~n17914 & ~n17924;
  assign n17926 = ~pi787 & ~n17925;
  assign n17927 = ~pi647 & n17815;
  assign n17928 = pi647 & n17925;
  assign n17929 = pi1157 & ~n17927;
  assign n17930 = ~n17928 & n17929;
  assign n17931 = ~pi647 & n17925;
  assign n17932 = pi647 & n17815;
  assign n17933 = ~pi1157 & ~n17932;
  assign n17934 = ~n17931 & n17933;
  assign n17935 = ~n17930 & ~n17934;
  assign n17936 = pi787 & ~n17935;
  assign n17937 = ~n17926 & ~n17936;
  assign n17938 = ~pi644 & n17937;
  assign n17939 = ~pi629 & n17918;
  assign n17940 = ~pi619 & n17815;
  assign n17941 = n2523 & n17592;
  assign n17942 = ~n17820 & ~n17941;
  assign n17943 = ~pi39 & ~n17942;
  assign n17944 = n17819 & ~n17943;
  assign n17945 = pi142 & ~pi743;
  assign n17946 = ~n16055 & n17945;
  assign n17947 = ~pi142 & ~n16519;
  assign n17948 = pi142 & ~n16445;
  assign n17949 = pi743 & ~n17947;
  assign n17950 = ~n17948 & n17949;
  assign n17951 = ~pi299 & ~n17946;
  assign n17952 = ~n17950 & n17951;
  assign n17953 = pi142 & n16433;
  assign n17954 = ~pi142 & ~n16524;
  assign n17955 = ~pi743 & n16051;
  assign n17956 = ~n17953 & ~n17955;
  assign n17957 = ~n17954 & n17956;
  assign n17958 = pi299 & ~n17957;
  assign n17959 = ~n17952 & ~n17958;
  assign n17960 = ~pi39 & n17959;
  assign n17961 = pi743 & n16538;
  assign n17962 = ~n17852 & ~n17961;
  assign n17963 = ~n6194 & ~n17962;
  assign n17964 = pi142 & ~n16467;
  assign n17965 = ~pi142 & ~n16544;
  assign n17966 = ~n17964 & ~n17965;
  assign n17967 = pi743 & ~n17966;
  assign n17968 = ~pi743 & ~n17860;
  assign n17969 = ~n17967 & ~n17968;
  assign n17970 = n6194 & n17969;
  assign n17971 = ~n2608 & ~n17963;
  assign n17972 = ~n17970 & n17971;
  assign n17973 = n16062 & n17592;
  assign n17974 = ~n17806 & ~n17973;
  assign n17975 = n2608 & n17974;
  assign n17976 = ~pi223 & ~n17975;
  assign n17977 = ~n17972 & n17976;
  assign n17978 = ~pi743 & ~n17800;
  assign n17979 = pi142 & ~n16493;
  assign n17980 = ~n16533 & ~n16701;
  assign n17981 = pi743 & n17980;
  assign n17982 = ~n17979 & n17981;
  assign n17983 = ~n17978 & ~n17982;
  assign n17984 = ~n6194 & ~n17983;
  assign n17985 = ~pi743 & ~n17798;
  assign n17986 = pi142 & n16484;
  assign n17987 = pi743 & n16534;
  assign n17988 = ~n17986 & n17987;
  assign n17989 = ~n17985 & ~n17988;
  assign n17990 = n6194 & ~n17989;
  assign n17991 = pi223 & ~n17990;
  assign n17992 = ~n17984 & n17991;
  assign n17993 = ~pi299 & ~n17992;
  assign n17994 = ~n17977 & n17993;
  assign n17995 = n6221 & n17969;
  assign n17996 = ~n6221 & ~n17962;
  assign n17997 = ~n3302 & ~n17996;
  assign n17998 = ~n17995 & n17997;
  assign n17999 = n3302 & n17974;
  assign n18000 = ~n17998 & ~n17999;
  assign n18001 = ~pi215 & ~n18000;
  assign n18002 = n6221 & n17989;
  assign n18003 = ~n6221 & n17983;
  assign n18004 = pi215 & ~n18002;
  assign n18005 = ~n18003 & n18004;
  assign n18006 = ~n18001 & ~n18005;
  assign n18007 = pi299 & ~n18006;
  assign n18008 = pi39 & ~n17994;
  assign n18009 = ~n18007 & n18008;
  assign n18010 = ~pi38 & ~n17960;
  assign n18011 = ~n18009 & n18010;
  assign n18012 = n9829 & ~n17944;
  assign n18013 = ~n18011 & n18012;
  assign n18014 = ~n17817 & ~n18013;
  assign n18015 = ~n15777 & ~n18014;
  assign n18016 = n15777 & ~n17815;
  assign n18017 = ~n18015 & ~n18016;
  assign n18018 = ~pi785 & ~n18017;
  assign n18019 = ~n15786 & ~n17815;
  assign n18020 = pi609 & n18015;
  assign n18021 = ~n18019 & ~n18020;
  assign n18022 = pi1155 & ~n18021;
  assign n18023 = ~n16585 & ~n17815;
  assign n18024 = ~pi609 & n18015;
  assign n18025 = ~n18023 & ~n18024;
  assign n18026 = ~pi1155 & ~n18025;
  assign n18027 = ~n18022 & ~n18026;
  assign n18028 = pi785 & ~n18027;
  assign n18029 = ~n18018 & ~n18028;
  assign n18030 = ~pi781 & ~n18029;
  assign n18031 = ~pi618 & n17815;
  assign n18032 = pi618 & n18029;
  assign n18033 = pi1154 & ~n18031;
  assign n18034 = ~n18032 & n18033;
  assign n18035 = ~pi618 & n18029;
  assign n18036 = pi618 & n17815;
  assign n18037 = ~pi1154 & ~n18036;
  assign n18038 = ~n18035 & n18037;
  assign n18039 = ~n18034 & ~n18038;
  assign n18040 = pi781 & ~n18039;
  assign n18041 = ~n18030 & ~n18040;
  assign n18042 = pi619 & n18041;
  assign n18043 = pi1159 & ~n17940;
  assign n18044 = ~n18042 & n18043;
  assign n18045 = pi619 & ~n17908;
  assign n18046 = pi609 & n17902;
  assign n18047 = ~pi625 & n18014;
  assign n18048 = ~pi735 & n17959;
  assign n18049 = pi142 & ~n16366;
  assign n18050 = ~n16524 & n18049;
  assign n18051 = n16433 & ~n16655;
  assign n18052 = n16351 & n18051;
  assign n18053 = ~pi142 & n18052;
  assign n18054 = pi299 & ~n18050;
  assign n18055 = ~n18053 & n18054;
  assign n18056 = pi142 & ~n16361;
  assign n18057 = ~n16519 & n18056;
  assign n18058 = n16345 & ~n16655;
  assign n18059 = ~n16445 & n18058;
  assign n18060 = pi680 & n18059;
  assign n18061 = ~pi142 & n18060;
  assign n18062 = ~pi299 & ~n18057;
  assign n18063 = ~n18061 & n18062;
  assign n18064 = ~n18055 & ~n18063;
  assign n18065 = ~pi743 & ~n18064;
  assign n18066 = n16361 & n17948;
  assign n18067 = ~n16346 & n17947;
  assign n18068 = ~pi299 & ~n18067;
  assign n18069 = ~n18066 & n18068;
  assign n18070 = ~n16351 & n17954;
  assign n18071 = ~n16365 & n17953;
  assign n18072 = pi299 & ~n18070;
  assign n18073 = ~n18071 & n18072;
  assign n18074 = pi743 & ~n18069;
  assign n18075 = ~n18073 & n18074;
  assign n18076 = pi735 & ~n18075;
  assign n18077 = ~n18065 & n18076;
  assign n18078 = ~pi39 & ~n18048;
  assign n18079 = ~n18077 & n18078;
  assign n18080 = pi142 & n16852;
  assign n18081 = ~pi142 & ~n16879;
  assign n18082 = pi743 & ~n18081;
  assign n18083 = ~n18080 & n18082;
  assign n18084 = ~pi142 & ~n16790;
  assign n18085 = pi142 & ~n16728;
  assign n18086 = ~pi743 & ~n18084;
  assign n18087 = ~n18085 & n18086;
  assign n18088 = ~n18083 & ~n18087;
  assign n18089 = pi735 & ~n18088;
  assign n18090 = ~pi735 & ~n17989;
  assign n18091 = ~n18089 & ~n18090;
  assign n18092 = n6194 & ~n18091;
  assign n18093 = pi142 & n16860;
  assign n18094 = ~pi142 & ~n17837;
  assign n18095 = n17980 & n18094;
  assign n18096 = ~n18093 & ~n18095;
  assign n18097 = pi743 & ~n18096;
  assign n18098 = ~pi142 & n16801;
  assign n18099 = pi142 & ~n16712;
  assign n18100 = ~pi743 & ~n18099;
  assign n18101 = ~n18098 & n18100;
  assign n18102 = ~n18097 & ~n18101;
  assign n18103 = pi735 & ~n18102;
  assign n18104 = ~pi735 & ~n17983;
  assign n18105 = ~n18103 & ~n18104;
  assign n18106 = ~n6194 & ~n18105;
  assign n18107 = pi223 & ~n18092;
  assign n18108 = ~n18106 & n18107;
  assign n18109 = ~pi735 & n17974;
  assign n18110 = n2523 & n16921;
  assign n18111 = n17942 & ~n18110;
  assign n18112 = ~n16060 & ~n18111;
  assign n18113 = pi735 & ~n18112;
  assign n18114 = ~n17806 & n18113;
  assign n18115 = ~n18109 & ~n18114;
  assign n18116 = n2608 & ~n18115;
  assign n18117 = ~pi142 & n16892;
  assign n18118 = pi142 & ~n16837;
  assign n18119 = pi743 & ~n18117;
  assign n18120 = ~n18118 & n18119;
  assign n18121 = ~pi142 & ~n16762;
  assign n18122 = pi142 & ~n16695;
  assign n18123 = ~pi743 & ~n18121;
  assign n18124 = ~n18122 & n18123;
  assign n18125 = ~n18120 & ~n18124;
  assign n18126 = pi735 & ~n18125;
  assign n18127 = ~pi735 & ~n17969;
  assign n18128 = ~n18126 & ~n18127;
  assign n18129 = n6194 & n18128;
  assign n18130 = ~pi142 & n16896;
  assign n18131 = pi142 & ~n16843;
  assign n18132 = pi743 & ~n18131;
  assign n18133 = ~n18130 & n18132;
  assign n18134 = ~pi142 & n16781;
  assign n18135 = pi142 & ~n16677;
  assign n18136 = ~pi743 & ~n18135;
  assign n18137 = ~n18134 & n18136;
  assign n18138 = ~n18133 & ~n18137;
  assign n18139 = pi735 & ~n18138;
  assign n18140 = ~pi735 & n17962;
  assign n18141 = ~n18139 & ~n18140;
  assign n18142 = ~n6194 & n18141;
  assign n18143 = ~n2608 & ~n18142;
  assign n18144 = ~n18129 & n18143;
  assign n18145 = ~pi223 & ~n18116;
  assign n18146 = ~n18144 & n18145;
  assign n18147 = ~n18108 & ~n18146;
  assign n18148 = ~pi299 & ~n18147;
  assign n18149 = n6221 & ~n18091;
  assign n18150 = ~n6221 & ~n18105;
  assign n18151 = pi215 & ~n18149;
  assign n18152 = ~n18150 & n18151;
  assign n18153 = n3302 & ~n18115;
  assign n18154 = n6221 & n18128;
  assign n18155 = ~n6221 & n18141;
  assign n18156 = ~n3302 & ~n18155;
  assign n18157 = ~n18154 & n18156;
  assign n18158 = ~pi215 & ~n18153;
  assign n18159 = ~n18157 & n18158;
  assign n18160 = ~n18152 & ~n18159;
  assign n18161 = pi299 & ~n18160;
  assign n18162 = pi39 & ~n18148;
  assign n18163 = ~n18161 & n18162;
  assign n18164 = ~n18079 & ~n18163;
  assign n18165 = ~pi38 & ~n18164;
  assign n18166 = n6081 & n17648;
  assign n18167 = n17944 & ~n18166;
  assign n18168 = n9829 & ~n18167;
  assign n18169 = ~n18165 & n18168;
  assign n18170 = ~n17817 & ~n18169;
  assign n18171 = pi625 & n18170;
  assign n18172 = pi1153 & ~n18047;
  assign n18173 = ~n18171 & n18172;
  assign n18174 = pi608 & ~n17895;
  assign n18175 = ~n18173 & n18174;
  assign n18176 = ~pi625 & n18170;
  assign n18177 = pi625 & n18014;
  assign n18178 = ~pi1153 & ~n18177;
  assign n18179 = ~n18176 & n18178;
  assign n18180 = ~pi608 & ~n17899;
  assign n18181 = ~n18179 & n18180;
  assign n18182 = ~n18175 & ~n18181;
  assign n18183 = pi778 & ~n18182;
  assign n18184 = ~pi778 & n18170;
  assign n18185 = ~n18183 & ~n18184;
  assign n18186 = ~pi609 & ~n18185;
  assign n18187 = ~pi1155 & ~n18046;
  assign n18188 = ~n18186 & n18187;
  assign n18189 = ~pi660 & ~n18022;
  assign n18190 = ~n18188 & n18189;
  assign n18191 = ~pi609 & n17902;
  assign n18192 = pi609 & ~n18185;
  assign n18193 = pi1155 & ~n18191;
  assign n18194 = ~n18192 & n18193;
  assign n18195 = pi660 & ~n18026;
  assign n18196 = ~n18194 & n18195;
  assign n18197 = ~n18190 & ~n18196;
  assign n18198 = pi785 & ~n18197;
  assign n18199 = ~pi785 & ~n18185;
  assign n18200 = ~n18198 & ~n18199;
  assign n18201 = ~pi618 & ~n18200;
  assign n18202 = pi618 & n17905;
  assign n18203 = ~pi1154 & ~n18202;
  assign n18204 = ~n18201 & n18203;
  assign n18205 = ~pi627 & ~n18034;
  assign n18206 = ~n18204 & n18205;
  assign n18207 = ~pi618 & n17905;
  assign n18208 = pi618 & ~n18200;
  assign n18209 = pi1154 & ~n18207;
  assign n18210 = ~n18208 & n18209;
  assign n18211 = pi627 & ~n18038;
  assign n18212 = ~n18210 & n18211;
  assign n18213 = ~n18206 & ~n18212;
  assign n18214 = pi781 & ~n18213;
  assign n18215 = ~pi781 & ~n18200;
  assign n18216 = ~n18214 & ~n18215;
  assign n18217 = ~pi619 & ~n18216;
  assign n18218 = ~pi1159 & ~n18045;
  assign n18219 = ~n18217 & n18218;
  assign n18220 = ~pi648 & ~n18044;
  assign n18221 = ~n18219 & n18220;
  assign n18222 = ~pi619 & n18041;
  assign n18223 = pi619 & n17815;
  assign n18224 = ~pi1159 & ~n18223;
  assign n18225 = ~n18222 & n18224;
  assign n18226 = ~pi619 & ~n17908;
  assign n18227 = pi619 & ~n18216;
  assign n18228 = pi1159 & ~n18226;
  assign n18229 = ~n18227 & n18228;
  assign n18230 = pi648 & ~n18225;
  assign n18231 = ~n18229 & n18230;
  assign n18232 = ~n18221 & ~n18231;
  assign n18233 = pi789 & ~n18232;
  assign n18234 = ~pi789 & ~n18216;
  assign n18235 = ~n18233 & ~n18234;
  assign n18236 = ~pi788 & n18235;
  assign n18237 = ~pi789 & ~n18041;
  assign n18238 = ~n18044 & ~n18225;
  assign n18239 = pi789 & ~n18238;
  assign n18240 = ~n18237 & ~n18239;
  assign n18241 = ~pi626 & n18240;
  assign n18242 = pi626 & n17815;
  assign n18243 = ~pi1158 & ~n18242;
  assign n18244 = ~n18241 & n18243;
  assign n18245 = ~n16995 & ~n18244;
  assign n18246 = ~pi626 & n18235;
  assign n18247 = pi626 & ~n17910;
  assign n18248 = ~pi641 & ~n18247;
  assign n18249 = ~n18246 & n18248;
  assign n18250 = ~n18245 & ~n18249;
  assign n18251 = ~pi626 & n17815;
  assign n18252 = pi626 & n18240;
  assign n18253 = pi1158 & ~n18251;
  assign n18254 = ~n18252 & n18253;
  assign n18255 = ~n17002 & ~n18254;
  assign n18256 = pi626 & n18235;
  assign n18257 = ~pi626 & ~n17910;
  assign n18258 = pi641 & ~n18257;
  assign n18259 = ~n18256 & n18258;
  assign n18260 = ~n18255 & ~n18259;
  assign n18261 = ~n18250 & ~n18260;
  assign n18262 = pi788 & ~n18261;
  assign n18263 = ~n18236 & ~n18262;
  assign n18264 = ~n16643 & ~n18263;
  assign n18265 = ~n18244 & ~n18254;
  assign n18266 = pi788 & ~n18265;
  assign n18267 = ~pi788 & ~n18240;
  assign n18268 = ~n18266 & ~n18267;
  assign n18269 = ~n16633 & ~n18268;
  assign n18270 = pi629 & n17922;
  assign n18271 = ~n17939 & ~n18270;
  assign n18272 = ~n18269 & n18271;
  assign n18273 = ~n18264 & n18272;
  assign n18274 = pi792 & ~n18273;
  assign n18275 = ~pi792 & ~n18263;
  assign n18276 = ~n18274 & ~n18275;
  assign n18277 = ~pi647 & n18276;
  assign n18278 = ~n15925 & n18268;
  assign n18279 = n15925 & n17815;
  assign n18280 = ~n18278 & ~n18279;
  assign n18281 = pi647 & ~n18280;
  assign n18282 = ~pi1157 & ~n18281;
  assign n18283 = ~n18277 & n18282;
  assign n18284 = ~pi630 & ~n17930;
  assign n18285 = ~n18283 & n18284;
  assign n18286 = ~pi647 & ~n18280;
  assign n18287 = pi647 & n18276;
  assign n18288 = pi1157 & ~n18286;
  assign n18289 = ~n18287 & n18288;
  assign n18290 = pi630 & ~n17934;
  assign n18291 = ~n18289 & n18290;
  assign n18292 = ~n18285 & ~n18291;
  assign n18293 = pi787 & ~n18292;
  assign n18294 = ~pi787 & n18276;
  assign n18295 = ~n18293 & ~n18294;
  assign n18296 = pi644 & ~n18295;
  assign n18297 = pi715 & ~n17938;
  assign n18298 = ~n18296 & n18297;
  assign n18299 = ~n15960 & ~n18280;
  assign n18300 = n15960 & n17815;
  assign n18301 = ~n18299 & ~n18300;
  assign n18302 = pi644 & ~n18301;
  assign n18303 = ~pi644 & n17815;
  assign n18304 = ~pi715 & ~n18303;
  assign n18305 = ~n18302 & n18304;
  assign n18306 = pi1160 & ~n18305;
  assign n18307 = ~n18298 & n18306;
  assign n18308 = pi644 & n17937;
  assign n18309 = ~pi715 & ~n18308;
  assign n18310 = ~pi644 & ~n18301;
  assign n18311 = pi644 & n17815;
  assign n18312 = pi715 & ~n18311;
  assign n18313 = ~n18310 & n18312;
  assign n18314 = ~pi1160 & ~n18313;
  assign n18315 = ~n18309 & n18314;
  assign n18316 = ~n18307 & ~n18315;
  assign n18317 = pi790 & ~n18316;
  assign n18318 = ~pi644 & n18314;
  assign n18319 = pi790 & ~n18318;
  assign n18320 = ~n18295 & ~n18319;
  assign n18321 = ~n18317 & ~n18320;
  assign n18322 = n6258 & ~n18321;
  assign n18323 = ~pi57 & ~n17792;
  assign n18324 = ~n18322 & n18323;
  assign n18325 = ~pi832 & ~n17791;
  assign n18326 = ~n18324 & n18325;
  assign po299 = ~n17790 & ~n18326;
  assign n18328 = ~pi143 & ~n2923;
  assign n18329 = ~pi647 & n18328;
  assign n18330 = pi687 & n15726;
  assign n18331 = ~n18328 & ~n18330;
  assign n18332 = ~pi778 & n18331;
  assign n18333 = ~pi625 & n18330;
  assign n18334 = ~n18331 & ~n18333;
  assign n18335 = pi1153 & ~n18334;
  assign n18336 = ~pi1153 & ~n18328;
  assign n18337 = ~n18333 & n18336;
  assign n18338 = ~n18335 & ~n18337;
  assign n18339 = pi778 & ~n18338;
  assign n18340 = ~n18332 & ~n18339;
  assign n18341 = ~n15742 & n18340;
  assign n18342 = ~n15748 & n18341;
  assign n18343 = ~n15754 & n18342;
  assign n18344 = ~n15760 & n18343;
  assign n18345 = ~n15766 & n18344;
  assign n18346 = pi647 & n18345;
  assign n18347 = pi1157 & ~n18329;
  assign n18348 = ~n18346 & n18347;
  assign n18349 = n15772 & n18344;
  assign n18350 = ~pi774 & n15781;
  assign n18351 = ~n18328 & ~n18350;
  assign n18352 = ~n15778 & ~n18351;
  assign n18353 = ~pi785 & ~n18352;
  assign n18354 = ~n15787 & ~n18351;
  assign n18355 = pi1155 & ~n18354;
  assign n18356 = ~n15790 & n18352;
  assign n18357 = ~pi1155 & ~n18356;
  assign n18358 = ~n18355 & ~n18357;
  assign n18359 = pi785 & ~n18358;
  assign n18360 = ~n18353 & ~n18359;
  assign n18361 = ~pi781 & ~n18360;
  assign n18362 = ~n15797 & n18360;
  assign n18363 = pi1154 & ~n18362;
  assign n18364 = ~n15800 & n18360;
  assign n18365 = ~pi1154 & ~n18364;
  assign n18366 = ~n18363 & ~n18365;
  assign n18367 = pi781 & ~n18366;
  assign n18368 = ~n18361 & ~n18367;
  assign n18369 = ~pi789 & ~n18368;
  assign n18370 = ~pi619 & n18328;
  assign n18371 = pi619 & n18368;
  assign n18372 = pi1159 & ~n18370;
  assign n18373 = ~n18371 & n18372;
  assign n18374 = ~pi619 & n18368;
  assign n18375 = pi619 & n18328;
  assign n18376 = ~pi1159 & ~n18375;
  assign n18377 = ~n18374 & n18376;
  assign n18378 = ~n18373 & ~n18377;
  assign n18379 = pi789 & ~n18378;
  assign n18380 = ~n18369 & ~n18379;
  assign n18381 = n15820 & n18380;
  assign n18382 = ~n15820 & n18328;
  assign n18383 = ~n18381 & ~n18382;
  assign n18384 = ~n15758 & ~n18383;
  assign n18385 = n15828 & n18343;
  assign n18386 = ~n18384 & ~n18385;
  assign n18387 = pi788 & ~n18386;
  assign n18388 = pi618 & n18341;
  assign n18389 = pi609 & n18340;
  assign n18390 = ~n15780 & ~n18331;
  assign n18391 = pi625 & n18390;
  assign n18392 = n18351 & ~n18390;
  assign n18393 = ~n18391 & ~n18392;
  assign n18394 = n18336 & ~n18393;
  assign n18395 = ~pi608 & ~n18335;
  assign n18396 = ~n18394 & n18395;
  assign n18397 = pi1153 & n18351;
  assign n18398 = ~n18391 & n18397;
  assign n18399 = pi608 & ~n18337;
  assign n18400 = ~n18398 & n18399;
  assign n18401 = ~n18396 & ~n18400;
  assign n18402 = pi778 & ~n18401;
  assign n18403 = ~pi778 & ~n18392;
  assign n18404 = ~n18402 & ~n18403;
  assign n18405 = ~pi609 & ~n18404;
  assign n18406 = ~pi1155 & ~n18389;
  assign n18407 = ~n18405 & n18406;
  assign n18408 = ~pi660 & ~n18355;
  assign n18409 = ~n18407 & n18408;
  assign n18410 = ~pi609 & n18340;
  assign n18411 = pi609 & ~n18404;
  assign n18412 = pi1155 & ~n18410;
  assign n18413 = ~n18411 & n18412;
  assign n18414 = pi660 & ~n18357;
  assign n18415 = ~n18413 & n18414;
  assign n18416 = ~n18409 & ~n18415;
  assign n18417 = pi785 & ~n18416;
  assign n18418 = ~pi785 & ~n18404;
  assign n18419 = ~n18417 & ~n18418;
  assign n18420 = ~pi618 & ~n18419;
  assign n18421 = ~pi1154 & ~n18388;
  assign n18422 = ~n18420 & n18421;
  assign n18423 = ~pi627 & ~n18363;
  assign n18424 = ~n18422 & n18423;
  assign n18425 = ~pi618 & n18341;
  assign n18426 = pi618 & ~n18419;
  assign n18427 = pi1154 & ~n18425;
  assign n18428 = ~n18426 & n18427;
  assign n18429 = pi627 & ~n18365;
  assign n18430 = ~n18428 & n18429;
  assign n18431 = ~n18424 & ~n18430;
  assign n18432 = pi781 & ~n18431;
  assign n18433 = ~pi781 & ~n18419;
  assign n18434 = ~n18432 & ~n18433;
  assign n18435 = ~pi789 & n18434;
  assign n18436 = ~pi619 & n18342;
  assign n18437 = pi619 & ~n18434;
  assign n18438 = pi1159 & ~n18436;
  assign n18439 = ~n18437 & n18438;
  assign n18440 = pi648 & ~n18377;
  assign n18441 = ~n18439 & n18440;
  assign n18442 = pi619 & n18342;
  assign n18443 = ~pi619 & ~n18434;
  assign n18444 = ~pi1159 & ~n18442;
  assign n18445 = ~n18443 & n18444;
  assign n18446 = ~pi648 & ~n18373;
  assign n18447 = ~n18445 & n18446;
  assign n18448 = pi789 & ~n18441;
  assign n18449 = ~n18447 & n18448;
  assign n18450 = n15833 & ~n18435;
  assign n18451 = ~n18449 & n18450;
  assign n18452 = ~n18387 & ~n18451;
  assign n18453 = ~pi628 & n18452;
  assign n18454 = pi788 & ~n18383;
  assign n18455 = ~pi788 & n18380;
  assign n18456 = ~n18454 & ~n18455;
  assign n18457 = pi628 & n18456;
  assign n18458 = ~pi1156 & ~n18457;
  assign n18459 = ~n18453 & n18458;
  assign n18460 = ~pi629 & ~n18349;
  assign n18461 = ~n18459 & n18460;
  assign n18462 = n15909 & n18344;
  assign n18463 = ~pi628 & n18456;
  assign n18464 = pi628 & n18452;
  assign n18465 = pi1156 & ~n18463;
  assign n18466 = ~n18464 & n18465;
  assign n18467 = pi629 & ~n18462;
  assign n18468 = ~n18466 & n18467;
  assign n18469 = ~n18461 & ~n18468;
  assign n18470 = pi792 & ~n18469;
  assign n18471 = ~pi792 & n18452;
  assign n18472 = ~n18470 & ~n18471;
  assign n18473 = ~pi647 & n18472;
  assign n18474 = n15925 & ~n18328;
  assign n18475 = ~n15925 & n18456;
  assign n18476 = ~n18474 & ~n18475;
  assign n18477 = pi647 & n18476;
  assign n18478 = ~pi1157 & ~n18477;
  assign n18479 = ~n18473 & n18478;
  assign n18480 = ~pi630 & ~n18348;
  assign n18481 = ~n18479 & n18480;
  assign n18482 = ~pi647 & n18345;
  assign n18483 = pi647 & n18328;
  assign n18484 = ~pi1157 & ~n18483;
  assign n18485 = ~n18482 & n18484;
  assign n18486 = ~pi647 & n18476;
  assign n18487 = pi647 & n18472;
  assign n18488 = pi1157 & ~n18486;
  assign n18489 = ~n18487 & n18488;
  assign n18490 = pi630 & ~n18485;
  assign n18491 = ~n18489 & n18490;
  assign n18492 = ~n18481 & ~n18491;
  assign n18493 = pi787 & ~n18492;
  assign n18494 = ~pi787 & n18472;
  assign n18495 = ~n18493 & ~n18494;
  assign n18496 = ~pi790 & ~n18495;
  assign n18497 = ~pi787 & ~n18345;
  assign n18498 = ~n18348 & ~n18485;
  assign n18499 = pi787 & ~n18498;
  assign n18500 = ~n18497 & ~n18499;
  assign n18501 = ~pi644 & n18500;
  assign n18502 = pi644 & ~n18495;
  assign n18503 = pi715 & ~n18501;
  assign n18504 = ~n18502 & n18503;
  assign n18505 = ~n15960 & n18476;
  assign n18506 = n15960 & n18328;
  assign n18507 = ~n18505 & ~n18506;
  assign n18508 = pi644 & ~n18507;
  assign n18509 = ~pi644 & n18328;
  assign n18510 = ~pi715 & ~n18509;
  assign n18511 = ~n18508 & n18510;
  assign n18512 = pi1160 & ~n18511;
  assign n18513 = ~n18504 & n18512;
  assign n18514 = ~pi644 & ~n18507;
  assign n18515 = pi644 & n18328;
  assign n18516 = pi715 & ~n18515;
  assign n18517 = ~n18514 & n18516;
  assign n18518 = pi644 & n18500;
  assign n18519 = ~pi644 & ~n18495;
  assign n18520 = ~pi715 & ~n18518;
  assign n18521 = ~n18519 & n18520;
  assign n18522 = ~pi1160 & ~n18517;
  assign n18523 = ~n18521 & n18522;
  assign n18524 = ~n18513 & ~n18523;
  assign n18525 = pi790 & ~n18524;
  assign n18526 = pi832 & ~n18496;
  assign n18527 = ~n18525 & n18526;
  assign n18528 = ~pi143 & po1038;
  assign n18529 = ~pi143 & ~n16219;
  assign n18530 = n15759 & ~n18529;
  assign n18531 = n15747 & ~n18529;
  assign n18532 = pi143 & ~n9829;
  assign n18533 = ~pi143 & ~n16218;
  assign n18534 = ~pi687 & n18533;
  assign n18535 = ~pi143 & ~n16228;
  assign n18536 = n16227 & ~n18535;
  assign n18537 = pi143 & n17272;
  assign n18538 = ~pi143 & ~n17276;
  assign n18539 = ~pi38 & ~n18537;
  assign n18540 = ~n18538 & n18539;
  assign n18541 = pi687 & ~n18536;
  assign n18542 = ~n18540 & n18541;
  assign n18543 = n9829 & ~n18542;
  assign n18544 = ~n18534 & n18543;
  assign n18545 = ~n18532 & ~n18544;
  assign n18546 = ~pi778 & ~n18545;
  assign n18547 = ~pi625 & n18529;
  assign n18548 = pi625 & n18545;
  assign n18549 = pi1153 & ~n18547;
  assign n18550 = ~n18548 & n18549;
  assign n18551 = ~pi625 & n18545;
  assign n18552 = pi625 & n18529;
  assign n18553 = ~pi1153 & ~n18552;
  assign n18554 = ~n18551 & n18553;
  assign n18555 = ~n18550 & ~n18554;
  assign n18556 = pi778 & ~n18555;
  assign n18557 = ~n18546 & ~n18556;
  assign n18558 = ~n15741 & n18557;
  assign n18559 = n15741 & n18529;
  assign n18560 = ~n18558 & ~n18559;
  assign n18561 = ~n15747 & n18560;
  assign n18562 = ~n18531 & ~n18561;
  assign n18563 = ~n15753 & n18562;
  assign n18564 = n15753 & n18529;
  assign n18565 = ~n18563 & ~n18564;
  assign n18566 = ~n15759 & n18565;
  assign n18567 = ~n18530 & ~n18566;
  assign n18568 = ~pi792 & ~n18567;
  assign n18569 = ~pi628 & ~n18529;
  assign n18570 = pi628 & ~n18567;
  assign n18571 = ~n18569 & ~n18570;
  assign n18572 = pi1156 & ~n18571;
  assign n18573 = ~pi628 & n18567;
  assign n18574 = pi628 & n18529;
  assign n18575 = ~pi1156 & ~n18574;
  assign n18576 = ~n18573 & n18575;
  assign n18577 = ~n18572 & ~n18576;
  assign n18578 = pi792 & ~n18577;
  assign n18579 = ~n18568 & ~n18578;
  assign n18580 = ~pi787 & ~n18579;
  assign n18581 = ~pi647 & n18529;
  assign n18582 = pi647 & n18579;
  assign n18583 = pi1157 & ~n18581;
  assign n18584 = ~n18582 & n18583;
  assign n18585 = ~pi647 & n18579;
  assign n18586 = pi647 & n18529;
  assign n18587 = ~pi1157 & ~n18586;
  assign n18588 = ~n18585 & n18587;
  assign n18589 = ~n18584 & ~n18588;
  assign n18590 = pi787 & ~n18589;
  assign n18591 = ~n18580 & ~n18590;
  assign n18592 = ~pi644 & n18591;
  assign n18593 = ~pi629 & n18572;
  assign n18594 = ~pi619 & n18529;
  assign n18595 = pi774 & ~n18533;
  assign n18596 = pi38 & ~pi39;
  assign n18597 = n15781 & n18596;
  assign n18598 = n2513 & n18597;
  assign n18599 = ~pi38 & n16565;
  assign n18600 = pi143 & ~n18599;
  assign n18601 = ~pi38 & ~n16514;
  assign n18602 = n6081 & n16486;
  assign n18603 = pi38 & ~n18602;
  assign n18604 = ~n18601 & ~n18603;
  assign n18605 = ~pi143 & ~pi774;
  assign n18606 = n18604 & n18605;
  assign n18607 = ~n18600 & ~n18606;
  assign n18608 = ~n18598 & ~n18607;
  assign n18609 = ~n18595 & ~n18608;
  assign n18610 = n9829 & ~n18609;
  assign n18611 = ~n18532 & ~n18610;
  assign n18612 = ~n15777 & ~n18611;
  assign n18613 = n15777 & ~n18529;
  assign n18614 = ~n18612 & ~n18613;
  assign n18615 = ~pi785 & ~n18614;
  assign n18616 = ~n15786 & ~n18529;
  assign n18617 = pi609 & n18612;
  assign n18618 = ~n18616 & ~n18617;
  assign n18619 = pi1155 & ~n18618;
  assign n18620 = ~n16585 & ~n18529;
  assign n18621 = ~pi609 & n18612;
  assign n18622 = ~n18620 & ~n18621;
  assign n18623 = ~pi1155 & ~n18622;
  assign n18624 = ~n18619 & ~n18623;
  assign n18625 = pi785 & ~n18624;
  assign n18626 = ~n18615 & ~n18625;
  assign n18627 = ~pi781 & ~n18626;
  assign n18628 = ~pi618 & n18529;
  assign n18629 = pi618 & n18626;
  assign n18630 = pi1154 & ~n18628;
  assign n18631 = ~n18629 & n18630;
  assign n18632 = ~pi618 & n18626;
  assign n18633 = pi618 & n18529;
  assign n18634 = ~pi1154 & ~n18633;
  assign n18635 = ~n18632 & n18634;
  assign n18636 = ~n18631 & ~n18635;
  assign n18637 = pi781 & ~n18636;
  assign n18638 = ~n18627 & ~n18637;
  assign n18639 = pi619 & n18638;
  assign n18640 = pi1159 & ~n18594;
  assign n18641 = ~n18639 & n18640;
  assign n18642 = pi618 & ~n18560;
  assign n18643 = pi609 & n18557;
  assign n18644 = ~pi687 & n18609;
  assign n18645 = ~pi39 & ~n16647;
  assign n18646 = ~pi38 & n18645;
  assign n18647 = pi39 & n16877;
  assign n18648 = ~pi39 & n16808;
  assign n18649 = pi38 & ~n18648;
  assign n18650 = ~n18646 & ~n18649;
  assign n18651 = ~n18647 & n18650;
  assign n18652 = ~pi143 & ~n18651;
  assign n18653 = n16228 & ~n16807;
  assign n18654 = pi38 & ~n18653;
  assign n18655 = pi39 & ~n16913;
  assign n18656 = ~n16526 & n17270;
  assign n18657 = ~n18655 & ~n18656;
  assign n18658 = ~pi38 & ~n18657;
  assign n18659 = ~n18654 & ~n18658;
  assign n18660 = pi143 & n18659;
  assign n18661 = ~pi774 & ~n18652;
  assign n18662 = ~n18660 & n18661;
  assign n18663 = pi39 & ~n16825;
  assign n18664 = ~pi39 & ~n16657;
  assign n18665 = ~n18663 & ~n18664;
  assign n18666 = ~pi38 & n18665;
  assign n18667 = pi143 & n18666;
  assign n18668 = n18110 & n18596;
  assign n18669 = n16228 & ~n16664;
  assign n18670 = pi38 & n18669;
  assign n18671 = pi39 & ~n16747;
  assign n18672 = ~pi39 & n16653;
  assign n18673 = ~n18671 & ~n18672;
  assign n18674 = ~pi38 & n18673;
  assign n18675 = ~n18670 & ~n18674;
  assign n18676 = ~pi143 & n18675;
  assign n18677 = pi774 & ~n18668;
  assign n18678 = ~n18667 & n18677;
  assign n18679 = ~n18676 & n18678;
  assign n18680 = pi687 & ~n18662;
  assign n18681 = ~n18679 & n18680;
  assign n18682 = n9829 & ~n18681;
  assign n18683 = ~n18644 & n18682;
  assign n18684 = ~n18532 & ~n18683;
  assign n18685 = ~pi625 & n18684;
  assign n18686 = pi625 & n18611;
  assign n18687 = ~pi1153 & ~n18686;
  assign n18688 = ~n18685 & n18687;
  assign n18689 = ~pi608 & ~n18550;
  assign n18690 = ~n18688 & n18689;
  assign n18691 = ~pi625 & n18611;
  assign n18692 = pi625 & n18684;
  assign n18693 = pi1153 & ~n18691;
  assign n18694 = ~n18692 & n18693;
  assign n18695 = pi608 & ~n18554;
  assign n18696 = ~n18694 & n18695;
  assign n18697 = ~n18690 & ~n18696;
  assign n18698 = pi778 & ~n18697;
  assign n18699 = ~pi778 & n18684;
  assign n18700 = ~n18698 & ~n18699;
  assign n18701 = ~pi609 & ~n18700;
  assign n18702 = ~pi1155 & ~n18643;
  assign n18703 = ~n18701 & n18702;
  assign n18704 = ~pi660 & ~n18619;
  assign n18705 = ~n18703 & n18704;
  assign n18706 = ~pi609 & n18557;
  assign n18707 = pi609 & ~n18700;
  assign n18708 = pi1155 & ~n18706;
  assign n18709 = ~n18707 & n18708;
  assign n18710 = pi660 & ~n18623;
  assign n18711 = ~n18709 & n18710;
  assign n18712 = ~n18705 & ~n18711;
  assign n18713 = pi785 & ~n18712;
  assign n18714 = ~pi785 & ~n18700;
  assign n18715 = ~n18713 & ~n18714;
  assign n18716 = ~pi618 & ~n18715;
  assign n18717 = ~pi1154 & ~n18642;
  assign n18718 = ~n18716 & n18717;
  assign n18719 = ~pi627 & ~n18631;
  assign n18720 = ~n18718 & n18719;
  assign n18721 = ~pi618 & ~n18560;
  assign n18722 = pi618 & ~n18715;
  assign n18723 = pi1154 & ~n18721;
  assign n18724 = ~n18722 & n18723;
  assign n18725 = pi627 & ~n18635;
  assign n18726 = ~n18724 & n18725;
  assign n18727 = ~n18720 & ~n18726;
  assign n18728 = pi781 & ~n18727;
  assign n18729 = ~pi781 & ~n18715;
  assign n18730 = ~n18728 & ~n18729;
  assign n18731 = ~pi619 & ~n18730;
  assign n18732 = pi619 & n18562;
  assign n18733 = ~pi1159 & ~n18732;
  assign n18734 = ~n18731 & n18733;
  assign n18735 = ~pi648 & ~n18641;
  assign n18736 = ~n18734 & n18735;
  assign n18737 = ~pi619 & n18638;
  assign n18738 = pi619 & n18529;
  assign n18739 = ~pi1159 & ~n18738;
  assign n18740 = ~n18737 & n18739;
  assign n18741 = ~pi619 & n18562;
  assign n18742 = pi619 & ~n18730;
  assign n18743 = pi1159 & ~n18741;
  assign n18744 = ~n18742 & n18743;
  assign n18745 = pi648 & ~n18740;
  assign n18746 = ~n18744 & n18745;
  assign n18747 = ~n18736 & ~n18746;
  assign n18748 = pi789 & ~n18747;
  assign n18749 = ~pi789 & ~n18730;
  assign n18750 = ~n18748 & ~n18749;
  assign n18751 = ~pi788 & n18750;
  assign n18752 = ~pi789 & ~n18638;
  assign n18753 = ~n18641 & ~n18740;
  assign n18754 = pi789 & ~n18753;
  assign n18755 = ~n18752 & ~n18754;
  assign n18756 = ~pi626 & n18755;
  assign n18757 = pi626 & n18529;
  assign n18758 = ~pi1158 & ~n18757;
  assign n18759 = ~n18756 & n18758;
  assign n18760 = ~n16995 & ~n18759;
  assign n18761 = ~pi626 & n18750;
  assign n18762 = pi626 & n18565;
  assign n18763 = ~pi641 & ~n18762;
  assign n18764 = ~n18761 & n18763;
  assign n18765 = ~n18760 & ~n18764;
  assign n18766 = ~pi626 & n18529;
  assign n18767 = pi626 & n18755;
  assign n18768 = pi1158 & ~n18766;
  assign n18769 = ~n18767 & n18768;
  assign n18770 = ~n17002 & ~n18769;
  assign n18771 = ~pi626 & n18565;
  assign n18772 = pi626 & n18750;
  assign n18773 = pi641 & ~n18771;
  assign n18774 = ~n18772 & n18773;
  assign n18775 = ~n18770 & ~n18774;
  assign n18776 = ~n18765 & ~n18775;
  assign n18777 = pi788 & ~n18776;
  assign n18778 = ~n18751 & ~n18777;
  assign n18779 = ~n16643 & ~n18778;
  assign n18780 = ~n18759 & ~n18769;
  assign n18781 = pi788 & ~n18780;
  assign n18782 = ~pi788 & ~n18755;
  assign n18783 = ~n18781 & ~n18782;
  assign n18784 = ~n16633 & ~n18783;
  assign n18785 = pi629 & n18576;
  assign n18786 = ~n18593 & ~n18785;
  assign n18787 = ~n18784 & n18786;
  assign n18788 = ~n18779 & n18787;
  assign n18789 = pi792 & ~n18788;
  assign n18790 = ~pi792 & ~n18778;
  assign n18791 = ~n18789 & ~n18790;
  assign n18792 = ~pi647 & n18791;
  assign n18793 = ~n15925 & n18783;
  assign n18794 = n15925 & n18529;
  assign n18795 = ~n18793 & ~n18794;
  assign n18796 = pi647 & ~n18795;
  assign n18797 = ~pi1157 & ~n18796;
  assign n18798 = ~n18792 & n18797;
  assign n18799 = ~pi630 & ~n18584;
  assign n18800 = ~n18798 & n18799;
  assign n18801 = ~pi647 & ~n18795;
  assign n18802 = pi647 & n18791;
  assign n18803 = pi1157 & ~n18801;
  assign n18804 = ~n18802 & n18803;
  assign n18805 = pi630 & ~n18588;
  assign n18806 = ~n18804 & n18805;
  assign n18807 = ~n18800 & ~n18806;
  assign n18808 = pi787 & ~n18807;
  assign n18809 = ~pi787 & n18791;
  assign n18810 = ~n18808 & ~n18809;
  assign n18811 = pi644 & ~n18810;
  assign n18812 = pi715 & ~n18592;
  assign n18813 = ~n18811 & n18812;
  assign n18814 = ~n15960 & ~n18795;
  assign n18815 = n15960 & n18529;
  assign n18816 = ~n18814 & ~n18815;
  assign n18817 = pi644 & ~n18816;
  assign n18818 = ~pi644 & n18529;
  assign n18819 = ~pi715 & ~n18818;
  assign n18820 = ~n18817 & n18819;
  assign n18821 = pi1160 & ~n18820;
  assign n18822 = ~n18813 & n18821;
  assign n18823 = pi644 & n18591;
  assign n18824 = ~pi715 & ~n18823;
  assign n18825 = ~pi644 & ~n18816;
  assign n18826 = pi644 & n18529;
  assign n18827 = pi715 & ~n18826;
  assign n18828 = ~n18825 & n18827;
  assign n18829 = ~pi1160 & ~n18828;
  assign n18830 = ~n18824 & n18829;
  assign n18831 = ~n18822 & ~n18830;
  assign n18832 = pi790 & ~n18831;
  assign n18833 = ~pi644 & n18829;
  assign n18834 = pi790 & ~n18833;
  assign n18835 = ~n18810 & ~n18834;
  assign n18836 = ~n18832 & ~n18835;
  assign n18837 = ~po1038 & ~n18836;
  assign n18838 = ~pi832 & ~n18528;
  assign n18839 = ~n18837 & n18838;
  assign po300 = ~n18527 & ~n18839;
  assign n18841 = ~n15960 & ~n17768;
  assign n18842 = pi144 & ~n2923;
  assign n18843 = pi736 & n15726;
  assign n18844 = ~n18842 & ~n18843;
  assign n18845 = ~pi778 & n18844;
  assign n18846 = pi625 & n18843;
  assign n18847 = ~n18844 & ~n18846;
  assign n18848 = ~pi1153 & ~n18847;
  assign n18849 = pi1153 & ~n18842;
  assign n18850 = ~n18846 & n18849;
  assign n18851 = ~n18848 & ~n18850;
  assign n18852 = pi778 & ~n18851;
  assign n18853 = ~n18845 & ~n18852;
  assign n18854 = n17584 & n18853;
  assign n18855 = n17585 & n18854;
  assign n18856 = ~pi628 & n18855;
  assign n18857 = pi629 & ~n18856;
  assign n18858 = ~pi609 & ~pi1155;
  assign n18859 = pi609 & pi1155;
  assign n18860 = pi785 & ~n18858;
  assign n18861 = ~n18859 & n18860;
  assign n18862 = ~pi619 & pi1159;
  assign n18863 = pi619 & ~pi1159;
  assign n18864 = ~n18862 & ~n18863;
  assign n18865 = pi789 & ~n18864;
  assign n18866 = ~pi618 & ~pi1154;
  assign n18867 = pi618 & pi1154;
  assign n18868 = pi781 & ~n18866;
  assign n18869 = ~n18867 & n18868;
  assign n18870 = ~n15777 & ~n18861;
  assign n18871 = ~n18865 & ~n18869;
  assign n18872 = n18870 & n18871;
  assign n18873 = pi758 & n15781;
  assign n18874 = n18872 & n18873;
  assign n18875 = ~n15832 & n18874;
  assign n18876 = pi628 & ~n18875;
  assign n18877 = ~n18857 & ~n18876;
  assign n18878 = ~pi1156 & ~n18877;
  assign n18879 = pi628 & n18855;
  assign n18880 = ~pi628 & ~n18875;
  assign n18881 = pi629 & ~n18880;
  assign n18882 = pi1156 & ~n18881;
  assign n18883 = ~n18879 & n18882;
  assign n18884 = ~n18878 & ~n18883;
  assign n18885 = ~n18842 & ~n18884;
  assign n18886 = pi792 & n18885;
  assign n18887 = pi618 & ~pi627;
  assign n18888 = ~pi1154 & n18887;
  assign n18889 = ~pi618 & pi627;
  assign n18890 = pi1154 & n18889;
  assign n18891 = ~n18888 & ~n18890;
  assign n18892 = pi781 & ~n18891;
  assign n18893 = ~n15747 & ~n18892;
  assign n18894 = ~n18842 & ~n18873;
  assign n18895 = ~n15780 & n18843;
  assign n18896 = n18894 & ~n18895;
  assign n18897 = pi625 & n18895;
  assign n18898 = ~n18896 & ~n18897;
  assign n18899 = ~pi1153 & ~n18898;
  assign n18900 = ~pi608 & ~n18850;
  assign n18901 = ~n18899 & n18900;
  assign n18902 = pi1153 & n18894;
  assign n18903 = ~n18897 & n18902;
  assign n18904 = pi608 & ~n18848;
  assign n18905 = ~n18903 & n18904;
  assign n18906 = ~n18901 & ~n18905;
  assign n18907 = pi778 & ~n18906;
  assign n18908 = ~pi778 & ~n18896;
  assign n18909 = ~n18907 & ~n18908;
  assign n18910 = pi660 & n18859;
  assign n18911 = pi785 & ~n18910;
  assign n18912 = n18909 & ~n18911;
  assign n18913 = ~n15787 & ~n18894;
  assign n18914 = pi1155 & ~n18913;
  assign n18915 = ~pi609 & ~n18909;
  assign n18916 = pi609 & n18853;
  assign n18917 = ~pi1155 & ~n18916;
  assign n18918 = ~n18915 & n18917;
  assign n18919 = ~pi660 & ~n18914;
  assign n18920 = ~n18918 & n18919;
  assign n18921 = n16585 & n18873;
  assign n18922 = ~pi1155 & ~n18842;
  assign n18923 = ~n18921 & n18922;
  assign n18924 = ~pi609 & pi1155;
  assign n18925 = ~n18853 & n18924;
  assign n18926 = pi660 & ~n18923;
  assign n18927 = ~n18925 & n18926;
  assign n18928 = pi785 & ~n18927;
  assign n18929 = ~n18920 & n18928;
  assign n18930 = ~n18912 & ~n18929;
  assign n18931 = n18893 & ~n18930;
  assign n18932 = ~n18861 & n18873;
  assign n18933 = ~n18869 & n18932;
  assign n18934 = ~pi619 & ~n15777;
  assign n18935 = n18933 & n18934;
  assign n18936 = n15751 & ~n18842;
  assign n18937 = ~n18935 & n18936;
  assign n18938 = pi619 & ~n15777;
  assign n18939 = n18933 & n18938;
  assign n18940 = n15750 & ~n18842;
  assign n18941 = ~n18939 & n18940;
  assign n18942 = pi648 & n18862;
  assign n18943 = ~pi648 & n18863;
  assign n18944 = ~n18942 & ~n18943;
  assign n18945 = ~n18842 & ~n18944;
  assign n18946 = ~n18854 & n18945;
  assign n18947 = ~n18937 & ~n18941;
  assign n18948 = ~n18946 & n18947;
  assign n18949 = pi789 & ~n18948;
  assign n18950 = pi618 & ~n15777;
  assign n18951 = n15745 & ~n18950;
  assign n18952 = ~n15741 & n18853;
  assign n18953 = ~n18891 & ~n18952;
  assign n18954 = ~n15746 & ~n18932;
  assign n18955 = ~pi618 & ~n15777;
  assign n18956 = n15744 & ~n18955;
  assign n18957 = ~n18951 & ~n18956;
  assign n18958 = ~n18954 & n18957;
  assign n18959 = ~n18953 & n18958;
  assign n18960 = pi781 & ~n18842;
  assign n18961 = ~n18959 & n18960;
  assign n18962 = ~n18949 & ~n18961;
  assign n18963 = ~n18931 & n18962;
  assign n18964 = ~pi619 & ~pi1159;
  assign n18965 = ~pi648 & n18964;
  assign n18966 = pi619 & pi1159;
  assign n18967 = pi648 & n18966;
  assign n18968 = ~n18965 & ~n18967;
  assign n18969 = pi789 & n18968;
  assign n18970 = n18948 & n18969;
  assign n18971 = ~n18963 & ~n18970;
  assign n18972 = n15833 & ~n18971;
  assign n18973 = ~n15753 & n18854;
  assign n18974 = ~n18842 & ~n18973;
  assign n18975 = n15818 & ~n18974;
  assign n18976 = ~pi626 & n18874;
  assign n18977 = ~n18842 & ~n18976;
  assign n18978 = ~pi1158 & ~n18977;
  assign n18979 = pi641 & ~n18978;
  assign n18980 = ~n18975 & n18979;
  assign n18981 = pi626 & n18874;
  assign n18982 = ~n18842 & ~n18981;
  assign n18983 = pi1158 & ~n18982;
  assign n18984 = n15819 & ~n18974;
  assign n18985 = ~pi641 & ~n18983;
  assign n18986 = ~n18984 & n18985;
  assign n18987 = pi788 & ~n18980;
  assign n18988 = ~n18986 & n18987;
  assign n18989 = ~n18972 & ~n18988;
  assign n18990 = ~n18886 & ~n18989;
  assign n18991 = n16644 & ~n18885;
  assign n18992 = n18841 & ~n18991;
  assign n18993 = ~n18990 & n18992;
  assign n18994 = ~n15925 & n18875;
  assign n18995 = pi630 & n18994;
  assign n18996 = ~n15765 & n18855;
  assign n18997 = ~pi630 & ~n18996;
  assign n18998 = pi647 & ~n18997;
  assign n18999 = pi1157 & ~n18995;
  assign n19000 = ~n18998 & n18999;
  assign n19001 = ~pi630 & n18994;
  assign n19002 = pi630 & ~n18996;
  assign n19003 = ~pi647 & ~n19002;
  assign n19004 = ~pi1157 & ~n19001;
  assign n19005 = ~n19003 & n19004;
  assign n19006 = ~n19000 & ~n19005;
  assign n19007 = pi787 & ~n18842;
  assign n19008 = ~n19006 & n19007;
  assign n19009 = ~n18993 & ~n19008;
  assign n19010 = ~pi790 & n19009;
  assign n19011 = ~n17768 & n18996;
  assign n19012 = ~n18842 & ~n19011;
  assign n19013 = ~pi644 & ~n19012;
  assign n19014 = pi644 & n19009;
  assign n19015 = pi715 & ~n19013;
  assign n19016 = ~n19014 & n19015;
  assign n19017 = ~n15960 & n18994;
  assign n19018 = pi644 & n19017;
  assign n19019 = ~pi715 & ~n18842;
  assign n19020 = ~n19018 & n19019;
  assign n19021 = pi1160 & ~n19020;
  assign n19022 = ~n19016 & n19021;
  assign n19023 = ~pi644 & n19017;
  assign n19024 = pi715 & ~n18842;
  assign n19025 = ~n19023 & n19024;
  assign n19026 = ~pi644 & n19009;
  assign n19027 = pi644 & ~n19012;
  assign n19028 = ~pi715 & ~n19027;
  assign n19029 = ~n19026 & n19028;
  assign n19030 = ~pi1160 & ~n19025;
  assign n19031 = ~n19029 & n19030;
  assign n19032 = ~n19022 & ~n19031;
  assign n19033 = pi790 & ~n19032;
  assign n19034 = pi832 & ~n19010;
  assign n19035 = ~n19033 & n19034;
  assign n19036 = pi57 & pi144;
  assign n19037 = ~pi144 & ~n6258;
  assign n19038 = pi144 & ~n16219;
  assign n19039 = n15759 & ~n19038;
  assign n19040 = n15747 & ~n19038;
  assign n19041 = pi736 & n9829;
  assign n19042 = ~n19038 & ~n19041;
  assign n19043 = ~pi144 & ~n17272;
  assign n19044 = pi144 & n17276;
  assign n19045 = ~pi38 & ~n19043;
  assign n19046 = ~n19044 & n19045;
  assign n19047 = ~pi144 & ~n16228;
  assign n19048 = ~n15725 & n16228;
  assign n19049 = pi38 & ~n19048;
  assign n19050 = ~n19047 & n19049;
  assign n19051 = n19041 & ~n19050;
  assign n19052 = ~n19046 & n19051;
  assign n19053 = ~n19042 & ~n19052;
  assign n19054 = ~pi778 & n19053;
  assign n19055 = ~pi625 & ~n19038;
  assign n19056 = pi625 & ~n19053;
  assign n19057 = pi1153 & ~n19055;
  assign n19058 = ~n19056 & n19057;
  assign n19059 = ~pi625 & ~n19053;
  assign n19060 = pi625 & ~n19038;
  assign n19061 = ~pi1153 & ~n19060;
  assign n19062 = ~n19059 & n19061;
  assign n19063 = ~n19058 & ~n19062;
  assign n19064 = pi778 & ~n19063;
  assign n19065 = ~n19054 & ~n19064;
  assign n19066 = ~n15741 & ~n19065;
  assign n19067 = n15741 & n19038;
  assign n19068 = ~n19066 & ~n19067;
  assign n19069 = ~n15747 & n19068;
  assign n19070 = ~n19040 & ~n19069;
  assign n19071 = ~n15753 & n19070;
  assign n19072 = n15753 & n19038;
  assign n19073 = ~n19071 & ~n19072;
  assign n19074 = ~n15759 & n19073;
  assign n19075 = ~n19039 & ~n19074;
  assign n19076 = ~pi792 & n19075;
  assign n19077 = pi628 & n19075;
  assign n19078 = ~pi628 & n19038;
  assign n19079 = ~n19077 & ~n19078;
  assign n19080 = pi1156 & ~n19079;
  assign n19081 = pi628 & ~n19038;
  assign n19082 = ~pi628 & ~n19075;
  assign n19083 = ~pi1156 & ~n19081;
  assign n19084 = ~n19082 & n19083;
  assign n19085 = ~n19080 & ~n19084;
  assign n19086 = pi792 & ~n19085;
  assign n19087 = ~n19076 & ~n19086;
  assign n19088 = ~pi787 & ~n19087;
  assign n19089 = ~pi647 & ~n19038;
  assign n19090 = pi647 & n19087;
  assign n19091 = pi1157 & ~n19089;
  assign n19092 = ~n19090 & n19091;
  assign n19093 = pi647 & ~n19038;
  assign n19094 = ~pi647 & n19087;
  assign n19095 = ~pi1157 & ~n19093;
  assign n19096 = ~n19094 & n19095;
  assign n19097 = ~n19092 & ~n19096;
  assign n19098 = pi787 & ~n19097;
  assign n19099 = ~n19088 & ~n19098;
  assign n19100 = ~pi644 & n19099;
  assign n19101 = ~pi629 & n19080;
  assign n19102 = ~pi619 & ~n19038;
  assign n19103 = pi144 & ~n9829;
  assign n19104 = ~pi758 & ~n16212;
  assign n19105 = pi758 & ~n16512;
  assign n19106 = ~n19104 & ~n19105;
  assign n19107 = pi39 & ~n19106;
  assign n19108 = ~pi758 & n16057;
  assign n19109 = n16448 & ~n19108;
  assign n19110 = ~n19107 & ~n19109;
  assign n19111 = pi144 & ~n19110;
  assign n19112 = ~pi144 & pi758;
  assign n19113 = n16565 & n19112;
  assign n19114 = ~n19111 & ~n19113;
  assign n19115 = ~pi38 & ~n19114;
  assign n19116 = pi758 & n15780;
  assign n19117 = n16228 & ~n19116;
  assign n19118 = pi38 & ~n19047;
  assign n19119 = ~n19117 & n19118;
  assign n19120 = ~n19115 & ~n19119;
  assign n19121 = n9829 & ~n19120;
  assign n19122 = ~n19103 & ~n19121;
  assign n19123 = ~n15777 & ~n19122;
  assign n19124 = n15777 & n19038;
  assign n19125 = ~n19123 & ~n19124;
  assign n19126 = ~pi785 & ~n19125;
  assign n19127 = pi609 & n19125;
  assign n19128 = ~pi609 & ~n19038;
  assign n19129 = pi1155 & ~n19128;
  assign n19130 = ~n19127 & n19129;
  assign n19131 = ~pi609 & n19125;
  assign n19132 = pi609 & ~n19038;
  assign n19133 = ~pi1155 & ~n19132;
  assign n19134 = ~n19131 & n19133;
  assign n19135 = ~n19130 & ~n19134;
  assign n19136 = pi785 & ~n19135;
  assign n19137 = ~n19126 & ~n19136;
  assign n19138 = ~pi781 & ~n19137;
  assign n19139 = ~pi618 & ~n19038;
  assign n19140 = pi618 & n19137;
  assign n19141 = pi1154 & ~n19139;
  assign n19142 = ~n19140 & n19141;
  assign n19143 = pi618 & ~n19038;
  assign n19144 = ~pi618 & n19137;
  assign n19145 = ~pi1154 & ~n19143;
  assign n19146 = ~n19144 & n19145;
  assign n19147 = ~n19142 & ~n19146;
  assign n19148 = pi781 & ~n19147;
  assign n19149 = ~n19138 & ~n19148;
  assign n19150 = pi619 & n19149;
  assign n19151 = pi1159 & ~n19102;
  assign n19152 = ~n19150 & n19151;
  assign n19153 = pi619 & ~n19070;
  assign n19154 = pi609 & n19065;
  assign n19155 = ~n19041 & ~n19121;
  assign n19156 = ~pi144 & ~n16657;
  assign n19157 = pi144 & ~n16653;
  assign n19158 = ~pi758 & ~n19156;
  assign n19159 = ~n19157 & n19158;
  assign n19160 = ~pi144 & n17397;
  assign n19161 = pi144 & n16647;
  assign n19162 = pi758 & ~n19160;
  assign n19163 = ~n19161 & n19162;
  assign n19164 = ~pi39 & ~n19163;
  assign n19165 = ~n19159 & n19164;
  assign n19166 = pi144 & ~n16877;
  assign n19167 = ~pi144 & ~n16913;
  assign n19168 = pi758 & ~n19166;
  assign n19169 = ~n19167 & n19168;
  assign n19170 = pi144 & n16747;
  assign n19171 = ~pi144 & ~n16825;
  assign n19172 = ~pi758 & ~n19171;
  assign n19173 = ~n19170 & n19172;
  assign n19174 = pi39 & ~n19169;
  assign n19175 = ~n19173 & n19174;
  assign n19176 = ~pi38 & ~n19165;
  assign n19177 = ~n19175 & n19176;
  assign n19178 = pi736 & ~n18668;
  assign n19179 = ~n19119 & n19178;
  assign n19180 = ~n19177 & n19179;
  assign n19181 = ~n19155 & ~n19180;
  assign n19182 = ~n19103 & ~n19181;
  assign n19183 = ~pi625 & n19182;
  assign n19184 = pi625 & n19122;
  assign n19185 = ~pi1153 & ~n19184;
  assign n19186 = ~n19183 & n19185;
  assign n19187 = ~pi608 & ~n19058;
  assign n19188 = ~n19186 & n19187;
  assign n19189 = ~pi625 & n19122;
  assign n19190 = pi625 & n19182;
  assign n19191 = pi1153 & ~n19189;
  assign n19192 = ~n19190 & n19191;
  assign n19193 = pi608 & ~n19062;
  assign n19194 = ~n19192 & n19193;
  assign n19195 = ~n19188 & ~n19194;
  assign n19196 = pi778 & ~n19195;
  assign n19197 = ~pi778 & n19182;
  assign n19198 = ~n19196 & ~n19197;
  assign n19199 = ~pi609 & ~n19198;
  assign n19200 = ~pi1155 & ~n19154;
  assign n19201 = ~n19199 & n19200;
  assign n19202 = ~pi660 & ~n19130;
  assign n19203 = ~n19201 & n19202;
  assign n19204 = ~pi609 & n19065;
  assign n19205 = pi609 & ~n19198;
  assign n19206 = pi1155 & ~n19204;
  assign n19207 = ~n19205 & n19206;
  assign n19208 = pi660 & ~n19134;
  assign n19209 = ~n19207 & n19208;
  assign n19210 = ~n19203 & ~n19209;
  assign n19211 = pi785 & ~n19210;
  assign n19212 = ~pi785 & ~n19198;
  assign n19213 = ~n19211 & ~n19212;
  assign n19214 = ~pi618 & ~n19213;
  assign n19215 = pi618 & n19068;
  assign n19216 = ~pi1154 & ~n19215;
  assign n19217 = ~n19214 & n19216;
  assign n19218 = ~pi627 & ~n19142;
  assign n19219 = ~n19217 & n19218;
  assign n19220 = ~pi618 & n19068;
  assign n19221 = pi618 & ~n19213;
  assign n19222 = pi1154 & ~n19220;
  assign n19223 = ~n19221 & n19222;
  assign n19224 = pi627 & ~n19146;
  assign n19225 = ~n19223 & n19224;
  assign n19226 = ~n19219 & ~n19225;
  assign n19227 = pi781 & ~n19226;
  assign n19228 = ~pi781 & ~n19213;
  assign n19229 = ~n19227 & ~n19228;
  assign n19230 = ~pi619 & ~n19229;
  assign n19231 = ~pi1159 & ~n19153;
  assign n19232 = ~n19230 & n19231;
  assign n19233 = ~pi648 & ~n19152;
  assign n19234 = ~n19232 & n19233;
  assign n19235 = pi619 & ~n19038;
  assign n19236 = ~pi619 & n19149;
  assign n19237 = ~pi1159 & ~n19235;
  assign n19238 = ~n19236 & n19237;
  assign n19239 = ~pi619 & ~n19070;
  assign n19240 = pi619 & ~n19229;
  assign n19241 = pi1159 & ~n19239;
  assign n19242 = ~n19240 & n19241;
  assign n19243 = pi648 & ~n19238;
  assign n19244 = ~n19242 & n19243;
  assign n19245 = ~n19234 & ~n19244;
  assign n19246 = pi789 & ~n19245;
  assign n19247 = ~pi789 & ~n19229;
  assign n19248 = ~n19246 & ~n19247;
  assign n19249 = ~pi788 & n19248;
  assign n19250 = ~pi789 & ~n19149;
  assign n19251 = ~n19152 & ~n19238;
  assign n19252 = pi789 & ~n19251;
  assign n19253 = ~n19250 & ~n19252;
  assign n19254 = ~pi626 & n19253;
  assign n19255 = pi626 & ~n19038;
  assign n19256 = ~pi1158 & ~n19255;
  assign n19257 = ~n19254 & n19256;
  assign n19258 = ~n16995 & ~n19257;
  assign n19259 = ~pi626 & n19248;
  assign n19260 = pi626 & ~n19073;
  assign n19261 = ~pi641 & ~n19260;
  assign n19262 = ~n19259 & n19261;
  assign n19263 = ~n19258 & ~n19262;
  assign n19264 = pi626 & n19253;
  assign n19265 = ~pi626 & ~n19038;
  assign n19266 = pi1158 & ~n19265;
  assign n19267 = ~n19264 & n19266;
  assign n19268 = ~n17002 & ~n19267;
  assign n19269 = pi626 & n19248;
  assign n19270 = ~pi626 & ~n19073;
  assign n19271 = pi641 & ~n19270;
  assign n19272 = ~n19269 & n19271;
  assign n19273 = ~n19268 & ~n19272;
  assign n19274 = ~n19263 & ~n19273;
  assign n19275 = pi788 & ~n19274;
  assign n19276 = ~n19249 & ~n19275;
  assign n19277 = ~n16643 & ~n19276;
  assign n19278 = ~n19257 & ~n19267;
  assign n19279 = pi788 & ~n19278;
  assign n19280 = ~pi788 & ~n19253;
  assign n19281 = ~n19279 & ~n19280;
  assign n19282 = ~n16633 & ~n19281;
  assign n19283 = pi629 & n19084;
  assign n19284 = ~n19101 & ~n19283;
  assign n19285 = ~n19282 & n19284;
  assign n19286 = ~n19277 & n19285;
  assign n19287 = pi792 & ~n19286;
  assign n19288 = ~pi792 & ~n19276;
  assign n19289 = ~n19287 & ~n19288;
  assign n19290 = ~pi647 & n19289;
  assign n19291 = ~n15925 & ~n19281;
  assign n19292 = n15925 & n19038;
  assign n19293 = ~n19291 & ~n19292;
  assign n19294 = pi647 & n19293;
  assign n19295 = ~pi1157 & ~n19294;
  assign n19296 = ~n19290 & n19295;
  assign n19297 = ~pi630 & ~n19092;
  assign n19298 = ~n19296 & n19297;
  assign n19299 = ~pi647 & n19293;
  assign n19300 = pi647 & n19289;
  assign n19301 = pi1157 & ~n19299;
  assign n19302 = ~n19300 & n19301;
  assign n19303 = pi630 & ~n19096;
  assign n19304 = ~n19302 & n19303;
  assign n19305 = ~n19298 & ~n19304;
  assign n19306 = pi787 & ~n19305;
  assign n19307 = ~pi787 & n19289;
  assign n19308 = ~n19306 & ~n19307;
  assign n19309 = pi644 & ~n19308;
  assign n19310 = pi715 & ~n19100;
  assign n19311 = ~n19309 & n19310;
  assign n19312 = ~n15960 & ~n19293;
  assign n19313 = n15960 & n19038;
  assign n19314 = ~n19312 & ~n19313;
  assign n19315 = pi644 & n19314;
  assign n19316 = ~pi644 & ~n19038;
  assign n19317 = ~pi715 & ~n19316;
  assign n19318 = ~n19315 & n19317;
  assign n19319 = pi1160 & ~n19318;
  assign n19320 = ~n19311 & n19319;
  assign n19321 = pi644 & n19099;
  assign n19322 = ~pi715 & ~n19321;
  assign n19323 = ~pi644 & n19314;
  assign n19324 = pi644 & ~n19038;
  assign n19325 = pi715 & ~n19324;
  assign n19326 = ~n19323 & n19325;
  assign n19327 = ~pi1160 & ~n19326;
  assign n19328 = ~n19322 & n19327;
  assign n19329 = ~n19320 & ~n19328;
  assign n19330 = pi790 & ~n19329;
  assign n19331 = ~pi644 & n19327;
  assign n19332 = pi790 & ~n19331;
  assign n19333 = ~n19308 & ~n19332;
  assign n19334 = ~n19330 & ~n19333;
  assign n19335 = n6258 & ~n19334;
  assign n19336 = ~pi57 & ~n19037;
  assign n19337 = ~n19335 & n19336;
  assign n19338 = ~pi832 & ~n19036;
  assign n19339 = ~n19337 & n19338;
  assign po301 = ~n19035 & ~n19339;
  assign n19341 = ~pi145 & po1038;
  assign n19342 = ~pi145 & ~n16219;
  assign n19343 = n15747 & ~n19342;
  assign n19344 = ~pi698 & n9829;
  assign n19345 = n19342 & ~n19344;
  assign n19346 = ~pi145 & ~n16228;
  assign n19347 = n16227 & ~n19346;
  assign n19348 = ~pi145 & ~n17276;
  assign n19349 = ~pi38 & ~n17272;
  assign n19350 = n9829 & ~n19349;
  assign n19351 = ~pi38 & ~pi145;
  assign n19352 = n19350 & ~n19351;
  assign n19353 = ~n19348 & ~n19352;
  assign n19354 = ~pi698 & ~n19347;
  assign n19355 = ~n19353 & n19354;
  assign n19356 = ~n19345 & ~n19355;
  assign n19357 = ~pi778 & n19356;
  assign n19358 = ~pi625 & n19342;
  assign n19359 = pi625 & ~n19356;
  assign n19360 = pi1153 & ~n19358;
  assign n19361 = ~n19359 & n19360;
  assign n19362 = pi625 & n19342;
  assign n19363 = ~pi625 & ~n19356;
  assign n19364 = ~pi1153 & ~n19362;
  assign n19365 = ~n19363 & n19364;
  assign n19366 = ~n19361 & ~n19365;
  assign n19367 = pi778 & ~n19366;
  assign n19368 = ~n19357 & ~n19367;
  assign n19369 = ~n15741 & n19368;
  assign n19370 = n15741 & n19342;
  assign n19371 = ~n19369 & ~n19370;
  assign n19372 = ~n15747 & n19371;
  assign n19373 = ~n19343 & ~n19372;
  assign n19374 = ~n15753 & n19373;
  assign n19375 = n15753 & n19342;
  assign n19376 = ~n19374 & ~n19375;
  assign n19377 = ~n15759 & ~n19376;
  assign n19378 = n15759 & n19342;
  assign n19379 = ~n19377 & ~n19378;
  assign n19380 = ~pi792 & n19379;
  assign n19381 = ~pi628 & n19342;
  assign n19382 = pi628 & ~n19379;
  assign n19383 = pi1156 & ~n19381;
  assign n19384 = ~n19382 & n19383;
  assign n19385 = pi628 & n19342;
  assign n19386 = ~pi628 & ~n19379;
  assign n19387 = ~pi1156 & ~n19385;
  assign n19388 = ~n19386 & n19387;
  assign n19389 = ~n19384 & ~n19388;
  assign n19390 = pi792 & ~n19389;
  assign n19391 = ~n19380 & ~n19390;
  assign n19392 = pi647 & ~pi1157;
  assign n19393 = ~pi647 & pi1157;
  assign n19394 = ~n19392 & ~n19393;
  assign n19395 = n19391 & n19394;
  assign n19396 = n19342 & ~n19394;
  assign n19397 = ~n19395 & ~n19396;
  assign n19398 = pi787 & ~n19397;
  assign n19399 = ~pi787 & n19391;
  assign n19400 = ~n19398 & ~n19399;
  assign n19401 = ~pi644 & ~n19400;
  assign n19402 = pi715 & ~n19401;
  assign n19403 = pi145 & ~n9829;
  assign n19404 = ~pi767 & n16570;
  assign n19405 = ~n19346 & ~n19404;
  assign n19406 = pi38 & ~n19405;
  assign n19407 = ~n18599 & ~n19351;
  assign n19408 = ~pi145 & ~n16214;
  assign n19409 = pi767 & ~n19408;
  assign n19410 = ~pi145 & ~pi767;
  assign n19411 = n16514 & n19410;
  assign n19412 = ~n19407 & ~n19411;
  assign n19413 = ~n19409 & n19412;
  assign n19414 = n9829 & ~n19406;
  assign n19415 = ~n19413 & n19414;
  assign n19416 = ~n19403 & ~n19415;
  assign n19417 = ~n15777 & ~n19416;
  assign n19418 = n15777 & ~n19342;
  assign n19419 = ~n19417 & ~n19418;
  assign n19420 = ~pi785 & ~n19419;
  assign n19421 = ~n15786 & ~n19342;
  assign n19422 = pi609 & n19417;
  assign n19423 = ~n19421 & ~n19422;
  assign n19424 = pi1155 & ~n19423;
  assign n19425 = ~n16585 & ~n19342;
  assign n19426 = ~pi609 & n19417;
  assign n19427 = ~n19425 & ~n19426;
  assign n19428 = ~pi1155 & ~n19427;
  assign n19429 = ~n19424 & ~n19428;
  assign n19430 = pi785 & ~n19429;
  assign n19431 = ~n19420 & ~n19430;
  assign n19432 = ~pi781 & ~n19431;
  assign n19433 = ~pi618 & n19342;
  assign n19434 = pi618 & n19431;
  assign n19435 = pi1154 & ~n19433;
  assign n19436 = ~n19434 & n19435;
  assign n19437 = ~pi618 & n19431;
  assign n19438 = pi618 & n19342;
  assign n19439 = ~pi1154 & ~n19438;
  assign n19440 = ~n19437 & n19439;
  assign n19441 = ~n19436 & ~n19440;
  assign n19442 = pi781 & ~n19441;
  assign n19443 = ~n19432 & ~n19442;
  assign n19444 = ~pi789 & ~n19443;
  assign n19445 = ~pi619 & n19342;
  assign n19446 = pi619 & n19443;
  assign n19447 = pi1159 & ~n19445;
  assign n19448 = ~n19446 & n19447;
  assign n19449 = ~pi619 & n19443;
  assign n19450 = pi619 & n19342;
  assign n19451 = ~pi1159 & ~n19450;
  assign n19452 = ~n19449 & n19451;
  assign n19453 = ~n19448 & ~n19452;
  assign n19454 = pi789 & ~n19453;
  assign n19455 = ~n19444 & ~n19454;
  assign n19456 = n15820 & n19455;
  assign n19457 = ~n15820 & n19342;
  assign n19458 = ~n19456 & ~n19457;
  assign n19459 = pi788 & ~n19458;
  assign n19460 = ~pi788 & n19455;
  assign n19461 = ~n19459 & ~n19460;
  assign n19462 = ~n15925 & ~n19461;
  assign n19463 = n15925 & n19342;
  assign n19464 = ~n19462 & ~n19463;
  assign n19465 = ~n15960 & ~n19464;
  assign n19466 = n15960 & n19342;
  assign n19467 = ~n19465 & ~n19466;
  assign n19468 = pi644 & ~n19467;
  assign n19469 = ~pi644 & n19342;
  assign n19470 = ~pi715 & ~n19469;
  assign n19471 = ~n19468 & n19470;
  assign n19472 = pi1160 & ~n19471;
  assign n19473 = ~n19402 & n19472;
  assign n19474 = pi644 & ~n19400;
  assign n19475 = pi630 & ~pi647;
  assign n19476 = ~pi630 & pi647;
  assign n19477 = ~n19475 & ~n19476;
  assign n19478 = n15959 & ~n19477;
  assign n19479 = n19464 & n19478;
  assign n19480 = ~n15959 & n19397;
  assign n19481 = ~n19479 & ~n19480;
  assign n19482 = pi787 & ~n19481;
  assign n19483 = ~n16633 & n19461;
  assign n19484 = ~pi629 & n19384;
  assign n19485 = pi629 & n19388;
  assign n19486 = ~n19484 & ~n19485;
  assign n19487 = ~n19483 & n19486;
  assign n19488 = pi792 & ~n19487;
  assign n19489 = n15828 & ~n19376;
  assign n19490 = ~n15758 & ~n19458;
  assign n19491 = ~n19489 & ~n19490;
  assign n19492 = pi788 & ~n19491;
  assign n19493 = pi618 & ~n19371;
  assign n19494 = pi609 & n19368;
  assign n19495 = ~n19344 & ~n19415;
  assign n19496 = ~pi767 & ~n16808;
  assign n19497 = n18669 & ~n19496;
  assign n19498 = ~pi145 & ~n19497;
  assign n19499 = ~pi767 & n15781;
  assign n19500 = ~n16921 & ~n19499;
  assign n19501 = pi145 & ~n19500;
  assign n19502 = n6081 & n19501;
  assign n19503 = pi38 & ~n19502;
  assign n19504 = ~n19498 & n19503;
  assign n19505 = ~pi145 & ~n16647;
  assign n19506 = pi145 & ~n17397;
  assign n19507 = ~pi767 & ~n19505;
  assign n19508 = ~n19506 & n19507;
  assign n19509 = ~pi145 & n16653;
  assign n19510 = pi145 & n16657;
  assign n19511 = pi767 & ~n19509;
  assign n19512 = ~n19510 & n19511;
  assign n19513 = ~pi39 & ~n19508;
  assign n19514 = ~n19512 & n19513;
  assign n19515 = pi145 & n16825;
  assign n19516 = ~pi145 & ~n16747;
  assign n19517 = pi767 & ~n19515;
  assign n19518 = ~n19516 & n19517;
  assign n19519 = ~pi145 & n16877;
  assign n19520 = pi145 & n16913;
  assign n19521 = ~pi767 & ~n19519;
  assign n19522 = ~n19520 & n19521;
  assign n19523 = pi39 & ~n19522;
  assign n19524 = ~n19518 & n19523;
  assign n19525 = ~pi38 & ~n19514;
  assign n19526 = ~n19524 & n19525;
  assign n19527 = ~pi698 & ~n19504;
  assign n19528 = ~n19526 & n19527;
  assign n19529 = ~n19495 & ~n19528;
  assign n19530 = ~n19403 & ~n19529;
  assign n19531 = ~pi625 & n19530;
  assign n19532 = pi625 & n19416;
  assign n19533 = ~pi1153 & ~n19532;
  assign n19534 = ~n19531 & n19533;
  assign n19535 = ~pi608 & ~n19361;
  assign n19536 = ~n19534 & n19535;
  assign n19537 = ~pi625 & n19416;
  assign n19538 = pi625 & n19530;
  assign n19539 = pi1153 & ~n19537;
  assign n19540 = ~n19538 & n19539;
  assign n19541 = pi608 & ~n19365;
  assign n19542 = ~n19540 & n19541;
  assign n19543 = ~n19536 & ~n19542;
  assign n19544 = pi778 & ~n19543;
  assign n19545 = ~pi778 & n19530;
  assign n19546 = ~n19544 & ~n19545;
  assign n19547 = ~pi609 & ~n19546;
  assign n19548 = ~pi1155 & ~n19494;
  assign n19549 = ~n19547 & n19548;
  assign n19550 = ~pi660 & ~n19424;
  assign n19551 = ~n19549 & n19550;
  assign n19552 = ~pi609 & n19368;
  assign n19553 = pi609 & ~n19546;
  assign n19554 = pi1155 & ~n19552;
  assign n19555 = ~n19553 & n19554;
  assign n19556 = pi660 & ~n19428;
  assign n19557 = ~n19555 & n19556;
  assign n19558 = ~n19551 & ~n19557;
  assign n19559 = pi785 & ~n19558;
  assign n19560 = ~pi785 & ~n19546;
  assign n19561 = ~n19559 & ~n19560;
  assign n19562 = ~pi618 & ~n19561;
  assign n19563 = ~pi1154 & ~n19493;
  assign n19564 = ~n19562 & n19563;
  assign n19565 = ~pi627 & ~n19436;
  assign n19566 = ~n19564 & n19565;
  assign n19567 = ~pi618 & ~n19371;
  assign n19568 = pi618 & ~n19561;
  assign n19569 = pi1154 & ~n19567;
  assign n19570 = ~n19568 & n19569;
  assign n19571 = pi627 & ~n19440;
  assign n19572 = ~n19570 & n19571;
  assign n19573 = ~n19566 & ~n19572;
  assign n19574 = pi781 & ~n19573;
  assign n19575 = ~pi781 & ~n19561;
  assign n19576 = ~n19574 & ~n19575;
  assign n19577 = ~pi789 & n19576;
  assign n19578 = ~pi619 & n19373;
  assign n19579 = pi619 & ~n19576;
  assign n19580 = pi1159 & ~n19578;
  assign n19581 = ~n19579 & n19580;
  assign n19582 = pi648 & ~n19452;
  assign n19583 = ~n19581 & n19582;
  assign n19584 = ~pi619 & ~n19576;
  assign n19585 = pi619 & n19373;
  assign n19586 = ~pi1159 & ~n19585;
  assign n19587 = ~n19584 & n19586;
  assign n19588 = ~pi648 & ~n19448;
  assign n19589 = ~n19587 & n19588;
  assign n19590 = pi789 & ~n19583;
  assign n19591 = ~n19589 & n19590;
  assign n19592 = n15833 & ~n19577;
  assign n19593 = ~n19591 & n19592;
  assign n19594 = ~n16644 & ~n19492;
  assign n19595 = ~n19593 & n19594;
  assign n19596 = ~n19488 & ~n19595;
  assign n19597 = n18841 & ~n19596;
  assign n19598 = ~n19482 & ~n19597;
  assign n19599 = ~pi644 & n19598;
  assign n19600 = ~pi715 & ~n19474;
  assign n19601 = ~n19599 & n19600;
  assign n19602 = pi644 & n19342;
  assign n19603 = ~pi644 & ~n19467;
  assign n19604 = pi715 & ~n19602;
  assign n19605 = ~n19603 & n19604;
  assign n19606 = ~pi1160 & ~n19605;
  assign n19607 = ~n19601 & n19606;
  assign n19608 = ~n19473 & ~n19607;
  assign n19609 = pi790 & ~n19608;
  assign n19610 = pi644 & n19472;
  assign n19611 = pi790 & ~n19610;
  assign n19612 = n19598 & ~n19611;
  assign n19613 = ~n19609 & ~n19612;
  assign n19614 = ~po1038 & ~n19613;
  assign n19615 = ~pi832 & ~n19341;
  assign n19616 = ~n19614 & n19615;
  assign n19617 = ~pi145 & ~n2923;
  assign n19618 = ~pi698 & n15726;
  assign n19619 = ~n19617 & ~n19618;
  assign n19620 = ~pi778 & n19619;
  assign n19621 = ~pi625 & n19618;
  assign n19622 = ~n19619 & ~n19621;
  assign n19623 = pi1153 & ~n19622;
  assign n19624 = ~pi1153 & ~n19617;
  assign n19625 = ~n19621 & n19624;
  assign n19626 = ~n19623 & ~n19625;
  assign n19627 = pi778 & ~n19626;
  assign n19628 = ~n19620 & ~n19627;
  assign n19629 = ~n15742 & n19628;
  assign n19630 = ~n15748 & n19629;
  assign n19631 = ~n15754 & n19630;
  assign n19632 = ~n15760 & n19631;
  assign n19633 = ~n15766 & n19632;
  assign n19634 = n19394 & n19633;
  assign n19635 = ~n19394 & n19617;
  assign n19636 = ~n19634 & ~n19635;
  assign n19637 = ~n15959 & n19636;
  assign n19638 = n15925 & n19617;
  assign n19639 = ~n19499 & ~n19617;
  assign n19640 = ~n15778 & ~n19639;
  assign n19641 = ~pi785 & ~n19640;
  assign n19642 = ~n15787 & ~n19639;
  assign n19643 = pi1155 & ~n19642;
  assign n19644 = ~n15790 & n19640;
  assign n19645 = ~pi1155 & ~n19644;
  assign n19646 = ~n19643 & ~n19645;
  assign n19647 = pi785 & ~n19646;
  assign n19648 = ~n19641 & ~n19647;
  assign n19649 = ~pi781 & ~n19648;
  assign n19650 = ~n15797 & n19648;
  assign n19651 = pi1154 & ~n19650;
  assign n19652 = ~n15800 & n19648;
  assign n19653 = ~pi1154 & ~n19652;
  assign n19654 = ~n19651 & ~n19653;
  assign n19655 = pi781 & ~n19654;
  assign n19656 = ~n19649 & ~n19655;
  assign n19657 = ~pi789 & ~n19656;
  assign n19658 = ~pi619 & n19617;
  assign n19659 = pi619 & n19656;
  assign n19660 = pi1159 & ~n19658;
  assign n19661 = ~n19659 & n19660;
  assign n19662 = ~pi619 & n19656;
  assign n19663 = pi619 & n19617;
  assign n19664 = ~pi1159 & ~n19663;
  assign n19665 = ~n19662 & n19664;
  assign n19666 = ~n19661 & ~n19665;
  assign n19667 = pi789 & ~n19666;
  assign n19668 = ~n19657 & ~n19667;
  assign n19669 = n15820 & n19668;
  assign n19670 = ~n15820 & n19617;
  assign n19671 = ~n19669 & ~n19670;
  assign n19672 = pi788 & ~n19671;
  assign n19673 = ~pi788 & n19668;
  assign n19674 = ~n19672 & ~n19673;
  assign n19675 = ~n15925 & ~n19674;
  assign n19676 = n19478 & ~n19638;
  assign n19677 = ~n19675 & n19676;
  assign n19678 = ~n19637 & ~n19677;
  assign n19679 = pi787 & ~n19678;
  assign n19680 = ~n15758 & ~n19671;
  assign n19681 = n15828 & n19631;
  assign n19682 = ~n19680 & ~n19681;
  assign n19683 = pi788 & ~n19682;
  assign n19684 = pi618 & n19629;
  assign n19685 = pi609 & n19628;
  assign n19686 = ~n15780 & ~n19619;
  assign n19687 = pi625 & n19686;
  assign n19688 = n19639 & ~n19686;
  assign n19689 = ~n19687 & ~n19688;
  assign n19690 = n19624 & ~n19689;
  assign n19691 = ~pi608 & ~n19623;
  assign n19692 = ~n19690 & n19691;
  assign n19693 = pi1153 & n19639;
  assign n19694 = ~n19687 & n19693;
  assign n19695 = pi608 & ~n19625;
  assign n19696 = ~n19694 & n19695;
  assign n19697 = ~n19692 & ~n19696;
  assign n19698 = pi778 & ~n19697;
  assign n19699 = ~pi778 & ~n19688;
  assign n19700 = ~n19698 & ~n19699;
  assign n19701 = ~pi609 & ~n19700;
  assign n19702 = ~pi1155 & ~n19685;
  assign n19703 = ~n19701 & n19702;
  assign n19704 = ~pi660 & ~n19643;
  assign n19705 = ~n19703 & n19704;
  assign n19706 = ~pi609 & n19628;
  assign n19707 = pi609 & ~n19700;
  assign n19708 = pi1155 & ~n19706;
  assign n19709 = ~n19707 & n19708;
  assign n19710 = pi660 & ~n19645;
  assign n19711 = ~n19709 & n19710;
  assign n19712 = ~n19705 & ~n19711;
  assign n19713 = pi785 & ~n19712;
  assign n19714 = ~pi785 & ~n19700;
  assign n19715 = ~n19713 & ~n19714;
  assign n19716 = ~pi618 & ~n19715;
  assign n19717 = ~pi1154 & ~n19684;
  assign n19718 = ~n19716 & n19717;
  assign n19719 = ~pi627 & ~n19651;
  assign n19720 = ~n19718 & n19719;
  assign n19721 = ~pi618 & n19629;
  assign n19722 = pi618 & ~n19715;
  assign n19723 = pi1154 & ~n19721;
  assign n19724 = ~n19722 & n19723;
  assign n19725 = pi627 & ~n19653;
  assign n19726 = ~n19724 & n19725;
  assign n19727 = ~n19720 & ~n19726;
  assign n19728 = pi781 & ~n19727;
  assign n19729 = ~pi781 & ~n19715;
  assign n19730 = ~n19728 & ~n19729;
  assign n19731 = ~pi789 & n19730;
  assign n19732 = ~pi619 & n19630;
  assign n19733 = pi619 & ~n19730;
  assign n19734 = pi1159 & ~n19732;
  assign n19735 = ~n19733 & n19734;
  assign n19736 = pi648 & ~n19665;
  assign n19737 = ~n19735 & n19736;
  assign n19738 = pi619 & n19630;
  assign n19739 = ~pi619 & ~n19730;
  assign n19740 = ~pi1159 & ~n19738;
  assign n19741 = ~n19739 & n19740;
  assign n19742 = ~pi648 & ~n19661;
  assign n19743 = ~n19741 & n19742;
  assign n19744 = pi789 & ~n19737;
  assign n19745 = ~n19743 & n19744;
  assign n19746 = n15833 & ~n19731;
  assign n19747 = ~n19745 & n19746;
  assign n19748 = ~n19683 & ~n19747;
  assign n19749 = ~n16644 & ~n19748;
  assign n19750 = n15763 & ~n19674;
  assign n19751 = n15772 & n19632;
  assign n19752 = ~pi629 & ~n19751;
  assign n19753 = ~n19750 & n19752;
  assign n19754 = n15762 & ~n19674;
  assign n19755 = n15909 & n19632;
  assign n19756 = pi629 & ~n19755;
  assign n19757 = ~n19754 & n19756;
  assign n19758 = pi792 & ~n19753;
  assign n19759 = ~n19757 & n19758;
  assign n19760 = n18841 & ~n19759;
  assign n19761 = ~n19749 & n19760;
  assign n19762 = ~n19679 & ~n19761;
  assign n19763 = ~pi790 & n19762;
  assign n19764 = pi787 & ~n19636;
  assign n19765 = ~pi787 & n19633;
  assign n19766 = ~n19764 & ~n19765;
  assign n19767 = ~pi644 & ~n19766;
  assign n19768 = pi644 & n19762;
  assign n19769 = pi715 & ~n19767;
  assign n19770 = ~n19768 & n19769;
  assign n19771 = ~n15925 & ~n15960;
  assign n19772 = n19617 & ~n19771;
  assign n19773 = ~n15960 & n19675;
  assign n19774 = ~n19772 & ~n19773;
  assign n19775 = pi644 & ~n19774;
  assign n19776 = ~pi644 & n19617;
  assign n19777 = ~pi715 & ~n19776;
  assign n19778 = ~n19775 & n19777;
  assign n19779 = pi1160 & ~n19778;
  assign n19780 = ~n19770 & n19779;
  assign n19781 = ~pi644 & ~n19774;
  assign n19782 = pi644 & n19617;
  assign n19783 = pi715 & ~n19782;
  assign n19784 = ~n19781 & n19783;
  assign n19785 = pi644 & ~n19766;
  assign n19786 = ~pi644 & n19762;
  assign n19787 = ~pi715 & ~n19785;
  assign n19788 = ~n19786 & n19787;
  assign n19789 = ~pi1160 & ~n19784;
  assign n19790 = ~n19788 & n19789;
  assign n19791 = ~n19780 & ~n19790;
  assign n19792 = pi790 & ~n19791;
  assign n19793 = pi832 & ~n19763;
  assign n19794 = ~n19792 & n19793;
  assign po302 = ~n19616 & ~n19794;
  assign n19796 = ~pi146 & ~n2923;
  assign n19797 = pi743 & pi947;
  assign n19798 = pi907 & ~pi947;
  assign n19799 = pi735 & n19798;
  assign n19800 = ~n19797 & ~n19799;
  assign n19801 = n2923 & n19800;
  assign n19802 = pi832 & ~n19796;
  assign n19803 = ~n19801 & n19802;
  assign n19804 = ~pi146 & ~n9830;
  assign n19805 = ~pi146 & ~n16228;
  assign n19806 = n16228 & n19800;
  assign n19807 = pi38 & ~n19805;
  assign n19808 = ~n19806 & n19807;
  assign n19809 = pi146 & ~n16051;
  assign n19810 = n16051 & ~n19800;
  assign n19811 = pi299 & ~n19809;
  assign n19812 = ~n19810 & n19811;
  assign n19813 = pi146 & ~n16055;
  assign n19814 = n16055 & ~n19800;
  assign n19815 = ~pi299 & ~n19813;
  assign n19816 = ~n19814 & n19815;
  assign n19817 = ~n19812 & ~n19816;
  assign n19818 = ~pi39 & ~n19817;
  assign n19819 = pi146 & ~n16184;
  assign n19820 = n16184 & ~n19800;
  assign n19821 = n6194 & ~n19819;
  assign n19822 = ~n19820 & n19821;
  assign n19823 = n16153 & ~n19800;
  assign n19824 = pi146 & ~n16153;
  assign n19825 = ~n6194 & ~n19823;
  assign n19826 = ~n19824 & n19825;
  assign n19827 = ~n2608 & ~n19826;
  assign n19828 = ~n19822 & n19827;
  assign n19829 = ~pi146 & ~n16063;
  assign n19830 = n16063 & n19800;
  assign n19831 = ~n19829 & ~n19830;
  assign n19832 = n2608 & n19831;
  assign n19833 = ~pi223 & ~n19832;
  assign n19834 = ~n19828 & n19833;
  assign n19835 = n16104 & ~n19800;
  assign n19836 = pi146 & ~n16104;
  assign n19837 = ~n19835 & ~n19836;
  assign n19838 = ~n6194 & ~n19837;
  assign n19839 = ~pi146 & ~n16122;
  assign n19840 = n16122 & n19800;
  assign n19841 = n6194 & ~n19839;
  assign n19842 = ~n19840 & n19841;
  assign n19843 = pi223 & ~n19842;
  assign n19844 = ~n19838 & n19843;
  assign n19845 = ~n19834 & ~n19844;
  assign n19846 = ~pi299 & ~n19845;
  assign n19847 = pi146 & n16208;
  assign n19848 = ~n19835 & ~n19847;
  assign n19849 = pi215 & ~n19848;
  assign n19850 = n3302 & ~n19831;
  assign n19851 = pi146 & n16196;
  assign n19852 = ~n3302 & ~n19823;
  assign n19853 = ~n19851 & n19852;
  assign n19854 = ~pi215 & ~n19850;
  assign n19855 = ~n19853 & n19854;
  assign n19856 = pi299 & ~n19849;
  assign n19857 = ~n19855 & n19856;
  assign n19858 = ~n19846 & ~n19857;
  assign n19859 = pi39 & ~n19858;
  assign n19860 = ~pi38 & ~n19818;
  assign n19861 = ~n19859 & n19860;
  assign n19862 = n9830 & ~n19808;
  assign n19863 = ~n19861 & n19862;
  assign n19864 = ~pi832 & ~n19804;
  assign n19865 = ~n19863 & n19864;
  assign po303 = n19803 | n19865;
  assign n19867 = ~pi147 & ~n2923;
  assign n19868 = ~pi770 & pi947;
  assign n19869 = pi726 & n19798;
  assign n19870 = ~n19868 & ~n19869;
  assign n19871 = n2923 & ~n19870;
  assign n19872 = pi832 & ~n19867;
  assign n19873 = ~n19871 & n19872;
  assign n19874 = ~pi147 & ~n9830;
  assign n19875 = ~pi947 & n16057;
  assign n19876 = ~pi39 & ~n19875;
  assign n19877 = ~pi947 & n16199;
  assign n19878 = n16153 & n19798;
  assign n19879 = ~n16197 & ~n19878;
  assign n19880 = ~n3302 & ~n19879;
  assign n19881 = ~pi215 & ~n19880;
  assign n19882 = ~n19877 & n19881;
  assign n19883 = n16104 & n19798;
  assign n19884 = pi215 & ~n16207;
  assign n19885 = ~n19883 & n19884;
  assign n19886 = ~n19882 & ~n19885;
  assign n19887 = pi299 & ~n19886;
  assign n19888 = ~n16191 & ~n19887;
  assign n19889 = pi947 & n16190;
  assign n19890 = ~pi299 & n19889;
  assign n19891 = n19888 & ~n19890;
  assign n19892 = pi39 & ~n19891;
  assign n19893 = ~n19876 & ~n19892;
  assign n19894 = ~pi38 & n19893;
  assign n19895 = pi38 & ~pi947;
  assign n19896 = n16216 & n19895;
  assign n19897 = ~n19894 & ~n19896;
  assign n19898 = ~pi770 & ~n19897;
  assign n19899 = pi770 & n16218;
  assign n19900 = ~pi147 & ~n19899;
  assign n19901 = ~n19898 & n19900;
  assign n19902 = ~n16217 & ~n19896;
  assign n19903 = pi947 & n16057;
  assign n19904 = ~pi39 & ~n19903;
  assign n19905 = ~pi299 & ~n19889;
  assign n19906 = pi215 & pi947;
  assign n19907 = n16104 & n19906;
  assign n19908 = pi299 & ~n19907;
  assign n19909 = pi947 & n16153;
  assign n19910 = ~n3302 & ~n19909;
  assign n19911 = pi947 & n16063;
  assign n19912 = n3302 & ~n19911;
  assign n19913 = ~pi215 & ~n19912;
  assign n19914 = ~n19910 & n19913;
  assign n19915 = n19908 & ~n19914;
  assign n19916 = ~n19905 & ~n19915;
  assign n19917 = pi39 & ~n19916;
  assign n19918 = ~n19904 & ~n19917;
  assign n19919 = ~pi38 & ~n19918;
  assign n19920 = n19902 & ~n19919;
  assign n19921 = pi147 & ~pi770;
  assign n19922 = n19920 & n19921;
  assign n19923 = ~pi726 & ~n19922;
  assign n19924 = ~n19901 & n19923;
  assign n19925 = ~pi147 & ~n16228;
  assign n19926 = n16228 & n19798;
  assign n19927 = pi38 & ~n19926;
  assign n19928 = ~n19925 & n19927;
  assign n19929 = n16199 & ~n19798;
  assign n19930 = ~n16197 & ~n19909;
  assign n19931 = ~n3302 & ~n19930;
  assign n19932 = ~pi215 & ~n19931;
  assign n19933 = ~n19929 & n19932;
  assign n19934 = ~n19884 & ~n19933;
  assign n19935 = ~n19907 & ~n19934;
  assign n19936 = pi299 & ~n19935;
  assign n19937 = ~pi299 & n16190;
  assign n19938 = ~n19798 & n19937;
  assign n19939 = ~n19936 & ~n19938;
  assign n19940 = pi39 & ~n19939;
  assign n19941 = n16057 & ~n19798;
  assign n19942 = ~pi39 & n19941;
  assign n19943 = ~n19940 & ~n19942;
  assign n19944 = ~pi147 & n19943;
  assign n19945 = pi215 & ~n19883;
  assign n19946 = ~n3302 & ~n19878;
  assign n19947 = pi907 & n16063;
  assign n19948 = ~pi947 & n19947;
  assign n19949 = n3302 & ~n19948;
  assign n19950 = ~n19946 & ~n19949;
  assign n19951 = ~pi215 & ~n19950;
  assign n19952 = ~n19945 & ~n19951;
  assign n19953 = pi299 & ~n19952;
  assign n19954 = n16190 & n19798;
  assign n19955 = ~pi299 & ~n19954;
  assign n19956 = ~n19953 & ~n19955;
  assign n19957 = pi39 & ~n19956;
  assign n19958 = n16057 & n19798;
  assign n19959 = ~pi39 & ~n19958;
  assign n19960 = ~n19957 & ~n19959;
  assign n19961 = pi147 & n19960;
  assign n19962 = ~pi38 & ~n19961;
  assign n19963 = ~n19944 & n19962;
  assign n19964 = pi770 & ~n19928;
  assign n19965 = ~n19963 & n19964;
  assign n19966 = n6220 & n16216;
  assign n19967 = ~pi147 & ~n19966;
  assign n19968 = ~n6220 & n16228;
  assign n19969 = pi38 & ~n19968;
  assign n19970 = ~n19967 & n19969;
  assign n19971 = ~n6220 & n19937;
  assign n19972 = pi299 & ~n19934;
  assign n19973 = pi299 & pi947;
  assign n19974 = ~n16191 & ~n19973;
  assign n19975 = ~n19971 & n19974;
  assign n19976 = ~n19972 & n19975;
  assign n19977 = pi39 & n19976;
  assign n19978 = ~n6220 & n16057;
  assign n19979 = ~pi39 & ~n19978;
  assign n19980 = n16057 & n19979;
  assign n19981 = ~n19977 & ~n19980;
  assign n19982 = ~pi147 & n19981;
  assign n19983 = pi215 & ~n16203;
  assign n19984 = ~n6220 & n16199;
  assign n19985 = ~pi215 & ~n19984;
  assign n19986 = ~n16193 & n19985;
  assign n19987 = pi299 & ~n19983;
  assign n19988 = ~n19986 & n19987;
  assign n19989 = ~n19971 & ~n19988;
  assign n19990 = pi39 & n19989;
  assign n19991 = ~n19979 & ~n19990;
  assign n19992 = pi147 & n19991;
  assign n19993 = ~pi38 & ~n19992;
  assign n19994 = ~n19982 & n19993;
  assign n19995 = ~pi770 & ~n19970;
  assign n19996 = ~n19994 & n19995;
  assign n19997 = pi726 & ~n19996;
  assign n19998 = ~n19965 & n19997;
  assign n19999 = n9830 & ~n19998;
  assign n20000 = ~n19924 & n19999;
  assign n20001 = ~pi832 & ~n19874;
  assign n20002 = ~n20000 & n20001;
  assign po304 = ~n19873 & ~n20002;
  assign n20004 = pi57 & pi148;
  assign n20005 = n6258 & n9829;
  assign n20006 = ~pi148 & ~n20005;
  assign n20007 = ~pi749 & pi947;
  assign n20008 = n19968 & ~n20007;
  assign n20009 = ~pi148 & ~n16228;
  assign n20010 = ~n20008 & ~n20009;
  assign n20011 = pi38 & ~n20010;
  assign n20012 = ~pi148 & ~n16057;
  assign n20013 = ~pi39 & ~n20012;
  assign n20014 = n19978 & ~n20007;
  assign n20015 = n20013 & ~n20014;
  assign n20016 = ~n9399 & ~n19939;
  assign n20017 = ~n16191 & ~n19953;
  assign n20018 = pi148 & ~n20017;
  assign n20019 = ~n20016 & ~n20018;
  assign n20020 = ~pi749 & ~n20019;
  assign n20021 = pi148 & ~n19989;
  assign n20022 = ~pi148 & ~n19976;
  assign n20023 = pi749 & ~n20021;
  assign n20024 = ~n20022 & n20023;
  assign n20025 = ~n20020 & ~n20024;
  assign n20026 = pi39 & ~n20025;
  assign n20027 = ~pi38 & ~n20015;
  assign n20028 = ~n20026 & n20027;
  assign n20029 = pi706 & ~n20011;
  assign n20030 = ~n20028 & n20029;
  assign n20031 = pi148 & ~n16216;
  assign n20032 = pi749 & pi947;
  assign n20033 = n16228 & ~n20032;
  assign n20034 = pi38 & ~n20033;
  assign n20035 = ~n20031 & n20034;
  assign n20036 = n16057 & n20032;
  assign n20037 = n20013 & ~n20036;
  assign n20038 = ~pi148 & ~pi749;
  assign n20039 = ~n16212 & n20038;
  assign n20040 = ~pi148 & ~n16190;
  assign n20041 = n19905 & ~n20040;
  assign n20042 = ~n19907 & ~n19914;
  assign n20043 = pi148 & ~n20042;
  assign n20044 = ~pi148 & ~n19886;
  assign n20045 = pi299 & ~n20043;
  assign n20046 = ~n20044 & n20045;
  assign n20047 = pi749 & ~n20041;
  assign n20048 = ~n20046 & n20047;
  assign n20049 = pi39 & ~n20039;
  assign n20050 = ~n20048 & n20049;
  assign n20051 = ~pi38 & ~n20037;
  assign n20052 = ~n20050 & n20051;
  assign n20053 = ~pi706 & ~n20035;
  assign n20054 = ~n20052 & n20053;
  assign n20055 = n20005 & ~n20054;
  assign n20056 = ~n20030 & n20055;
  assign n20057 = ~pi57 & ~n20006;
  assign n20058 = ~n20056 & n20057;
  assign n20059 = ~pi832 & ~n20004;
  assign n20060 = ~n20058 & n20059;
  assign n20061 = pi148 & ~n2923;
  assign n20062 = pi706 & n19798;
  assign n20063 = n2923 & ~n20032;
  assign n20064 = ~n20062 & n20063;
  assign n20065 = pi832 & ~n20061;
  assign n20066 = ~n20064 & n20065;
  assign po305 = n20060 | n20066;
  assign n20068 = ~pi149 & ~n2923;
  assign n20069 = ~pi755 & pi947;
  assign n20070 = ~pi725 & n19798;
  assign n20071 = ~n20069 & ~n20070;
  assign n20072 = n2923 & ~n20071;
  assign n20073 = pi832 & ~n20068;
  assign n20074 = ~n20072 & n20073;
  assign n20075 = ~pi149 & ~n9830;
  assign n20076 = n16228 & ~n20069;
  assign n20077 = pi149 & ~n16216;
  assign n20078 = pi38 & ~n20076;
  assign n20079 = ~n20077 & n20078;
  assign n20080 = ~pi149 & pi755;
  assign n20081 = ~n16212 & n20080;
  assign n20082 = ~pi149 & ~n16190;
  assign n20083 = n19905 & ~n20082;
  assign n20084 = ~pi149 & ~n19886;
  assign n20085 = ~n15198 & ~n19915;
  assign n20086 = ~n20084 & ~n20085;
  assign n20087 = ~pi755 & ~n20083;
  assign n20088 = ~n20086 & n20087;
  assign n20089 = pi39 & ~n20081;
  assign n20090 = ~n20088 & n20089;
  assign n20091 = ~pi149 & ~n16057;
  assign n20092 = n16057 & n20069;
  assign n20093 = ~pi39 & ~n20091;
  assign n20094 = ~n20092 & n20093;
  assign n20095 = ~pi38 & ~n20094;
  assign n20096 = ~n20090 & n20095;
  assign n20097 = ~n20079 & ~n20096;
  assign n20098 = pi725 & ~n20097;
  assign n20099 = ~n19958 & n20094;
  assign n20100 = pi149 & ~n20017;
  assign n20101 = ~pi149 & n19936;
  assign n20102 = ~n19938 & ~n20100;
  assign n20103 = ~n20101 & n20102;
  assign n20104 = pi755 & ~n20103;
  assign n20105 = ~pi149 & ~n19976;
  assign n20106 = pi149 & ~n19989;
  assign n20107 = ~pi755 & ~n20106;
  assign n20108 = ~n20105 & n20107;
  assign n20109 = ~n20104 & ~n20108;
  assign n20110 = pi39 & ~n20109;
  assign n20111 = ~n20099 & ~n20110;
  assign n20112 = ~pi38 & ~n20111;
  assign n20113 = ~pi149 & ~n16228;
  assign n20114 = ~n19798 & ~n20069;
  assign n20115 = n16228 & ~n20114;
  assign n20116 = pi38 & ~n20113;
  assign n20117 = ~n20115 & n20116;
  assign n20118 = ~pi725 & ~n20117;
  assign n20119 = ~n20112 & n20118;
  assign n20120 = ~n20098 & ~n20119;
  assign n20121 = n9830 & ~n20120;
  assign n20122 = ~pi832 & ~n20075;
  assign n20123 = ~n20121 & n20122;
  assign po306 = ~n20074 & ~n20123;
  assign n20125 = ~pi150 & ~n2923;
  assign n20126 = ~pi751 & pi947;
  assign n20127 = ~pi701 & n19798;
  assign n20128 = ~n20126 & ~n20127;
  assign n20129 = n2923 & ~n20128;
  assign n20130 = pi832 & ~n20125;
  assign n20131 = ~n20129 & n20130;
  assign n20132 = ~pi150 & ~n9830;
  assign n20133 = ~pi150 & ~n16228;
  assign n20134 = ~n19798 & ~n20126;
  assign n20135 = n16228 & ~n20134;
  assign n20136 = pi38 & ~n20133;
  assign n20137 = ~n20135 & n20136;
  assign n20138 = pi150 & ~n16057;
  assign n20139 = n19941 & ~n20126;
  assign n20140 = ~pi39 & ~n20138;
  assign n20141 = ~n20139 & n20140;
  assign n20142 = ~pi150 & n19939;
  assign n20143 = pi150 & n19956;
  assign n20144 = pi751 & ~n20143;
  assign n20145 = ~n20142 & n20144;
  assign n20146 = pi150 & ~n19989;
  assign n20147 = ~pi150 & ~n19976;
  assign n20148 = ~pi751 & ~n20146;
  assign n20149 = ~n20147 & n20148;
  assign n20150 = pi39 & ~n20149;
  assign n20151 = ~n20145 & n20150;
  assign n20152 = ~pi38 & ~n20141;
  assign n20153 = ~n20151 & n20152;
  assign n20154 = ~pi701 & ~n20137;
  assign n20155 = ~n20153 & n20154;
  assign n20156 = pi150 & ~n16216;
  assign n20157 = n16228 & ~n20126;
  assign n20158 = ~n20156 & ~n20157;
  assign n20159 = pi38 & ~n20158;
  assign n20160 = ~pi150 & n19891;
  assign n20161 = pi150 & ~n19916;
  assign n20162 = ~pi751 & ~n20161;
  assign n20163 = ~n20160 & n20162;
  assign n20164 = ~pi150 & pi751;
  assign n20165 = ~n16212 & n20164;
  assign n20166 = ~n20163 & ~n20165;
  assign n20167 = pi39 & ~n20166;
  assign n20168 = pi751 & n16057;
  assign n20169 = ~n20138 & ~n20168;
  assign n20170 = n19876 & n20169;
  assign n20171 = ~pi38 & ~n20170;
  assign n20172 = ~n20167 & n20171;
  assign n20173 = pi701 & ~n20159;
  assign n20174 = ~n20172 & n20173;
  assign n20175 = ~n20155 & ~n20174;
  assign n20176 = n9830 & ~n20175;
  assign n20177 = ~pi832 & ~n20132;
  assign n20178 = ~n20176 & n20177;
  assign po307 = ~n20131 & ~n20178;
  assign n20180 = ~pi151 & ~n2923;
  assign n20181 = ~pi745 & pi947;
  assign n20182 = ~pi723 & n19798;
  assign n20183 = ~n20181 & ~n20182;
  assign n20184 = n2923 & ~n20183;
  assign n20185 = pi832 & ~n20180;
  assign n20186 = ~n20184 & n20185;
  assign n20187 = ~pi151 & ~n9830;
  assign n20188 = pi151 & ~n16216;
  assign n20189 = n16228 & ~n20181;
  assign n20190 = ~n20188 & ~n20189;
  assign n20191 = pi38 & ~n20190;
  assign n20192 = ~pi151 & ~n16057;
  assign n20193 = ~pi745 & n19903;
  assign n20194 = ~n20192 & ~n20193;
  assign n20195 = ~pi39 & ~n20194;
  assign n20196 = ~pi745 & ~n16191;
  assign n20197 = ~pi151 & ~n16212;
  assign n20198 = ~n20196 & n20197;
  assign n20199 = ~pi151 & ~n16063;
  assign n20200 = n19912 & ~n20199;
  assign n20201 = ~n3302 & ~n16192;
  assign n20202 = pi151 & n20201;
  assign n20203 = ~n16198 & ~n20202;
  assign n20204 = ~n20200 & n20203;
  assign n20205 = n19881 & n20204;
  assign n20206 = ~n16207 & ~n19883;
  assign n20207 = ~pi151 & n20206;
  assign n20208 = ~n16203 & ~n20207;
  assign n20209 = n19945 & ~n20208;
  assign n20210 = pi299 & ~n20209;
  assign n20211 = ~n20205 & n20210;
  assign n20212 = ~pi745 & ~n19905;
  assign n20213 = ~n20211 & n20212;
  assign n20214 = ~n20198 & ~n20213;
  assign n20215 = pi39 & ~n20214;
  assign n20216 = ~pi38 & ~n20195;
  assign n20217 = ~n20215 & n20216;
  assign n20218 = pi723 & ~n20191;
  assign n20219 = ~n20217 & n20218;
  assign n20220 = ~pi151 & ~n16228;
  assign n20221 = ~n19798 & ~n20181;
  assign n20222 = n16228 & ~n20221;
  assign n20223 = pi38 & ~n20220;
  assign n20224 = ~n20222 & n20223;
  assign n20225 = n19959 & n20194;
  assign n20226 = pi215 & ~n20208;
  assign n20227 = n19949 & ~n20199;
  assign n20228 = n20203 & ~n20227;
  assign n20229 = n19932 & n20228;
  assign n20230 = ~n20226 & ~n20229;
  assign n20231 = ~n19907 & ~n20230;
  assign n20232 = pi299 & ~n20231;
  assign n20233 = ~pi151 & ~n16190;
  assign n20234 = n19955 & ~n20233;
  assign n20235 = ~n20232 & ~n20234;
  assign n20236 = pi745 & ~n20235;
  assign n20237 = ~n6220 & n16190;
  assign n20238 = ~n20233 & ~n20237;
  assign n20239 = ~pi299 & ~n20238;
  assign n20240 = ~n6220 & n16063;
  assign n20241 = n20227 & ~n20240;
  assign n20242 = ~pi215 & ~n20241;
  assign n20243 = n20203 & n20242;
  assign n20244 = ~n20226 & ~n20243;
  assign n20245 = pi299 & ~n20244;
  assign n20246 = ~pi745 & ~n20245;
  assign n20247 = ~n20239 & n20246;
  assign n20248 = ~n20236 & ~n20247;
  assign n20249 = pi39 & ~n20248;
  assign n20250 = ~n20225 & ~n20249;
  assign n20251 = ~pi38 & ~n20250;
  assign n20252 = ~pi723 & ~n20224;
  assign n20253 = ~n20251 & n20252;
  assign n20254 = ~n20219 & ~n20253;
  assign n20255 = n9830 & ~n20254;
  assign n20256 = ~pi832 & ~n20187;
  assign n20257 = ~n20255 & n20256;
  assign po308 = ~n20186 & ~n20257;
  assign n20259 = ~pi152 & ~n9830;
  assign n20260 = pi759 & pi947;
  assign n20261 = n16228 & ~n20260;
  assign n20262 = ~n19798 & n20261;
  assign n20263 = ~pi152 & ~n16228;
  assign n20264 = pi38 & ~n20263;
  assign n20265 = ~n20262 & n20264;
  assign n20266 = pi152 & ~n16057;
  assign n20267 = n16057 & n20260;
  assign n20268 = ~pi39 & ~n20266;
  assign n20269 = ~n20267 & n20268;
  assign n20270 = ~n19958 & n20269;
  assign n20271 = ~pi152 & ~n16203;
  assign n20272 = n19884 & ~n20271;
  assign n20273 = ~n19798 & ~n19983;
  assign n20274 = n20272 & ~n20273;
  assign n20275 = pi152 & n19930;
  assign n20276 = n19946 & ~n20275;
  assign n20277 = pi152 & ~n16063;
  assign n20278 = ~n20240 & ~n20277;
  assign n20279 = n3302 & n20278;
  assign n20280 = ~pi215 & ~n20279;
  assign n20281 = ~n19929 & n20280;
  assign n20282 = ~n20276 & n20281;
  assign n20283 = pi299 & ~n20274;
  assign n20284 = ~n20282 & n20283;
  assign n20285 = ~n19948 & ~n20277;
  assign n20286 = n2608 & ~n20285;
  assign n20287 = ~pi152 & n16186;
  assign n20288 = ~n16186 & ~n19798;
  assign n20289 = ~n2608 & ~n20288;
  assign n20290 = ~n20287 & n20289;
  assign n20291 = ~n20286 & ~n20290;
  assign n20292 = ~pi223 & ~n20291;
  assign n20293 = ~n16124 & ~n19798;
  assign n20294 = pi223 & ~n20293;
  assign n20295 = ~pi152 & n16124;
  assign n20296 = n20294 & ~n20295;
  assign n20297 = ~pi299 & ~n20296;
  assign n20298 = ~n20292 & n20297;
  assign n20299 = ~pi759 & ~n20284;
  assign n20300 = ~n20298 & n20299;
  assign n20301 = ~n16192 & n20276;
  assign n20302 = n20280 & ~n20301;
  assign n20303 = pi299 & ~n20272;
  assign n20304 = ~n20302 & n20303;
  assign n20305 = n2608 & n20278;
  assign n20306 = ~pi947 & ~n16186;
  assign n20307 = ~n2608 & ~n20306;
  assign n20308 = ~n20287 & n20307;
  assign n20309 = ~n2608 & n6220;
  assign n20310 = ~n16187 & ~n20309;
  assign n20311 = ~n20308 & ~n20310;
  assign n20312 = ~pi223 & ~n20305;
  assign n20313 = ~n20311 & n20312;
  assign n20314 = ~pi947 & ~n16124;
  assign n20315 = pi223 & ~n20314;
  assign n20316 = ~n20295 & n20315;
  assign n20317 = ~pi299 & ~n20316;
  assign n20318 = ~n20296 & n20317;
  assign n20319 = ~n20313 & n20318;
  assign n20320 = pi759 & ~n20319;
  assign n20321 = ~n20304 & n20320;
  assign n20322 = pi39 & ~n20300;
  assign n20323 = ~n20321 & n20322;
  assign n20324 = ~pi38 & ~n20270;
  assign n20325 = ~n20323 & n20324;
  assign n20326 = pi696 & ~n20265;
  assign n20327 = ~n20325 & n20326;
  assign n20328 = ~pi152 & ~n16216;
  assign n20329 = pi38 & ~n20261;
  assign n20330 = ~n20328 & n20329;
  assign n20331 = ~n19911 & ~n20277;
  assign n20332 = n2608 & ~n20331;
  assign n20333 = ~n20308 & ~n20332;
  assign n20334 = ~pi223 & ~n20333;
  assign n20335 = n20317 & ~n20334;
  assign n20336 = pi152 & n19885;
  assign n20337 = n3302 & n20331;
  assign n20338 = n19881 & ~n20337;
  assign n20339 = ~n20301 & n20338;
  assign n20340 = n19908 & ~n20336;
  assign n20341 = ~n20339 & n20340;
  assign n20342 = pi759 & ~n20335;
  assign n20343 = ~n20341 & n20342;
  assign n20344 = ~pi759 & ~n16212;
  assign n20345 = pi152 & n20344;
  assign n20346 = pi39 & ~n20343;
  assign n20347 = ~n20345 & n20346;
  assign n20348 = ~pi38 & ~n20269;
  assign n20349 = ~n20347 & n20348;
  assign n20350 = ~pi696 & ~n20330;
  assign n20351 = ~n20349 & n20350;
  assign n20352 = ~n20327 & ~n20351;
  assign n20353 = n9830 & ~n20352;
  assign n20354 = ~pi832 & ~n20259;
  assign n20355 = ~n20353 & n20354;
  assign n20356 = ~pi152 & ~n2923;
  assign n20357 = pi696 & n19798;
  assign n20358 = n2923 & ~n20260;
  assign n20359 = ~n20357 & n20358;
  assign n20360 = pi832 & ~n20356;
  assign n20361 = ~n20359 & n20360;
  assign po309 = n20355 | n20361;
  assign n20363 = pi700 & n19798;
  assign n20364 = pi766 & pi947;
  assign n20365 = n2923 & ~n20364;
  assign n20366 = ~n20363 & n20365;
  assign n20367 = pi153 & ~n2923;
  assign n20368 = pi832 & ~n20367;
  assign n20369 = ~n20366 & n20368;
  assign n20370 = pi57 & pi153;
  assign n20371 = ~pi153 & ~n20005;
  assign n20372 = pi153 & ~n16216;
  assign n20373 = n16228 & ~n20364;
  assign n20374 = pi38 & ~n20373;
  assign n20375 = ~n20372 & n20374;
  assign n20376 = ~pi153 & ~pi766;
  assign n20377 = ~n16212 & n20376;
  assign n20378 = ~pi153 & ~n16190;
  assign n20379 = n19905 & ~n20378;
  assign n20380 = pi153 & ~n16203;
  assign n20381 = n19884 & ~n20380;
  assign n20382 = ~n19883 & n20381;
  assign n20383 = ~pi153 & ~n16063;
  assign n20384 = n19912 & ~n20383;
  assign n20385 = pi153 & n20201;
  assign n20386 = ~n16198 & ~n20385;
  assign n20387 = ~n20384 & n20386;
  assign n20388 = n19881 & n20387;
  assign n20389 = pi299 & ~n20382;
  assign n20390 = ~n20388 & n20389;
  assign n20391 = pi766 & ~n20390;
  assign n20392 = ~n20379 & n20391;
  assign n20393 = pi39 & ~n20377;
  assign n20394 = ~n20392 & n20393;
  assign n20395 = ~pi153 & ~n16057;
  assign n20396 = ~pi766 & n17347;
  assign n20397 = ~n19904 & ~n20396;
  assign n20398 = ~n20395 & ~n20397;
  assign n20399 = ~pi38 & ~n20398;
  assign n20400 = ~n20394 & n20399;
  assign n20401 = ~n20375 & ~n20400;
  assign n20402 = ~pi700 & ~n20401;
  assign n20403 = ~n19958 & n20398;
  assign n20404 = n19955 & ~n20378;
  assign n20405 = n19983 & ~n20381;
  assign n20406 = n19949 & ~n20383;
  assign n20407 = ~n19931 & ~n20406;
  assign n20408 = n20386 & n20407;
  assign n20409 = ~pi215 & ~n20408;
  assign n20410 = ~n19907 & ~n20405;
  assign n20411 = ~n20409 & n20410;
  assign n20412 = pi299 & ~n20411;
  assign n20413 = ~n20404 & ~n20412;
  assign n20414 = ~pi766 & ~n20413;
  assign n20415 = ~n20237 & ~n20378;
  assign n20416 = ~pi299 & ~n20415;
  assign n20417 = ~n19947 & n20384;
  assign n20418 = ~pi215 & ~n20417;
  assign n20419 = n20386 & n20418;
  assign n20420 = ~n20381 & ~n20419;
  assign n20421 = pi299 & ~n20420;
  assign n20422 = pi766 & ~n20421;
  assign n20423 = ~n20416 & n20422;
  assign n20424 = ~n20414 & ~n20423;
  assign n20425 = pi39 & ~n20424;
  assign n20426 = ~n20403 & ~n20425;
  assign n20427 = ~pi38 & ~n20426;
  assign n20428 = ~pi153 & ~n16228;
  assign n20429 = ~n19798 & ~n20364;
  assign n20430 = n16228 & ~n20429;
  assign n20431 = pi38 & ~n20428;
  assign n20432 = ~n20430 & n20431;
  assign n20433 = pi700 & ~n20432;
  assign n20434 = ~n20427 & n20433;
  assign n20435 = ~n20402 & ~n20434;
  assign n20436 = n20005 & ~n20435;
  assign n20437 = ~pi57 & ~n20371;
  assign n20438 = ~n20436 & n20437;
  assign n20439 = ~pi832 & ~n20370;
  assign n20440 = ~n20438 & n20439;
  assign po310 = n20369 | n20440;
  assign n20442 = ~pi154 & ~n2923;
  assign n20443 = ~pi742 & pi947;
  assign n20444 = ~pi704 & n19798;
  assign n20445 = ~n20443 & ~n20444;
  assign n20446 = n2923 & ~n20445;
  assign n20447 = pi832 & ~n20442;
  assign n20448 = ~n20446 & n20447;
  assign n20449 = ~pi154 & ~n9830;
  assign n20450 = ~pi154 & ~n16228;
  assign n20451 = n19927 & ~n20450;
  assign n20452 = ~pi154 & ~n16057;
  assign n20453 = n19959 & ~n20452;
  assign n20454 = ~pi154 & n19939;
  assign n20455 = pi154 & n19956;
  assign n20456 = pi39 & ~n20455;
  assign n20457 = ~n20454 & n20456;
  assign n20458 = ~n20453 & ~n20457;
  assign n20459 = ~pi38 & ~n20458;
  assign n20460 = pi742 & ~n20451;
  assign n20461 = ~n20459 & n20460;
  assign n20462 = n19969 & ~n20450;
  assign n20463 = ~n19978 & n20453;
  assign n20464 = pi154 & ~n19989;
  assign n20465 = ~pi154 & ~n19976;
  assign n20466 = pi39 & ~n20464;
  assign n20467 = ~n20465 & n20466;
  assign n20468 = ~n20463 & ~n20467;
  assign n20469 = ~pi38 & ~n20468;
  assign n20470 = ~pi742 & ~n20462;
  assign n20471 = ~n20469 & n20470;
  assign n20472 = ~pi704 & ~n20471;
  assign n20473 = ~n20461 & n20472;
  assign n20474 = ~pi154 & ~n16216;
  assign n20475 = ~n19902 & ~n20474;
  assign n20476 = n19904 & ~n20452;
  assign n20477 = pi154 & n19916;
  assign n20478 = ~pi154 & ~n19891;
  assign n20479 = pi39 & ~n20477;
  assign n20480 = ~n20478 & n20479;
  assign n20481 = ~n20476 & ~n20480;
  assign n20482 = ~pi38 & ~n20481;
  assign n20483 = ~pi742 & ~n20475;
  assign n20484 = ~n20482 & n20483;
  assign n20485 = ~pi154 & pi742;
  assign n20486 = ~n16218 & n20485;
  assign n20487 = pi704 & ~n20486;
  assign n20488 = ~n20484 & n20487;
  assign n20489 = n9830 & ~n20473;
  assign n20490 = ~n20488 & n20489;
  assign n20491 = ~pi832 & ~n20449;
  assign n20492 = ~n20490 & n20491;
  assign po311 = ~n20448 & ~n20492;
  assign n20494 = ~pi757 & n19920;
  assign n20495 = pi686 & ~n20494;
  assign n20496 = ~pi38 & ~n19991;
  assign n20497 = ~n19969 & ~n20496;
  assign n20498 = ~pi757 & n20497;
  assign n20499 = ~pi38 & ~n19960;
  assign n20500 = ~n19927 & ~n20499;
  assign n20501 = pi757 & n20500;
  assign n20502 = ~pi686 & ~n20498;
  assign n20503 = ~n20501 & n20502;
  assign n20504 = n9830 & ~n20495;
  assign n20505 = ~n20503 & n20504;
  assign n20506 = pi155 & ~n20505;
  assign n20507 = ~pi38 & ~n19981;
  assign n20508 = pi38 & n19966;
  assign n20509 = ~n20507 & ~n20508;
  assign n20510 = ~pi757 & n20509;
  assign n20511 = ~pi38 & ~n19943;
  assign n20512 = n18596 & ~n19798;
  assign n20513 = n16065 & n20512;
  assign n20514 = ~n20511 & ~n20513;
  assign n20515 = pi757 & n20514;
  assign n20516 = ~pi686 & ~n20510;
  assign n20517 = ~n20515 & n20516;
  assign n20518 = ~pi757 & n19897;
  assign n20519 = pi757 & ~n16218;
  assign n20520 = pi686 & ~n20519;
  assign n20521 = ~n20518 & n20520;
  assign n20522 = ~n20517 & ~n20521;
  assign n20523 = ~pi155 & n9830;
  assign n20524 = ~n20522 & n20523;
  assign n20525 = ~n20506 & ~n20524;
  assign n20526 = ~pi832 & ~n20525;
  assign n20527 = ~pi155 & ~n2923;
  assign n20528 = ~pi757 & pi947;
  assign n20529 = ~pi686 & n19798;
  assign n20530 = ~n20528 & ~n20529;
  assign n20531 = n2923 & ~n20530;
  assign n20532 = pi832 & ~n20527;
  assign n20533 = ~n20531 & n20532;
  assign po312 = ~n20526 & ~n20533;
  assign n20535 = ~pi156 & ~n2923;
  assign n20536 = ~pi741 & pi947;
  assign n20537 = ~pi724 & n19798;
  assign n20538 = ~n20536 & ~n20537;
  assign n20539 = n2923 & ~n20538;
  assign n20540 = pi832 & ~n20535;
  assign n20541 = ~n20539 & n20540;
  assign n20542 = ~pi741 & ~n20509;
  assign n20543 = pi741 & ~n20514;
  assign n20544 = ~pi724 & ~n20542;
  assign n20545 = ~n20543 & n20544;
  assign n20546 = ~pi741 & ~n19897;
  assign n20547 = pi741 & n16218;
  assign n20548 = pi724 & ~n20547;
  assign n20549 = ~n20546 & n20548;
  assign n20550 = n9830 & ~n20545;
  assign n20551 = ~n20549 & n20550;
  assign n20552 = ~pi156 & ~n20551;
  assign n20553 = ~pi741 & ~n20497;
  assign n20554 = pi741 & ~n20500;
  assign n20555 = ~pi724 & ~n20553;
  assign n20556 = ~n20554 & n20555;
  assign n20557 = pi724 & ~pi741;
  assign n20558 = n19920 & n20557;
  assign n20559 = ~n20556 & ~n20558;
  assign n20560 = pi156 & n9830;
  assign n20561 = ~n20559 & n20560;
  assign n20562 = ~pi832 & ~n20561;
  assign n20563 = ~n20552 & n20562;
  assign po313 = ~n20541 & ~n20563;
  assign n20565 = ~pi157 & ~n2923;
  assign n20566 = ~pi760 & pi947;
  assign n20567 = ~pi688 & n19798;
  assign n20568 = ~n20566 & ~n20567;
  assign n20569 = n2923 & ~n20568;
  assign n20570 = pi832 & ~n20565;
  assign n20571 = ~n20569 & n20570;
  assign n20572 = ~pi157 & ~n9830;
  assign n20573 = n16228 & ~n20566;
  assign n20574 = pi157 & ~n16216;
  assign n20575 = pi38 & ~n20573;
  assign n20576 = ~n20574 & n20575;
  assign n20577 = ~pi157 & pi760;
  assign n20578 = ~n16212 & n20577;
  assign n20579 = ~pi157 & ~n16190;
  assign n20580 = n19905 & ~n20579;
  assign n20581 = ~pi157 & ~n19886;
  assign n20582 = ~n12970 & ~n19915;
  assign n20583 = ~n20581 & ~n20582;
  assign n20584 = ~pi760 & ~n20580;
  assign n20585 = ~n20583 & n20584;
  assign n20586 = pi39 & ~n20578;
  assign n20587 = ~n20585 & n20586;
  assign n20588 = ~pi157 & ~n16057;
  assign n20589 = n16057 & n20566;
  assign n20590 = ~pi39 & ~n20588;
  assign n20591 = ~n20589 & n20590;
  assign n20592 = ~pi38 & ~n20591;
  assign n20593 = ~n20587 & n20592;
  assign n20594 = ~n20576 & ~n20593;
  assign n20595 = pi688 & ~n20594;
  assign n20596 = ~n19958 & n20591;
  assign n20597 = pi760 & n19956;
  assign n20598 = ~pi760 & ~n19989;
  assign n20599 = pi157 & ~n20597;
  assign n20600 = ~n20598 & n20599;
  assign n20601 = pi760 & n19939;
  assign n20602 = ~pi760 & ~n19976;
  assign n20603 = ~pi157 & ~n20602;
  assign n20604 = ~n20601 & n20603;
  assign n20605 = ~n20600 & ~n20604;
  assign n20606 = pi39 & ~n20605;
  assign n20607 = ~n20596 & ~n20606;
  assign n20608 = ~pi38 & ~n20607;
  assign n20609 = ~pi157 & ~n16228;
  assign n20610 = ~n19798 & ~n20566;
  assign n20611 = n16228 & ~n20610;
  assign n20612 = pi38 & ~n20609;
  assign n20613 = ~n20611 & n20612;
  assign n20614 = ~pi688 & ~n20613;
  assign n20615 = ~n20608 & n20614;
  assign n20616 = ~n20595 & ~n20615;
  assign n20617 = n9830 & ~n20616;
  assign n20618 = ~pi832 & ~n20572;
  assign n20619 = ~n20617 & n20618;
  assign po314 = ~n20571 & ~n20619;
  assign n20621 = ~pi158 & ~n2923;
  assign n20622 = ~pi753 & pi947;
  assign n20623 = ~pi702 & n19798;
  assign n20624 = ~n20622 & ~n20623;
  assign n20625 = n2923 & ~n20624;
  assign n20626 = pi832 & ~n20621;
  assign n20627 = ~n20625 & n20626;
  assign n20628 = ~pi158 & ~n9830;
  assign n20629 = ~pi158 & ~n16228;
  assign n20630 = ~n19798 & ~n20622;
  assign n20631 = n16228 & ~n20630;
  assign n20632 = pi38 & ~n20629;
  assign n20633 = ~n20631 & n20632;
  assign n20634 = pi158 & ~n16057;
  assign n20635 = n19941 & ~n20622;
  assign n20636 = ~pi39 & ~n20634;
  assign n20637 = ~n20635 & n20636;
  assign n20638 = ~pi158 & n19939;
  assign n20639 = pi158 & n19956;
  assign n20640 = pi753 & ~n20639;
  assign n20641 = ~n20638 & n20640;
  assign n20642 = pi158 & ~n19989;
  assign n20643 = ~pi158 & ~n19976;
  assign n20644 = ~pi753 & ~n20642;
  assign n20645 = ~n20643 & n20644;
  assign n20646 = pi39 & ~n20645;
  assign n20647 = ~n20641 & n20646;
  assign n20648 = ~pi38 & ~n20637;
  assign n20649 = ~n20647 & n20648;
  assign n20650 = ~pi702 & ~n20633;
  assign n20651 = ~n20649 & n20650;
  assign n20652 = pi158 & ~n16216;
  assign n20653 = n16228 & ~n20622;
  assign n20654 = ~n20652 & ~n20653;
  assign n20655 = pi38 & ~n20654;
  assign n20656 = ~pi158 & n19891;
  assign n20657 = pi158 & ~n19916;
  assign n20658 = ~pi753 & ~n20657;
  assign n20659 = ~n20656 & n20658;
  assign n20660 = ~pi158 & pi753;
  assign n20661 = ~n16212 & n20660;
  assign n20662 = ~n20659 & ~n20661;
  assign n20663 = pi39 & ~n20662;
  assign n20664 = pi753 & n16057;
  assign n20665 = ~n20634 & ~n20664;
  assign n20666 = n19876 & n20665;
  assign n20667 = ~pi38 & ~n20666;
  assign n20668 = ~n20663 & n20667;
  assign n20669 = pi702 & ~n20655;
  assign n20670 = ~n20668 & n20669;
  assign n20671 = ~n20651 & ~n20670;
  assign n20672 = n9830 & ~n20671;
  assign n20673 = ~pi832 & ~n20628;
  assign n20674 = ~n20672 & n20673;
  assign po315 = ~n20627 & ~n20674;
  assign n20676 = ~pi159 & ~n2923;
  assign n20677 = ~pi754 & pi947;
  assign n20678 = ~pi709 & n19798;
  assign n20679 = ~n20677 & ~n20678;
  assign n20680 = n2923 & ~n20679;
  assign n20681 = pi832 & ~n20676;
  assign n20682 = ~n20680 & n20681;
  assign n20683 = ~pi159 & ~n9830;
  assign n20684 = ~pi159 & ~n16228;
  assign n20685 = ~n19798 & ~n20677;
  assign n20686 = n16228 & ~n20685;
  assign n20687 = pi38 & ~n20684;
  assign n20688 = ~n20686 & n20687;
  assign n20689 = pi159 & ~n16057;
  assign n20690 = n19941 & ~n20677;
  assign n20691 = ~pi39 & ~n20689;
  assign n20692 = ~n20690 & n20691;
  assign n20693 = ~pi159 & n19939;
  assign n20694 = pi159 & n19956;
  assign n20695 = pi754 & ~n20694;
  assign n20696 = ~n20693 & n20695;
  assign n20697 = pi159 & ~n19989;
  assign n20698 = ~pi159 & ~n19976;
  assign n20699 = ~pi754 & ~n20697;
  assign n20700 = ~n20698 & n20699;
  assign n20701 = pi39 & ~n20700;
  assign n20702 = ~n20696 & n20701;
  assign n20703 = ~pi38 & ~n20692;
  assign n20704 = ~n20702 & n20703;
  assign n20705 = ~pi709 & ~n20688;
  assign n20706 = ~n20704 & n20705;
  assign n20707 = pi159 & ~n16216;
  assign n20708 = n16228 & ~n20677;
  assign n20709 = ~n20707 & ~n20708;
  assign n20710 = pi38 & ~n20709;
  assign n20711 = ~pi159 & n19891;
  assign n20712 = pi159 & ~n19916;
  assign n20713 = ~pi754 & ~n20712;
  assign n20714 = ~n20711 & n20713;
  assign n20715 = ~pi159 & pi754;
  assign n20716 = ~n16212 & n20715;
  assign n20717 = ~n20714 & ~n20716;
  assign n20718 = pi39 & ~n20717;
  assign n20719 = pi754 & n16057;
  assign n20720 = ~n20689 & ~n20719;
  assign n20721 = n19876 & n20720;
  assign n20722 = ~pi38 & ~n20721;
  assign n20723 = ~n20718 & n20722;
  assign n20724 = pi709 & ~n20710;
  assign n20725 = ~n20723 & n20724;
  assign n20726 = ~n20706 & ~n20725;
  assign n20727 = n9830 & ~n20726;
  assign n20728 = ~pi832 & ~n20683;
  assign n20729 = ~n20727 & n20728;
  assign po316 = ~n20682 & ~n20729;
  assign n20731 = ~pi160 & ~n2923;
  assign n20732 = ~pi756 & pi947;
  assign n20733 = ~pi734 & n19798;
  assign n20734 = ~n20732 & ~n20733;
  assign n20735 = n2923 & ~n20734;
  assign n20736 = pi832 & ~n20731;
  assign n20737 = ~n20735 & n20736;
  assign n20738 = ~pi160 & ~n9830;
  assign n20739 = n16228 & ~n20732;
  assign n20740 = pi160 & ~n16216;
  assign n20741 = pi38 & ~n20739;
  assign n20742 = ~n20740 & n20741;
  assign n20743 = ~pi160 & pi756;
  assign n20744 = ~n16212 & n20743;
  assign n20745 = ~pi160 & ~n16190;
  assign n20746 = n19905 & ~n20745;
  assign n20747 = pi160 & ~n20042;
  assign n20748 = ~pi160 & ~n19886;
  assign n20749 = pi299 & ~n20747;
  assign n20750 = ~n20748 & n20749;
  assign n20751 = ~pi756 & ~n20746;
  assign n20752 = ~n20750 & n20751;
  assign n20753 = pi39 & ~n20744;
  assign n20754 = ~n20752 & n20753;
  assign n20755 = ~pi160 & ~n16057;
  assign n20756 = n16057 & n20732;
  assign n20757 = ~pi39 & ~n20755;
  assign n20758 = ~n20756 & n20757;
  assign n20759 = ~pi38 & ~n20758;
  assign n20760 = ~n20754 & n20759;
  assign n20761 = ~n20742 & ~n20760;
  assign n20762 = pi734 & ~n20761;
  assign n20763 = ~n19958 & n20758;
  assign n20764 = pi160 & ~n20017;
  assign n20765 = ~pi160 & n19936;
  assign n20766 = ~n19938 & ~n20764;
  assign n20767 = ~n20765 & n20766;
  assign n20768 = pi756 & ~n20767;
  assign n20769 = ~pi160 & ~n19976;
  assign n20770 = pi160 & ~n19989;
  assign n20771 = ~pi756 & ~n20770;
  assign n20772 = ~n20769 & n20771;
  assign n20773 = ~n20768 & ~n20772;
  assign n20774 = pi39 & ~n20773;
  assign n20775 = ~n20763 & ~n20774;
  assign n20776 = ~pi38 & ~n20775;
  assign n20777 = ~pi160 & ~n16228;
  assign n20778 = ~n19798 & ~n20732;
  assign n20779 = n16228 & ~n20778;
  assign n20780 = pi38 & ~n20777;
  assign n20781 = ~n20779 & n20780;
  assign n20782 = ~pi734 & ~n20781;
  assign n20783 = ~n20776 & n20782;
  assign n20784 = ~n20762 & ~n20783;
  assign n20785 = n9830 & ~n20784;
  assign n20786 = ~pi832 & ~n20738;
  assign n20787 = ~n20785 & n20786;
  assign po317 = ~n20737 & ~n20787;
  assign n20789 = ~pi161 & ~n9830;
  assign n20790 = pi758 & pi947;
  assign n20791 = n16228 & ~n20790;
  assign n20792 = ~n19798 & n20791;
  assign n20793 = ~pi161 & ~n16228;
  assign n20794 = pi38 & ~n20793;
  assign n20795 = ~n20792 & n20794;
  assign n20796 = pi161 & ~n16057;
  assign n20797 = n16057 & n20790;
  assign n20798 = ~pi39 & ~n20796;
  assign n20799 = ~n20797 & n20798;
  assign n20800 = ~n19958 & n20799;
  assign n20801 = ~pi161 & ~n16203;
  assign n20802 = n19884 & ~n20801;
  assign n20803 = ~n20273 & n20802;
  assign n20804 = pi161 & n19930;
  assign n20805 = n19946 & ~n20804;
  assign n20806 = pi161 & ~n16063;
  assign n20807 = ~n20240 & ~n20806;
  assign n20808 = n3302 & n20807;
  assign n20809 = ~pi215 & ~n20808;
  assign n20810 = ~n19929 & n20809;
  assign n20811 = ~n20805 & n20810;
  assign n20812 = pi299 & ~n20803;
  assign n20813 = ~n20811 & n20812;
  assign n20814 = ~n19948 & ~n20806;
  assign n20815 = n2608 & ~n20814;
  assign n20816 = ~pi161 & n16186;
  assign n20817 = n20289 & ~n20816;
  assign n20818 = ~n20815 & ~n20817;
  assign n20819 = ~pi223 & ~n20818;
  assign n20820 = ~pi161 & n16124;
  assign n20821 = n20294 & ~n20820;
  assign n20822 = ~pi299 & ~n20821;
  assign n20823 = ~n20819 & n20822;
  assign n20824 = ~pi758 & ~n20813;
  assign n20825 = ~n20823 & n20824;
  assign n20826 = ~n16192 & n20805;
  assign n20827 = n20809 & ~n20826;
  assign n20828 = pi299 & ~n20802;
  assign n20829 = ~n20827 & n20828;
  assign n20830 = n2608 & n20807;
  assign n20831 = n20307 & ~n20816;
  assign n20832 = ~n20310 & ~n20831;
  assign n20833 = ~pi223 & ~n20830;
  assign n20834 = ~n20832 & n20833;
  assign n20835 = n20315 & ~n20820;
  assign n20836 = ~pi299 & ~n20835;
  assign n20837 = ~n20821 & n20836;
  assign n20838 = ~n20834 & n20837;
  assign n20839 = pi758 & ~n20838;
  assign n20840 = ~n20829 & n20839;
  assign n20841 = pi39 & ~n20825;
  assign n20842 = ~n20840 & n20841;
  assign n20843 = ~pi38 & ~n20800;
  assign n20844 = ~n20842 & n20843;
  assign n20845 = pi736 & ~n20795;
  assign n20846 = ~n20844 & n20845;
  assign n20847 = ~pi161 & ~n16216;
  assign n20848 = pi38 & ~n20791;
  assign n20849 = ~n20847 & n20848;
  assign n20850 = ~n19911 & ~n20806;
  assign n20851 = n2608 & ~n20850;
  assign n20852 = ~n20831 & ~n20851;
  assign n20853 = ~pi223 & ~n20852;
  assign n20854 = n20836 & ~n20853;
  assign n20855 = pi161 & n19885;
  assign n20856 = n3302 & n20850;
  assign n20857 = n19881 & ~n20856;
  assign n20858 = ~n20826 & n20857;
  assign n20859 = n19908 & ~n20855;
  assign n20860 = ~n20858 & n20859;
  assign n20861 = pi758 & ~n20854;
  assign n20862 = ~n20860 & n20861;
  assign n20863 = pi161 & n19104;
  assign n20864 = pi39 & ~n20862;
  assign n20865 = ~n20863 & n20864;
  assign n20866 = ~pi38 & ~n20799;
  assign n20867 = ~n20865 & n20866;
  assign n20868 = ~pi736 & ~n20849;
  assign n20869 = ~n20867 & n20868;
  assign n20870 = ~n20846 & ~n20869;
  assign n20871 = n9830 & ~n20870;
  assign n20872 = ~pi832 & ~n20789;
  assign n20873 = ~n20871 & n20872;
  assign n20874 = ~pi161 & ~n2923;
  assign n20875 = pi736 & n19798;
  assign n20876 = n2923 & ~n20790;
  assign n20877 = ~n20875 & n20876;
  assign n20878 = pi832 & ~n20874;
  assign n20879 = ~n20877 & n20878;
  assign po318 = n20873 | n20879;
  assign n20881 = ~pi162 & ~n9830;
  assign n20882 = ~pi761 & pi947;
  assign n20883 = n16228 & ~n20882;
  assign n20884 = pi162 & ~n16216;
  assign n20885 = pi38 & ~n20883;
  assign n20886 = ~n20884 & n20885;
  assign n20887 = ~pi162 & ~n16057;
  assign n20888 = n16057 & n20882;
  assign n20889 = ~pi39 & ~n20887;
  assign n20890 = ~n20888 & n20889;
  assign n20891 = ~pi162 & ~n16212;
  assign n20892 = pi761 & ~n20891;
  assign n20893 = ~pi761 & n19888;
  assign n20894 = ~pi162 & ~n20893;
  assign n20895 = n14257 & ~n20042;
  assign n20896 = ~n19890 & ~n20895;
  assign n20897 = ~n20894 & n20896;
  assign n20898 = ~n20892 & ~n20897;
  assign n20899 = pi39 & ~n20898;
  assign n20900 = ~pi38 & ~n20890;
  assign n20901 = ~n20899 & n20900;
  assign n20902 = ~n20886 & ~n20901;
  assign n20903 = pi738 & ~n20902;
  assign n20904 = ~n19958 & n20890;
  assign n20905 = ~n14257 & ~n19939;
  assign n20906 = pi162 & ~n20017;
  assign n20907 = ~n20905 & ~n20906;
  assign n20908 = pi761 & ~n20907;
  assign n20909 = pi162 & ~n19989;
  assign n20910 = ~pi162 & ~n19976;
  assign n20911 = ~pi761 & ~n20909;
  assign n20912 = ~n20910 & n20911;
  assign n20913 = ~n20908 & ~n20912;
  assign n20914 = pi39 & ~n20913;
  assign n20915 = ~n20904 & ~n20914;
  assign n20916 = ~pi38 & ~n20915;
  assign n20917 = ~pi162 & ~n16228;
  assign n20918 = ~n19798 & ~n20882;
  assign n20919 = n16228 & ~n20918;
  assign n20920 = pi38 & ~n20917;
  assign n20921 = ~n20919 & n20920;
  assign n20922 = ~pi738 & ~n20921;
  assign n20923 = ~n20916 & n20922;
  assign n20924 = ~n20903 & ~n20923;
  assign n20925 = n9830 & ~n20924;
  assign n20926 = ~pi832 & ~n20881;
  assign n20927 = ~n20925 & n20926;
  assign n20928 = ~pi162 & ~n2923;
  assign n20929 = ~pi738 & n19798;
  assign n20930 = ~n20882 & ~n20929;
  assign n20931 = n2923 & ~n20930;
  assign n20932 = pi832 & ~n20928;
  assign n20933 = ~n20931 & n20932;
  assign po319 = ~n20927 & ~n20933;
  assign n20935 = ~pi163 & ~n2923;
  assign n20936 = ~pi777 & pi947;
  assign n20937 = ~pi737 & n19798;
  assign n20938 = ~n20936 & ~n20937;
  assign n20939 = n2923 & ~n20938;
  assign n20940 = pi832 & ~n20935;
  assign n20941 = ~n20939 & n20940;
  assign n20942 = ~pi163 & ~n9830;
  assign n20943 = n16228 & ~n20936;
  assign n20944 = pi163 & ~n16216;
  assign n20945 = pi38 & ~n20943;
  assign n20946 = ~n20944 & n20945;
  assign n20947 = ~pi163 & pi777;
  assign n20948 = ~n16212 & n20947;
  assign n20949 = ~pi163 & ~n16190;
  assign n20950 = n19905 & ~n20949;
  assign n20951 = ~pi163 & ~n19886;
  assign n20952 = ~n13632 & ~n19915;
  assign n20953 = ~n20951 & ~n20952;
  assign n20954 = ~pi777 & ~n20950;
  assign n20955 = ~n20953 & n20954;
  assign n20956 = pi39 & ~n20948;
  assign n20957 = ~n20955 & n20956;
  assign n20958 = ~pi163 & ~n16057;
  assign n20959 = n16057 & n20936;
  assign n20960 = ~pi39 & ~n20958;
  assign n20961 = ~n20959 & n20960;
  assign n20962 = ~pi38 & ~n20961;
  assign n20963 = ~n20957 & n20962;
  assign n20964 = ~n20946 & ~n20963;
  assign n20965 = pi737 & ~n20964;
  assign n20966 = ~n19958 & n20961;
  assign n20967 = pi163 & ~n20017;
  assign n20968 = ~pi163 & n19936;
  assign n20969 = ~n19938 & ~n20967;
  assign n20970 = ~n20968 & n20969;
  assign n20971 = pi777 & ~n20970;
  assign n20972 = ~pi163 & ~n19976;
  assign n20973 = pi163 & ~n19989;
  assign n20974 = ~pi777 & ~n20973;
  assign n20975 = ~n20972 & n20974;
  assign n20976 = ~n20971 & ~n20975;
  assign n20977 = pi39 & ~n20976;
  assign n20978 = ~n20966 & ~n20977;
  assign n20979 = ~pi38 & ~n20978;
  assign n20980 = ~pi163 & ~n16228;
  assign n20981 = ~n19798 & ~n20936;
  assign n20982 = n16228 & ~n20981;
  assign n20983 = pi38 & ~n20980;
  assign n20984 = ~n20982 & n20983;
  assign n20985 = ~pi737 & ~n20984;
  assign n20986 = ~n20979 & n20985;
  assign n20987 = ~n20965 & ~n20986;
  assign n20988 = n9830 & ~n20987;
  assign n20989 = ~pi832 & ~n20942;
  assign n20990 = ~n20988 & n20989;
  assign po320 = ~n20941 & ~n20990;
  assign n20992 = ~pi164 & ~n2923;
  assign n20993 = ~pi752 & pi947;
  assign n20994 = pi703 & n19798;
  assign n20995 = ~n20993 & ~n20994;
  assign n20996 = n2923 & ~n20995;
  assign n20997 = pi832 & ~n20992;
  assign n20998 = ~n20996 & n20997;
  assign n20999 = ~pi164 & ~n9830;
  assign n21000 = ~pi164 & ~n19966;
  assign n21001 = n19969 & ~n21000;
  assign n21002 = ~pi164 & n19981;
  assign n21003 = pi164 & n19991;
  assign n21004 = ~pi38 & ~n21003;
  assign n21005 = ~n21002 & n21004;
  assign n21006 = ~pi752 & ~n21001;
  assign n21007 = ~n21005 & n21006;
  assign n21008 = ~pi164 & ~n16228;
  assign n21009 = n19927 & ~n21008;
  assign n21010 = ~pi164 & n19943;
  assign n21011 = pi164 & n19960;
  assign n21012 = ~pi38 & ~n21011;
  assign n21013 = ~n21010 & n21012;
  assign n21014 = pi752 & ~n21009;
  assign n21015 = ~n21013 & n21014;
  assign n21016 = ~n21007 & ~n21015;
  assign n21017 = pi703 & ~n21016;
  assign n21018 = pi164 & ~n19920;
  assign n21019 = pi164 & ~n19896;
  assign n21020 = ~pi752 & ~n21019;
  assign n21021 = ~n19897 & n21020;
  assign n21022 = ~pi164 & ~n16218;
  assign n21023 = pi752 & ~n21022;
  assign n21024 = ~pi703 & ~n21018;
  assign n21025 = ~n21023 & n21024;
  assign n21026 = ~n21021 & n21025;
  assign n21027 = ~n21017 & ~n21026;
  assign n21028 = n9830 & ~n21027;
  assign n21029 = ~pi832 & ~n20999;
  assign n21030 = ~n21028 & n21029;
  assign po321 = ~n20998 & ~n21030;
  assign n21032 = ~pi165 & ~n2923;
  assign n21033 = ~pi774 & pi947;
  assign n21034 = pi687 & n19798;
  assign n21035 = ~n21033 & ~n21034;
  assign n21036 = n2923 & ~n21035;
  assign n21037 = pi832 & ~n21032;
  assign n21038 = ~n21036 & n21037;
  assign n21039 = ~pi165 & ~n9830;
  assign n21040 = ~pi165 & ~n19966;
  assign n21041 = n19969 & ~n21040;
  assign n21042 = ~pi165 & n19981;
  assign n21043 = pi165 & n19991;
  assign n21044 = ~pi38 & ~n21043;
  assign n21045 = ~n21042 & n21044;
  assign n21046 = ~pi774 & ~n21041;
  assign n21047 = ~n21045 & n21046;
  assign n21048 = ~pi165 & ~n16228;
  assign n21049 = n19927 & ~n21048;
  assign n21050 = ~pi165 & n19943;
  assign n21051 = pi165 & n19960;
  assign n21052 = ~pi38 & ~n21051;
  assign n21053 = ~n21050 & n21052;
  assign n21054 = pi774 & ~n21049;
  assign n21055 = ~n21053 & n21054;
  assign n21056 = ~n21047 & ~n21055;
  assign n21057 = pi687 & ~n21056;
  assign n21058 = pi165 & ~n19920;
  assign n21059 = pi165 & ~n19896;
  assign n21060 = ~pi774 & ~n21059;
  assign n21061 = ~n19897 & n21060;
  assign n21062 = ~pi165 & ~n16218;
  assign n21063 = pi774 & ~n21062;
  assign n21064 = ~pi687 & ~n21058;
  assign n21065 = ~n21063 & n21064;
  assign n21066 = ~n21061 & n21065;
  assign n21067 = ~n21057 & ~n21066;
  assign n21068 = n9830 & ~n21067;
  assign n21069 = ~pi832 & ~n21039;
  assign n21070 = ~n21068 & n21069;
  assign po322 = ~n21038 & ~n21070;
  assign n21072 = ~pi166 & ~n9830;
  assign n21073 = ~pi166 & ~n16216;
  assign n21074 = pi772 & pi947;
  assign n21075 = n16228 & ~n21074;
  assign n21076 = pi38 & ~n21075;
  assign n21077 = ~n21073 & n21076;
  assign n21078 = pi166 & ~n16057;
  assign n21079 = ~pi39 & ~n21074;
  assign n21080 = ~n16058 & ~n21079;
  assign n21081 = ~n21078 & ~n21080;
  assign n21082 = ~pi166 & n16124;
  assign n21083 = n20315 & ~n21082;
  assign n21084 = pi166 & ~n16063;
  assign n21085 = ~n19911 & ~n21084;
  assign n21086 = n2608 & ~n21085;
  assign n21087 = ~pi166 & n16186;
  assign n21088 = n20307 & ~n21087;
  assign n21089 = ~n21086 & ~n21088;
  assign n21090 = ~pi223 & ~n21089;
  assign n21091 = ~pi299 & ~n21083;
  assign n21092 = ~n21090 & n21091;
  assign n21093 = pi166 & n19885;
  assign n21094 = pi166 & n19930;
  assign n21095 = n19946 & ~n21094;
  assign n21096 = ~n16192 & n21095;
  assign n21097 = n3302 & n21085;
  assign n21098 = n19881 & ~n21097;
  assign n21099 = ~n21096 & n21098;
  assign n21100 = n19908 & ~n21093;
  assign n21101 = ~n21099 & n21100;
  assign n21102 = pi772 & ~n21092;
  assign n21103 = ~n21101 & n21102;
  assign n21104 = ~pi772 & ~n16212;
  assign n21105 = pi166 & n21104;
  assign n21106 = pi39 & ~n21103;
  assign n21107 = ~n21105 & n21106;
  assign n21108 = ~pi38 & ~n21081;
  assign n21109 = ~n21107 & n21108;
  assign n21110 = ~pi727 & ~n21077;
  assign n21111 = ~n21109 & n21110;
  assign n21112 = ~pi166 & ~n16228;
  assign n21113 = ~n19798 & n21075;
  assign n21114 = pi38 & ~n21112;
  assign n21115 = ~n21113 & n21114;
  assign n21116 = ~n19958 & n21081;
  assign n21117 = ~pi166 & ~n16203;
  assign n21118 = n19884 & ~n21117;
  assign n21119 = ~n20273 & n21118;
  assign n21120 = ~n20240 & ~n21084;
  assign n21121 = n3302 & n21120;
  assign n21122 = ~pi215 & ~n21121;
  assign n21123 = ~n19929 & n21122;
  assign n21124 = ~n21095 & n21123;
  assign n21125 = pi299 & ~n21119;
  assign n21126 = ~n21124 & n21125;
  assign n21127 = ~n6220 & ~n16124;
  assign n21128 = ~pi166 & ~n21127;
  assign n21129 = n20294 & ~n21128;
  assign n21130 = ~pi299 & ~n21129;
  assign n21131 = n2608 & n21120;
  assign n21132 = ~pi223 & ~n21131;
  assign n21133 = ~n20288 & ~n21087;
  assign n21134 = ~n2608 & ~n21133;
  assign n21135 = n2608 & n19911;
  assign n21136 = n21132 & ~n21135;
  assign n21137 = ~n21134 & n21136;
  assign n21138 = n21130 & ~n21137;
  assign n21139 = ~pi772 & ~n21138;
  assign n21140 = ~n21126 & n21139;
  assign n21141 = ~n21096 & n21122;
  assign n21142 = pi299 & ~n21118;
  assign n21143 = ~n21141 & n21142;
  assign n21144 = ~n20310 & ~n21133;
  assign n21145 = n21132 & ~n21144;
  assign n21146 = ~n21083 & n21130;
  assign n21147 = ~n21145 & n21146;
  assign n21148 = pi772 & ~n21147;
  assign n21149 = ~n21143 & n21148;
  assign n21150 = pi39 & ~n21140;
  assign n21151 = ~n21149 & n21150;
  assign n21152 = ~pi38 & ~n21116;
  assign n21153 = ~n21151 & n21152;
  assign n21154 = pi727 & ~n21115;
  assign n21155 = ~n21153 & n21154;
  assign n21156 = ~n21111 & ~n21155;
  assign n21157 = n9830 & ~n21156;
  assign n21158 = ~pi832 & ~n21072;
  assign n21159 = ~n21157 & n21158;
  assign n21160 = ~pi166 & ~n2923;
  assign n21161 = pi727 & n19798;
  assign n21162 = n2923 & ~n21074;
  assign n21163 = ~n21161 & n21162;
  assign n21164 = pi832 & ~n21160;
  assign n21165 = ~n21163 & n21164;
  assign po323 = n21159 | n21165;
  assign n21167 = ~pi167 & ~n2923;
  assign n21168 = ~pi768 & pi947;
  assign n21169 = pi705 & n19798;
  assign n21170 = ~n21168 & ~n21169;
  assign n21171 = n2923 & ~n21170;
  assign n21172 = pi832 & ~n21167;
  assign n21173 = ~n21171 & n21172;
  assign n21174 = ~pi167 & ~n9830;
  assign n21175 = ~pi167 & ~n16216;
  assign n21176 = ~n19902 & ~n21175;
  assign n21177 = pi167 & n19918;
  assign n21178 = ~pi167 & ~n19893;
  assign n21179 = ~pi38 & ~n21177;
  assign n21180 = ~n21178 & n21179;
  assign n21181 = ~pi768 & ~n21176;
  assign n21182 = ~n21180 & n21181;
  assign n21183 = ~pi167 & pi768;
  assign n21184 = ~n16218 & n21183;
  assign n21185 = ~pi705 & ~n21184;
  assign n21186 = ~n21182 & n21185;
  assign n21187 = ~pi167 & ~n19966;
  assign n21188 = n19969 & ~n21187;
  assign n21189 = ~pi167 & n19981;
  assign n21190 = pi167 & n19991;
  assign n21191 = ~pi38 & ~n21190;
  assign n21192 = ~n21189 & n21191;
  assign n21193 = ~pi768 & ~n21188;
  assign n21194 = ~n21192 & n21193;
  assign n21195 = ~pi167 & ~n16228;
  assign n21196 = n19927 & ~n21195;
  assign n21197 = ~pi167 & n19943;
  assign n21198 = pi167 & n19960;
  assign n21199 = ~pi38 & ~n21198;
  assign n21200 = ~n21197 & n21199;
  assign n21201 = pi768 & ~n21196;
  assign n21202 = ~n21200 & n21201;
  assign n21203 = pi705 & ~n21194;
  assign n21204 = ~n21202 & n21203;
  assign n21205 = n9830 & ~n21186;
  assign n21206 = ~n21204 & n21205;
  assign n21207 = ~pi832 & ~n21174;
  assign n21208 = ~n21206 & n21207;
  assign po324 = ~n21173 & ~n21208;
  assign n21210 = pi699 & n19798;
  assign n21211 = pi763 & pi947;
  assign n21212 = n2923 & ~n21211;
  assign n21213 = ~n21210 & n21212;
  assign n21214 = pi168 & ~n2923;
  assign n21215 = pi832 & ~n21214;
  assign n21216 = ~n21213 & n21215;
  assign n21217 = pi57 & pi168;
  assign n21218 = ~pi168 & ~n20005;
  assign n21219 = pi168 & ~n16216;
  assign n21220 = n16228 & ~n21211;
  assign n21221 = pi38 & ~n21220;
  assign n21222 = ~n21219 & n21221;
  assign n21223 = ~pi168 & ~pi763;
  assign n21224 = ~n16212 & n21223;
  assign n21225 = ~pi168 & ~n16190;
  assign n21226 = n19905 & ~n21225;
  assign n21227 = pi168 & ~n16203;
  assign n21228 = n19884 & ~n21227;
  assign n21229 = ~n19883 & n21228;
  assign n21230 = ~pi168 & ~n16063;
  assign n21231 = n19912 & ~n21230;
  assign n21232 = pi168 & n20201;
  assign n21233 = ~n16198 & ~n21232;
  assign n21234 = ~n21231 & n21233;
  assign n21235 = n19881 & n21234;
  assign n21236 = pi299 & ~n21229;
  assign n21237 = ~n21235 & n21236;
  assign n21238 = pi763 & ~n21237;
  assign n21239 = ~n21226 & n21238;
  assign n21240 = pi39 & ~n21224;
  assign n21241 = ~n21239 & n21240;
  assign n21242 = ~pi168 & ~n16057;
  assign n21243 = ~pi763 & n17347;
  assign n21244 = ~n19904 & ~n21243;
  assign n21245 = ~n21242 & ~n21244;
  assign n21246 = ~pi38 & ~n21245;
  assign n21247 = ~n21241 & n21246;
  assign n21248 = ~n21222 & ~n21247;
  assign n21249 = ~pi699 & ~n21248;
  assign n21250 = ~n19958 & n21245;
  assign n21251 = n19955 & ~n21225;
  assign n21252 = n19983 & ~n21228;
  assign n21253 = n19949 & ~n21230;
  assign n21254 = ~n19931 & ~n21253;
  assign n21255 = n21233 & n21254;
  assign n21256 = ~pi215 & ~n21255;
  assign n21257 = ~n19907 & ~n21252;
  assign n21258 = ~n21256 & n21257;
  assign n21259 = pi299 & ~n21258;
  assign n21260 = ~n21251 & ~n21259;
  assign n21261 = ~pi763 & ~n21260;
  assign n21262 = ~n20237 & ~n21225;
  assign n21263 = ~pi299 & ~n21262;
  assign n21264 = ~n19947 & n21231;
  assign n21265 = ~pi215 & ~n21264;
  assign n21266 = n21233 & n21265;
  assign n21267 = ~n21228 & ~n21266;
  assign n21268 = pi299 & ~n21267;
  assign n21269 = pi763 & ~n21268;
  assign n21270 = ~n21263 & n21269;
  assign n21271 = ~n21261 & ~n21270;
  assign n21272 = pi39 & ~n21271;
  assign n21273 = ~n21250 & ~n21272;
  assign n21274 = ~pi38 & ~n21273;
  assign n21275 = ~pi168 & ~n16228;
  assign n21276 = ~n19798 & ~n21211;
  assign n21277 = n16228 & ~n21276;
  assign n21278 = pi38 & ~n21275;
  assign n21279 = ~n21277 & n21278;
  assign n21280 = pi699 & ~n21279;
  assign n21281 = ~n21274 & n21280;
  assign n21282 = ~n21249 & ~n21281;
  assign n21283 = n20005 & ~n21282;
  assign n21284 = ~pi57 & ~n21218;
  assign n21285 = ~n21283 & n21284;
  assign n21286 = ~pi832 & ~n21217;
  assign n21287 = ~n21285 & n21286;
  assign po325 = n21216 | n21287;
  assign n21289 = pi729 & n19798;
  assign n21290 = pi746 & pi947;
  assign n21291 = n2923 & ~n21290;
  assign n21292 = ~n21289 & n21291;
  assign n21293 = pi169 & ~n2923;
  assign n21294 = pi832 & ~n21293;
  assign n21295 = ~n21292 & n21294;
  assign n21296 = pi57 & pi169;
  assign n21297 = ~pi169 & ~n20005;
  assign n21298 = pi169 & ~n16216;
  assign n21299 = n16228 & ~n21290;
  assign n21300 = pi38 & ~n21299;
  assign n21301 = ~n21298 & n21300;
  assign n21302 = ~pi169 & ~pi746;
  assign n21303 = ~n16212 & n21302;
  assign n21304 = ~pi169 & ~n16190;
  assign n21305 = n19905 & ~n21304;
  assign n21306 = pi169 & ~n16203;
  assign n21307 = n19884 & ~n21306;
  assign n21308 = ~n19883 & n21307;
  assign n21309 = ~pi169 & ~n16063;
  assign n21310 = n19912 & ~n21309;
  assign n21311 = pi169 & n20201;
  assign n21312 = ~n16198 & ~n21311;
  assign n21313 = ~n21310 & n21312;
  assign n21314 = n19881 & n21313;
  assign n21315 = pi299 & ~n21308;
  assign n21316 = ~n21314 & n21315;
  assign n21317 = pi746 & ~n21316;
  assign n21318 = ~n21305 & n21317;
  assign n21319 = pi39 & ~n21303;
  assign n21320 = ~n21318 & n21319;
  assign n21321 = ~pi169 & ~n16057;
  assign n21322 = ~pi746 & n17347;
  assign n21323 = ~n19904 & ~n21322;
  assign n21324 = ~n21321 & ~n21323;
  assign n21325 = ~pi38 & ~n21324;
  assign n21326 = ~n21320 & n21325;
  assign n21327 = ~n21301 & ~n21326;
  assign n21328 = ~pi729 & ~n21327;
  assign n21329 = ~n19958 & n21324;
  assign n21330 = n19955 & ~n21304;
  assign n21331 = n19983 & ~n21307;
  assign n21332 = n19949 & ~n21309;
  assign n21333 = ~n19931 & ~n21332;
  assign n21334 = n21312 & n21333;
  assign n21335 = ~pi215 & ~n21334;
  assign n21336 = ~n19907 & ~n21331;
  assign n21337 = ~n21335 & n21336;
  assign n21338 = pi299 & ~n21337;
  assign n21339 = ~n21330 & ~n21338;
  assign n21340 = ~pi746 & ~n21339;
  assign n21341 = ~n20237 & ~n21304;
  assign n21342 = ~pi299 & ~n21341;
  assign n21343 = ~n19947 & n21310;
  assign n21344 = ~pi215 & ~n21343;
  assign n21345 = n21312 & n21344;
  assign n21346 = ~n21307 & ~n21345;
  assign n21347 = pi299 & ~n21346;
  assign n21348 = pi746 & ~n21347;
  assign n21349 = ~n21342 & n21348;
  assign n21350 = ~n21340 & ~n21349;
  assign n21351 = pi39 & ~n21350;
  assign n21352 = ~n21329 & ~n21351;
  assign n21353 = ~pi38 & ~n21352;
  assign n21354 = ~pi169 & ~n16228;
  assign n21355 = ~n19798 & ~n21290;
  assign n21356 = n16228 & ~n21355;
  assign n21357 = pi38 & ~n21354;
  assign n21358 = ~n21356 & n21357;
  assign n21359 = pi729 & ~n21358;
  assign n21360 = ~n21353 & n21359;
  assign n21361 = ~n21328 & ~n21360;
  assign n21362 = n20005 & ~n21361;
  assign n21363 = ~pi57 & ~n21297;
  assign n21364 = ~n21362 & n21363;
  assign n21365 = ~pi832 & ~n21296;
  assign n21366 = ~n21364 & n21365;
  assign po326 = n21295 | n21366;
  assign n21368 = pi730 & n19798;
  assign n21369 = pi748 & pi947;
  assign n21370 = n2923 & ~n21369;
  assign n21371 = ~n21368 & n21370;
  assign n21372 = pi170 & ~n2923;
  assign n21373 = pi832 & ~n21372;
  assign n21374 = ~n21371 & n21373;
  assign n21375 = pi57 & pi170;
  assign n21376 = ~pi170 & ~n20005;
  assign n21377 = ~pi170 & ~n16228;
  assign n21378 = n19927 & ~n21377;
  assign n21379 = pi170 & ~n16203;
  assign n21380 = n19884 & ~n21379;
  assign n21381 = n19983 & ~n21380;
  assign n21382 = pi170 & n20201;
  assign n21383 = ~n16198 & ~n21382;
  assign n21384 = ~pi170 & ~n16063;
  assign n21385 = n19949 & ~n21384;
  assign n21386 = ~n19931 & ~n21385;
  assign n21387 = n21383 & n21386;
  assign n21388 = ~pi215 & ~n21387;
  assign n21389 = ~n19907 & ~n21381;
  assign n21390 = ~n21388 & n21389;
  assign n21391 = pi299 & ~n21390;
  assign n21392 = ~pi170 & ~n16190;
  assign n21393 = ~pi299 & ~n21392;
  assign n21394 = ~n19954 & n21393;
  assign n21395 = ~n21391 & ~n21394;
  assign n21396 = pi39 & ~n21395;
  assign n21397 = ~pi170 & ~n16057;
  assign n21398 = n19959 & ~n21397;
  assign n21399 = ~n21396 & ~n21398;
  assign n21400 = ~pi38 & ~n21399;
  assign n21401 = ~pi748 & ~n21378;
  assign n21402 = ~n21400 & n21401;
  assign n21403 = n19969 & ~n21377;
  assign n21404 = n19979 & ~n21397;
  assign n21405 = n19912 & ~n21384;
  assign n21406 = ~n19947 & n21405;
  assign n21407 = ~pi215 & ~n21406;
  assign n21408 = n21383 & n21407;
  assign n21409 = ~n21380 & ~n21408;
  assign n21410 = pi299 & ~n21409;
  assign n21411 = ~n20237 & ~n21392;
  assign n21412 = ~pi299 & ~n21411;
  assign n21413 = pi39 & ~n21410;
  assign n21414 = ~n21412 & n21413;
  assign n21415 = ~n21404 & ~n21414;
  assign n21416 = ~pi38 & ~n21415;
  assign n21417 = pi748 & ~n21403;
  assign n21418 = ~n21416 & n21417;
  assign n21419 = pi730 & ~n21418;
  assign n21420 = ~n21402 & n21419;
  assign n21421 = ~pi170 & ~n16216;
  assign n21422 = ~n19902 & ~n21421;
  assign n21423 = n19904 & ~n21397;
  assign n21424 = ~n19883 & n21380;
  assign n21425 = n21383 & ~n21405;
  assign n21426 = n19881 & n21425;
  assign n21427 = pi299 & ~n21424;
  assign n21428 = ~n21426 & n21427;
  assign n21429 = ~n19889 & n21393;
  assign n21430 = ~n21428 & ~n21429;
  assign n21431 = pi39 & ~n21430;
  assign n21432 = ~n21423 & ~n21431;
  assign n21433 = ~pi38 & ~n21432;
  assign n21434 = pi748 & ~n21422;
  assign n21435 = ~n21433 & n21434;
  assign n21436 = ~pi170 & ~pi748;
  assign n21437 = ~n16218 & n21436;
  assign n21438 = ~pi730 & ~n21437;
  assign n21439 = ~n21435 & n21438;
  assign n21440 = n20005 & ~n21439;
  assign n21441 = ~n21420 & n21440;
  assign n21442 = ~pi57 & ~n21376;
  assign n21443 = ~n21441 & n21442;
  assign n21444 = ~pi832 & ~n21375;
  assign n21445 = ~n21443 & n21444;
  assign po327 = n21374 | n21445;
  assign n21447 = pi691 & n19798;
  assign n21448 = pi764 & pi947;
  assign n21449 = n2923 & ~n21448;
  assign n21450 = ~n21447 & n21449;
  assign n21451 = pi171 & ~n2923;
  assign n21452 = pi832 & ~n21451;
  assign n21453 = ~n21450 & n21452;
  assign n21454 = pi57 & pi171;
  assign n21455 = ~pi171 & ~n20005;
  assign n21456 = pi171 & ~n16216;
  assign n21457 = n16228 & ~n21448;
  assign n21458 = pi38 & ~n21457;
  assign n21459 = ~n21456 & n21458;
  assign n21460 = ~pi171 & ~pi764;
  assign n21461 = ~n16212 & n21460;
  assign n21462 = ~pi171 & ~n16190;
  assign n21463 = n19905 & ~n21462;
  assign n21464 = pi171 & ~n16203;
  assign n21465 = n19884 & ~n21464;
  assign n21466 = ~n19883 & n21465;
  assign n21467 = ~pi171 & ~n16063;
  assign n21468 = n19912 & ~n21467;
  assign n21469 = pi171 & n20201;
  assign n21470 = ~n16198 & ~n21469;
  assign n21471 = ~n21468 & n21470;
  assign n21472 = n19881 & n21471;
  assign n21473 = pi299 & ~n21466;
  assign n21474 = ~n21472 & n21473;
  assign n21475 = pi764 & ~n21474;
  assign n21476 = ~n21463 & n21475;
  assign n21477 = pi39 & ~n21461;
  assign n21478 = ~n21476 & n21477;
  assign n21479 = ~pi171 & ~n16057;
  assign n21480 = ~pi764 & n17347;
  assign n21481 = ~n19904 & ~n21480;
  assign n21482 = ~n21479 & ~n21481;
  assign n21483 = ~pi38 & ~n21482;
  assign n21484 = ~n21478 & n21483;
  assign n21485 = ~n21459 & ~n21484;
  assign n21486 = ~pi691 & ~n21485;
  assign n21487 = ~n19958 & n21482;
  assign n21488 = n19955 & ~n21462;
  assign n21489 = n19983 & ~n21465;
  assign n21490 = n19949 & ~n21467;
  assign n21491 = ~n19931 & ~n21490;
  assign n21492 = n21470 & n21491;
  assign n21493 = ~pi215 & ~n21492;
  assign n21494 = ~n19907 & ~n21489;
  assign n21495 = ~n21493 & n21494;
  assign n21496 = pi299 & ~n21495;
  assign n21497 = ~n21488 & ~n21496;
  assign n21498 = ~pi764 & ~n21497;
  assign n21499 = ~n20237 & ~n21462;
  assign n21500 = ~pi299 & ~n21499;
  assign n21501 = ~n19947 & n21468;
  assign n21502 = ~pi215 & ~n21501;
  assign n21503 = n21470 & n21502;
  assign n21504 = ~n21465 & ~n21503;
  assign n21505 = pi299 & ~n21504;
  assign n21506 = pi764 & ~n21505;
  assign n21507 = ~n21500 & n21506;
  assign n21508 = ~n21498 & ~n21507;
  assign n21509 = pi39 & ~n21508;
  assign n21510 = ~n21487 & ~n21509;
  assign n21511 = ~pi38 & ~n21510;
  assign n21512 = ~pi171 & ~n16228;
  assign n21513 = ~n19798 & ~n21448;
  assign n21514 = n16228 & ~n21513;
  assign n21515 = pi38 & ~n21512;
  assign n21516 = ~n21514 & n21515;
  assign n21517 = pi691 & ~n21516;
  assign n21518 = ~n21511 & n21517;
  assign n21519 = ~n21486 & ~n21518;
  assign n21520 = n20005 & ~n21519;
  assign n21521 = ~pi57 & ~n21455;
  assign n21522 = ~n21520 & n21521;
  assign n21523 = ~pi832 & ~n21454;
  assign n21524 = ~n21522 & n21523;
  assign po328 = n21453 | n21524;
  assign n21526 = pi690 & n19798;
  assign n21527 = pi739 & pi947;
  assign n21528 = n2923 & ~n21527;
  assign n21529 = ~n21526 & n21528;
  assign n21530 = pi172 & ~n2923;
  assign n21531 = pi832 & ~n21530;
  assign n21532 = ~n21529 & n21531;
  assign n21533 = pi57 & pi172;
  assign n21534 = ~pi172 & ~n20005;
  assign n21535 = n16228 & ~n21527;
  assign n21536 = pi172 & ~n16216;
  assign n21537 = pi38 & ~n21535;
  assign n21538 = ~n21536 & n21537;
  assign n21539 = ~pi172 & ~pi739;
  assign n21540 = ~n16212 & n21539;
  assign n21541 = ~pi172 & ~n16190;
  assign n21542 = n19905 & ~n21541;
  assign n21543 = pi172 & ~n16203;
  assign n21544 = n19884 & ~n21543;
  assign n21545 = ~n19883 & n21544;
  assign n21546 = ~pi172 & ~n16063;
  assign n21547 = n19912 & ~n21546;
  assign n21548 = pi172 & n20201;
  assign n21549 = ~n16198 & ~n21548;
  assign n21550 = ~n21547 & n21549;
  assign n21551 = n19881 & n21550;
  assign n21552 = pi299 & ~n21545;
  assign n21553 = ~n21551 & n21552;
  assign n21554 = pi739 & ~n21553;
  assign n21555 = ~n21542 & n21554;
  assign n21556 = pi39 & ~n21540;
  assign n21557 = ~n21555 & n21556;
  assign n21558 = ~pi172 & ~n16057;
  assign n21559 = n16057 & n21527;
  assign n21560 = ~pi39 & ~n21558;
  assign n21561 = ~n21559 & n21560;
  assign n21562 = ~pi38 & ~n21561;
  assign n21563 = ~n21557 & n21562;
  assign n21564 = ~n21538 & ~n21563;
  assign n21565 = ~pi690 & ~n21564;
  assign n21566 = ~n19958 & n21561;
  assign n21567 = n19955 & ~n21541;
  assign n21568 = n19983 & ~n21544;
  assign n21569 = n19949 & ~n21546;
  assign n21570 = ~n19931 & ~n21569;
  assign n21571 = n21549 & n21570;
  assign n21572 = ~pi215 & ~n21571;
  assign n21573 = ~n19907 & ~n21568;
  assign n21574 = ~n21572 & n21573;
  assign n21575 = pi299 & ~n21574;
  assign n21576 = ~n21567 & ~n21575;
  assign n21577 = ~pi739 & ~n21576;
  assign n21578 = ~n20237 & ~n21541;
  assign n21579 = ~pi299 & ~n21578;
  assign n21580 = ~n19947 & n21547;
  assign n21581 = ~pi215 & ~n21580;
  assign n21582 = n21549 & n21581;
  assign n21583 = ~n21544 & ~n21582;
  assign n21584 = pi299 & ~n21583;
  assign n21585 = pi739 & ~n21584;
  assign n21586 = ~n21579 & n21585;
  assign n21587 = ~n21577 & ~n21586;
  assign n21588 = pi39 & ~n21587;
  assign n21589 = ~n21566 & ~n21588;
  assign n21590 = ~pi38 & ~n21589;
  assign n21591 = ~pi172 & ~n16228;
  assign n21592 = ~n19798 & ~n21527;
  assign n21593 = n16228 & ~n21592;
  assign n21594 = pi38 & ~n21591;
  assign n21595 = ~n21593 & n21594;
  assign n21596 = pi690 & ~n21595;
  assign n21597 = ~n21590 & n21596;
  assign n21598 = ~n21565 & ~n21597;
  assign n21599 = n20005 & ~n21598;
  assign n21600 = ~pi57 & ~n21534;
  assign n21601 = ~n21599 & n21600;
  assign n21602 = ~pi832 & ~n21533;
  assign n21603 = ~n21601 & n21602;
  assign po329 = n21532 | n21603;
  assign n21605 = ~pi173 & po1038;
  assign n21606 = ~pi173 & ~n16219;
  assign n21607 = n15747 & ~n21606;
  assign n21608 = ~pi723 & n9829;
  assign n21609 = n21606 & ~n21608;
  assign n21610 = ~pi173 & ~n16228;
  assign n21611 = n16227 & ~n21610;
  assign n21612 = ~pi173 & ~n17276;
  assign n21613 = ~pi38 & ~pi173;
  assign n21614 = n19350 & ~n21613;
  assign n21615 = ~n21612 & ~n21614;
  assign n21616 = ~pi723 & ~n21611;
  assign n21617 = ~n21615 & n21616;
  assign n21618 = ~n21609 & ~n21617;
  assign n21619 = ~pi778 & n21618;
  assign n21620 = ~pi625 & n21606;
  assign n21621 = pi625 & ~n21618;
  assign n21622 = pi1153 & ~n21620;
  assign n21623 = ~n21621 & n21622;
  assign n21624 = pi625 & n21606;
  assign n21625 = ~pi625 & ~n21618;
  assign n21626 = ~pi1153 & ~n21624;
  assign n21627 = ~n21625 & n21626;
  assign n21628 = ~n21623 & ~n21627;
  assign n21629 = pi778 & ~n21628;
  assign n21630 = ~n21619 & ~n21629;
  assign n21631 = ~n15741 & n21630;
  assign n21632 = n15741 & n21606;
  assign n21633 = ~n21631 & ~n21632;
  assign n21634 = ~n15747 & n21633;
  assign n21635 = ~n21607 & ~n21634;
  assign n21636 = ~n15753 & n21635;
  assign n21637 = n15753 & n21606;
  assign n21638 = ~n21636 & ~n21637;
  assign n21639 = ~n15759 & ~n21638;
  assign n21640 = n15759 & n21606;
  assign n21641 = ~n21639 & ~n21640;
  assign n21642 = ~pi792 & n21641;
  assign n21643 = ~pi628 & n21606;
  assign n21644 = pi628 & ~n21641;
  assign n21645 = pi1156 & ~n21643;
  assign n21646 = ~n21644 & n21645;
  assign n21647 = pi628 & n21606;
  assign n21648 = ~pi628 & ~n21641;
  assign n21649 = ~pi1156 & ~n21647;
  assign n21650 = ~n21648 & n21649;
  assign n21651 = ~n21646 & ~n21650;
  assign n21652 = pi792 & ~n21651;
  assign n21653 = ~n21642 & ~n21652;
  assign n21654 = n19394 & n21653;
  assign n21655 = ~n19394 & n21606;
  assign n21656 = ~n21654 & ~n21655;
  assign n21657 = pi787 & ~n21656;
  assign n21658 = ~pi787 & n21653;
  assign n21659 = ~n21657 & ~n21658;
  assign n21660 = ~pi644 & ~n21659;
  assign n21661 = pi715 & ~n21660;
  assign n21662 = pi173 & ~n9829;
  assign n21663 = ~pi745 & n16570;
  assign n21664 = ~n21610 & ~n21663;
  assign n21665 = pi38 & ~n21664;
  assign n21666 = ~n18599 & ~n21613;
  assign n21667 = ~pi173 & ~n16214;
  assign n21668 = pi745 & ~n21667;
  assign n21669 = ~pi173 & ~pi745;
  assign n21670 = n16514 & n21669;
  assign n21671 = ~n21666 & ~n21670;
  assign n21672 = ~n21668 & n21671;
  assign n21673 = n9829 & ~n21665;
  assign n21674 = ~n21672 & n21673;
  assign n21675 = ~n21662 & ~n21674;
  assign n21676 = ~n15777 & ~n21675;
  assign n21677 = n15777 & ~n21606;
  assign n21678 = ~n21676 & ~n21677;
  assign n21679 = ~pi785 & ~n21678;
  assign n21680 = ~n15786 & ~n21606;
  assign n21681 = pi609 & n21676;
  assign n21682 = ~n21680 & ~n21681;
  assign n21683 = pi1155 & ~n21682;
  assign n21684 = ~n16585 & ~n21606;
  assign n21685 = ~pi609 & n21676;
  assign n21686 = ~n21684 & ~n21685;
  assign n21687 = ~pi1155 & ~n21686;
  assign n21688 = ~n21683 & ~n21687;
  assign n21689 = pi785 & ~n21688;
  assign n21690 = ~n21679 & ~n21689;
  assign n21691 = ~pi781 & ~n21690;
  assign n21692 = ~pi618 & n21606;
  assign n21693 = pi618 & n21690;
  assign n21694 = pi1154 & ~n21692;
  assign n21695 = ~n21693 & n21694;
  assign n21696 = ~pi618 & n21690;
  assign n21697 = pi618 & n21606;
  assign n21698 = ~pi1154 & ~n21697;
  assign n21699 = ~n21696 & n21698;
  assign n21700 = ~n21695 & ~n21699;
  assign n21701 = pi781 & ~n21700;
  assign n21702 = ~n21691 & ~n21701;
  assign n21703 = ~pi789 & ~n21702;
  assign n21704 = ~pi619 & n21606;
  assign n21705 = pi619 & n21702;
  assign n21706 = pi1159 & ~n21704;
  assign n21707 = ~n21705 & n21706;
  assign n21708 = ~pi619 & n21702;
  assign n21709 = pi619 & n21606;
  assign n21710 = ~pi1159 & ~n21709;
  assign n21711 = ~n21708 & n21710;
  assign n21712 = ~n21707 & ~n21711;
  assign n21713 = pi789 & ~n21712;
  assign n21714 = ~n21703 & ~n21713;
  assign n21715 = n15820 & n21714;
  assign n21716 = ~n15820 & n21606;
  assign n21717 = ~n21715 & ~n21716;
  assign n21718 = pi788 & ~n21717;
  assign n21719 = ~pi788 & n21714;
  assign n21720 = ~n21718 & ~n21719;
  assign n21721 = ~n15925 & ~n21720;
  assign n21722 = n15925 & n21606;
  assign n21723 = ~n21721 & ~n21722;
  assign n21724 = ~n15960 & ~n21723;
  assign n21725 = n15960 & n21606;
  assign n21726 = ~n21724 & ~n21725;
  assign n21727 = pi644 & ~n21726;
  assign n21728 = ~pi644 & n21606;
  assign n21729 = ~pi715 & ~n21728;
  assign n21730 = ~n21727 & n21729;
  assign n21731 = pi1160 & ~n21730;
  assign n21732 = ~n21661 & n21731;
  assign n21733 = pi644 & ~n21659;
  assign n21734 = n19478 & n21723;
  assign n21735 = ~n15959 & n21656;
  assign n21736 = ~n21734 & ~n21735;
  assign n21737 = pi787 & ~n21736;
  assign n21738 = ~n16633 & n21720;
  assign n21739 = ~pi629 & n21646;
  assign n21740 = pi629 & n21650;
  assign n21741 = ~n21739 & ~n21740;
  assign n21742 = ~n21738 & n21741;
  assign n21743 = pi792 & ~n21742;
  assign n21744 = n15828 & ~n21638;
  assign n21745 = ~n15758 & ~n21717;
  assign n21746 = ~n21744 & ~n21745;
  assign n21747 = pi788 & ~n21746;
  assign n21748 = pi618 & ~n21633;
  assign n21749 = pi609 & n21630;
  assign n21750 = ~n21608 & ~n21674;
  assign n21751 = ~pi745 & ~n16808;
  assign n21752 = n18669 & ~n21751;
  assign n21753 = ~pi173 & ~n21752;
  assign n21754 = ~pi745 & n15781;
  assign n21755 = ~n16921 & ~n21754;
  assign n21756 = pi173 & ~n21755;
  assign n21757 = n6081 & n21756;
  assign n21758 = pi38 & ~n21757;
  assign n21759 = ~n21753 & n21758;
  assign n21760 = ~pi173 & ~n16647;
  assign n21761 = pi173 & ~n17397;
  assign n21762 = ~pi745 & ~n21760;
  assign n21763 = ~n21761 & n21762;
  assign n21764 = ~pi173 & n16653;
  assign n21765 = pi173 & n16657;
  assign n21766 = pi745 & ~n21764;
  assign n21767 = ~n21765 & n21766;
  assign n21768 = ~pi39 & ~n21763;
  assign n21769 = ~n21767 & n21768;
  assign n21770 = pi173 & n16825;
  assign n21771 = ~pi173 & ~n16747;
  assign n21772 = pi745 & ~n21770;
  assign n21773 = ~n21771 & n21772;
  assign n21774 = ~pi173 & n16877;
  assign n21775 = pi173 & n16913;
  assign n21776 = ~pi745 & ~n21774;
  assign n21777 = ~n21775 & n21776;
  assign n21778 = pi39 & ~n21777;
  assign n21779 = ~n21773 & n21778;
  assign n21780 = ~pi38 & ~n21769;
  assign n21781 = ~n21779 & n21780;
  assign n21782 = ~pi723 & ~n21759;
  assign n21783 = ~n21781 & n21782;
  assign n21784 = ~n21750 & ~n21783;
  assign n21785 = ~n21662 & ~n21784;
  assign n21786 = ~pi625 & n21785;
  assign n21787 = pi625 & n21675;
  assign n21788 = ~pi1153 & ~n21787;
  assign n21789 = ~n21786 & n21788;
  assign n21790 = ~pi608 & ~n21623;
  assign n21791 = ~n21789 & n21790;
  assign n21792 = ~pi625 & n21675;
  assign n21793 = pi625 & n21785;
  assign n21794 = pi1153 & ~n21792;
  assign n21795 = ~n21793 & n21794;
  assign n21796 = pi608 & ~n21627;
  assign n21797 = ~n21795 & n21796;
  assign n21798 = ~n21791 & ~n21797;
  assign n21799 = pi778 & ~n21798;
  assign n21800 = ~pi778 & n21785;
  assign n21801 = ~n21799 & ~n21800;
  assign n21802 = ~pi609 & ~n21801;
  assign n21803 = ~pi1155 & ~n21749;
  assign n21804 = ~n21802 & n21803;
  assign n21805 = ~pi660 & ~n21683;
  assign n21806 = ~n21804 & n21805;
  assign n21807 = ~pi609 & n21630;
  assign n21808 = pi609 & ~n21801;
  assign n21809 = pi1155 & ~n21807;
  assign n21810 = ~n21808 & n21809;
  assign n21811 = pi660 & ~n21687;
  assign n21812 = ~n21810 & n21811;
  assign n21813 = ~n21806 & ~n21812;
  assign n21814 = pi785 & ~n21813;
  assign n21815 = ~pi785 & ~n21801;
  assign n21816 = ~n21814 & ~n21815;
  assign n21817 = ~pi618 & ~n21816;
  assign n21818 = ~pi1154 & ~n21748;
  assign n21819 = ~n21817 & n21818;
  assign n21820 = ~pi627 & ~n21695;
  assign n21821 = ~n21819 & n21820;
  assign n21822 = ~pi618 & ~n21633;
  assign n21823 = pi618 & ~n21816;
  assign n21824 = pi1154 & ~n21822;
  assign n21825 = ~n21823 & n21824;
  assign n21826 = pi627 & ~n21699;
  assign n21827 = ~n21825 & n21826;
  assign n21828 = ~n21821 & ~n21827;
  assign n21829 = pi781 & ~n21828;
  assign n21830 = ~pi781 & ~n21816;
  assign n21831 = ~n21829 & ~n21830;
  assign n21832 = ~pi789 & n21831;
  assign n21833 = ~pi619 & n21635;
  assign n21834 = pi619 & ~n21831;
  assign n21835 = pi1159 & ~n21833;
  assign n21836 = ~n21834 & n21835;
  assign n21837 = pi648 & ~n21711;
  assign n21838 = ~n21836 & n21837;
  assign n21839 = ~pi619 & ~n21831;
  assign n21840 = pi619 & n21635;
  assign n21841 = ~pi1159 & ~n21840;
  assign n21842 = ~n21839 & n21841;
  assign n21843 = ~pi648 & ~n21707;
  assign n21844 = ~n21842 & n21843;
  assign n21845 = pi789 & ~n21838;
  assign n21846 = ~n21844 & n21845;
  assign n21847 = n15833 & ~n21832;
  assign n21848 = ~n21846 & n21847;
  assign n21849 = ~n16644 & ~n21747;
  assign n21850 = ~n21848 & n21849;
  assign n21851 = ~n21743 & ~n21850;
  assign n21852 = n18841 & ~n21851;
  assign n21853 = ~n21737 & ~n21852;
  assign n21854 = ~pi644 & n21853;
  assign n21855 = ~pi715 & ~n21733;
  assign n21856 = ~n21854 & n21855;
  assign n21857 = pi644 & n21606;
  assign n21858 = ~pi644 & ~n21726;
  assign n21859 = pi715 & ~n21857;
  assign n21860 = ~n21858 & n21859;
  assign n21861 = ~pi1160 & ~n21860;
  assign n21862 = ~n21856 & n21861;
  assign n21863 = ~n21732 & ~n21862;
  assign n21864 = pi790 & ~n21863;
  assign n21865 = pi644 & n21731;
  assign n21866 = pi790 & ~n21865;
  assign n21867 = n21853 & ~n21866;
  assign n21868 = ~n21864 & ~n21867;
  assign n21869 = ~po1038 & ~n21868;
  assign n21870 = ~pi832 & ~n21605;
  assign n21871 = ~n21869 & n21870;
  assign n21872 = ~pi173 & ~n2923;
  assign n21873 = ~pi723 & n15726;
  assign n21874 = ~n21872 & ~n21873;
  assign n21875 = ~pi778 & ~n21874;
  assign n21876 = ~pi625 & n21873;
  assign n21877 = ~n21874 & ~n21876;
  assign n21878 = pi1153 & ~n21877;
  assign n21879 = ~pi1153 & ~n21872;
  assign n21880 = ~n21876 & n21879;
  assign n21881 = pi778 & ~n21880;
  assign n21882 = ~n21878 & n21881;
  assign n21883 = ~n21875 & ~n21882;
  assign n21884 = ~n15742 & ~n21883;
  assign n21885 = ~n15748 & n21884;
  assign n21886 = ~n15754 & n21885;
  assign n21887 = ~n15760 & n21886;
  assign n21888 = ~n15766 & n21887;
  assign n21889 = n19394 & n21888;
  assign n21890 = ~n19394 & n21872;
  assign n21891 = ~n21889 & ~n21890;
  assign n21892 = ~n15959 & n21891;
  assign n21893 = n15925 & n21872;
  assign n21894 = ~n21754 & ~n21872;
  assign n21895 = ~n15778 & ~n21894;
  assign n21896 = ~pi785 & ~n21895;
  assign n21897 = n16585 & n21754;
  assign n21898 = n21895 & ~n21897;
  assign n21899 = pi1155 & ~n21898;
  assign n21900 = ~pi1155 & ~n21872;
  assign n21901 = ~n21897 & n21900;
  assign n21902 = ~n21899 & ~n21901;
  assign n21903 = pi785 & ~n21902;
  assign n21904 = ~n21896 & ~n21903;
  assign n21905 = ~pi781 & ~n21904;
  assign n21906 = ~n15797 & n21904;
  assign n21907 = pi1154 & ~n21906;
  assign n21908 = ~n15800 & n21904;
  assign n21909 = ~pi1154 & ~n21908;
  assign n21910 = ~n21907 & ~n21909;
  assign n21911 = pi781 & ~n21910;
  assign n21912 = ~n21905 & ~n21911;
  assign n21913 = pi789 & n2923;
  assign n21914 = ~n18964 & ~n18966;
  assign n21915 = n21913 & n21914;
  assign n21916 = n21912 & ~n21915;
  assign n21917 = n15820 & n21916;
  assign n21918 = ~n15820 & n21872;
  assign n21919 = ~n21917 & ~n21918;
  assign n21920 = pi788 & ~n21919;
  assign n21921 = ~pi788 & n21916;
  assign n21922 = ~n21920 & ~n21921;
  assign n21923 = ~n15925 & ~n21922;
  assign n21924 = n19478 & ~n21893;
  assign n21925 = ~n21923 & n21924;
  assign n21926 = ~n21892 & ~n21925;
  assign n21927 = pi787 & ~n21926;
  assign n21928 = ~n15758 & ~n21919;
  assign n21929 = n15828 & n21886;
  assign n21930 = ~n21928 & ~n21929;
  assign n21931 = pi788 & ~n21930;
  assign n21932 = pi619 & n2923;
  assign n21933 = n21912 & ~n21932;
  assign n21934 = pi648 & ~n21933;
  assign n21935 = pi619 & ~pi648;
  assign n21936 = ~n21885 & n21935;
  assign n21937 = ~n21934 & ~n21936;
  assign n21938 = ~pi1159 & ~n21937;
  assign n21939 = ~pi619 & ~n21885;
  assign n21940 = pi648 & ~n21939;
  assign n21941 = ~pi619 & n2923;
  assign n21942 = ~pi648 & ~n21941;
  assign n21943 = n21912 & n21942;
  assign n21944 = pi1159 & ~n21940;
  assign n21945 = ~n21943 & n21944;
  assign n21946 = ~n21938 & ~n21945;
  assign n21947 = pi789 & ~n21946;
  assign n21948 = pi609 & ~n21883;
  assign n21949 = ~n15780 & ~n21874;
  assign n21950 = pi625 & n21949;
  assign n21951 = n21894 & ~n21949;
  assign n21952 = ~n21950 & ~n21951;
  assign n21953 = n21879 & ~n21952;
  assign n21954 = ~pi608 & ~n21878;
  assign n21955 = ~n21953 & n21954;
  assign n21956 = pi1153 & n21894;
  assign n21957 = ~n21950 & n21956;
  assign n21958 = pi608 & ~n21880;
  assign n21959 = ~n21957 & n21958;
  assign n21960 = ~n21955 & ~n21959;
  assign n21961 = pi778 & ~n21960;
  assign n21962 = ~pi778 & ~n21951;
  assign n21963 = ~n21961 & ~n21962;
  assign n21964 = ~pi609 & ~n21963;
  assign n21965 = ~pi1155 & ~n21948;
  assign n21966 = ~n21964 & n21965;
  assign n21967 = ~pi660 & ~n21899;
  assign n21968 = ~n21966 & n21967;
  assign n21969 = ~pi609 & ~n21883;
  assign n21970 = pi609 & ~n21963;
  assign n21971 = pi1155 & ~n21969;
  assign n21972 = ~n21970 & n21971;
  assign n21973 = pi660 & ~n21901;
  assign n21974 = ~n21972 & n21973;
  assign n21975 = ~n21968 & ~n21974;
  assign n21976 = pi785 & ~n21975;
  assign n21977 = ~pi785 & ~n21963;
  assign n21978 = ~n21976 & ~n21977;
  assign n21979 = ~pi781 & n21978;
  assign n21980 = pi618 & n21884;
  assign n21981 = ~pi618 & ~n21978;
  assign n21982 = ~pi1154 & ~n21980;
  assign n21983 = ~n21981 & n21982;
  assign n21984 = ~pi627 & ~n21907;
  assign n21985 = ~n21983 & n21984;
  assign n21986 = ~pi618 & n21884;
  assign n21987 = pi618 & ~n21978;
  assign n21988 = pi1154 & ~n21986;
  assign n21989 = ~n21987 & n21988;
  assign n21990 = pi627 & ~n21909;
  assign n21991 = ~n21989 & n21990;
  assign n21992 = pi781 & ~n21985;
  assign n21993 = ~n21991 & n21992;
  assign n21994 = ~n21947 & ~n21979;
  assign n21995 = ~n21993 & n21994;
  assign n21996 = n18969 & n21946;
  assign n21997 = ~n21995 & ~n21996;
  assign n21998 = n15833 & ~n21997;
  assign n21999 = ~n21931 & ~n21998;
  assign n22000 = ~n16644 & ~n21999;
  assign n22001 = n15763 & ~n21922;
  assign n22002 = n15772 & n21887;
  assign n22003 = ~pi629 & ~n22002;
  assign n22004 = ~n22001 & n22003;
  assign n22005 = n15762 & ~n21922;
  assign n22006 = n15909 & n21887;
  assign n22007 = pi629 & ~n22006;
  assign n22008 = ~n22005 & n22007;
  assign n22009 = pi792 & ~n22004;
  assign n22010 = ~n22008 & n22009;
  assign n22011 = n18841 & ~n22010;
  assign n22012 = ~n22000 & n22011;
  assign n22013 = ~n21927 & ~n22012;
  assign n22014 = ~pi790 & n22013;
  assign n22015 = pi787 & ~n21891;
  assign n22016 = ~pi787 & n21888;
  assign n22017 = ~n22015 & ~n22016;
  assign n22018 = ~pi644 & ~n22017;
  assign n22019 = pi644 & n22013;
  assign n22020 = pi715 & ~n22018;
  assign n22021 = ~n22019 & n22020;
  assign n22022 = ~n19771 & n21872;
  assign n22023 = ~n15960 & n21923;
  assign n22024 = ~n22022 & ~n22023;
  assign n22025 = pi644 & ~n22024;
  assign n22026 = ~pi644 & n21872;
  assign n22027 = ~pi715 & ~n22026;
  assign n22028 = ~n22025 & n22027;
  assign n22029 = pi1160 & ~n22028;
  assign n22030 = ~n22021 & n22029;
  assign n22031 = ~pi644 & ~n22024;
  assign n22032 = pi644 & n21872;
  assign n22033 = pi715 & ~n22032;
  assign n22034 = ~n22031 & n22033;
  assign n22035 = pi644 & ~n22017;
  assign n22036 = ~pi644 & n22013;
  assign n22037 = ~pi715 & ~n22035;
  assign n22038 = ~n22036 & n22037;
  assign n22039 = ~pi1160 & ~n22034;
  assign n22040 = ~n22038 & n22039;
  assign n22041 = ~n22030 & ~n22040;
  assign n22042 = pi790 & ~n22041;
  assign n22043 = pi832 & ~n22014;
  assign n22044 = ~n22042 & n22043;
  assign po330 = ~n21871 & ~n22044;
  assign n22046 = pi174 & ~n2923;
  assign n22047 = pi759 & n15781;
  assign n22048 = n18872 & n22047;
  assign n22049 = ~pi626 & n22048;
  assign n22050 = ~n22046 & ~n22049;
  assign n22051 = ~pi1158 & ~n22050;
  assign n22052 = ~n15753 & n17584;
  assign n22053 = pi696 & n15726;
  assign n22054 = ~n22046 & ~n22053;
  assign n22055 = ~pi778 & n22054;
  assign n22056 = pi625 & n22053;
  assign n22057 = ~n22054 & ~n22056;
  assign n22058 = ~pi1153 & ~n22057;
  assign n22059 = pi1153 & ~n22046;
  assign n22060 = ~n22056 & n22059;
  assign n22061 = ~n22058 & ~n22060;
  assign n22062 = pi778 & ~n22061;
  assign n22063 = ~n22055 & ~n22062;
  assign n22064 = n22052 & n22063;
  assign n22065 = ~n22046 & ~n22064;
  assign n22066 = n15818 & ~n22065;
  assign n22067 = pi641 & ~n22051;
  assign n22068 = ~n22066 & n22067;
  assign n22069 = n15819 & ~n22065;
  assign n22070 = pi626 & n22048;
  assign n22071 = ~n22046 & ~n22070;
  assign n22072 = pi1158 & ~n22071;
  assign n22073 = ~pi641 & ~n22072;
  assign n22074 = ~n22069 & n22073;
  assign n22075 = pi788 & ~n22068;
  assign n22076 = ~n22074 & n22075;
  assign n22077 = ~n18861 & n22047;
  assign n22078 = ~n18869 & n22077;
  assign n22079 = ~n15752 & ~n22078;
  assign n22080 = n17584 & n22063;
  assign n22081 = ~n18944 & ~n22080;
  assign n22082 = ~n15777 & n18864;
  assign n22083 = ~n15752 & ~n22082;
  assign n22084 = ~n22079 & ~n22083;
  assign n22085 = ~n22081 & n22084;
  assign n22086 = pi789 & ~n22046;
  assign n22087 = ~n22085 & n22086;
  assign n22088 = ~n22046 & ~n22047;
  assign n22089 = ~n15780 & n22053;
  assign n22090 = n22088 & ~n22089;
  assign n22091 = pi625 & n22089;
  assign n22092 = ~n22090 & ~n22091;
  assign n22093 = ~pi1153 & ~n22092;
  assign n22094 = ~pi608 & ~n22060;
  assign n22095 = ~n22093 & n22094;
  assign n22096 = pi1153 & n22088;
  assign n22097 = ~n22091 & n22096;
  assign n22098 = pi608 & ~n22058;
  assign n22099 = ~n22097 & n22098;
  assign n22100 = ~n22095 & ~n22099;
  assign n22101 = pi778 & ~n22100;
  assign n22102 = ~pi778 & ~n22090;
  assign n22103 = ~n22101 & ~n22102;
  assign n22104 = ~pi609 & n22103;
  assign n22105 = pi609 & ~n22063;
  assign n22106 = ~pi1155 & ~n22105;
  assign n22107 = ~n22104 & n22106;
  assign n22108 = pi1155 & ~n15787;
  assign n22109 = ~n22088 & n22108;
  assign n22110 = ~n22107 & ~n22109;
  assign n22111 = ~pi660 & ~n22110;
  assign n22112 = n16585 & n22047;
  assign n22113 = ~pi1155 & ~n22046;
  assign n22114 = ~n22112 & n22113;
  assign n22115 = ~pi609 & n22063;
  assign n22116 = pi609 & ~n22103;
  assign n22117 = pi1155 & ~n22115;
  assign n22118 = ~n22116 & n22117;
  assign n22119 = pi660 & ~n22114;
  assign n22120 = ~n22118 & n22119;
  assign n22121 = ~n22111 & ~n22120;
  assign n22122 = pi785 & ~n22121;
  assign n22123 = ~pi785 & ~n22103;
  assign n22124 = ~n22122 & ~n22123;
  assign n22125 = ~pi781 & ~n22124;
  assign n22126 = n18950 & n22077;
  assign n22127 = pi1154 & ~n22046;
  assign n22128 = ~n22126 & n22127;
  assign n22129 = ~pi618 & ~n22124;
  assign n22130 = ~n15742 & n22063;
  assign n22131 = pi618 & n22130;
  assign n22132 = ~pi1154 & ~n22131;
  assign n22133 = ~n22129 & n22132;
  assign n22134 = ~pi627 & ~n22128;
  assign n22135 = ~n22133 & n22134;
  assign n22136 = n18955 & n22077;
  assign n22137 = ~pi1154 & ~n22046;
  assign n22138 = ~n22136 & n22137;
  assign n22139 = pi618 & ~n22124;
  assign n22140 = ~pi618 & n22130;
  assign n22141 = pi1154 & ~n22140;
  assign n22142 = ~n22139 & n22141;
  assign n22143 = pi627 & ~n22138;
  assign n22144 = ~n22142 & n22143;
  assign n22145 = ~n22135 & ~n22144;
  assign n22146 = pi781 & ~n22145;
  assign n22147 = n15752 & n18944;
  assign n22148 = pi789 & ~n22147;
  assign n22149 = ~n22125 & ~n22148;
  assign n22150 = ~n22146 & n22149;
  assign n22151 = n15833 & ~n22087;
  assign n22152 = ~n22150 & n22151;
  assign n22153 = ~n16644 & ~n22076;
  assign n22154 = ~n22152 & n22153;
  assign n22155 = ~n15759 & n22064;
  assign n22156 = ~pi628 & n22155;
  assign n22157 = pi629 & ~n22156;
  assign n22158 = ~n15832 & n22048;
  assign n22159 = pi628 & ~n22158;
  assign n22160 = ~n22157 & ~n22159;
  assign n22161 = ~pi1156 & ~n22160;
  assign n22162 = pi628 & n22155;
  assign n22163 = ~pi628 & ~n22158;
  assign n22164 = pi629 & ~n22163;
  assign n22165 = pi1156 & ~n22164;
  assign n22166 = ~n22162 & n22165;
  assign n22167 = ~n22161 & ~n22166;
  assign n22168 = pi792 & ~n22046;
  assign n22169 = ~n22167 & n22168;
  assign n22170 = ~n22154 & ~n22169;
  assign n22171 = n18841 & ~n22170;
  assign n22172 = ~n15765 & n22155;
  assign n22173 = ~pi647 & n22172;
  assign n22174 = pi630 & ~n22173;
  assign n22175 = ~n15925 & n22158;
  assign n22176 = pi647 & ~n22175;
  assign n22177 = ~n22174 & ~n22176;
  assign n22178 = ~pi1157 & ~n22177;
  assign n22179 = ~pi630 & ~n22172;
  assign n22180 = pi647 & ~n22179;
  assign n22181 = pi630 & n22175;
  assign n22182 = pi1157 & ~n22181;
  assign n22183 = ~n22180 & n22182;
  assign n22184 = ~n22178 & ~n22183;
  assign n22185 = pi787 & ~n22046;
  assign n22186 = ~n22184 & n22185;
  assign n22187 = ~n22171 & ~n22186;
  assign n22188 = ~pi790 & n22187;
  assign n22189 = ~n17768 & n22172;
  assign n22190 = ~n22046 & ~n22189;
  assign n22191 = ~pi644 & ~n22190;
  assign n22192 = pi644 & n22187;
  assign n22193 = pi715 & ~n22191;
  assign n22194 = ~n22192 & n22193;
  assign n22195 = n19771 & n22158;
  assign n22196 = pi644 & n22195;
  assign n22197 = ~pi715 & ~n22046;
  assign n22198 = ~n22196 & n22197;
  assign n22199 = pi1160 & ~n22198;
  assign n22200 = ~n22194 & n22199;
  assign n22201 = ~pi644 & n22195;
  assign n22202 = pi715 & ~n22046;
  assign n22203 = ~n22201 & n22202;
  assign n22204 = ~pi644 & n22187;
  assign n22205 = pi644 & ~n22190;
  assign n22206 = ~pi715 & ~n22205;
  assign n22207 = ~n22204 & n22206;
  assign n22208 = ~pi1160 & ~n22203;
  assign n22209 = ~n22207 & n22208;
  assign n22210 = ~n22200 & ~n22209;
  assign n22211 = pi790 & ~n22210;
  assign n22212 = pi832 & ~n22188;
  assign n22213 = ~n22211 & n22212;
  assign n22214 = pi57 & pi174;
  assign n22215 = ~pi174 & ~n6258;
  assign n22216 = pi174 & ~n16219;
  assign n22217 = n15759 & ~n22216;
  assign n22218 = n15747 & ~n22216;
  assign n22219 = pi696 & n9829;
  assign n22220 = ~n22216 & ~n22219;
  assign n22221 = ~pi174 & ~n17272;
  assign n22222 = pi174 & n17276;
  assign n22223 = ~pi38 & ~n22221;
  assign n22224 = ~n22222 & n22223;
  assign n22225 = ~pi174 & ~n16228;
  assign n22226 = n19049 & ~n22225;
  assign n22227 = n22219 & ~n22226;
  assign n22228 = ~n22224 & n22227;
  assign n22229 = ~n22220 & ~n22228;
  assign n22230 = ~pi778 & n22229;
  assign n22231 = ~pi625 & ~n22216;
  assign n22232 = pi625 & ~n22229;
  assign n22233 = pi1153 & ~n22231;
  assign n22234 = ~n22232 & n22233;
  assign n22235 = ~pi625 & ~n22229;
  assign n22236 = pi625 & ~n22216;
  assign n22237 = ~pi1153 & ~n22236;
  assign n22238 = ~n22235 & n22237;
  assign n22239 = ~n22234 & ~n22238;
  assign n22240 = pi778 & ~n22239;
  assign n22241 = ~n22230 & ~n22240;
  assign n22242 = ~n15741 & ~n22241;
  assign n22243 = n15741 & n22216;
  assign n22244 = ~n22242 & ~n22243;
  assign n22245 = ~n15747 & n22244;
  assign n22246 = ~n22218 & ~n22245;
  assign n22247 = ~n15753 & n22246;
  assign n22248 = n15753 & n22216;
  assign n22249 = ~n22247 & ~n22248;
  assign n22250 = ~n15759 & n22249;
  assign n22251 = ~n22217 & ~n22250;
  assign n22252 = ~pi792 & n22251;
  assign n22253 = pi628 & n22251;
  assign n22254 = ~pi628 & n22216;
  assign n22255 = ~n22253 & ~n22254;
  assign n22256 = pi1156 & ~n22255;
  assign n22257 = pi628 & ~n22216;
  assign n22258 = ~pi628 & ~n22251;
  assign n22259 = ~pi1156 & ~n22257;
  assign n22260 = ~n22258 & n22259;
  assign n22261 = ~n22256 & ~n22260;
  assign n22262 = pi792 & ~n22261;
  assign n22263 = ~n22252 & ~n22262;
  assign n22264 = ~pi787 & ~n22263;
  assign n22265 = ~pi647 & ~n22216;
  assign n22266 = pi647 & n22263;
  assign n22267 = pi1157 & ~n22265;
  assign n22268 = ~n22266 & n22267;
  assign n22269 = pi647 & ~n22216;
  assign n22270 = ~pi647 & n22263;
  assign n22271 = ~pi1157 & ~n22269;
  assign n22272 = ~n22270 & n22271;
  assign n22273 = ~n22268 & ~n22272;
  assign n22274 = pi787 & ~n22273;
  assign n22275 = ~n22264 & ~n22274;
  assign n22276 = ~pi644 & n22275;
  assign n22277 = ~pi629 & n22256;
  assign n22278 = pi174 & ~n9829;
  assign n22279 = pi759 & ~n16512;
  assign n22280 = ~n20344 & ~n22279;
  assign n22281 = pi39 & ~n22280;
  assign n22282 = ~pi759 & n16057;
  assign n22283 = n16448 & ~n22282;
  assign n22284 = ~n22281 & ~n22283;
  assign n22285 = pi174 & ~n22284;
  assign n22286 = ~pi174 & pi759;
  assign n22287 = n16565 & n22286;
  assign n22288 = ~n22285 & ~n22287;
  assign n22289 = ~pi38 & ~n22288;
  assign n22290 = pi759 & n15780;
  assign n22291 = n16228 & ~n22290;
  assign n22292 = pi38 & ~n22225;
  assign n22293 = ~n22291 & n22292;
  assign n22294 = ~n22289 & ~n22293;
  assign n22295 = n9829 & ~n22294;
  assign n22296 = ~n22278 & ~n22295;
  assign n22297 = ~n15777 & ~n22296;
  assign n22298 = n15777 & n22216;
  assign n22299 = ~n22297 & ~n22298;
  assign n22300 = ~pi785 & ~n22299;
  assign n22301 = pi609 & n22299;
  assign n22302 = ~pi609 & ~n22216;
  assign n22303 = pi1155 & ~n22302;
  assign n22304 = ~n22301 & n22303;
  assign n22305 = ~pi609 & n22299;
  assign n22306 = pi609 & ~n22216;
  assign n22307 = ~pi1155 & ~n22306;
  assign n22308 = ~n22305 & n22307;
  assign n22309 = ~n22304 & ~n22308;
  assign n22310 = pi785 & ~n22309;
  assign n22311 = ~n22300 & ~n22310;
  assign n22312 = ~pi781 & ~n22311;
  assign n22313 = ~pi618 & ~n22216;
  assign n22314 = pi618 & n22311;
  assign n22315 = pi1154 & ~n22313;
  assign n22316 = ~n22314 & n22315;
  assign n22317 = pi618 & ~n22216;
  assign n22318 = ~pi618 & n22311;
  assign n22319 = ~pi1154 & ~n22317;
  assign n22320 = ~n22318 & n22319;
  assign n22321 = ~n22316 & ~n22320;
  assign n22322 = pi781 & ~n22321;
  assign n22323 = ~n22312 & ~n22322;
  assign n22324 = ~pi789 & ~n22323;
  assign n22325 = ~pi619 & ~n22216;
  assign n22326 = pi619 & n22323;
  assign n22327 = pi1159 & ~n22325;
  assign n22328 = ~n22326 & n22327;
  assign n22329 = pi619 & ~n22216;
  assign n22330 = ~pi619 & n22323;
  assign n22331 = ~pi1159 & ~n22329;
  assign n22332 = ~n22330 & n22331;
  assign n22333 = ~n22328 & ~n22332;
  assign n22334 = pi789 & ~n22333;
  assign n22335 = ~n22324 & ~n22334;
  assign n22336 = ~n15832 & ~n22335;
  assign n22337 = n15832 & n22216;
  assign n22338 = ~n22336 & ~n22337;
  assign n22339 = ~n16633 & ~n22338;
  assign n22340 = pi629 & n22260;
  assign n22341 = ~n22277 & ~n22340;
  assign n22342 = ~n22339 & n22341;
  assign n22343 = pi792 & ~n22342;
  assign n22344 = pi641 & n22216;
  assign n22345 = ~pi641 & ~n22249;
  assign n22346 = n15819 & ~n22344;
  assign n22347 = ~n22345 & n22346;
  assign n22348 = ~n15758 & ~n15827;
  assign n22349 = n22335 & n22348;
  assign n22350 = ~pi641 & n22216;
  assign n22351 = pi641 & ~n22249;
  assign n22352 = n15818 & ~n22350;
  assign n22353 = ~n22351 & n22352;
  assign n22354 = ~n22347 & ~n22353;
  assign n22355 = ~n22349 & n22354;
  assign n22356 = pi788 & ~n22355;
  assign n22357 = pi609 & n22241;
  assign n22358 = ~n22219 & ~n22295;
  assign n22359 = ~pi174 & ~n16657;
  assign n22360 = pi174 & ~n16653;
  assign n22361 = ~pi759 & ~n22359;
  assign n22362 = ~n22360 & n22361;
  assign n22363 = ~pi174 & n17397;
  assign n22364 = pi174 & n16647;
  assign n22365 = pi759 & ~n22363;
  assign n22366 = ~n22364 & n22365;
  assign n22367 = ~pi39 & ~n22366;
  assign n22368 = ~n22362 & n22367;
  assign n22369 = pi174 & ~n16877;
  assign n22370 = ~pi174 & ~n16913;
  assign n22371 = pi759 & ~n22369;
  assign n22372 = ~n22370 & n22371;
  assign n22373 = pi174 & n16747;
  assign n22374 = ~pi174 & ~n16825;
  assign n22375 = ~pi759 & ~n22374;
  assign n22376 = ~n22373 & n22375;
  assign n22377 = pi39 & ~n22372;
  assign n22378 = ~n22376 & n22377;
  assign n22379 = ~pi38 & ~n22368;
  assign n22380 = ~n22378 & n22379;
  assign n22381 = pi696 & ~n18668;
  assign n22382 = ~n22293 & n22381;
  assign n22383 = ~n22380 & n22382;
  assign n22384 = ~n22358 & ~n22383;
  assign n22385 = ~n22278 & ~n22384;
  assign n22386 = ~pi625 & n22385;
  assign n22387 = pi625 & n22296;
  assign n22388 = ~pi1153 & ~n22387;
  assign n22389 = ~n22386 & n22388;
  assign n22390 = ~pi608 & ~n22234;
  assign n22391 = ~n22389 & n22390;
  assign n22392 = ~pi625 & n22296;
  assign n22393 = pi625 & n22385;
  assign n22394 = pi1153 & ~n22392;
  assign n22395 = ~n22393 & n22394;
  assign n22396 = pi608 & ~n22238;
  assign n22397 = ~n22395 & n22396;
  assign n22398 = ~n22391 & ~n22397;
  assign n22399 = pi778 & ~n22398;
  assign n22400 = ~pi778 & n22385;
  assign n22401 = ~n22399 & ~n22400;
  assign n22402 = ~pi609 & ~n22401;
  assign n22403 = ~pi1155 & ~n22357;
  assign n22404 = ~n22402 & n22403;
  assign n22405 = ~pi660 & ~n22304;
  assign n22406 = ~n22404 & n22405;
  assign n22407 = ~pi609 & n22241;
  assign n22408 = pi609 & ~n22401;
  assign n22409 = pi1155 & ~n22407;
  assign n22410 = ~n22408 & n22409;
  assign n22411 = pi660 & ~n22308;
  assign n22412 = ~n22410 & n22411;
  assign n22413 = ~n22406 & ~n22412;
  assign n22414 = pi785 & ~n22413;
  assign n22415 = ~pi785 & ~n22401;
  assign n22416 = ~n22414 & ~n22415;
  assign n22417 = ~pi618 & ~n22416;
  assign n22418 = pi618 & n22244;
  assign n22419 = ~pi1154 & ~n22418;
  assign n22420 = ~n22417 & n22419;
  assign n22421 = ~pi627 & ~n22316;
  assign n22422 = ~n22420 & n22421;
  assign n22423 = ~pi618 & n22244;
  assign n22424 = pi618 & ~n22416;
  assign n22425 = pi1154 & ~n22423;
  assign n22426 = ~n22424 & n22425;
  assign n22427 = pi627 & ~n22320;
  assign n22428 = ~n22426 & n22427;
  assign n22429 = ~n22422 & ~n22428;
  assign n22430 = pi781 & ~n22429;
  assign n22431 = ~pi781 & ~n22416;
  assign n22432 = ~n22430 & ~n22431;
  assign n22433 = ~pi789 & n22432;
  assign n22434 = ~pi619 & ~n22246;
  assign n22435 = pi619 & ~n22432;
  assign n22436 = pi1159 & ~n22434;
  assign n22437 = ~n22435 & n22436;
  assign n22438 = pi648 & ~n22332;
  assign n22439 = ~n22437 & n22438;
  assign n22440 = pi619 & ~n22246;
  assign n22441 = ~pi619 & ~n22432;
  assign n22442 = ~pi1159 & ~n22440;
  assign n22443 = ~n22441 & n22442;
  assign n22444 = ~pi648 & ~n22328;
  assign n22445 = ~n22443 & n22444;
  assign n22446 = pi789 & ~n22439;
  assign n22447 = ~n22445 & n22446;
  assign n22448 = n15833 & ~n22433;
  assign n22449 = ~n22447 & n22448;
  assign n22450 = ~n16644 & ~n22356;
  assign n22451 = ~n22449 & n22450;
  assign n22452 = ~n22343 & ~n22451;
  assign n22453 = ~pi647 & n22452;
  assign n22454 = ~n15925 & ~n22338;
  assign n22455 = n15925 & n22216;
  assign n22456 = ~n22454 & ~n22455;
  assign n22457 = pi647 & n22456;
  assign n22458 = ~pi1157 & ~n22457;
  assign n22459 = ~n22453 & n22458;
  assign n22460 = ~pi630 & ~n22268;
  assign n22461 = ~n22459 & n22460;
  assign n22462 = ~pi647 & n22456;
  assign n22463 = pi647 & n22452;
  assign n22464 = pi1157 & ~n22462;
  assign n22465 = ~n22463 & n22464;
  assign n22466 = pi630 & ~n22272;
  assign n22467 = ~n22465 & n22466;
  assign n22468 = ~n22461 & ~n22467;
  assign n22469 = pi787 & ~n22468;
  assign n22470 = ~pi787 & n22452;
  assign n22471 = ~n22469 & ~n22470;
  assign n22472 = pi644 & ~n22471;
  assign n22473 = pi715 & ~n22276;
  assign n22474 = ~n22472 & n22473;
  assign n22475 = ~n15960 & ~n22456;
  assign n22476 = n15960 & n22216;
  assign n22477 = ~n22475 & ~n22476;
  assign n22478 = pi644 & n22477;
  assign n22479 = ~pi644 & ~n22216;
  assign n22480 = ~pi715 & ~n22479;
  assign n22481 = ~n22478 & n22480;
  assign n22482 = pi1160 & ~n22481;
  assign n22483 = ~n22474 & n22482;
  assign n22484 = pi644 & n22275;
  assign n22485 = ~pi715 & ~n22484;
  assign n22486 = ~pi644 & n22477;
  assign n22487 = pi644 & ~n22216;
  assign n22488 = pi715 & ~n22487;
  assign n22489 = ~n22486 & n22488;
  assign n22490 = ~pi1160 & ~n22489;
  assign n22491 = ~n22485 & n22490;
  assign n22492 = ~n22483 & ~n22491;
  assign n22493 = pi790 & ~n22492;
  assign n22494 = ~pi644 & n22490;
  assign n22495 = pi790 & ~n22494;
  assign n22496 = ~n22471 & ~n22495;
  assign n22497 = ~n22493 & ~n22496;
  assign n22498 = n6258 & ~n22497;
  assign n22499 = ~pi57 & ~n22215;
  assign n22500 = ~n22498 & n22499;
  assign n22501 = ~pi832 & ~n22214;
  assign n22502 = ~n22500 & n22501;
  assign po331 = ~n22213 & ~n22502;
  assign n22504 = ~pi175 & ~n2923;
  assign n22505 = pi700 & n15726;
  assign n22506 = ~n22504 & ~n22505;
  assign n22507 = ~pi778 & ~n22506;
  assign n22508 = ~pi625 & n22505;
  assign n22509 = ~n22506 & ~n22508;
  assign n22510 = pi1153 & ~n22509;
  assign n22511 = ~pi1153 & ~n22504;
  assign n22512 = ~n22508 & n22511;
  assign n22513 = pi778 & ~n22512;
  assign n22514 = ~n22510 & n22513;
  assign n22515 = ~n22507 & ~n22514;
  assign n22516 = ~n15742 & ~n22515;
  assign n22517 = ~n15748 & n22516;
  assign n22518 = ~n15754 & n22517;
  assign n22519 = ~n15760 & n22518;
  assign n22520 = ~n15766 & n22519;
  assign n22521 = n19394 & n22520;
  assign n22522 = ~n19394 & n22504;
  assign n22523 = ~n22521 & ~n22522;
  assign n22524 = ~n15959 & n22523;
  assign n22525 = n15925 & n22504;
  assign n22526 = pi766 & n15781;
  assign n22527 = ~n22504 & ~n22526;
  assign n22528 = ~n15778 & ~n22527;
  assign n22529 = ~pi785 & ~n22528;
  assign n22530 = n16585 & n22526;
  assign n22531 = n22528 & ~n22530;
  assign n22532 = pi1155 & ~n22531;
  assign n22533 = ~pi1155 & ~n22504;
  assign n22534 = ~n22530 & n22533;
  assign n22535 = ~n22532 & ~n22534;
  assign n22536 = pi785 & ~n22535;
  assign n22537 = ~n22529 & ~n22536;
  assign n22538 = ~pi781 & ~n22537;
  assign n22539 = ~n15797 & n22537;
  assign n22540 = pi1154 & ~n22539;
  assign n22541 = ~n15800 & n22537;
  assign n22542 = ~pi1154 & ~n22541;
  assign n22543 = ~n22540 & ~n22542;
  assign n22544 = pi781 & ~n22543;
  assign n22545 = ~n22538 & ~n22544;
  assign n22546 = ~n21915 & n22545;
  assign n22547 = ~n15832 & ~n22546;
  assign n22548 = n15832 & ~n22504;
  assign n22549 = ~n22547 & ~n22548;
  assign n22550 = ~n15925 & n22549;
  assign n22551 = n19478 & ~n22525;
  assign n22552 = ~n22550 & n22551;
  assign n22553 = ~n22524 & ~n22552;
  assign n22554 = pi787 & ~n22553;
  assign n22555 = n15763 & n22549;
  assign n22556 = n15772 & n22519;
  assign n22557 = ~pi629 & ~n22556;
  assign n22558 = ~n22555 & n22557;
  assign n22559 = n15762 & n22549;
  assign n22560 = n15909 & n22519;
  assign n22561 = pi629 & ~n22560;
  assign n22562 = ~n22559 & n22561;
  assign n22563 = pi792 & ~n22558;
  assign n22564 = ~n22562 & n22563;
  assign n22565 = ~n21932 & n22545;
  assign n22566 = pi648 & ~n22565;
  assign n22567 = n21935 & ~n22517;
  assign n22568 = ~n22566 & ~n22567;
  assign n22569 = ~pi1159 & ~n22568;
  assign n22570 = ~pi619 & ~n22517;
  assign n22571 = pi648 & ~n22570;
  assign n22572 = n21942 & n22545;
  assign n22573 = pi1159 & ~n22571;
  assign n22574 = ~n22572 & n22573;
  assign n22575 = ~n22569 & ~n22574;
  assign n22576 = pi789 & ~n22575;
  assign n22577 = pi609 & ~n22515;
  assign n22578 = ~n15780 & ~n22506;
  assign n22579 = pi625 & n22578;
  assign n22580 = n22527 & ~n22578;
  assign n22581 = ~n22579 & ~n22580;
  assign n22582 = n22511 & ~n22581;
  assign n22583 = ~pi608 & ~n22510;
  assign n22584 = ~n22582 & n22583;
  assign n22585 = pi1153 & n22527;
  assign n22586 = ~n22579 & n22585;
  assign n22587 = pi608 & ~n22512;
  assign n22588 = ~n22586 & n22587;
  assign n22589 = ~n22584 & ~n22588;
  assign n22590 = pi778 & ~n22589;
  assign n22591 = ~pi778 & ~n22580;
  assign n22592 = ~n22590 & ~n22591;
  assign n22593 = ~pi609 & ~n22592;
  assign n22594 = ~pi1155 & ~n22577;
  assign n22595 = ~n22593 & n22594;
  assign n22596 = ~pi660 & ~n22532;
  assign n22597 = ~n22595 & n22596;
  assign n22598 = ~pi609 & ~n22515;
  assign n22599 = pi609 & ~n22592;
  assign n22600 = pi1155 & ~n22598;
  assign n22601 = ~n22599 & n22600;
  assign n22602 = pi660 & ~n22534;
  assign n22603 = ~n22601 & n22602;
  assign n22604 = ~n22597 & ~n22603;
  assign n22605 = pi785 & ~n22604;
  assign n22606 = ~pi785 & ~n22592;
  assign n22607 = ~n22605 & ~n22606;
  assign n22608 = ~pi781 & n22607;
  assign n22609 = pi618 & n22516;
  assign n22610 = ~pi618 & ~n22607;
  assign n22611 = ~pi1154 & ~n22609;
  assign n22612 = ~n22610 & n22611;
  assign n22613 = ~pi627 & ~n22540;
  assign n22614 = ~n22612 & n22613;
  assign n22615 = ~pi618 & n22516;
  assign n22616 = pi618 & ~n22607;
  assign n22617 = pi1154 & ~n22615;
  assign n22618 = ~n22616 & n22617;
  assign n22619 = pi627 & ~n22542;
  assign n22620 = ~n22618 & n22619;
  assign n22621 = pi781 & ~n22614;
  assign n22622 = ~n22620 & n22621;
  assign n22623 = ~n22576 & ~n22608;
  assign n22624 = ~n22622 & n22623;
  assign n22625 = n18969 & n22575;
  assign n22626 = ~n22624 & ~n22625;
  assign n22627 = n15833 & ~n22626;
  assign n22628 = n15828 & n22518;
  assign n22629 = ~pi626 & ~n22504;
  assign n22630 = pi626 & ~n22546;
  assign n22631 = n15756 & ~n22629;
  assign n22632 = ~n22630 & n22631;
  assign n22633 = pi626 & ~n22504;
  assign n22634 = ~pi626 & ~n22546;
  assign n22635 = n15757 & ~n22633;
  assign n22636 = ~n22634 & n22635;
  assign n22637 = ~n22628 & ~n22632;
  assign n22638 = ~n22636 & n22637;
  assign n22639 = pi788 & ~n22638;
  assign n22640 = ~n22627 & ~n22639;
  assign n22641 = ~n16644 & ~n22640;
  assign n22642 = n18841 & ~n22564;
  assign n22643 = ~n22641 & n22642;
  assign n22644 = ~n22554 & ~n22643;
  assign n22645 = ~pi790 & n22644;
  assign n22646 = pi787 & ~n22523;
  assign n22647 = ~pi787 & n22520;
  assign n22648 = ~n22646 & ~n22647;
  assign n22649 = ~pi644 & ~n22648;
  assign n22650 = pi644 & n22644;
  assign n22651 = pi715 & ~n22649;
  assign n22652 = ~n22650 & n22651;
  assign n22653 = ~n19771 & n22504;
  assign n22654 = ~n15960 & n22550;
  assign n22655 = ~n22653 & ~n22654;
  assign n22656 = pi644 & ~n22655;
  assign n22657 = ~pi644 & n22504;
  assign n22658 = ~pi715 & ~n22657;
  assign n22659 = ~n22656 & n22658;
  assign n22660 = pi1160 & ~n22659;
  assign n22661 = ~n22652 & n22660;
  assign n22662 = ~pi644 & ~n22655;
  assign n22663 = pi644 & n22504;
  assign n22664 = pi715 & ~n22663;
  assign n22665 = ~n22662 & n22664;
  assign n22666 = pi644 & ~n22648;
  assign n22667 = ~pi644 & n22644;
  assign n22668 = ~pi715 & ~n22666;
  assign n22669 = ~n22667 & n22668;
  assign n22670 = ~pi1160 & ~n22665;
  assign n22671 = ~n22669 & n22670;
  assign n22672 = ~n22661 & ~n22671;
  assign n22673 = pi790 & ~n22672;
  assign n22674 = pi832 & ~n22645;
  assign n22675 = ~n22673 & n22674;
  assign n22676 = ~pi175 & po1038;
  assign n22677 = ~pi175 & ~n16219;
  assign n22678 = n15747 & ~n22677;
  assign n22679 = pi175 & ~n9829;
  assign n22680 = ~pi175 & ~n16228;
  assign n22681 = n16227 & ~n22680;
  assign n22682 = pi175 & n17272;
  assign n22683 = ~pi175 & ~n17276;
  assign n22684 = ~pi38 & ~n22682;
  assign n22685 = ~n22683 & n22684;
  assign n22686 = pi700 & ~n22681;
  assign n22687 = ~n22685 & n22686;
  assign n22688 = ~pi175 & ~pi700;
  assign n22689 = ~n16218 & n22688;
  assign n22690 = n9829 & ~n22687;
  assign n22691 = ~n22689 & n22690;
  assign n22692 = ~n22679 & ~n22691;
  assign n22693 = ~pi778 & ~n22692;
  assign n22694 = ~pi625 & n22677;
  assign n22695 = pi625 & n22692;
  assign n22696 = pi1153 & ~n22694;
  assign n22697 = ~n22695 & n22696;
  assign n22698 = ~pi625 & n22692;
  assign n22699 = pi625 & n22677;
  assign n22700 = ~pi1153 & ~n22699;
  assign n22701 = ~n22698 & n22700;
  assign n22702 = ~n22697 & ~n22701;
  assign n22703 = pi778 & ~n22702;
  assign n22704 = ~n22693 & ~n22703;
  assign n22705 = ~n15741 & n22704;
  assign n22706 = n15741 & n22677;
  assign n22707 = ~n22705 & ~n22706;
  assign n22708 = ~n15747 & n22707;
  assign n22709 = ~n22678 & ~n22708;
  assign n22710 = ~n15753 & n22709;
  assign n22711 = n15753 & n22677;
  assign n22712 = ~n22710 & ~n22711;
  assign n22713 = ~n15759 & ~n22712;
  assign n22714 = n15759 & n22677;
  assign n22715 = ~n22713 & ~n22714;
  assign n22716 = ~n15765 & ~n22715;
  assign n22717 = n15765 & n22677;
  assign n22718 = ~n22716 & ~n22717;
  assign n22719 = ~n17768 & ~n22718;
  assign n22720 = n17768 & n22677;
  assign n22721 = ~n22719 & ~n22720;
  assign n22722 = ~pi644 & ~n22721;
  assign n22723 = pi715 & ~n22722;
  assign n22724 = ~pi766 & n16212;
  assign n22725 = pi175 & ~n16563;
  assign n22726 = ~n22724 & ~n22725;
  assign n22727 = pi39 & ~n22726;
  assign n22728 = pi766 & ~n16527;
  assign n22729 = pi175 & ~n22728;
  assign n22730 = ~pi175 & pi766;
  assign n22731 = n16514 & n22730;
  assign n22732 = ~n20396 & ~n22729;
  assign n22733 = ~n22731 & n22732;
  assign n22734 = ~n22727 & n22733;
  assign n22735 = ~pi38 & ~n22734;
  assign n22736 = pi766 & n16570;
  assign n22737 = pi38 & ~n22680;
  assign n22738 = ~n22736 & n22737;
  assign n22739 = ~n22735 & ~n22738;
  assign n22740 = n9829 & ~n22739;
  assign n22741 = ~n22679 & ~n22740;
  assign n22742 = ~n15777 & ~n22741;
  assign n22743 = n15777 & ~n22677;
  assign n22744 = ~n22742 & ~n22743;
  assign n22745 = ~pi785 & ~n22744;
  assign n22746 = ~n15786 & ~n22677;
  assign n22747 = pi609 & n22742;
  assign n22748 = ~n22746 & ~n22747;
  assign n22749 = pi1155 & ~n22748;
  assign n22750 = ~n16585 & ~n22677;
  assign n22751 = ~pi609 & n22742;
  assign n22752 = ~n22750 & ~n22751;
  assign n22753 = ~pi1155 & ~n22752;
  assign n22754 = ~n22749 & ~n22753;
  assign n22755 = pi785 & ~n22754;
  assign n22756 = ~n22745 & ~n22755;
  assign n22757 = ~pi781 & ~n22756;
  assign n22758 = ~pi618 & n22677;
  assign n22759 = pi618 & n22756;
  assign n22760 = pi1154 & ~n22758;
  assign n22761 = ~n22759 & n22760;
  assign n22762 = ~pi618 & n22756;
  assign n22763 = pi618 & n22677;
  assign n22764 = ~pi1154 & ~n22763;
  assign n22765 = ~n22762 & n22764;
  assign n22766 = ~n22761 & ~n22765;
  assign n22767 = pi781 & ~n22766;
  assign n22768 = ~n22757 & ~n22767;
  assign n22769 = ~pi789 & ~n22768;
  assign n22770 = ~pi619 & n22677;
  assign n22771 = pi619 & n22768;
  assign n22772 = pi1159 & ~n22770;
  assign n22773 = ~n22771 & n22772;
  assign n22774 = ~pi619 & n22768;
  assign n22775 = pi619 & n22677;
  assign n22776 = ~pi1159 & ~n22775;
  assign n22777 = ~n22774 & n22776;
  assign n22778 = ~n22773 & ~n22777;
  assign n22779 = pi789 & ~n22778;
  assign n22780 = ~n22769 & ~n22779;
  assign n22781 = ~n15832 & n22780;
  assign n22782 = n15832 & n22677;
  assign n22783 = ~n22781 & ~n22782;
  assign n22784 = ~n15925 & ~n22783;
  assign n22785 = n15925 & n22677;
  assign n22786 = ~n22784 & ~n22785;
  assign n22787 = ~n15960 & ~n22786;
  assign n22788 = n15960 & n22677;
  assign n22789 = ~n22787 & ~n22788;
  assign n22790 = pi644 & ~n22789;
  assign n22791 = ~pi644 & n22677;
  assign n22792 = ~pi715 & ~n22791;
  assign n22793 = ~n22790 & n22792;
  assign n22794 = pi1160 & ~n22723;
  assign n22795 = ~n22793 & n22794;
  assign n22796 = pi644 & ~n22721;
  assign n22797 = ~pi715 & ~n22796;
  assign n22798 = ~pi644 & ~n22789;
  assign n22799 = pi644 & n22677;
  assign n22800 = pi715 & ~n22799;
  assign n22801 = ~n22798 & n22800;
  assign n22802 = ~pi1160 & ~n22801;
  assign n22803 = ~n22797 & n22802;
  assign n22804 = ~n22795 & ~n22803;
  assign n22805 = pi790 & ~n22804;
  assign n22806 = ~pi647 & n22677;
  assign n22807 = pi647 & ~n22718;
  assign n22808 = n15957 & ~n22806;
  assign n22809 = ~n22807 & n22808;
  assign n22810 = n19478 & n22786;
  assign n22811 = pi647 & n22677;
  assign n22812 = ~pi647 & ~n22718;
  assign n22813 = n15958 & ~n22811;
  assign n22814 = ~n22812 & n22813;
  assign n22815 = ~n22809 & ~n22814;
  assign n22816 = ~n22810 & n22815;
  assign n22817 = pi787 & ~n22816;
  assign n22818 = pi628 & n22677;
  assign n22819 = ~pi628 & ~n22715;
  assign n22820 = n15923 & ~n22818;
  assign n22821 = ~n22819 & n22820;
  assign n22822 = ~n16633 & n22783;
  assign n22823 = ~pi628 & n22677;
  assign n22824 = pi628 & ~n22715;
  assign n22825 = n15922 & ~n22823;
  assign n22826 = ~n22824 & n22825;
  assign n22827 = ~n22821 & ~n22826;
  assign n22828 = ~n22822 & n22827;
  assign n22829 = pi792 & ~n22828;
  assign n22830 = n15828 & ~n22712;
  assign n22831 = ~pi626 & ~n22677;
  assign n22832 = pi626 & ~n22780;
  assign n22833 = n15756 & ~n22831;
  assign n22834 = ~n22832 & n22833;
  assign n22835 = pi626 & ~n22677;
  assign n22836 = ~pi626 & ~n22780;
  assign n22837 = n15757 & ~n22835;
  assign n22838 = ~n22836 & n22837;
  assign n22839 = ~n22830 & ~n22834;
  assign n22840 = ~n22838 & n22839;
  assign n22841 = pi788 & ~n22840;
  assign n22842 = pi618 & ~n22707;
  assign n22843 = pi609 & n22704;
  assign n22844 = ~pi700 & n22739;
  assign n22845 = ~n16921 & ~n22526;
  assign n22846 = pi175 & ~n22845;
  assign n22847 = n6081 & n22846;
  assign n22848 = n16065 & ~n16663;
  assign n22849 = ~pi766 & n22848;
  assign n22850 = ~n16808 & ~n22849;
  assign n22851 = ~pi39 & ~n22850;
  assign n22852 = ~pi175 & ~n22851;
  assign n22853 = pi38 & ~n22847;
  assign n22854 = ~n22852 & n22853;
  assign n22855 = ~pi175 & n16653;
  assign n22856 = pi175 & n16657;
  assign n22857 = ~pi766 & ~n22855;
  assign n22858 = ~n22856 & n22857;
  assign n22859 = ~pi175 & ~n16647;
  assign n22860 = pi175 & ~n17397;
  assign n22861 = pi766 & ~n22859;
  assign n22862 = ~n22860 & n22861;
  assign n22863 = ~pi39 & ~n22862;
  assign n22864 = ~n22858 & n22863;
  assign n22865 = ~pi175 & n16877;
  assign n22866 = pi175 & n16913;
  assign n22867 = pi766 & ~n22865;
  assign n22868 = ~n22866 & n22867;
  assign n22869 = pi175 & n16825;
  assign n22870 = ~pi175 & ~n16747;
  assign n22871 = ~pi766 & ~n22869;
  assign n22872 = ~n22870 & n22871;
  assign n22873 = pi39 & ~n22868;
  assign n22874 = ~n22872 & n22873;
  assign n22875 = ~pi38 & ~n22864;
  assign n22876 = ~n22874 & n22875;
  assign n22877 = pi700 & ~n22854;
  assign n22878 = ~n22876 & n22877;
  assign n22879 = n9829 & ~n22878;
  assign n22880 = ~n22844 & n22879;
  assign n22881 = ~n22679 & ~n22880;
  assign n22882 = ~pi625 & n22881;
  assign n22883 = pi625 & n22741;
  assign n22884 = ~pi1153 & ~n22883;
  assign n22885 = ~n22882 & n22884;
  assign n22886 = ~pi608 & ~n22697;
  assign n22887 = ~n22885 & n22886;
  assign n22888 = ~pi625 & n22741;
  assign n22889 = pi625 & n22881;
  assign n22890 = pi1153 & ~n22888;
  assign n22891 = ~n22889 & n22890;
  assign n22892 = pi608 & ~n22701;
  assign n22893 = ~n22891 & n22892;
  assign n22894 = ~n22887 & ~n22893;
  assign n22895 = pi778 & ~n22894;
  assign n22896 = ~pi778 & n22881;
  assign n22897 = ~n22895 & ~n22896;
  assign n22898 = ~pi609 & ~n22897;
  assign n22899 = ~pi1155 & ~n22843;
  assign n22900 = ~n22898 & n22899;
  assign n22901 = ~pi660 & ~n22749;
  assign n22902 = ~n22900 & n22901;
  assign n22903 = ~pi609 & n22704;
  assign n22904 = pi609 & ~n22897;
  assign n22905 = pi1155 & ~n22903;
  assign n22906 = ~n22904 & n22905;
  assign n22907 = pi660 & ~n22753;
  assign n22908 = ~n22906 & n22907;
  assign n22909 = ~n22902 & ~n22908;
  assign n22910 = pi785 & ~n22909;
  assign n22911 = ~pi785 & ~n22897;
  assign n22912 = ~n22910 & ~n22911;
  assign n22913 = ~pi618 & ~n22912;
  assign n22914 = ~pi1154 & ~n22842;
  assign n22915 = ~n22913 & n22914;
  assign n22916 = ~pi627 & ~n22761;
  assign n22917 = ~n22915 & n22916;
  assign n22918 = ~pi618 & ~n22707;
  assign n22919 = pi618 & ~n22912;
  assign n22920 = pi1154 & ~n22918;
  assign n22921 = ~n22919 & n22920;
  assign n22922 = pi627 & ~n22765;
  assign n22923 = ~n22921 & n22922;
  assign n22924 = ~n22917 & ~n22923;
  assign n22925 = pi781 & ~n22924;
  assign n22926 = ~pi781 & ~n22912;
  assign n22927 = ~n22925 & ~n22926;
  assign n22928 = ~pi789 & n22927;
  assign n22929 = ~pi619 & n22709;
  assign n22930 = pi619 & ~n22927;
  assign n22931 = pi1159 & ~n22929;
  assign n22932 = ~n22930 & n22931;
  assign n22933 = pi648 & ~n22777;
  assign n22934 = ~n22932 & n22933;
  assign n22935 = ~pi619 & ~n22927;
  assign n22936 = pi619 & n22709;
  assign n22937 = ~pi1159 & ~n22936;
  assign n22938 = ~n22935 & n22937;
  assign n22939 = ~pi648 & ~n22773;
  assign n22940 = ~n22938 & n22939;
  assign n22941 = pi789 & ~n22934;
  assign n22942 = ~n22940 & n22941;
  assign n22943 = n15833 & ~n22928;
  assign n22944 = ~n22942 & n22943;
  assign n22945 = ~n16644 & ~n22841;
  assign n22946 = ~n22944 & n22945;
  assign n22947 = ~n22829 & ~n22946;
  assign n22948 = n18841 & ~n22947;
  assign n22949 = pi644 & ~pi1160;
  assign n22950 = pi644 & ~n22793;
  assign n22951 = ~n22802 & ~n22950;
  assign n22952 = ~n22949 & ~n22951;
  assign n22953 = pi790 & ~n22952;
  assign n22954 = ~n22817 & ~n22948;
  assign n22955 = ~n22953 & n22954;
  assign n22956 = ~n22805 & ~n22955;
  assign n22957 = ~po1038 & ~n22956;
  assign n22958 = ~pi832 & ~n22676;
  assign n22959 = ~n22957 & n22958;
  assign po332 = ~n22675 & ~n22959;
  assign n22961 = ~pi176 & ~n2923;
  assign n22962 = ~pi704 & n15726;
  assign n22963 = ~n22961 & ~n22962;
  assign n22964 = ~pi778 & n22963;
  assign n22965 = ~pi625 & n22962;
  assign n22966 = ~n22963 & ~n22965;
  assign n22967 = pi1153 & ~n22966;
  assign n22968 = ~pi1153 & ~n22961;
  assign n22969 = ~n22965 & n22968;
  assign n22970 = ~n22967 & ~n22969;
  assign n22971 = pi778 & ~n22970;
  assign n22972 = ~n22964 & ~n22971;
  assign n22973 = ~n15742 & n22972;
  assign n22974 = ~n15748 & n22973;
  assign n22975 = ~n15754 & n22974;
  assign n22976 = ~n15760 & n22975;
  assign n22977 = ~n15766 & n22976;
  assign n22978 = n19394 & n22977;
  assign n22979 = ~n19394 & n22961;
  assign n22980 = ~n22978 & ~n22979;
  assign n22981 = ~n15959 & n22980;
  assign n22982 = n15925 & n22961;
  assign n22983 = ~pi742 & n15781;
  assign n22984 = ~n22961 & ~n22983;
  assign n22985 = ~n15778 & ~n22984;
  assign n22986 = ~pi785 & ~n22985;
  assign n22987 = ~n15787 & ~n22984;
  assign n22988 = pi1155 & ~n22987;
  assign n22989 = ~n15790 & n22985;
  assign n22990 = ~pi1155 & ~n22989;
  assign n22991 = ~n22988 & ~n22990;
  assign n22992 = pi785 & ~n22991;
  assign n22993 = ~n22986 & ~n22992;
  assign n22994 = ~pi781 & ~n22993;
  assign n22995 = ~n15797 & n22993;
  assign n22996 = pi1154 & ~n22995;
  assign n22997 = ~n15800 & n22993;
  assign n22998 = ~pi1154 & ~n22997;
  assign n22999 = ~n22996 & ~n22998;
  assign n23000 = pi781 & ~n22999;
  assign n23001 = ~n22994 & ~n23000;
  assign n23002 = ~pi789 & ~n23001;
  assign n23003 = ~pi619 & n22961;
  assign n23004 = pi619 & n23001;
  assign n23005 = pi1159 & ~n23003;
  assign n23006 = ~n23004 & n23005;
  assign n23007 = ~pi619 & n23001;
  assign n23008 = pi619 & n22961;
  assign n23009 = ~pi1159 & ~n23008;
  assign n23010 = ~n23007 & n23009;
  assign n23011 = ~n23006 & ~n23010;
  assign n23012 = pi789 & ~n23011;
  assign n23013 = ~n23002 & ~n23012;
  assign n23014 = ~n15832 & ~n23013;
  assign n23015 = n15832 & ~n22961;
  assign n23016 = ~n23014 & ~n23015;
  assign n23017 = ~n15925 & n23016;
  assign n23018 = n19478 & ~n22982;
  assign n23019 = ~n23017 & n23018;
  assign n23020 = ~n22981 & ~n23019;
  assign n23021 = pi787 & ~n23020;
  assign n23022 = n15828 & n22975;
  assign n23023 = ~pi626 & ~n22961;
  assign n23024 = pi626 & ~n23013;
  assign n23025 = n15756 & ~n23023;
  assign n23026 = ~n23024 & n23025;
  assign n23027 = pi626 & ~n22961;
  assign n23028 = ~pi626 & ~n23013;
  assign n23029 = n15757 & ~n23027;
  assign n23030 = ~n23028 & n23029;
  assign n23031 = ~n23022 & ~n23026;
  assign n23032 = ~n23030 & n23031;
  assign n23033 = pi788 & ~n23032;
  assign n23034 = pi618 & n22973;
  assign n23035 = pi609 & n22972;
  assign n23036 = ~n15780 & ~n22963;
  assign n23037 = pi625 & n23036;
  assign n23038 = n22984 & ~n23036;
  assign n23039 = ~n23037 & ~n23038;
  assign n23040 = n22968 & ~n23039;
  assign n23041 = ~pi608 & ~n22967;
  assign n23042 = ~n23040 & n23041;
  assign n23043 = pi1153 & n22984;
  assign n23044 = ~n23037 & n23043;
  assign n23045 = pi608 & ~n22969;
  assign n23046 = ~n23044 & n23045;
  assign n23047 = ~n23042 & ~n23046;
  assign n23048 = pi778 & ~n23047;
  assign n23049 = ~pi778 & ~n23038;
  assign n23050 = ~n23048 & ~n23049;
  assign n23051 = ~pi609 & ~n23050;
  assign n23052 = ~pi1155 & ~n23035;
  assign n23053 = ~n23051 & n23052;
  assign n23054 = ~pi660 & ~n22988;
  assign n23055 = ~n23053 & n23054;
  assign n23056 = ~pi609 & n22972;
  assign n23057 = pi609 & ~n23050;
  assign n23058 = pi1155 & ~n23056;
  assign n23059 = ~n23057 & n23058;
  assign n23060 = pi660 & ~n22990;
  assign n23061 = ~n23059 & n23060;
  assign n23062 = ~n23055 & ~n23061;
  assign n23063 = pi785 & ~n23062;
  assign n23064 = ~pi785 & ~n23050;
  assign n23065 = ~n23063 & ~n23064;
  assign n23066 = ~pi618 & ~n23065;
  assign n23067 = ~pi1154 & ~n23034;
  assign n23068 = ~n23066 & n23067;
  assign n23069 = ~pi627 & ~n22996;
  assign n23070 = ~n23068 & n23069;
  assign n23071 = ~pi618 & n22973;
  assign n23072 = pi618 & ~n23065;
  assign n23073 = pi1154 & ~n23071;
  assign n23074 = ~n23072 & n23073;
  assign n23075 = pi627 & ~n22998;
  assign n23076 = ~n23074 & n23075;
  assign n23077 = ~n23070 & ~n23076;
  assign n23078 = pi781 & ~n23077;
  assign n23079 = ~pi781 & ~n23065;
  assign n23080 = ~n23078 & ~n23079;
  assign n23081 = ~pi789 & n23080;
  assign n23082 = ~pi619 & n22974;
  assign n23083 = pi619 & ~n23080;
  assign n23084 = pi1159 & ~n23082;
  assign n23085 = ~n23083 & n23084;
  assign n23086 = pi648 & ~n23010;
  assign n23087 = ~n23085 & n23086;
  assign n23088 = pi619 & n22974;
  assign n23089 = ~pi619 & ~n23080;
  assign n23090 = ~pi1159 & ~n23088;
  assign n23091 = ~n23089 & n23090;
  assign n23092 = ~pi648 & ~n23006;
  assign n23093 = ~n23091 & n23092;
  assign n23094 = pi789 & ~n23087;
  assign n23095 = ~n23093 & n23094;
  assign n23096 = n15833 & ~n23081;
  assign n23097 = ~n23095 & n23096;
  assign n23098 = ~n23033 & ~n23097;
  assign n23099 = ~n16644 & ~n23098;
  assign n23100 = n15763 & n23016;
  assign n23101 = n15772 & n22976;
  assign n23102 = ~pi629 & ~n23101;
  assign n23103 = ~n23100 & n23102;
  assign n23104 = n15762 & n23016;
  assign n23105 = n15909 & n22976;
  assign n23106 = pi629 & ~n23105;
  assign n23107 = ~n23104 & n23106;
  assign n23108 = pi792 & ~n23103;
  assign n23109 = ~n23107 & n23108;
  assign n23110 = n18841 & ~n23109;
  assign n23111 = ~n23099 & n23110;
  assign n23112 = ~n23021 & ~n23111;
  assign n23113 = ~pi790 & n23112;
  assign n23114 = pi787 & ~n22980;
  assign n23115 = ~pi787 & n22977;
  assign n23116 = ~n23114 & ~n23115;
  assign n23117 = ~pi644 & ~n23116;
  assign n23118 = pi644 & n23112;
  assign n23119 = pi715 & ~n23117;
  assign n23120 = ~n23118 & n23119;
  assign n23121 = ~n19771 & n22961;
  assign n23122 = ~n15960 & n23017;
  assign n23123 = ~n23121 & ~n23122;
  assign n23124 = pi644 & ~n23123;
  assign n23125 = ~pi644 & n22961;
  assign n23126 = ~pi715 & ~n23125;
  assign n23127 = ~n23124 & n23126;
  assign n23128 = pi1160 & ~n23127;
  assign n23129 = ~n23120 & n23128;
  assign n23130 = ~pi644 & ~n23123;
  assign n23131 = pi644 & n22961;
  assign n23132 = pi715 & ~n23131;
  assign n23133 = ~n23130 & n23132;
  assign n23134 = pi644 & ~n23116;
  assign n23135 = ~pi644 & n23112;
  assign n23136 = ~pi715 & ~n23134;
  assign n23137 = ~n23135 & n23136;
  assign n23138 = ~pi1160 & ~n23133;
  assign n23139 = ~n23137 & n23138;
  assign n23140 = ~n23129 & ~n23139;
  assign n23141 = pi790 & ~n23140;
  assign n23142 = pi832 & ~n23113;
  assign n23143 = ~n23141 & n23142;
  assign n23144 = ~pi176 & po1038;
  assign n23145 = ~pi176 & ~n16219;
  assign n23146 = n15747 & ~n23145;
  assign n23147 = ~n16227 & n19350;
  assign n23148 = pi176 & ~n23147;
  assign n23149 = ~pi38 & ~n17276;
  assign n23150 = ~n19049 & ~n23149;
  assign n23151 = ~pi176 & n23150;
  assign n23152 = ~pi704 & ~n23151;
  assign n23153 = ~pi176 & ~n16218;
  assign n23154 = pi704 & n23153;
  assign n23155 = n9829 & ~n23152;
  assign n23156 = ~n23154 & n23155;
  assign n23157 = ~n23148 & ~n23156;
  assign n23158 = ~pi778 & ~n23157;
  assign n23159 = ~pi625 & n23145;
  assign n23160 = pi625 & n23157;
  assign n23161 = pi1153 & ~n23159;
  assign n23162 = ~n23160 & n23161;
  assign n23163 = ~pi625 & n23157;
  assign n23164 = pi625 & n23145;
  assign n23165 = ~pi1153 & ~n23164;
  assign n23166 = ~n23163 & n23165;
  assign n23167 = ~n23162 & ~n23166;
  assign n23168 = pi778 & ~n23167;
  assign n23169 = ~n23158 & ~n23168;
  assign n23170 = ~n15741 & n23169;
  assign n23171 = n15741 & n23145;
  assign n23172 = ~n23170 & ~n23171;
  assign n23173 = ~n15747 & n23172;
  assign n23174 = ~n23146 & ~n23173;
  assign n23175 = ~n15753 & n23174;
  assign n23176 = n15753 & n23145;
  assign n23177 = ~n23175 & ~n23176;
  assign n23178 = ~n15759 & ~n23177;
  assign n23179 = n15759 & n23145;
  assign n23180 = ~n23178 & ~n23179;
  assign n23181 = ~n15765 & ~n23180;
  assign n23182 = n15765 & n23145;
  assign n23183 = ~n23181 & ~n23182;
  assign n23184 = ~n17768 & ~n23183;
  assign n23185 = n17768 & n23145;
  assign n23186 = ~n23184 & ~n23185;
  assign n23187 = ~pi644 & ~n23186;
  assign n23188 = pi715 & ~n23187;
  assign n23189 = pi176 & ~n9829;
  assign n23190 = ~pi176 & n18604;
  assign n23191 = ~n18598 & ~n18599;
  assign n23192 = pi176 & n23191;
  assign n23193 = ~n23190 & ~n23192;
  assign n23194 = ~pi742 & ~n23193;
  assign n23195 = pi742 & ~n23153;
  assign n23196 = ~n23194 & ~n23195;
  assign n23197 = n9829 & ~n23196;
  assign n23198 = ~n23189 & ~n23197;
  assign n23199 = ~n15777 & ~n23198;
  assign n23200 = n15777 & ~n23145;
  assign n23201 = ~n23199 & ~n23200;
  assign n23202 = ~pi785 & ~n23201;
  assign n23203 = ~n15786 & ~n23145;
  assign n23204 = pi609 & n23199;
  assign n23205 = ~n23203 & ~n23204;
  assign n23206 = pi1155 & ~n23205;
  assign n23207 = ~n16585 & ~n23145;
  assign n23208 = ~pi609 & n23199;
  assign n23209 = ~n23207 & ~n23208;
  assign n23210 = ~pi1155 & ~n23209;
  assign n23211 = ~n23206 & ~n23210;
  assign n23212 = pi785 & ~n23211;
  assign n23213 = ~n23202 & ~n23212;
  assign n23214 = ~pi781 & ~n23213;
  assign n23215 = ~pi618 & n23145;
  assign n23216 = pi618 & n23213;
  assign n23217 = pi1154 & ~n23215;
  assign n23218 = ~n23216 & n23217;
  assign n23219 = ~pi618 & n23213;
  assign n23220 = pi618 & n23145;
  assign n23221 = ~pi1154 & ~n23220;
  assign n23222 = ~n23219 & n23221;
  assign n23223 = ~n23218 & ~n23222;
  assign n23224 = pi781 & ~n23223;
  assign n23225 = ~n23214 & ~n23224;
  assign n23226 = ~pi789 & ~n23225;
  assign n23227 = ~pi619 & n23145;
  assign n23228 = pi619 & n23225;
  assign n23229 = pi1159 & ~n23227;
  assign n23230 = ~n23228 & n23229;
  assign n23231 = ~pi619 & n23225;
  assign n23232 = pi619 & n23145;
  assign n23233 = ~pi1159 & ~n23232;
  assign n23234 = ~n23231 & n23233;
  assign n23235 = ~n23230 & ~n23234;
  assign n23236 = pi789 & ~n23235;
  assign n23237 = ~n23226 & ~n23236;
  assign n23238 = ~n15832 & n23237;
  assign n23239 = n15832 & n23145;
  assign n23240 = ~n23238 & ~n23239;
  assign n23241 = ~n15925 & ~n23240;
  assign n23242 = n15925 & n23145;
  assign n23243 = ~n23241 & ~n23242;
  assign n23244 = ~n15960 & ~n23243;
  assign n23245 = n15960 & n23145;
  assign n23246 = ~n23244 & ~n23245;
  assign n23247 = pi644 & ~n23246;
  assign n23248 = ~pi644 & n23145;
  assign n23249 = ~pi715 & ~n23248;
  assign n23250 = ~n23247 & n23249;
  assign n23251 = pi1160 & ~n23188;
  assign n23252 = ~n23250 & n23251;
  assign n23253 = pi644 & ~n23186;
  assign n23254 = ~pi715 & ~n23253;
  assign n23255 = ~pi644 & ~n23246;
  assign n23256 = pi644 & n23145;
  assign n23257 = pi715 & ~n23256;
  assign n23258 = ~n23255 & n23257;
  assign n23259 = ~pi1160 & ~n23258;
  assign n23260 = ~n23254 & n23259;
  assign n23261 = ~n23252 & ~n23260;
  assign n23262 = pi790 & ~n23261;
  assign n23263 = ~pi647 & n23145;
  assign n23264 = pi647 & ~n23183;
  assign n23265 = n15957 & ~n23263;
  assign n23266 = ~n23264 & n23265;
  assign n23267 = n19478 & n23243;
  assign n23268 = pi647 & n23145;
  assign n23269 = ~pi647 & ~n23183;
  assign n23270 = n15958 & ~n23268;
  assign n23271 = ~n23269 & n23270;
  assign n23272 = ~n23266 & ~n23271;
  assign n23273 = ~n23267 & n23272;
  assign n23274 = pi787 & ~n23273;
  assign n23275 = pi644 & ~n23250;
  assign n23276 = ~n23259 & ~n23275;
  assign n23277 = ~n22949 & ~n23276;
  assign n23278 = pi790 & ~n23277;
  assign n23279 = pi628 & n23145;
  assign n23280 = ~pi628 & ~n23180;
  assign n23281 = n15923 & ~n23279;
  assign n23282 = ~n23280 & n23281;
  assign n23283 = ~n16633 & n23240;
  assign n23284 = ~pi628 & n23145;
  assign n23285 = pi628 & ~n23180;
  assign n23286 = n15922 & ~n23284;
  assign n23287 = ~n23285 & n23286;
  assign n23288 = ~n23282 & ~n23287;
  assign n23289 = ~n23283 & n23288;
  assign n23290 = n16644 & n23289;
  assign n23291 = pi792 & ~n23289;
  assign n23292 = n15828 & ~n23177;
  assign n23293 = ~pi626 & ~n23145;
  assign n23294 = pi626 & ~n23237;
  assign n23295 = n15756 & ~n23293;
  assign n23296 = ~n23294 & n23295;
  assign n23297 = pi626 & ~n23145;
  assign n23298 = ~pi626 & ~n23237;
  assign n23299 = n15757 & ~n23297;
  assign n23300 = ~n23298 & n23299;
  assign n23301 = ~n23292 & ~n23296;
  assign n23302 = ~n23300 & n23301;
  assign n23303 = pi788 & ~n23302;
  assign n23304 = pi618 & ~n23172;
  assign n23305 = pi609 & n23169;
  assign n23306 = pi704 & n23196;
  assign n23307 = ~pi176 & ~n18675;
  assign n23308 = ~n18666 & ~n18668;
  assign n23309 = pi176 & n23308;
  assign n23310 = pi742 & ~n23309;
  assign n23311 = ~n23307 & n23310;
  assign n23312 = ~pi176 & n18651;
  assign n23313 = pi176 & ~n18659;
  assign n23314 = ~pi742 & ~n23312;
  assign n23315 = ~n23313 & n23314;
  assign n23316 = ~n23311 & ~n23315;
  assign n23317 = ~pi704 & ~n23316;
  assign n23318 = n9829 & ~n23306;
  assign n23319 = ~n23317 & n23318;
  assign n23320 = ~n23189 & ~n23319;
  assign n23321 = ~pi625 & n23320;
  assign n23322 = pi625 & n23198;
  assign n23323 = ~pi1153 & ~n23322;
  assign n23324 = ~n23321 & n23323;
  assign n23325 = ~pi608 & ~n23162;
  assign n23326 = ~n23324 & n23325;
  assign n23327 = ~pi625 & n23198;
  assign n23328 = pi625 & n23320;
  assign n23329 = pi1153 & ~n23327;
  assign n23330 = ~n23328 & n23329;
  assign n23331 = pi608 & ~n23166;
  assign n23332 = ~n23330 & n23331;
  assign n23333 = ~n23326 & ~n23332;
  assign n23334 = pi778 & ~n23333;
  assign n23335 = ~pi778 & n23320;
  assign n23336 = ~n23334 & ~n23335;
  assign n23337 = ~pi609 & ~n23336;
  assign n23338 = ~pi1155 & ~n23305;
  assign n23339 = ~n23337 & n23338;
  assign n23340 = ~pi660 & ~n23206;
  assign n23341 = ~n23339 & n23340;
  assign n23342 = ~pi609 & n23169;
  assign n23343 = pi609 & ~n23336;
  assign n23344 = pi1155 & ~n23342;
  assign n23345 = ~n23343 & n23344;
  assign n23346 = pi660 & ~n23210;
  assign n23347 = ~n23345 & n23346;
  assign n23348 = ~n23341 & ~n23347;
  assign n23349 = pi785 & ~n23348;
  assign n23350 = ~pi785 & ~n23336;
  assign n23351 = ~n23349 & ~n23350;
  assign n23352 = ~pi618 & ~n23351;
  assign n23353 = ~pi1154 & ~n23304;
  assign n23354 = ~n23352 & n23353;
  assign n23355 = ~pi627 & ~n23218;
  assign n23356 = ~n23354 & n23355;
  assign n23357 = ~pi618 & ~n23172;
  assign n23358 = pi618 & ~n23351;
  assign n23359 = pi1154 & ~n23357;
  assign n23360 = ~n23358 & n23359;
  assign n23361 = pi627 & ~n23222;
  assign n23362 = ~n23360 & n23361;
  assign n23363 = ~n23356 & ~n23362;
  assign n23364 = pi781 & ~n23363;
  assign n23365 = ~pi781 & ~n23351;
  assign n23366 = ~n23364 & ~n23365;
  assign n23367 = ~pi789 & n23366;
  assign n23368 = ~pi619 & n23174;
  assign n23369 = pi619 & ~n23366;
  assign n23370 = pi1159 & ~n23368;
  assign n23371 = ~n23369 & n23370;
  assign n23372 = pi648 & ~n23234;
  assign n23373 = ~n23371 & n23372;
  assign n23374 = ~pi619 & ~n23366;
  assign n23375 = pi619 & n23174;
  assign n23376 = ~pi1159 & ~n23375;
  assign n23377 = ~n23374 & n23376;
  assign n23378 = ~pi648 & ~n23230;
  assign n23379 = ~n23377 & n23378;
  assign n23380 = pi789 & ~n23373;
  assign n23381 = ~n23379 & n23380;
  assign n23382 = n15833 & ~n23367;
  assign n23383 = ~n23381 & n23382;
  assign n23384 = ~n23303 & ~n23383;
  assign n23385 = ~n23291 & ~n23384;
  assign n23386 = n18841 & ~n23290;
  assign n23387 = ~n23385 & n23386;
  assign n23388 = ~n23274 & ~n23278;
  assign n23389 = ~n23387 & n23388;
  assign n23390 = ~n23262 & ~n23389;
  assign n23391 = ~po1038 & ~n23390;
  assign n23392 = ~pi832 & ~n23144;
  assign n23393 = ~n23391 & n23392;
  assign po333 = ~n23143 & ~n23393;
  assign n23395 = ~pi177 & ~n2923;
  assign n23396 = ~pi686 & n15726;
  assign n23397 = ~n23395 & ~n23396;
  assign n23398 = ~pi778 & n23397;
  assign n23399 = ~pi625 & n23396;
  assign n23400 = ~n23397 & ~n23399;
  assign n23401 = pi1153 & ~n23400;
  assign n23402 = ~pi1153 & ~n23395;
  assign n23403 = ~n23399 & n23402;
  assign n23404 = ~n23401 & ~n23403;
  assign n23405 = pi778 & ~n23404;
  assign n23406 = ~n23398 & ~n23405;
  assign n23407 = ~n15742 & n23406;
  assign n23408 = ~n15748 & n23407;
  assign n23409 = ~n15754 & n23408;
  assign n23410 = ~n15760 & n23409;
  assign n23411 = ~n15766 & n23410;
  assign n23412 = n19394 & n23411;
  assign n23413 = ~n19394 & n23395;
  assign n23414 = ~n23412 & ~n23413;
  assign n23415 = ~n15959 & n23414;
  assign n23416 = n15925 & n23395;
  assign n23417 = ~pi757 & n15781;
  assign n23418 = ~n23395 & ~n23417;
  assign n23419 = ~n15778 & ~n23418;
  assign n23420 = ~pi785 & ~n23419;
  assign n23421 = ~n15787 & ~n23418;
  assign n23422 = pi1155 & ~n23421;
  assign n23423 = ~n15790 & n23419;
  assign n23424 = ~pi1155 & ~n23423;
  assign n23425 = ~n23422 & ~n23424;
  assign n23426 = pi785 & ~n23425;
  assign n23427 = ~n23420 & ~n23426;
  assign n23428 = ~pi781 & ~n23427;
  assign n23429 = ~n15797 & n23427;
  assign n23430 = pi1154 & ~n23429;
  assign n23431 = ~n15800 & n23427;
  assign n23432 = ~pi1154 & ~n23431;
  assign n23433 = ~n23430 & ~n23432;
  assign n23434 = pi781 & ~n23433;
  assign n23435 = ~n23428 & ~n23434;
  assign n23436 = ~pi789 & ~n23435;
  assign n23437 = ~pi619 & n23395;
  assign n23438 = pi619 & n23435;
  assign n23439 = pi1159 & ~n23437;
  assign n23440 = ~n23438 & n23439;
  assign n23441 = ~pi619 & n23435;
  assign n23442 = pi619 & n23395;
  assign n23443 = ~pi1159 & ~n23442;
  assign n23444 = ~n23441 & n23443;
  assign n23445 = ~n23440 & ~n23444;
  assign n23446 = pi789 & ~n23445;
  assign n23447 = ~n23436 & ~n23446;
  assign n23448 = ~n15832 & ~n23447;
  assign n23449 = n15832 & ~n23395;
  assign n23450 = ~n23448 & ~n23449;
  assign n23451 = ~n15925 & n23450;
  assign n23452 = n19478 & ~n23416;
  assign n23453 = ~n23451 & n23452;
  assign n23454 = ~n23415 & ~n23453;
  assign n23455 = pi787 & ~n23454;
  assign n23456 = n15828 & n23409;
  assign n23457 = ~pi626 & ~n23395;
  assign n23458 = pi626 & ~n23447;
  assign n23459 = n15756 & ~n23457;
  assign n23460 = ~n23458 & n23459;
  assign n23461 = pi626 & ~n23395;
  assign n23462 = ~pi626 & ~n23447;
  assign n23463 = n15757 & ~n23461;
  assign n23464 = ~n23462 & n23463;
  assign n23465 = ~n23456 & ~n23460;
  assign n23466 = ~n23464 & n23465;
  assign n23467 = pi788 & ~n23466;
  assign n23468 = pi618 & n23407;
  assign n23469 = pi609 & n23406;
  assign n23470 = ~n15780 & ~n23397;
  assign n23471 = pi625 & n23470;
  assign n23472 = n23418 & ~n23470;
  assign n23473 = ~n23471 & ~n23472;
  assign n23474 = n23402 & ~n23473;
  assign n23475 = ~pi608 & ~n23401;
  assign n23476 = ~n23474 & n23475;
  assign n23477 = pi1153 & n23418;
  assign n23478 = ~n23471 & n23477;
  assign n23479 = pi608 & ~n23403;
  assign n23480 = ~n23478 & n23479;
  assign n23481 = ~n23476 & ~n23480;
  assign n23482 = pi778 & ~n23481;
  assign n23483 = ~pi778 & ~n23472;
  assign n23484 = ~n23482 & ~n23483;
  assign n23485 = ~pi609 & ~n23484;
  assign n23486 = ~pi1155 & ~n23469;
  assign n23487 = ~n23485 & n23486;
  assign n23488 = ~pi660 & ~n23422;
  assign n23489 = ~n23487 & n23488;
  assign n23490 = ~pi609 & n23406;
  assign n23491 = pi609 & ~n23484;
  assign n23492 = pi1155 & ~n23490;
  assign n23493 = ~n23491 & n23492;
  assign n23494 = pi660 & ~n23424;
  assign n23495 = ~n23493 & n23494;
  assign n23496 = ~n23489 & ~n23495;
  assign n23497 = pi785 & ~n23496;
  assign n23498 = ~pi785 & ~n23484;
  assign n23499 = ~n23497 & ~n23498;
  assign n23500 = ~pi618 & ~n23499;
  assign n23501 = ~pi1154 & ~n23468;
  assign n23502 = ~n23500 & n23501;
  assign n23503 = ~pi627 & ~n23430;
  assign n23504 = ~n23502 & n23503;
  assign n23505 = ~pi618 & n23407;
  assign n23506 = pi618 & ~n23499;
  assign n23507 = pi1154 & ~n23505;
  assign n23508 = ~n23506 & n23507;
  assign n23509 = pi627 & ~n23432;
  assign n23510 = ~n23508 & n23509;
  assign n23511 = ~n23504 & ~n23510;
  assign n23512 = pi781 & ~n23511;
  assign n23513 = ~pi781 & ~n23499;
  assign n23514 = ~n23512 & ~n23513;
  assign n23515 = ~pi789 & n23514;
  assign n23516 = ~pi619 & n23408;
  assign n23517 = pi619 & ~n23514;
  assign n23518 = pi1159 & ~n23516;
  assign n23519 = ~n23517 & n23518;
  assign n23520 = pi648 & ~n23444;
  assign n23521 = ~n23519 & n23520;
  assign n23522 = pi619 & n23408;
  assign n23523 = ~pi619 & ~n23514;
  assign n23524 = ~pi1159 & ~n23522;
  assign n23525 = ~n23523 & n23524;
  assign n23526 = ~pi648 & ~n23440;
  assign n23527 = ~n23525 & n23526;
  assign n23528 = pi789 & ~n23521;
  assign n23529 = ~n23527 & n23528;
  assign n23530 = n15833 & ~n23515;
  assign n23531 = ~n23529 & n23530;
  assign n23532 = ~n23467 & ~n23531;
  assign n23533 = ~n16644 & ~n23532;
  assign n23534 = n15763 & n23450;
  assign n23535 = n15772 & n23410;
  assign n23536 = ~pi629 & ~n23535;
  assign n23537 = ~n23534 & n23536;
  assign n23538 = n15762 & n23450;
  assign n23539 = n15909 & n23410;
  assign n23540 = pi629 & ~n23539;
  assign n23541 = ~n23538 & n23540;
  assign n23542 = pi792 & ~n23537;
  assign n23543 = ~n23541 & n23542;
  assign n23544 = n18841 & ~n23543;
  assign n23545 = ~n23533 & n23544;
  assign n23546 = ~n23455 & ~n23545;
  assign n23547 = ~pi790 & n23546;
  assign n23548 = pi787 & ~n23414;
  assign n23549 = ~pi787 & n23411;
  assign n23550 = ~n23548 & ~n23549;
  assign n23551 = ~pi644 & ~n23550;
  assign n23552 = pi644 & n23546;
  assign n23553 = pi715 & ~n23551;
  assign n23554 = ~n23552 & n23553;
  assign n23555 = ~n19771 & n23395;
  assign n23556 = ~n15960 & n23451;
  assign n23557 = ~n23555 & ~n23556;
  assign n23558 = pi644 & ~n23557;
  assign n23559 = ~pi644 & n23395;
  assign n23560 = ~pi715 & ~n23559;
  assign n23561 = ~n23558 & n23560;
  assign n23562 = pi1160 & ~n23561;
  assign n23563 = ~n23554 & n23562;
  assign n23564 = ~pi644 & ~n23557;
  assign n23565 = pi644 & n23395;
  assign n23566 = pi715 & ~n23565;
  assign n23567 = ~n23564 & n23566;
  assign n23568 = pi644 & ~n23550;
  assign n23569 = ~pi644 & n23546;
  assign n23570 = ~pi715 & ~n23568;
  assign n23571 = ~n23569 & n23570;
  assign n23572 = ~pi1160 & ~n23567;
  assign n23573 = ~n23571 & n23572;
  assign n23574 = ~n23563 & ~n23573;
  assign n23575 = pi790 & ~n23574;
  assign n23576 = pi832 & ~n23547;
  assign n23577 = ~n23575 & n23576;
  assign n23578 = ~pi177 & po1038;
  assign n23579 = ~pi177 & ~n16219;
  assign n23580 = n15759 & ~n23579;
  assign n23581 = n15747 & ~n23579;
  assign n23582 = pi177 & ~n9829;
  assign n23583 = pi177 & n17272;
  assign n23584 = ~pi177 & ~n17276;
  assign n23585 = ~pi38 & ~n23583;
  assign n23586 = ~n23584 & n23585;
  assign n23587 = ~pi177 & ~n16228;
  assign n23588 = n16227 & ~n23587;
  assign n23589 = ~pi686 & ~n23588;
  assign n23590 = ~n23586 & n23589;
  assign n23591 = ~pi177 & pi686;
  assign n23592 = ~n16218 & n23591;
  assign n23593 = n9829 & ~n23590;
  assign n23594 = ~n23592 & n23593;
  assign n23595 = ~n23582 & ~n23594;
  assign n23596 = ~pi778 & ~n23595;
  assign n23597 = ~pi625 & n23579;
  assign n23598 = pi625 & n23595;
  assign n23599 = pi1153 & ~n23597;
  assign n23600 = ~n23598 & n23599;
  assign n23601 = ~pi625 & n23595;
  assign n23602 = pi625 & n23579;
  assign n23603 = ~pi1153 & ~n23602;
  assign n23604 = ~n23601 & n23603;
  assign n23605 = ~n23600 & ~n23604;
  assign n23606 = pi778 & ~n23605;
  assign n23607 = ~n23596 & ~n23606;
  assign n23608 = ~n15741 & n23607;
  assign n23609 = n15741 & n23579;
  assign n23610 = ~n23608 & ~n23609;
  assign n23611 = ~n15747 & n23610;
  assign n23612 = ~n23581 & ~n23611;
  assign n23613 = ~n15753 & n23612;
  assign n23614 = n15753 & n23579;
  assign n23615 = ~n23613 & ~n23614;
  assign n23616 = ~n15759 & n23615;
  assign n23617 = ~n23580 & ~n23616;
  assign n23618 = ~pi792 & ~n23617;
  assign n23619 = ~pi628 & ~n23579;
  assign n23620 = pi628 & ~n23617;
  assign n23621 = ~n23619 & ~n23620;
  assign n23622 = pi1156 & ~n23621;
  assign n23623 = ~pi628 & n23617;
  assign n23624 = pi628 & n23579;
  assign n23625 = ~pi1156 & ~n23624;
  assign n23626 = ~n23623 & n23625;
  assign n23627 = ~n23622 & ~n23626;
  assign n23628 = pi792 & ~n23627;
  assign n23629 = ~n23618 & ~n23628;
  assign n23630 = ~pi787 & ~n23629;
  assign n23631 = ~pi647 & n23579;
  assign n23632 = pi647 & n23629;
  assign n23633 = pi1157 & ~n23631;
  assign n23634 = ~n23632 & n23633;
  assign n23635 = ~pi647 & n23629;
  assign n23636 = pi647 & n23579;
  assign n23637 = ~pi1157 & ~n23636;
  assign n23638 = ~n23635 & n23637;
  assign n23639 = ~n23634 & ~n23638;
  assign n23640 = pi787 & ~n23639;
  assign n23641 = ~n23630 & ~n23640;
  assign n23642 = ~pi644 & n23641;
  assign n23643 = ~pi629 & n23622;
  assign n23644 = ~pi757 & ~n18604;
  assign n23645 = ~n20519 & ~n23644;
  assign n23646 = ~pi177 & ~n23645;
  assign n23647 = ~pi177 & ~n18598;
  assign n23648 = ~pi757 & ~n23647;
  assign n23649 = ~n23191 & n23648;
  assign n23650 = ~n23646 & ~n23649;
  assign n23651 = n9829 & n23650;
  assign n23652 = ~n23582 & ~n23651;
  assign n23653 = ~n15777 & ~n23652;
  assign n23654 = n15777 & ~n23579;
  assign n23655 = ~n23653 & ~n23654;
  assign n23656 = ~pi785 & ~n23655;
  assign n23657 = ~n15786 & ~n23579;
  assign n23658 = pi609 & n23653;
  assign n23659 = ~n23657 & ~n23658;
  assign n23660 = pi1155 & ~n23659;
  assign n23661 = ~n16585 & ~n23579;
  assign n23662 = ~pi609 & n23653;
  assign n23663 = ~n23661 & ~n23662;
  assign n23664 = ~pi1155 & ~n23663;
  assign n23665 = ~n23660 & ~n23664;
  assign n23666 = pi785 & ~n23665;
  assign n23667 = ~n23656 & ~n23666;
  assign n23668 = ~pi781 & ~n23667;
  assign n23669 = ~pi618 & n23579;
  assign n23670 = pi618 & n23667;
  assign n23671 = pi1154 & ~n23669;
  assign n23672 = ~n23670 & n23671;
  assign n23673 = ~pi618 & n23667;
  assign n23674 = pi618 & n23579;
  assign n23675 = ~pi1154 & ~n23674;
  assign n23676 = ~n23673 & n23675;
  assign n23677 = ~n23672 & ~n23676;
  assign n23678 = pi781 & ~n23677;
  assign n23679 = ~n23668 & ~n23678;
  assign n23680 = ~pi789 & ~n23679;
  assign n23681 = ~pi619 & n23579;
  assign n23682 = pi619 & n23679;
  assign n23683 = pi1159 & ~n23681;
  assign n23684 = ~n23682 & n23683;
  assign n23685 = ~pi619 & n23679;
  assign n23686 = pi619 & n23579;
  assign n23687 = ~pi1159 & ~n23686;
  assign n23688 = ~n23685 & n23687;
  assign n23689 = ~n23684 & ~n23688;
  assign n23690 = pi789 & ~n23689;
  assign n23691 = ~n23680 & ~n23690;
  assign n23692 = ~n15832 & n23691;
  assign n23693 = n15832 & n23579;
  assign n23694 = ~n23692 & ~n23693;
  assign n23695 = ~n16633 & n23694;
  assign n23696 = pi629 & n23626;
  assign n23697 = ~n23643 & ~n23696;
  assign n23698 = ~n23695 & n23697;
  assign n23699 = pi792 & ~n23698;
  assign n23700 = pi619 & n23612;
  assign n23701 = ~pi1159 & ~n23700;
  assign n23702 = ~pi648 & ~n23684;
  assign n23703 = ~n23701 & n23702;
  assign n23704 = pi618 & ~n23610;
  assign n23705 = pi609 & n23607;
  assign n23706 = n17390 & ~n23587;
  assign n23707 = pi177 & n18665;
  assign n23708 = ~pi177 & ~n18673;
  assign n23709 = ~pi38 & ~n23707;
  assign n23710 = ~n23708 & n23709;
  assign n23711 = pi757 & ~n23706;
  assign n23712 = ~n23710 & n23711;
  assign n23713 = n18654 & ~n23587;
  assign n23714 = ~n18645 & ~n18647;
  assign n23715 = ~pi177 & ~n23714;
  assign n23716 = pi177 & n18657;
  assign n23717 = ~pi38 & ~n23715;
  assign n23718 = ~n23716 & n23717;
  assign n23719 = ~pi757 & ~n23713;
  assign n23720 = ~n23718 & n23719;
  assign n23721 = ~n23712 & ~n23720;
  assign n23722 = ~pi686 & ~n23721;
  assign n23723 = pi686 & ~n23650;
  assign n23724 = n9829 & ~n23722;
  assign n23725 = ~n23723 & n23724;
  assign n23726 = ~n23582 & ~n23725;
  assign n23727 = ~pi625 & n23726;
  assign n23728 = pi625 & n23652;
  assign n23729 = ~pi1153 & ~n23728;
  assign n23730 = ~n23727 & n23729;
  assign n23731 = ~pi608 & ~n23600;
  assign n23732 = ~n23730 & n23731;
  assign n23733 = ~pi625 & n23652;
  assign n23734 = pi625 & n23726;
  assign n23735 = pi1153 & ~n23733;
  assign n23736 = ~n23734 & n23735;
  assign n23737 = pi608 & ~n23604;
  assign n23738 = ~n23736 & n23737;
  assign n23739 = ~n23732 & ~n23738;
  assign n23740 = pi778 & ~n23739;
  assign n23741 = ~pi778 & n23726;
  assign n23742 = ~n23740 & ~n23741;
  assign n23743 = ~pi609 & ~n23742;
  assign n23744 = ~pi1155 & ~n23705;
  assign n23745 = ~n23743 & n23744;
  assign n23746 = ~pi660 & ~n23660;
  assign n23747 = ~n23745 & n23746;
  assign n23748 = ~pi609 & n23607;
  assign n23749 = pi609 & ~n23742;
  assign n23750 = pi1155 & ~n23748;
  assign n23751 = ~n23749 & n23750;
  assign n23752 = pi660 & ~n23664;
  assign n23753 = ~n23751 & n23752;
  assign n23754 = ~n23747 & ~n23753;
  assign n23755 = pi785 & ~n23754;
  assign n23756 = ~pi785 & ~n23742;
  assign n23757 = ~n23755 & ~n23756;
  assign n23758 = ~pi618 & ~n23757;
  assign n23759 = ~pi1154 & ~n23704;
  assign n23760 = ~n23758 & n23759;
  assign n23761 = ~pi627 & ~n23672;
  assign n23762 = ~n23760 & n23761;
  assign n23763 = ~pi618 & ~n23610;
  assign n23764 = pi618 & ~n23757;
  assign n23765 = pi1154 & ~n23763;
  assign n23766 = ~n23764 & n23765;
  assign n23767 = pi627 & ~n23676;
  assign n23768 = ~n23766 & n23767;
  assign n23769 = ~n23762 & ~n23768;
  assign n23770 = pi781 & ~n23769;
  assign n23771 = ~pi781 & ~n23757;
  assign n23772 = ~n23770 & ~n23771;
  assign n23773 = pi619 & ~n23772;
  assign n23774 = ~pi619 & n23612;
  assign n23775 = pi1159 & ~n23774;
  assign n23776 = ~n23773 & n23775;
  assign n23777 = pi648 & ~n23688;
  assign n23778 = ~n23776 & n23777;
  assign n23779 = ~n23703 & ~n23778;
  assign n23780 = pi789 & ~n23779;
  assign n23781 = ~pi619 & n23702;
  assign n23782 = pi789 & ~n23781;
  assign n23783 = ~n23772 & ~n23782;
  assign n23784 = ~n23780 & ~n23783;
  assign n23785 = n15833 & ~n23784;
  assign n23786 = pi641 & ~n23579;
  assign n23787 = ~pi641 & n23615;
  assign n23788 = n15819 & ~n23786;
  assign n23789 = ~n23787 & n23788;
  assign n23790 = n22348 & n23691;
  assign n23791 = ~pi641 & ~n23579;
  assign n23792 = pi641 & n23615;
  assign n23793 = n15818 & ~n23791;
  assign n23794 = ~n23792 & n23793;
  assign n23795 = ~n23789 & ~n23794;
  assign n23796 = ~n23790 & n23795;
  assign n23797 = pi788 & ~n23796;
  assign n23798 = ~n16644 & ~n23797;
  assign n23799 = ~n23785 & n23798;
  assign n23800 = ~n23699 & ~n23799;
  assign n23801 = ~pi647 & n23800;
  assign n23802 = ~n15925 & ~n23694;
  assign n23803 = n15925 & n23579;
  assign n23804 = ~n23802 & ~n23803;
  assign n23805 = pi647 & ~n23804;
  assign n23806 = ~pi1157 & ~n23805;
  assign n23807 = ~n23801 & n23806;
  assign n23808 = ~pi630 & ~n23634;
  assign n23809 = ~n23807 & n23808;
  assign n23810 = ~pi647 & ~n23804;
  assign n23811 = pi647 & n23800;
  assign n23812 = pi1157 & ~n23810;
  assign n23813 = ~n23811 & n23812;
  assign n23814 = pi630 & ~n23638;
  assign n23815 = ~n23813 & n23814;
  assign n23816 = ~n23809 & ~n23815;
  assign n23817 = pi787 & ~n23816;
  assign n23818 = ~pi787 & n23800;
  assign n23819 = ~n23817 & ~n23818;
  assign n23820 = pi644 & ~n23819;
  assign n23821 = pi715 & ~n23642;
  assign n23822 = ~n23820 & n23821;
  assign n23823 = ~n15960 & ~n23804;
  assign n23824 = n15960 & n23579;
  assign n23825 = ~n23823 & ~n23824;
  assign n23826 = pi644 & ~n23825;
  assign n23827 = ~pi644 & n23579;
  assign n23828 = ~pi715 & ~n23827;
  assign n23829 = ~n23826 & n23828;
  assign n23830 = pi1160 & ~n23829;
  assign n23831 = ~n23822 & n23830;
  assign n23832 = pi644 & n23641;
  assign n23833 = ~pi715 & ~n23832;
  assign n23834 = ~pi644 & ~n23825;
  assign n23835 = pi644 & n23579;
  assign n23836 = pi715 & ~n23835;
  assign n23837 = ~n23834 & n23836;
  assign n23838 = ~pi1160 & ~n23837;
  assign n23839 = ~n23833 & n23838;
  assign n23840 = ~n23831 & ~n23839;
  assign n23841 = pi790 & ~n23840;
  assign n23842 = ~pi644 & n23838;
  assign n23843 = pi790 & ~n23842;
  assign n23844 = ~n23819 & ~n23843;
  assign n23845 = ~n23841 & ~n23844;
  assign n23846 = ~po1038 & ~n23845;
  assign n23847 = ~pi832 & ~n23578;
  assign n23848 = ~n23846 & n23847;
  assign po334 = ~n23577 & ~n23848;
  assign n23850 = ~pi178 & ~n2923;
  assign n23851 = ~pi688 & n15726;
  assign n23852 = ~n23850 & ~n23851;
  assign n23853 = ~pi778 & ~n23852;
  assign n23854 = ~pi625 & n23851;
  assign n23855 = ~n23852 & ~n23854;
  assign n23856 = pi1153 & ~n23855;
  assign n23857 = ~pi1153 & ~n23850;
  assign n23858 = ~n23854 & n23857;
  assign n23859 = pi778 & ~n23858;
  assign n23860 = ~n23856 & n23859;
  assign n23861 = ~n23853 & ~n23860;
  assign n23862 = ~n15742 & ~n23861;
  assign n23863 = ~n15748 & n23862;
  assign n23864 = ~n15754 & n23863;
  assign n23865 = ~n15760 & n23864;
  assign n23866 = ~n15766 & n23865;
  assign n23867 = n19394 & n23866;
  assign n23868 = ~n19394 & n23850;
  assign n23869 = ~n23867 & ~n23868;
  assign n23870 = ~n15959 & n23869;
  assign n23871 = n15925 & n23850;
  assign n23872 = ~pi760 & n15781;
  assign n23873 = ~n23850 & ~n23872;
  assign n23874 = ~n15778 & ~n23873;
  assign n23875 = ~pi785 & ~n23874;
  assign n23876 = n16585 & n23872;
  assign n23877 = n23874 & ~n23876;
  assign n23878 = pi1155 & ~n23877;
  assign n23879 = ~pi1155 & ~n23850;
  assign n23880 = ~n23876 & n23879;
  assign n23881 = ~n23878 & ~n23880;
  assign n23882 = pi785 & ~n23881;
  assign n23883 = ~n23875 & ~n23882;
  assign n23884 = ~pi781 & ~n23883;
  assign n23885 = ~n15797 & n23883;
  assign n23886 = pi1154 & ~n23885;
  assign n23887 = ~n15800 & n23883;
  assign n23888 = ~pi1154 & ~n23887;
  assign n23889 = ~n23886 & ~n23888;
  assign n23890 = pi781 & ~n23889;
  assign n23891 = ~n23884 & ~n23890;
  assign n23892 = ~n21915 & n23891;
  assign n23893 = ~n15832 & ~n23892;
  assign n23894 = n15832 & ~n23850;
  assign n23895 = ~n23893 & ~n23894;
  assign n23896 = ~n15925 & n23895;
  assign n23897 = n19478 & ~n23871;
  assign n23898 = ~n23896 & n23897;
  assign n23899 = ~n23870 & ~n23898;
  assign n23900 = pi787 & ~n23899;
  assign n23901 = n15763 & n23895;
  assign n23902 = n15772 & n23865;
  assign n23903 = ~pi629 & ~n23902;
  assign n23904 = ~n23901 & n23903;
  assign n23905 = n15762 & n23895;
  assign n23906 = n15909 & n23865;
  assign n23907 = pi629 & ~n23906;
  assign n23908 = ~n23905 & n23907;
  assign n23909 = pi792 & ~n23904;
  assign n23910 = ~n23908 & n23909;
  assign n23911 = ~n21932 & n23891;
  assign n23912 = pi648 & ~n23911;
  assign n23913 = n21935 & ~n23863;
  assign n23914 = ~n23912 & ~n23913;
  assign n23915 = ~pi1159 & ~n23914;
  assign n23916 = ~pi619 & ~n23863;
  assign n23917 = pi648 & ~n23916;
  assign n23918 = n21942 & n23891;
  assign n23919 = pi1159 & ~n23917;
  assign n23920 = ~n23918 & n23919;
  assign n23921 = ~n23915 & ~n23920;
  assign n23922 = pi789 & ~n23921;
  assign n23923 = pi609 & ~n23861;
  assign n23924 = ~n15780 & ~n23852;
  assign n23925 = pi625 & n23924;
  assign n23926 = n23873 & ~n23924;
  assign n23927 = ~n23925 & ~n23926;
  assign n23928 = n23857 & ~n23927;
  assign n23929 = ~pi608 & ~n23856;
  assign n23930 = ~n23928 & n23929;
  assign n23931 = pi1153 & n23873;
  assign n23932 = ~n23925 & n23931;
  assign n23933 = pi608 & ~n23858;
  assign n23934 = ~n23932 & n23933;
  assign n23935 = ~n23930 & ~n23934;
  assign n23936 = pi778 & ~n23935;
  assign n23937 = ~pi778 & ~n23926;
  assign n23938 = ~n23936 & ~n23937;
  assign n23939 = ~pi609 & ~n23938;
  assign n23940 = ~pi1155 & ~n23923;
  assign n23941 = ~n23939 & n23940;
  assign n23942 = ~pi660 & ~n23878;
  assign n23943 = ~n23941 & n23942;
  assign n23944 = ~pi609 & ~n23861;
  assign n23945 = pi609 & ~n23938;
  assign n23946 = pi1155 & ~n23944;
  assign n23947 = ~n23945 & n23946;
  assign n23948 = pi660 & ~n23880;
  assign n23949 = ~n23947 & n23948;
  assign n23950 = ~n23943 & ~n23949;
  assign n23951 = pi785 & ~n23950;
  assign n23952 = ~pi785 & ~n23938;
  assign n23953 = ~n23951 & ~n23952;
  assign n23954 = ~pi781 & n23953;
  assign n23955 = pi618 & n23862;
  assign n23956 = ~pi618 & ~n23953;
  assign n23957 = ~pi1154 & ~n23955;
  assign n23958 = ~n23956 & n23957;
  assign n23959 = ~pi627 & ~n23886;
  assign n23960 = ~n23958 & n23959;
  assign n23961 = ~pi618 & n23862;
  assign n23962 = pi618 & ~n23953;
  assign n23963 = pi1154 & ~n23961;
  assign n23964 = ~n23962 & n23963;
  assign n23965 = pi627 & ~n23888;
  assign n23966 = ~n23964 & n23965;
  assign n23967 = pi781 & ~n23960;
  assign n23968 = ~n23966 & n23967;
  assign n23969 = ~n23922 & ~n23954;
  assign n23970 = ~n23968 & n23969;
  assign n23971 = n18969 & n23921;
  assign n23972 = ~n23970 & ~n23971;
  assign n23973 = n15833 & ~n23972;
  assign n23974 = n15828 & n23864;
  assign n23975 = ~pi626 & ~n23850;
  assign n23976 = pi626 & ~n23892;
  assign n23977 = n15756 & ~n23975;
  assign n23978 = ~n23976 & n23977;
  assign n23979 = pi626 & ~n23850;
  assign n23980 = ~pi626 & ~n23892;
  assign n23981 = n15757 & ~n23979;
  assign n23982 = ~n23980 & n23981;
  assign n23983 = ~n23974 & ~n23978;
  assign n23984 = ~n23982 & n23983;
  assign n23985 = pi788 & ~n23984;
  assign n23986 = ~n23973 & ~n23985;
  assign n23987 = ~n16644 & ~n23986;
  assign n23988 = n18841 & ~n23910;
  assign n23989 = ~n23987 & n23988;
  assign n23990 = ~n23900 & ~n23989;
  assign n23991 = ~pi790 & n23990;
  assign n23992 = pi787 & ~n23869;
  assign n23993 = ~pi787 & n23866;
  assign n23994 = ~n23992 & ~n23993;
  assign n23995 = ~pi644 & ~n23994;
  assign n23996 = pi644 & n23990;
  assign n23997 = pi715 & ~n23995;
  assign n23998 = ~n23996 & n23997;
  assign n23999 = ~n19771 & n23850;
  assign n24000 = ~n15960 & n23896;
  assign n24001 = ~n23999 & ~n24000;
  assign n24002 = pi644 & ~n24001;
  assign n24003 = ~pi644 & n23850;
  assign n24004 = ~pi715 & ~n24003;
  assign n24005 = ~n24002 & n24004;
  assign n24006 = pi1160 & ~n24005;
  assign n24007 = ~n23998 & n24006;
  assign n24008 = ~pi644 & ~n24001;
  assign n24009 = pi644 & n23850;
  assign n24010 = pi715 & ~n24009;
  assign n24011 = ~n24008 & n24010;
  assign n24012 = pi644 & ~n23994;
  assign n24013 = ~pi644 & n23990;
  assign n24014 = ~pi715 & ~n24012;
  assign n24015 = ~n24013 & n24014;
  assign n24016 = ~pi1160 & ~n24011;
  assign n24017 = ~n24015 & n24016;
  assign n24018 = ~n24007 & ~n24017;
  assign n24019 = pi790 & ~n24018;
  assign n24020 = pi832 & ~n23991;
  assign n24021 = ~n24019 & n24020;
  assign n24022 = ~pi178 & po1038;
  assign n24023 = ~pi178 & ~n16219;
  assign n24024 = n15747 & ~n24023;
  assign n24025 = ~pi688 & n9829;
  assign n24026 = n24023 & ~n24025;
  assign n24027 = ~pi178 & ~n16228;
  assign n24028 = n16227 & ~n24027;
  assign n24029 = ~pi178 & ~n17276;
  assign n24030 = ~pi38 & ~pi178;
  assign n24031 = n19350 & ~n24030;
  assign n24032 = ~n24029 & ~n24031;
  assign n24033 = ~pi688 & ~n24028;
  assign n24034 = ~n24032 & n24033;
  assign n24035 = ~n24026 & ~n24034;
  assign n24036 = ~pi778 & n24035;
  assign n24037 = ~pi625 & n24023;
  assign n24038 = pi625 & ~n24035;
  assign n24039 = pi1153 & ~n24037;
  assign n24040 = ~n24038 & n24039;
  assign n24041 = pi625 & n24023;
  assign n24042 = ~pi625 & ~n24035;
  assign n24043 = ~pi1153 & ~n24041;
  assign n24044 = ~n24042 & n24043;
  assign n24045 = ~n24040 & ~n24044;
  assign n24046 = pi778 & ~n24045;
  assign n24047 = ~n24036 & ~n24046;
  assign n24048 = ~n15741 & n24047;
  assign n24049 = n15741 & n24023;
  assign n24050 = ~n24048 & ~n24049;
  assign n24051 = ~n15747 & n24050;
  assign n24052 = ~n24024 & ~n24051;
  assign n24053 = ~n15753 & n24052;
  assign n24054 = n15753 & n24023;
  assign n24055 = ~n24053 & ~n24054;
  assign n24056 = ~n15759 & ~n24055;
  assign n24057 = n15759 & n24023;
  assign n24058 = ~n24056 & ~n24057;
  assign n24059 = ~pi792 & n24058;
  assign n24060 = ~pi628 & n24023;
  assign n24061 = pi628 & ~n24058;
  assign n24062 = pi1156 & ~n24060;
  assign n24063 = ~n24061 & n24062;
  assign n24064 = pi628 & n24023;
  assign n24065 = ~pi628 & ~n24058;
  assign n24066 = ~pi1156 & ~n24064;
  assign n24067 = ~n24065 & n24066;
  assign n24068 = ~n24063 & ~n24067;
  assign n24069 = pi792 & ~n24068;
  assign n24070 = ~n24059 & ~n24069;
  assign n24071 = pi647 & n24070;
  assign n24072 = ~pi647 & n24023;
  assign n24073 = ~n24071 & ~n24072;
  assign n24074 = pi1157 & n24073;
  assign n24075 = ~pi647 & n24070;
  assign n24076 = pi647 & n24023;
  assign n24077 = ~pi1157 & ~n24076;
  assign n24078 = ~n24075 & n24077;
  assign n24079 = ~n24074 & ~n24078;
  assign n24080 = pi787 & ~n24079;
  assign n24081 = ~pi787 & ~n24070;
  assign n24082 = ~n24080 & ~n24081;
  assign n24083 = ~pi644 & n24082;
  assign n24084 = pi715 & ~n24083;
  assign n24085 = pi178 & ~n9829;
  assign n24086 = ~pi178 & n16514;
  assign n24087 = pi178 & ~n16565;
  assign n24088 = ~pi760 & ~n24086;
  assign n24089 = ~n24087 & n24088;
  assign n24090 = ~pi178 & pi760;
  assign n24091 = ~n16214 & n24090;
  assign n24092 = ~n24089 & ~n24091;
  assign n24093 = ~pi38 & ~n24092;
  assign n24094 = ~pi760 & n16570;
  assign n24095 = ~n24027 & ~n24094;
  assign n24096 = pi38 & ~n24095;
  assign n24097 = n9829 & ~n24096;
  assign n24098 = ~n24093 & n24097;
  assign n24099 = ~n24085 & ~n24098;
  assign n24100 = ~n15777 & ~n24099;
  assign n24101 = n15777 & ~n24023;
  assign n24102 = ~n24100 & ~n24101;
  assign n24103 = ~pi785 & ~n24102;
  assign n24104 = ~n15786 & ~n24023;
  assign n24105 = pi609 & n24100;
  assign n24106 = ~n24104 & ~n24105;
  assign n24107 = pi1155 & ~n24106;
  assign n24108 = ~n16585 & ~n24023;
  assign n24109 = ~pi609 & n24100;
  assign n24110 = ~n24108 & ~n24109;
  assign n24111 = ~pi1155 & ~n24110;
  assign n24112 = ~n24107 & ~n24111;
  assign n24113 = pi785 & ~n24112;
  assign n24114 = ~n24103 & ~n24113;
  assign n24115 = ~pi781 & ~n24114;
  assign n24116 = ~pi618 & n24023;
  assign n24117 = pi618 & n24114;
  assign n24118 = pi1154 & ~n24116;
  assign n24119 = ~n24117 & n24118;
  assign n24120 = ~pi618 & n24114;
  assign n24121 = pi618 & n24023;
  assign n24122 = ~pi1154 & ~n24121;
  assign n24123 = ~n24120 & n24122;
  assign n24124 = ~n24119 & ~n24123;
  assign n24125 = pi781 & ~n24124;
  assign n24126 = ~n24115 & ~n24125;
  assign n24127 = ~pi789 & ~n24126;
  assign n24128 = ~pi619 & n24023;
  assign n24129 = pi619 & n24126;
  assign n24130 = pi1159 & ~n24128;
  assign n24131 = ~n24129 & n24130;
  assign n24132 = ~pi619 & n24126;
  assign n24133 = pi619 & n24023;
  assign n24134 = ~pi1159 & ~n24133;
  assign n24135 = ~n24132 & n24134;
  assign n24136 = ~n24131 & ~n24135;
  assign n24137 = pi789 & ~n24136;
  assign n24138 = ~n24127 & ~n24137;
  assign n24139 = ~n15832 & n24138;
  assign n24140 = n15832 & n24023;
  assign n24141 = ~n24139 & ~n24140;
  assign n24142 = ~n15925 & ~n24141;
  assign n24143 = n15925 & n24023;
  assign n24144 = ~n24142 & ~n24143;
  assign n24145 = ~n15960 & ~n24144;
  assign n24146 = n15960 & n24023;
  assign n24147 = ~n24145 & ~n24146;
  assign n24148 = pi644 & ~n24147;
  assign n24149 = ~pi644 & n24023;
  assign n24150 = ~pi715 & ~n24149;
  assign n24151 = ~n24148 & n24150;
  assign n24152 = pi1160 & ~n24151;
  assign n24153 = ~n24084 & n24152;
  assign n24154 = pi644 & n24082;
  assign n24155 = ~pi715 & ~n24154;
  assign n24156 = ~pi644 & ~n24147;
  assign n24157 = pi644 & n24023;
  assign n24158 = pi715 & ~n24157;
  assign n24159 = ~n24156 & n24158;
  assign n24160 = ~pi1160 & ~n24159;
  assign n24161 = ~n24155 & n24160;
  assign n24162 = ~n24153 & ~n24161;
  assign n24163 = pi790 & ~n24162;
  assign n24164 = n15957 & n24073;
  assign n24165 = pi630 & n24078;
  assign n24166 = n19478 & n24144;
  assign n24167 = ~n24164 & ~n24165;
  assign n24168 = ~n24166 & n24167;
  assign n24169 = pi787 & ~n24168;
  assign n24170 = ~n16633 & n24141;
  assign n24171 = ~pi629 & n24063;
  assign n24172 = pi629 & n24067;
  assign n24173 = ~n24171 & ~n24172;
  assign n24174 = ~n24170 & n24173;
  assign n24175 = pi792 & ~n24174;
  assign n24176 = n15828 & ~n24055;
  assign n24177 = ~pi626 & ~n24023;
  assign n24178 = pi626 & ~n24138;
  assign n24179 = n15756 & ~n24177;
  assign n24180 = ~n24178 & n24179;
  assign n24181 = pi626 & ~n24023;
  assign n24182 = ~pi626 & ~n24138;
  assign n24183 = n15757 & ~n24181;
  assign n24184 = ~n24182 & n24183;
  assign n24185 = ~n24176 & ~n24180;
  assign n24186 = ~n24184 & n24185;
  assign n24187 = pi788 & ~n24186;
  assign n24188 = pi618 & ~n24050;
  assign n24189 = pi609 & n24047;
  assign n24190 = ~n24025 & ~n24098;
  assign n24191 = ~pi760 & ~n16808;
  assign n24192 = n18669 & ~n24191;
  assign n24193 = ~pi178 & ~n24192;
  assign n24194 = ~n16921 & ~n23872;
  assign n24195 = pi178 & ~n24194;
  assign n24196 = n6081 & n24195;
  assign n24197 = pi38 & ~n24196;
  assign n24198 = ~n24193 & n24197;
  assign n24199 = ~pi178 & ~n16647;
  assign n24200 = pi178 & ~n17397;
  assign n24201 = ~pi760 & ~n24199;
  assign n24202 = ~n24200 & n24201;
  assign n24203 = ~pi178 & n16653;
  assign n24204 = pi178 & n16657;
  assign n24205 = pi760 & ~n24203;
  assign n24206 = ~n24204 & n24205;
  assign n24207 = ~pi39 & ~n24202;
  assign n24208 = ~n24206 & n24207;
  assign n24209 = pi178 & n16825;
  assign n24210 = ~pi178 & ~n16747;
  assign n24211 = pi760 & ~n24209;
  assign n24212 = ~n24210 & n24211;
  assign n24213 = ~pi178 & n16877;
  assign n24214 = pi178 & n16913;
  assign n24215 = ~pi760 & ~n24213;
  assign n24216 = ~n24214 & n24215;
  assign n24217 = pi39 & ~n24216;
  assign n24218 = ~n24212 & n24217;
  assign n24219 = ~pi38 & ~n24208;
  assign n24220 = ~n24218 & n24219;
  assign n24221 = ~pi688 & ~n24198;
  assign n24222 = ~n24220 & n24221;
  assign n24223 = ~n24190 & ~n24222;
  assign n24224 = ~n24085 & ~n24223;
  assign n24225 = ~pi625 & n24224;
  assign n24226 = pi625 & n24099;
  assign n24227 = ~pi1153 & ~n24226;
  assign n24228 = ~n24225 & n24227;
  assign n24229 = ~pi608 & ~n24040;
  assign n24230 = ~n24228 & n24229;
  assign n24231 = ~pi625 & n24099;
  assign n24232 = pi625 & n24224;
  assign n24233 = pi1153 & ~n24231;
  assign n24234 = ~n24232 & n24233;
  assign n24235 = pi608 & ~n24044;
  assign n24236 = ~n24234 & n24235;
  assign n24237 = ~n24230 & ~n24236;
  assign n24238 = pi778 & ~n24237;
  assign n24239 = ~pi778 & n24224;
  assign n24240 = ~n24238 & ~n24239;
  assign n24241 = ~pi609 & ~n24240;
  assign n24242 = ~pi1155 & ~n24189;
  assign n24243 = ~n24241 & n24242;
  assign n24244 = ~pi660 & ~n24107;
  assign n24245 = ~n24243 & n24244;
  assign n24246 = ~pi609 & n24047;
  assign n24247 = pi609 & ~n24240;
  assign n24248 = pi1155 & ~n24246;
  assign n24249 = ~n24247 & n24248;
  assign n24250 = pi660 & ~n24111;
  assign n24251 = ~n24249 & n24250;
  assign n24252 = ~n24245 & ~n24251;
  assign n24253 = pi785 & ~n24252;
  assign n24254 = ~pi785 & ~n24240;
  assign n24255 = ~n24253 & ~n24254;
  assign n24256 = ~pi618 & ~n24255;
  assign n24257 = ~pi1154 & ~n24188;
  assign n24258 = ~n24256 & n24257;
  assign n24259 = ~pi627 & ~n24119;
  assign n24260 = ~n24258 & n24259;
  assign n24261 = ~pi618 & ~n24050;
  assign n24262 = pi618 & ~n24255;
  assign n24263 = pi1154 & ~n24261;
  assign n24264 = ~n24262 & n24263;
  assign n24265 = pi627 & ~n24123;
  assign n24266 = ~n24264 & n24265;
  assign n24267 = ~n24260 & ~n24266;
  assign n24268 = pi781 & ~n24267;
  assign n24269 = ~pi781 & ~n24255;
  assign n24270 = ~n24268 & ~n24269;
  assign n24271 = ~pi789 & n24270;
  assign n24272 = ~pi619 & n24052;
  assign n24273 = pi619 & ~n24270;
  assign n24274 = pi1159 & ~n24272;
  assign n24275 = ~n24273 & n24274;
  assign n24276 = pi648 & ~n24135;
  assign n24277 = ~n24275 & n24276;
  assign n24278 = ~pi619 & ~n24270;
  assign n24279 = pi619 & n24052;
  assign n24280 = ~pi1159 & ~n24279;
  assign n24281 = ~n24278 & n24280;
  assign n24282 = ~pi648 & ~n24131;
  assign n24283 = ~n24281 & n24282;
  assign n24284 = pi789 & ~n24277;
  assign n24285 = ~n24283 & n24284;
  assign n24286 = n15833 & ~n24271;
  assign n24287 = ~n24285 & n24286;
  assign n24288 = ~n16644 & ~n24187;
  assign n24289 = ~n24287 & n24288;
  assign n24290 = ~n24175 & ~n24289;
  assign n24291 = n18841 & ~n24290;
  assign n24292 = pi644 & ~n24151;
  assign n24293 = ~n24160 & ~n24292;
  assign n24294 = ~n22949 & ~n24293;
  assign n24295 = pi790 & ~n24294;
  assign n24296 = ~n24169 & ~n24291;
  assign n24297 = ~n24295 & n24296;
  assign n24298 = ~n24163 & ~n24297;
  assign n24299 = ~po1038 & ~n24298;
  assign n24300 = ~pi832 & ~n24022;
  assign n24301 = ~n24299 & n24300;
  assign po335 = ~n24021 & ~n24301;
  assign n24303 = ~pi179 & ~n2923;
  assign n24304 = ~pi724 & n15726;
  assign n24305 = ~n24303 & ~n24304;
  assign n24306 = ~pi778 & n24305;
  assign n24307 = ~pi625 & n24304;
  assign n24308 = ~n24305 & ~n24307;
  assign n24309 = pi1153 & ~n24308;
  assign n24310 = ~pi1153 & ~n24303;
  assign n24311 = ~n24307 & n24310;
  assign n24312 = ~n24309 & ~n24311;
  assign n24313 = pi778 & ~n24312;
  assign n24314 = ~n24306 & ~n24313;
  assign n24315 = ~n15742 & n24314;
  assign n24316 = ~n15748 & n24315;
  assign n24317 = ~n15754 & n24316;
  assign n24318 = ~n15760 & n24317;
  assign n24319 = ~n15766 & n24318;
  assign n24320 = n19394 & n24319;
  assign n24321 = ~n19394 & n24303;
  assign n24322 = ~n24320 & ~n24321;
  assign n24323 = ~n15959 & n24322;
  assign n24324 = n15925 & n24303;
  assign n24325 = ~pi741 & n15781;
  assign n24326 = ~n24303 & ~n24325;
  assign n24327 = ~n15778 & ~n24326;
  assign n24328 = ~pi785 & ~n24327;
  assign n24329 = ~n15787 & ~n24326;
  assign n24330 = pi1155 & ~n24329;
  assign n24331 = ~n15790 & n24327;
  assign n24332 = ~pi1155 & ~n24331;
  assign n24333 = ~n24330 & ~n24332;
  assign n24334 = pi785 & ~n24333;
  assign n24335 = ~n24328 & ~n24334;
  assign n24336 = ~pi781 & ~n24335;
  assign n24337 = ~n15797 & n24335;
  assign n24338 = pi1154 & ~n24337;
  assign n24339 = ~n15800 & n24335;
  assign n24340 = ~pi1154 & ~n24339;
  assign n24341 = ~n24338 & ~n24340;
  assign n24342 = pi781 & ~n24341;
  assign n24343 = ~n24336 & ~n24342;
  assign n24344 = ~pi789 & ~n24343;
  assign n24345 = ~pi619 & n24303;
  assign n24346 = pi619 & n24343;
  assign n24347 = pi1159 & ~n24345;
  assign n24348 = ~n24346 & n24347;
  assign n24349 = ~pi619 & n24343;
  assign n24350 = pi619 & n24303;
  assign n24351 = ~pi1159 & ~n24350;
  assign n24352 = ~n24349 & n24351;
  assign n24353 = ~n24348 & ~n24352;
  assign n24354 = pi789 & ~n24353;
  assign n24355 = ~n24344 & ~n24354;
  assign n24356 = ~n15832 & ~n24355;
  assign n24357 = n15832 & ~n24303;
  assign n24358 = ~n24356 & ~n24357;
  assign n24359 = ~n15925 & n24358;
  assign n24360 = n19478 & ~n24324;
  assign n24361 = ~n24359 & n24360;
  assign n24362 = ~n24323 & ~n24361;
  assign n24363 = pi787 & ~n24362;
  assign n24364 = n15828 & n24317;
  assign n24365 = ~pi626 & ~n24303;
  assign n24366 = pi626 & ~n24355;
  assign n24367 = n15756 & ~n24365;
  assign n24368 = ~n24366 & n24367;
  assign n24369 = pi626 & ~n24303;
  assign n24370 = ~pi626 & ~n24355;
  assign n24371 = n15757 & ~n24369;
  assign n24372 = ~n24370 & n24371;
  assign n24373 = ~n24364 & ~n24368;
  assign n24374 = ~n24372 & n24373;
  assign n24375 = pi788 & ~n24374;
  assign n24376 = pi618 & n24315;
  assign n24377 = pi609 & n24314;
  assign n24378 = ~n15780 & ~n24305;
  assign n24379 = pi625 & n24378;
  assign n24380 = n24326 & ~n24378;
  assign n24381 = ~n24379 & ~n24380;
  assign n24382 = n24310 & ~n24381;
  assign n24383 = ~pi608 & ~n24309;
  assign n24384 = ~n24382 & n24383;
  assign n24385 = pi1153 & n24326;
  assign n24386 = ~n24379 & n24385;
  assign n24387 = pi608 & ~n24311;
  assign n24388 = ~n24386 & n24387;
  assign n24389 = ~n24384 & ~n24388;
  assign n24390 = pi778 & ~n24389;
  assign n24391 = ~pi778 & ~n24380;
  assign n24392 = ~n24390 & ~n24391;
  assign n24393 = ~pi609 & ~n24392;
  assign n24394 = ~pi1155 & ~n24377;
  assign n24395 = ~n24393 & n24394;
  assign n24396 = ~pi660 & ~n24330;
  assign n24397 = ~n24395 & n24396;
  assign n24398 = ~pi609 & n24314;
  assign n24399 = pi609 & ~n24392;
  assign n24400 = pi1155 & ~n24398;
  assign n24401 = ~n24399 & n24400;
  assign n24402 = pi660 & ~n24332;
  assign n24403 = ~n24401 & n24402;
  assign n24404 = ~n24397 & ~n24403;
  assign n24405 = pi785 & ~n24404;
  assign n24406 = ~pi785 & ~n24392;
  assign n24407 = ~n24405 & ~n24406;
  assign n24408 = ~pi618 & ~n24407;
  assign n24409 = ~pi1154 & ~n24376;
  assign n24410 = ~n24408 & n24409;
  assign n24411 = ~pi627 & ~n24338;
  assign n24412 = ~n24410 & n24411;
  assign n24413 = ~pi618 & n24315;
  assign n24414 = pi618 & ~n24407;
  assign n24415 = pi1154 & ~n24413;
  assign n24416 = ~n24414 & n24415;
  assign n24417 = pi627 & ~n24340;
  assign n24418 = ~n24416 & n24417;
  assign n24419 = ~n24412 & ~n24418;
  assign n24420 = pi781 & ~n24419;
  assign n24421 = ~pi781 & ~n24407;
  assign n24422 = ~n24420 & ~n24421;
  assign n24423 = ~pi789 & n24422;
  assign n24424 = ~pi619 & n24316;
  assign n24425 = pi619 & ~n24422;
  assign n24426 = pi1159 & ~n24424;
  assign n24427 = ~n24425 & n24426;
  assign n24428 = pi648 & ~n24352;
  assign n24429 = ~n24427 & n24428;
  assign n24430 = pi619 & n24316;
  assign n24431 = ~pi619 & ~n24422;
  assign n24432 = ~pi1159 & ~n24430;
  assign n24433 = ~n24431 & n24432;
  assign n24434 = ~pi648 & ~n24348;
  assign n24435 = ~n24433 & n24434;
  assign n24436 = pi789 & ~n24429;
  assign n24437 = ~n24435 & n24436;
  assign n24438 = n15833 & ~n24423;
  assign n24439 = ~n24437 & n24438;
  assign n24440 = ~n24375 & ~n24439;
  assign n24441 = ~n16644 & ~n24440;
  assign n24442 = n15763 & n24358;
  assign n24443 = n15772 & n24318;
  assign n24444 = ~pi629 & ~n24443;
  assign n24445 = ~n24442 & n24444;
  assign n24446 = n15762 & n24358;
  assign n24447 = n15909 & n24318;
  assign n24448 = pi629 & ~n24447;
  assign n24449 = ~n24446 & n24448;
  assign n24450 = pi792 & ~n24445;
  assign n24451 = ~n24449 & n24450;
  assign n24452 = n18841 & ~n24451;
  assign n24453 = ~n24441 & n24452;
  assign n24454 = ~n24363 & ~n24453;
  assign n24455 = ~pi790 & n24454;
  assign n24456 = pi787 & ~n24322;
  assign n24457 = ~pi787 & n24319;
  assign n24458 = ~n24456 & ~n24457;
  assign n24459 = ~pi644 & ~n24458;
  assign n24460 = pi644 & n24454;
  assign n24461 = pi715 & ~n24459;
  assign n24462 = ~n24460 & n24461;
  assign n24463 = ~n19771 & n24303;
  assign n24464 = ~n15960 & n24359;
  assign n24465 = ~n24463 & ~n24464;
  assign n24466 = pi644 & ~n24465;
  assign n24467 = ~pi644 & n24303;
  assign n24468 = ~pi715 & ~n24467;
  assign n24469 = ~n24466 & n24468;
  assign n24470 = pi1160 & ~n24469;
  assign n24471 = ~n24462 & n24470;
  assign n24472 = ~pi644 & ~n24465;
  assign n24473 = pi644 & n24303;
  assign n24474 = pi715 & ~n24473;
  assign n24475 = ~n24472 & n24474;
  assign n24476 = pi644 & ~n24458;
  assign n24477 = ~pi644 & n24454;
  assign n24478 = ~pi715 & ~n24476;
  assign n24479 = ~n24477 & n24478;
  assign n24480 = ~pi1160 & ~n24475;
  assign n24481 = ~n24479 & n24480;
  assign n24482 = ~n24471 & ~n24481;
  assign n24483 = pi790 & ~n24482;
  assign n24484 = pi832 & ~n24455;
  assign n24485 = ~n24483 & n24484;
  assign n24486 = ~pi179 & po1038;
  assign n24487 = ~pi179 & ~n16219;
  assign n24488 = n15759 & ~n24487;
  assign n24489 = n15747 & ~n24487;
  assign n24490 = ~pi724 & n9829;
  assign n24491 = n24487 & ~n24490;
  assign n24492 = ~pi179 & ~n16228;
  assign n24493 = n16227 & ~n24492;
  assign n24494 = ~pi179 & ~n17276;
  assign n24495 = ~pi38 & ~pi179;
  assign n24496 = n19350 & ~n24495;
  assign n24497 = ~n24494 & ~n24496;
  assign n24498 = ~pi724 & ~n24493;
  assign n24499 = ~n24497 & n24498;
  assign n24500 = ~n24491 & ~n24499;
  assign n24501 = ~pi778 & n24500;
  assign n24502 = ~pi625 & n24487;
  assign n24503 = pi625 & ~n24500;
  assign n24504 = pi1153 & ~n24502;
  assign n24505 = ~n24503 & n24504;
  assign n24506 = pi625 & n24487;
  assign n24507 = ~pi625 & ~n24500;
  assign n24508 = ~pi1153 & ~n24506;
  assign n24509 = ~n24507 & n24508;
  assign n24510 = ~n24505 & ~n24509;
  assign n24511 = pi778 & ~n24510;
  assign n24512 = ~n24501 & ~n24511;
  assign n24513 = ~n15741 & n24512;
  assign n24514 = n15741 & n24487;
  assign n24515 = ~n24513 & ~n24514;
  assign n24516 = ~n15747 & n24515;
  assign n24517 = ~n24489 & ~n24516;
  assign n24518 = ~n15753 & n24517;
  assign n24519 = n15753 & n24487;
  assign n24520 = ~n24518 & ~n24519;
  assign n24521 = ~n15759 & n24520;
  assign n24522 = ~n24488 & ~n24521;
  assign n24523 = ~pi792 & ~n24522;
  assign n24524 = ~pi628 & ~n24487;
  assign n24525 = pi628 & ~n24522;
  assign n24526 = ~n24524 & ~n24525;
  assign n24527 = pi1156 & ~n24526;
  assign n24528 = ~pi628 & n24522;
  assign n24529 = pi628 & n24487;
  assign n24530 = ~pi1156 & ~n24529;
  assign n24531 = ~n24528 & n24530;
  assign n24532 = ~n24527 & ~n24531;
  assign n24533 = pi792 & ~n24532;
  assign n24534 = ~n24523 & ~n24533;
  assign n24535 = ~pi787 & ~n24534;
  assign n24536 = ~pi647 & n24487;
  assign n24537 = pi647 & n24534;
  assign n24538 = pi1157 & ~n24536;
  assign n24539 = ~n24537 & n24538;
  assign n24540 = ~pi647 & n24534;
  assign n24541 = pi647 & n24487;
  assign n24542 = ~pi1157 & ~n24541;
  assign n24543 = ~n24540 & n24542;
  assign n24544 = ~n24539 & ~n24543;
  assign n24545 = pi787 & ~n24544;
  assign n24546 = ~n24535 & ~n24545;
  assign n24547 = ~pi644 & n24546;
  assign n24548 = ~pi629 & n24527;
  assign n24549 = pi619 & n24517;
  assign n24550 = ~pi1159 & ~n24549;
  assign n24551 = ~pi619 & n24487;
  assign n24552 = pi179 & ~n9829;
  assign n24553 = ~pi741 & ~n23191;
  assign n24554 = pi179 & ~n24553;
  assign n24555 = ~n18598 & n18604;
  assign n24556 = ~pi179 & ~pi741;
  assign n24557 = n24555 & n24556;
  assign n24558 = ~n24554 & ~n24557;
  assign n24559 = ~n20547 & n24558;
  assign n24560 = n9829 & ~n24559;
  assign n24561 = ~n24552 & ~n24560;
  assign n24562 = ~n15777 & ~n24561;
  assign n24563 = n15777 & ~n24487;
  assign n24564 = ~n24562 & ~n24563;
  assign n24565 = ~pi785 & ~n24564;
  assign n24566 = ~n15786 & ~n24487;
  assign n24567 = pi609 & n24562;
  assign n24568 = ~n24566 & ~n24567;
  assign n24569 = pi1155 & ~n24568;
  assign n24570 = ~n16585 & ~n24487;
  assign n24571 = ~pi609 & n24562;
  assign n24572 = ~n24570 & ~n24571;
  assign n24573 = ~pi1155 & ~n24572;
  assign n24574 = ~n24569 & ~n24573;
  assign n24575 = pi785 & ~n24574;
  assign n24576 = ~n24565 & ~n24575;
  assign n24577 = ~pi781 & ~n24576;
  assign n24578 = ~pi618 & n24487;
  assign n24579 = pi618 & n24576;
  assign n24580 = pi1154 & ~n24578;
  assign n24581 = ~n24579 & n24580;
  assign n24582 = ~pi618 & n24576;
  assign n24583 = pi618 & n24487;
  assign n24584 = ~pi1154 & ~n24583;
  assign n24585 = ~n24582 & n24584;
  assign n24586 = ~n24581 & ~n24585;
  assign n24587 = pi781 & ~n24586;
  assign n24588 = ~n24577 & ~n24587;
  assign n24589 = pi619 & n24588;
  assign n24590 = pi1159 & ~n24551;
  assign n24591 = ~n24589 & n24590;
  assign n24592 = ~pi648 & ~n24591;
  assign n24593 = ~n24550 & n24592;
  assign n24594 = ~pi619 & n24517;
  assign n24595 = pi1159 & ~n24594;
  assign n24596 = ~pi619 & n24588;
  assign n24597 = pi619 & n24487;
  assign n24598 = ~pi1159 & ~n24597;
  assign n24599 = ~n24596 & n24598;
  assign n24600 = pi648 & ~n24599;
  assign n24601 = ~n24595 & n24600;
  assign n24602 = ~n24593 & ~n24601;
  assign n24603 = pi789 & ~n24602;
  assign n24604 = pi619 & n24600;
  assign n24605 = ~pi619 & n24592;
  assign n24606 = pi789 & ~n24604;
  assign n24607 = ~n24605 & n24606;
  assign n24608 = pi609 & n24512;
  assign n24609 = ~n24490 & ~n24560;
  assign n24610 = ~pi179 & ~n18651;
  assign n24611 = pi179 & n18659;
  assign n24612 = ~pi741 & ~n24610;
  assign n24613 = ~n24611 & n24612;
  assign n24614 = n17390 & ~n24492;
  assign n24615 = pi179 & n18665;
  assign n24616 = ~pi179 & ~n18673;
  assign n24617 = ~pi38 & ~n24615;
  assign n24618 = ~n24616 & n24617;
  assign n24619 = ~n24614 & ~n24618;
  assign n24620 = pi741 & ~n24619;
  assign n24621 = ~pi724 & ~n24613;
  assign n24622 = ~n24620 & n24621;
  assign n24623 = ~n24609 & ~n24622;
  assign n24624 = ~n24552 & ~n24623;
  assign n24625 = ~pi625 & n24624;
  assign n24626 = pi625 & n24561;
  assign n24627 = ~pi1153 & ~n24626;
  assign n24628 = ~n24625 & n24627;
  assign n24629 = ~pi608 & ~n24505;
  assign n24630 = ~n24628 & n24629;
  assign n24631 = ~pi625 & n24561;
  assign n24632 = pi625 & n24624;
  assign n24633 = pi1153 & ~n24631;
  assign n24634 = ~n24632 & n24633;
  assign n24635 = pi608 & ~n24509;
  assign n24636 = ~n24634 & n24635;
  assign n24637 = ~n24630 & ~n24636;
  assign n24638 = pi778 & ~n24637;
  assign n24639 = ~pi778 & n24624;
  assign n24640 = ~n24638 & ~n24639;
  assign n24641 = ~pi609 & ~n24640;
  assign n24642 = ~pi1155 & ~n24608;
  assign n24643 = ~n24641 & n24642;
  assign n24644 = ~pi660 & ~n24569;
  assign n24645 = ~n24643 & n24644;
  assign n24646 = ~pi609 & n24512;
  assign n24647 = pi609 & ~n24640;
  assign n24648 = pi1155 & ~n24646;
  assign n24649 = ~n24647 & n24648;
  assign n24650 = pi660 & ~n24573;
  assign n24651 = ~n24649 & n24650;
  assign n24652 = ~n24645 & ~n24651;
  assign n24653 = pi785 & ~n24652;
  assign n24654 = ~pi785 & ~n24640;
  assign n24655 = ~n24653 & ~n24654;
  assign n24656 = ~pi781 & n24655;
  assign n24657 = pi618 & ~n24515;
  assign n24658 = ~pi618 & ~n24655;
  assign n24659 = ~pi1154 & ~n24657;
  assign n24660 = ~n24658 & n24659;
  assign n24661 = ~pi627 & ~n24581;
  assign n24662 = ~n24660 & n24661;
  assign n24663 = ~pi618 & ~n24515;
  assign n24664 = pi618 & ~n24655;
  assign n24665 = pi1154 & ~n24663;
  assign n24666 = ~n24664 & n24665;
  assign n24667 = pi627 & ~n24585;
  assign n24668 = ~n24666 & n24667;
  assign n24669 = pi781 & ~n24662;
  assign n24670 = ~n24668 & n24669;
  assign n24671 = ~n24607 & ~n24656;
  assign n24672 = ~n24670 & n24671;
  assign n24673 = ~n24603 & ~n24672;
  assign n24674 = n15833 & ~n24673;
  assign n24675 = pi641 & ~n24487;
  assign n24676 = ~pi641 & n24520;
  assign n24677 = n15819 & ~n24675;
  assign n24678 = ~n24676 & n24677;
  assign n24679 = ~pi789 & ~n24588;
  assign n24680 = ~n24591 & ~n24599;
  assign n24681 = pi789 & ~n24680;
  assign n24682 = ~n24679 & ~n24681;
  assign n24683 = n22348 & n24682;
  assign n24684 = ~pi641 & ~n24487;
  assign n24685 = pi641 & n24520;
  assign n24686 = n15818 & ~n24684;
  assign n24687 = ~n24685 & n24686;
  assign n24688 = ~n24678 & ~n24687;
  assign n24689 = ~n24683 & n24688;
  assign n24690 = pi788 & ~n24689;
  assign n24691 = ~n24674 & ~n24690;
  assign n24692 = ~n16643 & n24691;
  assign n24693 = ~n15832 & n24682;
  assign n24694 = n15832 & n24487;
  assign n24695 = ~n24693 & ~n24694;
  assign n24696 = ~n16633 & n24695;
  assign n24697 = pi629 & n24531;
  assign n24698 = ~n24548 & ~n24697;
  assign n24699 = ~n24696 & n24698;
  assign n24700 = ~n24692 & n24699;
  assign n24701 = pi792 & ~n24700;
  assign n24702 = ~pi792 & n24691;
  assign n24703 = ~n24701 & ~n24702;
  assign n24704 = ~pi647 & n24703;
  assign n24705 = ~n15925 & ~n24695;
  assign n24706 = n15925 & n24487;
  assign n24707 = ~n24705 & ~n24706;
  assign n24708 = pi647 & ~n24707;
  assign n24709 = ~pi1157 & ~n24708;
  assign n24710 = ~n24704 & n24709;
  assign n24711 = ~pi630 & ~n24539;
  assign n24712 = ~n24710 & n24711;
  assign n24713 = ~pi647 & ~n24707;
  assign n24714 = pi647 & n24703;
  assign n24715 = pi1157 & ~n24713;
  assign n24716 = ~n24714 & n24715;
  assign n24717 = pi630 & ~n24543;
  assign n24718 = ~n24716 & n24717;
  assign n24719 = ~n24712 & ~n24718;
  assign n24720 = pi787 & ~n24719;
  assign n24721 = ~pi787 & n24703;
  assign n24722 = ~n24720 & ~n24721;
  assign n24723 = pi644 & ~n24722;
  assign n24724 = pi715 & ~n24547;
  assign n24725 = ~n24723 & n24724;
  assign n24726 = ~n15960 & ~n24707;
  assign n24727 = n15960 & n24487;
  assign n24728 = ~n24726 & ~n24727;
  assign n24729 = pi644 & ~n24728;
  assign n24730 = ~pi644 & n24487;
  assign n24731 = ~pi715 & ~n24730;
  assign n24732 = ~n24729 & n24731;
  assign n24733 = pi1160 & ~n24732;
  assign n24734 = ~n24725 & n24733;
  assign n24735 = pi644 & n24546;
  assign n24736 = ~pi715 & ~n24735;
  assign n24737 = ~pi644 & ~n24728;
  assign n24738 = pi644 & n24487;
  assign n24739 = pi715 & ~n24738;
  assign n24740 = ~n24737 & n24739;
  assign n24741 = ~pi1160 & ~n24740;
  assign n24742 = ~n24736 & n24741;
  assign n24743 = ~n24734 & ~n24742;
  assign n24744 = pi790 & ~n24743;
  assign n24745 = ~pi644 & n24741;
  assign n24746 = pi790 & ~n24745;
  assign n24747 = ~n24722 & ~n24746;
  assign n24748 = ~n24744 & ~n24747;
  assign n24749 = ~po1038 & ~n24748;
  assign n24750 = ~pi832 & ~n24486;
  assign n24751 = ~n24749 & n24750;
  assign po336 = ~n24485 & ~n24751;
  assign n24753 = ~pi180 & ~n2923;
  assign n24754 = ~pi702 & n15726;
  assign n24755 = ~n24753 & ~n24754;
  assign n24756 = ~pi778 & ~n24755;
  assign n24757 = ~pi625 & n24754;
  assign n24758 = ~n24755 & ~n24757;
  assign n24759 = pi1153 & ~n24758;
  assign n24760 = ~pi1153 & ~n24753;
  assign n24761 = ~n24757 & n24760;
  assign n24762 = pi778 & ~n24761;
  assign n24763 = ~n24759 & n24762;
  assign n24764 = ~n24756 & ~n24763;
  assign n24765 = ~n15742 & ~n24764;
  assign n24766 = ~n15748 & n24765;
  assign n24767 = ~n15754 & n24766;
  assign n24768 = ~n15760 & n24767;
  assign n24769 = ~n15766 & n24768;
  assign n24770 = n19394 & n24769;
  assign n24771 = ~n19394 & n24753;
  assign n24772 = ~n24770 & ~n24771;
  assign n24773 = ~n15959 & n24772;
  assign n24774 = n15925 & n24753;
  assign n24775 = ~pi753 & n15781;
  assign n24776 = ~n24753 & ~n24775;
  assign n24777 = ~n15778 & ~n24776;
  assign n24778 = ~pi785 & ~n24777;
  assign n24779 = n16585 & n24775;
  assign n24780 = n24777 & ~n24779;
  assign n24781 = pi1155 & ~n24780;
  assign n24782 = ~pi1155 & ~n24753;
  assign n24783 = ~n24779 & n24782;
  assign n24784 = ~n24781 & ~n24783;
  assign n24785 = pi785 & ~n24784;
  assign n24786 = ~n24778 & ~n24785;
  assign n24787 = ~pi781 & ~n24786;
  assign n24788 = ~n15797 & n24786;
  assign n24789 = pi1154 & ~n24788;
  assign n24790 = ~n15800 & n24786;
  assign n24791 = ~pi1154 & ~n24790;
  assign n24792 = ~n24789 & ~n24791;
  assign n24793 = pi781 & ~n24792;
  assign n24794 = ~n24787 & ~n24793;
  assign n24795 = ~n21915 & n24794;
  assign n24796 = ~n15832 & ~n24795;
  assign n24797 = n15832 & ~n24753;
  assign n24798 = ~n24796 & ~n24797;
  assign n24799 = ~n15925 & n24798;
  assign n24800 = n19478 & ~n24774;
  assign n24801 = ~n24799 & n24800;
  assign n24802 = ~n24773 & ~n24801;
  assign n24803 = pi787 & ~n24802;
  assign n24804 = n15763 & n24798;
  assign n24805 = n15772 & n24768;
  assign n24806 = ~pi629 & ~n24805;
  assign n24807 = ~n24804 & n24806;
  assign n24808 = n15762 & n24798;
  assign n24809 = n15909 & n24768;
  assign n24810 = pi629 & ~n24809;
  assign n24811 = ~n24808 & n24810;
  assign n24812 = pi792 & ~n24807;
  assign n24813 = ~n24811 & n24812;
  assign n24814 = ~n21932 & n24794;
  assign n24815 = pi648 & ~n24814;
  assign n24816 = n21935 & ~n24766;
  assign n24817 = ~n24815 & ~n24816;
  assign n24818 = ~pi1159 & ~n24817;
  assign n24819 = ~pi619 & ~n24766;
  assign n24820 = pi648 & ~n24819;
  assign n24821 = n21942 & n24794;
  assign n24822 = pi1159 & ~n24820;
  assign n24823 = ~n24821 & n24822;
  assign n24824 = ~n24818 & ~n24823;
  assign n24825 = pi789 & ~n24824;
  assign n24826 = pi609 & ~n24764;
  assign n24827 = ~n15780 & ~n24755;
  assign n24828 = pi625 & n24827;
  assign n24829 = n24776 & ~n24827;
  assign n24830 = ~n24828 & ~n24829;
  assign n24831 = n24760 & ~n24830;
  assign n24832 = ~pi608 & ~n24759;
  assign n24833 = ~n24831 & n24832;
  assign n24834 = pi1153 & n24776;
  assign n24835 = ~n24828 & n24834;
  assign n24836 = pi608 & ~n24761;
  assign n24837 = ~n24835 & n24836;
  assign n24838 = ~n24833 & ~n24837;
  assign n24839 = pi778 & ~n24838;
  assign n24840 = ~pi778 & ~n24829;
  assign n24841 = ~n24839 & ~n24840;
  assign n24842 = ~pi609 & ~n24841;
  assign n24843 = ~pi1155 & ~n24826;
  assign n24844 = ~n24842 & n24843;
  assign n24845 = ~pi660 & ~n24781;
  assign n24846 = ~n24844 & n24845;
  assign n24847 = ~pi609 & ~n24764;
  assign n24848 = pi609 & ~n24841;
  assign n24849 = pi1155 & ~n24847;
  assign n24850 = ~n24848 & n24849;
  assign n24851 = pi660 & ~n24783;
  assign n24852 = ~n24850 & n24851;
  assign n24853 = ~n24846 & ~n24852;
  assign n24854 = pi785 & ~n24853;
  assign n24855 = ~pi785 & ~n24841;
  assign n24856 = ~n24854 & ~n24855;
  assign n24857 = ~pi781 & n24856;
  assign n24858 = pi618 & n24765;
  assign n24859 = ~pi618 & ~n24856;
  assign n24860 = ~pi1154 & ~n24858;
  assign n24861 = ~n24859 & n24860;
  assign n24862 = ~pi627 & ~n24789;
  assign n24863 = ~n24861 & n24862;
  assign n24864 = ~pi618 & n24765;
  assign n24865 = pi618 & ~n24856;
  assign n24866 = pi1154 & ~n24864;
  assign n24867 = ~n24865 & n24866;
  assign n24868 = pi627 & ~n24791;
  assign n24869 = ~n24867 & n24868;
  assign n24870 = pi781 & ~n24863;
  assign n24871 = ~n24869 & n24870;
  assign n24872 = ~n24825 & ~n24857;
  assign n24873 = ~n24871 & n24872;
  assign n24874 = n18969 & n24824;
  assign n24875 = ~n24873 & ~n24874;
  assign n24876 = n15833 & ~n24875;
  assign n24877 = n15828 & n24767;
  assign n24878 = ~pi626 & ~n24753;
  assign n24879 = pi626 & ~n24795;
  assign n24880 = n15756 & ~n24878;
  assign n24881 = ~n24879 & n24880;
  assign n24882 = pi626 & ~n24753;
  assign n24883 = ~pi626 & ~n24795;
  assign n24884 = n15757 & ~n24882;
  assign n24885 = ~n24883 & n24884;
  assign n24886 = ~n24877 & ~n24881;
  assign n24887 = ~n24885 & n24886;
  assign n24888 = pi788 & ~n24887;
  assign n24889 = ~n24876 & ~n24888;
  assign n24890 = ~n16644 & ~n24889;
  assign n24891 = n18841 & ~n24813;
  assign n24892 = ~n24890 & n24891;
  assign n24893 = ~n24803 & ~n24892;
  assign n24894 = ~pi790 & n24893;
  assign n24895 = pi787 & ~n24772;
  assign n24896 = ~pi787 & n24769;
  assign n24897 = ~n24895 & ~n24896;
  assign n24898 = ~pi644 & ~n24897;
  assign n24899 = pi644 & n24893;
  assign n24900 = pi715 & ~n24898;
  assign n24901 = ~n24899 & n24900;
  assign n24902 = ~n19771 & n24753;
  assign n24903 = ~n15960 & n24799;
  assign n24904 = ~n24902 & ~n24903;
  assign n24905 = pi644 & ~n24904;
  assign n24906 = ~pi644 & n24753;
  assign n24907 = ~pi715 & ~n24906;
  assign n24908 = ~n24905 & n24907;
  assign n24909 = pi1160 & ~n24908;
  assign n24910 = ~n24901 & n24909;
  assign n24911 = ~pi644 & ~n24904;
  assign n24912 = pi644 & n24753;
  assign n24913 = pi715 & ~n24912;
  assign n24914 = ~n24911 & n24913;
  assign n24915 = pi644 & ~n24897;
  assign n24916 = ~pi644 & n24893;
  assign n24917 = ~pi715 & ~n24915;
  assign n24918 = ~n24916 & n24917;
  assign n24919 = ~pi1160 & ~n24914;
  assign n24920 = ~n24918 & n24919;
  assign n24921 = ~n24910 & ~n24920;
  assign n24922 = pi790 & ~n24921;
  assign n24923 = pi832 & ~n24894;
  assign n24924 = ~n24922 & n24923;
  assign n24925 = ~pi180 & po1038;
  assign n24926 = ~pi180 & ~n16219;
  assign n24927 = n15747 & ~n24926;
  assign n24928 = ~pi702 & n9829;
  assign n24929 = n24926 & ~n24928;
  assign n24930 = ~pi180 & ~n16228;
  assign n24931 = n16227 & ~n24930;
  assign n24932 = ~pi180 & ~n17276;
  assign n24933 = ~pi38 & ~pi180;
  assign n24934 = n19350 & ~n24933;
  assign n24935 = ~n24932 & ~n24934;
  assign n24936 = ~pi702 & ~n24931;
  assign n24937 = ~n24935 & n24936;
  assign n24938 = ~n24929 & ~n24937;
  assign n24939 = ~pi778 & n24938;
  assign n24940 = ~pi625 & n24926;
  assign n24941 = pi625 & ~n24938;
  assign n24942 = pi1153 & ~n24940;
  assign n24943 = ~n24941 & n24942;
  assign n24944 = pi625 & n24926;
  assign n24945 = ~pi625 & ~n24938;
  assign n24946 = ~pi1153 & ~n24944;
  assign n24947 = ~n24945 & n24946;
  assign n24948 = ~n24943 & ~n24947;
  assign n24949 = pi778 & ~n24948;
  assign n24950 = ~n24939 & ~n24949;
  assign n24951 = ~n15741 & n24950;
  assign n24952 = n15741 & n24926;
  assign n24953 = ~n24951 & ~n24952;
  assign n24954 = ~n15747 & n24953;
  assign n24955 = ~n24927 & ~n24954;
  assign n24956 = ~n15753 & n24955;
  assign n24957 = n15753 & n24926;
  assign n24958 = ~n24956 & ~n24957;
  assign n24959 = ~n15759 & ~n24958;
  assign n24960 = n15759 & n24926;
  assign n24961 = ~n24959 & ~n24960;
  assign n24962 = ~pi792 & n24961;
  assign n24963 = ~pi628 & n24926;
  assign n24964 = pi628 & ~n24961;
  assign n24965 = pi1156 & ~n24963;
  assign n24966 = ~n24964 & n24965;
  assign n24967 = pi628 & n24926;
  assign n24968 = ~pi628 & ~n24961;
  assign n24969 = ~pi1156 & ~n24967;
  assign n24970 = ~n24968 & n24969;
  assign n24971 = ~n24966 & ~n24970;
  assign n24972 = pi792 & ~n24971;
  assign n24973 = ~n24962 & ~n24972;
  assign n24974 = n19394 & n24973;
  assign n24975 = ~n19394 & n24926;
  assign n24976 = ~n24974 & ~n24975;
  assign n24977 = pi787 & ~n24976;
  assign n24978 = ~pi787 & n24973;
  assign n24979 = ~n24977 & ~n24978;
  assign n24980 = ~pi644 & ~n24979;
  assign n24981 = pi715 & ~n24980;
  assign n24982 = pi180 & ~n9829;
  assign n24983 = ~pi753 & n16570;
  assign n24984 = ~n24930 & ~n24983;
  assign n24985 = pi38 & ~n24984;
  assign n24986 = pi753 & n16212;
  assign n24987 = pi180 & ~n16563;
  assign n24988 = ~n24986 & ~n24987;
  assign n24989 = pi39 & ~n24988;
  assign n24990 = ~pi180 & ~pi753;
  assign n24991 = n16514 & n24990;
  assign n24992 = pi180 & pi753;
  assign n24993 = pi180 & ~n16526;
  assign n24994 = ~n20664 & ~n24993;
  assign n24995 = ~pi39 & ~n24994;
  assign n24996 = ~pi38 & ~n24992;
  assign n24997 = ~n24995 & n24996;
  assign n24998 = ~n24991 & n24997;
  assign n24999 = ~n24989 & n24998;
  assign n25000 = n9829 & ~n24985;
  assign n25001 = ~n24999 & n25000;
  assign n25002 = ~n24982 & ~n25001;
  assign n25003 = ~n15777 & ~n25002;
  assign n25004 = n15777 & ~n24926;
  assign n25005 = ~n25003 & ~n25004;
  assign n25006 = ~pi785 & ~n25005;
  assign n25007 = ~n15786 & ~n24926;
  assign n25008 = pi609 & n25003;
  assign n25009 = ~n25007 & ~n25008;
  assign n25010 = pi1155 & ~n25009;
  assign n25011 = ~n16585 & ~n24926;
  assign n25012 = ~pi609 & n25003;
  assign n25013 = ~n25011 & ~n25012;
  assign n25014 = ~pi1155 & ~n25013;
  assign n25015 = ~n25010 & ~n25014;
  assign n25016 = pi785 & ~n25015;
  assign n25017 = ~n25006 & ~n25016;
  assign n25018 = ~pi781 & ~n25017;
  assign n25019 = ~pi618 & n24926;
  assign n25020 = pi618 & n25017;
  assign n25021 = pi1154 & ~n25019;
  assign n25022 = ~n25020 & n25021;
  assign n25023 = ~pi618 & n25017;
  assign n25024 = pi618 & n24926;
  assign n25025 = ~pi1154 & ~n25024;
  assign n25026 = ~n25023 & n25025;
  assign n25027 = ~n25022 & ~n25026;
  assign n25028 = pi781 & ~n25027;
  assign n25029 = ~n25018 & ~n25028;
  assign n25030 = ~pi789 & ~n25029;
  assign n25031 = ~pi619 & n24926;
  assign n25032 = pi619 & n25029;
  assign n25033 = pi1159 & ~n25031;
  assign n25034 = ~n25032 & n25033;
  assign n25035 = ~pi619 & n25029;
  assign n25036 = pi619 & n24926;
  assign n25037 = ~pi1159 & ~n25036;
  assign n25038 = ~n25035 & n25037;
  assign n25039 = ~n25034 & ~n25038;
  assign n25040 = pi789 & ~n25039;
  assign n25041 = ~n25030 & ~n25040;
  assign n25042 = ~n15832 & n25041;
  assign n25043 = n15832 & n24926;
  assign n25044 = ~n25042 & ~n25043;
  assign n25045 = ~n15925 & ~n25044;
  assign n25046 = n15925 & n24926;
  assign n25047 = ~n25045 & ~n25046;
  assign n25048 = ~n15960 & ~n25047;
  assign n25049 = n15960 & n24926;
  assign n25050 = ~n25048 & ~n25049;
  assign n25051 = pi644 & ~n25050;
  assign n25052 = ~pi644 & n24926;
  assign n25053 = ~pi715 & ~n25052;
  assign n25054 = ~n25051 & n25053;
  assign n25055 = pi1160 & ~n25054;
  assign n25056 = ~n24981 & n25055;
  assign n25057 = pi644 & ~n24979;
  assign n25058 = ~pi715 & ~n25057;
  assign n25059 = ~pi644 & ~n25050;
  assign n25060 = pi644 & n24926;
  assign n25061 = pi715 & ~n25060;
  assign n25062 = ~n25059 & n25061;
  assign n25063 = ~pi1160 & ~n25062;
  assign n25064 = ~n25058 & n25063;
  assign n25065 = ~n25056 & ~n25064;
  assign n25066 = pi790 & ~n25065;
  assign n25067 = n19478 & n25047;
  assign n25068 = ~n15959 & n24976;
  assign n25069 = ~n25067 & ~n25068;
  assign n25070 = pi787 & ~n25069;
  assign n25071 = ~n16633 & n25044;
  assign n25072 = ~pi629 & n24966;
  assign n25073 = pi629 & n24970;
  assign n25074 = ~n25072 & ~n25073;
  assign n25075 = ~n25071 & n25074;
  assign n25076 = pi792 & ~n25075;
  assign n25077 = n15828 & ~n24958;
  assign n25078 = ~pi626 & ~n24926;
  assign n25079 = pi626 & ~n25041;
  assign n25080 = n15756 & ~n25078;
  assign n25081 = ~n25079 & n25080;
  assign n25082 = pi626 & ~n24926;
  assign n25083 = ~pi626 & ~n25041;
  assign n25084 = n15757 & ~n25082;
  assign n25085 = ~n25083 & n25084;
  assign n25086 = ~n25077 & ~n25081;
  assign n25087 = ~n25085 & n25086;
  assign n25088 = pi788 & ~n25087;
  assign n25089 = pi618 & ~n24953;
  assign n25090 = pi609 & n24950;
  assign n25091 = ~n24928 & ~n25001;
  assign n25092 = ~pi753 & ~n16808;
  assign n25093 = n18669 & ~n25092;
  assign n25094 = ~pi180 & ~n25093;
  assign n25095 = ~n16921 & ~n24775;
  assign n25096 = pi180 & ~n25095;
  assign n25097 = n6081 & n25096;
  assign n25098 = pi38 & ~n25097;
  assign n25099 = ~n25094 & n25098;
  assign n25100 = ~pi180 & ~n16647;
  assign n25101 = pi180 & ~n17397;
  assign n25102 = ~pi753 & ~n25100;
  assign n25103 = ~n25101 & n25102;
  assign n25104 = ~pi180 & n16653;
  assign n25105 = pi180 & n16657;
  assign n25106 = pi753 & ~n25104;
  assign n25107 = ~n25105 & n25106;
  assign n25108 = ~pi39 & ~n25103;
  assign n25109 = ~n25107 & n25108;
  assign n25110 = pi180 & n16825;
  assign n25111 = ~pi180 & ~n16747;
  assign n25112 = pi753 & ~n25110;
  assign n25113 = ~n25111 & n25112;
  assign n25114 = ~pi180 & n16877;
  assign n25115 = pi180 & n16913;
  assign n25116 = ~pi753 & ~n25114;
  assign n25117 = ~n25115 & n25116;
  assign n25118 = pi39 & ~n25117;
  assign n25119 = ~n25113 & n25118;
  assign n25120 = ~pi38 & ~n25109;
  assign n25121 = ~n25119 & n25120;
  assign n25122 = ~pi702 & ~n25099;
  assign n25123 = ~n25121 & n25122;
  assign n25124 = ~n25091 & ~n25123;
  assign n25125 = ~n24982 & ~n25124;
  assign n25126 = ~pi625 & n25125;
  assign n25127 = pi625 & n25002;
  assign n25128 = ~pi1153 & ~n25127;
  assign n25129 = ~n25126 & n25128;
  assign n25130 = ~pi608 & ~n24943;
  assign n25131 = ~n25129 & n25130;
  assign n25132 = ~pi625 & n25002;
  assign n25133 = pi625 & n25125;
  assign n25134 = pi1153 & ~n25132;
  assign n25135 = ~n25133 & n25134;
  assign n25136 = pi608 & ~n24947;
  assign n25137 = ~n25135 & n25136;
  assign n25138 = ~n25131 & ~n25137;
  assign n25139 = pi778 & ~n25138;
  assign n25140 = ~pi778 & n25125;
  assign n25141 = ~n25139 & ~n25140;
  assign n25142 = ~pi609 & ~n25141;
  assign n25143 = ~pi1155 & ~n25090;
  assign n25144 = ~n25142 & n25143;
  assign n25145 = ~pi660 & ~n25010;
  assign n25146 = ~n25144 & n25145;
  assign n25147 = ~pi609 & n24950;
  assign n25148 = pi609 & ~n25141;
  assign n25149 = pi1155 & ~n25147;
  assign n25150 = ~n25148 & n25149;
  assign n25151 = pi660 & ~n25014;
  assign n25152 = ~n25150 & n25151;
  assign n25153 = ~n25146 & ~n25152;
  assign n25154 = pi785 & ~n25153;
  assign n25155 = ~pi785 & ~n25141;
  assign n25156 = ~n25154 & ~n25155;
  assign n25157 = ~pi618 & ~n25156;
  assign n25158 = ~pi1154 & ~n25089;
  assign n25159 = ~n25157 & n25158;
  assign n25160 = ~pi627 & ~n25022;
  assign n25161 = ~n25159 & n25160;
  assign n25162 = ~pi618 & ~n24953;
  assign n25163 = pi618 & ~n25156;
  assign n25164 = pi1154 & ~n25162;
  assign n25165 = ~n25163 & n25164;
  assign n25166 = pi627 & ~n25026;
  assign n25167 = ~n25165 & n25166;
  assign n25168 = ~n25161 & ~n25167;
  assign n25169 = pi781 & ~n25168;
  assign n25170 = ~pi781 & ~n25156;
  assign n25171 = ~n25169 & ~n25170;
  assign n25172 = ~pi789 & n25171;
  assign n25173 = ~pi619 & n24955;
  assign n25174 = pi619 & ~n25171;
  assign n25175 = pi1159 & ~n25173;
  assign n25176 = ~n25174 & n25175;
  assign n25177 = pi648 & ~n25038;
  assign n25178 = ~n25176 & n25177;
  assign n25179 = ~pi619 & ~n25171;
  assign n25180 = pi619 & n24955;
  assign n25181 = ~pi1159 & ~n25180;
  assign n25182 = ~n25179 & n25181;
  assign n25183 = ~pi648 & ~n25034;
  assign n25184 = ~n25182 & n25183;
  assign n25185 = pi789 & ~n25178;
  assign n25186 = ~n25184 & n25185;
  assign n25187 = n15833 & ~n25172;
  assign n25188 = ~n25186 & n25187;
  assign n25189 = ~n16644 & ~n25088;
  assign n25190 = ~n25188 & n25189;
  assign n25191 = ~n25076 & ~n25190;
  assign n25192 = n18841 & ~n25191;
  assign n25193 = pi644 & ~n25054;
  assign n25194 = ~n25063 & ~n25193;
  assign n25195 = ~n22949 & ~n25194;
  assign n25196 = pi790 & ~n25195;
  assign n25197 = ~n25070 & ~n25196;
  assign n25198 = ~n25192 & n25197;
  assign n25199 = ~n25066 & ~n25198;
  assign n25200 = ~po1038 & ~n25199;
  assign n25201 = ~pi832 & ~n24925;
  assign n25202 = ~n25200 & n25201;
  assign po337 = ~n24924 & ~n25202;
  assign n25204 = ~pi181 & ~n2923;
  assign n25205 = ~pi709 & n15726;
  assign n25206 = ~n25204 & ~n25205;
  assign n25207 = ~pi778 & ~n25206;
  assign n25208 = ~pi625 & n25205;
  assign n25209 = ~n25206 & ~n25208;
  assign n25210 = pi1153 & ~n25209;
  assign n25211 = ~pi1153 & ~n25204;
  assign n25212 = ~n25208 & n25211;
  assign n25213 = pi778 & ~n25212;
  assign n25214 = ~n25210 & n25213;
  assign n25215 = ~n25207 & ~n25214;
  assign n25216 = ~n15742 & ~n25215;
  assign n25217 = ~n15748 & n25216;
  assign n25218 = ~n15754 & n25217;
  assign n25219 = ~n15760 & n25218;
  assign n25220 = ~n15766 & n25219;
  assign n25221 = n19394 & n25220;
  assign n25222 = ~n19394 & n25204;
  assign n25223 = ~n25221 & ~n25222;
  assign n25224 = ~n15959 & n25223;
  assign n25225 = n15925 & n25204;
  assign n25226 = ~pi754 & n15781;
  assign n25227 = ~n25204 & ~n25226;
  assign n25228 = ~n15778 & ~n25227;
  assign n25229 = ~pi785 & ~n25228;
  assign n25230 = n16585 & n25226;
  assign n25231 = n25228 & ~n25230;
  assign n25232 = pi1155 & ~n25231;
  assign n25233 = ~pi1155 & ~n25204;
  assign n25234 = ~n25230 & n25233;
  assign n25235 = ~n25232 & ~n25234;
  assign n25236 = pi785 & ~n25235;
  assign n25237 = ~n25229 & ~n25236;
  assign n25238 = ~pi781 & ~n25237;
  assign n25239 = ~n15797 & n25237;
  assign n25240 = pi1154 & ~n25239;
  assign n25241 = ~n15800 & n25237;
  assign n25242 = ~pi1154 & ~n25241;
  assign n25243 = ~n25240 & ~n25242;
  assign n25244 = pi781 & ~n25243;
  assign n25245 = ~n25238 & ~n25244;
  assign n25246 = ~n21915 & n25245;
  assign n25247 = ~n15832 & ~n25246;
  assign n25248 = n15832 & ~n25204;
  assign n25249 = ~n25247 & ~n25248;
  assign n25250 = ~n15925 & n25249;
  assign n25251 = n19478 & ~n25225;
  assign n25252 = ~n25250 & n25251;
  assign n25253 = ~n25224 & ~n25252;
  assign n25254 = pi787 & ~n25253;
  assign n25255 = n15763 & n25249;
  assign n25256 = n15772 & n25219;
  assign n25257 = ~pi629 & ~n25256;
  assign n25258 = ~n25255 & n25257;
  assign n25259 = n15762 & n25249;
  assign n25260 = n15909 & n25219;
  assign n25261 = pi629 & ~n25260;
  assign n25262 = ~n25259 & n25261;
  assign n25263 = pi792 & ~n25258;
  assign n25264 = ~n25262 & n25263;
  assign n25265 = ~n21932 & n25245;
  assign n25266 = pi648 & ~n25265;
  assign n25267 = n21935 & ~n25217;
  assign n25268 = ~n25266 & ~n25267;
  assign n25269 = ~pi1159 & ~n25268;
  assign n25270 = ~pi619 & ~n25217;
  assign n25271 = pi648 & ~n25270;
  assign n25272 = n21942 & n25245;
  assign n25273 = pi1159 & ~n25271;
  assign n25274 = ~n25272 & n25273;
  assign n25275 = ~n25269 & ~n25274;
  assign n25276 = pi789 & ~n25275;
  assign n25277 = pi609 & ~n25215;
  assign n25278 = ~n15780 & ~n25206;
  assign n25279 = pi625 & n25278;
  assign n25280 = n25227 & ~n25278;
  assign n25281 = ~n25279 & ~n25280;
  assign n25282 = n25211 & ~n25281;
  assign n25283 = ~pi608 & ~n25210;
  assign n25284 = ~n25282 & n25283;
  assign n25285 = pi1153 & n25227;
  assign n25286 = ~n25279 & n25285;
  assign n25287 = pi608 & ~n25212;
  assign n25288 = ~n25286 & n25287;
  assign n25289 = ~n25284 & ~n25288;
  assign n25290 = pi778 & ~n25289;
  assign n25291 = ~pi778 & ~n25280;
  assign n25292 = ~n25290 & ~n25291;
  assign n25293 = ~pi609 & ~n25292;
  assign n25294 = ~pi1155 & ~n25277;
  assign n25295 = ~n25293 & n25294;
  assign n25296 = ~pi660 & ~n25232;
  assign n25297 = ~n25295 & n25296;
  assign n25298 = ~pi609 & ~n25215;
  assign n25299 = pi609 & ~n25292;
  assign n25300 = pi1155 & ~n25298;
  assign n25301 = ~n25299 & n25300;
  assign n25302 = pi660 & ~n25234;
  assign n25303 = ~n25301 & n25302;
  assign n25304 = ~n25297 & ~n25303;
  assign n25305 = pi785 & ~n25304;
  assign n25306 = ~pi785 & ~n25292;
  assign n25307 = ~n25305 & ~n25306;
  assign n25308 = ~pi781 & n25307;
  assign n25309 = pi618 & n25216;
  assign n25310 = ~pi618 & ~n25307;
  assign n25311 = ~pi1154 & ~n25309;
  assign n25312 = ~n25310 & n25311;
  assign n25313 = ~pi627 & ~n25240;
  assign n25314 = ~n25312 & n25313;
  assign n25315 = ~pi618 & n25216;
  assign n25316 = pi618 & ~n25307;
  assign n25317 = pi1154 & ~n25315;
  assign n25318 = ~n25316 & n25317;
  assign n25319 = pi627 & ~n25242;
  assign n25320 = ~n25318 & n25319;
  assign n25321 = pi781 & ~n25314;
  assign n25322 = ~n25320 & n25321;
  assign n25323 = ~n25276 & ~n25308;
  assign n25324 = ~n25322 & n25323;
  assign n25325 = n18969 & n25275;
  assign n25326 = ~n25324 & ~n25325;
  assign n25327 = n15833 & ~n25326;
  assign n25328 = n15828 & n25218;
  assign n25329 = ~pi626 & ~n25204;
  assign n25330 = pi626 & ~n25246;
  assign n25331 = n15756 & ~n25329;
  assign n25332 = ~n25330 & n25331;
  assign n25333 = pi626 & ~n25204;
  assign n25334 = ~pi626 & ~n25246;
  assign n25335 = n15757 & ~n25333;
  assign n25336 = ~n25334 & n25335;
  assign n25337 = ~n25328 & ~n25332;
  assign n25338 = ~n25336 & n25337;
  assign n25339 = pi788 & ~n25338;
  assign n25340 = ~n25327 & ~n25339;
  assign n25341 = ~n16644 & ~n25340;
  assign n25342 = n18841 & ~n25264;
  assign n25343 = ~n25341 & n25342;
  assign n25344 = ~n25254 & ~n25343;
  assign n25345 = ~pi790 & n25344;
  assign n25346 = pi787 & ~n25223;
  assign n25347 = ~pi787 & n25220;
  assign n25348 = ~n25346 & ~n25347;
  assign n25349 = ~pi644 & ~n25348;
  assign n25350 = pi644 & n25344;
  assign n25351 = pi715 & ~n25349;
  assign n25352 = ~n25350 & n25351;
  assign n25353 = ~n19771 & n25204;
  assign n25354 = ~n15960 & n25250;
  assign n25355 = ~n25353 & ~n25354;
  assign n25356 = pi644 & ~n25355;
  assign n25357 = ~pi644 & n25204;
  assign n25358 = ~pi715 & ~n25357;
  assign n25359 = ~n25356 & n25358;
  assign n25360 = pi1160 & ~n25359;
  assign n25361 = ~n25352 & n25360;
  assign n25362 = ~pi644 & ~n25355;
  assign n25363 = pi644 & n25204;
  assign n25364 = pi715 & ~n25363;
  assign n25365 = ~n25362 & n25364;
  assign n25366 = pi644 & ~n25348;
  assign n25367 = ~pi644 & n25344;
  assign n25368 = ~pi715 & ~n25366;
  assign n25369 = ~n25367 & n25368;
  assign n25370 = ~pi1160 & ~n25365;
  assign n25371 = ~n25369 & n25370;
  assign n25372 = ~n25361 & ~n25371;
  assign n25373 = pi790 & ~n25372;
  assign n25374 = pi832 & ~n25345;
  assign n25375 = ~n25373 & n25374;
  assign n25376 = ~pi181 & po1038;
  assign n25377 = ~pi181 & ~n16219;
  assign n25378 = n15747 & ~n25377;
  assign n25379 = ~pi709 & n9829;
  assign n25380 = n25377 & ~n25379;
  assign n25381 = ~pi181 & ~n16228;
  assign n25382 = n16227 & ~n25381;
  assign n25383 = ~pi181 & ~n17276;
  assign n25384 = ~pi38 & ~pi181;
  assign n25385 = n19350 & ~n25384;
  assign n25386 = ~n25383 & ~n25385;
  assign n25387 = ~pi709 & ~n25382;
  assign n25388 = ~n25386 & n25387;
  assign n25389 = ~n25380 & ~n25388;
  assign n25390 = ~pi778 & n25389;
  assign n25391 = ~pi625 & n25377;
  assign n25392 = pi625 & ~n25389;
  assign n25393 = pi1153 & ~n25391;
  assign n25394 = ~n25392 & n25393;
  assign n25395 = pi625 & n25377;
  assign n25396 = ~pi625 & ~n25389;
  assign n25397 = ~pi1153 & ~n25395;
  assign n25398 = ~n25396 & n25397;
  assign n25399 = ~n25394 & ~n25398;
  assign n25400 = pi778 & ~n25399;
  assign n25401 = ~n25390 & ~n25400;
  assign n25402 = ~n15741 & n25401;
  assign n25403 = n15741 & n25377;
  assign n25404 = ~n25402 & ~n25403;
  assign n25405 = ~n15747 & n25404;
  assign n25406 = ~n25378 & ~n25405;
  assign n25407 = ~n15753 & n25406;
  assign n25408 = n15753 & n25377;
  assign n25409 = ~n25407 & ~n25408;
  assign n25410 = ~n15759 & ~n25409;
  assign n25411 = n15759 & n25377;
  assign n25412 = ~n25410 & ~n25411;
  assign n25413 = ~pi792 & n25412;
  assign n25414 = ~pi628 & n25377;
  assign n25415 = pi628 & ~n25412;
  assign n25416 = pi1156 & ~n25414;
  assign n25417 = ~n25415 & n25416;
  assign n25418 = pi628 & n25377;
  assign n25419 = ~pi628 & ~n25412;
  assign n25420 = ~pi1156 & ~n25418;
  assign n25421 = ~n25419 & n25420;
  assign n25422 = ~n25417 & ~n25421;
  assign n25423 = pi792 & ~n25422;
  assign n25424 = ~n25413 & ~n25423;
  assign n25425 = n19394 & n25424;
  assign n25426 = ~n19394 & n25377;
  assign n25427 = ~n25425 & ~n25426;
  assign n25428 = pi787 & ~n25427;
  assign n25429 = ~pi787 & n25424;
  assign n25430 = ~n25428 & ~n25429;
  assign n25431 = ~pi644 & ~n25430;
  assign n25432 = pi715 & ~n25431;
  assign n25433 = pi181 & ~n9829;
  assign n25434 = ~pi754 & n16570;
  assign n25435 = ~n25381 & ~n25434;
  assign n25436 = pi38 & ~n25435;
  assign n25437 = pi754 & n16212;
  assign n25438 = pi181 & ~n16563;
  assign n25439 = ~n25437 & ~n25438;
  assign n25440 = pi39 & ~n25439;
  assign n25441 = ~pi181 & ~pi754;
  assign n25442 = n16514 & n25441;
  assign n25443 = pi181 & pi754;
  assign n25444 = pi181 & ~n16526;
  assign n25445 = ~n20719 & ~n25444;
  assign n25446 = ~pi39 & ~n25445;
  assign n25447 = ~pi38 & ~n25443;
  assign n25448 = ~n25446 & n25447;
  assign n25449 = ~n25442 & n25448;
  assign n25450 = ~n25440 & n25449;
  assign n25451 = n9829 & ~n25436;
  assign n25452 = ~n25450 & n25451;
  assign n25453 = ~n25433 & ~n25452;
  assign n25454 = ~n15777 & ~n25453;
  assign n25455 = n15777 & ~n25377;
  assign n25456 = ~n25454 & ~n25455;
  assign n25457 = ~pi785 & ~n25456;
  assign n25458 = ~n15786 & ~n25377;
  assign n25459 = pi609 & n25454;
  assign n25460 = ~n25458 & ~n25459;
  assign n25461 = pi1155 & ~n25460;
  assign n25462 = ~n16585 & ~n25377;
  assign n25463 = ~pi609 & n25454;
  assign n25464 = ~n25462 & ~n25463;
  assign n25465 = ~pi1155 & ~n25464;
  assign n25466 = ~n25461 & ~n25465;
  assign n25467 = pi785 & ~n25466;
  assign n25468 = ~n25457 & ~n25467;
  assign n25469 = ~pi781 & ~n25468;
  assign n25470 = ~pi618 & n25377;
  assign n25471 = pi618 & n25468;
  assign n25472 = pi1154 & ~n25470;
  assign n25473 = ~n25471 & n25472;
  assign n25474 = ~pi618 & n25468;
  assign n25475 = pi618 & n25377;
  assign n25476 = ~pi1154 & ~n25475;
  assign n25477 = ~n25474 & n25476;
  assign n25478 = ~n25473 & ~n25477;
  assign n25479 = pi781 & ~n25478;
  assign n25480 = ~n25469 & ~n25479;
  assign n25481 = ~pi789 & ~n25480;
  assign n25482 = ~pi619 & n25377;
  assign n25483 = pi619 & n25480;
  assign n25484 = pi1159 & ~n25482;
  assign n25485 = ~n25483 & n25484;
  assign n25486 = ~pi619 & n25480;
  assign n25487 = pi619 & n25377;
  assign n25488 = ~pi1159 & ~n25487;
  assign n25489 = ~n25486 & n25488;
  assign n25490 = ~n25485 & ~n25489;
  assign n25491 = pi789 & ~n25490;
  assign n25492 = ~n25481 & ~n25491;
  assign n25493 = ~n15832 & n25492;
  assign n25494 = n15832 & n25377;
  assign n25495 = ~n25493 & ~n25494;
  assign n25496 = ~n15925 & ~n25495;
  assign n25497 = n15925 & n25377;
  assign n25498 = ~n25496 & ~n25497;
  assign n25499 = ~n15960 & ~n25498;
  assign n25500 = n15960 & n25377;
  assign n25501 = ~n25499 & ~n25500;
  assign n25502 = pi644 & ~n25501;
  assign n25503 = ~pi644 & n25377;
  assign n25504 = ~pi715 & ~n25503;
  assign n25505 = ~n25502 & n25504;
  assign n25506 = pi1160 & ~n25505;
  assign n25507 = ~n25432 & n25506;
  assign n25508 = pi644 & ~n25430;
  assign n25509 = ~pi715 & ~n25508;
  assign n25510 = ~pi644 & ~n25501;
  assign n25511 = pi644 & n25377;
  assign n25512 = pi715 & ~n25511;
  assign n25513 = ~n25510 & n25512;
  assign n25514 = ~pi1160 & ~n25513;
  assign n25515 = ~n25509 & n25514;
  assign n25516 = ~n25507 & ~n25515;
  assign n25517 = pi790 & ~n25516;
  assign n25518 = n19478 & n25498;
  assign n25519 = ~n15959 & n25427;
  assign n25520 = ~n25518 & ~n25519;
  assign n25521 = pi787 & ~n25520;
  assign n25522 = ~n16633 & n25495;
  assign n25523 = ~pi629 & n25417;
  assign n25524 = pi629 & n25421;
  assign n25525 = ~n25523 & ~n25524;
  assign n25526 = ~n25522 & n25525;
  assign n25527 = pi792 & ~n25526;
  assign n25528 = n15828 & ~n25409;
  assign n25529 = ~pi626 & ~n25377;
  assign n25530 = pi626 & ~n25492;
  assign n25531 = n15756 & ~n25529;
  assign n25532 = ~n25530 & n25531;
  assign n25533 = pi626 & ~n25377;
  assign n25534 = ~pi626 & ~n25492;
  assign n25535 = n15757 & ~n25533;
  assign n25536 = ~n25534 & n25535;
  assign n25537 = ~n25528 & ~n25532;
  assign n25538 = ~n25536 & n25537;
  assign n25539 = pi788 & ~n25538;
  assign n25540 = pi618 & ~n25404;
  assign n25541 = pi609 & n25401;
  assign n25542 = ~n25379 & ~n25452;
  assign n25543 = ~pi754 & ~n16808;
  assign n25544 = n18669 & ~n25543;
  assign n25545 = ~pi181 & ~n25544;
  assign n25546 = ~n16921 & ~n25226;
  assign n25547 = pi181 & ~n25546;
  assign n25548 = n6081 & n25547;
  assign n25549 = pi38 & ~n25548;
  assign n25550 = ~n25545 & n25549;
  assign n25551 = ~pi181 & ~n16647;
  assign n25552 = pi181 & ~n17397;
  assign n25553 = ~pi754 & ~n25551;
  assign n25554 = ~n25552 & n25553;
  assign n25555 = ~pi181 & n16653;
  assign n25556 = pi181 & n16657;
  assign n25557 = pi754 & ~n25555;
  assign n25558 = ~n25556 & n25557;
  assign n25559 = ~pi39 & ~n25554;
  assign n25560 = ~n25558 & n25559;
  assign n25561 = pi181 & n16825;
  assign n25562 = ~pi181 & ~n16747;
  assign n25563 = pi754 & ~n25561;
  assign n25564 = ~n25562 & n25563;
  assign n25565 = ~pi181 & n16877;
  assign n25566 = pi181 & n16913;
  assign n25567 = ~pi754 & ~n25565;
  assign n25568 = ~n25566 & n25567;
  assign n25569 = pi39 & ~n25568;
  assign n25570 = ~n25564 & n25569;
  assign n25571 = ~pi38 & ~n25560;
  assign n25572 = ~n25570 & n25571;
  assign n25573 = ~pi709 & ~n25550;
  assign n25574 = ~n25572 & n25573;
  assign n25575 = ~n25542 & ~n25574;
  assign n25576 = ~n25433 & ~n25575;
  assign n25577 = ~pi625 & n25576;
  assign n25578 = pi625 & n25453;
  assign n25579 = ~pi1153 & ~n25578;
  assign n25580 = ~n25577 & n25579;
  assign n25581 = ~pi608 & ~n25394;
  assign n25582 = ~n25580 & n25581;
  assign n25583 = ~pi625 & n25453;
  assign n25584 = pi625 & n25576;
  assign n25585 = pi1153 & ~n25583;
  assign n25586 = ~n25584 & n25585;
  assign n25587 = pi608 & ~n25398;
  assign n25588 = ~n25586 & n25587;
  assign n25589 = ~n25582 & ~n25588;
  assign n25590 = pi778 & ~n25589;
  assign n25591 = ~pi778 & n25576;
  assign n25592 = ~n25590 & ~n25591;
  assign n25593 = ~pi609 & ~n25592;
  assign n25594 = ~pi1155 & ~n25541;
  assign n25595 = ~n25593 & n25594;
  assign n25596 = ~pi660 & ~n25461;
  assign n25597 = ~n25595 & n25596;
  assign n25598 = ~pi609 & n25401;
  assign n25599 = pi609 & ~n25592;
  assign n25600 = pi1155 & ~n25598;
  assign n25601 = ~n25599 & n25600;
  assign n25602 = pi660 & ~n25465;
  assign n25603 = ~n25601 & n25602;
  assign n25604 = ~n25597 & ~n25603;
  assign n25605 = pi785 & ~n25604;
  assign n25606 = ~pi785 & ~n25592;
  assign n25607 = ~n25605 & ~n25606;
  assign n25608 = ~pi618 & ~n25607;
  assign n25609 = ~pi1154 & ~n25540;
  assign n25610 = ~n25608 & n25609;
  assign n25611 = ~pi627 & ~n25473;
  assign n25612 = ~n25610 & n25611;
  assign n25613 = ~pi618 & ~n25404;
  assign n25614 = pi618 & ~n25607;
  assign n25615 = pi1154 & ~n25613;
  assign n25616 = ~n25614 & n25615;
  assign n25617 = pi627 & ~n25477;
  assign n25618 = ~n25616 & n25617;
  assign n25619 = ~n25612 & ~n25618;
  assign n25620 = pi781 & ~n25619;
  assign n25621 = ~pi781 & ~n25607;
  assign n25622 = ~n25620 & ~n25621;
  assign n25623 = ~pi789 & n25622;
  assign n25624 = ~pi619 & n25406;
  assign n25625 = pi619 & ~n25622;
  assign n25626 = pi1159 & ~n25624;
  assign n25627 = ~n25625 & n25626;
  assign n25628 = pi648 & ~n25489;
  assign n25629 = ~n25627 & n25628;
  assign n25630 = ~pi619 & ~n25622;
  assign n25631 = pi619 & n25406;
  assign n25632 = ~pi1159 & ~n25631;
  assign n25633 = ~n25630 & n25632;
  assign n25634 = ~pi648 & ~n25485;
  assign n25635 = ~n25633 & n25634;
  assign n25636 = pi789 & ~n25629;
  assign n25637 = ~n25635 & n25636;
  assign n25638 = n15833 & ~n25623;
  assign n25639 = ~n25637 & n25638;
  assign n25640 = ~n16644 & ~n25539;
  assign n25641 = ~n25639 & n25640;
  assign n25642 = ~n25527 & ~n25641;
  assign n25643 = n18841 & ~n25642;
  assign n25644 = pi644 & ~n25505;
  assign n25645 = ~n25514 & ~n25644;
  assign n25646 = ~n22949 & ~n25645;
  assign n25647 = pi790 & ~n25646;
  assign n25648 = ~n25521 & ~n25647;
  assign n25649 = ~n25643 & n25648;
  assign n25650 = ~n25517 & ~n25649;
  assign n25651 = ~po1038 & ~n25650;
  assign n25652 = ~pi832 & ~n25376;
  assign n25653 = ~n25651 & n25652;
  assign po338 = ~n25375 & ~n25653;
  assign n25655 = ~pi182 & ~n2923;
  assign n25656 = ~pi734 & n15726;
  assign n25657 = ~n25655 & ~n25656;
  assign n25658 = ~pi778 & ~n25657;
  assign n25659 = ~pi625 & n25656;
  assign n25660 = ~n25657 & ~n25659;
  assign n25661 = pi1153 & ~n25660;
  assign n25662 = ~pi1153 & ~n25655;
  assign n25663 = ~n25659 & n25662;
  assign n25664 = pi778 & ~n25663;
  assign n25665 = ~n25661 & n25664;
  assign n25666 = ~n25658 & ~n25665;
  assign n25667 = ~n15742 & ~n25666;
  assign n25668 = ~n15748 & n25667;
  assign n25669 = ~n15754 & n25668;
  assign n25670 = ~n15760 & n25669;
  assign n25671 = ~n15766 & n25670;
  assign n25672 = n19394 & n25671;
  assign n25673 = ~n19394 & n25655;
  assign n25674 = ~n25672 & ~n25673;
  assign n25675 = ~n15959 & n25674;
  assign n25676 = n15925 & n25655;
  assign n25677 = ~pi756 & n15781;
  assign n25678 = ~n25655 & ~n25677;
  assign n25679 = ~n15778 & ~n25678;
  assign n25680 = ~pi785 & ~n25679;
  assign n25681 = n16585 & n25677;
  assign n25682 = n25679 & ~n25681;
  assign n25683 = pi1155 & ~n25682;
  assign n25684 = ~pi1155 & ~n25655;
  assign n25685 = ~n25681 & n25684;
  assign n25686 = ~n25683 & ~n25685;
  assign n25687 = pi785 & ~n25686;
  assign n25688 = ~n25680 & ~n25687;
  assign n25689 = ~pi781 & ~n25688;
  assign n25690 = ~n15797 & n25688;
  assign n25691 = pi1154 & ~n25690;
  assign n25692 = ~n15800 & n25688;
  assign n25693 = ~pi1154 & ~n25692;
  assign n25694 = ~n25691 & ~n25693;
  assign n25695 = pi781 & ~n25694;
  assign n25696 = ~n25689 & ~n25695;
  assign n25697 = ~n21915 & n25696;
  assign n25698 = ~n15832 & ~n25697;
  assign n25699 = n15832 & ~n25655;
  assign n25700 = ~n25698 & ~n25699;
  assign n25701 = ~n15925 & n25700;
  assign n25702 = n19478 & ~n25676;
  assign n25703 = ~n25701 & n25702;
  assign n25704 = ~n25675 & ~n25703;
  assign n25705 = pi787 & ~n25704;
  assign n25706 = n15763 & n25700;
  assign n25707 = n15772 & n25670;
  assign n25708 = ~pi629 & ~n25707;
  assign n25709 = ~n25706 & n25708;
  assign n25710 = n15762 & n25700;
  assign n25711 = n15909 & n25670;
  assign n25712 = pi629 & ~n25711;
  assign n25713 = ~n25710 & n25712;
  assign n25714 = pi792 & ~n25709;
  assign n25715 = ~n25713 & n25714;
  assign n25716 = ~n21932 & n25696;
  assign n25717 = pi648 & ~n25716;
  assign n25718 = n21935 & ~n25668;
  assign n25719 = ~n25717 & ~n25718;
  assign n25720 = ~pi1159 & ~n25719;
  assign n25721 = ~pi619 & ~n25668;
  assign n25722 = pi648 & ~n25721;
  assign n25723 = n21942 & n25696;
  assign n25724 = pi1159 & ~n25722;
  assign n25725 = ~n25723 & n25724;
  assign n25726 = ~n25720 & ~n25725;
  assign n25727 = pi789 & ~n25726;
  assign n25728 = pi609 & ~n25666;
  assign n25729 = ~n15780 & ~n25657;
  assign n25730 = pi625 & n25729;
  assign n25731 = n25678 & ~n25729;
  assign n25732 = ~n25730 & ~n25731;
  assign n25733 = n25662 & ~n25732;
  assign n25734 = ~pi608 & ~n25661;
  assign n25735 = ~n25733 & n25734;
  assign n25736 = pi1153 & n25678;
  assign n25737 = ~n25730 & n25736;
  assign n25738 = pi608 & ~n25663;
  assign n25739 = ~n25737 & n25738;
  assign n25740 = ~n25735 & ~n25739;
  assign n25741 = pi778 & ~n25740;
  assign n25742 = ~pi778 & ~n25731;
  assign n25743 = ~n25741 & ~n25742;
  assign n25744 = ~pi609 & ~n25743;
  assign n25745 = ~pi1155 & ~n25728;
  assign n25746 = ~n25744 & n25745;
  assign n25747 = ~pi660 & ~n25683;
  assign n25748 = ~n25746 & n25747;
  assign n25749 = ~pi609 & ~n25666;
  assign n25750 = pi609 & ~n25743;
  assign n25751 = pi1155 & ~n25749;
  assign n25752 = ~n25750 & n25751;
  assign n25753 = pi660 & ~n25685;
  assign n25754 = ~n25752 & n25753;
  assign n25755 = ~n25748 & ~n25754;
  assign n25756 = pi785 & ~n25755;
  assign n25757 = ~pi785 & ~n25743;
  assign n25758 = ~n25756 & ~n25757;
  assign n25759 = ~pi781 & n25758;
  assign n25760 = pi618 & n25667;
  assign n25761 = ~pi618 & ~n25758;
  assign n25762 = ~pi1154 & ~n25760;
  assign n25763 = ~n25761 & n25762;
  assign n25764 = ~pi627 & ~n25691;
  assign n25765 = ~n25763 & n25764;
  assign n25766 = ~pi618 & n25667;
  assign n25767 = pi618 & ~n25758;
  assign n25768 = pi1154 & ~n25766;
  assign n25769 = ~n25767 & n25768;
  assign n25770 = pi627 & ~n25693;
  assign n25771 = ~n25769 & n25770;
  assign n25772 = pi781 & ~n25765;
  assign n25773 = ~n25771 & n25772;
  assign n25774 = ~n25727 & ~n25759;
  assign n25775 = ~n25773 & n25774;
  assign n25776 = n18969 & n25726;
  assign n25777 = ~n25775 & ~n25776;
  assign n25778 = n15833 & ~n25777;
  assign n25779 = n15828 & n25669;
  assign n25780 = ~pi626 & ~n25655;
  assign n25781 = pi626 & ~n25697;
  assign n25782 = n15756 & ~n25780;
  assign n25783 = ~n25781 & n25782;
  assign n25784 = pi626 & ~n25655;
  assign n25785 = ~pi626 & ~n25697;
  assign n25786 = n15757 & ~n25784;
  assign n25787 = ~n25785 & n25786;
  assign n25788 = ~n25779 & ~n25783;
  assign n25789 = ~n25787 & n25788;
  assign n25790 = pi788 & ~n25789;
  assign n25791 = ~n25778 & ~n25790;
  assign n25792 = ~n16644 & ~n25791;
  assign n25793 = n18841 & ~n25715;
  assign n25794 = ~n25792 & n25793;
  assign n25795 = ~n25705 & ~n25794;
  assign n25796 = ~pi790 & n25795;
  assign n25797 = pi787 & ~n25674;
  assign n25798 = ~pi787 & n25671;
  assign n25799 = ~n25797 & ~n25798;
  assign n25800 = ~pi644 & ~n25799;
  assign n25801 = pi644 & n25795;
  assign n25802 = pi715 & ~n25800;
  assign n25803 = ~n25801 & n25802;
  assign n25804 = ~n19771 & n25655;
  assign n25805 = ~n15960 & n25701;
  assign n25806 = ~n25804 & ~n25805;
  assign n25807 = pi644 & ~n25806;
  assign n25808 = ~pi644 & n25655;
  assign n25809 = ~pi715 & ~n25808;
  assign n25810 = ~n25807 & n25809;
  assign n25811 = pi1160 & ~n25810;
  assign n25812 = ~n25803 & n25811;
  assign n25813 = ~pi644 & ~n25806;
  assign n25814 = pi644 & n25655;
  assign n25815 = pi715 & ~n25814;
  assign n25816 = ~n25813 & n25815;
  assign n25817 = pi644 & ~n25799;
  assign n25818 = ~pi644 & n25795;
  assign n25819 = ~pi715 & ~n25817;
  assign n25820 = ~n25818 & n25819;
  assign n25821 = ~pi1160 & ~n25816;
  assign n25822 = ~n25820 & n25821;
  assign n25823 = ~n25812 & ~n25822;
  assign n25824 = pi790 & ~n25823;
  assign n25825 = pi832 & ~n25796;
  assign n25826 = ~n25824 & n25825;
  assign n25827 = ~pi182 & po1038;
  assign n25828 = ~pi182 & ~n16219;
  assign n25829 = n15747 & ~n25828;
  assign n25830 = ~pi734 & n9829;
  assign n25831 = n25828 & ~n25830;
  assign n25832 = ~pi182 & ~n16228;
  assign n25833 = n16227 & ~n25832;
  assign n25834 = ~pi182 & ~n17276;
  assign n25835 = ~pi38 & ~pi182;
  assign n25836 = n19350 & ~n25835;
  assign n25837 = ~n25834 & ~n25836;
  assign n25838 = ~pi734 & ~n25833;
  assign n25839 = ~n25837 & n25838;
  assign n25840 = ~n25831 & ~n25839;
  assign n25841 = ~pi778 & n25840;
  assign n25842 = ~pi625 & n25828;
  assign n25843 = pi625 & ~n25840;
  assign n25844 = pi1153 & ~n25842;
  assign n25845 = ~n25843 & n25844;
  assign n25846 = pi625 & n25828;
  assign n25847 = ~pi625 & ~n25840;
  assign n25848 = ~pi1153 & ~n25846;
  assign n25849 = ~n25847 & n25848;
  assign n25850 = ~n25845 & ~n25849;
  assign n25851 = pi778 & ~n25850;
  assign n25852 = ~n25841 & ~n25851;
  assign n25853 = ~n15741 & n25852;
  assign n25854 = n15741 & n25828;
  assign n25855 = ~n25853 & ~n25854;
  assign n25856 = ~n15747 & n25855;
  assign n25857 = ~n25829 & ~n25856;
  assign n25858 = ~n15753 & n25857;
  assign n25859 = n15753 & n25828;
  assign n25860 = ~n25858 & ~n25859;
  assign n25861 = ~n15759 & ~n25860;
  assign n25862 = n15759 & n25828;
  assign n25863 = ~n25861 & ~n25862;
  assign n25864 = ~pi792 & n25863;
  assign n25865 = ~pi628 & n25828;
  assign n25866 = pi628 & ~n25863;
  assign n25867 = pi1156 & ~n25865;
  assign n25868 = ~n25866 & n25867;
  assign n25869 = pi628 & n25828;
  assign n25870 = ~pi628 & ~n25863;
  assign n25871 = ~pi1156 & ~n25869;
  assign n25872 = ~n25870 & n25871;
  assign n25873 = ~n25868 & ~n25872;
  assign n25874 = pi792 & ~n25873;
  assign n25875 = ~n25864 & ~n25874;
  assign n25876 = pi647 & n25875;
  assign n25877 = ~pi647 & n25828;
  assign n25878 = ~n25876 & ~n25877;
  assign n25879 = pi1157 & n25878;
  assign n25880 = ~pi647 & n25875;
  assign n25881 = pi647 & n25828;
  assign n25882 = ~pi1157 & ~n25881;
  assign n25883 = ~n25880 & n25882;
  assign n25884 = ~n25879 & ~n25883;
  assign n25885 = pi787 & ~n25884;
  assign n25886 = ~pi787 & ~n25875;
  assign n25887 = ~n25885 & ~n25886;
  assign n25888 = ~pi644 & n25887;
  assign n25889 = pi715 & ~n25888;
  assign n25890 = pi182 & ~n9829;
  assign n25891 = ~pi182 & n16514;
  assign n25892 = pi182 & ~n16565;
  assign n25893 = ~pi756 & ~n25891;
  assign n25894 = ~n25892 & n25893;
  assign n25895 = ~pi182 & pi756;
  assign n25896 = ~n16214 & n25895;
  assign n25897 = ~n25894 & ~n25896;
  assign n25898 = ~pi38 & ~n25897;
  assign n25899 = ~pi756 & n16570;
  assign n25900 = ~n25832 & ~n25899;
  assign n25901 = pi38 & ~n25900;
  assign n25902 = n9829 & ~n25901;
  assign n25903 = ~n25898 & n25902;
  assign n25904 = ~n25890 & ~n25903;
  assign n25905 = ~n15777 & ~n25904;
  assign n25906 = n15777 & ~n25828;
  assign n25907 = ~n25905 & ~n25906;
  assign n25908 = ~pi785 & ~n25907;
  assign n25909 = ~n15786 & ~n25828;
  assign n25910 = pi609 & n25905;
  assign n25911 = ~n25909 & ~n25910;
  assign n25912 = pi1155 & ~n25911;
  assign n25913 = ~n16585 & ~n25828;
  assign n25914 = ~pi609 & n25905;
  assign n25915 = ~n25913 & ~n25914;
  assign n25916 = ~pi1155 & ~n25915;
  assign n25917 = ~n25912 & ~n25916;
  assign n25918 = pi785 & ~n25917;
  assign n25919 = ~n25908 & ~n25918;
  assign n25920 = ~pi781 & ~n25919;
  assign n25921 = ~pi618 & n25828;
  assign n25922 = pi618 & n25919;
  assign n25923 = pi1154 & ~n25921;
  assign n25924 = ~n25922 & n25923;
  assign n25925 = ~pi618 & n25919;
  assign n25926 = pi618 & n25828;
  assign n25927 = ~pi1154 & ~n25926;
  assign n25928 = ~n25925 & n25927;
  assign n25929 = ~n25924 & ~n25928;
  assign n25930 = pi781 & ~n25929;
  assign n25931 = ~n25920 & ~n25930;
  assign n25932 = ~pi789 & ~n25931;
  assign n25933 = ~pi619 & n25828;
  assign n25934 = pi619 & n25931;
  assign n25935 = pi1159 & ~n25933;
  assign n25936 = ~n25934 & n25935;
  assign n25937 = ~pi619 & n25931;
  assign n25938 = pi619 & n25828;
  assign n25939 = ~pi1159 & ~n25938;
  assign n25940 = ~n25937 & n25939;
  assign n25941 = ~n25936 & ~n25940;
  assign n25942 = pi789 & ~n25941;
  assign n25943 = ~n25932 & ~n25942;
  assign n25944 = ~n15832 & n25943;
  assign n25945 = n15832 & n25828;
  assign n25946 = ~n25944 & ~n25945;
  assign n25947 = ~n15925 & ~n25946;
  assign n25948 = n15925 & n25828;
  assign n25949 = ~n25947 & ~n25948;
  assign n25950 = ~n15960 & ~n25949;
  assign n25951 = n15960 & n25828;
  assign n25952 = ~n25950 & ~n25951;
  assign n25953 = pi644 & ~n25952;
  assign n25954 = ~pi644 & n25828;
  assign n25955 = ~pi715 & ~n25954;
  assign n25956 = ~n25953 & n25955;
  assign n25957 = pi1160 & ~n25956;
  assign n25958 = ~n25889 & n25957;
  assign n25959 = pi644 & n25887;
  assign n25960 = ~pi715 & ~n25959;
  assign n25961 = ~pi644 & ~n25952;
  assign n25962 = pi644 & n25828;
  assign n25963 = pi715 & ~n25962;
  assign n25964 = ~n25961 & n25963;
  assign n25965 = ~pi1160 & ~n25964;
  assign n25966 = ~n25960 & n25965;
  assign n25967 = ~n25958 & ~n25966;
  assign n25968 = pi790 & ~n25967;
  assign n25969 = n15957 & n25878;
  assign n25970 = pi630 & n25883;
  assign n25971 = n19478 & n25949;
  assign n25972 = ~n25969 & ~n25970;
  assign n25973 = ~n25971 & n25972;
  assign n25974 = pi787 & ~n25973;
  assign n25975 = ~n16633 & n25946;
  assign n25976 = ~pi629 & n25868;
  assign n25977 = pi629 & n25872;
  assign n25978 = ~n25976 & ~n25977;
  assign n25979 = ~n25975 & n25978;
  assign n25980 = pi792 & ~n25979;
  assign n25981 = n15828 & ~n25860;
  assign n25982 = ~pi626 & ~n25828;
  assign n25983 = pi626 & ~n25943;
  assign n25984 = n15756 & ~n25982;
  assign n25985 = ~n25983 & n25984;
  assign n25986 = pi626 & ~n25828;
  assign n25987 = ~pi626 & ~n25943;
  assign n25988 = n15757 & ~n25986;
  assign n25989 = ~n25987 & n25988;
  assign n25990 = ~n25981 & ~n25985;
  assign n25991 = ~n25989 & n25990;
  assign n25992 = pi788 & ~n25991;
  assign n25993 = pi618 & ~n25855;
  assign n25994 = pi609 & n25852;
  assign n25995 = ~n25830 & ~n25903;
  assign n25996 = ~pi756 & ~n16808;
  assign n25997 = n18669 & ~n25996;
  assign n25998 = ~pi182 & ~n25997;
  assign n25999 = ~n16921 & ~n25677;
  assign n26000 = pi182 & ~n25999;
  assign n26001 = n6081 & n26000;
  assign n26002 = pi38 & ~n26001;
  assign n26003 = ~n25998 & n26002;
  assign n26004 = ~pi182 & ~n16647;
  assign n26005 = pi182 & ~n17397;
  assign n26006 = ~pi756 & ~n26004;
  assign n26007 = ~n26005 & n26006;
  assign n26008 = ~pi182 & n16653;
  assign n26009 = pi182 & n16657;
  assign n26010 = pi756 & ~n26008;
  assign n26011 = ~n26009 & n26010;
  assign n26012 = ~pi39 & ~n26007;
  assign n26013 = ~n26011 & n26012;
  assign n26014 = pi182 & n16825;
  assign n26015 = ~pi182 & ~n16747;
  assign n26016 = pi756 & ~n26014;
  assign n26017 = ~n26015 & n26016;
  assign n26018 = ~pi182 & n16877;
  assign n26019 = pi182 & n16913;
  assign n26020 = ~pi756 & ~n26018;
  assign n26021 = ~n26019 & n26020;
  assign n26022 = pi39 & ~n26021;
  assign n26023 = ~n26017 & n26022;
  assign n26024 = ~pi38 & ~n26013;
  assign n26025 = ~n26023 & n26024;
  assign n26026 = ~pi734 & ~n26003;
  assign n26027 = ~n26025 & n26026;
  assign n26028 = ~n25995 & ~n26027;
  assign n26029 = ~n25890 & ~n26028;
  assign n26030 = ~pi625 & n26029;
  assign n26031 = pi625 & n25904;
  assign n26032 = ~pi1153 & ~n26031;
  assign n26033 = ~n26030 & n26032;
  assign n26034 = ~pi608 & ~n25845;
  assign n26035 = ~n26033 & n26034;
  assign n26036 = ~pi625 & n25904;
  assign n26037 = pi625 & n26029;
  assign n26038 = pi1153 & ~n26036;
  assign n26039 = ~n26037 & n26038;
  assign n26040 = pi608 & ~n25849;
  assign n26041 = ~n26039 & n26040;
  assign n26042 = ~n26035 & ~n26041;
  assign n26043 = pi778 & ~n26042;
  assign n26044 = ~pi778 & n26029;
  assign n26045 = ~n26043 & ~n26044;
  assign n26046 = ~pi609 & ~n26045;
  assign n26047 = ~pi1155 & ~n25994;
  assign n26048 = ~n26046 & n26047;
  assign n26049 = ~pi660 & ~n25912;
  assign n26050 = ~n26048 & n26049;
  assign n26051 = ~pi609 & n25852;
  assign n26052 = pi609 & ~n26045;
  assign n26053 = pi1155 & ~n26051;
  assign n26054 = ~n26052 & n26053;
  assign n26055 = pi660 & ~n25916;
  assign n26056 = ~n26054 & n26055;
  assign n26057 = ~n26050 & ~n26056;
  assign n26058 = pi785 & ~n26057;
  assign n26059 = ~pi785 & ~n26045;
  assign n26060 = ~n26058 & ~n26059;
  assign n26061 = ~pi618 & ~n26060;
  assign n26062 = ~pi1154 & ~n25993;
  assign n26063 = ~n26061 & n26062;
  assign n26064 = ~pi627 & ~n25924;
  assign n26065 = ~n26063 & n26064;
  assign n26066 = ~pi618 & ~n25855;
  assign n26067 = pi618 & ~n26060;
  assign n26068 = pi1154 & ~n26066;
  assign n26069 = ~n26067 & n26068;
  assign n26070 = pi627 & ~n25928;
  assign n26071 = ~n26069 & n26070;
  assign n26072 = ~n26065 & ~n26071;
  assign n26073 = pi781 & ~n26072;
  assign n26074 = ~pi781 & ~n26060;
  assign n26075 = ~n26073 & ~n26074;
  assign n26076 = ~pi789 & n26075;
  assign n26077 = ~pi619 & n25857;
  assign n26078 = pi619 & ~n26075;
  assign n26079 = pi1159 & ~n26077;
  assign n26080 = ~n26078 & n26079;
  assign n26081 = pi648 & ~n25940;
  assign n26082 = ~n26080 & n26081;
  assign n26083 = ~pi619 & ~n26075;
  assign n26084 = pi619 & n25857;
  assign n26085 = ~pi1159 & ~n26084;
  assign n26086 = ~n26083 & n26085;
  assign n26087 = ~pi648 & ~n25936;
  assign n26088 = ~n26086 & n26087;
  assign n26089 = pi789 & ~n26082;
  assign n26090 = ~n26088 & n26089;
  assign n26091 = n15833 & ~n26076;
  assign n26092 = ~n26090 & n26091;
  assign n26093 = ~n16644 & ~n25992;
  assign n26094 = ~n26092 & n26093;
  assign n26095 = ~n25980 & ~n26094;
  assign n26096 = n18841 & ~n26095;
  assign n26097 = pi644 & ~n25956;
  assign n26098 = ~n25965 & ~n26097;
  assign n26099 = ~n22949 & ~n26098;
  assign n26100 = pi790 & ~n26099;
  assign n26101 = ~n25974 & ~n26096;
  assign n26102 = ~n26100 & n26101;
  assign n26103 = ~n25968 & ~n26102;
  assign n26104 = ~po1038 & ~n26103;
  assign n26105 = ~pi832 & ~n25827;
  assign n26106 = ~n26104 & n26105;
  assign po339 = ~n25826 & ~n26106;
  assign n26108 = ~pi183 & ~n2923;
  assign n26109 = ~pi725 & n15726;
  assign n26110 = ~n26108 & ~n26109;
  assign n26111 = ~pi778 & ~n26110;
  assign n26112 = ~pi625 & n26109;
  assign n26113 = ~n26110 & ~n26112;
  assign n26114 = pi1153 & ~n26113;
  assign n26115 = ~pi1153 & ~n26108;
  assign n26116 = ~n26112 & n26115;
  assign n26117 = pi778 & ~n26116;
  assign n26118 = ~n26114 & n26117;
  assign n26119 = ~n26111 & ~n26118;
  assign n26120 = ~n15742 & ~n26119;
  assign n26121 = ~n15748 & n26120;
  assign n26122 = ~n15754 & n26121;
  assign n26123 = ~n15760 & n26122;
  assign n26124 = ~n15766 & n26123;
  assign n26125 = n19394 & n26124;
  assign n26126 = ~n19394 & n26108;
  assign n26127 = ~n26125 & ~n26126;
  assign n26128 = ~n15959 & n26127;
  assign n26129 = n15925 & n26108;
  assign n26130 = ~pi755 & n15781;
  assign n26131 = ~n26108 & ~n26130;
  assign n26132 = ~n15778 & ~n26131;
  assign n26133 = ~pi785 & ~n26132;
  assign n26134 = n16585 & n26130;
  assign n26135 = n26132 & ~n26134;
  assign n26136 = pi1155 & ~n26135;
  assign n26137 = ~pi1155 & ~n26108;
  assign n26138 = ~n26134 & n26137;
  assign n26139 = ~n26136 & ~n26138;
  assign n26140 = pi785 & ~n26139;
  assign n26141 = ~n26133 & ~n26140;
  assign n26142 = ~pi781 & ~n26141;
  assign n26143 = ~n15797 & n26141;
  assign n26144 = pi1154 & ~n26143;
  assign n26145 = ~n15800 & n26141;
  assign n26146 = ~pi1154 & ~n26145;
  assign n26147 = ~n26144 & ~n26146;
  assign n26148 = pi781 & ~n26147;
  assign n26149 = ~n26142 & ~n26148;
  assign n26150 = ~n21915 & n26149;
  assign n26151 = ~n15832 & ~n26150;
  assign n26152 = n15832 & ~n26108;
  assign n26153 = ~n26151 & ~n26152;
  assign n26154 = ~n15925 & n26153;
  assign n26155 = n19478 & ~n26129;
  assign n26156 = ~n26154 & n26155;
  assign n26157 = ~n26128 & ~n26156;
  assign n26158 = pi787 & ~n26157;
  assign n26159 = n15763 & n26153;
  assign n26160 = n15772 & n26123;
  assign n26161 = ~pi629 & ~n26160;
  assign n26162 = ~n26159 & n26161;
  assign n26163 = n15762 & n26153;
  assign n26164 = n15909 & n26123;
  assign n26165 = pi629 & ~n26164;
  assign n26166 = ~n26163 & n26165;
  assign n26167 = pi792 & ~n26162;
  assign n26168 = ~n26166 & n26167;
  assign n26169 = ~n21932 & n26149;
  assign n26170 = pi648 & ~n26169;
  assign n26171 = n21935 & ~n26121;
  assign n26172 = ~n26170 & ~n26171;
  assign n26173 = ~pi1159 & ~n26172;
  assign n26174 = ~pi619 & ~n26121;
  assign n26175 = pi648 & ~n26174;
  assign n26176 = n21942 & n26149;
  assign n26177 = pi1159 & ~n26175;
  assign n26178 = ~n26176 & n26177;
  assign n26179 = ~n26173 & ~n26178;
  assign n26180 = pi789 & ~n26179;
  assign n26181 = pi609 & ~n26119;
  assign n26182 = ~n15780 & ~n26110;
  assign n26183 = pi625 & n26182;
  assign n26184 = n26131 & ~n26182;
  assign n26185 = ~n26183 & ~n26184;
  assign n26186 = n26115 & ~n26185;
  assign n26187 = ~pi608 & ~n26114;
  assign n26188 = ~n26186 & n26187;
  assign n26189 = pi1153 & n26131;
  assign n26190 = ~n26183 & n26189;
  assign n26191 = pi608 & ~n26116;
  assign n26192 = ~n26190 & n26191;
  assign n26193 = ~n26188 & ~n26192;
  assign n26194 = pi778 & ~n26193;
  assign n26195 = ~pi778 & ~n26184;
  assign n26196 = ~n26194 & ~n26195;
  assign n26197 = ~pi609 & ~n26196;
  assign n26198 = ~pi1155 & ~n26181;
  assign n26199 = ~n26197 & n26198;
  assign n26200 = ~pi660 & ~n26136;
  assign n26201 = ~n26199 & n26200;
  assign n26202 = ~pi609 & ~n26119;
  assign n26203 = pi609 & ~n26196;
  assign n26204 = pi1155 & ~n26202;
  assign n26205 = ~n26203 & n26204;
  assign n26206 = pi660 & ~n26138;
  assign n26207 = ~n26205 & n26206;
  assign n26208 = ~n26201 & ~n26207;
  assign n26209 = pi785 & ~n26208;
  assign n26210 = ~pi785 & ~n26196;
  assign n26211 = ~n26209 & ~n26210;
  assign n26212 = ~pi781 & n26211;
  assign n26213 = pi618 & n26120;
  assign n26214 = ~pi618 & ~n26211;
  assign n26215 = ~pi1154 & ~n26213;
  assign n26216 = ~n26214 & n26215;
  assign n26217 = ~pi627 & ~n26144;
  assign n26218 = ~n26216 & n26217;
  assign n26219 = ~pi618 & n26120;
  assign n26220 = pi618 & ~n26211;
  assign n26221 = pi1154 & ~n26219;
  assign n26222 = ~n26220 & n26221;
  assign n26223 = pi627 & ~n26146;
  assign n26224 = ~n26222 & n26223;
  assign n26225 = pi781 & ~n26218;
  assign n26226 = ~n26224 & n26225;
  assign n26227 = ~n26180 & ~n26212;
  assign n26228 = ~n26226 & n26227;
  assign n26229 = n18969 & n26179;
  assign n26230 = ~n26228 & ~n26229;
  assign n26231 = n15833 & ~n26230;
  assign n26232 = n15828 & n26122;
  assign n26233 = ~pi626 & ~n26108;
  assign n26234 = pi626 & ~n26150;
  assign n26235 = n15756 & ~n26233;
  assign n26236 = ~n26234 & n26235;
  assign n26237 = pi626 & ~n26108;
  assign n26238 = ~pi626 & ~n26150;
  assign n26239 = n15757 & ~n26237;
  assign n26240 = ~n26238 & n26239;
  assign n26241 = ~n26232 & ~n26236;
  assign n26242 = ~n26240 & n26241;
  assign n26243 = pi788 & ~n26242;
  assign n26244 = ~n26231 & ~n26243;
  assign n26245 = ~n16644 & ~n26244;
  assign n26246 = n18841 & ~n26168;
  assign n26247 = ~n26245 & n26246;
  assign n26248 = ~n26158 & ~n26247;
  assign n26249 = ~pi790 & n26248;
  assign n26250 = pi787 & ~n26127;
  assign n26251 = ~pi787 & n26124;
  assign n26252 = ~n26250 & ~n26251;
  assign n26253 = ~pi644 & ~n26252;
  assign n26254 = pi644 & n26248;
  assign n26255 = pi715 & ~n26253;
  assign n26256 = ~n26254 & n26255;
  assign n26257 = ~n19771 & n26108;
  assign n26258 = ~n15960 & n26154;
  assign n26259 = ~n26257 & ~n26258;
  assign n26260 = pi644 & ~n26259;
  assign n26261 = ~pi644 & n26108;
  assign n26262 = ~pi715 & ~n26261;
  assign n26263 = ~n26260 & n26262;
  assign n26264 = pi1160 & ~n26263;
  assign n26265 = ~n26256 & n26264;
  assign n26266 = ~pi644 & ~n26259;
  assign n26267 = pi644 & n26108;
  assign n26268 = pi715 & ~n26267;
  assign n26269 = ~n26266 & n26268;
  assign n26270 = pi644 & ~n26252;
  assign n26271 = ~pi644 & n26248;
  assign n26272 = ~pi715 & ~n26270;
  assign n26273 = ~n26271 & n26272;
  assign n26274 = ~pi1160 & ~n26269;
  assign n26275 = ~n26273 & n26274;
  assign n26276 = ~n26265 & ~n26275;
  assign n26277 = pi790 & ~n26276;
  assign n26278 = pi832 & ~n26249;
  assign n26279 = ~n26277 & n26278;
  assign n26280 = ~pi183 & po1038;
  assign n26281 = ~pi183 & ~n16219;
  assign n26282 = n15747 & ~n26281;
  assign n26283 = ~pi725 & n9829;
  assign n26284 = n26281 & ~n26283;
  assign n26285 = ~pi183 & ~n16228;
  assign n26286 = n16227 & ~n26285;
  assign n26287 = ~pi183 & ~n17276;
  assign n26288 = ~pi38 & ~pi183;
  assign n26289 = n19350 & ~n26288;
  assign n26290 = ~n26287 & ~n26289;
  assign n26291 = ~pi725 & ~n26286;
  assign n26292 = ~n26290 & n26291;
  assign n26293 = ~n26284 & ~n26292;
  assign n26294 = ~pi778 & n26293;
  assign n26295 = ~pi625 & n26281;
  assign n26296 = pi625 & ~n26293;
  assign n26297 = pi1153 & ~n26295;
  assign n26298 = ~n26296 & n26297;
  assign n26299 = pi625 & n26281;
  assign n26300 = ~pi625 & ~n26293;
  assign n26301 = ~pi1153 & ~n26299;
  assign n26302 = ~n26300 & n26301;
  assign n26303 = ~n26298 & ~n26302;
  assign n26304 = pi778 & ~n26303;
  assign n26305 = ~n26294 & ~n26304;
  assign n26306 = ~n15741 & n26305;
  assign n26307 = n15741 & n26281;
  assign n26308 = ~n26306 & ~n26307;
  assign n26309 = ~n15747 & n26308;
  assign n26310 = ~n26282 & ~n26309;
  assign n26311 = ~n15753 & n26310;
  assign n26312 = n15753 & n26281;
  assign n26313 = ~n26311 & ~n26312;
  assign n26314 = ~n15759 & ~n26313;
  assign n26315 = n15759 & n26281;
  assign n26316 = ~n26314 & ~n26315;
  assign n26317 = ~pi792 & n26316;
  assign n26318 = ~pi628 & n26281;
  assign n26319 = pi628 & ~n26316;
  assign n26320 = pi1156 & ~n26318;
  assign n26321 = ~n26319 & n26320;
  assign n26322 = pi628 & n26281;
  assign n26323 = ~pi628 & ~n26316;
  assign n26324 = ~pi1156 & ~n26322;
  assign n26325 = ~n26323 & n26324;
  assign n26326 = ~n26321 & ~n26325;
  assign n26327 = pi792 & ~n26326;
  assign n26328 = ~n26317 & ~n26327;
  assign n26329 = pi647 & n26328;
  assign n26330 = ~pi647 & n26281;
  assign n26331 = ~n26329 & ~n26330;
  assign n26332 = pi1157 & n26331;
  assign n26333 = ~pi647 & n26328;
  assign n26334 = pi647 & n26281;
  assign n26335 = ~pi1157 & ~n26334;
  assign n26336 = ~n26333 & n26335;
  assign n26337 = ~n26332 & ~n26336;
  assign n26338 = pi787 & ~n26337;
  assign n26339 = ~pi787 & ~n26328;
  assign n26340 = ~n26338 & ~n26339;
  assign n26341 = ~pi644 & n26340;
  assign n26342 = pi715 & ~n26341;
  assign n26343 = pi183 & ~n9829;
  assign n26344 = ~pi183 & n16514;
  assign n26345 = pi183 & ~n16565;
  assign n26346 = ~pi755 & ~n26344;
  assign n26347 = ~n26345 & n26346;
  assign n26348 = ~pi183 & pi755;
  assign n26349 = ~n16214 & n26348;
  assign n26350 = ~n26347 & ~n26349;
  assign n26351 = ~pi38 & ~n26350;
  assign n26352 = ~pi755 & n16570;
  assign n26353 = ~n26285 & ~n26352;
  assign n26354 = pi38 & ~n26353;
  assign n26355 = n9829 & ~n26354;
  assign n26356 = ~n26351 & n26355;
  assign n26357 = ~n26343 & ~n26356;
  assign n26358 = ~n15777 & ~n26357;
  assign n26359 = n15777 & ~n26281;
  assign n26360 = ~n26358 & ~n26359;
  assign n26361 = ~pi785 & ~n26360;
  assign n26362 = ~n15786 & ~n26281;
  assign n26363 = pi609 & n26358;
  assign n26364 = ~n26362 & ~n26363;
  assign n26365 = pi1155 & ~n26364;
  assign n26366 = ~n16585 & ~n26281;
  assign n26367 = ~pi609 & n26358;
  assign n26368 = ~n26366 & ~n26367;
  assign n26369 = ~pi1155 & ~n26368;
  assign n26370 = ~n26365 & ~n26369;
  assign n26371 = pi785 & ~n26370;
  assign n26372 = ~n26361 & ~n26371;
  assign n26373 = ~pi781 & ~n26372;
  assign n26374 = ~pi618 & n26281;
  assign n26375 = pi618 & n26372;
  assign n26376 = pi1154 & ~n26374;
  assign n26377 = ~n26375 & n26376;
  assign n26378 = ~pi618 & n26372;
  assign n26379 = pi618 & n26281;
  assign n26380 = ~pi1154 & ~n26379;
  assign n26381 = ~n26378 & n26380;
  assign n26382 = ~n26377 & ~n26381;
  assign n26383 = pi781 & ~n26382;
  assign n26384 = ~n26373 & ~n26383;
  assign n26385 = ~pi789 & ~n26384;
  assign n26386 = ~pi619 & n26281;
  assign n26387 = pi619 & n26384;
  assign n26388 = pi1159 & ~n26386;
  assign n26389 = ~n26387 & n26388;
  assign n26390 = ~pi619 & n26384;
  assign n26391 = pi619 & n26281;
  assign n26392 = ~pi1159 & ~n26391;
  assign n26393 = ~n26390 & n26392;
  assign n26394 = ~n26389 & ~n26393;
  assign n26395 = pi789 & ~n26394;
  assign n26396 = ~n26385 & ~n26395;
  assign n26397 = ~n15832 & n26396;
  assign n26398 = n15832 & n26281;
  assign n26399 = ~n26397 & ~n26398;
  assign n26400 = ~n15925 & ~n26399;
  assign n26401 = n15925 & n26281;
  assign n26402 = ~n26400 & ~n26401;
  assign n26403 = ~n15960 & ~n26402;
  assign n26404 = n15960 & n26281;
  assign n26405 = ~n26403 & ~n26404;
  assign n26406 = pi644 & ~n26405;
  assign n26407 = ~pi644 & n26281;
  assign n26408 = ~pi715 & ~n26407;
  assign n26409 = ~n26406 & n26408;
  assign n26410 = pi1160 & ~n26409;
  assign n26411 = ~n26342 & n26410;
  assign n26412 = pi644 & n26340;
  assign n26413 = ~pi715 & ~n26412;
  assign n26414 = ~pi644 & ~n26405;
  assign n26415 = pi644 & n26281;
  assign n26416 = pi715 & ~n26415;
  assign n26417 = ~n26414 & n26416;
  assign n26418 = ~pi1160 & ~n26417;
  assign n26419 = ~n26413 & n26418;
  assign n26420 = ~n26411 & ~n26419;
  assign n26421 = pi790 & ~n26420;
  assign n26422 = n15957 & n26331;
  assign n26423 = pi630 & n26336;
  assign n26424 = n19478 & n26402;
  assign n26425 = ~n26422 & ~n26423;
  assign n26426 = ~n26424 & n26425;
  assign n26427 = pi787 & ~n26426;
  assign n26428 = ~n16633 & n26399;
  assign n26429 = ~pi629 & n26321;
  assign n26430 = pi629 & n26325;
  assign n26431 = ~n26429 & ~n26430;
  assign n26432 = ~n26428 & n26431;
  assign n26433 = pi792 & ~n26432;
  assign n26434 = n15828 & ~n26313;
  assign n26435 = ~pi626 & ~n26281;
  assign n26436 = pi626 & ~n26396;
  assign n26437 = n15756 & ~n26435;
  assign n26438 = ~n26436 & n26437;
  assign n26439 = pi626 & ~n26281;
  assign n26440 = ~pi626 & ~n26396;
  assign n26441 = n15757 & ~n26439;
  assign n26442 = ~n26440 & n26441;
  assign n26443 = ~n26434 & ~n26438;
  assign n26444 = ~n26442 & n26443;
  assign n26445 = pi788 & ~n26444;
  assign n26446 = pi618 & ~n26308;
  assign n26447 = pi609 & n26305;
  assign n26448 = ~n26283 & ~n26356;
  assign n26449 = ~pi755 & ~n16808;
  assign n26450 = n18669 & ~n26449;
  assign n26451 = ~pi183 & ~n26450;
  assign n26452 = ~n16921 & ~n26130;
  assign n26453 = pi183 & ~n26452;
  assign n26454 = n6081 & n26453;
  assign n26455 = pi38 & ~n26454;
  assign n26456 = ~n26451 & n26455;
  assign n26457 = ~pi183 & ~n16647;
  assign n26458 = pi183 & ~n17397;
  assign n26459 = ~pi755 & ~n26457;
  assign n26460 = ~n26458 & n26459;
  assign n26461 = ~pi183 & n16653;
  assign n26462 = pi183 & n16657;
  assign n26463 = pi755 & ~n26461;
  assign n26464 = ~n26462 & n26463;
  assign n26465 = ~pi39 & ~n26460;
  assign n26466 = ~n26464 & n26465;
  assign n26467 = pi183 & n16825;
  assign n26468 = ~pi183 & ~n16747;
  assign n26469 = pi755 & ~n26467;
  assign n26470 = ~n26468 & n26469;
  assign n26471 = ~pi183 & n16877;
  assign n26472 = pi183 & n16913;
  assign n26473 = ~pi755 & ~n26471;
  assign n26474 = ~n26472 & n26473;
  assign n26475 = pi39 & ~n26474;
  assign n26476 = ~n26470 & n26475;
  assign n26477 = ~pi38 & ~n26466;
  assign n26478 = ~n26476 & n26477;
  assign n26479 = ~pi725 & ~n26456;
  assign n26480 = ~n26478 & n26479;
  assign n26481 = ~n26448 & ~n26480;
  assign n26482 = ~n26343 & ~n26481;
  assign n26483 = ~pi625 & n26482;
  assign n26484 = pi625 & n26357;
  assign n26485 = ~pi1153 & ~n26484;
  assign n26486 = ~n26483 & n26485;
  assign n26487 = ~pi608 & ~n26298;
  assign n26488 = ~n26486 & n26487;
  assign n26489 = ~pi625 & n26357;
  assign n26490 = pi625 & n26482;
  assign n26491 = pi1153 & ~n26489;
  assign n26492 = ~n26490 & n26491;
  assign n26493 = pi608 & ~n26302;
  assign n26494 = ~n26492 & n26493;
  assign n26495 = ~n26488 & ~n26494;
  assign n26496 = pi778 & ~n26495;
  assign n26497 = ~pi778 & n26482;
  assign n26498 = ~n26496 & ~n26497;
  assign n26499 = ~pi609 & ~n26498;
  assign n26500 = ~pi1155 & ~n26447;
  assign n26501 = ~n26499 & n26500;
  assign n26502 = ~pi660 & ~n26365;
  assign n26503 = ~n26501 & n26502;
  assign n26504 = ~pi609 & n26305;
  assign n26505 = pi609 & ~n26498;
  assign n26506 = pi1155 & ~n26504;
  assign n26507 = ~n26505 & n26506;
  assign n26508 = pi660 & ~n26369;
  assign n26509 = ~n26507 & n26508;
  assign n26510 = ~n26503 & ~n26509;
  assign n26511 = pi785 & ~n26510;
  assign n26512 = ~pi785 & ~n26498;
  assign n26513 = ~n26511 & ~n26512;
  assign n26514 = ~pi618 & ~n26513;
  assign n26515 = ~pi1154 & ~n26446;
  assign n26516 = ~n26514 & n26515;
  assign n26517 = ~pi627 & ~n26377;
  assign n26518 = ~n26516 & n26517;
  assign n26519 = ~pi618 & ~n26308;
  assign n26520 = pi618 & ~n26513;
  assign n26521 = pi1154 & ~n26519;
  assign n26522 = ~n26520 & n26521;
  assign n26523 = pi627 & ~n26381;
  assign n26524 = ~n26522 & n26523;
  assign n26525 = ~n26518 & ~n26524;
  assign n26526 = pi781 & ~n26525;
  assign n26527 = ~pi781 & ~n26513;
  assign n26528 = ~n26526 & ~n26527;
  assign n26529 = ~pi789 & n26528;
  assign n26530 = ~pi619 & n26310;
  assign n26531 = pi619 & ~n26528;
  assign n26532 = pi1159 & ~n26530;
  assign n26533 = ~n26531 & n26532;
  assign n26534 = pi648 & ~n26393;
  assign n26535 = ~n26533 & n26534;
  assign n26536 = ~pi619 & ~n26528;
  assign n26537 = pi619 & n26310;
  assign n26538 = ~pi1159 & ~n26537;
  assign n26539 = ~n26536 & n26538;
  assign n26540 = ~pi648 & ~n26389;
  assign n26541 = ~n26539 & n26540;
  assign n26542 = pi789 & ~n26535;
  assign n26543 = ~n26541 & n26542;
  assign n26544 = n15833 & ~n26529;
  assign n26545 = ~n26543 & n26544;
  assign n26546 = ~n16644 & ~n26445;
  assign n26547 = ~n26545 & n26546;
  assign n26548 = ~n26433 & ~n26547;
  assign n26549 = n18841 & ~n26548;
  assign n26550 = pi644 & ~n26409;
  assign n26551 = ~n26418 & ~n26550;
  assign n26552 = ~n22949 & ~n26551;
  assign n26553 = pi790 & ~n26552;
  assign n26554 = ~n26427 & ~n26549;
  assign n26555 = ~n26553 & n26554;
  assign n26556 = ~n26421 & ~n26555;
  assign n26557 = ~po1038 & ~n26556;
  assign n26558 = ~pi832 & ~n26280;
  assign n26559 = ~n26557 & n26558;
  assign po340 = ~n26279 & ~n26559;
  assign n26561 = ~pi184 & ~n2923;
  assign n26562 = ~pi737 & n15726;
  assign n26563 = ~n26561 & ~n26562;
  assign n26564 = ~pi778 & ~n26563;
  assign n26565 = ~pi625 & n26562;
  assign n26566 = ~n26563 & ~n26565;
  assign n26567 = pi1153 & ~n26566;
  assign n26568 = ~pi1153 & ~n26561;
  assign n26569 = ~n26565 & n26568;
  assign n26570 = pi778 & ~n26569;
  assign n26571 = ~n26567 & n26570;
  assign n26572 = ~n26564 & ~n26571;
  assign n26573 = ~n15742 & ~n26572;
  assign n26574 = ~n15748 & n26573;
  assign n26575 = ~n15754 & n26574;
  assign n26576 = ~n15760 & n26575;
  assign n26577 = ~n15766 & n26576;
  assign n26578 = n19394 & n26577;
  assign n26579 = ~n19394 & n26561;
  assign n26580 = ~n26578 & ~n26579;
  assign n26581 = ~n15959 & n26580;
  assign n26582 = n15925 & n26561;
  assign n26583 = ~pi777 & n15781;
  assign n26584 = ~n26561 & ~n26583;
  assign n26585 = ~n15778 & ~n26584;
  assign n26586 = ~pi785 & ~n26585;
  assign n26587 = n16585 & n26583;
  assign n26588 = n26585 & ~n26587;
  assign n26589 = pi1155 & ~n26588;
  assign n26590 = ~pi1155 & ~n26561;
  assign n26591 = ~n26587 & n26590;
  assign n26592 = ~n26589 & ~n26591;
  assign n26593 = pi785 & ~n26592;
  assign n26594 = ~n26586 & ~n26593;
  assign n26595 = ~pi781 & ~n26594;
  assign n26596 = ~n15797 & n26594;
  assign n26597 = pi1154 & ~n26596;
  assign n26598 = ~n15800 & n26594;
  assign n26599 = ~pi1154 & ~n26598;
  assign n26600 = ~n26597 & ~n26599;
  assign n26601 = pi781 & ~n26600;
  assign n26602 = ~n26595 & ~n26601;
  assign n26603 = ~n21915 & n26602;
  assign n26604 = ~n15832 & ~n26603;
  assign n26605 = n15832 & ~n26561;
  assign n26606 = ~n26604 & ~n26605;
  assign n26607 = ~n15925 & n26606;
  assign n26608 = n19478 & ~n26582;
  assign n26609 = ~n26607 & n26608;
  assign n26610 = ~n26581 & ~n26609;
  assign n26611 = pi787 & ~n26610;
  assign n26612 = n15763 & n26606;
  assign n26613 = n15772 & n26576;
  assign n26614 = ~pi629 & ~n26613;
  assign n26615 = ~n26612 & n26614;
  assign n26616 = n15762 & n26606;
  assign n26617 = n15909 & n26576;
  assign n26618 = pi629 & ~n26617;
  assign n26619 = ~n26616 & n26618;
  assign n26620 = pi792 & ~n26615;
  assign n26621 = ~n26619 & n26620;
  assign n26622 = ~n21932 & n26602;
  assign n26623 = pi648 & ~n26622;
  assign n26624 = n21935 & ~n26574;
  assign n26625 = ~n26623 & ~n26624;
  assign n26626 = ~pi1159 & ~n26625;
  assign n26627 = ~pi619 & ~n26574;
  assign n26628 = pi648 & ~n26627;
  assign n26629 = n21942 & n26602;
  assign n26630 = pi1159 & ~n26628;
  assign n26631 = ~n26629 & n26630;
  assign n26632 = ~n26626 & ~n26631;
  assign n26633 = pi789 & ~n26632;
  assign n26634 = pi609 & ~n26572;
  assign n26635 = ~n15780 & ~n26563;
  assign n26636 = pi625 & n26635;
  assign n26637 = n26584 & ~n26635;
  assign n26638 = ~n26636 & ~n26637;
  assign n26639 = n26568 & ~n26638;
  assign n26640 = ~pi608 & ~n26567;
  assign n26641 = ~n26639 & n26640;
  assign n26642 = pi1153 & n26584;
  assign n26643 = ~n26636 & n26642;
  assign n26644 = pi608 & ~n26569;
  assign n26645 = ~n26643 & n26644;
  assign n26646 = ~n26641 & ~n26645;
  assign n26647 = pi778 & ~n26646;
  assign n26648 = ~pi778 & ~n26637;
  assign n26649 = ~n26647 & ~n26648;
  assign n26650 = ~pi609 & ~n26649;
  assign n26651 = ~pi1155 & ~n26634;
  assign n26652 = ~n26650 & n26651;
  assign n26653 = ~pi660 & ~n26589;
  assign n26654 = ~n26652 & n26653;
  assign n26655 = ~pi609 & ~n26572;
  assign n26656 = pi609 & ~n26649;
  assign n26657 = pi1155 & ~n26655;
  assign n26658 = ~n26656 & n26657;
  assign n26659 = pi660 & ~n26591;
  assign n26660 = ~n26658 & n26659;
  assign n26661 = ~n26654 & ~n26660;
  assign n26662 = pi785 & ~n26661;
  assign n26663 = ~pi785 & ~n26649;
  assign n26664 = ~n26662 & ~n26663;
  assign n26665 = ~pi781 & n26664;
  assign n26666 = pi618 & n26573;
  assign n26667 = ~pi618 & ~n26664;
  assign n26668 = ~pi1154 & ~n26666;
  assign n26669 = ~n26667 & n26668;
  assign n26670 = ~pi627 & ~n26597;
  assign n26671 = ~n26669 & n26670;
  assign n26672 = ~pi618 & n26573;
  assign n26673 = pi618 & ~n26664;
  assign n26674 = pi1154 & ~n26672;
  assign n26675 = ~n26673 & n26674;
  assign n26676 = pi627 & ~n26599;
  assign n26677 = ~n26675 & n26676;
  assign n26678 = pi781 & ~n26671;
  assign n26679 = ~n26677 & n26678;
  assign n26680 = ~n26633 & ~n26665;
  assign n26681 = ~n26679 & n26680;
  assign n26682 = n18969 & n26632;
  assign n26683 = ~n26681 & ~n26682;
  assign n26684 = n15833 & ~n26683;
  assign n26685 = n15828 & n26575;
  assign n26686 = ~pi626 & ~n26561;
  assign n26687 = pi626 & ~n26603;
  assign n26688 = n15756 & ~n26686;
  assign n26689 = ~n26687 & n26688;
  assign n26690 = pi626 & ~n26561;
  assign n26691 = ~pi626 & ~n26603;
  assign n26692 = n15757 & ~n26690;
  assign n26693 = ~n26691 & n26692;
  assign n26694 = ~n26685 & ~n26689;
  assign n26695 = ~n26693 & n26694;
  assign n26696 = pi788 & ~n26695;
  assign n26697 = ~n26684 & ~n26696;
  assign n26698 = ~n16644 & ~n26697;
  assign n26699 = n18841 & ~n26621;
  assign n26700 = ~n26698 & n26699;
  assign n26701 = ~n26611 & ~n26700;
  assign n26702 = ~pi790 & n26701;
  assign n26703 = pi787 & ~n26580;
  assign n26704 = ~pi787 & n26577;
  assign n26705 = ~n26703 & ~n26704;
  assign n26706 = ~pi644 & ~n26705;
  assign n26707 = pi644 & n26701;
  assign n26708 = pi715 & ~n26706;
  assign n26709 = ~n26707 & n26708;
  assign n26710 = ~n19771 & n26561;
  assign n26711 = ~n15960 & n26607;
  assign n26712 = ~n26710 & ~n26711;
  assign n26713 = pi644 & ~n26712;
  assign n26714 = ~pi644 & n26561;
  assign n26715 = ~pi715 & ~n26714;
  assign n26716 = ~n26713 & n26715;
  assign n26717 = pi1160 & ~n26716;
  assign n26718 = ~n26709 & n26717;
  assign n26719 = ~pi644 & ~n26712;
  assign n26720 = pi644 & n26561;
  assign n26721 = pi715 & ~n26720;
  assign n26722 = ~n26719 & n26721;
  assign n26723 = pi644 & ~n26705;
  assign n26724 = ~pi644 & n26701;
  assign n26725 = ~pi715 & ~n26723;
  assign n26726 = ~n26724 & n26725;
  assign n26727 = ~pi1160 & ~n26722;
  assign n26728 = ~n26726 & n26727;
  assign n26729 = ~n26718 & ~n26728;
  assign n26730 = pi790 & ~n26729;
  assign n26731 = pi832 & ~n26702;
  assign n26732 = ~n26730 & n26731;
  assign n26733 = ~pi184 & po1038;
  assign n26734 = ~pi184 & ~n16219;
  assign n26735 = n15747 & ~n26734;
  assign n26736 = ~pi737 & n9829;
  assign n26737 = n26734 & ~n26736;
  assign n26738 = ~pi184 & ~n16228;
  assign n26739 = n16227 & ~n26738;
  assign n26740 = ~pi184 & ~n17276;
  assign n26741 = ~pi38 & ~pi184;
  assign n26742 = n19350 & ~n26741;
  assign n26743 = ~n26740 & ~n26742;
  assign n26744 = ~pi737 & ~n26739;
  assign n26745 = ~n26743 & n26744;
  assign n26746 = ~n26737 & ~n26745;
  assign n26747 = ~pi778 & n26746;
  assign n26748 = ~pi625 & n26734;
  assign n26749 = pi625 & ~n26746;
  assign n26750 = pi1153 & ~n26748;
  assign n26751 = ~n26749 & n26750;
  assign n26752 = pi625 & n26734;
  assign n26753 = ~pi625 & ~n26746;
  assign n26754 = ~pi1153 & ~n26752;
  assign n26755 = ~n26753 & n26754;
  assign n26756 = ~n26751 & ~n26755;
  assign n26757 = pi778 & ~n26756;
  assign n26758 = ~n26747 & ~n26757;
  assign n26759 = ~n15741 & n26758;
  assign n26760 = n15741 & n26734;
  assign n26761 = ~n26759 & ~n26760;
  assign n26762 = ~n15747 & n26761;
  assign n26763 = ~n26735 & ~n26762;
  assign n26764 = ~n15753 & n26763;
  assign n26765 = n15753 & n26734;
  assign n26766 = ~n26764 & ~n26765;
  assign n26767 = ~n15759 & ~n26766;
  assign n26768 = n15759 & n26734;
  assign n26769 = ~n26767 & ~n26768;
  assign n26770 = ~pi792 & n26769;
  assign n26771 = ~pi628 & n26734;
  assign n26772 = pi628 & ~n26769;
  assign n26773 = pi1156 & ~n26771;
  assign n26774 = ~n26772 & n26773;
  assign n26775 = pi628 & n26734;
  assign n26776 = ~pi628 & ~n26769;
  assign n26777 = ~pi1156 & ~n26775;
  assign n26778 = ~n26776 & n26777;
  assign n26779 = ~n26774 & ~n26778;
  assign n26780 = pi792 & ~n26779;
  assign n26781 = ~n26770 & ~n26780;
  assign n26782 = pi647 & n26781;
  assign n26783 = ~pi647 & n26734;
  assign n26784 = ~n26782 & ~n26783;
  assign n26785 = pi1157 & n26784;
  assign n26786 = ~pi647 & n26781;
  assign n26787 = pi647 & n26734;
  assign n26788 = ~pi1157 & ~n26787;
  assign n26789 = ~n26786 & n26788;
  assign n26790 = ~n26785 & ~n26789;
  assign n26791 = pi787 & ~n26790;
  assign n26792 = ~pi787 & ~n26781;
  assign n26793 = ~n26791 & ~n26792;
  assign n26794 = ~pi644 & n26793;
  assign n26795 = pi715 & ~n26794;
  assign n26796 = pi184 & ~n9829;
  assign n26797 = ~pi184 & n16514;
  assign n26798 = pi184 & ~n16565;
  assign n26799 = ~pi777 & ~n26797;
  assign n26800 = ~n26798 & n26799;
  assign n26801 = ~pi184 & pi777;
  assign n26802 = ~n16214 & n26801;
  assign n26803 = ~n26800 & ~n26802;
  assign n26804 = ~pi38 & ~n26803;
  assign n26805 = ~pi777 & n16570;
  assign n26806 = ~n26738 & ~n26805;
  assign n26807 = pi38 & ~n26806;
  assign n26808 = n9829 & ~n26807;
  assign n26809 = ~n26804 & n26808;
  assign n26810 = ~n26796 & ~n26809;
  assign n26811 = ~n15777 & ~n26810;
  assign n26812 = n15777 & ~n26734;
  assign n26813 = ~n26811 & ~n26812;
  assign n26814 = ~pi785 & ~n26813;
  assign n26815 = ~n15786 & ~n26734;
  assign n26816 = pi609 & n26811;
  assign n26817 = ~n26815 & ~n26816;
  assign n26818 = pi1155 & ~n26817;
  assign n26819 = ~n16585 & ~n26734;
  assign n26820 = ~pi609 & n26811;
  assign n26821 = ~n26819 & ~n26820;
  assign n26822 = ~pi1155 & ~n26821;
  assign n26823 = ~n26818 & ~n26822;
  assign n26824 = pi785 & ~n26823;
  assign n26825 = ~n26814 & ~n26824;
  assign n26826 = ~pi781 & ~n26825;
  assign n26827 = ~pi618 & n26734;
  assign n26828 = pi618 & n26825;
  assign n26829 = pi1154 & ~n26827;
  assign n26830 = ~n26828 & n26829;
  assign n26831 = ~pi618 & n26825;
  assign n26832 = pi618 & n26734;
  assign n26833 = ~pi1154 & ~n26832;
  assign n26834 = ~n26831 & n26833;
  assign n26835 = ~n26830 & ~n26834;
  assign n26836 = pi781 & ~n26835;
  assign n26837 = ~n26826 & ~n26836;
  assign n26838 = ~pi789 & ~n26837;
  assign n26839 = ~pi619 & n26734;
  assign n26840 = pi619 & n26837;
  assign n26841 = pi1159 & ~n26839;
  assign n26842 = ~n26840 & n26841;
  assign n26843 = ~pi619 & n26837;
  assign n26844 = pi619 & n26734;
  assign n26845 = ~pi1159 & ~n26844;
  assign n26846 = ~n26843 & n26845;
  assign n26847 = ~n26842 & ~n26846;
  assign n26848 = pi789 & ~n26847;
  assign n26849 = ~n26838 & ~n26848;
  assign n26850 = ~n15832 & n26849;
  assign n26851 = n15832 & n26734;
  assign n26852 = ~n26850 & ~n26851;
  assign n26853 = ~n15925 & ~n26852;
  assign n26854 = n15925 & n26734;
  assign n26855 = ~n26853 & ~n26854;
  assign n26856 = ~n15960 & ~n26855;
  assign n26857 = n15960 & n26734;
  assign n26858 = ~n26856 & ~n26857;
  assign n26859 = pi644 & ~n26858;
  assign n26860 = ~pi644 & n26734;
  assign n26861 = ~pi715 & ~n26860;
  assign n26862 = ~n26859 & n26861;
  assign n26863 = pi1160 & ~n26862;
  assign n26864 = ~n26795 & n26863;
  assign n26865 = pi644 & n26793;
  assign n26866 = ~pi715 & ~n26865;
  assign n26867 = ~pi644 & ~n26858;
  assign n26868 = pi644 & n26734;
  assign n26869 = pi715 & ~n26868;
  assign n26870 = ~n26867 & n26869;
  assign n26871 = ~pi1160 & ~n26870;
  assign n26872 = ~n26866 & n26871;
  assign n26873 = ~n26864 & ~n26872;
  assign n26874 = pi790 & ~n26873;
  assign n26875 = n15957 & n26784;
  assign n26876 = pi630 & n26789;
  assign n26877 = n19478 & n26855;
  assign n26878 = ~n26875 & ~n26876;
  assign n26879 = ~n26877 & n26878;
  assign n26880 = pi787 & ~n26879;
  assign n26881 = ~n16633 & n26852;
  assign n26882 = ~pi629 & n26774;
  assign n26883 = pi629 & n26778;
  assign n26884 = ~n26882 & ~n26883;
  assign n26885 = ~n26881 & n26884;
  assign n26886 = pi792 & ~n26885;
  assign n26887 = n15828 & ~n26766;
  assign n26888 = ~pi626 & ~n26734;
  assign n26889 = pi626 & ~n26849;
  assign n26890 = n15756 & ~n26888;
  assign n26891 = ~n26889 & n26890;
  assign n26892 = pi626 & ~n26734;
  assign n26893 = ~pi626 & ~n26849;
  assign n26894 = n15757 & ~n26892;
  assign n26895 = ~n26893 & n26894;
  assign n26896 = ~n26887 & ~n26891;
  assign n26897 = ~n26895 & n26896;
  assign n26898 = pi788 & ~n26897;
  assign n26899 = pi618 & ~n26761;
  assign n26900 = pi609 & n26758;
  assign n26901 = ~n26736 & ~n26809;
  assign n26902 = ~pi777 & ~n16808;
  assign n26903 = n18669 & ~n26902;
  assign n26904 = ~pi184 & ~n26903;
  assign n26905 = ~n16921 & ~n26583;
  assign n26906 = pi184 & ~n26905;
  assign n26907 = n6081 & n26906;
  assign n26908 = pi38 & ~n26907;
  assign n26909 = ~n26904 & n26908;
  assign n26910 = ~pi184 & ~n16647;
  assign n26911 = pi184 & ~n17397;
  assign n26912 = ~pi777 & ~n26910;
  assign n26913 = ~n26911 & n26912;
  assign n26914 = ~pi184 & n16653;
  assign n26915 = pi184 & n16657;
  assign n26916 = pi777 & ~n26914;
  assign n26917 = ~n26915 & n26916;
  assign n26918 = ~pi39 & ~n26913;
  assign n26919 = ~n26917 & n26918;
  assign n26920 = pi184 & n16825;
  assign n26921 = ~pi184 & ~n16747;
  assign n26922 = pi777 & ~n26920;
  assign n26923 = ~n26921 & n26922;
  assign n26924 = ~pi184 & n16877;
  assign n26925 = pi184 & n16913;
  assign n26926 = ~pi777 & ~n26924;
  assign n26927 = ~n26925 & n26926;
  assign n26928 = pi39 & ~n26927;
  assign n26929 = ~n26923 & n26928;
  assign n26930 = ~pi38 & ~n26919;
  assign n26931 = ~n26929 & n26930;
  assign n26932 = ~pi737 & ~n26909;
  assign n26933 = ~n26931 & n26932;
  assign n26934 = ~n26901 & ~n26933;
  assign n26935 = ~n26796 & ~n26934;
  assign n26936 = ~pi625 & n26935;
  assign n26937 = pi625 & n26810;
  assign n26938 = ~pi1153 & ~n26937;
  assign n26939 = ~n26936 & n26938;
  assign n26940 = ~pi608 & ~n26751;
  assign n26941 = ~n26939 & n26940;
  assign n26942 = ~pi625 & n26810;
  assign n26943 = pi625 & n26935;
  assign n26944 = pi1153 & ~n26942;
  assign n26945 = ~n26943 & n26944;
  assign n26946 = pi608 & ~n26755;
  assign n26947 = ~n26945 & n26946;
  assign n26948 = ~n26941 & ~n26947;
  assign n26949 = pi778 & ~n26948;
  assign n26950 = ~pi778 & n26935;
  assign n26951 = ~n26949 & ~n26950;
  assign n26952 = ~pi609 & ~n26951;
  assign n26953 = ~pi1155 & ~n26900;
  assign n26954 = ~n26952 & n26953;
  assign n26955 = ~pi660 & ~n26818;
  assign n26956 = ~n26954 & n26955;
  assign n26957 = ~pi609 & n26758;
  assign n26958 = pi609 & ~n26951;
  assign n26959 = pi1155 & ~n26957;
  assign n26960 = ~n26958 & n26959;
  assign n26961 = pi660 & ~n26822;
  assign n26962 = ~n26960 & n26961;
  assign n26963 = ~n26956 & ~n26962;
  assign n26964 = pi785 & ~n26963;
  assign n26965 = ~pi785 & ~n26951;
  assign n26966 = ~n26964 & ~n26965;
  assign n26967 = ~pi618 & ~n26966;
  assign n26968 = ~pi1154 & ~n26899;
  assign n26969 = ~n26967 & n26968;
  assign n26970 = ~pi627 & ~n26830;
  assign n26971 = ~n26969 & n26970;
  assign n26972 = ~pi618 & ~n26761;
  assign n26973 = pi618 & ~n26966;
  assign n26974 = pi1154 & ~n26972;
  assign n26975 = ~n26973 & n26974;
  assign n26976 = pi627 & ~n26834;
  assign n26977 = ~n26975 & n26976;
  assign n26978 = ~n26971 & ~n26977;
  assign n26979 = pi781 & ~n26978;
  assign n26980 = ~pi781 & ~n26966;
  assign n26981 = ~n26979 & ~n26980;
  assign n26982 = ~pi789 & n26981;
  assign n26983 = ~pi619 & n26763;
  assign n26984 = pi619 & ~n26981;
  assign n26985 = pi1159 & ~n26983;
  assign n26986 = ~n26984 & n26985;
  assign n26987 = pi648 & ~n26846;
  assign n26988 = ~n26986 & n26987;
  assign n26989 = ~pi619 & ~n26981;
  assign n26990 = pi619 & n26763;
  assign n26991 = ~pi1159 & ~n26990;
  assign n26992 = ~n26989 & n26991;
  assign n26993 = ~pi648 & ~n26842;
  assign n26994 = ~n26992 & n26993;
  assign n26995 = pi789 & ~n26988;
  assign n26996 = ~n26994 & n26995;
  assign n26997 = n15833 & ~n26982;
  assign n26998 = ~n26996 & n26997;
  assign n26999 = ~n16644 & ~n26898;
  assign n27000 = ~n26998 & n26999;
  assign n27001 = ~n26886 & ~n27000;
  assign n27002 = n18841 & ~n27001;
  assign n27003 = pi644 & ~n26862;
  assign n27004 = ~n26871 & ~n27003;
  assign n27005 = ~n22949 & ~n27004;
  assign n27006 = pi790 & ~n27005;
  assign n27007 = ~n26880 & ~n27002;
  assign n27008 = ~n27006 & n27007;
  assign n27009 = ~n26874 & ~n27008;
  assign n27010 = ~po1038 & ~n27009;
  assign n27011 = ~pi832 & ~n26733;
  assign n27012 = ~n27010 & n27011;
  assign po341 = ~n26732 & ~n27012;
  assign n27014 = ~pi185 & ~n2923;
  assign n27015 = ~pi701 & n15726;
  assign n27016 = ~n27014 & ~n27015;
  assign n27017 = ~pi778 & ~n27016;
  assign n27018 = ~pi625 & n27015;
  assign n27019 = ~n27016 & ~n27018;
  assign n27020 = pi1153 & ~n27019;
  assign n27021 = ~pi1153 & ~n27014;
  assign n27022 = ~n27018 & n27021;
  assign n27023 = pi778 & ~n27022;
  assign n27024 = ~n27020 & n27023;
  assign n27025 = ~n27017 & ~n27024;
  assign n27026 = ~n15742 & ~n27025;
  assign n27027 = ~n15748 & n27026;
  assign n27028 = ~n15754 & n27027;
  assign n27029 = ~n15760 & n27028;
  assign n27030 = ~n15766 & n27029;
  assign n27031 = n19394 & n27030;
  assign n27032 = ~n19394 & n27014;
  assign n27033 = ~n27031 & ~n27032;
  assign n27034 = ~n15959 & n27033;
  assign n27035 = n15925 & n27014;
  assign n27036 = ~pi751 & n15781;
  assign n27037 = ~n27014 & ~n27036;
  assign n27038 = ~n15778 & ~n27037;
  assign n27039 = ~pi785 & ~n27038;
  assign n27040 = n16585 & n27036;
  assign n27041 = n27038 & ~n27040;
  assign n27042 = pi1155 & ~n27041;
  assign n27043 = ~pi1155 & ~n27014;
  assign n27044 = ~n27040 & n27043;
  assign n27045 = ~n27042 & ~n27044;
  assign n27046 = pi785 & ~n27045;
  assign n27047 = ~n27039 & ~n27046;
  assign n27048 = ~pi781 & ~n27047;
  assign n27049 = ~n15797 & n27047;
  assign n27050 = pi1154 & ~n27049;
  assign n27051 = ~n15800 & n27047;
  assign n27052 = ~pi1154 & ~n27051;
  assign n27053 = ~n27050 & ~n27052;
  assign n27054 = pi781 & ~n27053;
  assign n27055 = ~n27048 & ~n27054;
  assign n27056 = ~n21915 & n27055;
  assign n27057 = ~n15832 & ~n27056;
  assign n27058 = n15832 & ~n27014;
  assign n27059 = ~n27057 & ~n27058;
  assign n27060 = ~n15925 & n27059;
  assign n27061 = n19478 & ~n27035;
  assign n27062 = ~n27060 & n27061;
  assign n27063 = ~n27034 & ~n27062;
  assign n27064 = pi787 & ~n27063;
  assign n27065 = n15763 & n27059;
  assign n27066 = n15772 & n27029;
  assign n27067 = ~pi629 & ~n27066;
  assign n27068 = ~n27065 & n27067;
  assign n27069 = n15762 & n27059;
  assign n27070 = n15909 & n27029;
  assign n27071 = pi629 & ~n27070;
  assign n27072 = ~n27069 & n27071;
  assign n27073 = pi792 & ~n27068;
  assign n27074 = ~n27072 & n27073;
  assign n27075 = ~n21932 & n27055;
  assign n27076 = pi648 & ~n27075;
  assign n27077 = n21935 & ~n27027;
  assign n27078 = ~n27076 & ~n27077;
  assign n27079 = ~pi1159 & ~n27078;
  assign n27080 = ~pi619 & ~n27027;
  assign n27081 = pi648 & ~n27080;
  assign n27082 = n21942 & n27055;
  assign n27083 = pi1159 & ~n27081;
  assign n27084 = ~n27082 & n27083;
  assign n27085 = ~n27079 & ~n27084;
  assign n27086 = pi789 & ~n27085;
  assign n27087 = pi609 & ~n27025;
  assign n27088 = ~n15780 & ~n27016;
  assign n27089 = pi625 & n27088;
  assign n27090 = n27037 & ~n27088;
  assign n27091 = ~n27089 & ~n27090;
  assign n27092 = n27021 & ~n27091;
  assign n27093 = ~pi608 & ~n27020;
  assign n27094 = ~n27092 & n27093;
  assign n27095 = pi1153 & n27037;
  assign n27096 = ~n27089 & n27095;
  assign n27097 = pi608 & ~n27022;
  assign n27098 = ~n27096 & n27097;
  assign n27099 = ~n27094 & ~n27098;
  assign n27100 = pi778 & ~n27099;
  assign n27101 = ~pi778 & ~n27090;
  assign n27102 = ~n27100 & ~n27101;
  assign n27103 = ~pi609 & ~n27102;
  assign n27104 = ~pi1155 & ~n27087;
  assign n27105 = ~n27103 & n27104;
  assign n27106 = ~pi660 & ~n27042;
  assign n27107 = ~n27105 & n27106;
  assign n27108 = ~pi609 & ~n27025;
  assign n27109 = pi609 & ~n27102;
  assign n27110 = pi1155 & ~n27108;
  assign n27111 = ~n27109 & n27110;
  assign n27112 = pi660 & ~n27044;
  assign n27113 = ~n27111 & n27112;
  assign n27114 = ~n27107 & ~n27113;
  assign n27115 = pi785 & ~n27114;
  assign n27116 = ~pi785 & ~n27102;
  assign n27117 = ~n27115 & ~n27116;
  assign n27118 = ~pi781 & n27117;
  assign n27119 = pi618 & n27026;
  assign n27120 = ~pi618 & ~n27117;
  assign n27121 = ~pi1154 & ~n27119;
  assign n27122 = ~n27120 & n27121;
  assign n27123 = ~pi627 & ~n27050;
  assign n27124 = ~n27122 & n27123;
  assign n27125 = ~pi618 & n27026;
  assign n27126 = pi618 & ~n27117;
  assign n27127 = pi1154 & ~n27125;
  assign n27128 = ~n27126 & n27127;
  assign n27129 = pi627 & ~n27052;
  assign n27130 = ~n27128 & n27129;
  assign n27131 = pi781 & ~n27124;
  assign n27132 = ~n27130 & n27131;
  assign n27133 = ~n27086 & ~n27118;
  assign n27134 = ~n27132 & n27133;
  assign n27135 = n18969 & n27085;
  assign n27136 = ~n27134 & ~n27135;
  assign n27137 = n15833 & ~n27136;
  assign n27138 = n15828 & n27028;
  assign n27139 = ~pi626 & ~n27014;
  assign n27140 = pi626 & ~n27056;
  assign n27141 = n15756 & ~n27139;
  assign n27142 = ~n27140 & n27141;
  assign n27143 = pi626 & ~n27014;
  assign n27144 = ~pi626 & ~n27056;
  assign n27145 = n15757 & ~n27143;
  assign n27146 = ~n27144 & n27145;
  assign n27147 = ~n27138 & ~n27142;
  assign n27148 = ~n27146 & n27147;
  assign n27149 = pi788 & ~n27148;
  assign n27150 = ~n27137 & ~n27149;
  assign n27151 = ~n16644 & ~n27150;
  assign n27152 = n18841 & ~n27074;
  assign n27153 = ~n27151 & n27152;
  assign n27154 = ~n27064 & ~n27153;
  assign n27155 = ~pi790 & n27154;
  assign n27156 = pi787 & ~n27033;
  assign n27157 = ~pi787 & n27030;
  assign n27158 = ~n27156 & ~n27157;
  assign n27159 = ~pi644 & ~n27158;
  assign n27160 = pi644 & n27154;
  assign n27161 = pi715 & ~n27159;
  assign n27162 = ~n27160 & n27161;
  assign n27163 = ~n19771 & n27014;
  assign n27164 = ~n15960 & n27060;
  assign n27165 = ~n27163 & ~n27164;
  assign n27166 = pi644 & ~n27165;
  assign n27167 = ~pi644 & n27014;
  assign n27168 = ~pi715 & ~n27167;
  assign n27169 = ~n27166 & n27168;
  assign n27170 = pi1160 & ~n27169;
  assign n27171 = ~n27162 & n27170;
  assign n27172 = ~pi644 & ~n27165;
  assign n27173 = pi644 & n27014;
  assign n27174 = pi715 & ~n27173;
  assign n27175 = ~n27172 & n27174;
  assign n27176 = pi644 & ~n27158;
  assign n27177 = ~pi644 & n27154;
  assign n27178 = ~pi715 & ~n27176;
  assign n27179 = ~n27177 & n27178;
  assign n27180 = ~pi1160 & ~n27175;
  assign n27181 = ~n27179 & n27180;
  assign n27182 = ~n27171 & ~n27181;
  assign n27183 = pi790 & ~n27182;
  assign n27184 = pi832 & ~n27155;
  assign n27185 = ~n27183 & n27184;
  assign n27186 = ~pi185 & po1038;
  assign n27187 = ~pi185 & ~n16219;
  assign n27188 = n15747 & ~n27187;
  assign n27189 = ~pi701 & n9829;
  assign n27190 = n27187 & ~n27189;
  assign n27191 = ~pi185 & ~n16228;
  assign n27192 = n16227 & ~n27191;
  assign n27193 = ~pi185 & ~n17276;
  assign n27194 = ~pi38 & ~pi185;
  assign n27195 = n19350 & ~n27194;
  assign n27196 = ~n27193 & ~n27195;
  assign n27197 = ~pi701 & ~n27192;
  assign n27198 = ~n27196 & n27197;
  assign n27199 = ~n27190 & ~n27198;
  assign n27200 = ~pi778 & n27199;
  assign n27201 = ~pi625 & n27187;
  assign n27202 = pi625 & ~n27199;
  assign n27203 = pi1153 & ~n27201;
  assign n27204 = ~n27202 & n27203;
  assign n27205 = pi625 & n27187;
  assign n27206 = ~pi625 & ~n27199;
  assign n27207 = ~pi1153 & ~n27205;
  assign n27208 = ~n27206 & n27207;
  assign n27209 = ~n27204 & ~n27208;
  assign n27210 = pi778 & ~n27209;
  assign n27211 = ~n27200 & ~n27210;
  assign n27212 = ~n15741 & n27211;
  assign n27213 = n15741 & n27187;
  assign n27214 = ~n27212 & ~n27213;
  assign n27215 = ~n15747 & n27214;
  assign n27216 = ~n27188 & ~n27215;
  assign n27217 = ~n15753 & n27216;
  assign n27218 = n15753 & n27187;
  assign n27219 = ~n27217 & ~n27218;
  assign n27220 = ~n15759 & ~n27219;
  assign n27221 = n15759 & n27187;
  assign n27222 = ~n27220 & ~n27221;
  assign n27223 = ~pi792 & n27222;
  assign n27224 = ~pi628 & n27187;
  assign n27225 = pi628 & ~n27222;
  assign n27226 = pi1156 & ~n27224;
  assign n27227 = ~n27225 & n27226;
  assign n27228 = pi628 & n27187;
  assign n27229 = ~pi628 & ~n27222;
  assign n27230 = ~pi1156 & ~n27228;
  assign n27231 = ~n27229 & n27230;
  assign n27232 = ~n27227 & ~n27231;
  assign n27233 = pi792 & ~n27232;
  assign n27234 = ~n27223 & ~n27233;
  assign n27235 = n19394 & n27234;
  assign n27236 = ~n19394 & n27187;
  assign n27237 = ~n27235 & ~n27236;
  assign n27238 = pi787 & ~n27237;
  assign n27239 = ~pi787 & n27234;
  assign n27240 = ~n27238 & ~n27239;
  assign n27241 = ~pi644 & ~n27240;
  assign n27242 = pi715 & ~n27241;
  assign n27243 = pi185 & ~n9829;
  assign n27244 = ~pi751 & n16570;
  assign n27245 = ~n27191 & ~n27244;
  assign n27246 = pi38 & ~n27245;
  assign n27247 = pi751 & n16212;
  assign n27248 = pi185 & ~n16563;
  assign n27249 = ~n27247 & ~n27248;
  assign n27250 = pi39 & ~n27249;
  assign n27251 = ~pi185 & ~pi751;
  assign n27252 = n16514 & n27251;
  assign n27253 = pi185 & pi751;
  assign n27254 = pi185 & ~n16526;
  assign n27255 = ~n20168 & ~n27254;
  assign n27256 = ~pi39 & ~n27255;
  assign n27257 = ~pi38 & ~n27253;
  assign n27258 = ~n27256 & n27257;
  assign n27259 = ~n27252 & n27258;
  assign n27260 = ~n27250 & n27259;
  assign n27261 = n9829 & ~n27246;
  assign n27262 = ~n27260 & n27261;
  assign n27263 = ~n27243 & ~n27262;
  assign n27264 = ~n15777 & ~n27263;
  assign n27265 = n15777 & ~n27187;
  assign n27266 = ~n27264 & ~n27265;
  assign n27267 = ~pi785 & ~n27266;
  assign n27268 = ~n15786 & ~n27187;
  assign n27269 = pi609 & n27264;
  assign n27270 = ~n27268 & ~n27269;
  assign n27271 = pi1155 & ~n27270;
  assign n27272 = ~n16585 & ~n27187;
  assign n27273 = ~pi609 & n27264;
  assign n27274 = ~n27272 & ~n27273;
  assign n27275 = ~pi1155 & ~n27274;
  assign n27276 = ~n27271 & ~n27275;
  assign n27277 = pi785 & ~n27276;
  assign n27278 = ~n27267 & ~n27277;
  assign n27279 = ~pi781 & ~n27278;
  assign n27280 = ~pi618 & n27187;
  assign n27281 = pi618 & n27278;
  assign n27282 = pi1154 & ~n27280;
  assign n27283 = ~n27281 & n27282;
  assign n27284 = ~pi618 & n27278;
  assign n27285 = pi618 & n27187;
  assign n27286 = ~pi1154 & ~n27285;
  assign n27287 = ~n27284 & n27286;
  assign n27288 = ~n27283 & ~n27287;
  assign n27289 = pi781 & ~n27288;
  assign n27290 = ~n27279 & ~n27289;
  assign n27291 = ~pi789 & ~n27290;
  assign n27292 = ~pi619 & n27187;
  assign n27293 = pi619 & n27290;
  assign n27294 = pi1159 & ~n27292;
  assign n27295 = ~n27293 & n27294;
  assign n27296 = ~pi619 & n27290;
  assign n27297 = pi619 & n27187;
  assign n27298 = ~pi1159 & ~n27297;
  assign n27299 = ~n27296 & n27298;
  assign n27300 = ~n27295 & ~n27299;
  assign n27301 = pi789 & ~n27300;
  assign n27302 = ~n27291 & ~n27301;
  assign n27303 = ~n15832 & n27302;
  assign n27304 = n15832 & n27187;
  assign n27305 = ~n27303 & ~n27304;
  assign n27306 = ~n15925 & ~n27305;
  assign n27307 = n15925 & n27187;
  assign n27308 = ~n27306 & ~n27307;
  assign n27309 = ~n15960 & ~n27308;
  assign n27310 = n15960 & n27187;
  assign n27311 = ~n27309 & ~n27310;
  assign n27312 = pi644 & ~n27311;
  assign n27313 = ~pi644 & n27187;
  assign n27314 = ~pi715 & ~n27313;
  assign n27315 = ~n27312 & n27314;
  assign n27316 = pi1160 & ~n27315;
  assign n27317 = ~n27242 & n27316;
  assign n27318 = pi644 & ~n27240;
  assign n27319 = ~pi715 & ~n27318;
  assign n27320 = ~pi644 & ~n27311;
  assign n27321 = pi644 & n27187;
  assign n27322 = pi715 & ~n27321;
  assign n27323 = ~n27320 & n27322;
  assign n27324 = ~pi1160 & ~n27323;
  assign n27325 = ~n27319 & n27324;
  assign n27326 = ~n27317 & ~n27325;
  assign n27327 = pi790 & ~n27326;
  assign n27328 = n19478 & n27308;
  assign n27329 = ~n15959 & n27237;
  assign n27330 = ~n27328 & ~n27329;
  assign n27331 = pi787 & ~n27330;
  assign n27332 = ~n16633 & n27305;
  assign n27333 = ~pi629 & n27227;
  assign n27334 = pi629 & n27231;
  assign n27335 = ~n27333 & ~n27334;
  assign n27336 = ~n27332 & n27335;
  assign n27337 = pi792 & ~n27336;
  assign n27338 = n15828 & ~n27219;
  assign n27339 = ~pi626 & ~n27187;
  assign n27340 = pi626 & ~n27302;
  assign n27341 = n15756 & ~n27339;
  assign n27342 = ~n27340 & n27341;
  assign n27343 = pi626 & ~n27187;
  assign n27344 = ~pi626 & ~n27302;
  assign n27345 = n15757 & ~n27343;
  assign n27346 = ~n27344 & n27345;
  assign n27347 = ~n27338 & ~n27342;
  assign n27348 = ~n27346 & n27347;
  assign n27349 = pi788 & ~n27348;
  assign n27350 = pi618 & ~n27214;
  assign n27351 = pi609 & n27211;
  assign n27352 = ~n27189 & ~n27262;
  assign n27353 = ~pi751 & ~n16808;
  assign n27354 = n18669 & ~n27353;
  assign n27355 = ~pi185 & ~n27354;
  assign n27356 = ~n16921 & ~n27036;
  assign n27357 = pi185 & ~n27356;
  assign n27358 = n6081 & n27357;
  assign n27359 = pi38 & ~n27358;
  assign n27360 = ~n27355 & n27359;
  assign n27361 = ~pi185 & ~n16647;
  assign n27362 = pi185 & ~n17397;
  assign n27363 = ~pi751 & ~n27361;
  assign n27364 = ~n27362 & n27363;
  assign n27365 = ~pi185 & n16653;
  assign n27366 = pi185 & n16657;
  assign n27367 = pi751 & ~n27365;
  assign n27368 = ~n27366 & n27367;
  assign n27369 = ~pi39 & ~n27364;
  assign n27370 = ~n27368 & n27369;
  assign n27371 = pi185 & n16825;
  assign n27372 = ~pi185 & ~n16747;
  assign n27373 = pi751 & ~n27371;
  assign n27374 = ~n27372 & n27373;
  assign n27375 = ~pi185 & n16877;
  assign n27376 = pi185 & n16913;
  assign n27377 = ~pi751 & ~n27375;
  assign n27378 = ~n27376 & n27377;
  assign n27379 = pi39 & ~n27378;
  assign n27380 = ~n27374 & n27379;
  assign n27381 = ~pi38 & ~n27370;
  assign n27382 = ~n27380 & n27381;
  assign n27383 = ~pi701 & ~n27360;
  assign n27384 = ~n27382 & n27383;
  assign n27385 = ~n27352 & ~n27384;
  assign n27386 = ~n27243 & ~n27385;
  assign n27387 = ~pi625 & n27386;
  assign n27388 = pi625 & n27263;
  assign n27389 = ~pi1153 & ~n27388;
  assign n27390 = ~n27387 & n27389;
  assign n27391 = ~pi608 & ~n27204;
  assign n27392 = ~n27390 & n27391;
  assign n27393 = ~pi625 & n27263;
  assign n27394 = pi625 & n27386;
  assign n27395 = pi1153 & ~n27393;
  assign n27396 = ~n27394 & n27395;
  assign n27397 = pi608 & ~n27208;
  assign n27398 = ~n27396 & n27397;
  assign n27399 = ~n27392 & ~n27398;
  assign n27400 = pi778 & ~n27399;
  assign n27401 = ~pi778 & n27386;
  assign n27402 = ~n27400 & ~n27401;
  assign n27403 = ~pi609 & ~n27402;
  assign n27404 = ~pi1155 & ~n27351;
  assign n27405 = ~n27403 & n27404;
  assign n27406 = ~pi660 & ~n27271;
  assign n27407 = ~n27405 & n27406;
  assign n27408 = ~pi609 & n27211;
  assign n27409 = pi609 & ~n27402;
  assign n27410 = pi1155 & ~n27408;
  assign n27411 = ~n27409 & n27410;
  assign n27412 = pi660 & ~n27275;
  assign n27413 = ~n27411 & n27412;
  assign n27414 = ~n27407 & ~n27413;
  assign n27415 = pi785 & ~n27414;
  assign n27416 = ~pi785 & ~n27402;
  assign n27417 = ~n27415 & ~n27416;
  assign n27418 = ~pi618 & ~n27417;
  assign n27419 = ~pi1154 & ~n27350;
  assign n27420 = ~n27418 & n27419;
  assign n27421 = ~pi627 & ~n27283;
  assign n27422 = ~n27420 & n27421;
  assign n27423 = ~pi618 & ~n27214;
  assign n27424 = pi618 & ~n27417;
  assign n27425 = pi1154 & ~n27423;
  assign n27426 = ~n27424 & n27425;
  assign n27427 = pi627 & ~n27287;
  assign n27428 = ~n27426 & n27427;
  assign n27429 = ~n27422 & ~n27428;
  assign n27430 = pi781 & ~n27429;
  assign n27431 = ~pi781 & ~n27417;
  assign n27432 = ~n27430 & ~n27431;
  assign n27433 = ~pi789 & n27432;
  assign n27434 = ~pi619 & n27216;
  assign n27435 = pi619 & ~n27432;
  assign n27436 = pi1159 & ~n27434;
  assign n27437 = ~n27435 & n27436;
  assign n27438 = pi648 & ~n27299;
  assign n27439 = ~n27437 & n27438;
  assign n27440 = ~pi619 & ~n27432;
  assign n27441 = pi619 & n27216;
  assign n27442 = ~pi1159 & ~n27441;
  assign n27443 = ~n27440 & n27442;
  assign n27444 = ~pi648 & ~n27295;
  assign n27445 = ~n27443 & n27444;
  assign n27446 = pi789 & ~n27439;
  assign n27447 = ~n27445 & n27446;
  assign n27448 = n15833 & ~n27433;
  assign n27449 = ~n27447 & n27448;
  assign n27450 = ~n16644 & ~n27349;
  assign n27451 = ~n27449 & n27450;
  assign n27452 = ~n27337 & ~n27451;
  assign n27453 = n18841 & ~n27452;
  assign n27454 = pi644 & ~n27315;
  assign n27455 = ~n27324 & ~n27454;
  assign n27456 = ~n22949 & ~n27455;
  assign n27457 = pi790 & ~n27456;
  assign n27458 = ~n27331 & ~n27457;
  assign n27459 = ~n27453 & n27458;
  assign n27460 = ~n27327 & ~n27459;
  assign n27461 = ~po1038 & ~n27460;
  assign n27462 = ~pi832 & ~n27186;
  assign n27463 = ~n27461 & n27462;
  assign po342 = ~n27185 & ~n27463;
  assign n27465 = ~pi186 & ~n2923;
  assign n27466 = pi703 & n15726;
  assign n27467 = ~n27465 & ~n27466;
  assign n27468 = ~pi778 & n27467;
  assign n27469 = ~pi625 & n27466;
  assign n27470 = ~n27467 & ~n27469;
  assign n27471 = pi1153 & ~n27470;
  assign n27472 = ~pi1153 & ~n27465;
  assign n27473 = ~n27469 & n27472;
  assign n27474 = ~n27471 & ~n27473;
  assign n27475 = pi778 & ~n27474;
  assign n27476 = ~n27468 & ~n27475;
  assign n27477 = ~n15742 & n27476;
  assign n27478 = ~n15748 & n27477;
  assign n27479 = ~n15754 & n27478;
  assign n27480 = ~n15760 & n27479;
  assign n27481 = ~n15766 & n27480;
  assign n27482 = n19394 & n27481;
  assign n27483 = ~n19394 & n27465;
  assign n27484 = ~n27482 & ~n27483;
  assign n27485 = ~n15959 & n27484;
  assign n27486 = n15925 & n27465;
  assign n27487 = ~pi752 & n15781;
  assign n27488 = ~n27465 & ~n27487;
  assign n27489 = ~n15778 & ~n27488;
  assign n27490 = ~pi785 & ~n27489;
  assign n27491 = ~n15787 & ~n27488;
  assign n27492 = pi1155 & ~n27491;
  assign n27493 = ~n15790 & n27489;
  assign n27494 = ~pi1155 & ~n27493;
  assign n27495 = ~n27492 & ~n27494;
  assign n27496 = pi785 & ~n27495;
  assign n27497 = ~n27490 & ~n27496;
  assign n27498 = ~pi781 & ~n27497;
  assign n27499 = ~n15797 & n27497;
  assign n27500 = pi1154 & ~n27499;
  assign n27501 = ~n15800 & n27497;
  assign n27502 = ~pi1154 & ~n27501;
  assign n27503 = ~n27500 & ~n27502;
  assign n27504 = pi781 & ~n27503;
  assign n27505 = ~n27498 & ~n27504;
  assign n27506 = ~pi789 & ~n27505;
  assign n27507 = ~pi619 & n27465;
  assign n27508 = pi619 & n27505;
  assign n27509 = pi1159 & ~n27507;
  assign n27510 = ~n27508 & n27509;
  assign n27511 = ~pi619 & n27505;
  assign n27512 = pi619 & n27465;
  assign n27513 = ~pi1159 & ~n27512;
  assign n27514 = ~n27511 & n27513;
  assign n27515 = ~n27510 & ~n27514;
  assign n27516 = pi789 & ~n27515;
  assign n27517 = ~n27506 & ~n27516;
  assign n27518 = ~n15832 & ~n27517;
  assign n27519 = n15832 & ~n27465;
  assign n27520 = ~n27518 & ~n27519;
  assign n27521 = ~n15925 & n27520;
  assign n27522 = n19478 & ~n27486;
  assign n27523 = ~n27521 & n27522;
  assign n27524 = ~n27485 & ~n27523;
  assign n27525 = pi787 & ~n27524;
  assign n27526 = n15828 & n27479;
  assign n27527 = ~pi626 & ~n27465;
  assign n27528 = pi626 & ~n27517;
  assign n27529 = n15756 & ~n27527;
  assign n27530 = ~n27528 & n27529;
  assign n27531 = pi626 & ~n27465;
  assign n27532 = ~pi626 & ~n27517;
  assign n27533 = n15757 & ~n27531;
  assign n27534 = ~n27532 & n27533;
  assign n27535 = ~n27526 & ~n27530;
  assign n27536 = ~n27534 & n27535;
  assign n27537 = pi788 & ~n27536;
  assign n27538 = pi618 & n27477;
  assign n27539 = pi609 & n27476;
  assign n27540 = ~n15780 & ~n27467;
  assign n27541 = pi625 & n27540;
  assign n27542 = n27488 & ~n27540;
  assign n27543 = ~n27541 & ~n27542;
  assign n27544 = n27472 & ~n27543;
  assign n27545 = ~pi608 & ~n27471;
  assign n27546 = ~n27544 & n27545;
  assign n27547 = pi1153 & n27488;
  assign n27548 = ~n27541 & n27547;
  assign n27549 = pi608 & ~n27473;
  assign n27550 = ~n27548 & n27549;
  assign n27551 = ~n27546 & ~n27550;
  assign n27552 = pi778 & ~n27551;
  assign n27553 = ~pi778 & ~n27542;
  assign n27554 = ~n27552 & ~n27553;
  assign n27555 = ~pi609 & ~n27554;
  assign n27556 = ~pi1155 & ~n27539;
  assign n27557 = ~n27555 & n27556;
  assign n27558 = ~pi660 & ~n27492;
  assign n27559 = ~n27557 & n27558;
  assign n27560 = ~pi609 & n27476;
  assign n27561 = pi609 & ~n27554;
  assign n27562 = pi1155 & ~n27560;
  assign n27563 = ~n27561 & n27562;
  assign n27564 = pi660 & ~n27494;
  assign n27565 = ~n27563 & n27564;
  assign n27566 = ~n27559 & ~n27565;
  assign n27567 = pi785 & ~n27566;
  assign n27568 = ~pi785 & ~n27554;
  assign n27569 = ~n27567 & ~n27568;
  assign n27570 = ~pi618 & ~n27569;
  assign n27571 = ~pi1154 & ~n27538;
  assign n27572 = ~n27570 & n27571;
  assign n27573 = ~pi627 & ~n27500;
  assign n27574 = ~n27572 & n27573;
  assign n27575 = ~pi618 & n27477;
  assign n27576 = pi618 & ~n27569;
  assign n27577 = pi1154 & ~n27575;
  assign n27578 = ~n27576 & n27577;
  assign n27579 = pi627 & ~n27502;
  assign n27580 = ~n27578 & n27579;
  assign n27581 = ~n27574 & ~n27580;
  assign n27582 = pi781 & ~n27581;
  assign n27583 = ~pi781 & ~n27569;
  assign n27584 = ~n27582 & ~n27583;
  assign n27585 = ~pi789 & n27584;
  assign n27586 = ~pi619 & n27478;
  assign n27587 = pi619 & ~n27584;
  assign n27588 = pi1159 & ~n27586;
  assign n27589 = ~n27587 & n27588;
  assign n27590 = pi648 & ~n27514;
  assign n27591 = ~n27589 & n27590;
  assign n27592 = pi619 & n27478;
  assign n27593 = ~pi619 & ~n27584;
  assign n27594 = ~pi1159 & ~n27592;
  assign n27595 = ~n27593 & n27594;
  assign n27596 = ~pi648 & ~n27510;
  assign n27597 = ~n27595 & n27596;
  assign n27598 = pi789 & ~n27591;
  assign n27599 = ~n27597 & n27598;
  assign n27600 = n15833 & ~n27585;
  assign n27601 = ~n27599 & n27600;
  assign n27602 = ~n27537 & ~n27601;
  assign n27603 = ~n16644 & ~n27602;
  assign n27604 = n15763 & n27520;
  assign n27605 = n15772 & n27480;
  assign n27606 = ~pi629 & ~n27605;
  assign n27607 = ~n27604 & n27606;
  assign n27608 = n15762 & n27520;
  assign n27609 = n15909 & n27480;
  assign n27610 = pi629 & ~n27609;
  assign n27611 = ~n27608 & n27610;
  assign n27612 = pi792 & ~n27607;
  assign n27613 = ~n27611 & n27612;
  assign n27614 = n18841 & ~n27613;
  assign n27615 = ~n27603 & n27614;
  assign n27616 = ~n27525 & ~n27615;
  assign n27617 = ~pi790 & n27616;
  assign n27618 = pi787 & ~n27484;
  assign n27619 = ~pi787 & n27481;
  assign n27620 = ~n27618 & ~n27619;
  assign n27621 = ~pi644 & ~n27620;
  assign n27622 = pi644 & n27616;
  assign n27623 = pi715 & ~n27621;
  assign n27624 = ~n27622 & n27623;
  assign n27625 = ~n19771 & n27465;
  assign n27626 = ~n15960 & n27521;
  assign n27627 = ~n27625 & ~n27626;
  assign n27628 = pi644 & ~n27627;
  assign n27629 = ~pi644 & n27465;
  assign n27630 = ~pi715 & ~n27629;
  assign n27631 = ~n27628 & n27630;
  assign n27632 = pi1160 & ~n27631;
  assign n27633 = ~n27624 & n27632;
  assign n27634 = ~pi644 & ~n27627;
  assign n27635 = pi644 & n27465;
  assign n27636 = pi715 & ~n27635;
  assign n27637 = ~n27634 & n27636;
  assign n27638 = pi644 & ~n27620;
  assign n27639 = ~pi644 & n27616;
  assign n27640 = ~pi715 & ~n27638;
  assign n27641 = ~n27639 & n27640;
  assign n27642 = ~pi1160 & ~n27637;
  assign n27643 = ~n27641 & n27642;
  assign n27644 = ~n27633 & ~n27643;
  assign n27645 = pi790 & ~n27644;
  assign n27646 = pi832 & ~n27617;
  assign n27647 = ~n27645 & n27646;
  assign n27648 = ~pi186 & po1038;
  assign n27649 = ~pi186 & ~n16219;
  assign n27650 = n15759 & ~n27649;
  assign n27651 = n15747 & ~n27649;
  assign n27652 = pi186 & ~n9829;
  assign n27653 = ~pi186 & ~n16218;
  assign n27654 = ~pi703 & n27653;
  assign n27655 = ~pi186 & ~n16228;
  assign n27656 = n16227 & ~n27655;
  assign n27657 = pi186 & n17272;
  assign n27658 = ~pi186 & ~n17276;
  assign n27659 = ~pi38 & ~n27657;
  assign n27660 = ~n27658 & n27659;
  assign n27661 = pi703 & ~n27656;
  assign n27662 = ~n27660 & n27661;
  assign n27663 = n9829 & ~n27662;
  assign n27664 = ~n27654 & n27663;
  assign n27665 = ~n27652 & ~n27664;
  assign n27666 = ~pi778 & ~n27665;
  assign n27667 = ~pi625 & n27649;
  assign n27668 = pi625 & n27665;
  assign n27669 = pi1153 & ~n27667;
  assign n27670 = ~n27668 & n27669;
  assign n27671 = ~pi625 & n27665;
  assign n27672 = pi625 & n27649;
  assign n27673 = ~pi1153 & ~n27672;
  assign n27674 = ~n27671 & n27673;
  assign n27675 = ~n27670 & ~n27674;
  assign n27676 = pi778 & ~n27675;
  assign n27677 = ~n27666 & ~n27676;
  assign n27678 = ~n15741 & n27677;
  assign n27679 = n15741 & n27649;
  assign n27680 = ~n27678 & ~n27679;
  assign n27681 = ~n15747 & n27680;
  assign n27682 = ~n27651 & ~n27681;
  assign n27683 = ~n15753 & n27682;
  assign n27684 = n15753 & n27649;
  assign n27685 = ~n27683 & ~n27684;
  assign n27686 = ~n15759 & n27685;
  assign n27687 = ~n27650 & ~n27686;
  assign n27688 = ~pi792 & ~n27687;
  assign n27689 = ~pi628 & ~n27649;
  assign n27690 = pi628 & ~n27687;
  assign n27691 = ~n27689 & ~n27690;
  assign n27692 = pi1156 & ~n27691;
  assign n27693 = ~pi628 & n27687;
  assign n27694 = pi628 & n27649;
  assign n27695 = ~pi1156 & ~n27694;
  assign n27696 = ~n27693 & n27695;
  assign n27697 = ~n27692 & ~n27696;
  assign n27698 = pi792 & ~n27697;
  assign n27699 = ~n27688 & ~n27698;
  assign n27700 = ~pi787 & ~n27699;
  assign n27701 = ~pi647 & n27649;
  assign n27702 = pi647 & n27699;
  assign n27703 = pi1157 & ~n27701;
  assign n27704 = ~n27702 & n27703;
  assign n27705 = ~pi647 & n27699;
  assign n27706 = pi647 & n27649;
  assign n27707 = ~pi1157 & ~n27706;
  assign n27708 = ~n27705 & n27707;
  assign n27709 = ~n27704 & ~n27708;
  assign n27710 = pi787 & ~n27709;
  assign n27711 = ~n27700 & ~n27710;
  assign n27712 = ~pi644 & n27711;
  assign n27713 = ~pi629 & n27692;
  assign n27714 = pi752 & ~n27653;
  assign n27715 = pi186 & ~n18599;
  assign n27716 = ~pi186 & ~pi752;
  assign n27717 = n18604 & n27716;
  assign n27718 = ~n27715 & ~n27717;
  assign n27719 = ~n18598 & ~n27718;
  assign n27720 = ~n27714 & ~n27719;
  assign n27721 = n9829 & ~n27720;
  assign n27722 = ~n27652 & ~n27721;
  assign n27723 = ~n15777 & ~n27722;
  assign n27724 = n15777 & ~n27649;
  assign n27725 = ~n27723 & ~n27724;
  assign n27726 = ~pi785 & ~n27725;
  assign n27727 = ~n15786 & ~n27649;
  assign n27728 = pi609 & n27723;
  assign n27729 = ~n27727 & ~n27728;
  assign n27730 = pi1155 & ~n27729;
  assign n27731 = ~n16585 & ~n27649;
  assign n27732 = ~pi609 & n27723;
  assign n27733 = ~n27731 & ~n27732;
  assign n27734 = ~pi1155 & ~n27733;
  assign n27735 = ~n27730 & ~n27734;
  assign n27736 = pi785 & ~n27735;
  assign n27737 = ~n27726 & ~n27736;
  assign n27738 = ~pi781 & ~n27737;
  assign n27739 = ~pi618 & n27649;
  assign n27740 = pi618 & n27737;
  assign n27741 = pi1154 & ~n27739;
  assign n27742 = ~n27740 & n27741;
  assign n27743 = ~pi618 & n27737;
  assign n27744 = pi618 & n27649;
  assign n27745 = ~pi1154 & ~n27744;
  assign n27746 = ~n27743 & n27745;
  assign n27747 = ~n27742 & ~n27746;
  assign n27748 = pi781 & ~n27747;
  assign n27749 = ~n27738 & ~n27748;
  assign n27750 = ~pi789 & ~n27749;
  assign n27751 = ~pi619 & n27649;
  assign n27752 = pi619 & n27749;
  assign n27753 = pi1159 & ~n27751;
  assign n27754 = ~n27752 & n27753;
  assign n27755 = ~pi619 & n27749;
  assign n27756 = pi619 & n27649;
  assign n27757 = ~pi1159 & ~n27756;
  assign n27758 = ~n27755 & n27757;
  assign n27759 = ~n27754 & ~n27758;
  assign n27760 = pi789 & ~n27759;
  assign n27761 = ~n27750 & ~n27760;
  assign n27762 = ~n15832 & n27761;
  assign n27763 = n15832 & n27649;
  assign n27764 = ~n27762 & ~n27763;
  assign n27765 = ~n16633 & n27764;
  assign n27766 = pi629 & n27696;
  assign n27767 = ~n27713 & ~n27766;
  assign n27768 = ~n27765 & n27767;
  assign n27769 = pi792 & ~n27768;
  assign n27770 = pi619 & n27682;
  assign n27771 = ~pi1159 & ~n27770;
  assign n27772 = ~pi648 & ~n27754;
  assign n27773 = ~n27771 & n27772;
  assign n27774 = pi618 & ~n27680;
  assign n27775 = pi609 & n27677;
  assign n27776 = ~pi703 & n27720;
  assign n27777 = ~pi186 & ~n18651;
  assign n27778 = pi186 & n18659;
  assign n27779 = ~pi752 & ~n27777;
  assign n27780 = ~n27778 & n27779;
  assign n27781 = pi186 & n18666;
  assign n27782 = ~pi186 & n18675;
  assign n27783 = pi752 & ~n18668;
  assign n27784 = ~n27781 & n27783;
  assign n27785 = ~n27782 & n27784;
  assign n27786 = pi703 & ~n27780;
  assign n27787 = ~n27785 & n27786;
  assign n27788 = n9829 & ~n27787;
  assign n27789 = ~n27776 & n27788;
  assign n27790 = ~n27652 & ~n27789;
  assign n27791 = ~pi625 & n27790;
  assign n27792 = pi625 & n27722;
  assign n27793 = ~pi1153 & ~n27792;
  assign n27794 = ~n27791 & n27793;
  assign n27795 = ~pi608 & ~n27670;
  assign n27796 = ~n27794 & n27795;
  assign n27797 = ~pi625 & n27722;
  assign n27798 = pi625 & n27790;
  assign n27799 = pi1153 & ~n27797;
  assign n27800 = ~n27798 & n27799;
  assign n27801 = pi608 & ~n27674;
  assign n27802 = ~n27800 & n27801;
  assign n27803 = ~n27796 & ~n27802;
  assign n27804 = pi778 & ~n27803;
  assign n27805 = ~pi778 & n27790;
  assign n27806 = ~n27804 & ~n27805;
  assign n27807 = ~pi609 & ~n27806;
  assign n27808 = ~pi1155 & ~n27775;
  assign n27809 = ~n27807 & n27808;
  assign n27810 = ~pi660 & ~n27730;
  assign n27811 = ~n27809 & n27810;
  assign n27812 = ~pi609 & n27677;
  assign n27813 = pi609 & ~n27806;
  assign n27814 = pi1155 & ~n27812;
  assign n27815 = ~n27813 & n27814;
  assign n27816 = pi660 & ~n27734;
  assign n27817 = ~n27815 & n27816;
  assign n27818 = ~n27811 & ~n27817;
  assign n27819 = pi785 & ~n27818;
  assign n27820 = ~pi785 & ~n27806;
  assign n27821 = ~n27819 & ~n27820;
  assign n27822 = ~pi618 & ~n27821;
  assign n27823 = ~pi1154 & ~n27774;
  assign n27824 = ~n27822 & n27823;
  assign n27825 = ~pi627 & ~n27742;
  assign n27826 = ~n27824 & n27825;
  assign n27827 = ~pi618 & ~n27680;
  assign n27828 = pi618 & ~n27821;
  assign n27829 = pi1154 & ~n27827;
  assign n27830 = ~n27828 & n27829;
  assign n27831 = pi627 & ~n27746;
  assign n27832 = ~n27830 & n27831;
  assign n27833 = ~n27826 & ~n27832;
  assign n27834 = pi781 & ~n27833;
  assign n27835 = ~pi781 & ~n27821;
  assign n27836 = ~n27834 & ~n27835;
  assign n27837 = pi619 & ~n27836;
  assign n27838 = ~pi619 & n27682;
  assign n27839 = pi1159 & ~n27838;
  assign n27840 = ~n27837 & n27839;
  assign n27841 = pi648 & ~n27758;
  assign n27842 = ~n27840 & n27841;
  assign n27843 = ~n27773 & ~n27842;
  assign n27844 = pi789 & ~n27843;
  assign n27845 = ~pi619 & n27772;
  assign n27846 = pi789 & ~n27845;
  assign n27847 = ~n27836 & ~n27846;
  assign n27848 = ~n27844 & ~n27847;
  assign n27849 = n15833 & ~n27848;
  assign n27850 = pi641 & ~n27649;
  assign n27851 = ~pi641 & n27685;
  assign n27852 = n15819 & ~n27850;
  assign n27853 = ~n27851 & n27852;
  assign n27854 = n22348 & n27761;
  assign n27855 = ~pi641 & ~n27649;
  assign n27856 = pi641 & n27685;
  assign n27857 = n15818 & ~n27855;
  assign n27858 = ~n27856 & n27857;
  assign n27859 = ~n27853 & ~n27858;
  assign n27860 = ~n27854 & n27859;
  assign n27861 = pi788 & ~n27860;
  assign n27862 = ~n16644 & ~n27861;
  assign n27863 = ~n27849 & n27862;
  assign n27864 = ~n27769 & ~n27863;
  assign n27865 = ~pi647 & n27864;
  assign n27866 = ~n15925 & ~n27764;
  assign n27867 = n15925 & n27649;
  assign n27868 = ~n27866 & ~n27867;
  assign n27869 = pi647 & ~n27868;
  assign n27870 = ~pi1157 & ~n27869;
  assign n27871 = ~n27865 & n27870;
  assign n27872 = ~pi630 & ~n27704;
  assign n27873 = ~n27871 & n27872;
  assign n27874 = ~pi647 & ~n27868;
  assign n27875 = pi647 & n27864;
  assign n27876 = pi1157 & ~n27874;
  assign n27877 = ~n27875 & n27876;
  assign n27878 = pi630 & ~n27708;
  assign n27879 = ~n27877 & n27878;
  assign n27880 = ~n27873 & ~n27879;
  assign n27881 = pi787 & ~n27880;
  assign n27882 = ~pi787 & n27864;
  assign n27883 = ~n27881 & ~n27882;
  assign n27884 = pi644 & ~n27883;
  assign n27885 = pi715 & ~n27712;
  assign n27886 = ~n27884 & n27885;
  assign n27887 = ~n15960 & ~n27868;
  assign n27888 = n15960 & n27649;
  assign n27889 = ~n27887 & ~n27888;
  assign n27890 = pi644 & ~n27889;
  assign n27891 = ~pi644 & n27649;
  assign n27892 = ~pi715 & ~n27891;
  assign n27893 = ~n27890 & n27892;
  assign n27894 = pi1160 & ~n27893;
  assign n27895 = ~n27886 & n27894;
  assign n27896 = pi644 & n27711;
  assign n27897 = ~pi715 & ~n27896;
  assign n27898 = ~pi644 & ~n27889;
  assign n27899 = pi644 & n27649;
  assign n27900 = pi715 & ~n27899;
  assign n27901 = ~n27898 & n27900;
  assign n27902 = ~pi1160 & ~n27901;
  assign n27903 = ~n27897 & n27902;
  assign n27904 = ~n27895 & ~n27903;
  assign n27905 = pi790 & ~n27904;
  assign n27906 = ~pi644 & n27902;
  assign n27907 = pi790 & ~n27906;
  assign n27908 = ~n27883 & ~n27907;
  assign n27909 = ~n27905 & ~n27908;
  assign n27910 = ~po1038 & ~n27909;
  assign n27911 = ~pi832 & ~n27648;
  assign n27912 = ~n27910 & n27911;
  assign po343 = ~n27647 & ~n27912;
  assign n27914 = ~pi187 & ~n2923;
  assign n27915 = pi726 & n15726;
  assign n27916 = ~n27914 & ~n27915;
  assign n27917 = ~pi778 & n27916;
  assign n27918 = ~pi625 & n27915;
  assign n27919 = ~n27916 & ~n27918;
  assign n27920 = pi1153 & ~n27919;
  assign n27921 = ~pi1153 & ~n27914;
  assign n27922 = ~n27918 & n27921;
  assign n27923 = ~n27920 & ~n27922;
  assign n27924 = pi778 & ~n27923;
  assign n27925 = ~n27917 & ~n27924;
  assign n27926 = ~n15742 & n27925;
  assign n27927 = ~n15748 & n27926;
  assign n27928 = ~n15754 & n27927;
  assign n27929 = ~n15760 & n27928;
  assign n27930 = ~n15766 & n27929;
  assign n27931 = n19394 & n27930;
  assign n27932 = ~n19394 & n27914;
  assign n27933 = ~n27931 & ~n27932;
  assign n27934 = ~n15959 & n27933;
  assign n27935 = n15925 & n27914;
  assign n27936 = ~pi770 & n15781;
  assign n27937 = ~n27914 & ~n27936;
  assign n27938 = ~n15778 & ~n27937;
  assign n27939 = ~pi785 & ~n27938;
  assign n27940 = ~n15787 & ~n27937;
  assign n27941 = pi1155 & ~n27940;
  assign n27942 = ~n15790 & n27938;
  assign n27943 = ~pi1155 & ~n27942;
  assign n27944 = ~n27941 & ~n27943;
  assign n27945 = pi785 & ~n27944;
  assign n27946 = ~n27939 & ~n27945;
  assign n27947 = ~pi781 & ~n27946;
  assign n27948 = ~n15797 & n27946;
  assign n27949 = pi1154 & ~n27948;
  assign n27950 = ~n15800 & n27946;
  assign n27951 = ~pi1154 & ~n27950;
  assign n27952 = ~n27949 & ~n27951;
  assign n27953 = pi781 & ~n27952;
  assign n27954 = ~n27947 & ~n27953;
  assign n27955 = ~pi789 & ~n27954;
  assign n27956 = ~pi619 & n27914;
  assign n27957 = pi619 & n27954;
  assign n27958 = pi1159 & ~n27956;
  assign n27959 = ~n27957 & n27958;
  assign n27960 = ~pi619 & n27954;
  assign n27961 = pi619 & n27914;
  assign n27962 = ~pi1159 & ~n27961;
  assign n27963 = ~n27960 & n27962;
  assign n27964 = ~n27959 & ~n27963;
  assign n27965 = pi789 & ~n27964;
  assign n27966 = ~n27955 & ~n27965;
  assign n27967 = ~n15832 & ~n27966;
  assign n27968 = n15832 & ~n27914;
  assign n27969 = ~n27967 & ~n27968;
  assign n27970 = ~n15925 & n27969;
  assign n27971 = n19478 & ~n27935;
  assign n27972 = ~n27970 & n27971;
  assign n27973 = ~n27934 & ~n27972;
  assign n27974 = pi787 & ~n27973;
  assign n27975 = n15828 & n27928;
  assign n27976 = ~pi626 & ~n27914;
  assign n27977 = pi626 & ~n27966;
  assign n27978 = n15756 & ~n27976;
  assign n27979 = ~n27977 & n27978;
  assign n27980 = pi626 & ~n27914;
  assign n27981 = ~pi626 & ~n27966;
  assign n27982 = n15757 & ~n27980;
  assign n27983 = ~n27981 & n27982;
  assign n27984 = ~n27975 & ~n27979;
  assign n27985 = ~n27983 & n27984;
  assign n27986 = pi788 & ~n27985;
  assign n27987 = pi618 & n27926;
  assign n27988 = pi609 & n27925;
  assign n27989 = ~n15780 & ~n27916;
  assign n27990 = pi625 & n27989;
  assign n27991 = n27937 & ~n27989;
  assign n27992 = ~n27990 & ~n27991;
  assign n27993 = n27921 & ~n27992;
  assign n27994 = ~pi608 & ~n27920;
  assign n27995 = ~n27993 & n27994;
  assign n27996 = pi1153 & n27937;
  assign n27997 = ~n27990 & n27996;
  assign n27998 = pi608 & ~n27922;
  assign n27999 = ~n27997 & n27998;
  assign n28000 = ~n27995 & ~n27999;
  assign n28001 = pi778 & ~n28000;
  assign n28002 = ~pi778 & ~n27991;
  assign n28003 = ~n28001 & ~n28002;
  assign n28004 = ~pi609 & ~n28003;
  assign n28005 = ~pi1155 & ~n27988;
  assign n28006 = ~n28004 & n28005;
  assign n28007 = ~pi660 & ~n27941;
  assign n28008 = ~n28006 & n28007;
  assign n28009 = ~pi609 & n27925;
  assign n28010 = pi609 & ~n28003;
  assign n28011 = pi1155 & ~n28009;
  assign n28012 = ~n28010 & n28011;
  assign n28013 = pi660 & ~n27943;
  assign n28014 = ~n28012 & n28013;
  assign n28015 = ~n28008 & ~n28014;
  assign n28016 = pi785 & ~n28015;
  assign n28017 = ~pi785 & ~n28003;
  assign n28018 = ~n28016 & ~n28017;
  assign n28019 = ~pi618 & ~n28018;
  assign n28020 = ~pi1154 & ~n27987;
  assign n28021 = ~n28019 & n28020;
  assign n28022 = ~pi627 & ~n27949;
  assign n28023 = ~n28021 & n28022;
  assign n28024 = ~pi618 & n27926;
  assign n28025 = pi618 & ~n28018;
  assign n28026 = pi1154 & ~n28024;
  assign n28027 = ~n28025 & n28026;
  assign n28028 = pi627 & ~n27951;
  assign n28029 = ~n28027 & n28028;
  assign n28030 = ~n28023 & ~n28029;
  assign n28031 = pi781 & ~n28030;
  assign n28032 = ~pi781 & ~n28018;
  assign n28033 = ~n28031 & ~n28032;
  assign n28034 = ~pi789 & n28033;
  assign n28035 = ~pi619 & n27927;
  assign n28036 = pi619 & ~n28033;
  assign n28037 = pi1159 & ~n28035;
  assign n28038 = ~n28036 & n28037;
  assign n28039 = pi648 & ~n27963;
  assign n28040 = ~n28038 & n28039;
  assign n28041 = pi619 & n27927;
  assign n28042 = ~pi619 & ~n28033;
  assign n28043 = ~pi1159 & ~n28041;
  assign n28044 = ~n28042 & n28043;
  assign n28045 = ~pi648 & ~n27959;
  assign n28046 = ~n28044 & n28045;
  assign n28047 = pi789 & ~n28040;
  assign n28048 = ~n28046 & n28047;
  assign n28049 = n15833 & ~n28034;
  assign n28050 = ~n28048 & n28049;
  assign n28051 = ~n27986 & ~n28050;
  assign n28052 = ~n16644 & ~n28051;
  assign n28053 = n15763 & n27969;
  assign n28054 = n15772 & n27929;
  assign n28055 = ~pi629 & ~n28054;
  assign n28056 = ~n28053 & n28055;
  assign n28057 = n15762 & n27969;
  assign n28058 = n15909 & n27929;
  assign n28059 = pi629 & ~n28058;
  assign n28060 = ~n28057 & n28059;
  assign n28061 = pi792 & ~n28056;
  assign n28062 = ~n28060 & n28061;
  assign n28063 = n18841 & ~n28062;
  assign n28064 = ~n28052 & n28063;
  assign n28065 = ~n27974 & ~n28064;
  assign n28066 = ~pi790 & n28065;
  assign n28067 = pi787 & ~n27933;
  assign n28068 = ~pi787 & n27930;
  assign n28069 = ~n28067 & ~n28068;
  assign n28070 = ~pi644 & ~n28069;
  assign n28071 = pi644 & n28065;
  assign n28072 = pi715 & ~n28070;
  assign n28073 = ~n28071 & n28072;
  assign n28074 = ~n19771 & n27914;
  assign n28075 = ~n15960 & n27970;
  assign n28076 = ~n28074 & ~n28075;
  assign n28077 = pi644 & ~n28076;
  assign n28078 = ~pi644 & n27914;
  assign n28079 = ~pi715 & ~n28078;
  assign n28080 = ~n28077 & n28079;
  assign n28081 = pi1160 & ~n28080;
  assign n28082 = ~n28073 & n28081;
  assign n28083 = ~pi644 & ~n28076;
  assign n28084 = pi644 & n27914;
  assign n28085 = pi715 & ~n28084;
  assign n28086 = ~n28083 & n28085;
  assign n28087 = pi644 & ~n28069;
  assign n28088 = ~pi644 & n28065;
  assign n28089 = ~pi715 & ~n28087;
  assign n28090 = ~n28088 & n28089;
  assign n28091 = ~pi1160 & ~n28086;
  assign n28092 = ~n28090 & n28091;
  assign n28093 = ~n28082 & ~n28092;
  assign n28094 = pi790 & ~n28093;
  assign n28095 = pi832 & ~n28066;
  assign n28096 = ~n28094 & n28095;
  assign n28097 = ~pi187 & po1038;
  assign n28098 = ~pi187 & ~n16219;
  assign n28099 = n15759 & ~n28098;
  assign n28100 = n15747 & ~n28098;
  assign n28101 = pi187 & ~n9829;
  assign n28102 = ~pi187 & ~n16228;
  assign n28103 = n16227 & ~n28102;
  assign n28104 = pi187 & n17272;
  assign n28105 = ~pi187 & ~n17276;
  assign n28106 = ~pi38 & ~n28104;
  assign n28107 = ~n28105 & n28106;
  assign n28108 = pi726 & ~n28103;
  assign n28109 = ~n28107 & n28108;
  assign n28110 = ~pi187 & ~pi726;
  assign n28111 = ~n16218 & n28110;
  assign n28112 = n9829 & ~n28109;
  assign n28113 = ~n28111 & n28112;
  assign n28114 = ~n28101 & ~n28113;
  assign n28115 = ~pi778 & ~n28114;
  assign n28116 = ~pi625 & n28098;
  assign n28117 = pi625 & n28114;
  assign n28118 = pi1153 & ~n28116;
  assign n28119 = ~n28117 & n28118;
  assign n28120 = ~pi625 & n28114;
  assign n28121 = pi625 & n28098;
  assign n28122 = ~pi1153 & ~n28121;
  assign n28123 = ~n28120 & n28122;
  assign n28124 = ~n28119 & ~n28123;
  assign n28125 = pi778 & ~n28124;
  assign n28126 = ~n28115 & ~n28125;
  assign n28127 = ~n15741 & n28126;
  assign n28128 = n15741 & n28098;
  assign n28129 = ~n28127 & ~n28128;
  assign n28130 = ~n15747 & n28129;
  assign n28131 = ~n28100 & ~n28130;
  assign n28132 = ~n15753 & n28131;
  assign n28133 = n15753 & n28098;
  assign n28134 = ~n28132 & ~n28133;
  assign n28135 = ~n15759 & n28134;
  assign n28136 = ~n28099 & ~n28135;
  assign n28137 = ~pi792 & ~n28136;
  assign n28138 = ~pi628 & ~n28098;
  assign n28139 = pi628 & ~n28136;
  assign n28140 = ~n28138 & ~n28139;
  assign n28141 = pi1156 & ~n28140;
  assign n28142 = ~pi628 & n28136;
  assign n28143 = pi628 & n28098;
  assign n28144 = ~pi1156 & ~n28143;
  assign n28145 = ~n28142 & n28144;
  assign n28146 = ~n28141 & ~n28145;
  assign n28147 = pi792 & ~n28146;
  assign n28148 = ~n28137 & ~n28147;
  assign n28149 = ~pi787 & ~n28148;
  assign n28150 = ~pi647 & n28098;
  assign n28151 = pi647 & n28148;
  assign n28152 = pi1157 & ~n28150;
  assign n28153 = ~n28151 & n28152;
  assign n28154 = ~pi647 & n28148;
  assign n28155 = pi647 & n28098;
  assign n28156 = ~pi1157 & ~n28155;
  assign n28157 = ~n28154 & n28156;
  assign n28158 = ~n28153 & ~n28157;
  assign n28159 = pi787 & ~n28158;
  assign n28160 = ~n28149 & ~n28159;
  assign n28161 = ~pi644 & n28160;
  assign n28162 = ~pi629 & n28141;
  assign n28163 = ~pi187 & ~pi770;
  assign n28164 = n24555 & n28163;
  assign n28165 = ~pi770 & ~n23191;
  assign n28166 = pi187 & ~n28165;
  assign n28167 = ~n28164 & ~n28166;
  assign n28168 = ~n19899 & n28167;
  assign n28169 = n9829 & ~n28168;
  assign n28170 = ~n28101 & ~n28169;
  assign n28171 = ~n15777 & ~n28170;
  assign n28172 = n15777 & ~n28098;
  assign n28173 = ~n28171 & ~n28172;
  assign n28174 = ~pi785 & ~n28173;
  assign n28175 = ~n15786 & ~n28098;
  assign n28176 = pi609 & n28171;
  assign n28177 = ~n28175 & ~n28176;
  assign n28178 = pi1155 & ~n28177;
  assign n28179 = ~n16585 & ~n28098;
  assign n28180 = ~pi609 & n28171;
  assign n28181 = ~n28179 & ~n28180;
  assign n28182 = ~pi1155 & ~n28181;
  assign n28183 = ~n28178 & ~n28182;
  assign n28184 = pi785 & ~n28183;
  assign n28185 = ~n28174 & ~n28184;
  assign n28186 = ~pi781 & ~n28185;
  assign n28187 = ~pi618 & n28098;
  assign n28188 = pi618 & n28185;
  assign n28189 = pi1154 & ~n28187;
  assign n28190 = ~n28188 & n28189;
  assign n28191 = ~pi618 & n28185;
  assign n28192 = pi618 & n28098;
  assign n28193 = ~pi1154 & ~n28192;
  assign n28194 = ~n28191 & n28193;
  assign n28195 = ~n28190 & ~n28194;
  assign n28196 = pi781 & ~n28195;
  assign n28197 = ~n28186 & ~n28196;
  assign n28198 = ~pi789 & ~n28197;
  assign n28199 = ~pi619 & n28098;
  assign n28200 = pi619 & n28197;
  assign n28201 = pi1159 & ~n28199;
  assign n28202 = ~n28200 & n28201;
  assign n28203 = ~pi619 & n28197;
  assign n28204 = pi619 & n28098;
  assign n28205 = ~pi1159 & ~n28204;
  assign n28206 = ~n28203 & n28205;
  assign n28207 = ~n28202 & ~n28206;
  assign n28208 = pi789 & ~n28207;
  assign n28209 = ~n28198 & ~n28208;
  assign n28210 = ~n15832 & n28209;
  assign n28211 = n15832 & n28098;
  assign n28212 = ~n28210 & ~n28211;
  assign n28213 = ~n16633 & n28212;
  assign n28214 = pi629 & n28145;
  assign n28215 = ~n28162 & ~n28214;
  assign n28216 = ~n28213 & n28215;
  assign n28217 = pi792 & ~n28216;
  assign n28218 = pi619 & n28131;
  assign n28219 = ~pi1159 & ~n28218;
  assign n28220 = ~pi648 & ~n28202;
  assign n28221 = ~n28219 & n28220;
  assign n28222 = pi618 & ~n28129;
  assign n28223 = pi609 & n28126;
  assign n28224 = ~pi726 & n28168;
  assign n28225 = ~pi187 & n18675;
  assign n28226 = pi187 & n18666;
  assign n28227 = ~n18668 & ~n28226;
  assign n28228 = ~n28225 & n28227;
  assign n28229 = pi770 & ~n28228;
  assign n28230 = pi187 & ~n18659;
  assign n28231 = ~pi187 & n18651;
  assign n28232 = ~pi770 & ~n28231;
  assign n28233 = ~n28230 & n28232;
  assign n28234 = ~n28229 & ~n28233;
  assign n28235 = pi726 & ~n28234;
  assign n28236 = n9829 & ~n28224;
  assign n28237 = ~n28235 & n28236;
  assign n28238 = ~n28101 & ~n28237;
  assign n28239 = ~pi625 & n28238;
  assign n28240 = pi625 & n28170;
  assign n28241 = ~pi1153 & ~n28240;
  assign n28242 = ~n28239 & n28241;
  assign n28243 = ~pi608 & ~n28119;
  assign n28244 = ~n28242 & n28243;
  assign n28245 = ~pi625 & n28170;
  assign n28246 = pi625 & n28238;
  assign n28247 = pi1153 & ~n28245;
  assign n28248 = ~n28246 & n28247;
  assign n28249 = pi608 & ~n28123;
  assign n28250 = ~n28248 & n28249;
  assign n28251 = ~n28244 & ~n28250;
  assign n28252 = pi778 & ~n28251;
  assign n28253 = ~pi778 & n28238;
  assign n28254 = ~n28252 & ~n28253;
  assign n28255 = ~pi609 & ~n28254;
  assign n28256 = ~pi1155 & ~n28223;
  assign n28257 = ~n28255 & n28256;
  assign n28258 = ~pi660 & ~n28178;
  assign n28259 = ~n28257 & n28258;
  assign n28260 = ~pi609 & n28126;
  assign n28261 = pi609 & ~n28254;
  assign n28262 = pi1155 & ~n28260;
  assign n28263 = ~n28261 & n28262;
  assign n28264 = pi660 & ~n28182;
  assign n28265 = ~n28263 & n28264;
  assign n28266 = ~n28259 & ~n28265;
  assign n28267 = pi785 & ~n28266;
  assign n28268 = ~pi785 & ~n28254;
  assign n28269 = ~n28267 & ~n28268;
  assign n28270 = ~pi618 & ~n28269;
  assign n28271 = ~pi1154 & ~n28222;
  assign n28272 = ~n28270 & n28271;
  assign n28273 = ~pi627 & ~n28190;
  assign n28274 = ~n28272 & n28273;
  assign n28275 = ~pi618 & ~n28129;
  assign n28276 = pi618 & ~n28269;
  assign n28277 = pi1154 & ~n28275;
  assign n28278 = ~n28276 & n28277;
  assign n28279 = pi627 & ~n28194;
  assign n28280 = ~n28278 & n28279;
  assign n28281 = ~n28274 & ~n28280;
  assign n28282 = pi781 & ~n28281;
  assign n28283 = ~pi781 & ~n28269;
  assign n28284 = ~n28282 & ~n28283;
  assign n28285 = pi619 & ~n28284;
  assign n28286 = ~pi619 & n28131;
  assign n28287 = pi1159 & ~n28286;
  assign n28288 = ~n28285 & n28287;
  assign n28289 = pi648 & ~n28206;
  assign n28290 = ~n28288 & n28289;
  assign n28291 = ~n28221 & ~n28290;
  assign n28292 = pi789 & ~n28291;
  assign n28293 = ~pi619 & n28220;
  assign n28294 = pi789 & ~n28293;
  assign n28295 = ~n28284 & ~n28294;
  assign n28296 = ~n28292 & ~n28295;
  assign n28297 = n15833 & ~n28296;
  assign n28298 = pi641 & ~n28098;
  assign n28299 = ~pi641 & n28134;
  assign n28300 = n15819 & ~n28298;
  assign n28301 = ~n28299 & n28300;
  assign n28302 = n22348 & n28209;
  assign n28303 = ~pi641 & ~n28098;
  assign n28304 = pi641 & n28134;
  assign n28305 = n15818 & ~n28303;
  assign n28306 = ~n28304 & n28305;
  assign n28307 = ~n28301 & ~n28306;
  assign n28308 = ~n28302 & n28307;
  assign n28309 = pi788 & ~n28308;
  assign n28310 = ~n16644 & ~n28309;
  assign n28311 = ~n28297 & n28310;
  assign n28312 = ~n28217 & ~n28311;
  assign n28313 = ~pi647 & n28312;
  assign n28314 = ~n15925 & ~n28212;
  assign n28315 = n15925 & n28098;
  assign n28316 = ~n28314 & ~n28315;
  assign n28317 = pi647 & ~n28316;
  assign n28318 = ~pi1157 & ~n28317;
  assign n28319 = ~n28313 & n28318;
  assign n28320 = ~pi630 & ~n28153;
  assign n28321 = ~n28319 & n28320;
  assign n28322 = ~pi647 & ~n28316;
  assign n28323 = pi647 & n28312;
  assign n28324 = pi1157 & ~n28322;
  assign n28325 = ~n28323 & n28324;
  assign n28326 = pi630 & ~n28157;
  assign n28327 = ~n28325 & n28326;
  assign n28328 = ~n28321 & ~n28327;
  assign n28329 = pi787 & ~n28328;
  assign n28330 = ~pi787 & n28312;
  assign n28331 = ~n28329 & ~n28330;
  assign n28332 = pi644 & ~n28331;
  assign n28333 = pi715 & ~n28161;
  assign n28334 = ~n28332 & n28333;
  assign n28335 = ~n15960 & ~n28316;
  assign n28336 = n15960 & n28098;
  assign n28337 = ~n28335 & ~n28336;
  assign n28338 = pi644 & ~n28337;
  assign n28339 = ~pi644 & n28098;
  assign n28340 = ~pi715 & ~n28339;
  assign n28341 = ~n28338 & n28340;
  assign n28342 = pi1160 & ~n28341;
  assign n28343 = ~n28334 & n28342;
  assign n28344 = pi644 & n28160;
  assign n28345 = ~pi715 & ~n28344;
  assign n28346 = ~pi644 & ~n28337;
  assign n28347 = pi644 & n28098;
  assign n28348 = pi715 & ~n28347;
  assign n28349 = ~n28346 & n28348;
  assign n28350 = ~pi1160 & ~n28349;
  assign n28351 = ~n28345 & n28350;
  assign n28352 = ~n28343 & ~n28351;
  assign n28353 = pi790 & ~n28352;
  assign n28354 = ~pi644 & n28350;
  assign n28355 = pi790 & ~n28354;
  assign n28356 = ~n28331 & ~n28355;
  assign n28357 = ~n28353 & ~n28356;
  assign n28358 = ~po1038 & ~n28357;
  assign n28359 = ~pi832 & ~n28097;
  assign n28360 = ~n28358 & n28359;
  assign po344 = ~n28096 & ~n28360;
  assign n28362 = ~pi188 & ~n2923;
  assign n28363 = pi705 & n15726;
  assign n28364 = ~n28362 & ~n28363;
  assign n28365 = ~pi778 & n28364;
  assign n28366 = ~pi625 & n28363;
  assign n28367 = ~n28364 & ~n28366;
  assign n28368 = pi1153 & ~n28367;
  assign n28369 = ~pi1153 & ~n28362;
  assign n28370 = ~n28366 & n28369;
  assign n28371 = ~n28368 & ~n28370;
  assign n28372 = pi778 & ~n28371;
  assign n28373 = ~n28365 & ~n28372;
  assign n28374 = ~n15742 & n28373;
  assign n28375 = ~n15748 & n28374;
  assign n28376 = ~n15754 & n28375;
  assign n28377 = ~n15760 & n28376;
  assign n28378 = ~n15766 & n28377;
  assign n28379 = n19394 & n28378;
  assign n28380 = ~n19394 & n28362;
  assign n28381 = ~n28379 & ~n28380;
  assign n28382 = ~n15959 & n28381;
  assign n28383 = n15925 & n28362;
  assign n28384 = ~pi768 & n15781;
  assign n28385 = ~n28362 & ~n28384;
  assign n28386 = ~n15778 & ~n28385;
  assign n28387 = ~pi785 & ~n28386;
  assign n28388 = ~n15787 & ~n28385;
  assign n28389 = pi1155 & ~n28388;
  assign n28390 = ~n15790 & n28386;
  assign n28391 = ~pi1155 & ~n28390;
  assign n28392 = ~n28389 & ~n28391;
  assign n28393 = pi785 & ~n28392;
  assign n28394 = ~n28387 & ~n28393;
  assign n28395 = ~pi781 & ~n28394;
  assign n28396 = ~n15797 & n28394;
  assign n28397 = pi1154 & ~n28396;
  assign n28398 = ~n15800 & n28394;
  assign n28399 = ~pi1154 & ~n28398;
  assign n28400 = ~n28397 & ~n28399;
  assign n28401 = pi781 & ~n28400;
  assign n28402 = ~n28395 & ~n28401;
  assign n28403 = ~pi789 & ~n28402;
  assign n28404 = ~pi619 & n28362;
  assign n28405 = pi619 & n28402;
  assign n28406 = pi1159 & ~n28404;
  assign n28407 = ~n28405 & n28406;
  assign n28408 = ~pi619 & n28402;
  assign n28409 = pi619 & n28362;
  assign n28410 = ~pi1159 & ~n28409;
  assign n28411 = ~n28408 & n28410;
  assign n28412 = ~n28407 & ~n28411;
  assign n28413 = pi789 & ~n28412;
  assign n28414 = ~n28403 & ~n28413;
  assign n28415 = ~n15832 & ~n28414;
  assign n28416 = n15832 & ~n28362;
  assign n28417 = ~n28415 & ~n28416;
  assign n28418 = ~n15925 & n28417;
  assign n28419 = n19478 & ~n28383;
  assign n28420 = ~n28418 & n28419;
  assign n28421 = ~n28382 & ~n28420;
  assign n28422 = pi787 & ~n28421;
  assign n28423 = n15828 & n28376;
  assign n28424 = ~pi626 & ~n28362;
  assign n28425 = pi626 & ~n28414;
  assign n28426 = n15756 & ~n28424;
  assign n28427 = ~n28425 & n28426;
  assign n28428 = pi626 & ~n28362;
  assign n28429 = ~pi626 & ~n28414;
  assign n28430 = n15757 & ~n28428;
  assign n28431 = ~n28429 & n28430;
  assign n28432 = ~n28423 & ~n28427;
  assign n28433 = ~n28431 & n28432;
  assign n28434 = pi788 & ~n28433;
  assign n28435 = pi618 & n28374;
  assign n28436 = pi609 & n28373;
  assign n28437 = ~n15780 & ~n28364;
  assign n28438 = pi625 & n28437;
  assign n28439 = n28385 & ~n28437;
  assign n28440 = ~n28438 & ~n28439;
  assign n28441 = n28369 & ~n28440;
  assign n28442 = ~pi608 & ~n28368;
  assign n28443 = ~n28441 & n28442;
  assign n28444 = pi1153 & n28385;
  assign n28445 = ~n28438 & n28444;
  assign n28446 = pi608 & ~n28370;
  assign n28447 = ~n28445 & n28446;
  assign n28448 = ~n28443 & ~n28447;
  assign n28449 = pi778 & ~n28448;
  assign n28450 = ~pi778 & ~n28439;
  assign n28451 = ~n28449 & ~n28450;
  assign n28452 = ~pi609 & ~n28451;
  assign n28453 = ~pi1155 & ~n28436;
  assign n28454 = ~n28452 & n28453;
  assign n28455 = ~pi660 & ~n28389;
  assign n28456 = ~n28454 & n28455;
  assign n28457 = ~pi609 & n28373;
  assign n28458 = pi609 & ~n28451;
  assign n28459 = pi1155 & ~n28457;
  assign n28460 = ~n28458 & n28459;
  assign n28461 = pi660 & ~n28391;
  assign n28462 = ~n28460 & n28461;
  assign n28463 = ~n28456 & ~n28462;
  assign n28464 = pi785 & ~n28463;
  assign n28465 = ~pi785 & ~n28451;
  assign n28466 = ~n28464 & ~n28465;
  assign n28467 = ~pi618 & ~n28466;
  assign n28468 = ~pi1154 & ~n28435;
  assign n28469 = ~n28467 & n28468;
  assign n28470 = ~pi627 & ~n28397;
  assign n28471 = ~n28469 & n28470;
  assign n28472 = ~pi618 & n28374;
  assign n28473 = pi618 & ~n28466;
  assign n28474 = pi1154 & ~n28472;
  assign n28475 = ~n28473 & n28474;
  assign n28476 = pi627 & ~n28399;
  assign n28477 = ~n28475 & n28476;
  assign n28478 = ~n28471 & ~n28477;
  assign n28479 = pi781 & ~n28478;
  assign n28480 = ~pi781 & ~n28466;
  assign n28481 = ~n28479 & ~n28480;
  assign n28482 = ~pi789 & n28481;
  assign n28483 = ~pi619 & n28375;
  assign n28484 = pi619 & ~n28481;
  assign n28485 = pi1159 & ~n28483;
  assign n28486 = ~n28484 & n28485;
  assign n28487 = pi648 & ~n28411;
  assign n28488 = ~n28486 & n28487;
  assign n28489 = pi619 & n28375;
  assign n28490 = ~pi619 & ~n28481;
  assign n28491 = ~pi1159 & ~n28489;
  assign n28492 = ~n28490 & n28491;
  assign n28493 = ~pi648 & ~n28407;
  assign n28494 = ~n28492 & n28493;
  assign n28495 = pi789 & ~n28488;
  assign n28496 = ~n28494 & n28495;
  assign n28497 = n15833 & ~n28482;
  assign n28498 = ~n28496 & n28497;
  assign n28499 = ~n28434 & ~n28498;
  assign n28500 = ~n16644 & ~n28499;
  assign n28501 = n15763 & n28417;
  assign n28502 = n15772 & n28377;
  assign n28503 = ~pi629 & ~n28502;
  assign n28504 = ~n28501 & n28503;
  assign n28505 = n15762 & n28417;
  assign n28506 = n15909 & n28377;
  assign n28507 = pi629 & ~n28506;
  assign n28508 = ~n28505 & n28507;
  assign n28509 = pi792 & ~n28504;
  assign n28510 = ~n28508 & n28509;
  assign n28511 = n18841 & ~n28510;
  assign n28512 = ~n28500 & n28511;
  assign n28513 = ~n28422 & ~n28512;
  assign n28514 = ~pi790 & n28513;
  assign n28515 = pi787 & ~n28381;
  assign n28516 = ~pi787 & n28378;
  assign n28517 = ~n28515 & ~n28516;
  assign n28518 = ~pi644 & ~n28517;
  assign n28519 = pi644 & n28513;
  assign n28520 = pi715 & ~n28518;
  assign n28521 = ~n28519 & n28520;
  assign n28522 = ~n19771 & n28362;
  assign n28523 = ~n15960 & n28418;
  assign n28524 = ~n28522 & ~n28523;
  assign n28525 = pi644 & ~n28524;
  assign n28526 = ~pi644 & n28362;
  assign n28527 = ~pi715 & ~n28526;
  assign n28528 = ~n28525 & n28527;
  assign n28529 = pi1160 & ~n28528;
  assign n28530 = ~n28521 & n28529;
  assign n28531 = ~pi644 & ~n28524;
  assign n28532 = pi644 & n28362;
  assign n28533 = pi715 & ~n28532;
  assign n28534 = ~n28531 & n28533;
  assign n28535 = pi644 & ~n28517;
  assign n28536 = ~pi644 & n28513;
  assign n28537 = ~pi715 & ~n28535;
  assign n28538 = ~n28536 & n28537;
  assign n28539 = ~pi1160 & ~n28534;
  assign n28540 = ~n28538 & n28539;
  assign n28541 = ~n28530 & ~n28540;
  assign n28542 = pi790 & ~n28541;
  assign n28543 = pi832 & ~n28514;
  assign n28544 = ~n28542 & n28543;
  assign n28545 = ~pi188 & po1038;
  assign n28546 = ~pi188 & ~n16219;
  assign n28547 = n15759 & ~n28546;
  assign n28548 = n15747 & ~n28546;
  assign n28549 = pi188 & ~n9829;
  assign n28550 = ~pi188 & ~n16228;
  assign n28551 = n16227 & ~n28550;
  assign n28552 = pi188 & n17272;
  assign n28553 = ~pi188 & ~n17276;
  assign n28554 = ~pi38 & ~n28552;
  assign n28555 = ~n28553 & n28554;
  assign n28556 = pi705 & ~n28551;
  assign n28557 = ~n28555 & n28556;
  assign n28558 = ~pi188 & ~pi705;
  assign n28559 = ~n16218 & n28558;
  assign n28560 = n9829 & ~n28557;
  assign n28561 = ~n28559 & n28560;
  assign n28562 = ~n28549 & ~n28561;
  assign n28563 = ~pi778 & ~n28562;
  assign n28564 = ~pi625 & n28546;
  assign n28565 = pi625 & n28562;
  assign n28566 = pi1153 & ~n28564;
  assign n28567 = ~n28565 & n28566;
  assign n28568 = ~pi625 & n28562;
  assign n28569 = pi625 & n28546;
  assign n28570 = ~pi1153 & ~n28569;
  assign n28571 = ~n28568 & n28570;
  assign n28572 = ~n28567 & ~n28571;
  assign n28573 = pi778 & ~n28572;
  assign n28574 = ~n28563 & ~n28573;
  assign n28575 = ~n15741 & n28574;
  assign n28576 = n15741 & n28546;
  assign n28577 = ~n28575 & ~n28576;
  assign n28578 = ~n15747 & n28577;
  assign n28579 = ~n28548 & ~n28578;
  assign n28580 = ~n15753 & n28579;
  assign n28581 = n15753 & n28546;
  assign n28582 = ~n28580 & ~n28581;
  assign n28583 = ~n15759 & n28582;
  assign n28584 = ~n28547 & ~n28583;
  assign n28585 = ~pi792 & ~n28584;
  assign n28586 = ~pi628 & ~n28546;
  assign n28587 = pi628 & ~n28584;
  assign n28588 = ~n28586 & ~n28587;
  assign n28589 = pi1156 & ~n28588;
  assign n28590 = ~pi628 & n28584;
  assign n28591 = pi628 & n28546;
  assign n28592 = ~pi1156 & ~n28591;
  assign n28593 = ~n28590 & n28592;
  assign n28594 = ~n28589 & ~n28593;
  assign n28595 = pi792 & ~n28594;
  assign n28596 = ~n28585 & ~n28595;
  assign n28597 = ~pi787 & ~n28596;
  assign n28598 = ~pi647 & n28546;
  assign n28599 = pi647 & n28596;
  assign n28600 = pi1157 & ~n28598;
  assign n28601 = ~n28599 & n28600;
  assign n28602 = ~pi647 & n28596;
  assign n28603 = pi647 & n28546;
  assign n28604 = ~pi1157 & ~n28603;
  assign n28605 = ~n28602 & n28604;
  assign n28606 = ~n28601 & ~n28605;
  assign n28607 = pi787 & ~n28606;
  assign n28608 = ~n28597 & ~n28607;
  assign n28609 = ~pi644 & n28608;
  assign n28610 = ~pi629 & n28589;
  assign n28611 = pi768 & n16218;
  assign n28612 = ~pi768 & ~n23191;
  assign n28613 = pi188 & ~n28612;
  assign n28614 = ~pi188 & ~pi768;
  assign n28615 = n24555 & n28614;
  assign n28616 = ~n28613 & ~n28615;
  assign n28617 = ~n28611 & n28616;
  assign n28618 = n9829 & ~n28617;
  assign n28619 = ~n28549 & ~n28618;
  assign n28620 = ~n15777 & ~n28619;
  assign n28621 = n15777 & ~n28546;
  assign n28622 = ~n28620 & ~n28621;
  assign n28623 = ~pi785 & ~n28622;
  assign n28624 = ~n15786 & ~n28546;
  assign n28625 = pi609 & n28620;
  assign n28626 = ~n28624 & ~n28625;
  assign n28627 = pi1155 & ~n28626;
  assign n28628 = ~n16585 & ~n28546;
  assign n28629 = ~pi609 & n28620;
  assign n28630 = ~n28628 & ~n28629;
  assign n28631 = ~pi1155 & ~n28630;
  assign n28632 = ~n28627 & ~n28631;
  assign n28633 = pi785 & ~n28632;
  assign n28634 = ~n28623 & ~n28633;
  assign n28635 = ~pi781 & ~n28634;
  assign n28636 = ~pi618 & n28546;
  assign n28637 = pi618 & n28634;
  assign n28638 = pi1154 & ~n28636;
  assign n28639 = ~n28637 & n28638;
  assign n28640 = ~pi618 & n28634;
  assign n28641 = pi618 & n28546;
  assign n28642 = ~pi1154 & ~n28641;
  assign n28643 = ~n28640 & n28642;
  assign n28644 = ~n28639 & ~n28643;
  assign n28645 = pi781 & ~n28644;
  assign n28646 = ~n28635 & ~n28645;
  assign n28647 = ~pi789 & ~n28646;
  assign n28648 = ~pi619 & n28546;
  assign n28649 = pi619 & n28646;
  assign n28650 = pi1159 & ~n28648;
  assign n28651 = ~n28649 & n28650;
  assign n28652 = ~pi619 & n28646;
  assign n28653 = pi619 & n28546;
  assign n28654 = ~pi1159 & ~n28653;
  assign n28655 = ~n28652 & n28654;
  assign n28656 = ~n28651 & ~n28655;
  assign n28657 = pi789 & ~n28656;
  assign n28658 = ~n28647 & ~n28657;
  assign n28659 = ~n15832 & n28658;
  assign n28660 = n15832 & n28546;
  assign n28661 = ~n28659 & ~n28660;
  assign n28662 = ~n16633 & n28661;
  assign n28663 = pi629 & n28593;
  assign n28664 = ~n28610 & ~n28663;
  assign n28665 = ~n28662 & n28664;
  assign n28666 = pi792 & ~n28665;
  assign n28667 = pi619 & n28579;
  assign n28668 = ~pi1159 & ~n28667;
  assign n28669 = ~pi648 & ~n28651;
  assign n28670 = ~n28668 & n28669;
  assign n28671 = pi618 & ~n28577;
  assign n28672 = pi609 & n28574;
  assign n28673 = ~pi705 & n28617;
  assign n28674 = ~pi188 & n18675;
  assign n28675 = pi188 & n18666;
  assign n28676 = ~n18668 & ~n28675;
  assign n28677 = ~n28674 & n28676;
  assign n28678 = pi768 & ~n28677;
  assign n28679 = pi188 & ~n18659;
  assign n28680 = ~pi188 & n18651;
  assign n28681 = ~pi768 & ~n28680;
  assign n28682 = ~n28679 & n28681;
  assign n28683 = ~n28678 & ~n28682;
  assign n28684 = pi705 & ~n28683;
  assign n28685 = n9829 & ~n28673;
  assign n28686 = ~n28684 & n28685;
  assign n28687 = ~n28549 & ~n28686;
  assign n28688 = ~pi625 & n28687;
  assign n28689 = pi625 & n28619;
  assign n28690 = ~pi1153 & ~n28689;
  assign n28691 = ~n28688 & n28690;
  assign n28692 = ~pi608 & ~n28567;
  assign n28693 = ~n28691 & n28692;
  assign n28694 = ~pi625 & n28619;
  assign n28695 = pi625 & n28687;
  assign n28696 = pi1153 & ~n28694;
  assign n28697 = ~n28695 & n28696;
  assign n28698 = pi608 & ~n28571;
  assign n28699 = ~n28697 & n28698;
  assign n28700 = ~n28693 & ~n28699;
  assign n28701 = pi778 & ~n28700;
  assign n28702 = ~pi778 & n28687;
  assign n28703 = ~n28701 & ~n28702;
  assign n28704 = ~pi609 & ~n28703;
  assign n28705 = ~pi1155 & ~n28672;
  assign n28706 = ~n28704 & n28705;
  assign n28707 = ~pi660 & ~n28627;
  assign n28708 = ~n28706 & n28707;
  assign n28709 = ~pi609 & n28574;
  assign n28710 = pi609 & ~n28703;
  assign n28711 = pi1155 & ~n28709;
  assign n28712 = ~n28710 & n28711;
  assign n28713 = pi660 & ~n28631;
  assign n28714 = ~n28712 & n28713;
  assign n28715 = ~n28708 & ~n28714;
  assign n28716 = pi785 & ~n28715;
  assign n28717 = ~pi785 & ~n28703;
  assign n28718 = ~n28716 & ~n28717;
  assign n28719 = ~pi618 & ~n28718;
  assign n28720 = ~pi1154 & ~n28671;
  assign n28721 = ~n28719 & n28720;
  assign n28722 = ~pi627 & ~n28639;
  assign n28723 = ~n28721 & n28722;
  assign n28724 = ~pi618 & ~n28577;
  assign n28725 = pi618 & ~n28718;
  assign n28726 = pi1154 & ~n28724;
  assign n28727 = ~n28725 & n28726;
  assign n28728 = pi627 & ~n28643;
  assign n28729 = ~n28727 & n28728;
  assign n28730 = ~n28723 & ~n28729;
  assign n28731 = pi781 & ~n28730;
  assign n28732 = ~pi781 & ~n28718;
  assign n28733 = ~n28731 & ~n28732;
  assign n28734 = pi619 & ~n28733;
  assign n28735 = ~pi619 & n28579;
  assign n28736 = pi1159 & ~n28735;
  assign n28737 = ~n28734 & n28736;
  assign n28738 = pi648 & ~n28655;
  assign n28739 = ~n28737 & n28738;
  assign n28740 = ~n28670 & ~n28739;
  assign n28741 = pi789 & ~n28740;
  assign n28742 = ~pi619 & n28669;
  assign n28743 = pi789 & ~n28742;
  assign n28744 = ~n28733 & ~n28743;
  assign n28745 = ~n28741 & ~n28744;
  assign n28746 = n15833 & ~n28745;
  assign n28747 = pi641 & ~n28546;
  assign n28748 = ~pi641 & n28582;
  assign n28749 = n15819 & ~n28747;
  assign n28750 = ~n28748 & n28749;
  assign n28751 = n22348 & n28658;
  assign n28752 = ~pi641 & ~n28546;
  assign n28753 = pi641 & n28582;
  assign n28754 = n15818 & ~n28752;
  assign n28755 = ~n28753 & n28754;
  assign n28756 = ~n28750 & ~n28755;
  assign n28757 = ~n28751 & n28756;
  assign n28758 = pi788 & ~n28757;
  assign n28759 = ~n16644 & ~n28758;
  assign n28760 = ~n28746 & n28759;
  assign n28761 = ~n28666 & ~n28760;
  assign n28762 = ~pi647 & n28761;
  assign n28763 = ~n15925 & ~n28661;
  assign n28764 = n15925 & n28546;
  assign n28765 = ~n28763 & ~n28764;
  assign n28766 = pi647 & ~n28765;
  assign n28767 = ~pi1157 & ~n28766;
  assign n28768 = ~n28762 & n28767;
  assign n28769 = ~pi630 & ~n28601;
  assign n28770 = ~n28768 & n28769;
  assign n28771 = ~pi647 & ~n28765;
  assign n28772 = pi647 & n28761;
  assign n28773 = pi1157 & ~n28771;
  assign n28774 = ~n28772 & n28773;
  assign n28775 = pi630 & ~n28605;
  assign n28776 = ~n28774 & n28775;
  assign n28777 = ~n28770 & ~n28776;
  assign n28778 = pi787 & ~n28777;
  assign n28779 = ~pi787 & n28761;
  assign n28780 = ~n28778 & ~n28779;
  assign n28781 = pi644 & ~n28780;
  assign n28782 = pi715 & ~n28609;
  assign n28783 = ~n28781 & n28782;
  assign n28784 = ~n15960 & ~n28765;
  assign n28785 = n15960 & n28546;
  assign n28786 = ~n28784 & ~n28785;
  assign n28787 = pi644 & ~n28786;
  assign n28788 = ~pi644 & n28546;
  assign n28789 = ~pi715 & ~n28788;
  assign n28790 = ~n28787 & n28789;
  assign n28791 = pi1160 & ~n28790;
  assign n28792 = ~n28783 & n28791;
  assign n28793 = pi644 & n28608;
  assign n28794 = ~pi715 & ~n28793;
  assign n28795 = ~pi644 & ~n28786;
  assign n28796 = pi644 & n28546;
  assign n28797 = pi715 & ~n28796;
  assign n28798 = ~n28795 & n28797;
  assign n28799 = ~pi1160 & ~n28798;
  assign n28800 = ~n28794 & n28799;
  assign n28801 = ~n28792 & ~n28800;
  assign n28802 = pi790 & ~n28801;
  assign n28803 = ~pi644 & n28799;
  assign n28804 = pi790 & ~n28803;
  assign n28805 = ~n28780 & ~n28804;
  assign n28806 = ~n28802 & ~n28805;
  assign n28807 = ~po1038 & ~n28806;
  assign n28808 = ~pi832 & ~n28545;
  assign n28809 = ~n28807 & n28808;
  assign po345 = ~n28544 & ~n28809;
  assign n28811 = pi189 & ~n2923;
  assign n28812 = pi772 & n15781;
  assign n28813 = n18872 & n28812;
  assign n28814 = ~pi626 & n28813;
  assign n28815 = ~n28811 & ~n28814;
  assign n28816 = ~pi1158 & ~n28815;
  assign n28817 = pi727 & n15726;
  assign n28818 = ~n28811 & ~n28817;
  assign n28819 = ~pi778 & n28818;
  assign n28820 = pi625 & n28817;
  assign n28821 = ~n28818 & ~n28820;
  assign n28822 = ~pi1153 & ~n28821;
  assign n28823 = pi1153 & ~n28811;
  assign n28824 = ~n28820 & n28823;
  assign n28825 = ~n28822 & ~n28824;
  assign n28826 = pi778 & ~n28825;
  assign n28827 = ~n28819 & ~n28826;
  assign n28828 = n17584 & n28827;
  assign n28829 = ~n15753 & n28828;
  assign n28830 = ~n28811 & ~n28829;
  assign n28831 = n15818 & ~n28830;
  assign n28832 = pi641 & ~n28816;
  assign n28833 = ~n28831 & n28832;
  assign n28834 = n15819 & ~n28830;
  assign n28835 = pi626 & n28813;
  assign n28836 = ~n28811 & ~n28835;
  assign n28837 = pi1158 & ~n28836;
  assign n28838 = ~pi641 & ~n28837;
  assign n28839 = ~n28834 & n28838;
  assign n28840 = pi788 & ~n28833;
  assign n28841 = ~n28839 & n28840;
  assign n28842 = ~n18944 & ~n28828;
  assign n28843 = ~n18861 & n28812;
  assign n28844 = ~n18869 & n28843;
  assign n28845 = ~n15752 & ~n28844;
  assign n28846 = ~n22083 & ~n28845;
  assign n28847 = ~n28842 & n28846;
  assign n28848 = pi789 & ~n28811;
  assign n28849 = ~n28847 & n28848;
  assign n28850 = ~n28811 & ~n28812;
  assign n28851 = ~n15780 & n28817;
  assign n28852 = n28850 & ~n28851;
  assign n28853 = pi625 & n28851;
  assign n28854 = ~n28852 & ~n28853;
  assign n28855 = ~pi1153 & ~n28854;
  assign n28856 = ~pi608 & ~n28824;
  assign n28857 = ~n28855 & n28856;
  assign n28858 = pi1153 & n28850;
  assign n28859 = ~n28853 & n28858;
  assign n28860 = pi608 & ~n28822;
  assign n28861 = ~n28859 & n28860;
  assign n28862 = ~n28857 & ~n28861;
  assign n28863 = pi778 & ~n28862;
  assign n28864 = ~pi778 & ~n28852;
  assign n28865 = ~n28863 & ~n28864;
  assign n28866 = ~pi609 & n28865;
  assign n28867 = pi609 & ~n28827;
  assign n28868 = ~pi1155 & ~n28867;
  assign n28869 = ~n28866 & n28868;
  assign n28870 = n22108 & ~n28850;
  assign n28871 = ~n28869 & ~n28870;
  assign n28872 = ~pi660 & ~n28871;
  assign n28873 = n16585 & n28812;
  assign n28874 = ~pi1155 & ~n28811;
  assign n28875 = ~n28873 & n28874;
  assign n28876 = ~pi609 & n28827;
  assign n28877 = pi609 & ~n28865;
  assign n28878 = pi1155 & ~n28876;
  assign n28879 = ~n28877 & n28878;
  assign n28880 = pi660 & ~n28875;
  assign n28881 = ~n28879 & n28880;
  assign n28882 = ~n28872 & ~n28881;
  assign n28883 = pi785 & ~n28882;
  assign n28884 = ~pi785 & ~n28865;
  assign n28885 = ~n28883 & ~n28884;
  assign n28886 = ~pi781 & ~n28885;
  assign n28887 = n18955 & n28843;
  assign n28888 = ~pi1154 & ~n28811;
  assign n28889 = ~n28887 & n28888;
  assign n28890 = pi618 & ~n28885;
  assign n28891 = ~n15742 & n28827;
  assign n28892 = ~pi618 & n28891;
  assign n28893 = pi1154 & ~n28892;
  assign n28894 = ~n28890 & n28893;
  assign n28895 = pi627 & ~n28889;
  assign n28896 = ~n28894 & n28895;
  assign n28897 = n18950 & n28843;
  assign n28898 = pi1154 & ~n28811;
  assign n28899 = ~n28897 & n28898;
  assign n28900 = ~pi618 & ~n28885;
  assign n28901 = pi618 & n28891;
  assign n28902 = ~pi1154 & ~n28901;
  assign n28903 = ~n28900 & n28902;
  assign n28904 = ~pi627 & ~n28899;
  assign n28905 = ~n28903 & n28904;
  assign n28906 = ~n28896 & ~n28905;
  assign n28907 = pi781 & ~n28906;
  assign n28908 = ~n22148 & ~n28886;
  assign n28909 = ~n28907 & n28908;
  assign n28910 = n15833 & ~n28849;
  assign n28911 = ~n28909 & n28910;
  assign n28912 = ~n16644 & ~n28841;
  assign n28913 = ~n28911 & n28912;
  assign n28914 = n17586 & n28827;
  assign n28915 = ~pi628 & n28914;
  assign n28916 = pi629 & ~n28915;
  assign n28917 = ~n15832 & n28813;
  assign n28918 = pi628 & ~n28917;
  assign n28919 = ~n28916 & ~n28918;
  assign n28920 = ~pi1156 & ~n28919;
  assign n28921 = pi628 & n28914;
  assign n28922 = ~pi628 & ~n28917;
  assign n28923 = pi629 & ~n28922;
  assign n28924 = pi1156 & ~n28923;
  assign n28925 = ~n28921 & n28924;
  assign n28926 = ~n28920 & ~n28925;
  assign n28927 = pi792 & ~n28811;
  assign n28928 = ~n28926 & n28927;
  assign n28929 = ~n28913 & ~n28928;
  assign n28930 = n18841 & ~n28929;
  assign n28931 = ~n15925 & n28917;
  assign n28932 = pi630 & n28931;
  assign n28933 = ~n15765 & n28914;
  assign n28934 = ~pi630 & ~n28933;
  assign n28935 = pi647 & ~n28934;
  assign n28936 = pi1157 & ~n28932;
  assign n28937 = ~n28935 & n28936;
  assign n28938 = ~pi630 & n28931;
  assign n28939 = pi630 & ~n28933;
  assign n28940 = ~pi647 & ~n28939;
  assign n28941 = ~pi1157 & ~n28938;
  assign n28942 = ~n28940 & n28941;
  assign n28943 = ~n28937 & ~n28942;
  assign n28944 = pi787 & ~n28811;
  assign n28945 = ~n28943 & n28944;
  assign n28946 = ~n28930 & ~n28945;
  assign n28947 = ~pi790 & n28946;
  assign n28948 = ~n17768 & n28933;
  assign n28949 = ~n28811 & ~n28948;
  assign n28950 = ~pi644 & ~n28949;
  assign n28951 = pi644 & n28946;
  assign n28952 = pi715 & ~n28950;
  assign n28953 = ~n28951 & n28952;
  assign n28954 = ~n15832 & n19771;
  assign n28955 = n28813 & n28954;
  assign n28956 = pi644 & n28955;
  assign n28957 = ~pi715 & ~n28811;
  assign n28958 = ~n28956 & n28957;
  assign n28959 = pi1160 & ~n28958;
  assign n28960 = ~n28953 & n28959;
  assign n28961 = ~pi644 & n28955;
  assign n28962 = pi715 & ~n28811;
  assign n28963 = ~n28961 & n28962;
  assign n28964 = ~pi644 & n28946;
  assign n28965 = pi644 & ~n28949;
  assign n28966 = ~pi715 & ~n28965;
  assign n28967 = ~n28964 & n28966;
  assign n28968 = ~pi1160 & ~n28963;
  assign n28969 = ~n28967 & n28968;
  assign n28970 = ~n28960 & ~n28969;
  assign n28971 = pi790 & ~n28970;
  assign n28972 = pi832 & ~n28947;
  assign n28973 = ~n28971 & n28972;
  assign n28974 = pi57 & pi189;
  assign n28975 = ~pi189 & ~n6258;
  assign n28976 = pi189 & ~n16219;
  assign n28977 = n15759 & ~n28976;
  assign n28978 = n15747 & ~n28976;
  assign n28979 = pi727 & n9829;
  assign n28980 = ~n28976 & ~n28979;
  assign n28981 = ~pi189 & ~n17272;
  assign n28982 = pi189 & n17276;
  assign n28983 = ~pi38 & ~n28981;
  assign n28984 = ~n28982 & n28983;
  assign n28985 = ~pi189 & ~n16228;
  assign n28986 = n19049 & ~n28985;
  assign n28987 = n28979 & ~n28986;
  assign n28988 = ~n28984 & n28987;
  assign n28989 = ~n28980 & ~n28988;
  assign n28990 = ~pi778 & n28989;
  assign n28991 = ~pi625 & ~n28976;
  assign n28992 = pi625 & ~n28989;
  assign n28993 = pi1153 & ~n28991;
  assign n28994 = ~n28992 & n28993;
  assign n28995 = ~pi625 & ~n28989;
  assign n28996 = pi625 & ~n28976;
  assign n28997 = ~pi1153 & ~n28996;
  assign n28998 = ~n28995 & n28997;
  assign n28999 = ~n28994 & ~n28998;
  assign n29000 = pi778 & ~n28999;
  assign n29001 = ~n28990 & ~n29000;
  assign n29002 = ~n15741 & ~n29001;
  assign n29003 = n15741 & n28976;
  assign n29004 = ~n29002 & ~n29003;
  assign n29005 = ~n15747 & n29004;
  assign n29006 = ~n28978 & ~n29005;
  assign n29007 = ~n15753 & n29006;
  assign n29008 = n15753 & n28976;
  assign n29009 = ~n29007 & ~n29008;
  assign n29010 = ~n15759 & n29009;
  assign n29011 = ~n28977 & ~n29010;
  assign n29012 = ~pi792 & n29011;
  assign n29013 = pi628 & n29011;
  assign n29014 = ~pi628 & n28976;
  assign n29015 = ~n29013 & ~n29014;
  assign n29016 = pi1156 & ~n29015;
  assign n29017 = pi628 & ~n28976;
  assign n29018 = ~pi628 & ~n29011;
  assign n29019 = ~pi1156 & ~n29017;
  assign n29020 = ~n29018 & n29019;
  assign n29021 = ~n29016 & ~n29020;
  assign n29022 = pi792 & ~n29021;
  assign n29023 = ~n29012 & ~n29022;
  assign n29024 = ~pi787 & ~n29023;
  assign n29025 = ~pi647 & ~n28976;
  assign n29026 = pi647 & n29023;
  assign n29027 = pi1157 & ~n29025;
  assign n29028 = ~n29026 & n29027;
  assign n29029 = pi647 & ~n28976;
  assign n29030 = ~pi647 & n29023;
  assign n29031 = ~pi1157 & ~n29029;
  assign n29032 = ~n29030 & n29031;
  assign n29033 = ~n29028 & ~n29032;
  assign n29034 = pi787 & ~n29033;
  assign n29035 = ~n29024 & ~n29034;
  assign n29036 = ~pi644 & n29035;
  assign n29037 = ~pi629 & n29016;
  assign n29038 = pi619 & ~n29006;
  assign n29039 = ~pi1159 & ~n29038;
  assign n29040 = ~pi619 & ~n28976;
  assign n29041 = pi189 & ~n9829;
  assign n29042 = pi772 & ~n16512;
  assign n29043 = ~n21104 & ~n29042;
  assign n29044 = pi39 & ~n29043;
  assign n29045 = ~pi772 & n16057;
  assign n29046 = n16448 & ~n29045;
  assign n29047 = ~n29044 & ~n29046;
  assign n29048 = pi189 & ~n29047;
  assign n29049 = ~pi189 & pi772;
  assign n29050 = n16565 & n29049;
  assign n29051 = ~n29048 & ~n29050;
  assign n29052 = ~pi38 & ~n29051;
  assign n29053 = pi772 & n15780;
  assign n29054 = n16228 & ~n29053;
  assign n29055 = pi38 & ~n28985;
  assign n29056 = ~n29054 & n29055;
  assign n29057 = ~n29052 & ~n29056;
  assign n29058 = n9829 & ~n29057;
  assign n29059 = ~n29041 & ~n29058;
  assign n29060 = ~n15777 & ~n29059;
  assign n29061 = n15777 & n28976;
  assign n29062 = ~n29060 & ~n29061;
  assign n29063 = ~pi785 & ~n29062;
  assign n29064 = pi609 & n29062;
  assign n29065 = ~pi609 & ~n28976;
  assign n29066 = pi1155 & ~n29065;
  assign n29067 = ~n29064 & n29066;
  assign n29068 = ~pi609 & n29062;
  assign n29069 = pi609 & ~n28976;
  assign n29070 = ~pi1155 & ~n29069;
  assign n29071 = ~n29068 & n29070;
  assign n29072 = ~n29067 & ~n29071;
  assign n29073 = pi785 & ~n29072;
  assign n29074 = ~n29063 & ~n29073;
  assign n29075 = ~pi781 & ~n29074;
  assign n29076 = ~pi618 & ~n28976;
  assign n29077 = pi618 & n29074;
  assign n29078 = pi1154 & ~n29076;
  assign n29079 = ~n29077 & n29078;
  assign n29080 = pi618 & ~n28976;
  assign n29081 = ~pi618 & n29074;
  assign n29082 = ~pi1154 & ~n29080;
  assign n29083 = ~n29081 & n29082;
  assign n29084 = ~n29079 & ~n29083;
  assign n29085 = pi781 & ~n29084;
  assign n29086 = ~n29075 & ~n29085;
  assign n29087 = pi619 & n29086;
  assign n29088 = pi1159 & ~n29040;
  assign n29089 = ~n29087 & n29088;
  assign n29090 = ~pi648 & ~n29089;
  assign n29091 = ~n29039 & n29090;
  assign n29092 = ~pi619 & ~n29006;
  assign n29093 = pi1159 & ~n29092;
  assign n29094 = pi619 & ~n28976;
  assign n29095 = ~pi619 & n29086;
  assign n29096 = ~pi1159 & ~n29094;
  assign n29097 = ~n29095 & n29096;
  assign n29098 = pi648 & ~n29097;
  assign n29099 = ~n29093 & n29098;
  assign n29100 = ~n29091 & ~n29099;
  assign n29101 = pi789 & ~n29100;
  assign n29102 = pi619 & n29098;
  assign n29103 = ~pi619 & n29090;
  assign n29104 = pi789 & ~n29102;
  assign n29105 = ~n29103 & n29104;
  assign n29106 = pi609 & n29001;
  assign n29107 = ~n28979 & ~n29058;
  assign n29108 = ~pi189 & ~n16657;
  assign n29109 = pi189 & ~n16653;
  assign n29110 = ~pi772 & ~n29108;
  assign n29111 = ~n29109 & n29110;
  assign n29112 = ~pi189 & n17397;
  assign n29113 = pi189 & n16647;
  assign n29114 = pi772 & ~n29112;
  assign n29115 = ~n29113 & n29114;
  assign n29116 = ~pi39 & ~n29115;
  assign n29117 = ~n29111 & n29116;
  assign n29118 = pi189 & ~n16877;
  assign n29119 = ~pi189 & ~n16913;
  assign n29120 = pi772 & ~n29118;
  assign n29121 = ~n29119 & n29120;
  assign n29122 = pi189 & n16747;
  assign n29123 = ~pi189 & ~n16825;
  assign n29124 = ~pi772 & ~n29123;
  assign n29125 = ~n29122 & n29124;
  assign n29126 = pi39 & ~n29121;
  assign n29127 = ~n29125 & n29126;
  assign n29128 = ~pi38 & ~n29117;
  assign n29129 = ~n29127 & n29128;
  assign n29130 = pi727 & ~n18668;
  assign n29131 = ~n29056 & n29130;
  assign n29132 = ~n29129 & n29131;
  assign n29133 = ~n29107 & ~n29132;
  assign n29134 = ~n29041 & ~n29133;
  assign n29135 = ~pi625 & n29134;
  assign n29136 = pi625 & n29059;
  assign n29137 = ~pi1153 & ~n29136;
  assign n29138 = ~n29135 & n29137;
  assign n29139 = ~pi608 & ~n28994;
  assign n29140 = ~n29138 & n29139;
  assign n29141 = ~pi625 & n29059;
  assign n29142 = pi625 & n29134;
  assign n29143 = pi1153 & ~n29141;
  assign n29144 = ~n29142 & n29143;
  assign n29145 = pi608 & ~n28998;
  assign n29146 = ~n29144 & n29145;
  assign n29147 = ~n29140 & ~n29146;
  assign n29148 = pi778 & ~n29147;
  assign n29149 = ~pi778 & n29134;
  assign n29150 = ~n29148 & ~n29149;
  assign n29151 = ~pi609 & ~n29150;
  assign n29152 = ~pi1155 & ~n29106;
  assign n29153 = ~n29151 & n29152;
  assign n29154 = ~pi660 & ~n29067;
  assign n29155 = ~n29153 & n29154;
  assign n29156 = ~pi609 & n29001;
  assign n29157 = pi609 & ~n29150;
  assign n29158 = pi1155 & ~n29156;
  assign n29159 = ~n29157 & n29158;
  assign n29160 = pi660 & ~n29071;
  assign n29161 = ~n29159 & n29160;
  assign n29162 = ~n29155 & ~n29161;
  assign n29163 = pi785 & ~n29162;
  assign n29164 = ~pi785 & ~n29150;
  assign n29165 = ~n29163 & ~n29164;
  assign n29166 = ~pi781 & n29165;
  assign n29167 = ~pi618 & ~n29165;
  assign n29168 = pi618 & n29004;
  assign n29169 = ~pi1154 & ~n29168;
  assign n29170 = ~n29167 & n29169;
  assign n29171 = ~pi627 & ~n29079;
  assign n29172 = ~n29170 & n29171;
  assign n29173 = ~pi618 & n29004;
  assign n29174 = pi618 & ~n29165;
  assign n29175 = pi1154 & ~n29173;
  assign n29176 = ~n29174 & n29175;
  assign n29177 = pi627 & ~n29083;
  assign n29178 = ~n29176 & n29177;
  assign n29179 = pi781 & ~n29172;
  assign n29180 = ~n29178 & n29179;
  assign n29181 = ~n29105 & ~n29166;
  assign n29182 = ~n29180 & n29181;
  assign n29183 = ~n29101 & ~n29182;
  assign n29184 = n15833 & ~n29183;
  assign n29185 = pi641 & n28976;
  assign n29186 = ~pi641 & ~n29009;
  assign n29187 = n15819 & ~n29185;
  assign n29188 = ~n29186 & n29187;
  assign n29189 = ~pi789 & ~n29086;
  assign n29190 = ~n29089 & ~n29097;
  assign n29191 = pi789 & ~n29190;
  assign n29192 = ~n29189 & ~n29191;
  assign n29193 = n22348 & n29192;
  assign n29194 = ~pi641 & n28976;
  assign n29195 = pi641 & ~n29009;
  assign n29196 = n15818 & ~n29194;
  assign n29197 = ~n29195 & n29196;
  assign n29198 = ~n29188 & ~n29197;
  assign n29199 = ~n29193 & n29198;
  assign n29200 = pi788 & ~n29199;
  assign n29201 = ~n29184 & ~n29200;
  assign n29202 = ~n16643 & n29201;
  assign n29203 = ~n15832 & ~n29192;
  assign n29204 = n15832 & n28976;
  assign n29205 = ~n29203 & ~n29204;
  assign n29206 = ~n16633 & ~n29205;
  assign n29207 = pi629 & n29020;
  assign n29208 = ~n29037 & ~n29207;
  assign n29209 = ~n29206 & n29208;
  assign n29210 = ~n29202 & n29209;
  assign n29211 = pi792 & ~n29210;
  assign n29212 = ~pi792 & n29201;
  assign n29213 = ~n29211 & ~n29212;
  assign n29214 = ~pi647 & n29213;
  assign n29215 = ~n15925 & ~n29205;
  assign n29216 = n15925 & n28976;
  assign n29217 = ~n29215 & ~n29216;
  assign n29218 = pi647 & n29217;
  assign n29219 = ~pi1157 & ~n29218;
  assign n29220 = ~n29214 & n29219;
  assign n29221 = ~pi630 & ~n29028;
  assign n29222 = ~n29220 & n29221;
  assign n29223 = ~pi647 & n29217;
  assign n29224 = pi647 & n29213;
  assign n29225 = pi1157 & ~n29223;
  assign n29226 = ~n29224 & n29225;
  assign n29227 = pi630 & ~n29032;
  assign n29228 = ~n29226 & n29227;
  assign n29229 = ~n29222 & ~n29228;
  assign n29230 = pi787 & ~n29229;
  assign n29231 = ~pi787 & n29213;
  assign n29232 = ~n29230 & ~n29231;
  assign n29233 = pi644 & ~n29232;
  assign n29234 = pi715 & ~n29036;
  assign n29235 = ~n29233 & n29234;
  assign n29236 = ~n15960 & ~n29217;
  assign n29237 = n15960 & n28976;
  assign n29238 = ~n29236 & ~n29237;
  assign n29239 = pi644 & n29238;
  assign n29240 = ~pi644 & ~n28976;
  assign n29241 = ~pi715 & ~n29240;
  assign n29242 = ~n29239 & n29241;
  assign n29243 = pi1160 & ~n29242;
  assign n29244 = ~n29235 & n29243;
  assign n29245 = pi644 & n29035;
  assign n29246 = ~pi715 & ~n29245;
  assign n29247 = ~pi644 & n29238;
  assign n29248 = pi644 & ~n28976;
  assign n29249 = pi715 & ~n29248;
  assign n29250 = ~n29247 & n29249;
  assign n29251 = ~pi1160 & ~n29250;
  assign n29252 = ~n29246 & n29251;
  assign n29253 = ~n29244 & ~n29252;
  assign n29254 = pi790 & ~n29253;
  assign n29255 = ~pi644 & n29251;
  assign n29256 = pi790 & ~n29255;
  assign n29257 = ~n29232 & ~n29256;
  assign n29258 = ~n29254 & ~n29257;
  assign n29259 = n6258 & ~n29258;
  assign n29260 = ~pi57 & ~n28975;
  assign n29261 = ~n29259 & n29260;
  assign n29262 = ~pi832 & ~n28974;
  assign n29263 = ~n29261 & n29262;
  assign po346 = ~n28973 & ~n29263;
  assign n29265 = ~pi190 & ~n2923;
  assign n29266 = pi699 & n15726;
  assign n29267 = ~n29265 & ~n29266;
  assign n29268 = ~pi778 & ~n29267;
  assign n29269 = ~pi625 & n29266;
  assign n29270 = ~n29267 & ~n29269;
  assign n29271 = pi1153 & ~n29270;
  assign n29272 = ~pi1153 & ~n29265;
  assign n29273 = ~n29269 & n29272;
  assign n29274 = pi778 & ~n29273;
  assign n29275 = ~n29271 & n29274;
  assign n29276 = ~n29268 & ~n29275;
  assign n29277 = ~n15742 & ~n29276;
  assign n29278 = ~n15748 & n29277;
  assign n29279 = ~n15754 & n29278;
  assign n29280 = ~n15760 & n29279;
  assign n29281 = ~n15766 & n29280;
  assign n29282 = n19394 & n29281;
  assign n29283 = ~n19394 & n29265;
  assign n29284 = ~n29282 & ~n29283;
  assign n29285 = ~n15959 & n29284;
  assign n29286 = n15925 & n29265;
  assign n29287 = pi763 & n15781;
  assign n29288 = ~n29265 & ~n29287;
  assign n29289 = ~n15778 & ~n29288;
  assign n29290 = ~pi785 & ~n29289;
  assign n29291 = n16585 & n29287;
  assign n29292 = n29289 & ~n29291;
  assign n29293 = pi1155 & ~n29292;
  assign n29294 = ~pi1155 & ~n29265;
  assign n29295 = ~n29291 & n29294;
  assign n29296 = ~n29293 & ~n29295;
  assign n29297 = pi785 & ~n29296;
  assign n29298 = ~n29290 & ~n29297;
  assign n29299 = ~pi781 & ~n29298;
  assign n29300 = ~n15797 & n29298;
  assign n29301 = pi1154 & ~n29300;
  assign n29302 = ~n15800 & n29298;
  assign n29303 = ~pi1154 & ~n29302;
  assign n29304 = ~n29301 & ~n29303;
  assign n29305 = pi781 & ~n29304;
  assign n29306 = ~n29299 & ~n29305;
  assign n29307 = ~n21915 & n29306;
  assign n29308 = ~n15832 & ~n29307;
  assign n29309 = n15832 & ~n29265;
  assign n29310 = ~n29308 & ~n29309;
  assign n29311 = ~n15925 & n29310;
  assign n29312 = n19478 & ~n29286;
  assign n29313 = ~n29311 & n29312;
  assign n29314 = ~n29285 & ~n29313;
  assign n29315 = pi787 & ~n29314;
  assign n29316 = n15763 & n29310;
  assign n29317 = n15772 & n29280;
  assign n29318 = ~pi629 & ~n29317;
  assign n29319 = ~n29316 & n29318;
  assign n29320 = n15762 & n29310;
  assign n29321 = n15909 & n29280;
  assign n29322 = pi629 & ~n29321;
  assign n29323 = ~n29320 & n29322;
  assign n29324 = pi792 & ~n29319;
  assign n29325 = ~n29323 & n29324;
  assign n29326 = ~n21932 & n29306;
  assign n29327 = pi648 & ~n29326;
  assign n29328 = n21935 & ~n29278;
  assign n29329 = ~n29327 & ~n29328;
  assign n29330 = ~pi1159 & ~n29329;
  assign n29331 = ~pi619 & ~n29278;
  assign n29332 = pi648 & ~n29331;
  assign n29333 = n21942 & n29306;
  assign n29334 = pi1159 & ~n29332;
  assign n29335 = ~n29333 & n29334;
  assign n29336 = ~n29330 & ~n29335;
  assign n29337 = pi789 & ~n29336;
  assign n29338 = pi609 & ~n29276;
  assign n29339 = ~n15780 & ~n29267;
  assign n29340 = pi625 & n29339;
  assign n29341 = n29288 & ~n29339;
  assign n29342 = ~n29340 & ~n29341;
  assign n29343 = n29272 & ~n29342;
  assign n29344 = ~pi608 & ~n29271;
  assign n29345 = ~n29343 & n29344;
  assign n29346 = pi1153 & n29288;
  assign n29347 = ~n29340 & n29346;
  assign n29348 = pi608 & ~n29273;
  assign n29349 = ~n29347 & n29348;
  assign n29350 = ~n29345 & ~n29349;
  assign n29351 = pi778 & ~n29350;
  assign n29352 = ~pi778 & ~n29341;
  assign n29353 = ~n29351 & ~n29352;
  assign n29354 = ~pi609 & ~n29353;
  assign n29355 = ~pi1155 & ~n29338;
  assign n29356 = ~n29354 & n29355;
  assign n29357 = ~pi660 & ~n29293;
  assign n29358 = ~n29356 & n29357;
  assign n29359 = ~pi609 & ~n29276;
  assign n29360 = pi609 & ~n29353;
  assign n29361 = pi1155 & ~n29359;
  assign n29362 = ~n29360 & n29361;
  assign n29363 = pi660 & ~n29295;
  assign n29364 = ~n29362 & n29363;
  assign n29365 = ~n29358 & ~n29364;
  assign n29366 = pi785 & ~n29365;
  assign n29367 = ~pi785 & ~n29353;
  assign n29368 = ~n29366 & ~n29367;
  assign n29369 = ~pi781 & n29368;
  assign n29370 = pi618 & n29277;
  assign n29371 = ~pi618 & ~n29368;
  assign n29372 = ~pi1154 & ~n29370;
  assign n29373 = ~n29371 & n29372;
  assign n29374 = ~pi627 & ~n29301;
  assign n29375 = ~n29373 & n29374;
  assign n29376 = ~pi618 & n29277;
  assign n29377 = pi618 & ~n29368;
  assign n29378 = pi1154 & ~n29376;
  assign n29379 = ~n29377 & n29378;
  assign n29380 = pi627 & ~n29303;
  assign n29381 = ~n29379 & n29380;
  assign n29382 = pi781 & ~n29375;
  assign n29383 = ~n29381 & n29382;
  assign n29384 = ~n29337 & ~n29369;
  assign n29385 = ~n29383 & n29384;
  assign n29386 = n18969 & n29336;
  assign n29387 = ~n29385 & ~n29386;
  assign n29388 = n15833 & ~n29387;
  assign n29389 = n15828 & n29279;
  assign n29390 = ~pi626 & ~n29265;
  assign n29391 = pi626 & ~n29307;
  assign n29392 = n15756 & ~n29390;
  assign n29393 = ~n29391 & n29392;
  assign n29394 = pi626 & ~n29265;
  assign n29395 = ~pi626 & ~n29307;
  assign n29396 = n15757 & ~n29394;
  assign n29397 = ~n29395 & n29396;
  assign n29398 = ~n29389 & ~n29393;
  assign n29399 = ~n29397 & n29398;
  assign n29400 = pi788 & ~n29399;
  assign n29401 = ~n29388 & ~n29400;
  assign n29402 = ~n16644 & ~n29401;
  assign n29403 = n18841 & ~n29325;
  assign n29404 = ~n29402 & n29403;
  assign n29405 = ~n29315 & ~n29404;
  assign n29406 = ~pi790 & n29405;
  assign n29407 = pi787 & ~n29284;
  assign n29408 = ~pi787 & n29281;
  assign n29409 = ~n29407 & ~n29408;
  assign n29410 = ~pi644 & ~n29409;
  assign n29411 = pi644 & n29405;
  assign n29412 = pi715 & ~n29410;
  assign n29413 = ~n29411 & n29412;
  assign n29414 = ~n19771 & n29265;
  assign n29415 = ~n15960 & n29311;
  assign n29416 = ~n29414 & ~n29415;
  assign n29417 = pi644 & ~n29416;
  assign n29418 = ~pi644 & n29265;
  assign n29419 = ~pi715 & ~n29418;
  assign n29420 = ~n29417 & n29419;
  assign n29421 = pi1160 & ~n29420;
  assign n29422 = ~n29413 & n29421;
  assign n29423 = ~pi644 & ~n29416;
  assign n29424 = pi644 & n29265;
  assign n29425 = pi715 & ~n29424;
  assign n29426 = ~n29423 & n29425;
  assign n29427 = pi644 & ~n29409;
  assign n29428 = ~pi644 & n29405;
  assign n29429 = ~pi715 & ~n29427;
  assign n29430 = ~n29428 & n29429;
  assign n29431 = ~pi1160 & ~n29426;
  assign n29432 = ~n29430 & n29431;
  assign n29433 = ~n29422 & ~n29432;
  assign n29434 = pi790 & ~n29433;
  assign n29435 = pi832 & ~n29406;
  assign n29436 = ~n29434 & n29435;
  assign n29437 = ~pi190 & po1038;
  assign n29438 = ~pi190 & ~n16219;
  assign n29439 = n15747 & ~n29438;
  assign n29440 = pi190 & ~n9829;
  assign n29441 = ~pi190 & ~n16228;
  assign n29442 = n16227 & ~n29441;
  assign n29443 = pi190 & n17272;
  assign n29444 = ~pi190 & ~n17276;
  assign n29445 = ~pi38 & ~n29443;
  assign n29446 = ~n29444 & n29445;
  assign n29447 = pi699 & ~n29442;
  assign n29448 = ~n29446 & n29447;
  assign n29449 = ~pi190 & ~pi699;
  assign n29450 = ~n16218 & n29449;
  assign n29451 = n9829 & ~n29448;
  assign n29452 = ~n29450 & n29451;
  assign n29453 = ~n29440 & ~n29452;
  assign n29454 = ~pi778 & ~n29453;
  assign n29455 = ~pi625 & n29438;
  assign n29456 = pi625 & n29453;
  assign n29457 = pi1153 & ~n29455;
  assign n29458 = ~n29456 & n29457;
  assign n29459 = ~pi625 & n29453;
  assign n29460 = pi625 & n29438;
  assign n29461 = ~pi1153 & ~n29460;
  assign n29462 = ~n29459 & n29461;
  assign n29463 = ~n29458 & ~n29462;
  assign n29464 = pi778 & ~n29463;
  assign n29465 = ~n29454 & ~n29464;
  assign n29466 = ~n15741 & n29465;
  assign n29467 = n15741 & n29438;
  assign n29468 = ~n29466 & ~n29467;
  assign n29469 = ~n15747 & n29468;
  assign n29470 = ~n29439 & ~n29469;
  assign n29471 = ~n15753 & n29470;
  assign n29472 = n15753 & n29438;
  assign n29473 = ~n29471 & ~n29472;
  assign n29474 = ~n15759 & ~n29473;
  assign n29475 = n15759 & n29438;
  assign n29476 = ~n29474 & ~n29475;
  assign n29477 = ~n15765 & ~n29476;
  assign n29478 = n15765 & n29438;
  assign n29479 = ~n29477 & ~n29478;
  assign n29480 = ~n17768 & ~n29479;
  assign n29481 = n17768 & n29438;
  assign n29482 = ~n29480 & ~n29481;
  assign n29483 = ~pi644 & ~n29482;
  assign n29484 = pi715 & ~n29483;
  assign n29485 = ~pi763 & n16212;
  assign n29486 = pi190 & ~n16563;
  assign n29487 = ~n29485 & ~n29486;
  assign n29488 = pi39 & ~n29487;
  assign n29489 = pi763 & ~n16527;
  assign n29490 = pi190 & ~n29489;
  assign n29491 = ~pi190 & pi763;
  assign n29492 = n16514 & n29491;
  assign n29493 = ~n21243 & ~n29490;
  assign n29494 = ~n29492 & n29493;
  assign n29495 = ~n29488 & n29494;
  assign n29496 = ~pi38 & ~n29495;
  assign n29497 = pi763 & n16570;
  assign n29498 = pi38 & ~n29441;
  assign n29499 = ~n29497 & n29498;
  assign n29500 = ~n29496 & ~n29499;
  assign n29501 = n9829 & ~n29500;
  assign n29502 = ~n29440 & ~n29501;
  assign n29503 = ~n15777 & ~n29502;
  assign n29504 = n15777 & ~n29438;
  assign n29505 = ~n29503 & ~n29504;
  assign n29506 = ~pi785 & ~n29505;
  assign n29507 = ~n15786 & ~n29438;
  assign n29508 = pi609 & n29503;
  assign n29509 = ~n29507 & ~n29508;
  assign n29510 = pi1155 & ~n29509;
  assign n29511 = ~n16585 & ~n29438;
  assign n29512 = ~pi609 & n29503;
  assign n29513 = ~n29511 & ~n29512;
  assign n29514 = ~pi1155 & ~n29513;
  assign n29515 = ~n29510 & ~n29514;
  assign n29516 = pi785 & ~n29515;
  assign n29517 = ~n29506 & ~n29516;
  assign n29518 = ~pi781 & ~n29517;
  assign n29519 = ~pi618 & n29438;
  assign n29520 = pi618 & n29517;
  assign n29521 = pi1154 & ~n29519;
  assign n29522 = ~n29520 & n29521;
  assign n29523 = ~pi618 & n29517;
  assign n29524 = pi618 & n29438;
  assign n29525 = ~pi1154 & ~n29524;
  assign n29526 = ~n29523 & n29525;
  assign n29527 = ~n29522 & ~n29526;
  assign n29528 = pi781 & ~n29527;
  assign n29529 = ~n29518 & ~n29528;
  assign n29530 = ~pi789 & ~n29529;
  assign n29531 = ~pi619 & n29438;
  assign n29532 = pi619 & n29529;
  assign n29533 = pi1159 & ~n29531;
  assign n29534 = ~n29532 & n29533;
  assign n29535 = ~pi619 & n29529;
  assign n29536 = pi619 & n29438;
  assign n29537 = ~pi1159 & ~n29536;
  assign n29538 = ~n29535 & n29537;
  assign n29539 = ~n29534 & ~n29538;
  assign n29540 = pi789 & ~n29539;
  assign n29541 = ~n29530 & ~n29540;
  assign n29542 = ~n15832 & n29541;
  assign n29543 = n15832 & n29438;
  assign n29544 = ~n29542 & ~n29543;
  assign n29545 = ~n15925 & ~n29544;
  assign n29546 = n15925 & n29438;
  assign n29547 = ~n29545 & ~n29546;
  assign n29548 = ~n15960 & ~n29547;
  assign n29549 = n15960 & n29438;
  assign n29550 = ~n29548 & ~n29549;
  assign n29551 = pi644 & ~n29550;
  assign n29552 = ~pi644 & n29438;
  assign n29553 = ~pi715 & ~n29552;
  assign n29554 = ~n29551 & n29553;
  assign n29555 = pi1160 & ~n29484;
  assign n29556 = ~n29554 & n29555;
  assign n29557 = pi644 & ~n29482;
  assign n29558 = ~pi715 & ~n29557;
  assign n29559 = ~pi644 & ~n29550;
  assign n29560 = pi644 & n29438;
  assign n29561 = pi715 & ~n29560;
  assign n29562 = ~n29559 & n29561;
  assign n29563 = ~pi1160 & ~n29562;
  assign n29564 = ~n29558 & n29563;
  assign n29565 = ~n29556 & ~n29564;
  assign n29566 = pi790 & ~n29565;
  assign n29567 = ~pi647 & n29438;
  assign n29568 = pi647 & ~n29479;
  assign n29569 = n15957 & ~n29567;
  assign n29570 = ~n29568 & n29569;
  assign n29571 = n19478 & n29547;
  assign n29572 = pi647 & n29438;
  assign n29573 = ~pi647 & ~n29479;
  assign n29574 = n15958 & ~n29572;
  assign n29575 = ~n29573 & n29574;
  assign n29576 = ~n29570 & ~n29575;
  assign n29577 = ~n29571 & n29576;
  assign n29578 = pi787 & ~n29577;
  assign n29579 = pi628 & n29438;
  assign n29580 = ~pi628 & ~n29476;
  assign n29581 = n15923 & ~n29579;
  assign n29582 = ~n29580 & n29581;
  assign n29583 = ~n16633 & n29544;
  assign n29584 = ~pi628 & n29438;
  assign n29585 = pi628 & ~n29476;
  assign n29586 = n15922 & ~n29584;
  assign n29587 = ~n29585 & n29586;
  assign n29588 = ~n29582 & ~n29587;
  assign n29589 = ~n29583 & n29588;
  assign n29590 = pi792 & ~n29589;
  assign n29591 = n15828 & ~n29473;
  assign n29592 = ~pi626 & ~n29438;
  assign n29593 = pi626 & ~n29541;
  assign n29594 = n15756 & ~n29592;
  assign n29595 = ~n29593 & n29594;
  assign n29596 = pi626 & ~n29438;
  assign n29597 = ~pi626 & ~n29541;
  assign n29598 = n15757 & ~n29596;
  assign n29599 = ~n29597 & n29598;
  assign n29600 = ~n29591 & ~n29595;
  assign n29601 = ~n29599 & n29600;
  assign n29602 = pi788 & ~n29601;
  assign n29603 = pi618 & ~n29468;
  assign n29604 = pi609 & n29465;
  assign n29605 = ~pi699 & n29500;
  assign n29606 = ~n16921 & ~n29287;
  assign n29607 = pi190 & ~n29606;
  assign n29608 = n6081 & n29607;
  assign n29609 = ~pi763 & n22848;
  assign n29610 = ~n16808 & ~n29609;
  assign n29611 = ~pi39 & ~n29610;
  assign n29612 = ~pi190 & ~n29611;
  assign n29613 = pi38 & ~n29608;
  assign n29614 = ~n29612 & n29613;
  assign n29615 = ~pi190 & n16653;
  assign n29616 = pi190 & n16657;
  assign n29617 = ~pi763 & ~n29615;
  assign n29618 = ~n29616 & n29617;
  assign n29619 = ~pi190 & ~n16647;
  assign n29620 = pi190 & ~n17397;
  assign n29621 = pi763 & ~n29619;
  assign n29622 = ~n29620 & n29621;
  assign n29623 = ~pi39 & ~n29622;
  assign n29624 = ~n29618 & n29623;
  assign n29625 = ~pi190 & n16877;
  assign n29626 = pi190 & n16913;
  assign n29627 = pi763 & ~n29625;
  assign n29628 = ~n29626 & n29627;
  assign n29629 = pi190 & n16825;
  assign n29630 = ~pi190 & ~n16747;
  assign n29631 = ~pi763 & ~n29629;
  assign n29632 = ~n29630 & n29631;
  assign n29633 = pi39 & ~n29628;
  assign n29634 = ~n29632 & n29633;
  assign n29635 = ~pi38 & ~n29624;
  assign n29636 = ~n29634 & n29635;
  assign n29637 = pi699 & ~n29614;
  assign n29638 = ~n29636 & n29637;
  assign n29639 = n9829 & ~n29638;
  assign n29640 = ~n29605 & n29639;
  assign n29641 = ~n29440 & ~n29640;
  assign n29642 = ~pi625 & n29641;
  assign n29643 = pi625 & n29502;
  assign n29644 = ~pi1153 & ~n29643;
  assign n29645 = ~n29642 & n29644;
  assign n29646 = ~pi608 & ~n29458;
  assign n29647 = ~n29645 & n29646;
  assign n29648 = ~pi625 & n29502;
  assign n29649 = pi625 & n29641;
  assign n29650 = pi1153 & ~n29648;
  assign n29651 = ~n29649 & n29650;
  assign n29652 = pi608 & ~n29462;
  assign n29653 = ~n29651 & n29652;
  assign n29654 = ~n29647 & ~n29653;
  assign n29655 = pi778 & ~n29654;
  assign n29656 = ~pi778 & n29641;
  assign n29657 = ~n29655 & ~n29656;
  assign n29658 = ~pi609 & ~n29657;
  assign n29659 = ~pi1155 & ~n29604;
  assign n29660 = ~n29658 & n29659;
  assign n29661 = ~pi660 & ~n29510;
  assign n29662 = ~n29660 & n29661;
  assign n29663 = ~pi609 & n29465;
  assign n29664 = pi609 & ~n29657;
  assign n29665 = pi1155 & ~n29663;
  assign n29666 = ~n29664 & n29665;
  assign n29667 = pi660 & ~n29514;
  assign n29668 = ~n29666 & n29667;
  assign n29669 = ~n29662 & ~n29668;
  assign n29670 = pi785 & ~n29669;
  assign n29671 = ~pi785 & ~n29657;
  assign n29672 = ~n29670 & ~n29671;
  assign n29673 = ~pi618 & ~n29672;
  assign n29674 = ~pi1154 & ~n29603;
  assign n29675 = ~n29673 & n29674;
  assign n29676 = ~pi627 & ~n29522;
  assign n29677 = ~n29675 & n29676;
  assign n29678 = ~pi618 & ~n29468;
  assign n29679 = pi618 & ~n29672;
  assign n29680 = pi1154 & ~n29678;
  assign n29681 = ~n29679 & n29680;
  assign n29682 = pi627 & ~n29526;
  assign n29683 = ~n29681 & n29682;
  assign n29684 = ~n29677 & ~n29683;
  assign n29685 = pi781 & ~n29684;
  assign n29686 = ~pi781 & ~n29672;
  assign n29687 = ~n29685 & ~n29686;
  assign n29688 = ~pi789 & n29687;
  assign n29689 = ~pi619 & n29470;
  assign n29690 = pi619 & ~n29687;
  assign n29691 = pi1159 & ~n29689;
  assign n29692 = ~n29690 & n29691;
  assign n29693 = pi648 & ~n29538;
  assign n29694 = ~n29692 & n29693;
  assign n29695 = ~pi619 & ~n29687;
  assign n29696 = pi619 & n29470;
  assign n29697 = ~pi1159 & ~n29696;
  assign n29698 = ~n29695 & n29697;
  assign n29699 = ~pi648 & ~n29534;
  assign n29700 = ~n29698 & n29699;
  assign n29701 = pi789 & ~n29694;
  assign n29702 = ~n29700 & n29701;
  assign n29703 = n15833 & ~n29688;
  assign n29704 = ~n29702 & n29703;
  assign n29705 = ~n16644 & ~n29602;
  assign n29706 = ~n29704 & n29705;
  assign n29707 = ~n29590 & ~n29706;
  assign n29708 = n18841 & ~n29707;
  assign n29709 = pi644 & ~n29554;
  assign n29710 = ~n29563 & ~n29709;
  assign n29711 = ~n22949 & ~n29710;
  assign n29712 = pi790 & ~n29711;
  assign n29713 = ~n29578 & ~n29708;
  assign n29714 = ~n29712 & n29713;
  assign n29715 = ~n29566 & ~n29714;
  assign n29716 = ~po1038 & ~n29715;
  assign n29717 = ~pi832 & ~n29437;
  assign n29718 = ~n29716 & n29717;
  assign po347 = ~n29436 & ~n29718;
  assign n29720 = ~pi191 & ~n2923;
  assign n29721 = pi729 & n15726;
  assign n29722 = ~n29720 & ~n29721;
  assign n29723 = ~pi778 & ~n29722;
  assign n29724 = ~pi625 & n29721;
  assign n29725 = ~n29722 & ~n29724;
  assign n29726 = pi1153 & ~n29725;
  assign n29727 = ~pi1153 & ~n29720;
  assign n29728 = ~n29724 & n29727;
  assign n29729 = pi778 & ~n29728;
  assign n29730 = ~n29726 & n29729;
  assign n29731 = ~n29723 & ~n29730;
  assign n29732 = ~n15742 & ~n29731;
  assign n29733 = ~n15748 & n29732;
  assign n29734 = ~n15754 & n29733;
  assign n29735 = ~n15760 & n29734;
  assign n29736 = ~n15766 & n29735;
  assign n29737 = n19394 & n29736;
  assign n29738 = ~n19394 & n29720;
  assign n29739 = ~n29737 & ~n29738;
  assign n29740 = ~n15959 & n29739;
  assign n29741 = n15925 & n29720;
  assign n29742 = pi746 & n15781;
  assign n29743 = ~n29720 & ~n29742;
  assign n29744 = ~n15778 & ~n29743;
  assign n29745 = ~pi785 & ~n29744;
  assign n29746 = n16585 & n29742;
  assign n29747 = n29744 & ~n29746;
  assign n29748 = pi1155 & ~n29747;
  assign n29749 = ~pi1155 & ~n29720;
  assign n29750 = ~n29746 & n29749;
  assign n29751 = ~n29748 & ~n29750;
  assign n29752 = pi785 & ~n29751;
  assign n29753 = ~n29745 & ~n29752;
  assign n29754 = ~pi781 & ~n29753;
  assign n29755 = ~n15797 & n29753;
  assign n29756 = pi1154 & ~n29755;
  assign n29757 = ~n15800 & n29753;
  assign n29758 = ~pi1154 & ~n29757;
  assign n29759 = ~n29756 & ~n29758;
  assign n29760 = pi781 & ~n29759;
  assign n29761 = ~n29754 & ~n29760;
  assign n29762 = ~n21915 & n29761;
  assign n29763 = ~n15832 & ~n29762;
  assign n29764 = n15832 & ~n29720;
  assign n29765 = ~n29763 & ~n29764;
  assign n29766 = ~n15925 & n29765;
  assign n29767 = n19478 & ~n29741;
  assign n29768 = ~n29766 & n29767;
  assign n29769 = ~n29740 & ~n29768;
  assign n29770 = pi787 & ~n29769;
  assign n29771 = n15763 & n29765;
  assign n29772 = n15772 & n29735;
  assign n29773 = ~pi629 & ~n29772;
  assign n29774 = ~n29771 & n29773;
  assign n29775 = n15762 & n29765;
  assign n29776 = n15909 & n29735;
  assign n29777 = pi629 & ~n29776;
  assign n29778 = ~n29775 & n29777;
  assign n29779 = pi792 & ~n29774;
  assign n29780 = ~n29778 & n29779;
  assign n29781 = ~n21932 & n29761;
  assign n29782 = pi648 & ~n29781;
  assign n29783 = n21935 & ~n29733;
  assign n29784 = ~n29782 & ~n29783;
  assign n29785 = ~pi1159 & ~n29784;
  assign n29786 = ~pi619 & ~n29733;
  assign n29787 = pi648 & ~n29786;
  assign n29788 = n21942 & n29761;
  assign n29789 = pi1159 & ~n29787;
  assign n29790 = ~n29788 & n29789;
  assign n29791 = ~n29785 & ~n29790;
  assign n29792 = pi789 & ~n29791;
  assign n29793 = pi609 & ~n29731;
  assign n29794 = ~n15780 & ~n29722;
  assign n29795 = pi625 & n29794;
  assign n29796 = n29743 & ~n29794;
  assign n29797 = ~n29795 & ~n29796;
  assign n29798 = n29727 & ~n29797;
  assign n29799 = ~pi608 & ~n29726;
  assign n29800 = ~n29798 & n29799;
  assign n29801 = pi1153 & n29743;
  assign n29802 = ~n29795 & n29801;
  assign n29803 = pi608 & ~n29728;
  assign n29804 = ~n29802 & n29803;
  assign n29805 = ~n29800 & ~n29804;
  assign n29806 = pi778 & ~n29805;
  assign n29807 = ~pi778 & ~n29796;
  assign n29808 = ~n29806 & ~n29807;
  assign n29809 = ~pi609 & ~n29808;
  assign n29810 = ~pi1155 & ~n29793;
  assign n29811 = ~n29809 & n29810;
  assign n29812 = ~pi660 & ~n29748;
  assign n29813 = ~n29811 & n29812;
  assign n29814 = ~pi609 & ~n29731;
  assign n29815 = pi609 & ~n29808;
  assign n29816 = pi1155 & ~n29814;
  assign n29817 = ~n29815 & n29816;
  assign n29818 = pi660 & ~n29750;
  assign n29819 = ~n29817 & n29818;
  assign n29820 = ~n29813 & ~n29819;
  assign n29821 = pi785 & ~n29820;
  assign n29822 = ~pi785 & ~n29808;
  assign n29823 = ~n29821 & ~n29822;
  assign n29824 = ~pi781 & n29823;
  assign n29825 = pi618 & n29732;
  assign n29826 = ~pi618 & ~n29823;
  assign n29827 = ~pi1154 & ~n29825;
  assign n29828 = ~n29826 & n29827;
  assign n29829 = ~pi627 & ~n29756;
  assign n29830 = ~n29828 & n29829;
  assign n29831 = ~pi618 & n29732;
  assign n29832 = pi618 & ~n29823;
  assign n29833 = pi1154 & ~n29831;
  assign n29834 = ~n29832 & n29833;
  assign n29835 = pi627 & ~n29758;
  assign n29836 = ~n29834 & n29835;
  assign n29837 = pi781 & ~n29830;
  assign n29838 = ~n29836 & n29837;
  assign n29839 = ~n29792 & ~n29824;
  assign n29840 = ~n29838 & n29839;
  assign n29841 = n18969 & n29791;
  assign n29842 = ~n29840 & ~n29841;
  assign n29843 = n15833 & ~n29842;
  assign n29844 = n15828 & n29734;
  assign n29845 = ~pi626 & ~n29720;
  assign n29846 = pi626 & ~n29762;
  assign n29847 = n15756 & ~n29845;
  assign n29848 = ~n29846 & n29847;
  assign n29849 = pi626 & ~n29720;
  assign n29850 = ~pi626 & ~n29762;
  assign n29851 = n15757 & ~n29849;
  assign n29852 = ~n29850 & n29851;
  assign n29853 = ~n29844 & ~n29848;
  assign n29854 = ~n29852 & n29853;
  assign n29855 = pi788 & ~n29854;
  assign n29856 = ~n29843 & ~n29855;
  assign n29857 = ~n16644 & ~n29856;
  assign n29858 = n18841 & ~n29780;
  assign n29859 = ~n29857 & n29858;
  assign n29860 = ~n29770 & ~n29859;
  assign n29861 = ~pi790 & n29860;
  assign n29862 = pi787 & ~n29739;
  assign n29863 = ~pi787 & n29736;
  assign n29864 = ~n29862 & ~n29863;
  assign n29865 = ~pi644 & ~n29864;
  assign n29866 = pi644 & n29860;
  assign n29867 = pi715 & ~n29865;
  assign n29868 = ~n29866 & n29867;
  assign n29869 = ~n19771 & n29720;
  assign n29870 = ~n15960 & n29766;
  assign n29871 = ~n29869 & ~n29870;
  assign n29872 = pi644 & ~n29871;
  assign n29873 = ~pi644 & n29720;
  assign n29874 = ~pi715 & ~n29873;
  assign n29875 = ~n29872 & n29874;
  assign n29876 = pi1160 & ~n29875;
  assign n29877 = ~n29868 & n29876;
  assign n29878 = ~pi644 & ~n29871;
  assign n29879 = pi644 & n29720;
  assign n29880 = pi715 & ~n29879;
  assign n29881 = ~n29878 & n29880;
  assign n29882 = pi644 & ~n29864;
  assign n29883 = ~pi644 & n29860;
  assign n29884 = ~pi715 & ~n29882;
  assign n29885 = ~n29883 & n29884;
  assign n29886 = ~pi1160 & ~n29881;
  assign n29887 = ~n29885 & n29886;
  assign n29888 = ~n29877 & ~n29887;
  assign n29889 = pi790 & ~n29888;
  assign n29890 = pi832 & ~n29861;
  assign n29891 = ~n29889 & n29890;
  assign n29892 = ~pi191 & po1038;
  assign n29893 = ~pi191 & ~n16219;
  assign n29894 = n15747 & ~n29893;
  assign n29895 = pi191 & ~n9829;
  assign n29896 = ~pi191 & ~n16228;
  assign n29897 = n16227 & ~n29896;
  assign n29898 = pi191 & n17272;
  assign n29899 = ~pi191 & ~n17276;
  assign n29900 = ~pi38 & ~n29898;
  assign n29901 = ~n29899 & n29900;
  assign n29902 = pi729 & ~n29897;
  assign n29903 = ~n29901 & n29902;
  assign n29904 = ~pi191 & ~pi729;
  assign n29905 = ~n16218 & n29904;
  assign n29906 = n9829 & ~n29903;
  assign n29907 = ~n29905 & n29906;
  assign n29908 = ~n29895 & ~n29907;
  assign n29909 = ~pi778 & ~n29908;
  assign n29910 = ~pi625 & n29893;
  assign n29911 = pi625 & n29908;
  assign n29912 = pi1153 & ~n29910;
  assign n29913 = ~n29911 & n29912;
  assign n29914 = ~pi625 & n29908;
  assign n29915 = pi625 & n29893;
  assign n29916 = ~pi1153 & ~n29915;
  assign n29917 = ~n29914 & n29916;
  assign n29918 = ~n29913 & ~n29917;
  assign n29919 = pi778 & ~n29918;
  assign n29920 = ~n29909 & ~n29919;
  assign n29921 = ~n15741 & n29920;
  assign n29922 = n15741 & n29893;
  assign n29923 = ~n29921 & ~n29922;
  assign n29924 = ~n15747 & n29923;
  assign n29925 = ~n29894 & ~n29924;
  assign n29926 = ~n15753 & n29925;
  assign n29927 = n15753 & n29893;
  assign n29928 = ~n29926 & ~n29927;
  assign n29929 = ~n15759 & ~n29928;
  assign n29930 = n15759 & n29893;
  assign n29931 = ~n29929 & ~n29930;
  assign n29932 = ~n15765 & ~n29931;
  assign n29933 = n15765 & n29893;
  assign n29934 = ~n29932 & ~n29933;
  assign n29935 = ~n17768 & ~n29934;
  assign n29936 = n17768 & n29893;
  assign n29937 = ~n29935 & ~n29936;
  assign n29938 = ~pi644 & ~n29937;
  assign n29939 = pi715 & ~n29938;
  assign n29940 = ~pi746 & n16212;
  assign n29941 = pi191 & ~n16563;
  assign n29942 = ~n29940 & ~n29941;
  assign n29943 = pi39 & ~n29942;
  assign n29944 = pi746 & ~n16527;
  assign n29945 = pi191 & ~n29944;
  assign n29946 = ~pi191 & pi746;
  assign n29947 = n16514 & n29946;
  assign n29948 = ~n21322 & ~n29945;
  assign n29949 = ~n29947 & n29948;
  assign n29950 = ~n29943 & n29949;
  assign n29951 = ~pi38 & ~n29950;
  assign n29952 = pi746 & n16570;
  assign n29953 = pi38 & ~n29896;
  assign n29954 = ~n29952 & n29953;
  assign n29955 = ~n29951 & ~n29954;
  assign n29956 = n9829 & ~n29955;
  assign n29957 = ~n29895 & ~n29956;
  assign n29958 = ~n15777 & ~n29957;
  assign n29959 = n15777 & ~n29893;
  assign n29960 = ~n29958 & ~n29959;
  assign n29961 = ~pi785 & ~n29960;
  assign n29962 = ~n15786 & ~n29893;
  assign n29963 = pi609 & n29958;
  assign n29964 = ~n29962 & ~n29963;
  assign n29965 = pi1155 & ~n29964;
  assign n29966 = ~n16585 & ~n29893;
  assign n29967 = ~pi609 & n29958;
  assign n29968 = ~n29966 & ~n29967;
  assign n29969 = ~pi1155 & ~n29968;
  assign n29970 = ~n29965 & ~n29969;
  assign n29971 = pi785 & ~n29970;
  assign n29972 = ~n29961 & ~n29971;
  assign n29973 = ~pi781 & ~n29972;
  assign n29974 = ~pi618 & n29893;
  assign n29975 = pi618 & n29972;
  assign n29976 = pi1154 & ~n29974;
  assign n29977 = ~n29975 & n29976;
  assign n29978 = ~pi618 & n29972;
  assign n29979 = pi618 & n29893;
  assign n29980 = ~pi1154 & ~n29979;
  assign n29981 = ~n29978 & n29980;
  assign n29982 = ~n29977 & ~n29981;
  assign n29983 = pi781 & ~n29982;
  assign n29984 = ~n29973 & ~n29983;
  assign n29985 = ~pi789 & ~n29984;
  assign n29986 = ~pi619 & n29893;
  assign n29987 = pi619 & n29984;
  assign n29988 = pi1159 & ~n29986;
  assign n29989 = ~n29987 & n29988;
  assign n29990 = ~pi619 & n29984;
  assign n29991 = pi619 & n29893;
  assign n29992 = ~pi1159 & ~n29991;
  assign n29993 = ~n29990 & n29992;
  assign n29994 = ~n29989 & ~n29993;
  assign n29995 = pi789 & ~n29994;
  assign n29996 = ~n29985 & ~n29995;
  assign n29997 = ~n15832 & n29996;
  assign n29998 = n15832 & n29893;
  assign n29999 = ~n29997 & ~n29998;
  assign n30000 = ~n15925 & ~n29999;
  assign n30001 = n15925 & n29893;
  assign n30002 = ~n30000 & ~n30001;
  assign n30003 = ~n15960 & ~n30002;
  assign n30004 = n15960 & n29893;
  assign n30005 = ~n30003 & ~n30004;
  assign n30006 = pi644 & ~n30005;
  assign n30007 = ~pi644 & n29893;
  assign n30008 = ~pi715 & ~n30007;
  assign n30009 = ~n30006 & n30008;
  assign n30010 = pi1160 & ~n29939;
  assign n30011 = ~n30009 & n30010;
  assign n30012 = pi644 & ~n29937;
  assign n30013 = ~pi715 & ~n30012;
  assign n30014 = ~pi644 & ~n30005;
  assign n30015 = pi644 & n29893;
  assign n30016 = pi715 & ~n30015;
  assign n30017 = ~n30014 & n30016;
  assign n30018 = ~pi1160 & ~n30017;
  assign n30019 = ~n30013 & n30018;
  assign n30020 = ~n30011 & ~n30019;
  assign n30021 = pi790 & ~n30020;
  assign n30022 = ~pi647 & n29893;
  assign n30023 = pi647 & ~n29934;
  assign n30024 = n15957 & ~n30022;
  assign n30025 = ~n30023 & n30024;
  assign n30026 = n19478 & n30002;
  assign n30027 = pi647 & n29893;
  assign n30028 = ~pi647 & ~n29934;
  assign n30029 = n15958 & ~n30027;
  assign n30030 = ~n30028 & n30029;
  assign n30031 = ~n30025 & ~n30030;
  assign n30032 = ~n30026 & n30031;
  assign n30033 = pi787 & ~n30032;
  assign n30034 = pi628 & n29893;
  assign n30035 = ~pi628 & ~n29931;
  assign n30036 = n15923 & ~n30034;
  assign n30037 = ~n30035 & n30036;
  assign n30038 = ~n16633 & n29999;
  assign n30039 = ~pi628 & n29893;
  assign n30040 = pi628 & ~n29931;
  assign n30041 = n15922 & ~n30039;
  assign n30042 = ~n30040 & n30041;
  assign n30043 = ~n30037 & ~n30042;
  assign n30044 = ~n30038 & n30043;
  assign n30045 = pi792 & ~n30044;
  assign n30046 = n15828 & ~n29928;
  assign n30047 = ~pi626 & ~n29893;
  assign n30048 = pi626 & ~n29996;
  assign n30049 = n15756 & ~n30047;
  assign n30050 = ~n30048 & n30049;
  assign n30051 = pi626 & ~n29893;
  assign n30052 = ~pi626 & ~n29996;
  assign n30053 = n15757 & ~n30051;
  assign n30054 = ~n30052 & n30053;
  assign n30055 = ~n30046 & ~n30050;
  assign n30056 = ~n30054 & n30055;
  assign n30057 = pi788 & ~n30056;
  assign n30058 = pi618 & ~n29923;
  assign n30059 = pi609 & n29920;
  assign n30060 = ~pi729 & n29955;
  assign n30061 = ~n16921 & ~n29742;
  assign n30062 = pi191 & ~n30061;
  assign n30063 = n6081 & n30062;
  assign n30064 = ~pi746 & n22848;
  assign n30065 = ~n16808 & ~n30064;
  assign n30066 = ~pi39 & ~n30065;
  assign n30067 = ~pi191 & ~n30066;
  assign n30068 = pi38 & ~n30063;
  assign n30069 = ~n30067 & n30068;
  assign n30070 = ~pi191 & n16653;
  assign n30071 = pi191 & n16657;
  assign n30072 = ~pi746 & ~n30070;
  assign n30073 = ~n30071 & n30072;
  assign n30074 = ~pi191 & ~n16647;
  assign n30075 = pi191 & ~n17397;
  assign n30076 = pi746 & ~n30074;
  assign n30077 = ~n30075 & n30076;
  assign n30078 = ~pi39 & ~n30077;
  assign n30079 = ~n30073 & n30078;
  assign n30080 = ~pi191 & n16877;
  assign n30081 = pi191 & n16913;
  assign n30082 = pi746 & ~n30080;
  assign n30083 = ~n30081 & n30082;
  assign n30084 = pi191 & n16825;
  assign n30085 = ~pi191 & ~n16747;
  assign n30086 = ~pi746 & ~n30084;
  assign n30087 = ~n30085 & n30086;
  assign n30088 = pi39 & ~n30083;
  assign n30089 = ~n30087 & n30088;
  assign n30090 = ~pi38 & ~n30079;
  assign n30091 = ~n30089 & n30090;
  assign n30092 = pi729 & ~n30069;
  assign n30093 = ~n30091 & n30092;
  assign n30094 = n9829 & ~n30093;
  assign n30095 = ~n30060 & n30094;
  assign n30096 = ~n29895 & ~n30095;
  assign n30097 = ~pi625 & n30096;
  assign n30098 = pi625 & n29957;
  assign n30099 = ~pi1153 & ~n30098;
  assign n30100 = ~n30097 & n30099;
  assign n30101 = ~pi608 & ~n29913;
  assign n30102 = ~n30100 & n30101;
  assign n30103 = ~pi625 & n29957;
  assign n30104 = pi625 & n30096;
  assign n30105 = pi1153 & ~n30103;
  assign n30106 = ~n30104 & n30105;
  assign n30107 = pi608 & ~n29917;
  assign n30108 = ~n30106 & n30107;
  assign n30109 = ~n30102 & ~n30108;
  assign n30110 = pi778 & ~n30109;
  assign n30111 = ~pi778 & n30096;
  assign n30112 = ~n30110 & ~n30111;
  assign n30113 = ~pi609 & ~n30112;
  assign n30114 = ~pi1155 & ~n30059;
  assign n30115 = ~n30113 & n30114;
  assign n30116 = ~pi660 & ~n29965;
  assign n30117 = ~n30115 & n30116;
  assign n30118 = ~pi609 & n29920;
  assign n30119 = pi609 & ~n30112;
  assign n30120 = pi1155 & ~n30118;
  assign n30121 = ~n30119 & n30120;
  assign n30122 = pi660 & ~n29969;
  assign n30123 = ~n30121 & n30122;
  assign n30124 = ~n30117 & ~n30123;
  assign n30125 = pi785 & ~n30124;
  assign n30126 = ~pi785 & ~n30112;
  assign n30127 = ~n30125 & ~n30126;
  assign n30128 = ~pi618 & ~n30127;
  assign n30129 = ~pi1154 & ~n30058;
  assign n30130 = ~n30128 & n30129;
  assign n30131 = ~pi627 & ~n29977;
  assign n30132 = ~n30130 & n30131;
  assign n30133 = ~pi618 & ~n29923;
  assign n30134 = pi618 & ~n30127;
  assign n30135 = pi1154 & ~n30133;
  assign n30136 = ~n30134 & n30135;
  assign n30137 = pi627 & ~n29981;
  assign n30138 = ~n30136 & n30137;
  assign n30139 = ~n30132 & ~n30138;
  assign n30140 = pi781 & ~n30139;
  assign n30141 = ~pi781 & ~n30127;
  assign n30142 = ~n30140 & ~n30141;
  assign n30143 = ~pi789 & n30142;
  assign n30144 = ~pi619 & n29925;
  assign n30145 = pi619 & ~n30142;
  assign n30146 = pi1159 & ~n30144;
  assign n30147 = ~n30145 & n30146;
  assign n30148 = pi648 & ~n29993;
  assign n30149 = ~n30147 & n30148;
  assign n30150 = ~pi619 & ~n30142;
  assign n30151 = pi619 & n29925;
  assign n30152 = ~pi1159 & ~n30151;
  assign n30153 = ~n30150 & n30152;
  assign n30154 = ~pi648 & ~n29989;
  assign n30155 = ~n30153 & n30154;
  assign n30156 = pi789 & ~n30149;
  assign n30157 = ~n30155 & n30156;
  assign n30158 = n15833 & ~n30143;
  assign n30159 = ~n30157 & n30158;
  assign n30160 = ~n16644 & ~n30057;
  assign n30161 = ~n30159 & n30160;
  assign n30162 = ~n30045 & ~n30161;
  assign n30163 = n18841 & ~n30162;
  assign n30164 = pi644 & ~n30009;
  assign n30165 = ~n30018 & ~n30164;
  assign n30166 = ~n22949 & ~n30165;
  assign n30167 = pi790 & ~n30166;
  assign n30168 = ~n30033 & ~n30163;
  assign n30169 = ~n30167 & n30168;
  assign n30170 = ~n30021 & ~n30169;
  assign n30171 = ~po1038 & ~n30170;
  assign n30172 = ~pi832 & ~n29892;
  assign n30173 = ~n30171 & n30172;
  assign po348 = ~n29891 & ~n30173;
  assign n30175 = ~pi192 & ~n2923;
  assign n30176 = pi691 & n15726;
  assign n30177 = ~n30175 & ~n30176;
  assign n30178 = ~pi778 & ~n30177;
  assign n30179 = ~pi625 & n30176;
  assign n30180 = ~n30177 & ~n30179;
  assign n30181 = pi1153 & ~n30180;
  assign n30182 = ~pi1153 & ~n30175;
  assign n30183 = ~n30179 & n30182;
  assign n30184 = pi778 & ~n30183;
  assign n30185 = ~n30181 & n30184;
  assign n30186 = ~n30178 & ~n30185;
  assign n30187 = ~n15742 & ~n30186;
  assign n30188 = ~n15748 & n30187;
  assign n30189 = ~n15754 & n30188;
  assign n30190 = ~n15760 & n30189;
  assign n30191 = ~n15766 & n30190;
  assign n30192 = n19394 & n30191;
  assign n30193 = ~n19394 & n30175;
  assign n30194 = ~n30192 & ~n30193;
  assign n30195 = ~n15959 & n30194;
  assign n30196 = n15925 & n30175;
  assign n30197 = pi764 & n15781;
  assign n30198 = ~n30175 & ~n30197;
  assign n30199 = ~n15778 & ~n30198;
  assign n30200 = ~pi785 & ~n30199;
  assign n30201 = n16585 & n30197;
  assign n30202 = n30199 & ~n30201;
  assign n30203 = pi1155 & ~n30202;
  assign n30204 = ~pi1155 & ~n30175;
  assign n30205 = ~n30201 & n30204;
  assign n30206 = ~n30203 & ~n30205;
  assign n30207 = pi785 & ~n30206;
  assign n30208 = ~n30200 & ~n30207;
  assign n30209 = ~pi781 & ~n30208;
  assign n30210 = ~n15797 & n30208;
  assign n30211 = pi1154 & ~n30210;
  assign n30212 = ~n15800 & n30208;
  assign n30213 = ~pi1154 & ~n30212;
  assign n30214 = ~n30211 & ~n30213;
  assign n30215 = pi781 & ~n30214;
  assign n30216 = ~n30209 & ~n30215;
  assign n30217 = ~n21915 & n30216;
  assign n30218 = ~n15832 & ~n30217;
  assign n30219 = n15832 & ~n30175;
  assign n30220 = ~n30218 & ~n30219;
  assign n30221 = ~n15925 & n30220;
  assign n30222 = n19478 & ~n30196;
  assign n30223 = ~n30221 & n30222;
  assign n30224 = ~n30195 & ~n30223;
  assign n30225 = pi787 & ~n30224;
  assign n30226 = n15763 & n30220;
  assign n30227 = n15772 & n30190;
  assign n30228 = ~pi629 & ~n30227;
  assign n30229 = ~n30226 & n30228;
  assign n30230 = n15762 & n30220;
  assign n30231 = n15909 & n30190;
  assign n30232 = pi629 & ~n30231;
  assign n30233 = ~n30230 & n30232;
  assign n30234 = pi792 & ~n30229;
  assign n30235 = ~n30233 & n30234;
  assign n30236 = ~n21932 & n30216;
  assign n30237 = pi648 & ~n30236;
  assign n30238 = n21935 & ~n30188;
  assign n30239 = ~n30237 & ~n30238;
  assign n30240 = ~pi1159 & ~n30239;
  assign n30241 = ~pi619 & ~n30188;
  assign n30242 = pi648 & ~n30241;
  assign n30243 = n21942 & n30216;
  assign n30244 = pi1159 & ~n30242;
  assign n30245 = ~n30243 & n30244;
  assign n30246 = ~n30240 & ~n30245;
  assign n30247 = pi789 & ~n30246;
  assign n30248 = pi609 & ~n30186;
  assign n30249 = ~n15780 & ~n30177;
  assign n30250 = pi625 & n30249;
  assign n30251 = n30198 & ~n30249;
  assign n30252 = ~n30250 & ~n30251;
  assign n30253 = n30182 & ~n30252;
  assign n30254 = ~pi608 & ~n30181;
  assign n30255 = ~n30253 & n30254;
  assign n30256 = pi1153 & n30198;
  assign n30257 = ~n30250 & n30256;
  assign n30258 = pi608 & ~n30183;
  assign n30259 = ~n30257 & n30258;
  assign n30260 = ~n30255 & ~n30259;
  assign n30261 = pi778 & ~n30260;
  assign n30262 = ~pi778 & ~n30251;
  assign n30263 = ~n30261 & ~n30262;
  assign n30264 = ~pi609 & ~n30263;
  assign n30265 = ~pi1155 & ~n30248;
  assign n30266 = ~n30264 & n30265;
  assign n30267 = ~pi660 & ~n30203;
  assign n30268 = ~n30266 & n30267;
  assign n30269 = ~pi609 & ~n30186;
  assign n30270 = pi609 & ~n30263;
  assign n30271 = pi1155 & ~n30269;
  assign n30272 = ~n30270 & n30271;
  assign n30273 = pi660 & ~n30205;
  assign n30274 = ~n30272 & n30273;
  assign n30275 = ~n30268 & ~n30274;
  assign n30276 = pi785 & ~n30275;
  assign n30277 = ~pi785 & ~n30263;
  assign n30278 = ~n30276 & ~n30277;
  assign n30279 = ~pi781 & n30278;
  assign n30280 = pi618 & n30187;
  assign n30281 = ~pi618 & ~n30278;
  assign n30282 = ~pi1154 & ~n30280;
  assign n30283 = ~n30281 & n30282;
  assign n30284 = ~pi627 & ~n30211;
  assign n30285 = ~n30283 & n30284;
  assign n30286 = ~pi618 & n30187;
  assign n30287 = pi618 & ~n30278;
  assign n30288 = pi1154 & ~n30286;
  assign n30289 = ~n30287 & n30288;
  assign n30290 = pi627 & ~n30213;
  assign n30291 = ~n30289 & n30290;
  assign n30292 = pi781 & ~n30285;
  assign n30293 = ~n30291 & n30292;
  assign n30294 = ~n30247 & ~n30279;
  assign n30295 = ~n30293 & n30294;
  assign n30296 = n18969 & n30246;
  assign n30297 = ~n30295 & ~n30296;
  assign n30298 = n15833 & ~n30297;
  assign n30299 = n15828 & n30189;
  assign n30300 = ~pi626 & ~n30175;
  assign n30301 = pi626 & ~n30217;
  assign n30302 = n15756 & ~n30300;
  assign n30303 = ~n30301 & n30302;
  assign n30304 = pi626 & ~n30175;
  assign n30305 = ~pi626 & ~n30217;
  assign n30306 = n15757 & ~n30304;
  assign n30307 = ~n30305 & n30306;
  assign n30308 = ~n30299 & ~n30303;
  assign n30309 = ~n30307 & n30308;
  assign n30310 = pi788 & ~n30309;
  assign n30311 = ~n30298 & ~n30310;
  assign n30312 = ~n16644 & ~n30311;
  assign n30313 = n18841 & ~n30235;
  assign n30314 = ~n30312 & n30313;
  assign n30315 = ~n30225 & ~n30314;
  assign n30316 = ~pi790 & n30315;
  assign n30317 = pi787 & ~n30194;
  assign n30318 = ~pi787 & n30191;
  assign n30319 = ~n30317 & ~n30318;
  assign n30320 = ~pi644 & ~n30319;
  assign n30321 = pi644 & n30315;
  assign n30322 = pi715 & ~n30320;
  assign n30323 = ~n30321 & n30322;
  assign n30324 = ~n19771 & n30175;
  assign n30325 = ~n15960 & n30221;
  assign n30326 = ~n30324 & ~n30325;
  assign n30327 = pi644 & ~n30326;
  assign n30328 = ~pi644 & n30175;
  assign n30329 = ~pi715 & ~n30328;
  assign n30330 = ~n30327 & n30329;
  assign n30331 = pi1160 & ~n30330;
  assign n30332 = ~n30323 & n30331;
  assign n30333 = ~pi644 & ~n30326;
  assign n30334 = pi644 & n30175;
  assign n30335 = pi715 & ~n30334;
  assign n30336 = ~n30333 & n30335;
  assign n30337 = pi644 & ~n30319;
  assign n30338 = ~pi644 & n30315;
  assign n30339 = ~pi715 & ~n30337;
  assign n30340 = ~n30338 & n30339;
  assign n30341 = ~pi1160 & ~n30336;
  assign n30342 = ~n30340 & n30341;
  assign n30343 = ~n30332 & ~n30342;
  assign n30344 = pi790 & ~n30343;
  assign n30345 = pi832 & ~n30316;
  assign n30346 = ~n30344 & n30345;
  assign n30347 = ~pi192 & po1038;
  assign n30348 = ~pi192 & ~n16219;
  assign n30349 = n15747 & ~n30348;
  assign n30350 = pi192 & ~n9829;
  assign n30351 = ~pi192 & ~n16228;
  assign n30352 = n16227 & ~n30351;
  assign n30353 = pi192 & n17272;
  assign n30354 = ~pi192 & ~n17276;
  assign n30355 = ~pi38 & ~n30353;
  assign n30356 = ~n30354 & n30355;
  assign n30357 = pi691 & ~n30352;
  assign n30358 = ~n30356 & n30357;
  assign n30359 = ~pi192 & ~pi691;
  assign n30360 = ~n16218 & n30359;
  assign n30361 = n9829 & ~n30358;
  assign n30362 = ~n30360 & n30361;
  assign n30363 = ~n30350 & ~n30362;
  assign n30364 = ~pi778 & ~n30363;
  assign n30365 = ~pi625 & n30348;
  assign n30366 = pi625 & n30363;
  assign n30367 = pi1153 & ~n30365;
  assign n30368 = ~n30366 & n30367;
  assign n30369 = ~pi625 & n30363;
  assign n30370 = pi625 & n30348;
  assign n30371 = ~pi1153 & ~n30370;
  assign n30372 = ~n30369 & n30371;
  assign n30373 = ~n30368 & ~n30372;
  assign n30374 = pi778 & ~n30373;
  assign n30375 = ~n30364 & ~n30374;
  assign n30376 = ~n15741 & n30375;
  assign n30377 = n15741 & n30348;
  assign n30378 = ~n30376 & ~n30377;
  assign n30379 = ~n15747 & n30378;
  assign n30380 = ~n30349 & ~n30379;
  assign n30381 = ~n15753 & n30380;
  assign n30382 = n15753 & n30348;
  assign n30383 = ~n30381 & ~n30382;
  assign n30384 = ~n15759 & ~n30383;
  assign n30385 = n15759 & n30348;
  assign n30386 = ~n30384 & ~n30385;
  assign n30387 = ~n15765 & ~n30386;
  assign n30388 = n15765 & n30348;
  assign n30389 = ~n30387 & ~n30388;
  assign n30390 = ~n17768 & ~n30389;
  assign n30391 = n17768 & n30348;
  assign n30392 = ~n30390 & ~n30391;
  assign n30393 = ~pi644 & ~n30392;
  assign n30394 = pi715 & ~n30393;
  assign n30395 = ~pi764 & n16212;
  assign n30396 = pi192 & ~n16563;
  assign n30397 = ~n30395 & ~n30396;
  assign n30398 = pi39 & ~n30397;
  assign n30399 = pi764 & ~n16527;
  assign n30400 = pi192 & ~n30399;
  assign n30401 = ~pi192 & pi764;
  assign n30402 = n16514 & n30401;
  assign n30403 = ~n21480 & ~n30400;
  assign n30404 = ~n30402 & n30403;
  assign n30405 = ~n30398 & n30404;
  assign n30406 = ~pi38 & ~n30405;
  assign n30407 = pi764 & n16570;
  assign n30408 = pi38 & ~n30351;
  assign n30409 = ~n30407 & n30408;
  assign n30410 = ~n30406 & ~n30409;
  assign n30411 = n9829 & ~n30410;
  assign n30412 = ~n30350 & ~n30411;
  assign n30413 = ~n15777 & ~n30412;
  assign n30414 = n15777 & ~n30348;
  assign n30415 = ~n30413 & ~n30414;
  assign n30416 = ~pi785 & ~n30415;
  assign n30417 = ~n15786 & ~n30348;
  assign n30418 = pi609 & n30413;
  assign n30419 = ~n30417 & ~n30418;
  assign n30420 = pi1155 & ~n30419;
  assign n30421 = ~n16585 & ~n30348;
  assign n30422 = ~pi609 & n30413;
  assign n30423 = ~n30421 & ~n30422;
  assign n30424 = ~pi1155 & ~n30423;
  assign n30425 = ~n30420 & ~n30424;
  assign n30426 = pi785 & ~n30425;
  assign n30427 = ~n30416 & ~n30426;
  assign n30428 = ~pi781 & ~n30427;
  assign n30429 = ~pi618 & n30348;
  assign n30430 = pi618 & n30427;
  assign n30431 = pi1154 & ~n30429;
  assign n30432 = ~n30430 & n30431;
  assign n30433 = ~pi618 & n30427;
  assign n30434 = pi618 & n30348;
  assign n30435 = ~pi1154 & ~n30434;
  assign n30436 = ~n30433 & n30435;
  assign n30437 = ~n30432 & ~n30436;
  assign n30438 = pi781 & ~n30437;
  assign n30439 = ~n30428 & ~n30438;
  assign n30440 = ~pi789 & ~n30439;
  assign n30441 = ~pi619 & n30348;
  assign n30442 = pi619 & n30439;
  assign n30443 = pi1159 & ~n30441;
  assign n30444 = ~n30442 & n30443;
  assign n30445 = ~pi619 & n30439;
  assign n30446 = pi619 & n30348;
  assign n30447 = ~pi1159 & ~n30446;
  assign n30448 = ~n30445 & n30447;
  assign n30449 = ~n30444 & ~n30448;
  assign n30450 = pi789 & ~n30449;
  assign n30451 = ~n30440 & ~n30450;
  assign n30452 = ~n15832 & n30451;
  assign n30453 = n15832 & n30348;
  assign n30454 = ~n30452 & ~n30453;
  assign n30455 = ~n15925 & ~n30454;
  assign n30456 = n15925 & n30348;
  assign n30457 = ~n30455 & ~n30456;
  assign n30458 = ~n15960 & ~n30457;
  assign n30459 = n15960 & n30348;
  assign n30460 = ~n30458 & ~n30459;
  assign n30461 = pi644 & ~n30460;
  assign n30462 = ~pi644 & n30348;
  assign n30463 = ~pi715 & ~n30462;
  assign n30464 = ~n30461 & n30463;
  assign n30465 = pi1160 & ~n30394;
  assign n30466 = ~n30464 & n30465;
  assign n30467 = pi644 & ~n30392;
  assign n30468 = ~pi715 & ~n30467;
  assign n30469 = ~pi644 & ~n30460;
  assign n30470 = pi644 & n30348;
  assign n30471 = pi715 & ~n30470;
  assign n30472 = ~n30469 & n30471;
  assign n30473 = ~pi1160 & ~n30472;
  assign n30474 = ~n30468 & n30473;
  assign n30475 = ~n30466 & ~n30474;
  assign n30476 = pi790 & ~n30475;
  assign n30477 = ~pi647 & n30348;
  assign n30478 = pi647 & ~n30389;
  assign n30479 = n15957 & ~n30477;
  assign n30480 = ~n30478 & n30479;
  assign n30481 = n19478 & n30457;
  assign n30482 = pi647 & n30348;
  assign n30483 = ~pi647 & ~n30389;
  assign n30484 = n15958 & ~n30482;
  assign n30485 = ~n30483 & n30484;
  assign n30486 = ~n30480 & ~n30485;
  assign n30487 = ~n30481 & n30486;
  assign n30488 = pi787 & ~n30487;
  assign n30489 = pi628 & n30348;
  assign n30490 = ~pi628 & ~n30386;
  assign n30491 = n15923 & ~n30489;
  assign n30492 = ~n30490 & n30491;
  assign n30493 = ~n16633 & n30454;
  assign n30494 = ~pi628 & n30348;
  assign n30495 = pi628 & ~n30386;
  assign n30496 = n15922 & ~n30494;
  assign n30497 = ~n30495 & n30496;
  assign n30498 = ~n30492 & ~n30497;
  assign n30499 = ~n30493 & n30498;
  assign n30500 = pi792 & ~n30499;
  assign n30501 = n15828 & ~n30383;
  assign n30502 = ~pi626 & ~n30348;
  assign n30503 = pi626 & ~n30451;
  assign n30504 = n15756 & ~n30502;
  assign n30505 = ~n30503 & n30504;
  assign n30506 = pi626 & ~n30348;
  assign n30507 = ~pi626 & ~n30451;
  assign n30508 = n15757 & ~n30506;
  assign n30509 = ~n30507 & n30508;
  assign n30510 = ~n30501 & ~n30505;
  assign n30511 = ~n30509 & n30510;
  assign n30512 = pi788 & ~n30511;
  assign n30513 = pi618 & ~n30378;
  assign n30514 = pi609 & n30375;
  assign n30515 = ~pi691 & n30410;
  assign n30516 = ~n16921 & ~n30197;
  assign n30517 = pi192 & ~n30516;
  assign n30518 = n6081 & n30517;
  assign n30519 = ~pi764 & n22848;
  assign n30520 = ~n16808 & ~n30519;
  assign n30521 = ~pi39 & ~n30520;
  assign n30522 = ~pi192 & ~n30521;
  assign n30523 = pi38 & ~n30518;
  assign n30524 = ~n30522 & n30523;
  assign n30525 = ~pi192 & n16653;
  assign n30526 = pi192 & n16657;
  assign n30527 = ~pi764 & ~n30525;
  assign n30528 = ~n30526 & n30527;
  assign n30529 = ~pi192 & ~n16647;
  assign n30530 = pi192 & ~n17397;
  assign n30531 = pi764 & ~n30529;
  assign n30532 = ~n30530 & n30531;
  assign n30533 = ~pi39 & ~n30532;
  assign n30534 = ~n30528 & n30533;
  assign n30535 = ~pi192 & n16877;
  assign n30536 = pi192 & n16913;
  assign n30537 = pi764 & ~n30535;
  assign n30538 = ~n30536 & n30537;
  assign n30539 = pi192 & n16825;
  assign n30540 = ~pi192 & ~n16747;
  assign n30541 = ~pi764 & ~n30539;
  assign n30542 = ~n30540 & n30541;
  assign n30543 = pi39 & ~n30538;
  assign n30544 = ~n30542 & n30543;
  assign n30545 = ~pi38 & ~n30534;
  assign n30546 = ~n30544 & n30545;
  assign n30547 = pi691 & ~n30524;
  assign n30548 = ~n30546 & n30547;
  assign n30549 = n9829 & ~n30548;
  assign n30550 = ~n30515 & n30549;
  assign n30551 = ~n30350 & ~n30550;
  assign n30552 = ~pi625 & n30551;
  assign n30553 = pi625 & n30412;
  assign n30554 = ~pi1153 & ~n30553;
  assign n30555 = ~n30552 & n30554;
  assign n30556 = ~pi608 & ~n30368;
  assign n30557 = ~n30555 & n30556;
  assign n30558 = ~pi625 & n30412;
  assign n30559 = pi625 & n30551;
  assign n30560 = pi1153 & ~n30558;
  assign n30561 = ~n30559 & n30560;
  assign n30562 = pi608 & ~n30372;
  assign n30563 = ~n30561 & n30562;
  assign n30564 = ~n30557 & ~n30563;
  assign n30565 = pi778 & ~n30564;
  assign n30566 = ~pi778 & n30551;
  assign n30567 = ~n30565 & ~n30566;
  assign n30568 = ~pi609 & ~n30567;
  assign n30569 = ~pi1155 & ~n30514;
  assign n30570 = ~n30568 & n30569;
  assign n30571 = ~pi660 & ~n30420;
  assign n30572 = ~n30570 & n30571;
  assign n30573 = ~pi609 & n30375;
  assign n30574 = pi609 & ~n30567;
  assign n30575 = pi1155 & ~n30573;
  assign n30576 = ~n30574 & n30575;
  assign n30577 = pi660 & ~n30424;
  assign n30578 = ~n30576 & n30577;
  assign n30579 = ~n30572 & ~n30578;
  assign n30580 = pi785 & ~n30579;
  assign n30581 = ~pi785 & ~n30567;
  assign n30582 = ~n30580 & ~n30581;
  assign n30583 = ~pi618 & ~n30582;
  assign n30584 = ~pi1154 & ~n30513;
  assign n30585 = ~n30583 & n30584;
  assign n30586 = ~pi627 & ~n30432;
  assign n30587 = ~n30585 & n30586;
  assign n30588 = ~pi618 & ~n30378;
  assign n30589 = pi618 & ~n30582;
  assign n30590 = pi1154 & ~n30588;
  assign n30591 = ~n30589 & n30590;
  assign n30592 = pi627 & ~n30436;
  assign n30593 = ~n30591 & n30592;
  assign n30594 = ~n30587 & ~n30593;
  assign n30595 = pi781 & ~n30594;
  assign n30596 = ~pi781 & ~n30582;
  assign n30597 = ~n30595 & ~n30596;
  assign n30598 = ~pi789 & n30597;
  assign n30599 = ~pi619 & n30380;
  assign n30600 = pi619 & ~n30597;
  assign n30601 = pi1159 & ~n30599;
  assign n30602 = ~n30600 & n30601;
  assign n30603 = pi648 & ~n30448;
  assign n30604 = ~n30602 & n30603;
  assign n30605 = ~pi619 & ~n30597;
  assign n30606 = pi619 & n30380;
  assign n30607 = ~pi1159 & ~n30606;
  assign n30608 = ~n30605 & n30607;
  assign n30609 = ~pi648 & ~n30444;
  assign n30610 = ~n30608 & n30609;
  assign n30611 = pi789 & ~n30604;
  assign n30612 = ~n30610 & n30611;
  assign n30613 = n15833 & ~n30598;
  assign n30614 = ~n30612 & n30613;
  assign n30615 = ~n16644 & ~n30512;
  assign n30616 = ~n30614 & n30615;
  assign n30617 = ~n30500 & ~n30616;
  assign n30618 = n18841 & ~n30617;
  assign n30619 = pi644 & ~n30464;
  assign n30620 = ~n30473 & ~n30619;
  assign n30621 = ~n22949 & ~n30620;
  assign n30622 = pi790 & ~n30621;
  assign n30623 = ~n30488 & ~n30618;
  assign n30624 = ~n30622 & n30623;
  assign n30625 = ~n30476 & ~n30624;
  assign n30626 = ~po1038 & ~n30625;
  assign n30627 = ~pi832 & ~n30347;
  assign n30628 = ~n30626 & n30627;
  assign po349 = ~n30346 & ~n30628;
  assign n30630 = ~pi193 & ~n2923;
  assign n30631 = pi690 & n15726;
  assign n30632 = ~n30630 & ~n30631;
  assign n30633 = ~pi778 & ~n30632;
  assign n30634 = ~pi625 & n30631;
  assign n30635 = ~n30632 & ~n30634;
  assign n30636 = pi1153 & ~n30635;
  assign n30637 = ~pi1153 & ~n30630;
  assign n30638 = ~n30634 & n30637;
  assign n30639 = pi778 & ~n30638;
  assign n30640 = ~n30636 & n30639;
  assign n30641 = ~n30633 & ~n30640;
  assign n30642 = ~n15742 & ~n30641;
  assign n30643 = ~n15748 & n30642;
  assign n30644 = ~n15754 & n30643;
  assign n30645 = ~n15760 & n30644;
  assign n30646 = ~n15766 & n30645;
  assign n30647 = n19394 & n30646;
  assign n30648 = ~n19394 & n30630;
  assign n30649 = ~n30647 & ~n30648;
  assign n30650 = ~n15959 & n30649;
  assign n30651 = n15925 & n30630;
  assign n30652 = pi739 & n15781;
  assign n30653 = ~n30630 & ~n30652;
  assign n30654 = ~n15778 & ~n30653;
  assign n30655 = ~pi785 & ~n30654;
  assign n30656 = n16585 & n30652;
  assign n30657 = n30654 & ~n30656;
  assign n30658 = pi1155 & ~n30657;
  assign n30659 = ~pi1155 & ~n30630;
  assign n30660 = ~n30656 & n30659;
  assign n30661 = ~n30658 & ~n30660;
  assign n30662 = pi785 & ~n30661;
  assign n30663 = ~n30655 & ~n30662;
  assign n30664 = ~pi781 & ~n30663;
  assign n30665 = ~n15797 & n30663;
  assign n30666 = pi1154 & ~n30665;
  assign n30667 = ~n15800 & n30663;
  assign n30668 = ~pi1154 & ~n30667;
  assign n30669 = ~n30666 & ~n30668;
  assign n30670 = pi781 & ~n30669;
  assign n30671 = ~n30664 & ~n30670;
  assign n30672 = ~n21915 & n30671;
  assign n30673 = ~n15832 & ~n30672;
  assign n30674 = n15832 & ~n30630;
  assign n30675 = ~n30673 & ~n30674;
  assign n30676 = ~n15925 & n30675;
  assign n30677 = n19478 & ~n30651;
  assign n30678 = ~n30676 & n30677;
  assign n30679 = ~n30650 & ~n30678;
  assign n30680 = pi787 & ~n30679;
  assign n30681 = n15763 & n30675;
  assign n30682 = n15772 & n30645;
  assign n30683 = ~pi629 & ~n30682;
  assign n30684 = ~n30681 & n30683;
  assign n30685 = n15762 & n30675;
  assign n30686 = n15909 & n30645;
  assign n30687 = pi629 & ~n30686;
  assign n30688 = ~n30685 & n30687;
  assign n30689 = pi792 & ~n30684;
  assign n30690 = ~n30688 & n30689;
  assign n30691 = ~n21932 & n30671;
  assign n30692 = pi648 & ~n30691;
  assign n30693 = n21935 & ~n30643;
  assign n30694 = ~n30692 & ~n30693;
  assign n30695 = ~pi1159 & ~n30694;
  assign n30696 = ~pi619 & ~n30643;
  assign n30697 = pi648 & ~n30696;
  assign n30698 = n21942 & n30671;
  assign n30699 = pi1159 & ~n30697;
  assign n30700 = ~n30698 & n30699;
  assign n30701 = ~n30695 & ~n30700;
  assign n30702 = pi789 & ~n30701;
  assign n30703 = pi609 & ~n30641;
  assign n30704 = ~n15780 & ~n30632;
  assign n30705 = pi625 & n30704;
  assign n30706 = n30653 & ~n30704;
  assign n30707 = ~n30705 & ~n30706;
  assign n30708 = n30637 & ~n30707;
  assign n30709 = ~pi608 & ~n30636;
  assign n30710 = ~n30708 & n30709;
  assign n30711 = pi1153 & n30653;
  assign n30712 = ~n30705 & n30711;
  assign n30713 = pi608 & ~n30638;
  assign n30714 = ~n30712 & n30713;
  assign n30715 = ~n30710 & ~n30714;
  assign n30716 = pi778 & ~n30715;
  assign n30717 = ~pi778 & ~n30706;
  assign n30718 = ~n30716 & ~n30717;
  assign n30719 = ~pi609 & ~n30718;
  assign n30720 = ~pi1155 & ~n30703;
  assign n30721 = ~n30719 & n30720;
  assign n30722 = ~pi660 & ~n30658;
  assign n30723 = ~n30721 & n30722;
  assign n30724 = ~pi609 & ~n30641;
  assign n30725 = pi609 & ~n30718;
  assign n30726 = pi1155 & ~n30724;
  assign n30727 = ~n30725 & n30726;
  assign n30728 = pi660 & ~n30660;
  assign n30729 = ~n30727 & n30728;
  assign n30730 = ~n30723 & ~n30729;
  assign n30731 = pi785 & ~n30730;
  assign n30732 = ~pi785 & ~n30718;
  assign n30733 = ~n30731 & ~n30732;
  assign n30734 = ~pi781 & n30733;
  assign n30735 = pi618 & n30642;
  assign n30736 = ~pi618 & ~n30733;
  assign n30737 = ~pi1154 & ~n30735;
  assign n30738 = ~n30736 & n30737;
  assign n30739 = ~pi627 & ~n30666;
  assign n30740 = ~n30738 & n30739;
  assign n30741 = ~pi618 & n30642;
  assign n30742 = pi618 & ~n30733;
  assign n30743 = pi1154 & ~n30741;
  assign n30744 = ~n30742 & n30743;
  assign n30745 = pi627 & ~n30668;
  assign n30746 = ~n30744 & n30745;
  assign n30747 = pi781 & ~n30740;
  assign n30748 = ~n30746 & n30747;
  assign n30749 = ~n30702 & ~n30734;
  assign n30750 = ~n30748 & n30749;
  assign n30751 = n18969 & n30701;
  assign n30752 = ~n30750 & ~n30751;
  assign n30753 = n15833 & ~n30752;
  assign n30754 = n15828 & n30644;
  assign n30755 = ~pi626 & ~n30630;
  assign n30756 = pi626 & ~n30672;
  assign n30757 = n15756 & ~n30755;
  assign n30758 = ~n30756 & n30757;
  assign n30759 = pi626 & ~n30630;
  assign n30760 = ~pi626 & ~n30672;
  assign n30761 = n15757 & ~n30759;
  assign n30762 = ~n30760 & n30761;
  assign n30763 = ~n30754 & ~n30758;
  assign n30764 = ~n30762 & n30763;
  assign n30765 = pi788 & ~n30764;
  assign n30766 = ~n30753 & ~n30765;
  assign n30767 = ~n16644 & ~n30766;
  assign n30768 = n18841 & ~n30690;
  assign n30769 = ~n30767 & n30768;
  assign n30770 = ~n30680 & ~n30769;
  assign n30771 = ~pi790 & n30770;
  assign n30772 = pi787 & ~n30649;
  assign n30773 = ~pi787 & n30646;
  assign n30774 = ~n30772 & ~n30773;
  assign n30775 = ~pi644 & ~n30774;
  assign n30776 = pi644 & n30770;
  assign n30777 = pi715 & ~n30775;
  assign n30778 = ~n30776 & n30777;
  assign n30779 = ~n19771 & n30630;
  assign n30780 = ~n15960 & n30676;
  assign n30781 = ~n30779 & ~n30780;
  assign n30782 = pi644 & ~n30781;
  assign n30783 = ~pi644 & n30630;
  assign n30784 = ~pi715 & ~n30783;
  assign n30785 = ~n30782 & n30784;
  assign n30786 = pi1160 & ~n30785;
  assign n30787 = ~n30778 & n30786;
  assign n30788 = ~pi644 & ~n30781;
  assign n30789 = pi644 & n30630;
  assign n30790 = pi715 & ~n30789;
  assign n30791 = ~n30788 & n30790;
  assign n30792 = pi644 & ~n30774;
  assign n30793 = ~pi644 & n30770;
  assign n30794 = ~pi715 & ~n30792;
  assign n30795 = ~n30793 & n30794;
  assign n30796 = ~pi1160 & ~n30791;
  assign n30797 = ~n30795 & n30796;
  assign n30798 = ~n30787 & ~n30797;
  assign n30799 = pi790 & ~n30798;
  assign n30800 = pi832 & ~n30771;
  assign n30801 = ~n30799 & n30800;
  assign n30802 = ~pi193 & po1038;
  assign n30803 = ~pi193 & ~n16219;
  assign n30804 = n15747 & ~n30803;
  assign n30805 = pi690 & n9829;
  assign n30806 = n30803 & ~n30805;
  assign n30807 = ~pi193 & ~n16228;
  assign n30808 = n16227 & ~n30807;
  assign n30809 = ~pi193 & ~n17276;
  assign n30810 = ~pi38 & ~pi193;
  assign n30811 = n19350 & ~n30810;
  assign n30812 = ~n30809 & ~n30811;
  assign n30813 = pi690 & ~n30808;
  assign n30814 = ~n30812 & n30813;
  assign n30815 = ~n30806 & ~n30814;
  assign n30816 = ~pi778 & n30815;
  assign n30817 = ~pi625 & n30803;
  assign n30818 = pi625 & ~n30815;
  assign n30819 = pi1153 & ~n30817;
  assign n30820 = ~n30818 & n30819;
  assign n30821 = pi625 & n30803;
  assign n30822 = ~pi625 & ~n30815;
  assign n30823 = ~pi1153 & ~n30821;
  assign n30824 = ~n30822 & n30823;
  assign n30825 = ~n30820 & ~n30824;
  assign n30826 = pi778 & ~n30825;
  assign n30827 = ~n30816 & ~n30826;
  assign n30828 = ~n15741 & n30827;
  assign n30829 = n15741 & n30803;
  assign n30830 = ~n30828 & ~n30829;
  assign n30831 = ~n15747 & n30830;
  assign n30832 = ~n30804 & ~n30831;
  assign n30833 = ~n15753 & n30832;
  assign n30834 = n15753 & n30803;
  assign n30835 = ~n30833 & ~n30834;
  assign n30836 = ~n15759 & ~n30835;
  assign n30837 = n15759 & n30803;
  assign n30838 = ~n30836 & ~n30837;
  assign n30839 = ~pi792 & n30838;
  assign n30840 = ~pi628 & n30803;
  assign n30841 = pi628 & ~n30838;
  assign n30842 = pi1156 & ~n30840;
  assign n30843 = ~n30841 & n30842;
  assign n30844 = pi628 & n30803;
  assign n30845 = ~pi628 & ~n30838;
  assign n30846 = ~pi1156 & ~n30844;
  assign n30847 = ~n30845 & n30846;
  assign n30848 = ~n30843 & ~n30847;
  assign n30849 = pi792 & ~n30848;
  assign n30850 = ~n30839 & ~n30849;
  assign n30851 = n19394 & n30850;
  assign n30852 = ~n19394 & n30803;
  assign n30853 = ~n30851 & ~n30852;
  assign n30854 = pi787 & ~n30853;
  assign n30855 = ~pi787 & n30850;
  assign n30856 = ~n30854 & ~n30855;
  assign n30857 = ~pi644 & ~n30856;
  assign n30858 = pi715 & ~n30857;
  assign n30859 = pi193 & ~n9829;
  assign n30860 = pi739 & n16570;
  assign n30861 = ~n30807 & ~n30860;
  assign n30862 = pi38 & ~n30861;
  assign n30863 = ~pi193 & n16514;
  assign n30864 = pi193 & ~n16565;
  assign n30865 = pi739 & ~n30863;
  assign n30866 = ~n30864 & n30865;
  assign n30867 = ~pi193 & ~pi739;
  assign n30868 = ~n16214 & n30867;
  assign n30869 = ~n30866 & ~n30868;
  assign n30870 = ~pi38 & ~n30869;
  assign n30871 = ~n30862 & ~n30870;
  assign n30872 = n9829 & n30871;
  assign n30873 = ~n30859 & ~n30872;
  assign n30874 = ~n15777 & ~n30873;
  assign n30875 = n15777 & ~n30803;
  assign n30876 = ~n30874 & ~n30875;
  assign n30877 = ~pi785 & ~n30876;
  assign n30878 = ~n15786 & ~n30803;
  assign n30879 = pi609 & n30874;
  assign n30880 = ~n30878 & ~n30879;
  assign n30881 = pi1155 & ~n30880;
  assign n30882 = ~n16585 & ~n30803;
  assign n30883 = ~pi609 & n30874;
  assign n30884 = ~n30882 & ~n30883;
  assign n30885 = ~pi1155 & ~n30884;
  assign n30886 = ~n30881 & ~n30885;
  assign n30887 = pi785 & ~n30886;
  assign n30888 = ~n30877 & ~n30887;
  assign n30889 = ~pi781 & ~n30888;
  assign n30890 = ~pi618 & n30803;
  assign n30891 = pi618 & n30888;
  assign n30892 = pi1154 & ~n30890;
  assign n30893 = ~n30891 & n30892;
  assign n30894 = ~pi618 & n30888;
  assign n30895 = pi618 & n30803;
  assign n30896 = ~pi1154 & ~n30895;
  assign n30897 = ~n30894 & n30896;
  assign n30898 = ~n30893 & ~n30897;
  assign n30899 = pi781 & ~n30898;
  assign n30900 = ~n30889 & ~n30899;
  assign n30901 = ~pi789 & ~n30900;
  assign n30902 = ~pi619 & n30803;
  assign n30903 = pi619 & n30900;
  assign n30904 = pi1159 & ~n30902;
  assign n30905 = ~n30903 & n30904;
  assign n30906 = ~pi619 & n30900;
  assign n30907 = pi619 & n30803;
  assign n30908 = ~pi1159 & ~n30907;
  assign n30909 = ~n30906 & n30908;
  assign n30910 = ~n30905 & ~n30909;
  assign n30911 = pi789 & ~n30910;
  assign n30912 = ~n30901 & ~n30911;
  assign n30913 = ~n15832 & n30912;
  assign n30914 = n15832 & n30803;
  assign n30915 = ~n30913 & ~n30914;
  assign n30916 = ~n15925 & ~n30915;
  assign n30917 = n15925 & n30803;
  assign n30918 = ~n30916 & ~n30917;
  assign n30919 = ~n15960 & ~n30918;
  assign n30920 = n15960 & n30803;
  assign n30921 = ~n30919 & ~n30920;
  assign n30922 = pi644 & ~n30921;
  assign n30923 = ~pi644 & n30803;
  assign n30924 = ~pi715 & ~n30923;
  assign n30925 = ~n30922 & n30924;
  assign n30926 = pi1160 & ~n30858;
  assign n30927 = ~n30925 & n30926;
  assign n30928 = pi644 & ~n30856;
  assign n30929 = ~pi715 & ~n30928;
  assign n30930 = ~pi644 & ~n30921;
  assign n30931 = pi644 & n30803;
  assign n30932 = pi715 & ~n30931;
  assign n30933 = ~n30930 & n30932;
  assign n30934 = ~pi1160 & ~n30933;
  assign n30935 = ~n30929 & n30934;
  assign n30936 = ~n30927 & ~n30935;
  assign n30937 = pi790 & ~n30936;
  assign n30938 = n19478 & n30918;
  assign n30939 = ~n15959 & n30853;
  assign n30940 = ~n30938 & ~n30939;
  assign n30941 = pi787 & ~n30940;
  assign n30942 = ~n16633 & n30915;
  assign n30943 = ~pi629 & n30843;
  assign n30944 = pi629 & n30847;
  assign n30945 = ~n30943 & ~n30944;
  assign n30946 = ~n30942 & n30945;
  assign n30947 = pi792 & ~n30946;
  assign n30948 = n15828 & ~n30835;
  assign n30949 = ~pi626 & ~n30803;
  assign n30950 = pi626 & ~n30912;
  assign n30951 = n15756 & ~n30949;
  assign n30952 = ~n30950 & n30951;
  assign n30953 = pi626 & ~n30803;
  assign n30954 = ~pi626 & ~n30912;
  assign n30955 = n15757 & ~n30953;
  assign n30956 = ~n30954 & n30955;
  assign n30957 = ~n30948 & ~n30952;
  assign n30958 = ~n30956 & n30957;
  assign n30959 = pi788 & ~n30958;
  assign n30960 = pi618 & ~n30830;
  assign n30961 = pi609 & n30827;
  assign n30962 = ~pi193 & n16653;
  assign n30963 = pi193 & n16657;
  assign n30964 = ~pi739 & ~n30962;
  assign n30965 = ~n30963 & n30964;
  assign n30966 = ~pi193 & ~n16647;
  assign n30967 = pi193 & ~n17397;
  assign n30968 = pi739 & ~n30966;
  assign n30969 = ~n30967 & n30968;
  assign n30970 = ~pi39 & ~n30969;
  assign n30971 = ~n30965 & n30970;
  assign n30972 = ~pi193 & n16877;
  assign n30973 = pi193 & n16913;
  assign n30974 = pi739 & ~n30972;
  assign n30975 = ~n30973 & n30974;
  assign n30976 = pi193 & n16825;
  assign n30977 = ~pi193 & ~n16747;
  assign n30978 = ~pi739 & ~n30976;
  assign n30979 = ~n30977 & n30978;
  assign n30980 = pi39 & ~n30975;
  assign n30981 = ~n30979 & n30980;
  assign n30982 = ~pi38 & ~n30971;
  assign n30983 = ~n30981 & n30982;
  assign n30984 = ~n16921 & ~n30652;
  assign n30985 = pi193 & ~n30984;
  assign n30986 = n6081 & n30985;
  assign n30987 = ~pi739 & n22848;
  assign n30988 = ~n16808 & ~n30987;
  assign n30989 = ~pi39 & ~n30988;
  assign n30990 = ~pi193 & ~n30989;
  assign n30991 = pi38 & ~n30986;
  assign n30992 = ~n30990 & n30991;
  assign n30993 = pi690 & ~n30992;
  assign n30994 = ~n30983 & n30993;
  assign n30995 = ~pi690 & ~n30871;
  assign n30996 = n9829 & ~n30994;
  assign n30997 = ~n30995 & n30996;
  assign n30998 = ~n30859 & ~n30997;
  assign n30999 = ~pi625 & n30998;
  assign n31000 = pi625 & n30873;
  assign n31001 = ~pi1153 & ~n31000;
  assign n31002 = ~n30999 & n31001;
  assign n31003 = ~pi608 & ~n30820;
  assign n31004 = ~n31002 & n31003;
  assign n31005 = ~pi625 & n30873;
  assign n31006 = pi625 & n30998;
  assign n31007 = pi1153 & ~n31005;
  assign n31008 = ~n31006 & n31007;
  assign n31009 = pi608 & ~n30824;
  assign n31010 = ~n31008 & n31009;
  assign n31011 = ~n31004 & ~n31010;
  assign n31012 = pi778 & ~n31011;
  assign n31013 = ~pi778 & n30998;
  assign n31014 = ~n31012 & ~n31013;
  assign n31015 = ~pi609 & ~n31014;
  assign n31016 = ~pi1155 & ~n30961;
  assign n31017 = ~n31015 & n31016;
  assign n31018 = ~pi660 & ~n30881;
  assign n31019 = ~n31017 & n31018;
  assign n31020 = ~pi609 & n30827;
  assign n31021 = pi609 & ~n31014;
  assign n31022 = pi1155 & ~n31020;
  assign n31023 = ~n31021 & n31022;
  assign n31024 = pi660 & ~n30885;
  assign n31025 = ~n31023 & n31024;
  assign n31026 = ~n31019 & ~n31025;
  assign n31027 = pi785 & ~n31026;
  assign n31028 = ~pi785 & ~n31014;
  assign n31029 = ~n31027 & ~n31028;
  assign n31030 = ~pi618 & ~n31029;
  assign n31031 = ~pi1154 & ~n30960;
  assign n31032 = ~n31030 & n31031;
  assign n31033 = ~pi627 & ~n30893;
  assign n31034 = ~n31032 & n31033;
  assign n31035 = ~pi618 & ~n30830;
  assign n31036 = pi618 & ~n31029;
  assign n31037 = pi1154 & ~n31035;
  assign n31038 = ~n31036 & n31037;
  assign n31039 = pi627 & ~n30897;
  assign n31040 = ~n31038 & n31039;
  assign n31041 = ~n31034 & ~n31040;
  assign n31042 = pi781 & ~n31041;
  assign n31043 = ~pi781 & ~n31029;
  assign n31044 = ~n31042 & ~n31043;
  assign n31045 = ~pi789 & n31044;
  assign n31046 = ~pi619 & n30832;
  assign n31047 = pi619 & ~n31044;
  assign n31048 = pi1159 & ~n31046;
  assign n31049 = ~n31047 & n31048;
  assign n31050 = pi648 & ~n30909;
  assign n31051 = ~n31049 & n31050;
  assign n31052 = ~pi619 & ~n31044;
  assign n31053 = pi619 & n30832;
  assign n31054 = ~pi1159 & ~n31053;
  assign n31055 = ~n31052 & n31054;
  assign n31056 = ~pi648 & ~n30905;
  assign n31057 = ~n31055 & n31056;
  assign n31058 = pi789 & ~n31051;
  assign n31059 = ~n31057 & n31058;
  assign n31060 = n15833 & ~n31045;
  assign n31061 = ~n31059 & n31060;
  assign n31062 = ~n16644 & ~n30959;
  assign n31063 = ~n31061 & n31062;
  assign n31064 = ~n30947 & ~n31063;
  assign n31065 = n18841 & ~n31064;
  assign n31066 = pi644 & ~n30925;
  assign n31067 = ~n30934 & ~n31066;
  assign n31068 = ~n22949 & ~n31067;
  assign n31069 = pi790 & ~n31068;
  assign n31070 = ~n30941 & ~n31065;
  assign n31071 = ~n31069 & n31070;
  assign n31072 = ~n30937 & ~n31071;
  assign n31073 = ~po1038 & ~n31072;
  assign n31074 = ~pi832 & ~n30802;
  assign n31075 = ~n31073 & n31074;
  assign po350 = ~n30801 & ~n31075;
  assign n31077 = ~pi194 & ~n2923;
  assign n31078 = pi730 & n15726;
  assign n31079 = ~n31077 & ~n31078;
  assign n31080 = ~pi778 & n31079;
  assign n31081 = ~pi625 & n31078;
  assign n31082 = ~n31079 & ~n31081;
  assign n31083 = pi1153 & ~n31082;
  assign n31084 = ~pi1153 & ~n31077;
  assign n31085 = ~n31081 & n31084;
  assign n31086 = ~n31083 & ~n31085;
  assign n31087 = pi778 & ~n31086;
  assign n31088 = ~n31080 & ~n31087;
  assign n31089 = ~n15742 & n31088;
  assign n31090 = ~n15748 & n31089;
  assign n31091 = ~n15754 & n31090;
  assign n31092 = ~n15760 & n31091;
  assign n31093 = ~n15766 & n31092;
  assign n31094 = n19394 & n31093;
  assign n31095 = ~n19394 & n31077;
  assign n31096 = ~n31094 & ~n31095;
  assign n31097 = ~n15959 & n31096;
  assign n31098 = n15925 & n31077;
  assign n31099 = pi748 & n15781;
  assign n31100 = ~n31077 & ~n31099;
  assign n31101 = ~n15778 & ~n31100;
  assign n31102 = ~pi785 & ~n31101;
  assign n31103 = ~n15787 & ~n31100;
  assign n31104 = pi1155 & ~n31103;
  assign n31105 = ~n15790 & n31101;
  assign n31106 = ~pi1155 & ~n31105;
  assign n31107 = ~n31104 & ~n31106;
  assign n31108 = pi785 & ~n31107;
  assign n31109 = ~n31102 & ~n31108;
  assign n31110 = ~pi781 & ~n31109;
  assign n31111 = ~n15797 & n31109;
  assign n31112 = pi1154 & ~n31111;
  assign n31113 = ~n15800 & n31109;
  assign n31114 = ~pi1154 & ~n31113;
  assign n31115 = ~n31112 & ~n31114;
  assign n31116 = pi781 & ~n31115;
  assign n31117 = ~n31110 & ~n31116;
  assign n31118 = ~pi789 & ~n31117;
  assign n31119 = ~pi619 & n31077;
  assign n31120 = pi619 & n31117;
  assign n31121 = pi1159 & ~n31119;
  assign n31122 = ~n31120 & n31121;
  assign n31123 = ~pi619 & n31117;
  assign n31124 = pi619 & n31077;
  assign n31125 = ~pi1159 & ~n31124;
  assign n31126 = ~n31123 & n31125;
  assign n31127 = ~n31122 & ~n31126;
  assign n31128 = pi789 & ~n31127;
  assign n31129 = ~n31118 & ~n31128;
  assign n31130 = ~n15832 & ~n31129;
  assign n31131 = n15832 & ~n31077;
  assign n31132 = ~n31130 & ~n31131;
  assign n31133 = ~n15925 & n31132;
  assign n31134 = n19478 & ~n31098;
  assign n31135 = ~n31133 & n31134;
  assign n31136 = ~n31097 & ~n31135;
  assign n31137 = pi787 & ~n31136;
  assign n31138 = n15828 & n31091;
  assign n31139 = ~pi626 & ~n31077;
  assign n31140 = pi626 & ~n31129;
  assign n31141 = n15756 & ~n31139;
  assign n31142 = ~n31140 & n31141;
  assign n31143 = pi626 & ~n31077;
  assign n31144 = ~pi626 & ~n31129;
  assign n31145 = n15757 & ~n31143;
  assign n31146 = ~n31144 & n31145;
  assign n31147 = ~n31138 & ~n31142;
  assign n31148 = ~n31146 & n31147;
  assign n31149 = pi788 & ~n31148;
  assign n31150 = pi618 & n31089;
  assign n31151 = pi609 & n31088;
  assign n31152 = ~n15780 & ~n31079;
  assign n31153 = pi625 & n31152;
  assign n31154 = n31100 & ~n31152;
  assign n31155 = ~n31153 & ~n31154;
  assign n31156 = n31084 & ~n31155;
  assign n31157 = ~pi608 & ~n31083;
  assign n31158 = ~n31156 & n31157;
  assign n31159 = pi1153 & n31100;
  assign n31160 = ~n31153 & n31159;
  assign n31161 = pi608 & ~n31085;
  assign n31162 = ~n31160 & n31161;
  assign n31163 = ~n31158 & ~n31162;
  assign n31164 = pi778 & ~n31163;
  assign n31165 = ~pi778 & ~n31154;
  assign n31166 = ~n31164 & ~n31165;
  assign n31167 = ~pi609 & ~n31166;
  assign n31168 = ~pi1155 & ~n31151;
  assign n31169 = ~n31167 & n31168;
  assign n31170 = ~pi660 & ~n31104;
  assign n31171 = ~n31169 & n31170;
  assign n31172 = ~pi609 & n31088;
  assign n31173 = pi609 & ~n31166;
  assign n31174 = pi1155 & ~n31172;
  assign n31175 = ~n31173 & n31174;
  assign n31176 = pi660 & ~n31106;
  assign n31177 = ~n31175 & n31176;
  assign n31178 = ~n31171 & ~n31177;
  assign n31179 = pi785 & ~n31178;
  assign n31180 = ~pi785 & ~n31166;
  assign n31181 = ~n31179 & ~n31180;
  assign n31182 = ~pi618 & ~n31181;
  assign n31183 = ~pi1154 & ~n31150;
  assign n31184 = ~n31182 & n31183;
  assign n31185 = ~pi627 & ~n31112;
  assign n31186 = ~n31184 & n31185;
  assign n31187 = ~pi618 & n31089;
  assign n31188 = pi618 & ~n31181;
  assign n31189 = pi1154 & ~n31187;
  assign n31190 = ~n31188 & n31189;
  assign n31191 = pi627 & ~n31114;
  assign n31192 = ~n31190 & n31191;
  assign n31193 = ~n31186 & ~n31192;
  assign n31194 = pi781 & ~n31193;
  assign n31195 = ~pi781 & ~n31181;
  assign n31196 = ~n31194 & ~n31195;
  assign n31197 = ~pi789 & n31196;
  assign n31198 = ~pi619 & n31090;
  assign n31199 = pi619 & ~n31196;
  assign n31200 = pi1159 & ~n31198;
  assign n31201 = ~n31199 & n31200;
  assign n31202 = pi648 & ~n31126;
  assign n31203 = ~n31201 & n31202;
  assign n31204 = pi619 & n31090;
  assign n31205 = ~pi619 & ~n31196;
  assign n31206 = ~pi1159 & ~n31204;
  assign n31207 = ~n31205 & n31206;
  assign n31208 = ~pi648 & ~n31122;
  assign n31209 = ~n31207 & n31208;
  assign n31210 = pi789 & ~n31203;
  assign n31211 = ~n31209 & n31210;
  assign n31212 = n15833 & ~n31197;
  assign n31213 = ~n31211 & n31212;
  assign n31214 = ~n31149 & ~n31213;
  assign n31215 = ~n16644 & ~n31214;
  assign n31216 = n15763 & n31132;
  assign n31217 = n15772 & n31092;
  assign n31218 = ~pi629 & ~n31217;
  assign n31219 = ~n31216 & n31218;
  assign n31220 = n15762 & n31132;
  assign n31221 = n15909 & n31092;
  assign n31222 = pi629 & ~n31221;
  assign n31223 = ~n31220 & n31222;
  assign n31224 = pi792 & ~n31219;
  assign n31225 = ~n31223 & n31224;
  assign n31226 = n18841 & ~n31225;
  assign n31227 = ~n31215 & n31226;
  assign n31228 = ~n31137 & ~n31227;
  assign n31229 = ~pi790 & n31228;
  assign n31230 = pi787 & ~n31096;
  assign n31231 = ~pi787 & n31093;
  assign n31232 = ~n31230 & ~n31231;
  assign n31233 = ~pi644 & ~n31232;
  assign n31234 = pi644 & n31228;
  assign n31235 = pi715 & ~n31233;
  assign n31236 = ~n31234 & n31235;
  assign n31237 = ~n19771 & n31077;
  assign n31238 = ~n15960 & n31133;
  assign n31239 = ~n31237 & ~n31238;
  assign n31240 = pi644 & ~n31239;
  assign n31241 = ~pi644 & n31077;
  assign n31242 = ~pi715 & ~n31241;
  assign n31243 = ~n31240 & n31242;
  assign n31244 = pi1160 & ~n31243;
  assign n31245 = ~n31236 & n31244;
  assign n31246 = ~pi644 & ~n31239;
  assign n31247 = pi644 & n31077;
  assign n31248 = pi715 & ~n31247;
  assign n31249 = ~n31246 & n31248;
  assign n31250 = pi644 & ~n31232;
  assign n31251 = ~pi644 & n31228;
  assign n31252 = ~pi715 & ~n31250;
  assign n31253 = ~n31251 & n31252;
  assign n31254 = ~pi1160 & ~n31249;
  assign n31255 = ~n31253 & n31254;
  assign n31256 = ~n31245 & ~n31255;
  assign n31257 = pi790 & ~n31256;
  assign n31258 = pi832 & ~n31229;
  assign n31259 = ~n31257 & n31258;
  assign n31260 = ~pi194 & po1038;
  assign n31261 = ~pi194 & ~n16219;
  assign n31262 = n15759 & ~n31261;
  assign n31263 = n15747 & ~n31261;
  assign n31264 = pi194 & ~n23147;
  assign n31265 = ~pi194 & n23150;
  assign n31266 = pi730 & ~n31265;
  assign n31267 = ~pi194 & ~n16218;
  assign n31268 = ~pi730 & n31267;
  assign n31269 = n9829 & ~n31266;
  assign n31270 = ~n31268 & n31269;
  assign n31271 = ~n31264 & ~n31270;
  assign n31272 = ~pi778 & ~n31271;
  assign n31273 = ~pi625 & n31261;
  assign n31274 = pi625 & n31271;
  assign n31275 = pi1153 & ~n31273;
  assign n31276 = ~n31274 & n31275;
  assign n31277 = ~pi625 & n31271;
  assign n31278 = pi625 & n31261;
  assign n31279 = ~pi1153 & ~n31278;
  assign n31280 = ~n31277 & n31279;
  assign n31281 = ~n31276 & ~n31280;
  assign n31282 = pi778 & ~n31281;
  assign n31283 = ~n31272 & ~n31282;
  assign n31284 = ~n15741 & n31283;
  assign n31285 = n15741 & n31261;
  assign n31286 = ~n31284 & ~n31285;
  assign n31287 = ~n15747 & n31286;
  assign n31288 = ~n31263 & ~n31287;
  assign n31289 = ~n15753 & n31288;
  assign n31290 = n15753 & n31261;
  assign n31291 = ~n31289 & ~n31290;
  assign n31292 = ~n15759 & n31291;
  assign n31293 = ~n31262 & ~n31292;
  assign n31294 = ~pi792 & ~n31293;
  assign n31295 = ~pi628 & ~n31261;
  assign n31296 = pi628 & ~n31293;
  assign n31297 = ~n31295 & ~n31296;
  assign n31298 = pi1156 & ~n31297;
  assign n31299 = ~pi628 & n31293;
  assign n31300 = pi628 & n31261;
  assign n31301 = ~pi1156 & ~n31300;
  assign n31302 = ~n31299 & n31301;
  assign n31303 = ~n31298 & ~n31302;
  assign n31304 = pi792 & ~n31303;
  assign n31305 = ~n31294 & ~n31304;
  assign n31306 = ~pi787 & ~n31305;
  assign n31307 = ~pi647 & n31261;
  assign n31308 = pi647 & n31305;
  assign n31309 = pi1157 & ~n31307;
  assign n31310 = ~n31308 & n31309;
  assign n31311 = ~pi647 & n31305;
  assign n31312 = pi647 & n31261;
  assign n31313 = ~pi1157 & ~n31312;
  assign n31314 = ~n31311 & n31313;
  assign n31315 = ~n31310 & ~n31314;
  assign n31316 = pi787 & ~n31315;
  assign n31317 = ~n31306 & ~n31316;
  assign n31318 = ~pi644 & n31317;
  assign n31319 = ~pi629 & n31298;
  assign n31320 = pi194 & ~n9829;
  assign n31321 = ~pi194 & n18604;
  assign n31322 = pi194 & n23191;
  assign n31323 = ~n31321 & ~n31322;
  assign n31324 = pi748 & ~n31323;
  assign n31325 = ~pi748 & ~n31267;
  assign n31326 = ~n31324 & ~n31325;
  assign n31327 = n9829 & ~n31326;
  assign n31328 = ~n31320 & ~n31327;
  assign n31329 = ~n15777 & ~n31328;
  assign n31330 = n15777 & ~n31261;
  assign n31331 = ~n31329 & ~n31330;
  assign n31332 = ~pi785 & ~n31331;
  assign n31333 = ~n15786 & ~n31261;
  assign n31334 = pi609 & n31329;
  assign n31335 = ~n31333 & ~n31334;
  assign n31336 = pi1155 & ~n31335;
  assign n31337 = ~n16585 & ~n31261;
  assign n31338 = ~pi609 & n31329;
  assign n31339 = ~n31337 & ~n31338;
  assign n31340 = ~pi1155 & ~n31339;
  assign n31341 = ~n31336 & ~n31340;
  assign n31342 = pi785 & ~n31341;
  assign n31343 = ~n31332 & ~n31342;
  assign n31344 = ~pi781 & ~n31343;
  assign n31345 = ~pi618 & n31261;
  assign n31346 = pi618 & n31343;
  assign n31347 = pi1154 & ~n31345;
  assign n31348 = ~n31346 & n31347;
  assign n31349 = ~pi618 & n31343;
  assign n31350 = pi618 & n31261;
  assign n31351 = ~pi1154 & ~n31350;
  assign n31352 = ~n31349 & n31351;
  assign n31353 = ~n31348 & ~n31352;
  assign n31354 = pi781 & ~n31353;
  assign n31355 = ~n31344 & ~n31354;
  assign n31356 = ~pi789 & ~n31355;
  assign n31357 = ~pi619 & n31261;
  assign n31358 = pi619 & n31355;
  assign n31359 = pi1159 & ~n31357;
  assign n31360 = ~n31358 & n31359;
  assign n31361 = ~pi619 & n31355;
  assign n31362 = pi619 & n31261;
  assign n31363 = ~pi1159 & ~n31362;
  assign n31364 = ~n31361 & n31363;
  assign n31365 = ~n31360 & ~n31364;
  assign n31366 = pi789 & ~n31365;
  assign n31367 = ~n31356 & ~n31366;
  assign n31368 = ~n15832 & n31367;
  assign n31369 = n15832 & n31261;
  assign n31370 = ~n31368 & ~n31369;
  assign n31371 = ~n16633 & n31370;
  assign n31372 = pi629 & n31302;
  assign n31373 = ~n31319 & ~n31372;
  assign n31374 = ~n31371 & n31373;
  assign n31375 = pi792 & ~n31374;
  assign n31376 = pi619 & n31288;
  assign n31377 = ~pi1159 & ~n31376;
  assign n31378 = ~pi648 & ~n31360;
  assign n31379 = ~n31377 & n31378;
  assign n31380 = pi618 & ~n31286;
  assign n31381 = pi609 & n31283;
  assign n31382 = ~pi730 & n31326;
  assign n31383 = ~pi194 & n18651;
  assign n31384 = pi194 & ~n18659;
  assign n31385 = pi748 & ~n31383;
  assign n31386 = ~n31384 & n31385;
  assign n31387 = ~pi194 & ~n18675;
  assign n31388 = pi194 & n23308;
  assign n31389 = ~pi748 & ~n31388;
  assign n31390 = ~n31387 & n31389;
  assign n31391 = ~n31386 & ~n31390;
  assign n31392 = pi730 & ~n31391;
  assign n31393 = n9829 & ~n31382;
  assign n31394 = ~n31392 & n31393;
  assign n31395 = ~n31320 & ~n31394;
  assign n31396 = ~pi625 & n31395;
  assign n31397 = pi625 & n31328;
  assign n31398 = ~pi1153 & ~n31397;
  assign n31399 = ~n31396 & n31398;
  assign n31400 = ~pi608 & ~n31276;
  assign n31401 = ~n31399 & n31400;
  assign n31402 = ~pi625 & n31328;
  assign n31403 = pi625 & n31395;
  assign n31404 = pi1153 & ~n31402;
  assign n31405 = ~n31403 & n31404;
  assign n31406 = pi608 & ~n31280;
  assign n31407 = ~n31405 & n31406;
  assign n31408 = ~n31401 & ~n31407;
  assign n31409 = pi778 & ~n31408;
  assign n31410 = ~pi778 & n31395;
  assign n31411 = ~n31409 & ~n31410;
  assign n31412 = ~pi609 & ~n31411;
  assign n31413 = ~pi1155 & ~n31381;
  assign n31414 = ~n31412 & n31413;
  assign n31415 = ~pi660 & ~n31336;
  assign n31416 = ~n31414 & n31415;
  assign n31417 = ~pi609 & n31283;
  assign n31418 = pi609 & ~n31411;
  assign n31419 = pi1155 & ~n31417;
  assign n31420 = ~n31418 & n31419;
  assign n31421 = pi660 & ~n31340;
  assign n31422 = ~n31420 & n31421;
  assign n31423 = ~n31416 & ~n31422;
  assign n31424 = pi785 & ~n31423;
  assign n31425 = ~pi785 & ~n31411;
  assign n31426 = ~n31424 & ~n31425;
  assign n31427 = ~pi618 & ~n31426;
  assign n31428 = ~pi1154 & ~n31380;
  assign n31429 = ~n31427 & n31428;
  assign n31430 = ~pi627 & ~n31348;
  assign n31431 = ~n31429 & n31430;
  assign n31432 = ~pi618 & ~n31286;
  assign n31433 = pi618 & ~n31426;
  assign n31434 = pi1154 & ~n31432;
  assign n31435 = ~n31433 & n31434;
  assign n31436 = pi627 & ~n31352;
  assign n31437 = ~n31435 & n31436;
  assign n31438 = ~n31431 & ~n31437;
  assign n31439 = pi781 & ~n31438;
  assign n31440 = ~pi781 & ~n31426;
  assign n31441 = ~n31439 & ~n31440;
  assign n31442 = pi619 & ~n31441;
  assign n31443 = ~pi619 & n31288;
  assign n31444 = pi1159 & ~n31443;
  assign n31445 = ~n31442 & n31444;
  assign n31446 = pi648 & ~n31364;
  assign n31447 = ~n31445 & n31446;
  assign n31448 = ~n31379 & ~n31447;
  assign n31449 = pi789 & ~n31448;
  assign n31450 = ~pi619 & n31378;
  assign n31451 = pi789 & ~n31450;
  assign n31452 = ~n31441 & ~n31451;
  assign n31453 = ~n31449 & ~n31452;
  assign n31454 = n15833 & ~n31453;
  assign n31455 = pi641 & ~n31261;
  assign n31456 = ~pi641 & n31291;
  assign n31457 = n15819 & ~n31455;
  assign n31458 = ~n31456 & n31457;
  assign n31459 = n22348 & n31367;
  assign n31460 = ~pi641 & ~n31261;
  assign n31461 = pi641 & n31291;
  assign n31462 = n15818 & ~n31460;
  assign n31463 = ~n31461 & n31462;
  assign n31464 = ~n31458 & ~n31463;
  assign n31465 = ~n31459 & n31464;
  assign n31466 = pi788 & ~n31465;
  assign n31467 = ~n16644 & ~n31466;
  assign n31468 = ~n31454 & n31467;
  assign n31469 = ~n31375 & ~n31468;
  assign n31470 = ~pi647 & n31469;
  assign n31471 = ~n15925 & ~n31370;
  assign n31472 = n15925 & n31261;
  assign n31473 = ~n31471 & ~n31472;
  assign n31474 = pi647 & ~n31473;
  assign n31475 = ~pi1157 & ~n31474;
  assign n31476 = ~n31470 & n31475;
  assign n31477 = ~pi630 & ~n31310;
  assign n31478 = ~n31476 & n31477;
  assign n31479 = ~pi647 & ~n31473;
  assign n31480 = pi647 & n31469;
  assign n31481 = pi1157 & ~n31479;
  assign n31482 = ~n31480 & n31481;
  assign n31483 = pi630 & ~n31314;
  assign n31484 = ~n31482 & n31483;
  assign n31485 = ~n31478 & ~n31484;
  assign n31486 = pi787 & ~n31485;
  assign n31487 = ~pi787 & n31469;
  assign n31488 = ~n31486 & ~n31487;
  assign n31489 = pi644 & ~n31488;
  assign n31490 = pi715 & ~n31318;
  assign n31491 = ~n31489 & n31490;
  assign n31492 = ~n15960 & ~n31473;
  assign n31493 = n15960 & n31261;
  assign n31494 = ~n31492 & ~n31493;
  assign n31495 = pi644 & ~n31494;
  assign n31496 = ~pi644 & n31261;
  assign n31497 = ~pi715 & ~n31496;
  assign n31498 = ~n31495 & n31497;
  assign n31499 = pi1160 & ~n31498;
  assign n31500 = ~n31491 & n31499;
  assign n31501 = pi644 & n31317;
  assign n31502 = ~pi715 & ~n31501;
  assign n31503 = ~pi644 & ~n31494;
  assign n31504 = pi644 & n31261;
  assign n31505 = pi715 & ~n31504;
  assign n31506 = ~n31503 & n31505;
  assign n31507 = ~pi1160 & ~n31506;
  assign n31508 = ~n31502 & n31507;
  assign n31509 = ~n31500 & ~n31508;
  assign n31510 = pi790 & ~n31509;
  assign n31511 = ~pi644 & n31507;
  assign n31512 = pi790 & ~n31511;
  assign n31513 = ~n31488 & ~n31512;
  assign n31514 = ~n31510 & ~n31513;
  assign n31515 = ~po1038 & ~n31514;
  assign n31516 = ~pi832 & ~n31260;
  assign n31517 = ~n31515 & n31516;
  assign po351 = ~n31259 & ~n31517;
  assign n31519 = ~pi138 & n15656;
  assign n31520 = ~pi196 & n31519;
  assign n31521 = pi195 & ~n31520;
  assign n31522 = ~n11063 & n15296;
  assign n31523 = ~n6205 & n15264;
  assign n31524 = n15263 & ~n15587;
  assign n31525 = ~n11066 & ~n31523;
  assign n31526 = ~n31522 & ~n31524;
  assign n31527 = n31525 & n31526;
  assign n31528 = pi232 & ~n31527;
  assign n31529 = ~n15667 & ~n31528;
  assign n31530 = pi39 & ~n31529;
  assign n31531 = n11070 & ~n15266;
  assign n31532 = ~pi39 & ~n31531;
  assign n31533 = n9833 & ~n31521;
  assign n31534 = ~n31532 & n31533;
  assign n31535 = ~n31530 & n31534;
  assign n31536 = ~pi192 & n15625;
  assign n31537 = n15263 & ~n15631;
  assign n31538 = ~n9219 & ~n15258;
  assign n31539 = pi171 & n13005;
  assign n31540 = ~n31538 & ~n31539;
  assign n31541 = pi299 & ~n31540;
  assign n31542 = pi232 & ~n31536;
  assign n31543 = ~n31537 & n31542;
  assign n31544 = ~n31541 & n31543;
  assign n31545 = n15628 & ~n31544;
  assign n31546 = ~pi192 & n15605;
  assign n31547 = ~pi171 & n9008;
  assign n31548 = ~n15612 & ~n31547;
  assign n31549 = n8739 & ~n31548;
  assign n31550 = n8979 & ~n31549;
  assign n31551 = pi192 & n15696;
  assign n31552 = ~n31550 & ~n31551;
  assign n31553 = pi232 & ~n31552;
  assign n31554 = ~n15611 & ~n31546;
  assign n31555 = ~n31553 & n31554;
  assign n31556 = pi39 & ~n31555;
  assign n31557 = n2613 & ~n31556;
  assign n31558 = ~n31545 & n31557;
  assign n31559 = ~pi87 & ~n31558;
  assign n31560 = n15601 & ~n31559;
  assign n31561 = ~pi92 & ~n31560;
  assign n31562 = n15600 & ~n31561;
  assign n31563 = ~pi55 & ~n31562;
  assign n31564 = ~n15650 & ~n31563;
  assign n31565 = n2530 & ~n31564;
  assign n31566 = n9532 & n31521;
  assign n31567 = ~n31565 & n31566;
  assign po352 = n31535 | n31567;
  assign n31569 = ~pi170 & n8740;
  assign n31570 = ~n15586 & ~n31569;
  assign n31571 = n12407 & ~n31570;
  assign n31572 = n12409 & n15586;
  assign n31573 = pi232 & ~n31572;
  assign n31574 = ~n31571 & n31573;
  assign n31575 = ~n15667 & ~n31574;
  assign n31576 = pi39 & ~n31575;
  assign n31577 = n11070 & n15381;
  assign n31578 = ~pi39 & ~n31577;
  assign n31579 = ~pi38 & ~n31578;
  assign n31580 = ~n31576 & n31579;
  assign n31581 = pi194 & ~n31580;
  assign n31582 = pi299 & ~n31575;
  assign n31583 = ~n11064 & ~n31582;
  assign n31584 = pi39 & ~n31583;
  assign n31585 = n11070 & ~n15370;
  assign n31586 = ~pi39 & ~n31585;
  assign n31587 = ~pi38 & ~n31586;
  assign n31588 = ~n31584 & n31587;
  assign n31589 = ~pi194 & ~n31588;
  assign n31590 = n9830 & ~n31581;
  assign n31591 = ~n31589 & n31590;
  assign n31592 = ~pi196 & ~n31591;
  assign n31593 = ~pi170 & n9008;
  assign n31594 = ~n15612 & ~n31593;
  assign n31595 = n8739 & ~n31594;
  assign n31596 = n8979 & ~n31595;
  assign n31597 = ~n15605 & ~n31596;
  assign n31598 = pi232 & ~n31597;
  assign n31599 = ~n15611 & ~n31598;
  assign n31600 = pi232 & n15696;
  assign n31601 = n31599 & ~n31600;
  assign n31602 = pi39 & ~n31601;
  assign n31603 = ~pi38 & pi194;
  assign n31604 = ~n31602 & n31603;
  assign n31605 = pi39 & ~n31599;
  assign n31606 = ~pi38 & ~pi194;
  assign n31607 = ~n31605 & n31606;
  assign n31608 = ~n31604 & ~n31607;
  assign n31609 = ~n9219 & ~n15369;
  assign n31610 = pi170 & n13005;
  assign n31611 = n10277 & ~n31609;
  assign n31612 = ~n31610 & n31611;
  assign n31613 = n15628 & ~n31612;
  assign n31614 = ~n31608 & ~n31613;
  assign n31615 = n9634 & n31607;
  assign n31616 = n15631 & n31604;
  assign n31617 = ~n31615 & ~n31616;
  assign n31618 = n10439 & ~n31617;
  assign n31619 = ~n31614 & ~n31618;
  assign n31620 = ~pi100 & ~n31619;
  assign n31621 = ~pi87 & ~n31620;
  assign n31622 = n15601 & ~n31621;
  assign n31623 = ~pi92 & ~n31622;
  assign n31624 = n15600 & ~n31623;
  assign n31625 = ~pi55 & ~n31624;
  assign n31626 = ~n15650 & ~n31625;
  assign n31627 = n2530 & ~n31626;
  assign n31628 = n9532 & ~n31627;
  assign n31629 = pi196 & ~n31628;
  assign n31630 = ~n31519 & ~n31592;
  assign n31631 = ~n31629 & n31630;
  assign n31632 = pi195 & ~pi196;
  assign n31633 = ~n31591 & ~n31632;
  assign n31634 = ~n31628 & n31632;
  assign n31635 = n31519 & ~n31633;
  assign n31636 = ~n31634 & n31635;
  assign po353 = n31631 | n31636;
  assign n31638 = ~pi197 & ~n2923;
  assign n31639 = ~pi767 & pi947;
  assign n31640 = ~pi698 & n19798;
  assign n31641 = ~n31639 & ~n31640;
  assign n31642 = n2923 & ~n31641;
  assign n31643 = pi832 & ~n31638;
  assign n31644 = ~n31642 & n31643;
  assign n31645 = ~pi197 & ~n9830;
  assign n31646 = n16228 & ~n31639;
  assign n31647 = pi197 & ~n16216;
  assign n31648 = pi38 & ~n31646;
  assign n31649 = ~n31647 & n31648;
  assign n31650 = ~pi197 & ~n16057;
  assign n31651 = n16057 & n31639;
  assign n31652 = ~pi39 & ~n31650;
  assign n31653 = ~n31651 & n31652;
  assign n31654 = ~pi197 & pi767;
  assign n31655 = ~n16212 & n31654;
  assign n31656 = ~pi197 & ~n16190;
  assign n31657 = n19905 & ~n31656;
  assign n31658 = pi197 & ~n20042;
  assign n31659 = ~pi197 & ~n19886;
  assign n31660 = pi299 & ~n31658;
  assign n31661 = ~n31659 & n31660;
  assign n31662 = ~pi767 & ~n31657;
  assign n31663 = ~n31661 & n31662;
  assign n31664 = pi39 & ~n31655;
  assign n31665 = ~n31663 & n31664;
  assign n31666 = ~pi38 & ~n31653;
  assign n31667 = ~n31665 & n31666;
  assign n31668 = ~n31649 & ~n31667;
  assign n31669 = pi698 & ~n31668;
  assign n31670 = ~n19958 & n31653;
  assign n31671 = n19955 & ~n31656;
  assign n31672 = pi197 & n19952;
  assign n31673 = ~pi197 & n19935;
  assign n31674 = pi299 & ~n31672;
  assign n31675 = ~n31673 & n31674;
  assign n31676 = pi767 & ~n31671;
  assign n31677 = ~n31675 & n31676;
  assign n31678 = ~pi197 & n19976;
  assign n31679 = pi197 & n19989;
  assign n31680 = ~pi767 & ~n31679;
  assign n31681 = ~n31678 & n31680;
  assign n31682 = pi39 & ~n31677;
  assign n31683 = ~n31681 & n31682;
  assign n31684 = ~n31670 & ~n31683;
  assign n31685 = ~pi38 & ~n31684;
  assign n31686 = ~pi197 & ~n16228;
  assign n31687 = ~n19798 & ~n31639;
  assign n31688 = n16228 & ~n31687;
  assign n31689 = pi38 & ~n31686;
  assign n31690 = ~n31688 & n31689;
  assign n31691 = ~pi698 & ~n31690;
  assign n31692 = ~n31685 & n31691;
  assign n31693 = ~n31669 & ~n31692;
  assign n31694 = n9830 & ~n31693;
  assign n31695 = ~pi832 & ~n31645;
  assign n31696 = ~n31694 & n31695;
  assign po354 = ~n31644 & ~n31696;
  assign n31698 = n2531 & ~n16057;
  assign n31699 = n17793 & ~n31698;
  assign n31700 = pi198 & ~n31699;
  assign n31701 = pi198 & ~n16085;
  assign n31702 = pi198 & ~n16063;
  assign n31703 = ~po1101 & ~n31702;
  assign n31704 = n31701 & ~n31703;
  assign n31705 = n6161 & ~n16079;
  assign n31706 = ~n6161 & ~n16081;
  assign n31707 = pi198 & ~n31705;
  assign n31708 = ~n31706 & n31707;
  assign n31709 = ~n6221 & n31708;
  assign n31710 = ~n31704 & ~n31709;
  assign n31711 = pi215 & ~n31710;
  assign n31712 = n3302 & ~n31702;
  assign n31713 = pi198 & ~n16153;
  assign n31714 = ~n6221 & n31713;
  assign n31715 = pi198 & ~n16157;
  assign n31716 = po1101 & ~n31715;
  assign n31717 = ~n31703 & ~n31716;
  assign n31718 = n6221 & n31717;
  assign n31719 = ~n3302 & ~n31718;
  assign n31720 = ~n31714 & n31719;
  assign n31721 = ~pi215 & ~n31712;
  assign n31722 = ~n31720 & n31721;
  assign n31723 = pi299 & ~n31711;
  assign n31724 = ~n31722 & n31723;
  assign n31725 = ~n6194 & n31708;
  assign n31726 = ~n31704 & ~n31725;
  assign n31727 = pi223 & ~n31726;
  assign n31728 = n2608 & ~n31702;
  assign n31729 = ~n6194 & n31713;
  assign n31730 = n6194 & n31717;
  assign n31731 = ~n2608 & ~n31730;
  assign n31732 = ~n31729 & n31731;
  assign n31733 = ~pi223 & ~n31728;
  assign n31734 = ~n31732 & n31733;
  assign n31735 = ~pi299 & ~n31727;
  assign n31736 = ~n31734 & n31735;
  assign n31737 = pi39 & n2576;
  assign n31738 = ~n31724 & n31737;
  assign n31739 = ~n31736 & n31738;
  assign n31740 = ~n31700 & ~n31739;
  assign n31741 = ~n17585 & n31740;
  assign n31742 = pi198 & ~n9829;
  assign n31743 = pi634 & pi680;
  assign n31744 = pi198 & n16355;
  assign n31745 = ~n16341 & n31743;
  assign n31746 = ~n31744 & n31745;
  assign n31747 = ~n16054 & ~n31746;
  assign n31748 = ~pi299 & ~n31747;
  assign n31749 = ~pi198 & n16350;
  assign n31750 = pi198 & ~n16364;
  assign n31751 = ~n31749 & ~n31750;
  assign n31752 = n31743 & ~n31751;
  assign n31753 = pi198 & ~n16051;
  assign n31754 = ~n31743 & n31753;
  assign n31755 = ~n31752 & ~n31754;
  assign n31756 = pi299 & ~n31755;
  assign n31757 = ~pi39 & ~n31748;
  assign n31758 = ~n31756 & n31757;
  assign n31759 = ~n16294 & ~n31702;
  assign n31760 = n31743 & ~n31759;
  assign n31761 = ~n31702 & ~n31760;
  assign n31762 = n2608 & n31761;
  assign n31763 = pi634 & ~n31759;
  assign n31764 = ~n31702 & ~n31763;
  assign n31765 = n6166 & ~n31764;
  assign n31766 = pi198 & n16144;
  assign n31767 = pi634 & n16777;
  assign n31768 = ~n31766 & ~n31767;
  assign n31769 = ~n6166 & ~n31768;
  assign n31770 = ~n31765 & ~n31769;
  assign n31771 = n6164 & ~n31770;
  assign n31772 = n6161 & n31770;
  assign n31773 = ~n6161 & n31764;
  assign n31774 = n16672 & ~n31773;
  assign n31775 = ~n31772 & n31774;
  assign n31776 = ~n6161 & ~n31702;
  assign n31777 = n6161 & ~n31715;
  assign n31778 = ~pi680 & ~n31776;
  assign n31779 = ~n31777 & n31778;
  assign n31780 = ~n31771 & ~n31779;
  assign n31781 = ~n31775 & n31780;
  assign n31782 = n6194 & ~n31781;
  assign n31783 = pi198 & n16675;
  assign n31784 = n6164 & ~n31768;
  assign n31785 = n6161 & n31768;
  assign n31786 = ~n6166 & n31764;
  assign n31787 = n6166 & n31768;
  assign n31788 = ~n31786 & ~n31787;
  assign n31789 = ~n6161 & ~n31788;
  assign n31790 = n16672 & ~n31785;
  assign n31791 = ~n31789 & n31790;
  assign n31792 = ~n31783 & ~n31784;
  assign n31793 = ~n31791 & n31792;
  assign n31794 = ~n6194 & ~n31793;
  assign n31795 = ~n2608 & ~n31782;
  assign n31796 = ~n31794 & n31795;
  assign n31797 = ~pi223 & ~n31762;
  assign n31798 = ~n31796 & n31797;
  assign n31799 = ~pi680 & n31708;
  assign n31800 = n31701 & n31799;
  assign n31801 = pi198 & n16079;
  assign n31802 = pi634 & ~n16079;
  assign n31803 = n16294 & n31802;
  assign n31804 = ~n31801 & ~n31803;
  assign n31805 = ~n6166 & ~n31804;
  assign n31806 = ~n31765 & ~n31805;
  assign n31807 = n6161 & n31806;
  assign n31808 = n31774 & ~n31807;
  assign n31809 = n6164 & ~n31806;
  assign n31810 = ~n31800 & ~n31809;
  assign n31811 = ~n31808 & n31810;
  assign n31812 = n6194 & n31811;
  assign n31813 = n6164 & ~n31804;
  assign n31814 = n6161 & n31804;
  assign n31815 = n6166 & n31804;
  assign n31816 = ~n31786 & ~n31815;
  assign n31817 = ~n6161 & ~n31816;
  assign n31818 = n16672 & ~n31814;
  assign n31819 = ~n31817 & n31818;
  assign n31820 = ~n31799 & ~n31813;
  assign n31821 = ~n31819 & n31820;
  assign n31822 = ~n6194 & n31821;
  assign n31823 = pi223 & ~n31812;
  assign n31824 = ~n31822 & n31823;
  assign n31825 = ~n31798 & ~n31824;
  assign n31826 = ~pi299 & ~n31825;
  assign n31827 = n3302 & n31761;
  assign n31828 = ~n6221 & ~n31793;
  assign n31829 = n6221 & ~n31781;
  assign n31830 = ~n3302 & ~n31828;
  assign n31831 = ~n31829 & n31830;
  assign n31832 = ~pi215 & ~n31827;
  assign n31833 = ~n31831 & n31832;
  assign n31834 = n6221 & n31811;
  assign n31835 = ~n6221 & n31821;
  assign n31836 = pi215 & ~n31834;
  assign n31837 = ~n31835 & n31836;
  assign n31838 = ~n31833 & ~n31837;
  assign n31839 = pi299 & ~n31838;
  assign n31840 = pi39 & ~n31826;
  assign n31841 = ~n31839 & n31840;
  assign n31842 = ~n31758 & ~n31841;
  assign n31843 = ~pi38 & ~n31842;
  assign n31844 = pi198 & ~n16228;
  assign n31845 = pi38 & ~n31844;
  assign n31846 = pi634 & n15725;
  assign n31847 = n16228 & n31846;
  assign n31848 = n31845 & ~n31847;
  assign n31849 = n9829 & ~n31848;
  assign n31850 = ~n31843 & n31849;
  assign n31851 = ~n31742 & ~n31850;
  assign n31852 = ~pi778 & ~n31851;
  assign n31853 = ~pi625 & n31740;
  assign n31854 = pi625 & n31851;
  assign n31855 = pi1153 & ~n31853;
  assign n31856 = ~n31854 & n31855;
  assign n31857 = ~pi625 & n31851;
  assign n31858 = pi625 & n31740;
  assign n31859 = ~pi1153 & ~n31858;
  assign n31860 = ~n31857 & n31859;
  assign n31861 = ~n31856 & ~n31860;
  assign n31862 = pi778 & ~n31861;
  assign n31863 = ~n31852 & ~n31862;
  assign n31864 = ~n15741 & ~n31863;
  assign n31865 = n15741 & ~n31740;
  assign n31866 = ~n31864 & ~n31865;
  assign n31867 = ~n15747 & n31866;
  assign n31868 = n15747 & n31740;
  assign n31869 = ~n31867 & ~n31868;
  assign n31870 = ~n15753 & ~n31869;
  assign n31871 = ~n15759 & n31870;
  assign n31872 = ~n31741 & ~n31871;
  assign n31873 = ~pi792 & n31872;
  assign n31874 = ~pi628 & n31740;
  assign n31875 = pi628 & ~n31872;
  assign n31876 = pi1156 & ~n31874;
  assign n31877 = ~n31875 & n31876;
  assign n31878 = pi628 & n31740;
  assign n31879 = ~pi628 & ~n31872;
  assign n31880 = ~pi1156 & ~n31878;
  assign n31881 = ~n31879 & n31880;
  assign n31882 = ~n31877 & ~n31881;
  assign n31883 = pi792 & ~n31882;
  assign n31884 = ~n31873 & ~n31883;
  assign n31885 = n19394 & n31884;
  assign n31886 = ~n19394 & n31740;
  assign n31887 = ~n31885 & ~n31886;
  assign n31888 = ~n15959 & n31887;
  assign n31889 = n15832 & n31740;
  assign n31890 = ~n16435 & ~n16439;
  assign n31891 = pi633 & ~n31890;
  assign n31892 = ~n16054 & ~n31891;
  assign n31893 = ~n16444 & ~n31892;
  assign n31894 = ~pi299 & n31893;
  assign n31895 = pi603 & pi633;
  assign n31896 = ~n31753 & ~n31895;
  assign n31897 = pi198 & ~n16431;
  assign n31898 = ~pi198 & n16523;
  assign n31899 = ~n31897 & ~n31898;
  assign n31900 = n31895 & n31899;
  assign n31901 = ~n31896 & ~n31900;
  assign n31902 = pi299 & n31901;
  assign n31903 = ~pi39 & ~n31894;
  assign n31904 = ~n31902 & n31903;
  assign n31905 = pi633 & n16532;
  assign n31906 = ~n31708 & ~n31905;
  assign n31907 = ~n6164 & ~n31906;
  assign n31908 = pi633 & n16063;
  assign n31909 = ~n15779 & n31908;
  assign n31910 = ~n16079 & n31909;
  assign n31911 = ~n31801 & ~n31910;
  assign n31912 = n16492 & ~n31911;
  assign n31913 = ~n31907 & ~n31912;
  assign n31914 = ~n6194 & n31913;
  assign n31915 = ~n31702 & ~n31909;
  assign n31916 = pi603 & ~n31915;
  assign n31917 = pi198 & ~pi603;
  assign n31918 = ~n16063 & n31917;
  assign n31919 = ~n31916 & ~n31918;
  assign n31920 = ~n16452 & n31919;
  assign n31921 = n6166 & ~n31915;
  assign n31922 = ~n31701 & ~n31910;
  assign n31923 = ~n31921 & n31922;
  assign n31924 = pi603 & ~n31923;
  assign n31925 = n16452 & ~n31918;
  assign n31926 = ~n31924 & n31925;
  assign n31927 = ~n31920 & ~n31926;
  assign n31928 = ~n6164 & n31927;
  assign n31929 = ~n31701 & ~n31924;
  assign n31930 = n6164 & ~n31929;
  assign n31931 = ~n31928 & ~n31930;
  assign n31932 = n6194 & n31931;
  assign n31933 = pi223 & ~n31914;
  assign n31934 = ~n31932 & n31933;
  assign n31935 = pi642 & ~n31916;
  assign n31936 = ~n15779 & ~n16144;
  assign n31937 = pi633 & n31936;
  assign n31938 = ~n31766 & ~n31937;
  assign n31939 = ~n6166 & ~n31938;
  assign n31940 = ~n31921 & ~n31939;
  assign n31941 = pi603 & ~n31940;
  assign n31942 = ~pi642 & ~n31941;
  assign n31943 = n6160 & ~n31935;
  assign n31944 = ~n31942 & n31943;
  assign n31945 = ~n6160 & n31916;
  assign n31946 = ~n31918 & ~n31945;
  assign n31947 = ~n31944 & n31946;
  assign n31948 = ~n6164 & n31947;
  assign n31949 = ~pi603 & n31715;
  assign n31950 = n6164 & ~n31949;
  assign n31951 = ~n31941 & n31950;
  assign n31952 = ~n31948 & ~n31951;
  assign n31953 = n6194 & n31952;
  assign n31954 = n6161 & ~n31938;
  assign n31955 = n16146 & n31917;
  assign n31956 = n6166 & n31938;
  assign n31957 = ~n6166 & n31915;
  assign n31958 = pi603 & ~n16452;
  assign n31959 = ~n31957 & n31958;
  assign n31960 = ~n31956 & n31959;
  assign n31961 = ~n31954 & ~n31955;
  assign n31962 = ~n31960 & n31961;
  assign n31963 = ~n6164 & n31962;
  assign n31964 = pi603 & ~n31938;
  assign n31965 = n6164 & ~n31766;
  assign n31966 = ~n31964 & n31965;
  assign n31967 = ~n31963 & ~n31966;
  assign n31968 = ~n6194 & n31967;
  assign n31969 = ~n2608 & ~n31968;
  assign n31970 = ~n31953 & n31969;
  assign n31971 = n2608 & n31919;
  assign n31972 = ~pi223 & ~n31971;
  assign n31973 = ~n31970 & n31972;
  assign n31974 = ~n31934 & ~n31973;
  assign n31975 = ~pi299 & ~n31974;
  assign n31976 = ~n6221 & n31913;
  assign n31977 = n6221 & n31931;
  assign n31978 = pi215 & ~n31976;
  assign n31979 = ~n31977 & n31978;
  assign n31980 = n6221 & n31952;
  assign n31981 = ~n6221 & n31967;
  assign n31982 = ~n3302 & ~n31981;
  assign n31983 = ~n31980 & n31982;
  assign n31984 = n3302 & n31919;
  assign n31985 = ~pi215 & ~n31984;
  assign n31986 = ~n31983 & n31985;
  assign n31987 = ~n31979 & ~n31986;
  assign n31988 = pi299 & ~n31987;
  assign n31989 = pi39 & ~n31975;
  assign n31990 = ~n31988 & n31989;
  assign n31991 = ~n31904 & ~n31990;
  assign n31992 = ~pi38 & ~n31991;
  assign n31993 = pi633 & n15780;
  assign n31994 = n16228 & n31993;
  assign n31995 = n31845 & ~n31994;
  assign n31996 = n9829 & ~n31995;
  assign n31997 = ~n31992 & n31996;
  assign n31998 = ~n31742 & ~n31997;
  assign n31999 = ~n15777 & ~n31998;
  assign n32000 = n15777 & ~n31740;
  assign n32001 = ~n31999 & ~n32000;
  assign n32002 = ~pi785 & ~n32001;
  assign n32003 = ~n15786 & ~n31740;
  assign n32004 = pi609 & n31999;
  assign n32005 = ~n32003 & ~n32004;
  assign n32006 = pi1155 & ~n32005;
  assign n32007 = ~n16585 & ~n31740;
  assign n32008 = ~pi609 & n31999;
  assign n32009 = ~n32007 & ~n32008;
  assign n32010 = ~pi1155 & ~n32009;
  assign n32011 = ~n32006 & ~n32010;
  assign n32012 = pi785 & ~n32011;
  assign n32013 = ~n32002 & ~n32012;
  assign n32014 = ~pi781 & ~n32013;
  assign n32015 = ~pi618 & n31740;
  assign n32016 = pi618 & n32013;
  assign n32017 = pi1154 & ~n32015;
  assign n32018 = ~n32016 & n32017;
  assign n32019 = ~pi618 & n32013;
  assign n32020 = pi618 & n31740;
  assign n32021 = ~pi1154 & ~n32020;
  assign n32022 = ~n32019 & n32021;
  assign n32023 = ~n32018 & ~n32022;
  assign n32024 = pi781 & ~n32023;
  assign n32025 = ~n32014 & ~n32024;
  assign n32026 = ~pi789 & ~n32025;
  assign n32027 = ~pi619 & n31740;
  assign n32028 = pi619 & n32025;
  assign n32029 = pi1159 & ~n32027;
  assign n32030 = ~n32028 & n32029;
  assign n32031 = ~pi619 & n32025;
  assign n32032 = pi619 & n31740;
  assign n32033 = ~pi1159 & ~n32032;
  assign n32034 = ~n32031 & n32033;
  assign n32035 = ~n32030 & ~n32034;
  assign n32036 = pi789 & ~n32035;
  assign n32037 = ~n32026 & ~n32036;
  assign n32038 = ~n15832 & n32037;
  assign n32039 = ~n31889 & ~n32038;
  assign n32040 = ~n15925 & ~n32039;
  assign n32041 = n15925 & n31740;
  assign n32042 = n19478 & ~n32041;
  assign n32043 = ~n32040 & n32042;
  assign n32044 = ~n31888 & ~n32043;
  assign n32045 = pi787 & ~n32044;
  assign n32046 = ~n16633 & n32039;
  assign n32047 = ~pi629 & n31877;
  assign n32048 = pi629 & n31881;
  assign n32049 = ~n32047 & ~n32048;
  assign n32050 = ~n32046 & n32049;
  assign n32051 = n16644 & n32050;
  assign n32052 = pi792 & ~n32050;
  assign n32053 = n15753 & n31740;
  assign n32054 = ~n31870 & ~n32053;
  assign n32055 = n15828 & ~n32054;
  assign n32056 = pi626 & ~n31740;
  assign n32057 = ~pi626 & ~n32037;
  assign n32058 = n15757 & ~n32056;
  assign n32059 = ~n32057 & n32058;
  assign n32060 = ~pi626 & ~n31740;
  assign n32061 = pi626 & ~n32037;
  assign n32062 = n15756 & ~n32060;
  assign n32063 = ~n32061 & n32062;
  assign n32064 = ~n32055 & ~n32059;
  assign n32065 = ~n32063 & n32064;
  assign n32066 = pi788 & ~n32065;
  assign n32067 = pi609 & n31863;
  assign n32068 = pi634 & n17389;
  assign n32069 = n31995 & ~n32068;
  assign n32070 = ~pi680 & ~n31893;
  assign n32071 = ~pi603 & n31747;
  assign n32072 = pi634 & ~pi665;
  assign n32073 = pi198 & ~pi633;
  assign n32074 = n32072 & ~n32073;
  assign n32075 = ~n16434 & n32074;
  assign n32076 = ~pi634 & n16054;
  assign n32077 = pi634 & n16356;
  assign n32078 = ~n16441 & n32077;
  assign n32079 = ~n32076 & ~n32078;
  assign n32080 = ~pi633 & ~n32079;
  assign n32081 = pi603 & ~n32075;
  assign n32082 = ~n31891 & n32081;
  assign n32083 = ~n32080 & n32082;
  assign n32084 = ~n32071 & ~n32083;
  assign n32085 = pi680 & ~n32084;
  assign n32086 = ~pi299 & ~n32070;
  assign n32087 = ~n32085 & n32086;
  assign n32088 = ~n31743 & ~n31901;
  assign n32089 = ~pi603 & ~n31751;
  assign n32090 = ~n16523 & n31750;
  assign n32091 = ~pi198 & ~pi665;
  assign n32092 = n16431 & n32091;
  assign n32093 = ~pi633 & ~n32092;
  assign n32094 = ~n32090 & n32093;
  assign n32095 = pi198 & ~pi665;
  assign n32096 = pi633 & ~n32095;
  assign n32097 = ~n31749 & n32096;
  assign n32098 = n31899 & n32097;
  assign n32099 = pi603 & ~n32094;
  assign n32100 = ~n32098 & n32099;
  assign n32101 = n31743 & ~n32089;
  assign n32102 = ~n32100 & n32101;
  assign n32103 = pi299 & ~n32088;
  assign n32104 = ~n32102 & n32103;
  assign n32105 = ~pi39 & ~n32087;
  assign n32106 = ~n32104 & n32105;
  assign n32107 = n16664 & n31763;
  assign n32108 = n31971 & ~n32107;
  assign n32109 = ~pi680 & n31947;
  assign n32110 = ~pi603 & ~n31764;
  assign n32111 = n16454 & n32072;
  assign n32112 = n31915 & ~n32111;
  assign n32113 = pi603 & ~n32112;
  assign n32114 = ~n32110 & ~n32113;
  assign n32115 = ~n6160 & ~n32114;
  assign n32116 = n6166 & ~n32112;
  assign n32117 = pi634 & n16764;
  assign n32118 = n31938 & ~n32117;
  assign n32119 = ~n6166 & ~n32118;
  assign n32120 = ~n32116 & ~n32119;
  assign n32121 = pi603 & ~n32120;
  assign n32122 = ~pi642 & n32121;
  assign n32123 = pi642 & n32113;
  assign n32124 = ~n32110 & ~n32123;
  assign n32125 = ~n32122 & n32124;
  assign n32126 = n6160 & ~n32125;
  assign n32127 = ~n16108 & ~n32115;
  assign n32128 = ~n32126 & n32127;
  assign n32129 = ~pi603 & ~n31770;
  assign n32130 = n16108 & ~n32129;
  assign n32131 = ~n32121 & n32130;
  assign n32132 = ~n32128 & ~n32131;
  assign n32133 = pi680 & ~n32132;
  assign n32134 = ~n32109 & ~n32133;
  assign n32135 = n6194 & n32134;
  assign n32136 = ~pi680 & ~n31962;
  assign n32137 = ~pi603 & n31788;
  assign n32138 = ~n16452 & n32113;
  assign n32139 = ~n31959 & ~n32138;
  assign n32140 = ~n6161 & n32139;
  assign n32141 = ~n6166 & ~n32139;
  assign n32142 = n32118 & ~n32141;
  assign n32143 = ~n32140 & ~n32142;
  assign n32144 = ~n32137 & ~n32143;
  assign n32145 = n16672 & ~n32144;
  assign n32146 = ~n15780 & ~n31768;
  assign n32147 = ~n31964 & ~n32146;
  assign n32148 = n6164 & ~n32147;
  assign n32149 = ~n32136 & ~n32148;
  assign n32150 = ~n32145 & n32149;
  assign n32151 = ~n6194 & ~n32150;
  assign n32152 = ~n2608 & ~n32151;
  assign n32153 = ~n32135 & n32152;
  assign n32154 = ~pi223 & ~n32108;
  assign n32155 = ~n32153 & n32154;
  assign n32156 = ~pi680 & ~n31906;
  assign n32157 = n16475 & n32072;
  assign n32158 = n31911 & ~n32157;
  assign n32159 = ~n32140 & ~n32158;
  assign n32160 = ~pi603 & n31816;
  assign n32161 = ~n32141 & ~n32160;
  assign n32162 = ~n32159 & n32161;
  assign n32163 = n16672 & ~n32162;
  assign n32164 = ~pi603 & n31804;
  assign n32165 = pi603 & n32158;
  assign n32166 = n6164 & ~n32164;
  assign n32167 = ~n32165 & n32166;
  assign n32168 = ~n32156 & ~n32167;
  assign n32169 = ~n32163 & n32168;
  assign n32170 = ~n6194 & n32169;
  assign n32171 = pi634 & n16789;
  assign n32172 = ~n16452 & n32114;
  assign n32173 = ~n6166 & ~n32158;
  assign n32174 = ~n32116 & ~n32173;
  assign n32175 = pi603 & ~n32174;
  assign n32176 = n16452 & ~n32110;
  assign n32177 = ~n32175 & n32176;
  assign n32178 = n16672 & ~n32172;
  assign n32179 = ~n32177 & n32178;
  assign n32180 = ~pi680 & n31927;
  assign n32181 = ~n31930 & ~n32171;
  assign n32182 = ~n32179 & n32181;
  assign n32183 = ~n32180 & n32182;
  assign n32184 = n6194 & n32183;
  assign n32185 = pi223 & ~n32170;
  assign n32186 = ~n32184 & n32185;
  assign n32187 = ~n32155 & ~n32186;
  assign n32188 = ~pi299 & ~n32187;
  assign n32189 = n31984 & ~n32107;
  assign n32190 = n6221 & n32134;
  assign n32191 = ~n6221 & ~n32150;
  assign n32192 = ~n3302 & ~n32191;
  assign n32193 = ~n32190 & n32192;
  assign n32194 = ~pi215 & ~n32189;
  assign n32195 = ~n32193 & n32194;
  assign n32196 = ~n6221 & n32169;
  assign n32197 = n6221 & n32183;
  assign n32198 = pi215 & ~n32196;
  assign n32199 = ~n32197 & n32198;
  assign n32200 = ~n32195 & ~n32199;
  assign n32201 = pi299 & ~n32200;
  assign n32202 = pi39 & ~n32188;
  assign n32203 = ~n32201 & n32202;
  assign n32204 = ~n32106 & ~n32203;
  assign n32205 = ~pi38 & ~n32204;
  assign n32206 = n9829 & ~n32069;
  assign n32207 = ~n32205 & n32206;
  assign n32208 = ~n31742 & ~n32207;
  assign n32209 = ~pi625 & n32208;
  assign n32210 = pi625 & n31998;
  assign n32211 = ~pi1153 & ~n32210;
  assign n32212 = ~n32209 & n32211;
  assign n32213 = ~pi608 & ~n31856;
  assign n32214 = ~n32212 & n32213;
  assign n32215 = ~pi625 & n31998;
  assign n32216 = pi625 & n32208;
  assign n32217 = pi1153 & ~n32215;
  assign n32218 = ~n32216 & n32217;
  assign n32219 = pi608 & ~n31860;
  assign n32220 = ~n32218 & n32219;
  assign n32221 = ~n32214 & ~n32220;
  assign n32222 = pi778 & ~n32221;
  assign n32223 = ~pi778 & n32208;
  assign n32224 = ~n32222 & ~n32223;
  assign n32225 = ~pi609 & ~n32224;
  assign n32226 = ~pi1155 & ~n32067;
  assign n32227 = ~n32225 & n32226;
  assign n32228 = ~pi660 & ~n32006;
  assign n32229 = ~n32227 & n32228;
  assign n32230 = ~pi609 & n31863;
  assign n32231 = pi609 & ~n32224;
  assign n32232 = pi1155 & ~n32230;
  assign n32233 = ~n32231 & n32232;
  assign n32234 = pi660 & ~n32010;
  assign n32235 = ~n32233 & n32234;
  assign n32236 = ~n32229 & ~n32235;
  assign n32237 = pi785 & ~n32236;
  assign n32238 = ~pi785 & ~n32224;
  assign n32239 = ~n32237 & ~n32238;
  assign n32240 = ~pi618 & ~n32239;
  assign n32241 = pi618 & n31866;
  assign n32242 = ~pi1154 & ~n32241;
  assign n32243 = ~n32240 & n32242;
  assign n32244 = ~pi627 & ~n32018;
  assign n32245 = ~n32243 & n32244;
  assign n32246 = ~pi618 & n31866;
  assign n32247 = pi618 & ~n32239;
  assign n32248 = pi1154 & ~n32246;
  assign n32249 = ~n32247 & n32248;
  assign n32250 = pi627 & ~n32022;
  assign n32251 = ~n32249 & n32250;
  assign n32252 = ~n32245 & ~n32251;
  assign n32253 = pi781 & ~n32252;
  assign n32254 = ~pi781 & ~n32239;
  assign n32255 = ~n32253 & ~n32254;
  assign n32256 = ~pi789 & n32255;
  assign n32257 = ~pi619 & ~n31869;
  assign n32258 = pi619 & ~n32255;
  assign n32259 = pi1159 & ~n32257;
  assign n32260 = ~n32258 & n32259;
  assign n32261 = pi648 & ~n32034;
  assign n32262 = ~n32260 & n32261;
  assign n32263 = pi619 & ~n31869;
  assign n32264 = ~pi619 & ~n32255;
  assign n32265 = ~pi1159 & ~n32263;
  assign n32266 = ~n32264 & n32265;
  assign n32267 = ~pi648 & ~n32030;
  assign n32268 = ~n32266 & n32267;
  assign n32269 = pi789 & ~n32262;
  assign n32270 = ~n32268 & n32269;
  assign n32271 = n15833 & ~n32256;
  assign n32272 = ~n32270 & n32271;
  assign n32273 = ~n32066 & ~n32272;
  assign n32274 = ~n32052 & ~n32273;
  assign n32275 = n18841 & ~n32051;
  assign n32276 = ~n32274 & n32275;
  assign n32277 = ~n32045 & ~n32276;
  assign n32278 = ~pi790 & ~n32277;
  assign n32279 = pi787 & ~n31887;
  assign n32280 = ~pi787 & n31884;
  assign n32281 = ~n32279 & ~n32280;
  assign n32282 = ~pi644 & ~n32281;
  assign n32283 = pi644 & n32277;
  assign n32284 = pi715 & ~n32282;
  assign n32285 = ~n32283 & n32284;
  assign n32286 = ~n28954 & n31740;
  assign n32287 = n19771 & n32038;
  assign n32288 = ~n32286 & ~n32287;
  assign n32289 = pi644 & ~n32288;
  assign n32290 = ~pi644 & n31740;
  assign n32291 = ~pi715 & ~n32290;
  assign n32292 = ~n32289 & n32291;
  assign n32293 = pi1160 & ~n32292;
  assign n32294 = ~n32285 & n32293;
  assign n32295 = ~pi644 & ~n32288;
  assign n32296 = pi644 & n31740;
  assign n32297 = pi715 & ~n32296;
  assign n32298 = ~n32295 & n32297;
  assign n32299 = pi644 & ~n32281;
  assign n32300 = ~pi644 & n32277;
  assign n32301 = ~pi715 & ~n32299;
  assign n32302 = ~n32300 & n32301;
  assign n32303 = ~pi1160 & ~n32298;
  assign n32304 = ~n32302 & n32303;
  assign n32305 = pi790 & ~n32294;
  assign n32306 = ~n32304 & n32305;
  assign n32307 = ~n32278 & ~n32306;
  assign n32308 = ~po1038 & ~n32307;
  assign n32309 = pi198 & po1038;
  assign po355 = n32308 | n32309;
  assign n32311 = pi199 & ~n16219;
  assign n32312 = ~pi647 & ~n32311;
  assign n32313 = n15759 & ~n32311;
  assign n32314 = n15747 & ~n32311;
  assign n32315 = ~pi637 & ~n32311;
  assign n32316 = ~pi199 & ~n16228;
  assign n32317 = n19049 & ~n32316;
  assign n32318 = ~pi199 & ~n16335;
  assign n32319 = pi199 & n16291;
  assign n32320 = pi39 & ~n32318;
  assign n32321 = ~n32319 & n32320;
  assign n32322 = ~pi199 & ~n16353;
  assign n32323 = pi199 & n16368;
  assign n32324 = ~pi39 & ~n32322;
  assign n32325 = ~n32323 & n32324;
  assign n32326 = ~n32321 & ~n32325;
  assign n32327 = ~pi38 & ~n32326;
  assign n32328 = ~n32317 & ~n32327;
  assign n32329 = n9829 & ~n32328;
  assign n32330 = pi199 & ~n9829;
  assign n32331 = pi637 & ~n32330;
  assign n32332 = ~n32329 & n32331;
  assign n32333 = ~n32315 & ~n32332;
  assign n32334 = ~pi778 & n32333;
  assign n32335 = ~pi625 & ~n32311;
  assign n32336 = pi625 & ~n32333;
  assign n32337 = pi1153 & ~n32335;
  assign n32338 = ~n32336 & n32337;
  assign n32339 = ~pi625 & ~n32333;
  assign n32340 = pi625 & ~n32311;
  assign n32341 = ~pi1153 & ~n32340;
  assign n32342 = ~n32339 & n32341;
  assign n32343 = ~n32338 & ~n32342;
  assign n32344 = pi778 & ~n32343;
  assign n32345 = ~n32334 & ~n32344;
  assign n32346 = ~n15741 & ~n32345;
  assign n32347 = n15741 & n32311;
  assign n32348 = ~n32346 & ~n32347;
  assign n32349 = ~n15747 & n32348;
  assign n32350 = ~n32314 & ~n32349;
  assign n32351 = ~n15753 & n32350;
  assign n32352 = n15753 & n32311;
  assign n32353 = ~n32351 & ~n32352;
  assign n32354 = ~n15759 & n32353;
  assign n32355 = ~n32313 & ~n32354;
  assign n32356 = ~pi792 & n32355;
  assign n32357 = pi628 & n32355;
  assign n32358 = ~pi628 & n32311;
  assign n32359 = ~n32357 & ~n32358;
  assign n32360 = pi1156 & ~n32359;
  assign n32361 = pi628 & ~n32311;
  assign n32362 = ~pi628 & ~n32355;
  assign n32363 = ~pi1156 & ~n32361;
  assign n32364 = ~n32362 & n32363;
  assign n32365 = ~n32360 & ~n32364;
  assign n32366 = pi792 & ~n32365;
  assign n32367 = ~n32356 & ~n32366;
  assign n32368 = pi647 & n32367;
  assign n32369 = pi1157 & ~n32312;
  assign n32370 = ~n32368 & n32369;
  assign n32371 = ~pi629 & n32360;
  assign n32372 = pi619 & ~n32350;
  assign n32373 = ~pi1159 & ~n32372;
  assign n32374 = ~pi619 & ~n32311;
  assign n32375 = ~pi617 & ~n32311;
  assign n32376 = n9829 & n18604;
  assign n32377 = pi199 & ~n32376;
  assign n32378 = n9829 & ~n23191;
  assign n32379 = pi199 & ~n18598;
  assign n32380 = n32378 & ~n32379;
  assign n32381 = pi617 & ~n32377;
  assign n32382 = ~n32380 & n32381;
  assign n32383 = ~n32375 & ~n32382;
  assign n32384 = ~n15777 & n32383;
  assign n32385 = n15777 & n32311;
  assign n32386 = ~n32384 & ~n32385;
  assign n32387 = ~pi785 & ~n32386;
  assign n32388 = pi609 & n32386;
  assign n32389 = ~pi609 & ~n32311;
  assign n32390 = pi1155 & ~n32389;
  assign n32391 = ~n32388 & n32390;
  assign n32392 = ~pi609 & n32386;
  assign n32393 = pi609 & ~n32311;
  assign n32394 = ~pi1155 & ~n32393;
  assign n32395 = ~n32392 & n32394;
  assign n32396 = ~n32391 & ~n32395;
  assign n32397 = pi785 & ~n32396;
  assign n32398 = ~n32387 & ~n32397;
  assign n32399 = ~pi781 & ~n32398;
  assign n32400 = ~pi618 & ~n32311;
  assign n32401 = pi618 & n32398;
  assign n32402 = pi1154 & ~n32400;
  assign n32403 = ~n32401 & n32402;
  assign n32404 = pi618 & ~n32311;
  assign n32405 = ~pi618 & n32398;
  assign n32406 = ~pi1154 & ~n32404;
  assign n32407 = ~n32405 & n32406;
  assign n32408 = ~n32403 & ~n32407;
  assign n32409 = pi781 & ~n32408;
  assign n32410 = ~n32399 & ~n32409;
  assign n32411 = pi619 & n32410;
  assign n32412 = pi1159 & ~n32374;
  assign n32413 = ~n32411 & n32412;
  assign n32414 = ~pi648 & ~n32413;
  assign n32415 = ~n32373 & n32414;
  assign n32416 = ~pi619 & ~n32350;
  assign n32417 = pi1159 & ~n32416;
  assign n32418 = pi619 & ~n32311;
  assign n32419 = ~pi619 & n32410;
  assign n32420 = ~pi1159 & ~n32418;
  assign n32421 = ~n32419 & n32420;
  assign n32422 = pi648 & ~n32421;
  assign n32423 = ~n32417 & n32422;
  assign n32424 = ~n32415 & ~n32423;
  assign n32425 = pi789 & ~n32424;
  assign n32426 = pi619 & n32422;
  assign n32427 = ~pi619 & n32414;
  assign n32428 = pi789 & ~n32426;
  assign n32429 = ~n32427 & n32428;
  assign n32430 = pi609 & n32345;
  assign n32431 = ~pi637 & n32383;
  assign n32432 = n9829 & n18659;
  assign n32433 = ~pi199 & ~n32432;
  assign n32434 = pi199 & n18651;
  assign n32435 = pi617 & ~n32434;
  assign n32436 = ~n32433 & n32435;
  assign n32437 = n9829 & ~n23308;
  assign n32438 = ~pi199 & ~n32437;
  assign n32439 = pi199 & n18674;
  assign n32440 = ~pi617 & ~n18670;
  assign n32441 = ~n32438 & n32440;
  assign n32442 = ~n32439 & n32441;
  assign n32443 = ~n32330 & ~n32436;
  assign n32444 = ~n32442 & n32443;
  assign n32445 = pi637 & ~n32444;
  assign n32446 = ~n32431 & ~n32445;
  assign n32447 = ~pi625 & n32446;
  assign n32448 = pi625 & ~n32383;
  assign n32449 = ~pi1153 & ~n32448;
  assign n32450 = ~n32447 & n32449;
  assign n32451 = ~pi608 & ~n32338;
  assign n32452 = ~n32450 & n32451;
  assign n32453 = pi625 & n32446;
  assign n32454 = ~pi625 & ~n32383;
  assign n32455 = pi1153 & ~n32454;
  assign n32456 = ~n32453 & n32455;
  assign n32457 = pi608 & ~n32342;
  assign n32458 = ~n32456 & n32457;
  assign n32459 = ~n32452 & ~n32458;
  assign n32460 = pi778 & ~n32459;
  assign n32461 = ~pi778 & n32446;
  assign n32462 = ~n32460 & ~n32461;
  assign n32463 = ~pi609 & ~n32462;
  assign n32464 = ~pi1155 & ~n32430;
  assign n32465 = ~n32463 & n32464;
  assign n32466 = ~pi660 & ~n32391;
  assign n32467 = ~n32465 & n32466;
  assign n32468 = ~pi609 & n32345;
  assign n32469 = pi609 & ~n32462;
  assign n32470 = pi1155 & ~n32468;
  assign n32471 = ~n32469 & n32470;
  assign n32472 = pi660 & ~n32395;
  assign n32473 = ~n32471 & n32472;
  assign n32474 = ~n32467 & ~n32473;
  assign n32475 = pi785 & ~n32474;
  assign n32476 = ~pi785 & ~n32462;
  assign n32477 = ~n32475 & ~n32476;
  assign n32478 = ~pi781 & n32477;
  assign n32479 = ~pi618 & ~n32477;
  assign n32480 = pi618 & n32348;
  assign n32481 = ~pi1154 & ~n32480;
  assign n32482 = ~n32479 & n32481;
  assign n32483 = ~pi627 & ~n32403;
  assign n32484 = ~n32482 & n32483;
  assign n32485 = ~pi618 & n32348;
  assign n32486 = pi618 & ~n32477;
  assign n32487 = pi1154 & ~n32485;
  assign n32488 = ~n32486 & n32487;
  assign n32489 = pi627 & ~n32407;
  assign n32490 = ~n32488 & n32489;
  assign n32491 = pi781 & ~n32484;
  assign n32492 = ~n32490 & n32491;
  assign n32493 = ~n32429 & ~n32478;
  assign n32494 = ~n32492 & n32493;
  assign n32495 = ~n32425 & ~n32494;
  assign n32496 = n15833 & ~n32495;
  assign n32497 = pi641 & n32311;
  assign n32498 = ~pi641 & ~n32353;
  assign n32499 = n15819 & ~n32497;
  assign n32500 = ~n32498 & n32499;
  assign n32501 = ~pi789 & ~n32410;
  assign n32502 = ~n32413 & ~n32421;
  assign n32503 = pi789 & ~n32502;
  assign n32504 = ~n32501 & ~n32503;
  assign n32505 = n22348 & n32504;
  assign n32506 = ~pi641 & n32311;
  assign n32507 = pi641 & ~n32353;
  assign n32508 = n15818 & ~n32506;
  assign n32509 = ~n32507 & n32508;
  assign n32510 = ~n32500 & ~n32509;
  assign n32511 = ~n32505 & n32510;
  assign n32512 = pi788 & ~n32511;
  assign n32513 = ~n32496 & ~n32512;
  assign n32514 = ~n16643 & n32513;
  assign n32515 = ~n15832 & ~n32504;
  assign n32516 = n15832 & n32311;
  assign n32517 = ~n32515 & ~n32516;
  assign n32518 = ~n16633 & ~n32517;
  assign n32519 = pi629 & n32364;
  assign n32520 = ~n32371 & ~n32519;
  assign n32521 = ~n32518 & n32520;
  assign n32522 = ~n32514 & n32521;
  assign n32523 = pi792 & ~n32522;
  assign n32524 = ~pi792 & n32513;
  assign n32525 = ~n32523 & ~n32524;
  assign n32526 = ~pi647 & n32525;
  assign n32527 = ~n15925 & ~n32517;
  assign n32528 = n15925 & n32311;
  assign n32529 = ~n32527 & ~n32528;
  assign n32530 = pi647 & n32529;
  assign n32531 = ~pi1157 & ~n32530;
  assign n32532 = ~n32526 & n32531;
  assign n32533 = ~pi630 & ~n32370;
  assign n32534 = ~n32532 & n32533;
  assign n32535 = pi647 & ~n32311;
  assign n32536 = ~pi647 & n32367;
  assign n32537 = ~pi1157 & ~n32535;
  assign n32538 = ~n32536 & n32537;
  assign n32539 = ~pi647 & n32529;
  assign n32540 = pi647 & n32525;
  assign n32541 = pi1157 & ~n32539;
  assign n32542 = ~n32540 & n32541;
  assign n32543 = pi630 & ~n32538;
  assign n32544 = ~n32542 & n32543;
  assign n32545 = ~n32534 & ~n32544;
  assign n32546 = pi787 & ~n32545;
  assign n32547 = ~pi787 & n32525;
  assign n32548 = ~n32546 & ~n32547;
  assign n32549 = ~pi790 & n32548;
  assign n32550 = ~pi787 & ~n32367;
  assign n32551 = ~n32370 & ~n32538;
  assign n32552 = pi787 & ~n32551;
  assign n32553 = ~n32550 & ~n32552;
  assign n32554 = ~pi644 & n32553;
  assign n32555 = pi644 & ~n32548;
  assign n32556 = pi715 & ~n32554;
  assign n32557 = ~n32555 & n32556;
  assign n32558 = ~n15960 & ~n32529;
  assign n32559 = n15960 & n32311;
  assign n32560 = ~n32558 & ~n32559;
  assign n32561 = pi644 & n32560;
  assign n32562 = ~pi644 & ~n32311;
  assign n32563 = ~pi715 & ~n32562;
  assign n32564 = ~n32561 & n32563;
  assign n32565 = pi1160 & ~n32564;
  assign n32566 = ~n32557 & n32565;
  assign n32567 = ~pi644 & n32560;
  assign n32568 = pi644 & ~n32311;
  assign n32569 = pi715 & ~n32568;
  assign n32570 = ~n32567 & n32569;
  assign n32571 = pi644 & n32553;
  assign n32572 = ~pi644 & ~n32548;
  assign n32573 = ~pi715 & ~n32571;
  assign n32574 = ~n32572 & n32573;
  assign n32575 = ~pi1160 & ~n32570;
  assign n32576 = ~n32574 & n32575;
  assign n32577 = pi790 & ~n32566;
  assign n32578 = ~n32576 & n32577;
  assign n32579 = ~n32549 & ~n32578;
  assign n32580 = ~po1038 & ~n32579;
  assign n32581 = pi199 & po1038;
  assign po356 = n32580 | n32581;
  assign n32583 = pi200 & ~n16219;
  assign n32584 = ~pi606 & ~n32583;
  assign n32585 = pi200 & ~n32376;
  assign n32586 = pi200 & ~n18598;
  assign n32587 = n32378 & ~n32586;
  assign n32588 = pi606 & ~n32585;
  assign n32589 = ~n32587 & n32588;
  assign n32590 = ~n32584 & ~n32589;
  assign n32591 = ~n15777 & n32590;
  assign n32592 = n15777 & n32583;
  assign n32593 = ~n32591 & ~n32592;
  assign n32594 = ~pi785 & ~n32593;
  assign n32595 = pi609 & n32593;
  assign n32596 = ~pi609 & ~n32583;
  assign n32597 = pi1155 & ~n32596;
  assign n32598 = ~n32595 & n32597;
  assign n32599 = ~pi609 & n32593;
  assign n32600 = pi609 & ~n32583;
  assign n32601 = ~pi1155 & ~n32600;
  assign n32602 = ~n32599 & n32601;
  assign n32603 = ~n32598 & ~n32602;
  assign n32604 = pi785 & ~n32603;
  assign n32605 = ~n32594 & ~n32604;
  assign n32606 = ~pi781 & ~n32605;
  assign n32607 = ~pi618 & ~n32583;
  assign n32608 = pi618 & n32605;
  assign n32609 = pi1154 & ~n32607;
  assign n32610 = ~n32608 & n32609;
  assign n32611 = pi618 & ~n32583;
  assign n32612 = ~pi618 & n32605;
  assign n32613 = ~pi1154 & ~n32611;
  assign n32614 = ~n32612 & n32613;
  assign n32615 = ~n32610 & ~n32614;
  assign n32616 = pi781 & ~n32615;
  assign n32617 = ~n32606 & ~n32616;
  assign n32618 = ~pi789 & ~n32617;
  assign n32619 = ~pi619 & ~n32583;
  assign n32620 = pi619 & n32617;
  assign n32621 = pi1159 & ~n32619;
  assign n32622 = ~n32620 & n32621;
  assign n32623 = pi619 & ~n32583;
  assign n32624 = ~pi619 & n32617;
  assign n32625 = ~pi1159 & ~n32623;
  assign n32626 = ~n32624 & n32625;
  assign n32627 = ~n32622 & ~n32626;
  assign n32628 = pi789 & ~n32627;
  assign n32629 = ~n32618 & ~n32628;
  assign n32630 = ~n15832 & ~n32629;
  assign n32631 = n15832 & n32583;
  assign n32632 = ~n32630 & ~n32631;
  assign n32633 = ~n15925 & ~n32632;
  assign n32634 = n15925 & n32583;
  assign n32635 = ~n32633 & ~n32634;
  assign n32636 = ~n15960 & ~n32635;
  assign n32637 = n15960 & n32583;
  assign n32638 = ~n32636 & ~n32637;
  assign n32639 = ~pi644 & n32638;
  assign n32640 = pi644 & ~n32583;
  assign n32641 = pi715 & ~n32640;
  assign n32642 = ~n32639 & n32641;
  assign n32643 = n19478 & ~n32635;
  assign n32644 = ~n19394 & n32583;
  assign n32645 = n15747 & ~n32583;
  assign n32646 = ~pi643 & ~n32583;
  assign n32647 = ~pi200 & ~n16228;
  assign n32648 = n19049 & ~n32647;
  assign n32649 = ~pi200 & n16333;
  assign n32650 = pi200 & n16276;
  assign n32651 = ~pi299 & ~n32649;
  assign n32652 = ~n32650 & n32651;
  assign n32653 = ~pi200 & ~n16320;
  assign n32654 = pi200 & n16289;
  assign n32655 = pi299 & ~n32653;
  assign n32656 = ~n32654 & n32655;
  assign n32657 = ~n32652 & ~n32656;
  assign n32658 = pi39 & ~n32657;
  assign n32659 = ~pi200 & ~n16353;
  assign n32660 = pi200 & n16368;
  assign n32661 = ~pi39 & ~n32659;
  assign n32662 = ~n32660 & n32661;
  assign n32663 = ~n32658 & ~n32662;
  assign n32664 = ~pi38 & ~n32663;
  assign n32665 = ~n32648 & ~n32664;
  assign n32666 = n9829 & ~n32665;
  assign n32667 = pi200 & ~n9829;
  assign n32668 = pi643 & ~n32667;
  assign n32669 = ~n32666 & n32668;
  assign n32670 = ~n32646 & ~n32669;
  assign n32671 = ~pi778 & n32670;
  assign n32672 = ~pi625 & ~n32583;
  assign n32673 = pi625 & ~n32670;
  assign n32674 = pi1153 & ~n32672;
  assign n32675 = ~n32673 & n32674;
  assign n32676 = ~pi625 & ~n32670;
  assign n32677 = pi625 & ~n32583;
  assign n32678 = ~pi1153 & ~n32677;
  assign n32679 = ~n32676 & n32678;
  assign n32680 = ~n32675 & ~n32679;
  assign n32681 = pi778 & ~n32680;
  assign n32682 = ~n32671 & ~n32681;
  assign n32683 = ~n15741 & ~n32682;
  assign n32684 = n15741 & n32583;
  assign n32685 = ~n32683 & ~n32684;
  assign n32686 = ~n15747 & n32685;
  assign n32687 = ~n32645 & ~n32686;
  assign n32688 = ~n15753 & n32687;
  assign n32689 = n15753 & n32583;
  assign n32690 = ~n32688 & ~n32689;
  assign n32691 = ~n15759 & ~n32690;
  assign n32692 = n15759 & n32583;
  assign n32693 = ~n32691 & ~n32692;
  assign n32694 = ~pi792 & ~n32693;
  assign n32695 = ~pi628 & ~n32583;
  assign n32696 = pi628 & n32693;
  assign n32697 = pi1156 & ~n32695;
  assign n32698 = ~n32696 & n32697;
  assign n32699 = ~pi628 & n32693;
  assign n32700 = pi628 & ~n32583;
  assign n32701 = ~pi1156 & ~n32700;
  assign n32702 = ~n32699 & n32701;
  assign n32703 = ~n32698 & ~n32702;
  assign n32704 = pi792 & ~n32703;
  assign n32705 = ~n32694 & ~n32704;
  assign n32706 = n19394 & ~n32705;
  assign n32707 = ~n32644 & ~n32706;
  assign n32708 = ~n15959 & ~n32707;
  assign n32709 = ~n32643 & ~n32708;
  assign n32710 = pi787 & ~n32709;
  assign n32711 = ~n16633 & ~n32632;
  assign n32712 = ~pi629 & n32698;
  assign n32713 = pi629 & n32702;
  assign n32714 = ~n32712 & ~n32713;
  assign n32715 = ~n32711 & n32714;
  assign n32716 = pi792 & ~n32715;
  assign n32717 = n15828 & n32690;
  assign n32718 = ~pi626 & n32583;
  assign n32719 = pi626 & ~n32629;
  assign n32720 = n15756 & ~n32718;
  assign n32721 = ~n32719 & n32720;
  assign n32722 = pi626 & n32583;
  assign n32723 = ~pi626 & ~n32629;
  assign n32724 = n15757 & ~n32722;
  assign n32725 = ~n32723 & n32724;
  assign n32726 = ~n32717 & ~n32721;
  assign n32727 = ~n32725 & n32726;
  assign n32728 = pi788 & ~n32727;
  assign n32729 = pi609 & n32682;
  assign n32730 = ~pi643 & n32590;
  assign n32731 = ~n18669 & n32648;
  assign n32732 = ~pi200 & ~n18665;
  assign n32733 = pi200 & n18673;
  assign n32734 = ~pi38 & ~n32732;
  assign n32735 = ~n32733 & n32734;
  assign n32736 = ~n32731 & ~n32735;
  assign n32737 = ~pi606 & n9829;
  assign n32738 = ~n32736 & n32737;
  assign n32739 = ~n18654 & ~n18655;
  assign n32740 = ~pi200 & ~n32739;
  assign n32741 = pi200 & n18596;
  assign n32742 = n16808 & n32741;
  assign n32743 = ~pi200 & ~n18656;
  assign n32744 = pi200 & ~n23714;
  assign n32745 = ~pi38 & ~n32743;
  assign n32746 = ~n32744 & n32745;
  assign n32747 = pi606 & n9829;
  assign n32748 = ~n32742 & n32747;
  assign n32749 = ~n32740 & n32748;
  assign n32750 = ~n32746 & n32749;
  assign n32751 = ~n32667 & ~n32750;
  assign n32752 = ~n32738 & n32751;
  assign n32753 = pi643 & ~n32752;
  assign n32754 = ~n32730 & ~n32753;
  assign n32755 = ~pi625 & n32754;
  assign n32756 = pi625 & ~n32590;
  assign n32757 = ~pi1153 & ~n32756;
  assign n32758 = ~n32755 & n32757;
  assign n32759 = ~pi608 & ~n32675;
  assign n32760 = ~n32758 & n32759;
  assign n32761 = pi625 & n32754;
  assign n32762 = ~pi625 & ~n32590;
  assign n32763 = pi1153 & ~n32762;
  assign n32764 = ~n32761 & n32763;
  assign n32765 = pi608 & ~n32679;
  assign n32766 = ~n32764 & n32765;
  assign n32767 = ~n32760 & ~n32766;
  assign n32768 = pi778 & ~n32767;
  assign n32769 = ~pi778 & n32754;
  assign n32770 = ~n32768 & ~n32769;
  assign n32771 = ~pi609 & ~n32770;
  assign n32772 = ~pi1155 & ~n32729;
  assign n32773 = ~n32771 & n32772;
  assign n32774 = ~pi660 & ~n32598;
  assign n32775 = ~n32773 & n32774;
  assign n32776 = ~pi609 & n32682;
  assign n32777 = pi609 & ~n32770;
  assign n32778 = pi1155 & ~n32776;
  assign n32779 = ~n32777 & n32778;
  assign n32780 = pi660 & ~n32602;
  assign n32781 = ~n32779 & n32780;
  assign n32782 = ~n32775 & ~n32781;
  assign n32783 = pi785 & ~n32782;
  assign n32784 = ~pi785 & ~n32770;
  assign n32785 = ~n32783 & ~n32784;
  assign n32786 = ~pi618 & ~n32785;
  assign n32787 = pi618 & n32685;
  assign n32788 = ~pi1154 & ~n32787;
  assign n32789 = ~n32786 & n32788;
  assign n32790 = ~pi627 & ~n32610;
  assign n32791 = ~n32789 & n32790;
  assign n32792 = ~pi618 & n32685;
  assign n32793 = pi618 & ~n32785;
  assign n32794 = pi1154 & ~n32792;
  assign n32795 = ~n32793 & n32794;
  assign n32796 = pi627 & ~n32614;
  assign n32797 = ~n32795 & n32796;
  assign n32798 = ~n32791 & ~n32797;
  assign n32799 = pi781 & ~n32798;
  assign n32800 = ~pi781 & ~n32785;
  assign n32801 = ~n32799 & ~n32800;
  assign n32802 = ~pi789 & n32801;
  assign n32803 = ~pi619 & ~n32687;
  assign n32804 = pi619 & ~n32801;
  assign n32805 = pi1159 & ~n32803;
  assign n32806 = ~n32804 & n32805;
  assign n32807 = pi648 & ~n32626;
  assign n32808 = ~n32806 & n32807;
  assign n32809 = pi619 & ~n32687;
  assign n32810 = ~pi619 & ~n32801;
  assign n32811 = ~pi1159 & ~n32809;
  assign n32812 = ~n32810 & n32811;
  assign n32813 = ~pi648 & ~n32622;
  assign n32814 = ~n32812 & n32813;
  assign n32815 = pi789 & ~n32808;
  assign n32816 = ~n32814 & n32815;
  assign n32817 = n15833 & ~n32802;
  assign n32818 = ~n32816 & n32817;
  assign n32819 = ~n16644 & ~n32728;
  assign n32820 = ~n32818 & n32819;
  assign n32821 = ~n32716 & ~n32820;
  assign n32822 = n18841 & ~n32821;
  assign n32823 = ~n32710 & ~n32822;
  assign n32824 = ~pi644 & n32823;
  assign n32825 = ~n17768 & ~n32705;
  assign n32826 = pi787 & n32644;
  assign n32827 = ~n32825 & ~n32826;
  assign n32828 = pi644 & n32827;
  assign n32829 = ~pi715 & ~n32828;
  assign n32830 = ~n32824 & n32829;
  assign n32831 = ~pi1160 & ~n32642;
  assign n32832 = ~n32830 & n32831;
  assign n32833 = pi644 & n32638;
  assign n32834 = ~pi644 & ~n32583;
  assign n32835 = ~pi715 & ~n32834;
  assign n32836 = ~n32833 & n32835;
  assign n32837 = ~pi644 & n32827;
  assign n32838 = pi644 & n32823;
  assign n32839 = pi715 & ~n32837;
  assign n32840 = ~n32838 & n32839;
  assign n32841 = pi1160 & ~n32836;
  assign n32842 = ~n32840 & n32841;
  assign n32843 = ~n32832 & ~n32842;
  assign n32844 = pi790 & ~n32843;
  assign n32845 = ~pi790 & n32823;
  assign n32846 = ~n32844 & ~n32845;
  assign n32847 = ~po1038 & ~n32846;
  assign n32848 = ~pi200 & po1038;
  assign po357 = ~n32847 & ~n32848;
  assign n32850 = pi233 & pi237;
  assign n32851 = ~pi332 & ~n6161;
  assign n32852 = ~pi947 & ~n32851;
  assign n32853 = pi96 & pi210;
  assign n32854 = pi332 & n32853;
  assign n32855 = ~pi70 & ~pi841;
  assign n32856 = pi32 & ~n32855;
  assign n32857 = ~pi32 & ~pi70;
  assign n32858 = ~n32856 & ~n32857;
  assign n32859 = ~pi210 & n32858;
  assign n32860 = ~pi32 & ~pi96;
  assign n32861 = pi70 & n32860;
  assign n32862 = ~pi332 & ~n32861;
  assign n32863 = ~n32859 & n32862;
  assign n32864 = ~n32854 & ~n32863;
  assign n32865 = ~n6166 & n32864;
  assign n32866 = n6161 & ~n32865;
  assign n32867 = n32852 & ~n32866;
  assign n32868 = n6161 & ~n32864;
  assign n32869 = pi332 & pi468;
  assign n32870 = ~pi468 & ~n32863;
  assign n32871 = ~n32869 & ~n32870;
  assign n32872 = ~n6161 & n32871;
  assign n32873 = pi947 & ~n32868;
  assign n32874 = ~n32872 & n32873;
  assign n32875 = ~n32867 & ~n32874;
  assign n32876 = pi57 & ~n32875;
  assign n32877 = ~n6257 & n32875;
  assign n32878 = ~n2577 & n32875;
  assign n32879 = ~pi95 & n2701;
  assign n32880 = ~pi96 & ~n32856;
  assign n32881 = n32879 & n32880;
  assign n32882 = n2966 & n32881;
  assign n32883 = ~n32858 & ~n32882;
  assign n32884 = ~pi210 & ~n32883;
  assign n32885 = ~pi95 & n2967;
  assign n32886 = ~pi70 & ~n32885;
  assign n32887 = n32860 & ~n32886;
  assign n32888 = pi210 & n32887;
  assign n32889 = ~pi332 & ~n32884;
  assign n32890 = ~n32888 & n32889;
  assign n32891 = ~n32854 & ~n32890;
  assign n32892 = ~n6166 & n32891;
  assign n32893 = n6161 & ~n32892;
  assign n32894 = n32852 & ~n32893;
  assign n32895 = n6161 & ~n32891;
  assign n32896 = ~pi468 & ~n32890;
  assign n32897 = ~n32869 & ~n32896;
  assign n32898 = ~n6161 & n32897;
  assign n32899 = pi947 & ~n32895;
  assign n32900 = ~n32898 & n32899;
  assign n32901 = ~n32894 & ~n32900;
  assign n32902 = n2577 & n32901;
  assign n32903 = ~n32878 & ~n32902;
  assign n32904 = n6257 & ~n32903;
  assign n32905 = pi59 & ~n32877;
  assign n32906 = ~n32904 & n32905;
  assign n32907 = ~n2530 & n32875;
  assign n32908 = pi55 & n32903;
  assign n32909 = ~pi74 & n2616;
  assign n32910 = pi299 & ~n32875;
  assign n32911 = pi96 & pi198;
  assign n32912 = pi332 & n32911;
  assign n32913 = ~pi198 & n32858;
  assign n32914 = n32862 & ~n32913;
  assign n32915 = ~n32912 & ~n32914;
  assign n32916 = n6161 & ~n32915;
  assign n32917 = n6535 & ~n32914;
  assign n32918 = n32851 & ~n32917;
  assign n32919 = ~pi299 & ~n6534;
  assign n32920 = ~n32916 & n32919;
  assign n32921 = ~n32918 & n32920;
  assign n32922 = ~n32909 & ~n32921;
  assign n32923 = ~n32910 & n32922;
  assign n32924 = n2509 & n2726;
  assign n32925 = n32881 & n32924;
  assign n32926 = ~n32858 & ~n32925;
  assign n32927 = ~pi198 & ~n32926;
  assign n32928 = n32879 & n32924;
  assign n32929 = ~pi70 & ~n32928;
  assign n32930 = n32860 & ~n32929;
  assign n32931 = pi198 & n32930;
  assign n32932 = ~pi332 & ~n32927;
  assign n32933 = ~n32931 & n32932;
  assign n32934 = ~n32912 & ~n32933;
  assign n32935 = n6161 & ~n32934;
  assign n32936 = ~pi468 & ~n32933;
  assign n32937 = ~n6161 & ~n32869;
  assign n32938 = ~n32936 & n32937;
  assign n32939 = pi587 & ~n32938;
  assign n32940 = pi468 & n6161;
  assign n32941 = ~pi332 & ~n32940;
  assign n32942 = ~pi587 & ~n32941;
  assign n32943 = ~n32939 & ~n32942;
  assign n32944 = ~n32935 & ~n32943;
  assign n32945 = ~pi299 & ~n32944;
  assign n32946 = ~pi210 & ~n32926;
  assign n32947 = pi210 & n32930;
  assign n32948 = ~pi332 & ~n32946;
  assign n32949 = ~n32947 & n32948;
  assign n32950 = ~n32854 & ~n32949;
  assign n32951 = ~n6166 & n32950;
  assign n32952 = n6161 & ~n32951;
  assign n32953 = n32852 & ~n32952;
  assign n32954 = n6161 & ~n32950;
  assign n32955 = ~pi468 & ~n32949;
  assign n32956 = n32937 & ~n32955;
  assign n32957 = pi947 & ~n32954;
  assign n32958 = ~n32956 & n32957;
  assign n32959 = pi299 & ~n32953;
  assign n32960 = ~n32958 & n32959;
  assign n32961 = ~n32945 & ~n32960;
  assign n32962 = n9779 & ~n32961;
  assign n32963 = pi299 & ~n32901;
  assign n32964 = ~pi198 & ~n32883;
  assign n32965 = pi198 & n32887;
  assign n32966 = ~pi332 & ~n32964;
  assign n32967 = ~n32965 & n32966;
  assign n32968 = ~n32912 & ~n32967;
  assign n32969 = n6161 & ~n32968;
  assign n32970 = ~pi468 & ~n32967;
  assign n32971 = n32937 & ~n32970;
  assign n32972 = pi587 & ~n32971;
  assign n32973 = ~n32942 & ~n32972;
  assign n32974 = ~pi299 & ~n32969;
  assign n32975 = ~n32973 & n32974;
  assign n32976 = n14757 & ~n32975;
  assign n32977 = ~n32963 & n32976;
  assign n32978 = ~n32962 & ~n32977;
  assign n32979 = ~pi74 & ~n32978;
  assign n32980 = ~pi55 & ~n32923;
  assign n32981 = ~n32979 & n32980;
  assign n32982 = n2530 & ~n32908;
  assign n32983 = ~n32981 & n32982;
  assign n32984 = ~pi59 & ~n32907;
  assign n32985 = ~n32983 & n32984;
  assign n32986 = ~n32906 & ~n32985;
  assign n32987 = ~pi57 & ~n32986;
  assign n32988 = ~n32876 & ~n32987;
  assign n32989 = n32850 & ~n32988;
  assign n32990 = pi57 & pi332;
  assign n32991 = n2577 & n6525;
  assign n32992 = n2523 & n32991;
  assign n32993 = ~pi332 & ~n32992;
  assign n32994 = n6257 & ~n32993;
  assign n32995 = pi332 & ~n6257;
  assign n32996 = pi59 & ~n32995;
  assign n32997 = ~n32994 & n32996;
  assign n32998 = pi332 & ~n2530;
  assign n32999 = ~pi59 & ~n32998;
  assign n33000 = pi74 & pi332;
  assign n33001 = ~pi55 & ~n33000;
  assign n33002 = n2523 & n6537;
  assign n33003 = ~pi332 & ~n33002;
  assign n33004 = n14757 & ~n33003;
  assign n33005 = ~pi299 & pi587;
  assign n33006 = ~n19973 & ~n33005;
  assign n33007 = ~pi468 & ~n33006;
  assign n33008 = ~n32940 & ~n33007;
  assign n33009 = n2726 & n10688;
  assign n33010 = ~n33008 & n33009;
  assign n33011 = ~pi332 & ~n33010;
  assign n33012 = n9779 & ~n33011;
  assign n33013 = pi332 & ~n2616;
  assign n33014 = ~n33004 & ~n33013;
  assign n33015 = ~n33012 & n33014;
  assign n33016 = ~pi74 & ~n33015;
  assign n33017 = n33001 & ~n33016;
  assign n33018 = pi55 & n32993;
  assign n33019 = n2530 & ~n33018;
  assign n33020 = ~n33017 & n33019;
  assign n33021 = n32999 & ~n33020;
  assign n33022 = ~pi57 & ~n32997;
  assign n33023 = ~n33021 & n33022;
  assign n33024 = ~n32990 & ~n33023;
  assign n33025 = ~n32850 & ~n33024;
  assign n33026 = ~n32989 & ~n33025;
  assign n33027 = ~pi201 & ~n33026;
  assign n33028 = ~n6525 & ~n15574;
  assign n33029 = n6535 & n32911;
  assign n33030 = n15574 & ~n33029;
  assign n33031 = ~n15574 & ~n32853;
  assign n33032 = ~n33028 & ~n33030;
  assign n33033 = ~n33031 & n33032;
  assign n33034 = n32850 & n33033;
  assign n33035 = pi201 & ~n33034;
  assign po358 = ~n33027 & ~n33035;
  assign n33037 = ~pi233 & pi237;
  assign n33038 = ~n32988 & n33037;
  assign n33039 = ~n33024 & ~n33037;
  assign n33040 = ~n33038 & ~n33039;
  assign n33041 = ~pi202 & ~n33040;
  assign n33042 = n33033 & n33037;
  assign n33043 = pi202 & ~n33042;
  assign po359 = ~n33041 & ~n33043;
  assign n33045 = ~pi233 & ~pi237;
  assign n33046 = ~n32988 & n33045;
  assign n33047 = ~n33024 & ~n33045;
  assign n33048 = ~n33046 & ~n33047;
  assign n33049 = ~pi203 & ~n33048;
  assign n33050 = n33033 & n33045;
  assign n33051 = pi203 & ~n33050;
  assign po360 = ~n33049 & ~n33051;
  assign n33053 = ~pi332 & ~n6164;
  assign n33054 = ~pi907 & ~n33053;
  assign n33055 = n6164 & ~n32865;
  assign n33056 = n33054 & ~n33055;
  assign n33057 = n6164 & ~n32864;
  assign n33058 = ~n6164 & n32871;
  assign n33059 = pi907 & ~n33057;
  assign n33060 = ~n33058 & n33059;
  assign n33061 = ~n33056 & ~n33060;
  assign n33062 = pi57 & ~n33061;
  assign n33063 = ~n6257 & n33061;
  assign n33064 = ~n2577 & n33061;
  assign n33065 = n6164 & ~n32891;
  assign n33066 = ~n6164 & n32897;
  assign n33067 = pi907 & ~n33065;
  assign n33068 = ~n33066 & n33067;
  assign n33069 = pi332 & ~n16108;
  assign n33070 = pi680 & ~n33069;
  assign n33071 = ~n32892 & n33070;
  assign n33072 = n33054 & ~n33071;
  assign n33073 = ~n33068 & ~n33072;
  assign n33074 = n2577 & n33073;
  assign n33075 = ~n33064 & ~n33074;
  assign n33076 = n6257 & ~n33075;
  assign n33077 = pi59 & ~n33063;
  assign n33078 = ~n33076 & n33077;
  assign n33079 = ~n2530 & n33061;
  assign n33080 = pi55 & n33075;
  assign n33081 = pi299 & n33073;
  assign n33082 = n6164 & n32911;
  assign n33083 = pi332 & ~n33082;
  assign n33084 = ~pi299 & ~n33083;
  assign n33085 = n6279 & n32968;
  assign n33086 = n33084 & ~n33085;
  assign n33087 = ~n33081 & ~n33086;
  assign n33088 = n14757 & ~n33087;
  assign n33089 = n6279 & n32934;
  assign n33090 = n33084 & ~n33089;
  assign n33091 = n6263 & n32930;
  assign n33092 = pi299 & n33061;
  assign n33093 = ~n33091 & n33092;
  assign n33094 = ~n33090 & ~n33093;
  assign n33095 = n9779 & ~n33094;
  assign n33096 = ~n33088 & ~n33095;
  assign n33097 = ~pi74 & ~n33096;
  assign n33098 = pi299 & ~n33061;
  assign n33099 = ~pi468 & pi602;
  assign n33100 = pi468 & n6164;
  assign n33101 = ~n33099 & ~n33100;
  assign n33102 = n32915 & ~n33101;
  assign n33103 = ~n33083 & ~n33102;
  assign n33104 = ~pi299 & ~n33103;
  assign n33105 = ~n32909 & ~n33104;
  assign n33106 = ~n33098 & n33105;
  assign n33107 = ~pi55 & ~n33106;
  assign n33108 = ~n33097 & n33107;
  assign n33109 = n2530 & ~n33080;
  assign n33110 = ~n33108 & n33109;
  assign n33111 = ~pi59 & ~n33079;
  assign n33112 = ~n33110 & n33111;
  assign n33113 = ~n33078 & ~n33112;
  assign n33114 = ~pi57 & ~n33113;
  assign n33115 = ~n33062 & ~n33114;
  assign n33116 = n32850 & ~n33115;
  assign n33117 = n2577 & n6263;
  assign n33118 = n2523 & n33117;
  assign n33119 = ~pi332 & ~n33118;
  assign n33120 = n6257 & ~n33119;
  assign n33121 = n32996 & ~n33120;
  assign n33122 = pi55 & n33119;
  assign n33123 = ~pi299 & ~n33101;
  assign n33124 = ~n6277 & ~n33123;
  assign n33125 = n2523 & ~n33124;
  assign n33126 = ~pi332 & ~n33125;
  assign n33127 = n14757 & ~n33126;
  assign n33128 = ~pi299 & ~pi602;
  assign n33129 = pi299 & ~pi907;
  assign n33130 = ~pi468 & ~n33128;
  assign n33131 = ~n33129 & n33130;
  assign n33132 = ~n33100 & ~n33131;
  assign n33133 = n33009 & ~n33132;
  assign n33134 = ~pi332 & ~n33133;
  assign n33135 = n9779 & ~n33134;
  assign n33136 = ~n33127 & ~n33135;
  assign n33137 = ~pi74 & ~n33136;
  assign n33138 = n33001 & ~n33013;
  assign n33139 = ~n33137 & n33138;
  assign n33140 = n2530 & ~n33122;
  assign n33141 = ~n33139 & n33140;
  assign n33142 = n32999 & ~n33141;
  assign n33143 = ~pi57 & ~n33121;
  assign n33144 = ~n33142 & n33143;
  assign n33145 = ~n32990 & ~n33144;
  assign n33146 = ~n32850 & ~n33145;
  assign n33147 = ~n33116 & ~n33146;
  assign n33148 = ~pi204 & ~n33147;
  assign n33149 = ~n6263 & ~n15574;
  assign n33150 = n6279 & n32911;
  assign n33151 = n15574 & ~n33150;
  assign n33152 = ~n33031 & ~n33149;
  assign n33153 = ~n33151 & n33152;
  assign n33154 = n32850 & n33153;
  assign n33155 = pi204 & ~n33154;
  assign po361 = ~n33148 & ~n33155;
  assign n33157 = n33037 & ~n33115;
  assign n33158 = ~n33037 & ~n33145;
  assign n33159 = ~n33157 & ~n33158;
  assign n33160 = ~pi205 & ~n33159;
  assign n33161 = n33037 & n33153;
  assign n33162 = pi205 & ~n33161;
  assign po362 = ~n33160 & ~n33162;
  assign n33164 = pi233 & ~pi237;
  assign n33165 = ~n33115 & n33164;
  assign n33166 = ~n33145 & ~n33164;
  assign n33167 = ~n33165 & ~n33166;
  assign n33168 = ~pi206 & ~n33167;
  assign n33169 = n33153 & n33164;
  assign n33170 = pi206 & ~n33169;
  assign po363 = ~n33168 & ~n33170;
  assign n33172 = ~n15777 & n32378;
  assign n33173 = ~n18861 & n33172;
  assign n33174 = ~n18869 & n33173;
  assign n33175 = ~n18865 & n33174;
  assign n33176 = ~n15832 & n33175;
  assign n33177 = ~n15925 & n33176;
  assign n33178 = pi207 & ~n33177;
  assign n33179 = n15777 & ~n16219;
  assign n33180 = ~n15777 & ~n32376;
  assign n33181 = ~n33179 & ~n33180;
  assign n33182 = ~pi785 & ~n33181;
  assign n33183 = ~n16219 & ~n16585;
  assign n33184 = ~pi609 & n33180;
  assign n33185 = ~n33183 & ~n33184;
  assign n33186 = ~pi1155 & ~n33185;
  assign n33187 = ~n15786 & ~n16219;
  assign n33188 = pi609 & n33180;
  assign n33189 = ~n33187 & ~n33188;
  assign n33190 = pi1155 & ~n33189;
  assign n33191 = ~n33186 & ~n33190;
  assign n33192 = pi785 & ~n33191;
  assign n33193 = ~n33182 & ~n33192;
  assign n33194 = ~pi781 & ~n33193;
  assign n33195 = ~pi618 & n33193;
  assign n33196 = pi618 & n16219;
  assign n33197 = ~pi1154 & ~n33196;
  assign n33198 = ~n33195 & n33197;
  assign n33199 = ~pi618 & n16219;
  assign n33200 = pi618 & n33193;
  assign n33201 = pi1154 & ~n33199;
  assign n33202 = ~n33200 & n33201;
  assign n33203 = ~n33198 & ~n33202;
  assign n33204 = pi781 & ~n33203;
  assign n33205 = ~n33194 & ~n33204;
  assign n33206 = ~pi789 & ~n33205;
  assign n33207 = ~pi619 & n33205;
  assign n33208 = pi619 & n16219;
  assign n33209 = ~pi1159 & ~n33208;
  assign n33210 = ~n33207 & n33209;
  assign n33211 = ~pi619 & n16219;
  assign n33212 = pi619 & n33205;
  assign n33213 = pi1159 & ~n33211;
  assign n33214 = ~n33212 & n33213;
  assign n33215 = ~n33210 & ~n33214;
  assign n33216 = pi789 & ~n33215;
  assign n33217 = ~n33206 & ~n33216;
  assign n33218 = ~n15832 & n33217;
  assign n33219 = n15832 & n16219;
  assign n33220 = ~n33218 & ~n33219;
  assign n33221 = ~n15925 & ~n33220;
  assign n33222 = n15925 & n16219;
  assign n33223 = ~n33221 & ~n33222;
  assign n33224 = ~pi207 & ~n33223;
  assign n33225 = pi623 & ~n33178;
  assign n33226 = ~n33224 & n33225;
  assign n33227 = ~pi207 & ~n16219;
  assign n33228 = ~pi623 & n33227;
  assign n33229 = ~n33226 & ~n33228;
  assign n33230 = ~n15960 & ~n33229;
  assign n33231 = n15960 & n33227;
  assign n33232 = ~n33230 & ~n33231;
  assign n33233 = ~pi644 & ~n33232;
  assign n33234 = pi644 & n33227;
  assign n33235 = pi715 & ~n33234;
  assign n33236 = ~n33233 & n33235;
  assign n33237 = ~n17581 & n23147;
  assign n33238 = n17586 & n33237;
  assign n33239 = ~n15765 & n33238;
  assign n33240 = pi207 & ~n33239;
  assign n33241 = n15759 & ~n16219;
  assign n33242 = n15747 & ~n16219;
  assign n33243 = n9829 & n23150;
  assign n33244 = ~pi778 & ~n33243;
  assign n33245 = ~pi625 & ~n16219;
  assign n33246 = pi625 & ~n33243;
  assign n33247 = ~n33245 & ~n33246;
  assign n33248 = pi1153 & ~n33247;
  assign n33249 = pi625 & ~n16219;
  assign n33250 = ~pi625 & ~n33243;
  assign n33251 = ~n33249 & ~n33250;
  assign n33252 = ~pi1153 & ~n33251;
  assign n33253 = ~n33248 & ~n33252;
  assign n33254 = pi778 & ~n33253;
  assign n33255 = ~n33244 & ~n33254;
  assign n33256 = ~n15741 & n33255;
  assign n33257 = n15741 & n16219;
  assign n33258 = ~n33256 & ~n33257;
  assign n33259 = ~n15747 & n33258;
  assign n33260 = ~n33242 & ~n33259;
  assign n33261 = ~n15753 & n33260;
  assign n33262 = n15753 & n16219;
  assign n33263 = ~n33261 & ~n33262;
  assign n33264 = ~n15759 & n33263;
  assign n33265 = ~n33241 & ~n33264;
  assign n33266 = ~n15765 & ~n33265;
  assign n33267 = n15765 & ~n16219;
  assign n33268 = ~n33266 & ~n33267;
  assign n33269 = ~pi207 & n33268;
  assign n33270 = ~n33240 & ~n33269;
  assign n33271 = pi710 & ~n33270;
  assign n33272 = ~pi710 & ~n33227;
  assign n33273 = ~n33271 & ~n33272;
  assign n33274 = ~pi787 & ~n33273;
  assign n33275 = ~pi647 & n33273;
  assign n33276 = pi647 & n33227;
  assign n33277 = ~pi1157 & ~n33276;
  assign n33278 = ~n33275 & n33277;
  assign n33279 = ~pi647 & n33227;
  assign n33280 = pi647 & n33273;
  assign n33281 = pi1157 & ~n33279;
  assign n33282 = ~n33280 & n33281;
  assign n33283 = ~n33278 & ~n33282;
  assign n33284 = pi787 & ~n33283;
  assign n33285 = ~n33274 & ~n33284;
  assign n33286 = pi644 & n33285;
  assign n33287 = ~pi630 & n33282;
  assign n33288 = pi630 & n33278;
  assign n33289 = n19478 & n33229;
  assign n33290 = ~n33287 & ~n33288;
  assign n33291 = ~n33289 & n33290;
  assign n33292 = pi787 & ~n33291;
  assign n33293 = ~pi710 & ~n33229;
  assign n33294 = n17584 & n33237;
  assign n33295 = ~pi1159 & ~n33294;
  assign n33296 = pi1159 & ~n33174;
  assign n33297 = n21935 & ~n33295;
  assign n33298 = ~n33296 & n33297;
  assign n33299 = pi1159 & ~n33294;
  assign n33300 = ~pi1159 & ~n33174;
  assign n33301 = ~pi619 & pi648;
  assign n33302 = ~n33299 & n33301;
  assign n33303 = ~n33300 & n33302;
  assign n33304 = pi789 & ~n33298;
  assign n33305 = ~n33303 & n33304;
  assign n33306 = ~pi778 & ~n32432;
  assign n33307 = ~pi625 & n23147;
  assign n33308 = ~pi1153 & ~n33307;
  assign n33309 = pi608 & ~n33308;
  assign n33310 = ~pi625 & n32378;
  assign n33311 = pi625 & n32432;
  assign n33312 = pi1153 & ~n33310;
  assign n33313 = ~n33311 & n33312;
  assign n33314 = n33309 & ~n33313;
  assign n33315 = pi625 & n23147;
  assign n33316 = pi1153 & ~n33315;
  assign n33317 = ~pi608 & ~n33316;
  assign n33318 = ~pi625 & n32432;
  assign n33319 = pi625 & n32378;
  assign n33320 = ~pi1153 & ~n33319;
  assign n33321 = ~n33318 & n33320;
  assign n33322 = n33317 & ~n33321;
  assign n33323 = pi778 & ~n33314;
  assign n33324 = ~n33322 & n33323;
  assign n33325 = ~n33306 & ~n33324;
  assign n33326 = ~pi785 & ~n33325;
  assign n33327 = n18859 & n33172;
  assign n33328 = pi609 & ~n33237;
  assign n33329 = ~pi1155 & ~n33328;
  assign n33330 = ~pi609 & ~n33325;
  assign n33331 = n33329 & ~n33330;
  assign n33332 = ~pi660 & ~n33327;
  assign n33333 = ~n33331 & n33332;
  assign n33334 = n18858 & n33172;
  assign n33335 = ~pi609 & ~n33237;
  assign n33336 = pi1155 & ~n33335;
  assign n33337 = pi609 & ~n33325;
  assign n33338 = n33336 & ~n33337;
  assign n33339 = pi660 & ~n33334;
  assign n33340 = ~n33338 & n33339;
  assign n33341 = ~n33333 & ~n33340;
  assign n33342 = pi785 & ~n33341;
  assign n33343 = ~n33326 & ~n33342;
  assign n33344 = ~pi618 & ~pi627;
  assign n33345 = pi781 & ~n33344;
  assign n33346 = ~n33343 & ~n33345;
  assign n33347 = n18867 & n33173;
  assign n33348 = ~n15741 & n33237;
  assign n33349 = pi618 & ~n33348;
  assign n33350 = ~pi1154 & ~n33349;
  assign n33351 = ~pi627 & ~n33347;
  assign n33352 = ~n33350 & n33351;
  assign n33353 = n18866 & n33173;
  assign n33354 = ~pi618 & ~n33348;
  assign n33355 = pi618 & ~n33343;
  assign n33356 = pi1154 & ~n33354;
  assign n33357 = ~n33355 & n33356;
  assign n33358 = pi627 & ~n33353;
  assign n33359 = ~n33357 & n33358;
  assign n33360 = ~n33352 & ~n33359;
  assign n33361 = pi781 & ~n33360;
  assign n33362 = ~n33346 & ~n33361;
  assign n33363 = ~pi789 & ~n33362;
  assign n33364 = ~n33305 & ~n33363;
  assign n33365 = n22147 & n33362;
  assign n33366 = ~n33364 & ~n33365;
  assign n33367 = n15833 & ~n33366;
  assign n33368 = ~n15753 & n33294;
  assign n33369 = n15826 & n33368;
  assign n33370 = n15825 & n33175;
  assign n33371 = ~pi1158 & ~n33369;
  assign n33372 = ~n33370 & n33371;
  assign n33373 = n15826 & n33175;
  assign n33374 = n15825 & n33368;
  assign n33375 = pi1158 & ~n33373;
  assign n33376 = ~n33374 & n33375;
  assign n33377 = pi788 & ~n33372;
  assign n33378 = ~n33376 & n33377;
  assign n33379 = ~n33367 & ~n33378;
  assign n33380 = ~n16644 & ~n33379;
  assign n33381 = n16631 & n33176;
  assign n33382 = n16629 & n33238;
  assign n33383 = ~pi1156 & ~n33382;
  assign n33384 = ~n33381 & n33383;
  assign n33385 = n16631 & n33238;
  assign n33386 = n16629 & n33176;
  assign n33387 = pi1156 & ~n33385;
  assign n33388 = ~n33386 & n33387;
  assign n33389 = pi792 & ~n33384;
  assign n33390 = ~n33388 & n33389;
  assign n33391 = ~n33380 & ~n33390;
  assign n33392 = pi207 & ~n33391;
  assign n33393 = ~pi628 & ~n16219;
  assign n33394 = pi628 & ~n33265;
  assign n33395 = ~n33393 & ~n33394;
  assign n33396 = ~pi629 & ~n33395;
  assign n33397 = pi1156 & n33396;
  assign n33398 = ~n16633 & n33220;
  assign n33399 = pi628 & n16219;
  assign n33400 = ~pi628 & n33265;
  assign n33401 = n15923 & ~n33399;
  assign n33402 = ~n33400 & n33401;
  assign n33403 = ~n33397 & ~n33402;
  assign n33404 = ~n33398 & n33403;
  assign n33405 = pi792 & ~n33404;
  assign n33406 = pi641 & n33263;
  assign n33407 = ~pi641 & ~n16219;
  assign n33408 = pi1158 & ~n33407;
  assign n33409 = ~pi626 & n33408;
  assign n33410 = ~n33406 & n33409;
  assign n33411 = n22348 & n33217;
  assign n33412 = pi641 & ~n16219;
  assign n33413 = ~pi1158 & ~n33412;
  assign n33414 = ~pi641 & n33263;
  assign n33415 = pi626 & n33413;
  assign n33416 = ~n33414 & n33415;
  assign n33417 = ~n33410 & ~n33416;
  assign n33418 = ~n33411 & n33417;
  assign n33419 = pi788 & ~n33418;
  assign n33420 = pi618 & n33258;
  assign n33421 = pi609 & ~n33255;
  assign n33422 = n9829 & n18651;
  assign n33423 = ~pi778 & ~n33422;
  assign n33424 = ~pi608 & ~n33248;
  assign n33425 = ~pi625 & n33422;
  assign n33426 = pi625 & n32376;
  assign n33427 = ~pi1153 & ~n33425;
  assign n33428 = ~n33426 & n33427;
  assign n33429 = n33424 & ~n33428;
  assign n33430 = pi608 & ~n33252;
  assign n33431 = ~pi625 & n32376;
  assign n33432 = pi625 & n33422;
  assign n33433 = pi1153 & ~n33432;
  assign n33434 = ~n33431 & n33433;
  assign n33435 = n33430 & ~n33434;
  assign n33436 = pi778 & ~n33429;
  assign n33437 = ~n33435 & n33436;
  assign n33438 = ~n33423 & ~n33437;
  assign n33439 = ~pi609 & ~n33438;
  assign n33440 = ~n33421 & ~n33439;
  assign n33441 = ~pi1155 & ~n33440;
  assign n33442 = ~pi660 & ~n33190;
  assign n33443 = ~n33441 & n33442;
  assign n33444 = ~pi609 & ~n33255;
  assign n33445 = pi609 & ~n33438;
  assign n33446 = ~n33444 & ~n33445;
  assign n33447 = pi1155 & ~n33446;
  assign n33448 = pi660 & ~n33186;
  assign n33449 = ~n33447 & n33448;
  assign n33450 = ~n33443 & ~n33449;
  assign n33451 = pi785 & ~n33450;
  assign n33452 = ~pi785 & n33438;
  assign n33453 = ~n33451 & ~n33452;
  assign n33454 = ~pi618 & n33453;
  assign n33455 = ~n33420 & ~n33454;
  assign n33456 = ~pi1154 & ~n33455;
  assign n33457 = ~pi627 & ~n33202;
  assign n33458 = ~n33456 & n33457;
  assign n33459 = ~pi618 & n33258;
  assign n33460 = pi618 & n33453;
  assign n33461 = ~n33459 & ~n33460;
  assign n33462 = pi1154 & ~n33461;
  assign n33463 = pi627 & ~n33198;
  assign n33464 = ~n33462 & n33463;
  assign n33465 = ~n33458 & ~n33464;
  assign n33466 = pi781 & ~n33465;
  assign n33467 = ~pi781 & ~n33453;
  assign n33468 = ~n33466 & ~n33467;
  assign n33469 = ~pi789 & n33468;
  assign n33470 = pi619 & ~n33260;
  assign n33471 = ~pi619 & n33468;
  assign n33472 = ~n33470 & ~n33471;
  assign n33473 = ~pi1159 & ~n33472;
  assign n33474 = ~pi648 & ~n33214;
  assign n33475 = ~n33473 & n33474;
  assign n33476 = ~pi619 & ~n33260;
  assign n33477 = pi619 & n33468;
  assign n33478 = ~n33476 & ~n33477;
  assign n33479 = pi1159 & ~n33478;
  assign n33480 = pi648 & ~n33210;
  assign n33481 = ~n33479 & n33480;
  assign n33482 = pi789 & ~n33475;
  assign n33483 = ~n33481 & n33482;
  assign n33484 = n15833 & ~n33469;
  assign n33485 = ~n33483 & n33484;
  assign n33486 = ~n16644 & ~n33419;
  assign n33487 = ~n33485 & n33486;
  assign n33488 = ~n33405 & ~n33487;
  assign n33489 = ~pi207 & ~n33488;
  assign n33490 = pi623 & ~n33392;
  assign n33491 = ~n33489 & n33490;
  assign n33492 = n18892 & n33348;
  assign n33493 = ~pi660 & n33329;
  assign n33494 = pi609 & ~n33493;
  assign n33495 = pi660 & n33336;
  assign n33496 = ~pi609 & ~n33495;
  assign n33497 = pi785 & ~n33494;
  assign n33498 = ~n33496 & n33497;
  assign n33499 = ~pi778 & ~n32437;
  assign n33500 = pi625 & n32437;
  assign n33501 = pi1153 & ~n33500;
  assign n33502 = n33309 & ~n33501;
  assign n33503 = ~pi625 & n32437;
  assign n33504 = ~pi1153 & ~n33503;
  assign n33505 = n33317 & ~n33504;
  assign n33506 = pi778 & ~n33502;
  assign n33507 = ~n33505 & n33506;
  assign n33508 = pi785 & ~n33493;
  assign n33509 = ~n33495 & n33508;
  assign n33510 = ~n33499 & ~n33509;
  assign n33511 = ~n33507 & n33510;
  assign n33512 = ~n33498 & ~n33511;
  assign n33513 = n18893 & ~n33512;
  assign n33514 = ~n33492 & ~n33513;
  assign n33515 = ~n22148 & ~n33514;
  assign n33516 = n15752 & n18865;
  assign n33517 = n33294 & n33516;
  assign n33518 = ~n33515 & ~n33517;
  assign n33519 = n15833 & ~n33518;
  assign n33520 = ~n15827 & n15832;
  assign n33521 = n33368 & n33520;
  assign n33522 = ~n33519 & ~n33521;
  assign n33523 = ~n16644 & ~n33522;
  assign n33524 = n15764 & n15925;
  assign n33525 = n33238 & n33524;
  assign n33526 = ~n33523 & ~n33525;
  assign n33527 = pi207 & ~n33526;
  assign n33528 = ~n33393 & ~n33396;
  assign n33529 = pi1156 & ~n33528;
  assign n33530 = n15763 & ~n33399;
  assign n33531 = ~n33402 & ~n33530;
  assign n33532 = ~n33529 & n33531;
  assign n33533 = pi792 & ~n33532;
  assign n33534 = pi1159 & ~n16219;
  assign n33535 = pi1154 & ~n16219;
  assign n33536 = pi1155 & ~n16219;
  assign n33537 = n9829 & ~n18675;
  assign n33538 = ~pi778 & ~n33537;
  assign n33539 = pi625 & ~n33537;
  assign n33540 = ~n33245 & ~n33539;
  assign n33541 = pi1153 & ~n33540;
  assign n33542 = n33430 & ~n33541;
  assign n33543 = ~pi625 & ~n33537;
  assign n33544 = ~n33249 & ~n33543;
  assign n33545 = ~pi1153 & ~n33544;
  assign n33546 = n33424 & ~n33545;
  assign n33547 = pi778 & ~n33542;
  assign n33548 = ~n33546 & n33547;
  assign n33549 = ~n33538 & ~n33548;
  assign n33550 = ~pi609 & ~n33549;
  assign n33551 = ~n33421 & ~n33550;
  assign n33552 = ~pi1155 & ~n33551;
  assign n33553 = ~pi660 & ~n33536;
  assign n33554 = ~n33552 & n33553;
  assign n33555 = ~pi1155 & ~n16219;
  assign n33556 = pi609 & ~n33549;
  assign n33557 = ~n33444 & ~n33556;
  assign n33558 = pi1155 & ~n33557;
  assign n33559 = pi660 & ~n33555;
  assign n33560 = ~n33558 & n33559;
  assign n33561 = ~n33554 & ~n33560;
  assign n33562 = pi785 & ~n33561;
  assign n33563 = ~pi785 & n33549;
  assign n33564 = ~n33562 & ~n33563;
  assign n33565 = ~pi618 & n33564;
  assign n33566 = ~n33420 & ~n33565;
  assign n33567 = ~pi1154 & ~n33566;
  assign n33568 = ~pi627 & ~n33535;
  assign n33569 = ~n33567 & n33568;
  assign n33570 = ~pi1154 & ~n16219;
  assign n33571 = pi618 & n33564;
  assign n33572 = ~n33459 & ~n33571;
  assign n33573 = pi1154 & ~n33572;
  assign n33574 = pi627 & ~n33570;
  assign n33575 = ~n33573 & n33574;
  assign n33576 = ~n33569 & ~n33575;
  assign n33577 = pi781 & ~n33576;
  assign n33578 = ~pi781 & ~n33564;
  assign n33579 = ~n33577 & ~n33578;
  assign n33580 = ~pi619 & n33579;
  assign n33581 = ~n33470 & ~n33580;
  assign n33582 = ~pi1159 & ~n33581;
  assign n33583 = ~pi648 & ~n33534;
  assign n33584 = ~n33582 & n33583;
  assign n33585 = ~pi1159 & ~n16219;
  assign n33586 = pi619 & n33579;
  assign n33587 = ~n33476 & ~n33586;
  assign n33588 = pi1159 & ~n33587;
  assign n33589 = pi648 & ~n33585;
  assign n33590 = ~n33588 & n33589;
  assign n33591 = ~n33584 & ~n33590;
  assign n33592 = pi789 & ~n33591;
  assign n33593 = ~pi789 & ~n33579;
  assign n33594 = ~n33592 & ~n33593;
  assign n33595 = ~pi788 & ~n33594;
  assign n33596 = ~pi626 & ~n33594;
  assign n33597 = pi626 & ~n33263;
  assign n33598 = ~pi641 & ~n33597;
  assign n33599 = ~n33596 & n33598;
  assign n33600 = n33413 & ~n33599;
  assign n33601 = pi626 & ~n33594;
  assign n33602 = ~pi626 & ~n33263;
  assign n33603 = pi641 & ~n33602;
  assign n33604 = ~n33601 & n33603;
  assign n33605 = n33408 & ~n33604;
  assign n33606 = ~n33600 & ~n33605;
  assign n33607 = pi788 & ~n33606;
  assign n33608 = ~n16644 & ~n33595;
  assign n33609 = ~n33607 & n33608;
  assign n33610 = ~n33533 & ~n33609;
  assign n33611 = ~pi207 & ~n33610;
  assign n33612 = ~pi623 & ~n33527;
  assign n33613 = ~n33611 & n33612;
  assign n33614 = pi710 & ~n33491;
  assign n33615 = ~n33613 & n33614;
  assign n33616 = n18841 & ~n33293;
  assign n33617 = ~n33615 & n33616;
  assign n33618 = ~n33292 & ~n33617;
  assign n33619 = ~pi644 & n33618;
  assign n33620 = ~pi715 & ~n33286;
  assign n33621 = ~n33619 & n33620;
  assign n33622 = ~pi1160 & ~n33236;
  assign n33623 = ~n33621 & n33622;
  assign n33624 = ~pi644 & n33285;
  assign n33625 = pi644 & n33618;
  assign n33626 = pi715 & ~n33624;
  assign n33627 = ~n33625 & n33626;
  assign n33628 = pi644 & ~n33232;
  assign n33629 = ~pi644 & n33227;
  assign n33630 = ~pi715 & ~n33629;
  assign n33631 = ~n33628 & n33630;
  assign n33632 = pi1160 & ~n33631;
  assign n33633 = ~n33627 & n33632;
  assign n33634 = ~n33623 & ~n33633;
  assign n33635 = pi790 & ~n33634;
  assign n33636 = ~pi790 & n33618;
  assign n33637 = ~n33635 & ~n33636;
  assign n33638 = ~po1038 & ~n33637;
  assign n33639 = ~pi207 & po1038;
  assign po364 = n33638 | n33639;
  assign n33641 = pi208 & ~n33177;
  assign n33642 = ~pi208 & ~n33223;
  assign n33643 = pi607 & ~n33641;
  assign n33644 = ~n33642 & n33643;
  assign n33645 = ~pi208 & ~n16219;
  assign n33646 = ~pi607 & n33645;
  assign n33647 = ~n33644 & ~n33646;
  assign n33648 = ~n15960 & ~n33647;
  assign n33649 = n15960 & n33645;
  assign n33650 = ~n33648 & ~n33649;
  assign n33651 = ~pi644 & ~n33650;
  assign n33652 = pi644 & n33645;
  assign n33653 = pi715 & ~n33652;
  assign n33654 = ~n33651 & n33653;
  assign n33655 = pi208 & ~n33239;
  assign n33656 = ~pi208 & n33268;
  assign n33657 = ~n33655 & ~n33656;
  assign n33658 = pi638 & ~n33657;
  assign n33659 = ~pi638 & ~n33645;
  assign n33660 = ~n33658 & ~n33659;
  assign n33661 = ~pi787 & ~n33660;
  assign n33662 = ~pi647 & n33660;
  assign n33663 = pi647 & n33645;
  assign n33664 = ~pi1157 & ~n33663;
  assign n33665 = ~n33662 & n33664;
  assign n33666 = ~pi647 & n33645;
  assign n33667 = pi647 & n33660;
  assign n33668 = pi1157 & ~n33666;
  assign n33669 = ~n33667 & n33668;
  assign n33670 = ~n33665 & ~n33669;
  assign n33671 = pi787 & ~n33670;
  assign n33672 = ~n33661 & ~n33671;
  assign n33673 = pi644 & n33672;
  assign n33674 = ~pi630 & n33669;
  assign n33675 = pi630 & n33665;
  assign n33676 = n19478 & n33647;
  assign n33677 = ~n33674 & ~n33675;
  assign n33678 = ~n33676 & n33677;
  assign n33679 = pi787 & ~n33678;
  assign n33680 = ~pi638 & ~n33647;
  assign n33681 = pi208 & ~n33391;
  assign n33682 = ~pi208 & ~n33488;
  assign n33683 = pi607 & ~n33681;
  assign n33684 = ~n33682 & n33683;
  assign n33685 = pi208 & ~n33526;
  assign n33686 = ~pi208 & ~n33610;
  assign n33687 = ~pi607 & ~n33685;
  assign n33688 = ~n33686 & n33687;
  assign n33689 = pi638 & ~n33684;
  assign n33690 = ~n33688 & n33689;
  assign n33691 = n18841 & ~n33680;
  assign n33692 = ~n33690 & n33691;
  assign n33693 = ~n33679 & ~n33692;
  assign n33694 = ~pi644 & n33693;
  assign n33695 = ~pi715 & ~n33673;
  assign n33696 = ~n33694 & n33695;
  assign n33697 = ~pi1160 & ~n33654;
  assign n33698 = ~n33696 & n33697;
  assign n33699 = ~pi644 & n33672;
  assign n33700 = pi644 & n33693;
  assign n33701 = pi715 & ~n33699;
  assign n33702 = ~n33700 & n33701;
  assign n33703 = pi644 & ~n33650;
  assign n33704 = ~pi644 & n33645;
  assign n33705 = ~pi715 & ~n33704;
  assign n33706 = ~n33703 & n33705;
  assign n33707 = pi1160 & ~n33706;
  assign n33708 = ~n33702 & n33707;
  assign n33709 = ~n33698 & ~n33708;
  assign n33710 = pi790 & ~n33709;
  assign n33711 = ~pi790 & n33693;
  assign n33712 = ~n33710 & ~n33711;
  assign n33713 = ~po1038 & ~n33712;
  assign n33714 = ~pi208 & po1038;
  assign po365 = n33713 | n33714;
  assign n33716 = ~po1038 & n16219;
  assign n33717 = ~pi639 & n33716;
  assign n33718 = pi715 & n16219;
  assign n33719 = n18841 & ~n33610;
  assign n33720 = ~pi647 & ~n16219;
  assign n33721 = n19476 & ~n33268;
  assign n33722 = ~n33720 & ~n33721;
  assign n33723 = pi1157 & ~n33722;
  assign n33724 = pi647 & ~n16219;
  assign n33725 = n19475 & ~n33268;
  assign n33726 = ~n33724 & ~n33725;
  assign n33727 = ~pi1157 & ~n33726;
  assign n33728 = ~n33723 & ~n33727;
  assign n33729 = pi787 & ~n33728;
  assign n33730 = ~n33719 & ~n33729;
  assign n33731 = ~pi644 & ~n33730;
  assign n33732 = ~n17768 & n33268;
  assign n33733 = n16219 & n17768;
  assign n33734 = ~n33732 & ~n33733;
  assign n33735 = pi644 & n33734;
  assign n33736 = ~pi715 & ~n33735;
  assign n33737 = ~n33731 & n33736;
  assign n33738 = ~pi1160 & ~n33718;
  assign n33739 = ~n33737 & n33738;
  assign n33740 = ~pi715 & n16219;
  assign n33741 = pi644 & ~n33730;
  assign n33742 = ~pi644 & n33734;
  assign n33743 = pi715 & ~n33742;
  assign n33744 = ~n33741 & n33743;
  assign n33745 = pi1160 & ~n33740;
  assign n33746 = ~n33744 & n33745;
  assign n33747 = ~n33739 & ~n33746;
  assign n33748 = pi790 & ~n33747;
  assign n33749 = ~pi790 & ~n33730;
  assign n33750 = ~po1038 & ~n33749;
  assign n33751 = ~n33748 & n33750;
  assign n33752 = pi639 & n33751;
  assign n33753 = ~pi622 & ~n33717;
  assign n33754 = ~n33752 & n33753;
  assign n33755 = ~n15960 & ~n33223;
  assign n33756 = n15960 & n16219;
  assign n33757 = ~n33755 & ~n33756;
  assign n33758 = ~pi790 & n33757;
  assign n33759 = pi644 & ~n33757;
  assign n33760 = ~pi644 & n16219;
  assign n33761 = ~n33759 & ~n33760;
  assign n33762 = pi1160 & ~n33761;
  assign n33763 = ~pi644 & ~n33757;
  assign n33764 = pi644 & n16219;
  assign n33765 = ~n33763 & ~n33764;
  assign n33766 = ~pi1160 & ~n33765;
  assign n33767 = pi790 & ~n33762;
  assign n33768 = ~n33766 & n33767;
  assign n33769 = ~po1038 & ~n33758;
  assign n33770 = ~n33768 & n33769;
  assign n33771 = ~pi639 & n33770;
  assign n33772 = pi715 & ~n33765;
  assign n33773 = n18841 & ~n33488;
  assign n33774 = n19478 & n33223;
  assign n33775 = ~n15959 & ~n33728;
  assign n33776 = ~n33774 & ~n33775;
  assign n33777 = pi787 & ~n33776;
  assign n33778 = ~n33773 & ~n33777;
  assign n33779 = ~pi644 & ~n33778;
  assign n33780 = n33736 & ~n33779;
  assign n33781 = ~pi1160 & ~n33772;
  assign n33782 = ~n33780 & n33781;
  assign n33783 = ~pi715 & ~n33761;
  assign n33784 = pi644 & ~n33778;
  assign n33785 = n33743 & ~n33784;
  assign n33786 = pi1160 & ~n33783;
  assign n33787 = ~n33785 & n33786;
  assign n33788 = ~n33782 & ~n33787;
  assign n33789 = pi790 & ~n33788;
  assign n33790 = ~pi790 & ~n33778;
  assign n33791 = ~po1038 & ~n33790;
  assign n33792 = ~n33789 & n33791;
  assign n33793 = pi639 & n33792;
  assign n33794 = pi622 & ~n33771;
  assign n33795 = ~n33793 & n33794;
  assign n33796 = ~n33754 & ~n33795;
  assign n33797 = ~pi209 & ~n33796;
  assign n33798 = ~pi644 & pi1160;
  assign n33799 = ~n22949 & ~n33798;
  assign n33800 = pi790 & ~n33799;
  assign n33801 = n19771 & n33176;
  assign n33802 = ~po1038 & ~n33800;
  assign n33803 = n33801 & n33802;
  assign n33804 = pi622 & n33803;
  assign n33805 = ~pi639 & ~n33804;
  assign n33806 = n18841 & ~n33526;
  assign n33807 = n15960 & n19394;
  assign n33808 = n33239 & n33807;
  assign n33809 = ~n33806 & ~n33808;
  assign n33810 = ~pi790 & n33809;
  assign n33811 = ~n17768 & n33239;
  assign n33812 = ~pi644 & ~n33811;
  assign n33813 = pi715 & ~n33812;
  assign n33814 = pi644 & n33809;
  assign n33815 = pi1160 & n33813;
  assign n33816 = ~n33814 & n33815;
  assign n33817 = pi644 & ~n33811;
  assign n33818 = ~pi715 & ~n33817;
  assign n33819 = ~pi644 & n33809;
  assign n33820 = ~pi1160 & n33818;
  assign n33821 = ~n33819 & n33820;
  assign n33822 = pi790 & ~n33816;
  assign n33823 = ~n33821 & n33822;
  assign n33824 = ~po1038 & ~n33810;
  assign n33825 = ~n33823 & n33824;
  assign n33826 = ~pi622 & ~n33825;
  assign n33827 = ~pi644 & pi715;
  assign n33828 = n33801 & n33827;
  assign n33829 = ~pi1157 & ~n33239;
  assign n33830 = pi1157 & ~n33177;
  assign n33831 = n19475 & ~n33829;
  assign n33832 = ~n33830 & n33831;
  assign n33833 = pi1157 & ~n33239;
  assign n33834 = ~pi1157 & ~n33177;
  assign n33835 = n19476 & ~n33833;
  assign n33836 = ~n33834 & n33835;
  assign n33837 = ~n33832 & ~n33836;
  assign n33838 = pi787 & ~n33837;
  assign n33839 = n18841 & ~n33391;
  assign n33840 = ~n33838 & ~n33839;
  assign n33841 = ~pi644 & n33840;
  assign n33842 = n33818 & ~n33841;
  assign n33843 = ~pi1160 & ~n33828;
  assign n33844 = ~n33842 & n33843;
  assign n33845 = pi644 & ~pi715;
  assign n33846 = n33801 & n33845;
  assign n33847 = pi644 & n33840;
  assign n33848 = n33813 & ~n33847;
  assign n33849 = pi1160 & ~n33846;
  assign n33850 = ~n33848 & n33849;
  assign n33851 = ~n33844 & ~n33850;
  assign n33852 = pi790 & ~n33851;
  assign n33853 = ~pi790 & n33840;
  assign n33854 = ~po1038 & ~n33853;
  assign n33855 = ~n33852 & n33854;
  assign n33856 = pi622 & pi639;
  assign n33857 = ~n33855 & n33856;
  assign n33858 = pi209 & ~n33805;
  assign n33859 = ~n33826 & n33858;
  assign n33860 = ~n33857 & n33859;
  assign po366 = n33797 | n33860;
  assign n33862 = pi634 & n19798;
  assign n33863 = pi633 & pi947;
  assign n33864 = ~n33862 & ~n33863;
  assign n33865 = ~n16033 & ~n33864;
  assign n33866 = pi299 & ~n16050;
  assign n33867 = ~n33865 & n33866;
  assign n33868 = pi210 & ~n16055;
  assign n33869 = n16055 & ~n33864;
  assign n33870 = ~pi299 & ~n33868;
  assign n33871 = ~n33869 & n33870;
  assign n33872 = ~pi39 & ~n33867;
  assign n33873 = ~n33871 & n33872;
  assign n33874 = pi210 & ~n16063;
  assign n33875 = ~n31908 & ~n33874;
  assign n33876 = n6197 & n33875;
  assign n33877 = pi947 & ~n33876;
  assign n33878 = pi210 & n16079;
  assign n33879 = pi633 & ~n16079;
  assign n33880 = ~n33878 & ~n33879;
  assign n33881 = ~n6197 & n33880;
  assign n33882 = n33877 & ~n33881;
  assign n33883 = pi634 & n16063;
  assign n33884 = ~n33874 & ~n33883;
  assign n33885 = n6197 & n33884;
  assign n33886 = pi907 & ~n33885;
  assign n33887 = ~n31802 & ~n33878;
  assign n33888 = ~n6197 & n33887;
  assign n33889 = n33886 & ~n33888;
  assign n33890 = ~po1101 & n33874;
  assign n33891 = pi210 & po1101;
  assign n33892 = ~n16085 & n33891;
  assign n33893 = ~n33890 & ~n33892;
  assign n33894 = n6219 & n33893;
  assign n33895 = n6197 & n16062;
  assign n33896 = n2923 & n33895;
  assign n33897 = n33878 & ~n33896;
  assign n33898 = ~n6219 & ~n33897;
  assign n33899 = ~pi907 & ~n33898;
  assign n33900 = ~n33894 & n33899;
  assign n33901 = ~n33889 & ~n33900;
  assign n33902 = ~pi947 & ~n33901;
  assign n33903 = ~n33882 & ~n33902;
  assign n33904 = pi215 & ~n33903;
  assign n33905 = n16063 & ~n33864;
  assign n33906 = ~n33874 & ~n33905;
  assign n33907 = n3302 & n33906;
  assign n33908 = pi210 & n16144;
  assign n33909 = pi634 & ~n16144;
  assign n33910 = ~n33908 & ~n33909;
  assign n33911 = ~n6197 & n33910;
  assign n33912 = n33886 & ~n33911;
  assign n33913 = pi210 & ~n16153;
  assign n33914 = ~n6219 & ~n33913;
  assign n33915 = ~n16157 & n33891;
  assign n33916 = ~n33890 & ~n33915;
  assign n33917 = n6219 & n33916;
  assign n33918 = ~pi907 & ~n33917;
  assign n33919 = ~n33914 & n33918;
  assign n33920 = ~n33912 & ~n33919;
  assign n33921 = ~pi947 & ~n33920;
  assign n33922 = pi633 & ~n16144;
  assign n33923 = ~n33908 & ~n33922;
  assign n33924 = ~n6197 & n33923;
  assign n33925 = n33877 & ~n33924;
  assign n33926 = ~n3302 & ~n33925;
  assign n33927 = ~n33921 & n33926;
  assign n33928 = ~pi215 & ~n33907;
  assign n33929 = ~n33927 & n33928;
  assign n33930 = pi299 & ~n33904;
  assign n33931 = ~n33929 & n33930;
  assign n33932 = n2608 & n33906;
  assign n33933 = ~po1101 & n33875;
  assign n33934 = pi947 & ~n33933;
  assign n33935 = ~n6166 & ~n33923;
  assign n33936 = po1101 & n33875;
  assign n33937 = ~n6205 & ~n33936;
  assign n33938 = ~n33935 & ~n33937;
  assign n33939 = n33934 & ~n33938;
  assign n33940 = ~n6205 & ~n33884;
  assign n33941 = pi907 & ~n33940;
  assign n33942 = n6205 & ~n33910;
  assign n33943 = n33941 & ~n33942;
  assign n33944 = ~pi907 & n33916;
  assign n33945 = ~pi947 & ~n33943;
  assign n33946 = ~n33944 & n33945;
  assign n33947 = n6194 & ~n33939;
  assign n33948 = ~n33946 & n33947;
  assign n33949 = ~pi907 & n33913;
  assign n33950 = ~n33912 & ~n33949;
  assign n33951 = ~pi947 & ~n33950;
  assign n33952 = ~n6194 & ~n33925;
  assign n33953 = ~n33951 & n33952;
  assign n33954 = ~n33948 & ~n33953;
  assign n33955 = ~n2608 & ~n33954;
  assign n33956 = ~pi223 & ~n33932;
  assign n33957 = ~n33955 & n33956;
  assign n33958 = ~n33889 & ~n33897;
  assign n33959 = ~pi947 & ~n33958;
  assign n33960 = ~n6194 & ~n33882;
  assign n33961 = ~n33959 & n33960;
  assign n33962 = ~n6166 & ~n33880;
  assign n33963 = ~n33937 & ~n33962;
  assign n33964 = n33934 & ~n33963;
  assign n33965 = n6205 & ~n33887;
  assign n33966 = n33941 & ~n33965;
  assign n33967 = ~pi907 & n33893;
  assign n33968 = ~pi947 & ~n33966;
  assign n33969 = ~n33967 & n33968;
  assign n33970 = n6194 & ~n33964;
  assign n33971 = ~n33969 & n33970;
  assign n33972 = pi223 & ~n33961;
  assign n33973 = ~n33971 & n33972;
  assign n33974 = ~pi299 & ~n33973;
  assign n33975 = ~n33957 & n33974;
  assign n33976 = pi39 & ~n33931;
  assign n33977 = ~n33975 & n33976;
  assign n33978 = ~pi38 & ~n33873;
  assign n33979 = ~n33977 & n33978;
  assign n33980 = n16228 & ~n33864;
  assign n33981 = pi210 & ~n16228;
  assign n33982 = pi38 & ~n33980;
  assign n33983 = ~n33981 & n33982;
  assign n33984 = ~n33979 & ~n33983;
  assign n33985 = n9830 & ~n33984;
  assign n33986 = ~pi210 & ~n9830;
  assign po367 = ~n33985 & ~n33986;
  assign n33988 = n9829 & ~n20514;
  assign n33989 = ~pi606 & n33988;
  assign n33990 = n9829 & ~n20509;
  assign n33991 = pi606 & n33990;
  assign n33992 = pi643 & ~n33991;
  assign n33993 = ~n33989 & n33992;
  assign n33994 = n9829 & ~n19897;
  assign n33995 = pi606 & n33994;
  assign n33996 = n16218 & n32737;
  assign n33997 = ~pi643 & ~n33996;
  assign n33998 = ~n33995 & n33997;
  assign n33999 = ~po1038 & ~n33993;
  assign n34000 = ~n33998 & n33999;
  assign n34001 = pi211 & ~n34000;
  assign n34002 = n9829 & n20500;
  assign n34003 = ~pi606 & ~n34002;
  assign n34004 = n9829 & n20497;
  assign n34005 = pi606 & ~n34004;
  assign n34006 = pi643 & ~n34003;
  assign n34007 = ~n34005 & n34006;
  assign n34008 = n9829 & n19920;
  assign n34009 = pi606 & ~pi643;
  assign n34010 = n34008 & n34009;
  assign n34011 = ~n34007 & ~n34010;
  assign n34012 = ~pi211 & ~po1038;
  assign n34013 = ~n34011 & n34012;
  assign po368 = n34001 | n34013;
  assign n34015 = ~pi607 & n33988;
  assign n34016 = pi607 & n33990;
  assign n34017 = pi638 & ~n34016;
  assign n34018 = ~n34015 & n34017;
  assign n34019 = ~pi607 & n16219;
  assign n34020 = pi607 & n33994;
  assign n34021 = ~pi638 & ~n34019;
  assign n34022 = ~n34020 & n34021;
  assign n34023 = ~po1038 & ~n34018;
  assign n34024 = ~n34022 & n34023;
  assign n34025 = ~pi212 & ~n34024;
  assign n34026 = pi607 & ~n34004;
  assign n34027 = ~pi607 & ~n34002;
  assign n34028 = pi638 & ~n34026;
  assign n34029 = ~n34027 & n34028;
  assign n34030 = pi607 & ~pi638;
  assign n34031 = n34008 & n34030;
  assign n34032 = ~n34029 & ~n34031;
  assign n34033 = pi212 & ~po1038;
  assign n34034 = ~n34032 & n34033;
  assign po369 = n34025 | n34034;
  assign n34036 = pi213 & ~po1038;
  assign n34037 = pi622 & ~n34004;
  assign n34038 = ~pi622 & ~n34002;
  assign n34039 = pi639 & ~n34037;
  assign n34040 = ~n34038 & n34039;
  assign n34041 = pi622 & ~pi639;
  assign n34042 = n34008 & n34041;
  assign n34043 = ~n34040 & ~n34042;
  assign n34044 = n34036 & ~n34043;
  assign n34045 = ~pi639 & ~n33994;
  assign n34046 = pi639 & ~n33990;
  assign n34047 = pi622 & ~n34046;
  assign n34048 = ~n34045 & n34047;
  assign n34049 = ~pi639 & ~n16219;
  assign n34050 = pi639 & ~n33988;
  assign n34051 = ~pi622 & ~n34049;
  assign n34052 = ~n34050 & n34051;
  assign n34053 = ~n34048 & ~n34052;
  assign n34054 = ~po1038 & ~n34053;
  assign n34055 = ~pi213 & ~n34054;
  assign po370 = n34044 | n34055;
  assign n34057 = ~pi623 & n33988;
  assign n34058 = pi623 & n33990;
  assign n34059 = pi710 & ~n34058;
  assign n34060 = ~n34057 & n34059;
  assign n34061 = ~pi623 & n16219;
  assign n34062 = pi623 & n33994;
  assign n34063 = ~pi710 & ~n34061;
  assign n34064 = ~n34062 & n34063;
  assign n34065 = ~po1038 & ~n34060;
  assign n34066 = ~n34064 & n34065;
  assign n34067 = ~pi214 & ~n34066;
  assign n34068 = pi623 & ~n34004;
  assign n34069 = ~pi623 & ~n34002;
  assign n34070 = pi710 & ~n34068;
  assign n34071 = ~n34069 & n34070;
  assign n34072 = pi623 & ~pi710;
  assign n34073 = n34008 & n34072;
  assign n34074 = ~n34071 & ~n34073;
  assign n34075 = pi214 & ~po1038;
  assign n34076 = ~n34074 & n34075;
  assign po371 = n34067 | n34076;
  assign n34078 = pi215 & ~n9830;
  assign n34079 = pi215 & ~n16228;
  assign n34080 = pi681 & pi907;
  assign n34081 = ~pi947 & n34080;
  assign n34082 = pi642 & pi947;
  assign n34083 = ~n34081 & ~n34082;
  assign n34084 = n16228 & ~n34083;
  assign n34085 = pi38 & ~n34079;
  assign n34086 = ~n34084 & n34085;
  assign n34087 = ~pi215 & ~n16051;
  assign n34088 = n16051 & n34083;
  assign n34089 = pi299 & ~n34087;
  assign n34090 = ~n34088 & n34089;
  assign n34091 = ~pi215 & ~n16055;
  assign n34092 = n16055 & n34083;
  assign n34093 = ~pi299 & ~n34091;
  assign n34094 = ~n34092 & n34093;
  assign n34095 = ~n34090 & ~n34094;
  assign n34096 = ~pi39 & ~n34095;
  assign n34097 = n6162 & n16097;
  assign n34098 = ~n6164 & ~n16089;
  assign n34099 = ~pi642 & ~n34097;
  assign n34100 = ~n34098 & n34099;
  assign n34101 = ~n6194 & ~n34100;
  assign n34102 = ~pi642 & ~n16116;
  assign n34103 = ~n16117 & n34102;
  assign n34104 = n6194 & ~n34103;
  assign n34105 = pi947 & ~n34101;
  assign n34106 = ~n34104 & n34105;
  assign n34107 = ~n20314 & ~n34106;
  assign n34108 = pi223 & ~n34081;
  assign n34109 = ~n34107 & n34108;
  assign n34110 = ~pi642 & n16153;
  assign n34111 = ~n6194 & ~n34110;
  assign n34112 = ~n6164 & n16887;
  assign n34113 = ~n6160 & n16063;
  assign n34114 = ~n6164 & ~n34113;
  assign n34115 = n6164 & ~n16157;
  assign n34116 = ~pi642 & ~n34114;
  assign n34117 = ~n34115 & n34116;
  assign n34118 = n6194 & ~n34117;
  assign n34119 = ~n34112 & n34118;
  assign n34120 = pi947 & ~n34119;
  assign n34121 = ~n34111 & n34120;
  assign n34122 = n20306 & ~n34080;
  assign n34123 = ~n2608 & ~n34121;
  assign n34124 = ~n34122 & n34123;
  assign n34125 = n2608 & ~n34083;
  assign n34126 = ~pi223 & ~n34125;
  assign n34127 = ~n16126 & n34126;
  assign n34128 = ~n34124 & n34127;
  assign n34129 = ~pi299 & ~n34109;
  assign n34130 = ~n34128 & n34129;
  assign n34131 = ~pi947 & n20206;
  assign n34132 = pi947 & ~n34100;
  assign n34133 = ~n34081 & ~n34132;
  assign n34134 = ~n34131 & n34133;
  assign n34135 = pi299 & ~n34134;
  assign n34136 = ~n34130 & ~n34135;
  assign n34137 = pi215 & ~n34136;
  assign n34138 = n16063 & n34125;
  assign n34139 = ~n16149 & n34080;
  assign n34140 = ~pi947 & ~n34139;
  assign n34141 = pi642 & n16108;
  assign n34142 = ~n6164 & n16146;
  assign n34143 = ~n16152 & ~n34142;
  assign n34144 = n34141 & n34143;
  assign n34145 = pi642 & ~n16108;
  assign n34146 = ~n16146 & n34145;
  assign n34147 = pi947 & ~n34146;
  assign n34148 = ~n34144 & n34147;
  assign n34149 = ~n34140 & ~n34148;
  assign n34150 = ~n6194 & ~n34149;
  assign n34151 = n16063 & n34145;
  assign n34152 = ~n16109 & n34141;
  assign n34153 = ~n16169 & n34152;
  assign n34154 = ~n34151 & ~n34153;
  assign n34155 = pi947 & ~n34154;
  assign n34156 = n16165 & n34081;
  assign n34157 = n6194 & ~n34155;
  assign n34158 = ~n34156 & n34157;
  assign n34159 = ~n2608 & ~n34150;
  assign n34160 = ~n34158 & n34159;
  assign n34161 = ~pi223 & ~n34138;
  assign n34162 = ~n34160 & n34161;
  assign n34163 = pi947 & ~n16081;
  assign n34164 = ~n16089 & ~n34163;
  assign n34165 = ~n6194 & n34164;
  assign n34166 = n6194 & ~n16095;
  assign n34167 = n34080 & ~n34166;
  assign n34168 = ~pi947 & ~n34167;
  assign n34169 = ~n16107 & n34152;
  assign n34170 = pi947 & ~n34151;
  assign n34171 = ~n34169 & n34170;
  assign n34172 = ~n34165 & ~n34171;
  assign n34173 = ~n34168 & n34172;
  assign n34174 = pi223 & ~n34173;
  assign n34175 = ~n34162 & ~n34174;
  assign n34176 = ~pi299 & ~n34175;
  assign n34177 = n16199 & ~n34083;
  assign n34178 = ~n3302 & n34149;
  assign n34179 = pi299 & ~n34177;
  assign n34180 = ~n34178 & n34179;
  assign n34181 = ~pi215 & ~n34180;
  assign n34182 = ~n34176 & n34181;
  assign n34183 = ~n34137 & ~n34182;
  assign n34184 = pi39 & ~n34183;
  assign n34185 = ~pi38 & ~n34096;
  assign n34186 = ~n34184 & n34185;
  assign n34187 = n9830 & ~n34086;
  assign n34188 = ~n34186 & n34187;
  assign po372 = n34078 | n34188;
  assign n34190 = pi216 & ~n16228;
  assign n34191 = pi662 & pi907;
  assign n34192 = ~pi947 & n34191;
  assign n34193 = pi614 & pi947;
  assign n34194 = ~n34192 & ~n34193;
  assign n34195 = n16228 & ~n34194;
  assign n34196 = pi38 & ~n34190;
  assign n34197 = ~n34195 & n34196;
  assign n34198 = ~pi216 & ~n16051;
  assign n34199 = n16051 & n34194;
  assign n34200 = pi299 & ~n34198;
  assign n34201 = ~n34199 & n34200;
  assign n34202 = ~pi216 & ~n16055;
  assign n34203 = n16055 & n34194;
  assign n34204 = ~pi299 & ~n34202;
  assign n34205 = ~n34203 & n34204;
  assign n34206 = ~n34201 & ~n34205;
  assign n34207 = ~pi39 & ~n34206;
  assign n34208 = ~pi614 & ~n16079;
  assign n34209 = n6164 & n34208;
  assign n34210 = ~n31705 & ~n31706;
  assign n34211 = n16173 & ~n34210;
  assign n34212 = ~n34209 & ~n34211;
  assign n34213 = ~n6194 & ~n34212;
  assign n34214 = ~pi614 & n6194;
  assign n34215 = ~n16116 & n34214;
  assign n34216 = ~n16117 & n34215;
  assign n34217 = ~n34213 & ~n34216;
  assign n34218 = pi947 & ~n34217;
  assign n34219 = ~n20314 & ~n34218;
  assign n34220 = pi223 & ~n34192;
  assign n34221 = ~n34219 & n34220;
  assign n34222 = n16154 & n34194;
  assign n34223 = pi947 & ~n16180;
  assign n34224 = ~pi947 & ~n34191;
  assign n34225 = n16184 & n34224;
  assign n34226 = ~n34223 & ~n34225;
  assign n34227 = n6194 & ~n34226;
  assign n34228 = ~n2608 & ~n34222;
  assign n34229 = ~n34227 & n34228;
  assign n34230 = n2608 & ~n34194;
  assign n34231 = ~pi223 & ~n34230;
  assign n34232 = ~n16126 & n34231;
  assign n34233 = ~n34229 & n34232;
  assign n34234 = pi216 & ~n34221;
  assign n34235 = ~n34233 & n34234;
  assign n34236 = ~n34166 & n34191;
  assign n34237 = ~pi947 & ~n34236;
  assign n34238 = ~n16107 & n16171;
  assign n34239 = pi947 & ~n16168;
  assign n34240 = ~n34238 & n34239;
  assign n34241 = ~n34165 & ~n34240;
  assign n34242 = ~n34237 & n34241;
  assign n34243 = pi223 & ~n34242;
  assign n34244 = n16063 & n34230;
  assign n34245 = n34143 & n34193;
  assign n34246 = ~n16149 & n34192;
  assign n34247 = ~n34245 & ~n34246;
  assign n34248 = ~n6194 & n34247;
  assign n34249 = ~n16168 & ~n16172;
  assign n34250 = pi947 & ~n34249;
  assign n34251 = n16165 & n34192;
  assign n34252 = n6194 & ~n34250;
  assign n34253 = ~n34251 & n34252;
  assign n34254 = ~n2608 & ~n34248;
  assign n34255 = ~n34253 & n34254;
  assign n34256 = ~pi223 & ~n34244;
  assign n34257 = ~n34255 & n34256;
  assign n34258 = ~pi216 & ~n34243;
  assign n34259 = ~n34257 & n34258;
  assign n34260 = ~pi299 & ~n34259;
  assign n34261 = ~n34235 & n34260;
  assign n34262 = ~n34163 & ~n34192;
  assign n34263 = ~n34240 & ~n34262;
  assign n34264 = ~n34164 & n34263;
  assign n34265 = ~pi216 & ~n34264;
  assign n34266 = pi947 & n34212;
  assign n34267 = pi216 & ~n34192;
  assign n34268 = ~n34266 & n34267;
  assign n34269 = ~n34131 & n34268;
  assign n34270 = ~n34265 & ~n34269;
  assign n34271 = pi215 & ~n34270;
  assign n34272 = n5724 & ~n34247;
  assign n34273 = ~n16196 & n34194;
  assign n34274 = pi216 & ~n34273;
  assign n34275 = n16199 & ~n34194;
  assign n34276 = ~pi215 & ~n34275;
  assign n34277 = ~n34272 & n34276;
  assign n34278 = ~n34274 & n34277;
  assign n34279 = ~n34271 & ~n34278;
  assign n34280 = pi299 & ~n34279;
  assign n34281 = pi39 & ~n34261;
  assign n34282 = ~n34280 & n34281;
  assign n34283 = ~pi38 & ~n34207;
  assign n34284 = ~n34282 & n34283;
  assign n34285 = ~n34197 & ~n34284;
  assign n34286 = n9830 & ~n34285;
  assign n34287 = ~pi216 & ~n9830;
  assign po373 = ~n34286 & ~n34287;
  assign n34289 = pi695 & ~n33770;
  assign n34290 = ~pi695 & ~n33792;
  assign n34291 = ~pi217 & ~n34289;
  assign n34292 = ~n34290 & n34291;
  assign n34293 = pi695 & n33803;
  assign n34294 = ~pi695 & n33855;
  assign n34295 = pi217 & ~n34293;
  assign n34296 = ~n34294 & n34295;
  assign n34297 = pi612 & ~n34296;
  assign n34298 = ~n34292 & n34297;
  assign n34299 = ~pi695 & n33825;
  assign n34300 = pi217 & ~n34299;
  assign n34301 = pi695 & ~n33716;
  assign n34302 = ~pi695 & ~n33751;
  assign n34303 = ~pi217 & ~n34301;
  assign n34304 = ~n34302 & n34303;
  assign n34305 = ~pi612 & ~n34300;
  assign n34306 = ~n34304 & n34305;
  assign po374 = n34298 | n34306;
  assign n34308 = n33045 & ~n33115;
  assign n34309 = ~n33045 & ~n33145;
  assign n34310 = ~n34308 & ~n34309;
  assign n34311 = ~pi218 & ~n34310;
  assign n34312 = n33045 & n33153;
  assign n34313 = pi218 & ~n34312;
  assign po375 = ~n34311 & ~n34313;
  assign n34315 = ~pi219 & ~po1038;
  assign n34316 = pi617 & ~n34004;
  assign n34317 = ~pi617 & ~n34002;
  assign n34318 = pi637 & ~n34316;
  assign n34319 = ~n34317 & n34318;
  assign n34320 = pi617 & ~pi637;
  assign n34321 = n34008 & n34320;
  assign n34322 = ~n34319 & ~n34321;
  assign n34323 = n34315 & ~n34322;
  assign n34324 = ~pi617 & ~n33988;
  assign n34325 = pi617 & ~n33990;
  assign n34326 = pi637 & ~n34325;
  assign n34327 = ~n34324 & n34326;
  assign n34328 = ~pi617 & ~n16219;
  assign n34329 = pi617 & ~n33994;
  assign n34330 = ~pi637 & ~n34328;
  assign n34331 = ~n34329 & n34330;
  assign n34332 = ~n34327 & ~n34331;
  assign n34333 = ~po1038 & ~n34332;
  assign n34334 = pi219 & ~n34333;
  assign po376 = n34323 | n34334;
  assign n34336 = ~n32988 & n33164;
  assign n34337 = ~n33024 & ~n33164;
  assign n34338 = ~n34336 & ~n34337;
  assign n34339 = ~pi220 & ~n34338;
  assign n34340 = n33033 & n33164;
  assign n34341 = pi220 & ~n34340;
  assign po377 = ~n34339 & ~n34341;
  assign n34343 = pi221 & ~n16228;
  assign n34344 = pi661 & n19798;
  assign n34345 = pi616 & pi947;
  assign n34346 = ~n34344 & ~n34345;
  assign n34347 = n16228 & ~n34346;
  assign n34348 = pi38 & ~n34343;
  assign n34349 = ~n34347 & n34348;
  assign n34350 = ~pi221 & ~n16051;
  assign n34351 = n16051 & n34346;
  assign n34352 = pi299 & ~n34350;
  assign n34353 = ~n34351 & n34352;
  assign n34354 = ~pi221 & ~n16055;
  assign n34355 = n16055 & n34346;
  assign n34356 = ~pi299 & ~n34354;
  assign n34357 = ~n34355 & n34356;
  assign n34358 = ~n34353 & ~n34357;
  assign n34359 = ~pi39 & ~n34358;
  assign n34360 = n16063 & ~n34346;
  assign n34361 = ~pi216 & n34360;
  assign n34362 = n34143 & n34345;
  assign n34363 = ~n16149 & n34344;
  assign n34364 = ~n34362 & ~n34363;
  assign n34365 = pi216 & ~n34364;
  assign n34366 = ~pi221 & ~n34361;
  assign n34367 = ~n34365 & n34366;
  assign n34368 = ~pi947 & n19879;
  assign n34369 = pi221 & ~n34344;
  assign n34370 = ~pi616 & ~n16108;
  assign n34371 = ~n6166 & n16163;
  assign n34372 = ~n16145 & ~n34371;
  assign n34373 = n34370 & ~n34372;
  assign n34374 = ~pi616 & n16108;
  assign n34375 = ~n34110 & ~n34144;
  assign n34376 = n34374 & ~n34375;
  assign n34377 = ~n34373 & ~n34376;
  assign n34378 = pi947 & n34377;
  assign n34379 = n34369 & ~n34378;
  assign n34380 = ~n34368 & n34379;
  assign n34381 = ~pi215 & ~n34367;
  assign n34382 = ~n34380 & n34381;
  assign n34383 = pi947 & ~n16115;
  assign n34384 = ~n34344 & ~n34383;
  assign n34385 = ~n34164 & ~n34384;
  assign n34386 = ~pi221 & ~n34385;
  assign n34387 = ~pi616 & ~n34097;
  assign n34388 = ~n34098 & n34387;
  assign n34389 = pi947 & ~n34388;
  assign n34390 = n34369 & ~n34389;
  assign n34391 = ~n34131 & n34390;
  assign n34392 = pi215 & ~n34386;
  assign n34393 = ~n34391 & n34392;
  assign n34394 = pi299 & ~n34393;
  assign n34395 = ~n34382 & n34394;
  assign n34396 = ~pi947 & ~n16104;
  assign n34397 = ~n34389 & ~n34396;
  assign n34398 = ~n6194 & ~n34397;
  assign n34399 = pi947 & n16119;
  assign n34400 = ~pi947 & n16122;
  assign n34401 = n6194 & ~n34399;
  assign n34402 = ~n34400 & n34401;
  assign n34403 = pi223 & ~n34344;
  assign n34404 = ~n34402 & n34403;
  assign n34405 = ~n34398 & n34404;
  assign n34406 = n2608 & n34360;
  assign n34407 = ~pi223 & ~n34406;
  assign n34408 = ~n6194 & n34377;
  assign n34409 = n16163 & n34370;
  assign n34410 = ~n16181 & n34374;
  assign n34411 = n6194 & ~n34409;
  assign n34412 = ~n34410 & n34411;
  assign n34413 = pi947 & ~n34412;
  assign n34414 = ~n34408 & n34413;
  assign n34415 = ~n20306 & ~n34414;
  assign n34416 = ~n34344 & ~n34415;
  assign n34417 = ~n2608 & ~n34416;
  assign n34418 = ~n16126 & n34407;
  assign n34419 = ~n34417 & n34418;
  assign n34420 = pi221 & ~n34405;
  assign n34421 = ~n34419 & n34420;
  assign n34422 = ~n6194 & n34364;
  assign n34423 = n16165 & n34344;
  assign n34424 = n16111 & ~n16169;
  assign n34425 = ~n16114 & ~n34424;
  assign n34426 = pi947 & ~n34425;
  assign n34427 = n6194 & ~n34426;
  assign n34428 = ~n34423 & n34427;
  assign n34429 = ~n2608 & ~n34422;
  assign n34430 = ~n34428 & n34429;
  assign n34431 = n34407 & ~n34430;
  assign n34432 = n34166 & ~n34383;
  assign n34433 = ~n34165 & ~n34384;
  assign n34434 = ~n34432 & n34433;
  assign n34435 = pi223 & ~n34434;
  assign n34436 = ~pi221 & ~n34435;
  assign n34437 = ~n34431 & n34436;
  assign n34438 = ~pi299 & ~n34437;
  assign n34439 = ~n34421 & n34438;
  assign n34440 = pi39 & ~n34395;
  assign n34441 = ~n34439 & n34440;
  assign n34442 = ~pi38 & ~n34359;
  assign n34443 = ~n34441 & n34442;
  assign n34444 = ~n34349 & ~n34443;
  assign n34445 = n9830 & ~n34444;
  assign n34446 = ~pi221 & ~n9830;
  assign po378 = ~n34445 & ~n34446;
  assign n34448 = ~pi223 & n16186;
  assign n34449 = ~n16125 & ~n34448;
  assign n34450 = ~pi299 & ~n34449;
  assign n34451 = pi39 & ~n34450;
  assign n34452 = ~n16211 & n34451;
  assign n34453 = ~pi38 & ~n17347;
  assign n34454 = ~n34452 & n34453;
  assign n34455 = n17793 & ~n34454;
  assign n34456 = pi222 & ~n34455;
  assign n34457 = ~n28954 & ~n34456;
  assign n34458 = n15777 & ~n34456;
  assign n34459 = pi222 & ~n9829;
  assign n34460 = pi222 & ~n16228;
  assign n34461 = pi38 & ~n34460;
  assign n34462 = pi616 & n16570;
  assign n34463 = n34461 & ~n34462;
  assign n34464 = pi222 & n16447;
  assign n34465 = ~pi222 & ~n16526;
  assign n34466 = ~pi616 & n16526;
  assign n34467 = ~pi39 & ~n34465;
  assign n34468 = ~n34466 & n34467;
  assign n34469 = ~n34464 & n34468;
  assign n34470 = ~n16149 & ~n16767;
  assign n34471 = ~n6162 & ~n34470;
  assign n34472 = ~n16767 & n31936;
  assign n34473 = ~n16456 & ~n34472;
  assign n34474 = n6163 & ~n34473;
  assign n34475 = ~n6163 & n34470;
  assign n34476 = n6162 & ~n34474;
  assign n34477 = ~n34475 & n34476;
  assign n34478 = ~n34471 & ~n34477;
  assign n34479 = ~n6194 & n34478;
  assign n34480 = pi616 & ~n16449;
  assign n34481 = ~n16164 & ~n34480;
  assign n34482 = ~n6162 & ~n34481;
  assign n34483 = n6163 & ~n16767;
  assign n34484 = n16157 & n34483;
  assign n34485 = ~n6163 & n34481;
  assign n34486 = n6162 & ~n34484;
  assign n34487 = ~n34485 & n34486;
  assign n34488 = ~n34482 & ~n34487;
  assign n34489 = n6194 & n34488;
  assign n34490 = pi222 & ~n34479;
  assign n34491 = ~n34489 & n34490;
  assign n34492 = n15780 & n34143;
  assign n34493 = pi616 & n34492;
  assign n34494 = ~n6194 & n34493;
  assign n34495 = ~n6164 & ~n16528;
  assign n34496 = ~n16465 & ~n34495;
  assign n34497 = n6194 & n34496;
  assign n34498 = pi616 & n34497;
  assign n34499 = pi224 & ~n34494;
  assign n34500 = ~n34498 & n34499;
  assign n34501 = n15780 & n16113;
  assign n34502 = ~pi224 & ~n34501;
  assign n34503 = ~pi222 & ~n34502;
  assign n34504 = ~n34500 & n34503;
  assign n34505 = ~pi223 & ~n34504;
  assign n34506 = ~n34491 & n34505;
  assign n34507 = ~n6166 & n34097;
  assign n34508 = n34501 & ~n34507;
  assign n34509 = ~pi222 & n34508;
  assign n34510 = ~n16329 & n34509;
  assign n34511 = pi616 & ~n16486;
  assign n34512 = n16089 & ~n34511;
  assign n34513 = ~n6162 & ~n34512;
  assign n34514 = ~n6163 & ~n16089;
  assign n34515 = ~n16097 & ~n34511;
  assign n34516 = ~n34514 & n34515;
  assign n34517 = n6162 & ~n34516;
  assign n34518 = ~n34513 & ~n34517;
  assign n34519 = ~n6194 & n34518;
  assign n34520 = ~pi616 & ~n16095;
  assign n34521 = ~n34480 & ~n34520;
  assign n34522 = ~n6162 & ~n34521;
  assign n34523 = n16085 & n34483;
  assign n34524 = ~n6163 & n34521;
  assign n34525 = n6162 & ~n34523;
  assign n34526 = ~n34524 & n34525;
  assign n34527 = ~n34522 & ~n34526;
  assign n34528 = n6194 & n34527;
  assign n34529 = pi222 & ~n34519;
  assign n34530 = ~n34528 & n34529;
  assign n34531 = pi223 & ~n34510;
  assign n34532 = ~n34530 & n34531;
  assign n34533 = ~n34506 & ~n34532;
  assign n34534 = ~pi299 & ~n34533;
  assign n34535 = ~n16293 & n34509;
  assign n34536 = n6221 & n34527;
  assign n34537 = ~n6221 & n34518;
  assign n34538 = pi222 & ~n34537;
  assign n34539 = ~n34536 & n34538;
  assign n34540 = ~n34535 & ~n34539;
  assign n34541 = pi215 & ~n34540;
  assign n34542 = pi222 & ~n16063;
  assign n34543 = n3302 & ~n34542;
  assign n34544 = ~n34501 & n34543;
  assign n34545 = ~n6221 & n34478;
  assign n34546 = n6221 & n34488;
  assign n34547 = pi222 & ~n34545;
  assign n34548 = ~n34546 & n34547;
  assign n34549 = pi616 & n34496;
  assign n34550 = n6221 & ~n34549;
  assign n34551 = ~n6221 & ~n34493;
  assign n34552 = ~pi222 & ~n34550;
  assign n34553 = ~n34551 & n34552;
  assign n34554 = ~n3302 & ~n34553;
  assign n34555 = ~n34548 & n34554;
  assign n34556 = ~pi215 & ~n34544;
  assign n34557 = ~n34555 & n34556;
  assign n34558 = pi299 & ~n34541;
  assign n34559 = ~n34557 & n34558;
  assign n34560 = pi39 & ~n34534;
  assign n34561 = ~n34559 & n34560;
  assign n34562 = ~pi38 & ~n34469;
  assign n34563 = ~n34561 & n34562;
  assign n34564 = n9829 & ~n34463;
  assign n34565 = ~n34563 & n34564;
  assign n34566 = ~n34459 & ~n34565;
  assign n34567 = ~n15777 & n34566;
  assign n34568 = ~n34458 & ~n34567;
  assign n34569 = ~pi785 & n34568;
  assign n34570 = ~pi609 & ~n34456;
  assign n34571 = pi609 & ~n34568;
  assign n34572 = pi1155 & ~n34570;
  assign n34573 = ~n34571 & n34572;
  assign n34574 = pi609 & ~n34456;
  assign n34575 = ~pi609 & ~n34568;
  assign n34576 = ~pi1155 & ~n34574;
  assign n34577 = ~n34575 & n34576;
  assign n34578 = ~n34573 & ~n34577;
  assign n34579 = pi785 & ~n34578;
  assign n34580 = ~n34569 & ~n34579;
  assign n34581 = ~pi781 & ~n34580;
  assign n34582 = pi618 & n34580;
  assign n34583 = ~pi618 & ~n34456;
  assign n34584 = pi1154 & ~n34583;
  assign n34585 = ~n34582 & n34584;
  assign n34586 = ~pi618 & n34580;
  assign n34587 = pi618 & ~n34456;
  assign n34588 = ~pi1154 & ~n34587;
  assign n34589 = ~n34586 & n34588;
  assign n34590 = ~n34585 & ~n34589;
  assign n34591 = pi781 & ~n34590;
  assign n34592 = ~n34581 & ~n34591;
  assign n34593 = ~pi789 & ~n34592;
  assign n34594 = pi619 & n34592;
  assign n34595 = ~pi619 & ~n34456;
  assign n34596 = pi1159 & ~n34595;
  assign n34597 = ~n34594 & n34596;
  assign n34598 = ~pi619 & n34592;
  assign n34599 = pi619 & ~n34456;
  assign n34600 = ~pi1159 & ~n34599;
  assign n34601 = ~n34598 & n34600;
  assign n34602 = ~n34597 & ~n34601;
  assign n34603 = pi789 & ~n34602;
  assign n34604 = ~n34593 & ~n34603;
  assign n34605 = ~n15832 & n34604;
  assign n34606 = n19771 & n34605;
  assign n34607 = ~n34457 & ~n34606;
  assign n34608 = ~pi644 & ~n34607;
  assign n34609 = pi644 & ~n34456;
  assign n34610 = pi715 & ~n34609;
  assign n34611 = ~n34608 & n34610;
  assign n34612 = n15765 & ~n34456;
  assign n34613 = ~n17585 & ~n34456;
  assign n34614 = n15741 & ~n34456;
  assign n34615 = pi661 & n16226;
  assign n34616 = n34461 & ~n34615;
  assign n34617 = pi661 & pi680;
  assign n34618 = n16345 & ~n34617;
  assign n34619 = ~pi222 & ~n16345;
  assign n34620 = pi222 & n16359;
  assign n34621 = ~pi299 & ~n34620;
  assign n34622 = ~n34618 & n34621;
  assign n34623 = ~n34619 & n34622;
  assign n34624 = pi222 & n16364;
  assign n34625 = n16350 & ~n34617;
  assign n34626 = ~pi222 & ~n16350;
  assign n34627 = pi299 & ~n34624;
  assign n34628 = ~n34625 & n34627;
  assign n34629 = ~n34626 & n34628;
  assign n34630 = ~pi39 & ~n34623;
  assign n34631 = ~n34629 & n34630;
  assign n34632 = ~pi661 & ~n16153;
  assign n34633 = ~n15725 & ~n16149;
  assign n34634 = pi661 & ~n34633;
  assign n34635 = ~n34632 & ~n34634;
  assign n34636 = ~n6194 & n34635;
  assign n34637 = pi661 & ~n16246;
  assign n34638 = ~pi661 & ~n16184;
  assign n34639 = ~n34637 & ~n34638;
  assign n34640 = n6194 & n34639;
  assign n34641 = pi222 & ~n34636;
  assign n34642 = ~n34640 & n34641;
  assign n34643 = pi661 & n16298;
  assign n34644 = ~pi224 & ~n34643;
  assign n34645 = ~n16308 & n34617;
  assign n34646 = n6194 & n34645;
  assign n34647 = n15725 & ~n16149;
  assign n34648 = pi661 & n34647;
  assign n34649 = ~n6194 & n34648;
  assign n34650 = pi224 & ~n34646;
  assign n34651 = ~n34649 & n34650;
  assign n34652 = ~pi222 & ~n34644;
  assign n34653 = ~n34651 & n34652;
  assign n34654 = ~pi223 & ~n34653;
  assign n34655 = ~n34642 & n34654;
  assign n34656 = ~pi222 & pi661;
  assign n34657 = n16330 & n34656;
  assign n34658 = ~pi661 & n16090;
  assign n34659 = n6162 & n16100;
  assign n34660 = pi661 & ~n16271;
  assign n34661 = ~n34658 & ~n34660;
  assign n34662 = ~n34659 & n34661;
  assign n34663 = ~n6194 & n34662;
  assign n34664 = ~pi661 & ~n16122;
  assign n34665 = ~n16257 & ~n16262;
  assign n34666 = pi661 & ~n34665;
  assign n34667 = ~n34664 & ~n34666;
  assign n34668 = n6194 & n34667;
  assign n34669 = pi222 & ~n34663;
  assign n34670 = ~n34668 & n34669;
  assign n34671 = pi223 & ~n34657;
  assign n34672 = ~n34670 & n34671;
  assign n34673 = ~n34655 & ~n34672;
  assign n34674 = ~pi299 & ~n34673;
  assign n34675 = ~n16293 & n16299;
  assign n34676 = n34656 & n34675;
  assign n34677 = ~n6221 & n34662;
  assign n34678 = n6221 & n34667;
  assign n34679 = pi222 & ~n34677;
  assign n34680 = ~n34678 & n34679;
  assign n34681 = ~n34676 & ~n34680;
  assign n34682 = pi215 & ~n34681;
  assign n34683 = ~n6221 & n34635;
  assign n34684 = n6221 & n34639;
  assign n34685 = pi222 & ~n34683;
  assign n34686 = ~n34684 & n34685;
  assign n34687 = ~n6221 & ~n34648;
  assign n34688 = n6221 & ~n34645;
  assign n34689 = ~pi222 & ~n34687;
  assign n34690 = ~n34688 & n34689;
  assign n34691 = ~n3302 & ~n34690;
  assign n34692 = ~n34686 & n34691;
  assign n34693 = n34543 & ~n34643;
  assign n34694 = ~pi215 & ~n34693;
  assign n34695 = ~n34692 & n34694;
  assign n34696 = pi299 & ~n34682;
  assign n34697 = ~n34695 & n34696;
  assign n34698 = ~n34674 & ~n34697;
  assign n34699 = pi39 & ~n34698;
  assign n34700 = ~n34631 & ~n34699;
  assign n34701 = ~pi38 & ~n34700;
  assign n34702 = n9829 & ~n34616;
  assign n34703 = ~n34701 & n34702;
  assign n34704 = ~n34459 & ~n34703;
  assign n34705 = ~pi778 & ~n34704;
  assign n34706 = pi625 & n34704;
  assign n34707 = ~pi625 & ~n34456;
  assign n34708 = pi1153 & ~n34707;
  assign n34709 = ~n34706 & n34708;
  assign n34710 = ~pi625 & n34704;
  assign n34711 = pi625 & ~n34456;
  assign n34712 = ~pi1153 & ~n34711;
  assign n34713 = ~n34710 & n34712;
  assign n34714 = ~n34709 & ~n34713;
  assign n34715 = pi778 & ~n34714;
  assign n34716 = ~n34705 & ~n34715;
  assign n34717 = ~n15741 & n34716;
  assign n34718 = ~n34614 & ~n34717;
  assign n34719 = ~n15747 & ~n34718;
  assign n34720 = n15747 & ~n34456;
  assign n34721 = ~n34719 & ~n34720;
  assign n34722 = ~n15753 & ~n34721;
  assign n34723 = ~n15759 & n34722;
  assign n34724 = ~n34613 & ~n34723;
  assign n34725 = ~n15765 & ~n34724;
  assign n34726 = ~n34612 & ~n34725;
  assign n34727 = ~pi787 & n34726;
  assign n34728 = n19394 & n34726;
  assign n34729 = ~n19394 & n34456;
  assign n34730 = ~n34728 & ~n34729;
  assign n34731 = pi787 & ~n34730;
  assign n34732 = ~n34727 & ~n34731;
  assign n34733 = pi644 & n34732;
  assign n34734 = n15832 & ~n34456;
  assign n34735 = ~n34605 & ~n34734;
  assign n34736 = ~n15925 & ~n34735;
  assign n34737 = n15925 & ~n34456;
  assign n34738 = n19478 & ~n34737;
  assign n34739 = ~n34736 & n34738;
  assign n34740 = ~n15959 & ~n34612;
  assign n34741 = ~n34730 & n34740;
  assign n34742 = ~n34739 & ~n34741;
  assign n34743 = pi787 & ~n34742;
  assign n34744 = pi628 & ~n34456;
  assign n34745 = ~pi628 & ~n34724;
  assign n34746 = n15923 & ~n34744;
  assign n34747 = ~n34745 & n34746;
  assign n34748 = ~n16633 & n34735;
  assign n34749 = ~pi628 & ~n34456;
  assign n34750 = pi628 & ~n34724;
  assign n34751 = n15922 & ~n34749;
  assign n34752 = ~n34750 & n34751;
  assign n34753 = ~n34747 & ~n34752;
  assign n34754 = ~n34748 & n34753;
  assign n34755 = pi792 & ~n34754;
  assign n34756 = pi626 & n34604;
  assign n34757 = ~pi626 & ~n34456;
  assign n34758 = n15756 & ~n34757;
  assign n34759 = ~n34756 & n34758;
  assign n34760 = n15753 & ~n34456;
  assign n34761 = n15828 & ~n34760;
  assign n34762 = ~n34722 & n34761;
  assign n34763 = ~pi626 & n34604;
  assign n34764 = pi626 & ~n34456;
  assign n34765 = n15757 & ~n34764;
  assign n34766 = ~n34763 & n34765;
  assign n34767 = ~n34759 & ~n34762;
  assign n34768 = ~n34766 & n34767;
  assign n34769 = ~n15833 & n34768;
  assign n34770 = pi618 & ~n34718;
  assign n34771 = pi609 & n34716;
  assign n34772 = n16065 & n16679;
  assign n34773 = ~pi222 & ~pi616;
  assign n34774 = ~pi39 & pi616;
  assign n34775 = n34617 & n34774;
  assign n34776 = ~n34773 & ~n34775;
  assign n34777 = n34772 & ~n34776;
  assign n34778 = ~n16767 & ~n34617;
  assign n34779 = ~pi616 & ~n16664;
  assign n34780 = ~n34778 & ~n34779;
  assign n34781 = n16228 & n34780;
  assign n34782 = ~n34460 & ~n34781;
  assign n34783 = ~n34777 & ~n34782;
  assign n34784 = pi38 & ~n34783;
  assign n34785 = pi616 & ~n16716;
  assign n34786 = ~n16724 & ~n34785;
  assign n34787 = n34617 & ~n34786;
  assign n34788 = n34522 & ~n34617;
  assign n34789 = ~n34526 & ~n34787;
  assign n34790 = ~n34788 & n34789;
  assign n34791 = n6194 & ~n34790;
  assign n34792 = ~pi661 & pi681;
  assign n34793 = ~n34512 & n34792;
  assign n34794 = ~pi680 & n34512;
  assign n34795 = pi680 & ~n16708;
  assign n34796 = ~n16705 & ~n16767;
  assign n34797 = n34795 & n34796;
  assign n34798 = pi661 & ~n34797;
  assign n34799 = ~n34794 & n34798;
  assign n34800 = ~n34517 & ~n34793;
  assign n34801 = ~n34799 & n34800;
  assign n34802 = ~n6194 & ~n34801;
  assign n34803 = pi222 & ~n34802;
  assign n34804 = ~n34791 & n34803;
  assign n34805 = n16786 & n34617;
  assign n34806 = ~n34508 & ~n34805;
  assign n34807 = n6194 & ~n34806;
  assign n34808 = ~n16081 & n34501;
  assign n34809 = ~pi661 & ~n34808;
  assign n34810 = pi616 & n16701;
  assign n34811 = n6164 & ~n34810;
  assign n34812 = ~pi680 & n34808;
  assign n34813 = ~n16530 & ~n17835;
  assign n34814 = pi616 & n34813;
  assign n34815 = pi614 & ~pi616;
  assign n34816 = ~n16792 & n34815;
  assign n34817 = pi680 & ~n34814;
  assign n34818 = ~n34816 & n34817;
  assign n34819 = ~n16796 & n34818;
  assign n34820 = pi661 & ~n34812;
  assign n34821 = ~n34819 & n34820;
  assign n34822 = ~n34809 & ~n34811;
  assign n34823 = ~n34821 & n34822;
  assign n34824 = ~n6194 & n34823;
  assign n34825 = ~pi222 & ~n34807;
  assign n34826 = ~n34824 & n34825;
  assign n34827 = pi223 & ~n34826;
  assign n34828 = ~n34804 & n34827;
  assign n34829 = n6166 & n16239;
  assign n34830 = ~n16268 & ~n34829;
  assign n34831 = n15780 & ~n16146;
  assign n34832 = n34830 & ~n34831;
  assign n34833 = n34815 & n34832;
  assign n34834 = n16679 & ~n34830;
  assign n34835 = pi616 & ~n34834;
  assign n34836 = ~pi603 & ~n34830;
  assign n34837 = pi603 & ~n16663;
  assign n34838 = ~n16144 & n34837;
  assign n34839 = ~n34836 & ~n34838;
  assign n34840 = ~pi642 & ~n34839;
  assign n34841 = pi642 & ~n34832;
  assign n34842 = n6160 & ~n34840;
  assign n34843 = ~n34841 & n34842;
  assign n34844 = ~n34833 & ~n34835;
  assign n34845 = ~n34843 & n34844;
  assign n34846 = pi680 & ~n34845;
  assign n34847 = pi661 & n34846;
  assign n34848 = n34471 & ~n34617;
  assign n34849 = ~n34477 & ~n34848;
  assign n34850 = ~n34847 & n34849;
  assign n34851 = ~n6194 & n34850;
  assign n34852 = ~n34481 & n34792;
  assign n34853 = ~pi680 & n34481;
  assign n34854 = pi680 & ~n34785;
  assign n34855 = ~n16691 & n34854;
  assign n34856 = pi661 & ~n34853;
  assign n34857 = ~n34855 & n34856;
  assign n34858 = ~n34487 & ~n34852;
  assign n34859 = ~n34857 & n34858;
  assign n34860 = n6194 & n34859;
  assign n34861 = pi222 & ~n34851;
  assign n34862 = ~n34860 & n34861;
  assign n34863 = n34501 & ~n34617;
  assign n34864 = ~pi616 & ~n16750;
  assign n34865 = pi616 & ~n16885;
  assign n34866 = ~n34778 & ~n34865;
  assign n34867 = ~n34864 & n34866;
  assign n34868 = ~pi224 & ~n34863;
  assign n34869 = ~n34867 & n34868;
  assign n34870 = pi616 & n6163;
  assign n34871 = n16464 & n34870;
  assign n34872 = ~pi681 & n34871;
  assign n34873 = ~pi661 & ~n34872;
  assign n34874 = ~n16146 & n16767;
  assign n34875 = n34873 & ~n34874;
  assign n34876 = ~pi680 & n34874;
  assign n34877 = pi680 & n16774;
  assign n34878 = pi661 & ~n34876;
  assign n34879 = ~n34877 & n34878;
  assign n34880 = ~n16152 & ~n34875;
  assign n34881 = ~n34879 & n34880;
  assign n34882 = ~n6194 & n34881;
  assign n34883 = ~n34501 & n34873;
  assign n34884 = n6164 & ~n34871;
  assign n34885 = pi680 & ~n16759;
  assign n34886 = ~n34865 & n34885;
  assign n34887 = pi661 & ~n34863;
  assign n34888 = ~n34886 & n34887;
  assign n34889 = ~n34883 & ~n34884;
  assign n34890 = ~n34888 & n34889;
  assign n34891 = n6194 & n34890;
  assign n34892 = pi224 & ~n34882;
  assign n34893 = ~n34891 & n34892;
  assign n34894 = ~pi222 & ~n34869;
  assign n34895 = ~n34893 & n34894;
  assign n34896 = ~n34862 & ~n34895;
  assign n34897 = ~pi223 & ~n34896;
  assign n34898 = ~pi299 & ~n34828;
  assign n34899 = ~n34897 & n34898;
  assign n34900 = n6221 & ~n34790;
  assign n34901 = ~n6221 & ~n34801;
  assign n34902 = pi222 & ~n34901;
  assign n34903 = ~n34900 & n34902;
  assign n34904 = n6221 & ~n34806;
  assign n34905 = ~n6221 & n34823;
  assign n34906 = ~pi222 & ~n34904;
  assign n34907 = ~n34905 & n34906;
  assign n34908 = pi215 & ~n34907;
  assign n34909 = ~n34903 & n34908;
  assign n34910 = n34543 & ~n34867;
  assign n34911 = ~pi222 & n34890;
  assign n34912 = pi222 & ~n34859;
  assign n34913 = n6221 & ~n34911;
  assign n34914 = ~n34912 & n34913;
  assign n34915 = ~pi222 & n34881;
  assign n34916 = pi222 & ~n34850;
  assign n34917 = ~n6221 & ~n34915;
  assign n34918 = ~n34916 & n34917;
  assign n34919 = ~n34914 & ~n34918;
  assign n34920 = ~n3302 & ~n34919;
  assign n34921 = ~pi215 & ~n34910;
  assign n34922 = ~n34920 & n34921;
  assign n34923 = pi299 & ~n34909;
  assign n34924 = ~n34922 & n34923;
  assign n34925 = ~n34899 & ~n34924;
  assign n34926 = pi39 & ~n34925;
  assign n34927 = pi616 & n16519;
  assign n34928 = pi661 & n18060;
  assign n34929 = ~n34927 & ~n34928;
  assign n34930 = ~pi222 & ~n34929;
  assign n34931 = n16359 & ~n16667;
  assign n34932 = n18059 & ~n34617;
  assign n34933 = ~pi616 & n16519;
  assign n34934 = pi222 & ~n34931;
  assign n34935 = ~n34933 & n34934;
  assign n34936 = ~n34932 & n34935;
  assign n34937 = ~n34930 & ~n34936;
  assign n34938 = ~pi299 & ~n34937;
  assign n34939 = pi616 & n16524;
  assign n34940 = n16350 & n18051;
  assign n34941 = n34617 & n34940;
  assign n34942 = ~n34939 & ~n34941;
  assign n34943 = ~pi222 & ~n34942;
  assign n34944 = n16364 & ~n16432;
  assign n34945 = ~pi616 & n16524;
  assign n34946 = ~n34617 & n34940;
  assign n34947 = pi222 & ~n34944;
  assign n34948 = ~n34945 & n34947;
  assign n34949 = ~n34946 & n34948;
  assign n34950 = ~n34943 & ~n34949;
  assign n34951 = pi299 & ~n34950;
  assign n34952 = ~pi39 & ~n34951;
  assign n34953 = ~n34938 & n34952;
  assign n34954 = ~n34926 & ~n34953;
  assign n34955 = ~pi38 & ~n34954;
  assign n34956 = n9829 & ~n34784;
  assign n34957 = ~n34955 & n34956;
  assign n34958 = ~n34459 & ~n34957;
  assign n34959 = ~pi625 & n34958;
  assign n34960 = pi625 & n34566;
  assign n34961 = ~pi1153 & ~n34960;
  assign n34962 = ~n34959 & n34961;
  assign n34963 = ~pi608 & ~n34709;
  assign n34964 = ~n34962 & n34963;
  assign n34965 = ~pi625 & n34566;
  assign n34966 = pi625 & n34958;
  assign n34967 = pi1153 & ~n34965;
  assign n34968 = ~n34966 & n34967;
  assign n34969 = pi608 & ~n34713;
  assign n34970 = ~n34968 & n34969;
  assign n34971 = ~n34964 & ~n34970;
  assign n34972 = pi778 & ~n34971;
  assign n34973 = ~pi778 & n34958;
  assign n34974 = ~n34972 & ~n34973;
  assign n34975 = ~pi609 & ~n34974;
  assign n34976 = ~pi1155 & ~n34771;
  assign n34977 = ~n34975 & n34976;
  assign n34978 = ~pi660 & ~n34573;
  assign n34979 = ~n34977 & n34978;
  assign n34980 = ~pi609 & n34716;
  assign n34981 = pi609 & ~n34974;
  assign n34982 = pi1155 & ~n34980;
  assign n34983 = ~n34981 & n34982;
  assign n34984 = pi660 & ~n34577;
  assign n34985 = ~n34983 & n34984;
  assign n34986 = ~n34979 & ~n34985;
  assign n34987 = pi785 & ~n34986;
  assign n34988 = ~pi785 & ~n34974;
  assign n34989 = ~n34987 & ~n34988;
  assign n34990 = ~pi618 & ~n34989;
  assign n34991 = ~pi1154 & ~n34770;
  assign n34992 = ~n34990 & n34991;
  assign n34993 = ~pi627 & ~n34585;
  assign n34994 = ~n34992 & n34993;
  assign n34995 = ~pi618 & ~n34718;
  assign n34996 = pi618 & ~n34989;
  assign n34997 = pi1154 & ~n34995;
  assign n34998 = ~n34996 & n34997;
  assign n34999 = pi627 & ~n34589;
  assign n35000 = ~n34998 & n34999;
  assign n35001 = ~n34994 & ~n35000;
  assign n35002 = pi781 & ~n35001;
  assign n35003 = ~pi781 & ~n34989;
  assign n35004 = ~n35002 & ~n35003;
  assign n35005 = ~pi789 & n35004;
  assign n35006 = pi788 & ~n34768;
  assign n35007 = ~pi619 & ~n34721;
  assign n35008 = pi619 & ~n35004;
  assign n35009 = pi1159 & ~n35007;
  assign n35010 = ~n35008 & n35009;
  assign n35011 = pi648 & ~n34601;
  assign n35012 = ~n35010 & n35011;
  assign n35013 = pi619 & ~n34721;
  assign n35014 = ~pi619 & ~n35004;
  assign n35015 = ~pi1159 & ~n35013;
  assign n35016 = ~n35014 & n35015;
  assign n35017 = ~pi648 & ~n34597;
  assign n35018 = ~n35016 & n35017;
  assign n35019 = pi789 & ~n35012;
  assign n35020 = ~n35018 & n35019;
  assign n35021 = ~n35005 & ~n35006;
  assign n35022 = ~n35020 & n35021;
  assign n35023 = ~n16644 & ~n34769;
  assign n35024 = ~n35022 & n35023;
  assign n35025 = ~n34755 & ~n35024;
  assign n35026 = n18841 & ~n35025;
  assign n35027 = ~n34743 & ~n35026;
  assign n35028 = ~pi644 & n35027;
  assign n35029 = ~pi715 & ~n34733;
  assign n35030 = ~n35028 & n35029;
  assign n35031 = ~pi1160 & ~n34611;
  assign n35032 = ~n35030 & n35031;
  assign n35033 = ~pi644 & n34732;
  assign n35034 = pi644 & n35027;
  assign n35035 = pi715 & ~n35033;
  assign n35036 = ~n35034 & n35035;
  assign n35037 = pi644 & ~n34607;
  assign n35038 = ~pi644 & ~n34456;
  assign n35039 = ~pi715 & ~n35038;
  assign n35040 = ~n35037 & n35039;
  assign n35041 = pi1160 & ~n35040;
  assign n35042 = ~n35036 & n35041;
  assign n35043 = ~n35032 & ~n35042;
  assign n35044 = pi790 & ~n35043;
  assign n35045 = ~pi790 & n35027;
  assign n35046 = ~n35044 & ~n35045;
  assign n35047 = ~po1038 & ~n35046;
  assign n35048 = ~pi222 & po1038;
  assign po379 = ~n35047 & ~n35048;
  assign n35050 = ~pi299 & n16124;
  assign n35051 = pi39 & ~n35050;
  assign n35052 = ~n16211 & n35051;
  assign n35053 = n2576 & ~n17347;
  assign n35054 = ~n35052 & n35053;
  assign n35055 = n17793 & ~n35054;
  assign n35056 = pi223 & ~n35055;
  assign n35057 = ~n28954 & ~n35056;
  assign n35058 = pi223 & ~n9829;
  assign n35059 = pi39 & pi223;
  assign n35060 = pi38 & ~n35059;
  assign n35061 = pi642 & n15780;
  assign n35062 = n16065 & ~n35061;
  assign n35063 = ~pi223 & ~n16065;
  assign n35064 = ~pi39 & ~n35063;
  assign n35065 = ~n35062 & n35064;
  assign n35066 = n35060 & ~n35065;
  assign n35067 = ~pi223 & pi642;
  assign n35068 = n16524 & n35067;
  assign n35069 = pi299 & ~n35068;
  assign n35070 = n6159 & n16523;
  assign n35071 = pi223 & ~n35070;
  assign n35072 = ~n16433 & n35071;
  assign n35073 = n35069 & ~n35072;
  assign n35074 = n16519 & n35067;
  assign n35075 = ~pi299 & ~n35074;
  assign n35076 = ~pi642 & n16519;
  assign n35077 = pi223 & ~n35076;
  assign n35078 = n16445 & n35077;
  assign n35079 = n35075 & ~n35078;
  assign n35080 = ~pi39 & ~n35073;
  assign n35081 = ~n35079 & n35080;
  assign n35082 = ~n6194 & n34492;
  assign n35083 = ~n34497 & ~n35082;
  assign n35084 = ~n2608 & ~n35083;
  assign n35085 = ~n16537 & ~n35084;
  assign n35086 = pi642 & ~n35085;
  assign n35087 = ~pi223 & ~n35086;
  assign n35088 = ~pi661 & n6163;
  assign n35089 = pi642 & ~n16486;
  assign n35090 = ~n16087 & n16452;
  assign n35091 = ~n16081 & ~n35089;
  assign n35092 = ~n35090 & n35091;
  assign n35093 = ~n35088 & n35092;
  assign n35094 = n35088 & ~n35089;
  assign n35095 = ~n16079 & n35094;
  assign n35096 = ~pi681 & ~n35095;
  assign n35097 = ~n35093 & n35096;
  assign n35098 = pi681 & ~n35092;
  assign n35099 = ~n35097 & ~n35098;
  assign n35100 = ~n6194 & ~n35099;
  assign n35101 = pi642 & n16528;
  assign n35102 = n16095 & ~n35101;
  assign n35103 = pi681 & ~n35102;
  assign n35104 = ~n35061 & n35088;
  assign n35105 = n16085 & n35104;
  assign n35106 = ~n35088 & n35102;
  assign n35107 = ~pi681 & ~n35105;
  assign n35108 = ~n35106 & n35107;
  assign n35109 = ~n35103 & ~n35108;
  assign n35110 = n6194 & ~n35109;
  assign n35111 = pi223 & ~n35100;
  assign n35112 = ~n35110 & n35111;
  assign n35113 = ~n35087 & ~n35112;
  assign n35114 = ~pi299 & ~n35113;
  assign n35115 = n6221 & ~n35109;
  assign n35116 = ~n6221 & ~n35099;
  assign n35117 = pi223 & ~n35116;
  assign n35118 = ~n35115 & n35117;
  assign n35119 = ~n35088 & n35101;
  assign n35120 = ~pi681 & ~n35119;
  assign n35121 = pi642 & n35088;
  assign n35122 = n16529 & n35121;
  assign n35123 = n35120 & ~n35122;
  assign n35124 = n16081 & n35096;
  assign n35125 = ~n35123 & ~n35124;
  assign n35126 = pi642 & n16530;
  assign n35127 = pi681 & ~n35126;
  assign n35128 = ~n6221 & n35125;
  assign n35129 = ~n35127 & n35128;
  assign n35130 = n6221 & ~n35123;
  assign n35131 = ~pi947 & n35101;
  assign n35132 = n35130 & n35131;
  assign n35133 = ~pi223 & ~n35132;
  assign n35134 = ~n35129 & n35133;
  assign n35135 = pi215 & ~n35134;
  assign n35136 = ~n35118 & n35135;
  assign n35137 = pi223 & ~n16063;
  assign n35138 = n3302 & ~n35137;
  assign n35139 = ~n35101 & n35138;
  assign n35140 = n34113 & ~n35061;
  assign n35141 = pi642 & ~n16449;
  assign n35142 = n6160 & ~n35141;
  assign n35143 = ~n16160 & n35142;
  assign n35144 = ~n35140 & ~n35143;
  assign n35145 = pi681 & n35144;
  assign n35146 = ~n35088 & ~n35144;
  assign n35147 = n16157 & n35104;
  assign n35148 = ~pi681 & ~n35147;
  assign n35149 = ~n35146 & n35148;
  assign n35150 = n6221 & ~n35149;
  assign n35151 = ~n35145 & n35150;
  assign n35152 = ~pi642 & ~n16149;
  assign n35153 = pi642 & ~n15780;
  assign n35154 = ~n16146 & n35153;
  assign n35155 = ~n35152 & ~n35154;
  assign n35156 = pi681 & n35155;
  assign n35157 = ~n35088 & ~n35155;
  assign n35158 = ~n16144 & n35104;
  assign n35159 = ~pi681 & ~n35158;
  assign n35160 = ~n35157 & n35159;
  assign n35161 = ~n6221 & ~n35160;
  assign n35162 = ~n35156 & n35161;
  assign n35163 = ~n35151 & ~n35162;
  assign n35164 = pi223 & ~n35163;
  assign n35165 = pi642 & n34492;
  assign n35166 = ~n6221 & n35165;
  assign n35167 = pi642 & n6221;
  assign n35168 = n34496 & n35167;
  assign n35169 = ~pi223 & ~n35168;
  assign n35170 = ~n35166 & n35169;
  assign n35171 = ~n35164 & ~n35170;
  assign n35172 = ~n3302 & ~n35171;
  assign n35173 = ~pi215 & ~n35139;
  assign n35174 = ~n35172 & n35173;
  assign n35175 = pi299 & ~n35136;
  assign n35176 = ~n35174 & n35175;
  assign n35177 = pi39 & ~n35114;
  assign n35178 = ~n35176 & n35177;
  assign n35179 = ~pi38 & ~n35081;
  assign n35180 = ~n35178 & n35179;
  assign n35181 = n9829 & ~n35066;
  assign n35182 = ~n35180 & n35181;
  assign n35183 = ~n35058 & ~n35182;
  assign n35184 = ~n15777 & ~n35183;
  assign n35185 = n15777 & n35056;
  assign n35186 = ~n35184 & ~n35185;
  assign n35187 = ~pi785 & ~n35186;
  assign n35188 = pi609 & n35186;
  assign n35189 = ~pi609 & ~n35056;
  assign n35190 = pi1155 & ~n35189;
  assign n35191 = ~n35188 & n35190;
  assign n35192 = ~pi609 & n35186;
  assign n35193 = pi609 & ~n35056;
  assign n35194 = ~pi1155 & ~n35193;
  assign n35195 = ~n35192 & n35194;
  assign n35196 = ~n35191 & ~n35195;
  assign n35197 = pi785 & ~n35196;
  assign n35198 = ~n35187 & ~n35197;
  assign n35199 = ~pi781 & ~n35198;
  assign n35200 = pi618 & n35198;
  assign n35201 = ~pi618 & ~n35056;
  assign n35202 = pi1154 & ~n35201;
  assign n35203 = ~n35200 & n35202;
  assign n35204 = ~pi618 & n35198;
  assign n35205 = pi618 & ~n35056;
  assign n35206 = ~pi1154 & ~n35205;
  assign n35207 = ~n35204 & n35206;
  assign n35208 = ~n35203 & ~n35207;
  assign n35209 = pi781 & ~n35208;
  assign n35210 = ~n35199 & ~n35209;
  assign n35211 = ~pi789 & ~n35210;
  assign n35212 = pi619 & n35210;
  assign n35213 = ~pi619 & ~n35056;
  assign n35214 = pi1159 & ~n35213;
  assign n35215 = ~n35212 & n35214;
  assign n35216 = ~pi619 & n35210;
  assign n35217 = pi619 & ~n35056;
  assign n35218 = ~pi1159 & ~n35217;
  assign n35219 = ~n35216 & n35218;
  assign n35220 = ~n35215 & ~n35219;
  assign n35221 = pi789 & ~n35220;
  assign n35222 = ~n35211 & ~n35221;
  assign n35223 = ~n15832 & n35222;
  assign n35224 = n19771 & n35223;
  assign n35225 = ~n35057 & ~n35224;
  assign n35226 = ~pi644 & ~n35225;
  assign n35227 = pi644 & ~n35056;
  assign n35228 = pi715 & ~n35227;
  assign n35229 = ~n35226 & n35228;
  assign n35230 = n15765 & ~n35056;
  assign n35231 = ~n17585 & ~n35056;
  assign n35232 = n15747 & ~n35056;
  assign n35233 = pi680 & pi681;
  assign n35234 = n16345 & ~n35233;
  assign n35235 = ~pi223 & ~n16345;
  assign n35236 = pi223 & n16359;
  assign n35237 = ~pi299 & ~n35236;
  assign n35238 = ~n35234 & n35237;
  assign n35239 = ~n35235 & n35238;
  assign n35240 = pi223 & n16364;
  assign n35241 = n16350 & ~n35233;
  assign n35242 = ~pi223 & ~n16350;
  assign n35243 = pi299 & ~n35240;
  assign n35244 = ~n35241 & n35243;
  assign n35245 = ~n35242 & n35244;
  assign n35246 = ~pi39 & ~n35239;
  assign n35247 = ~n35245 & n35246;
  assign n35248 = pi681 & ~n34665;
  assign n35249 = ~n16121 & ~n35248;
  assign n35250 = n6194 & n35249;
  assign n35251 = pi681 & ~n16271;
  assign n35252 = ~n16103 & ~n35251;
  assign n35253 = ~n6194 & n35252;
  assign n35254 = pi223 & ~n35250;
  assign n35255 = ~n35253 & n35254;
  assign n35256 = pi681 & n16298;
  assign n35257 = n2608 & ~n35256;
  assign n35258 = ~n16308 & n35233;
  assign n35259 = n6194 & ~n35258;
  assign n35260 = pi681 & n34647;
  assign n35261 = ~n6194 & ~n35260;
  assign n35262 = ~n35259 & ~n35261;
  assign n35263 = ~n2608 & ~n35262;
  assign n35264 = ~pi223 & ~n35257;
  assign n35265 = ~n35263 & n35264;
  assign n35266 = ~n35255 & ~n35265;
  assign n35267 = ~pi299 & ~n35266;
  assign n35268 = ~pi223 & pi681;
  assign n35269 = n34675 & n35268;
  assign n35270 = n6221 & n35249;
  assign n35271 = ~n6221 & n35252;
  assign n35272 = pi223 & ~n35270;
  assign n35273 = ~n35271 & n35272;
  assign n35274 = pi215 & ~n35269;
  assign n35275 = ~n35273 & n35274;
  assign n35276 = n35138 & ~n35256;
  assign n35277 = ~n6221 & ~n35260;
  assign n35278 = n6221 & ~n35258;
  assign n35279 = ~pi223 & ~n35277;
  assign n35280 = ~n35278 & n35279;
  assign n35281 = pi681 & ~n16246;
  assign n35282 = n6221 & ~n16183;
  assign n35283 = ~n35281 & n35282;
  assign n35284 = pi681 & ~n34633;
  assign n35285 = ~pi681 & ~n16153;
  assign n35286 = ~n6221 & ~n35284;
  assign n35287 = ~n35285 & n35286;
  assign n35288 = pi223 & ~n35287;
  assign n35289 = ~n35283 & n35288;
  assign n35290 = ~n3302 & ~n35280;
  assign n35291 = ~n35289 & n35290;
  assign n35292 = ~n35276 & ~n35291;
  assign n35293 = ~pi215 & ~n35292;
  assign n35294 = pi299 & ~n35275;
  assign n35295 = ~n35293 & n35294;
  assign n35296 = pi39 & ~n35267;
  assign n35297 = ~n35295 & n35296;
  assign n35298 = ~n35247 & ~n35297;
  assign n35299 = ~pi38 & ~n35298;
  assign n35300 = pi681 & n16226;
  assign n35301 = pi223 & ~n16228;
  assign n35302 = pi38 & ~n35300;
  assign n35303 = ~n35301 & n35302;
  assign n35304 = n9829 & ~n35303;
  assign n35305 = ~n35299 & n35304;
  assign n35306 = ~n35058 & ~n35305;
  assign n35307 = ~pi778 & ~n35306;
  assign n35308 = pi625 & n35306;
  assign n35309 = ~pi625 & ~n35056;
  assign n35310 = pi1153 & ~n35309;
  assign n35311 = ~n35308 & n35310;
  assign n35312 = ~pi625 & n35306;
  assign n35313 = pi625 & ~n35056;
  assign n35314 = ~pi1153 & ~n35313;
  assign n35315 = ~n35312 & n35314;
  assign n35316 = ~n35311 & ~n35315;
  assign n35317 = pi778 & ~n35316;
  assign n35318 = ~n35307 & ~n35317;
  assign n35319 = ~n15741 & ~n35318;
  assign n35320 = n15741 & n35056;
  assign n35321 = ~n35319 & ~n35320;
  assign n35322 = ~n15747 & n35321;
  assign n35323 = ~n35232 & ~n35322;
  assign n35324 = ~n15753 & ~n35323;
  assign n35325 = ~n15759 & n35324;
  assign n35326 = ~n35231 & ~n35325;
  assign n35327 = ~n15765 & ~n35326;
  assign n35328 = ~n35230 & ~n35327;
  assign n35329 = ~pi787 & n35328;
  assign n35330 = n19394 & n35328;
  assign n35331 = ~n19394 & n35056;
  assign n35332 = ~n35330 & ~n35331;
  assign n35333 = pi787 & ~n35332;
  assign n35334 = ~n35329 & ~n35333;
  assign n35335 = pi644 & n35334;
  assign n35336 = n15832 & ~n35056;
  assign n35337 = ~n35223 & ~n35336;
  assign n35338 = ~n15925 & ~n35337;
  assign n35339 = n15925 & ~n35056;
  assign n35340 = n19478 & ~n35339;
  assign n35341 = ~n35338 & n35340;
  assign n35342 = ~n15959 & ~n35230;
  assign n35343 = ~n35332 & n35342;
  assign n35344 = ~n35341 & ~n35343;
  assign n35345 = pi787 & ~n35344;
  assign n35346 = pi628 & ~n35056;
  assign n35347 = ~pi628 & ~n35326;
  assign n35348 = n15923 & ~n35346;
  assign n35349 = ~n35347 & n35348;
  assign n35350 = ~n16633 & n35337;
  assign n35351 = ~pi628 & ~n35056;
  assign n35352 = pi628 & ~n35326;
  assign n35353 = n15922 & ~n35351;
  assign n35354 = ~n35352 & n35353;
  assign n35355 = ~n35349 & ~n35354;
  assign n35356 = ~n35350 & n35355;
  assign n35357 = pi792 & ~n35356;
  assign n35358 = n15753 & ~n35056;
  assign n35359 = ~n35324 & ~n35358;
  assign n35360 = n15828 & ~n35359;
  assign n35361 = ~pi626 & n35056;
  assign n35362 = pi626 & ~n35222;
  assign n35363 = n15756 & ~n35361;
  assign n35364 = ~n35362 & n35363;
  assign n35365 = pi626 & n35056;
  assign n35366 = ~pi626 & ~n35222;
  assign n35367 = n15757 & ~n35365;
  assign n35368 = ~n35366 & n35367;
  assign n35369 = ~n35360 & ~n35364;
  assign n35370 = ~n35368 & n35369;
  assign n35371 = pi788 & ~n35370;
  assign n35372 = pi609 & n35318;
  assign n35373 = n35061 & ~n35233;
  assign n35374 = ~pi642 & ~n16663;
  assign n35375 = n35233 & ~n35374;
  assign n35376 = ~n34772 & n35375;
  assign n35377 = ~n35373 & ~n35376;
  assign n35378 = n35062 & ~n35233;
  assign n35379 = ~n16679 & ~n35374;
  assign n35380 = n35233 & ~n35379;
  assign n35381 = n16065 & n35380;
  assign n35382 = pi223 & ~n35381;
  assign n35383 = ~n35378 & n35382;
  assign n35384 = n35377 & ~n35383;
  assign n35385 = n35064 & ~n35384;
  assign n35386 = n35060 & ~n35385;
  assign n35387 = n18052 & n35268;
  assign n35388 = n34940 & ~n35233;
  assign n35389 = ~n34944 & n35071;
  assign n35390 = ~n35388 & n35389;
  assign n35391 = n35069 & ~n35387;
  assign n35392 = ~n35390 & n35391;
  assign n35393 = n18060 & n35268;
  assign n35394 = n18059 & ~n35233;
  assign n35395 = ~n34931 & n35077;
  assign n35396 = ~n35394 & n35395;
  assign n35397 = n35075 & ~n35393;
  assign n35398 = ~n35396 & n35397;
  assign n35399 = ~pi39 & ~n35392;
  assign n35400 = ~n35398 & n35399;
  assign n35401 = ~n35103 & ~n35233;
  assign n35402 = n34113 & n35379;
  assign n35403 = pi680 & ~n35402;
  assign n35404 = n16094 & n35403;
  assign n35405 = pi642 & ~n16716;
  assign n35406 = ~n16720 & ~n35405;
  assign n35407 = ~pi616 & ~n35406;
  assign n35408 = n35404 & ~n35407;
  assign n35409 = ~n35401 & ~n35408;
  assign n35410 = ~n35108 & ~n35409;
  assign n35411 = n6194 & n35410;
  assign n35412 = ~n35098 & ~n35233;
  assign n35413 = ~n6160 & n16705;
  assign n35414 = n16679 & ~n16704;
  assign n35415 = pi642 & ~n35414;
  assign n35416 = n34795 & ~n35415;
  assign n35417 = ~n35413 & n35416;
  assign n35418 = ~n35412 & ~n35417;
  assign n35419 = ~n35097 & ~n35418;
  assign n35420 = ~n6194 & n35419;
  assign n35421 = pi223 & ~n35420;
  assign n35422 = ~n35411 & n35421;
  assign n35423 = n16063 & ~n35377;
  assign n35424 = n2608 & ~n35423;
  assign n35425 = ~n15724 & ~n16146;
  assign n35426 = ~pi603 & ~n35425;
  assign n35427 = ~n16765 & ~n35426;
  assign n35428 = n16452 & ~n35427;
  assign n35429 = pi642 & ~n34831;
  assign n35430 = ~n35425 & n35429;
  assign n35431 = ~pi642 & ~n6160;
  assign n35432 = ~n16768 & n35431;
  assign n35433 = pi680 & ~n35432;
  assign n35434 = ~n35430 & n35433;
  assign n35435 = ~n35428 & n35434;
  assign n35436 = pi642 & ~pi680;
  assign n35437 = n34831 & n35436;
  assign n35438 = ~n35435 & ~n35437;
  assign n35439 = pi681 & ~n35438;
  assign n35440 = ~pi681 & n35165;
  assign n35441 = ~n35439 & ~n35440;
  assign n35442 = ~n6194 & ~n35441;
  assign n35443 = n16464 & n35121;
  assign n35444 = n35120 & ~n35443;
  assign n35445 = ~pi680 & ~n35101;
  assign n35446 = pi642 & ~n16885;
  assign n35447 = n6160 & ~n35446;
  assign n35448 = ~pi642 & ~n16755;
  assign n35449 = n35447 & ~n35448;
  assign n35450 = n35403 & ~n35449;
  assign n35451 = ~n35445 & ~n35450;
  assign n35452 = pi681 & ~n35451;
  assign n35453 = ~n35444 & ~n35452;
  assign n35454 = n6194 & n35453;
  assign n35455 = ~n2608 & ~n35442;
  assign n35456 = ~n35454 & n35455;
  assign n35457 = ~pi223 & ~n35424;
  assign n35458 = ~n35456 & n35457;
  assign n35459 = ~pi299 & ~n35422;
  assign n35460 = ~n35458 & n35459;
  assign n35461 = n6221 & ~n35410;
  assign n35462 = ~n6221 & ~n35419;
  assign n35463 = pi223 & ~n35462;
  assign n35464 = ~n35461 & n35463;
  assign n35465 = ~n16794 & n35447;
  assign n35466 = n35403 & ~n35465;
  assign n35467 = ~n35445 & ~n35466;
  assign n35468 = pi681 & ~n35467;
  assign n35469 = n35130 & ~n35468;
  assign n35470 = ~n35127 & ~n35233;
  assign n35471 = ~n16792 & n35431;
  assign n35472 = n16793 & n17835;
  assign n35473 = n16452 & ~n35472;
  assign n35474 = pi642 & n34813;
  assign n35475 = pi680 & ~n35471;
  assign n35476 = ~n35474 & n35475;
  assign n35477 = ~n35473 & n35476;
  assign n35478 = ~n35470 & ~n35477;
  assign n35479 = n35128 & ~n35478;
  assign n35480 = ~pi223 & ~n35469;
  assign n35481 = ~n35479 & n35480;
  assign n35482 = pi215 & ~n35481;
  assign n35483 = ~n35464 & n35482;
  assign n35484 = n35138 & ~n35423;
  assign n35485 = ~n35145 & ~n35233;
  assign n35486 = ~n16687 & ~n35405;
  assign n35487 = n6160 & ~n35486;
  assign n35488 = n35404 & ~n35487;
  assign n35489 = ~n35485 & ~n35488;
  assign n35490 = n35150 & ~n35489;
  assign n35491 = ~n35156 & ~n35233;
  assign n35492 = pi642 & ~n34834;
  assign n35493 = n16452 & n34839;
  assign n35494 = n34832 & n35431;
  assign n35495 = pi680 & ~n35492;
  assign n35496 = ~n35493 & n35495;
  assign n35497 = ~n35494 & n35496;
  assign n35498 = ~n35491 & ~n35497;
  assign n35499 = n35161 & ~n35498;
  assign n35500 = ~n35490 & ~n35499;
  assign n35501 = pi223 & ~n35500;
  assign n35502 = n6221 & n35453;
  assign n35503 = ~n6221 & ~n35441;
  assign n35504 = ~pi223 & ~n35502;
  assign n35505 = ~n35503 & n35504;
  assign n35506 = ~n35501 & ~n35505;
  assign n35507 = ~n3302 & ~n35506;
  assign n35508 = ~pi215 & ~n35484;
  assign n35509 = ~n35507 & n35508;
  assign n35510 = pi299 & ~n35483;
  assign n35511 = ~n35509 & n35510;
  assign n35512 = pi39 & ~n35460;
  assign n35513 = ~n35511 & n35512;
  assign n35514 = ~pi38 & ~n35400;
  assign n35515 = ~n35513 & n35514;
  assign n35516 = n9829 & ~n35386;
  assign n35517 = ~n35515 & n35516;
  assign n35518 = ~n35058 & ~n35517;
  assign n35519 = ~pi625 & n35518;
  assign n35520 = pi625 & n35183;
  assign n35521 = ~pi1153 & ~n35519;
  assign n35522 = ~n35520 & n35521;
  assign n35523 = ~pi608 & ~n35522;
  assign n35524 = ~n35311 & n35523;
  assign n35525 = ~pi625 & n35183;
  assign n35526 = pi625 & n35518;
  assign n35527 = pi1153 & ~n35525;
  assign n35528 = ~n35526 & n35527;
  assign n35529 = pi608 & ~n35528;
  assign n35530 = ~n35315 & n35529;
  assign n35531 = ~n35524 & ~n35530;
  assign n35532 = pi778 & ~n35531;
  assign n35533 = ~pi778 & n35518;
  assign n35534 = ~n35532 & ~n35533;
  assign n35535 = ~pi609 & ~n35534;
  assign n35536 = ~pi1155 & ~n35372;
  assign n35537 = ~n35535 & n35536;
  assign n35538 = ~pi660 & ~n35191;
  assign n35539 = ~n35537 & n35538;
  assign n35540 = ~pi609 & n35318;
  assign n35541 = pi609 & ~n35534;
  assign n35542 = pi1155 & ~n35540;
  assign n35543 = ~n35541 & n35542;
  assign n35544 = pi660 & ~n35195;
  assign n35545 = ~n35543 & n35544;
  assign n35546 = ~n35539 & ~n35545;
  assign n35547 = pi785 & ~n35546;
  assign n35548 = ~pi785 & ~n35534;
  assign n35549 = ~n35547 & ~n35548;
  assign n35550 = ~pi618 & ~n35549;
  assign n35551 = pi618 & n35321;
  assign n35552 = ~pi1154 & ~n35551;
  assign n35553 = ~n35550 & n35552;
  assign n35554 = ~pi627 & ~n35203;
  assign n35555 = ~n35553 & n35554;
  assign n35556 = ~pi618 & n35321;
  assign n35557 = pi618 & ~n35549;
  assign n35558 = pi1154 & ~n35556;
  assign n35559 = ~n35557 & n35558;
  assign n35560 = pi627 & ~n35207;
  assign n35561 = ~n35559 & n35560;
  assign n35562 = ~n35555 & ~n35561;
  assign n35563 = pi781 & ~n35562;
  assign n35564 = ~pi781 & ~n35549;
  assign n35565 = ~n35563 & ~n35564;
  assign n35566 = ~pi789 & n35565;
  assign n35567 = ~pi619 & ~n35323;
  assign n35568 = pi619 & ~n35565;
  assign n35569 = pi1159 & ~n35567;
  assign n35570 = ~n35568 & n35569;
  assign n35571 = pi648 & ~n35219;
  assign n35572 = ~n35570 & n35571;
  assign n35573 = pi619 & ~n35323;
  assign n35574 = ~pi619 & ~n35565;
  assign n35575 = ~pi1159 & ~n35573;
  assign n35576 = ~n35574 & n35575;
  assign n35577 = ~pi648 & ~n35215;
  assign n35578 = ~n35576 & n35577;
  assign n35579 = pi789 & ~n35572;
  assign n35580 = ~n35578 & n35579;
  assign n35581 = n15833 & ~n35566;
  assign n35582 = ~n35580 & n35581;
  assign n35583 = ~n16644 & ~n35371;
  assign n35584 = ~n35582 & n35583;
  assign n35585 = ~n35357 & ~n35584;
  assign n35586 = n18841 & ~n35585;
  assign n35587 = ~n35345 & ~n35586;
  assign n35588 = ~pi644 & n35587;
  assign n35589 = ~pi715 & ~n35335;
  assign n35590 = ~n35588 & n35589;
  assign n35591 = ~pi1160 & ~n35229;
  assign n35592 = ~n35590 & n35591;
  assign n35593 = ~pi644 & n35334;
  assign n35594 = pi644 & n35587;
  assign n35595 = pi715 & ~n35593;
  assign n35596 = ~n35594 & n35595;
  assign n35597 = pi644 & ~n35225;
  assign n35598 = ~pi644 & ~n35056;
  assign n35599 = ~pi715 & ~n35598;
  assign n35600 = ~n35597 & n35599;
  assign n35601 = pi1160 & ~n35600;
  assign n35602 = ~n35596 & n35601;
  assign n35603 = ~n35592 & ~n35602;
  assign n35604 = pi790 & ~n35603;
  assign n35605 = ~pi790 & n35587;
  assign n35606 = ~n35604 & ~n35605;
  assign n35607 = ~po1038 & ~n35606;
  assign n35608 = ~pi223 & po1038;
  assign po380 = ~n35607 & ~n35608;
  assign n35610 = pi224 & ~n34455;
  assign n35611 = ~n28954 & ~n35610;
  assign n35612 = n15777 & ~n35610;
  assign n35613 = pi224 & ~n9829;
  assign n35614 = pi224 & ~n16228;
  assign n35615 = pi38 & ~n35614;
  assign n35616 = pi614 & n16570;
  assign n35617 = n35615 & ~n35616;
  assign n35618 = ~pi614 & n16519;
  assign n35619 = pi224 & ~n35618;
  assign n35620 = n16445 & n35619;
  assign n35621 = pi614 & n16519;
  assign n35622 = ~pi224 & n35621;
  assign n35623 = ~pi299 & ~n35622;
  assign n35624 = ~n35620 & n35623;
  assign n35625 = pi614 & n16524;
  assign n35626 = pi224 & n16431;
  assign n35627 = n35625 & ~n35626;
  assign n35628 = pi224 & ~n16051;
  assign n35629 = ~n35627 & ~n35628;
  assign n35630 = pi299 & n35629;
  assign n35631 = ~pi39 & ~n35624;
  assign n35632 = ~n35630 & n35631;
  assign n35633 = n16715 & ~n34507;
  assign n35634 = ~pi224 & n35633;
  assign n35635 = ~n16329 & n35634;
  assign n35636 = pi614 & ~n16487;
  assign n35637 = n34210 & ~n34815;
  assign n35638 = ~n35636 & ~n35637;
  assign n35639 = ~pi680 & ~n35638;
  assign n35640 = pi680 & ~n16491;
  assign n35641 = ~n34208 & n35640;
  assign n35642 = ~n35639 & ~n35641;
  assign n35643 = n16108 & ~n35642;
  assign n35644 = ~n16108 & ~n35638;
  assign n35645 = ~n35643 & ~n35644;
  assign n35646 = ~n6194 & n35645;
  assign n35647 = pi614 & n15780;
  assign n35648 = n16063 & ~n35647;
  assign n35649 = ~n6161 & ~n35648;
  assign n35650 = ~n34520 & ~n35649;
  assign n35651 = ~n16108 & ~n35650;
  assign n35652 = pi680 & n35647;
  assign n35653 = ~pi680 & ~n35650;
  assign n35654 = ~n16107 & ~n35652;
  assign n35655 = ~n35653 & n35654;
  assign n35656 = n16108 & ~n35655;
  assign n35657 = ~n35651 & ~n35656;
  assign n35658 = n6194 & n35657;
  assign n35659 = pi224 & ~n35646;
  assign n35660 = ~n35658 & n35659;
  assign n35661 = pi223 & ~n35635;
  assign n35662 = ~n35660 & n35661;
  assign n35663 = n5754 & ~n35083;
  assign n35664 = ~n16537 & ~n35663;
  assign n35665 = pi614 & ~n35664;
  assign n35666 = ~n16149 & ~n35647;
  assign n35667 = ~n16108 & ~n35666;
  assign n35668 = ~pi680 & ~n35666;
  assign n35669 = ~n16151 & ~n35652;
  assign n35670 = ~n35668 & n35669;
  assign n35671 = n16108 & ~n35670;
  assign n35672 = ~n35667 & ~n35671;
  assign n35673 = ~n6194 & n35672;
  assign n35674 = ~n16164 & ~n35649;
  assign n35675 = ~n16108 & ~n35674;
  assign n35676 = ~pi680 & ~n35674;
  assign n35677 = ~n16169 & ~n35652;
  assign n35678 = ~n35676 & n35677;
  assign n35679 = n16108 & ~n35678;
  assign n35680 = ~n35675 & ~n35679;
  assign n35681 = n6194 & n35680;
  assign n35682 = pi224 & ~n35673;
  assign n35683 = ~n35681 & n35682;
  assign n35684 = ~pi223 & ~n35665;
  assign n35685 = ~n35683 & n35684;
  assign n35686 = ~n35662 & ~n35685;
  assign n35687 = ~pi299 & ~n35686;
  assign n35688 = ~n16293 & n35634;
  assign n35689 = ~n6221 & n35645;
  assign n35690 = n6221 & n35657;
  assign n35691 = pi224 & ~n35689;
  assign n35692 = ~n35690 & n35691;
  assign n35693 = ~n35688 & ~n35692;
  assign n35694 = pi215 & ~n35693;
  assign n35695 = pi224 & ~n16063;
  assign n35696 = n3302 & ~n35695;
  assign n35697 = ~n16715 & n35696;
  assign n35698 = ~n6221 & n35672;
  assign n35699 = n6221 & n35680;
  assign n35700 = pi224 & ~n35698;
  assign n35701 = ~n35699 & n35700;
  assign n35702 = n34143 & n35647;
  assign n35703 = ~n6221 & ~n35702;
  assign n35704 = pi614 & n34496;
  assign n35705 = n6221 & ~n35704;
  assign n35706 = ~pi224 & ~n35703;
  assign n35707 = ~n35705 & n35706;
  assign n35708 = ~n3302 & ~n35707;
  assign n35709 = ~n35701 & n35708;
  assign n35710 = ~pi215 & ~n35697;
  assign n35711 = ~n35709 & n35710;
  assign n35712 = pi299 & ~n35694;
  assign n35713 = ~n35711 & n35712;
  assign n35714 = pi39 & ~n35687;
  assign n35715 = ~n35713 & n35714;
  assign n35716 = ~pi38 & ~n35632;
  assign n35717 = ~n35715 & n35716;
  assign n35718 = n9829 & ~n35617;
  assign n35719 = ~n35717 & n35718;
  assign n35720 = ~n35613 & ~n35719;
  assign n35721 = ~n15777 & n35720;
  assign n35722 = ~n35612 & ~n35721;
  assign n35723 = ~pi785 & n35722;
  assign n35724 = ~pi609 & ~n35610;
  assign n35725 = pi609 & ~n35722;
  assign n35726 = pi1155 & ~n35724;
  assign n35727 = ~n35725 & n35726;
  assign n35728 = pi609 & ~n35610;
  assign n35729 = ~pi609 & ~n35722;
  assign n35730 = ~pi1155 & ~n35728;
  assign n35731 = ~n35729 & n35730;
  assign n35732 = ~n35727 & ~n35731;
  assign n35733 = pi785 & ~n35732;
  assign n35734 = ~n35723 & ~n35733;
  assign n35735 = ~pi781 & ~n35734;
  assign n35736 = pi618 & n35734;
  assign n35737 = ~pi618 & ~n35610;
  assign n35738 = pi1154 & ~n35737;
  assign n35739 = ~n35736 & n35738;
  assign n35740 = ~pi618 & n35734;
  assign n35741 = pi618 & ~n35610;
  assign n35742 = ~pi1154 & ~n35741;
  assign n35743 = ~n35740 & n35742;
  assign n35744 = ~n35739 & ~n35743;
  assign n35745 = pi781 & ~n35744;
  assign n35746 = ~n35735 & ~n35745;
  assign n35747 = ~pi789 & ~n35746;
  assign n35748 = pi619 & n35746;
  assign n35749 = ~pi619 & ~n35610;
  assign n35750 = pi1159 & ~n35749;
  assign n35751 = ~n35748 & n35750;
  assign n35752 = ~pi619 & n35746;
  assign n35753 = pi619 & ~n35610;
  assign n35754 = ~pi1159 & ~n35753;
  assign n35755 = ~n35752 & n35754;
  assign n35756 = ~n35751 & ~n35755;
  assign n35757 = pi789 & ~n35756;
  assign n35758 = ~n35747 & ~n35757;
  assign n35759 = ~n15832 & n35758;
  assign n35760 = n19771 & n35759;
  assign n35761 = ~n35611 & ~n35760;
  assign n35762 = ~pi644 & ~n35761;
  assign n35763 = pi644 & ~n35610;
  assign n35764 = pi715 & ~n35763;
  assign n35765 = ~n35762 & n35764;
  assign n35766 = n15765 & ~n35610;
  assign n35767 = ~n17585 & ~n35610;
  assign n35768 = n15741 & ~n35610;
  assign n35769 = pi662 & n16226;
  assign n35770 = n35615 & ~n35769;
  assign n35771 = pi662 & pi680;
  assign n35772 = n16345 & ~n35771;
  assign n35773 = ~pi224 & ~n16345;
  assign n35774 = pi224 & n16359;
  assign n35775 = ~pi299 & ~n35774;
  assign n35776 = ~n35772 & n35775;
  assign n35777 = ~n35773 & n35776;
  assign n35778 = pi224 & n16364;
  assign n35779 = n16350 & ~n35771;
  assign n35780 = ~pi224 & ~n16350;
  assign n35781 = pi299 & ~n35778;
  assign n35782 = ~n35779 & n35781;
  assign n35783 = ~n35780 & n35782;
  assign n35784 = ~pi39 & ~n35777;
  assign n35785 = ~n35783 & n35784;
  assign n35786 = pi662 & n16322;
  assign n35787 = pi662 & n34647;
  assign n35788 = ~n6194 & ~n35787;
  assign n35789 = ~n16308 & n35771;
  assign n35790 = n6194 & ~n35789;
  assign n35791 = n5754 & ~n35788;
  assign n35792 = ~n35790 & n35791;
  assign n35793 = ~n6163 & ~n34633;
  assign n35794 = n16153 & ~n35793;
  assign n35795 = ~n6194 & n35794;
  assign n35796 = pi662 & ~n16246;
  assign n35797 = ~pi662 & ~n16184;
  assign n35798 = ~n35796 & ~n35797;
  assign n35799 = n6194 & n35798;
  assign n35800 = pi224 & ~n35795;
  assign n35801 = ~n35799 & n35800;
  assign n35802 = ~pi223 & ~n35786;
  assign n35803 = ~n35792 & n35802;
  assign n35804 = ~n35801 & n35803;
  assign n35805 = ~pi224 & pi662;
  assign n35806 = n16330 & n35805;
  assign n35807 = ~pi662 & ~n16122;
  assign n35808 = pi662 & ~n34665;
  assign n35809 = ~n35807 & ~n35808;
  assign n35810 = n6194 & n35809;
  assign n35811 = ~pi662 & ~n16104;
  assign n35812 = pi662 & ~n16271;
  assign n35813 = ~n35811 & ~n35812;
  assign n35814 = ~n6194 & n35813;
  assign n35815 = pi224 & ~n35810;
  assign n35816 = ~n35814 & n35815;
  assign n35817 = pi223 & ~n35806;
  assign n35818 = ~n35816 & n35817;
  assign n35819 = ~pi299 & ~n35818;
  assign n35820 = ~n35804 & n35819;
  assign n35821 = pi662 & n16298;
  assign n35822 = n35696 & ~n35821;
  assign n35823 = ~n6221 & n35794;
  assign n35824 = n6221 & n35798;
  assign n35825 = pi224 & ~n35823;
  assign n35826 = ~n35824 & n35825;
  assign n35827 = ~n6221 & ~n35787;
  assign n35828 = n6221 & ~n35789;
  assign n35829 = ~pi224 & ~n35827;
  assign n35830 = ~n35828 & n35829;
  assign n35831 = ~n3302 & ~n35830;
  assign n35832 = ~n35826 & n35831;
  assign n35833 = ~n35822 & ~n35832;
  assign n35834 = ~pi215 & ~n35833;
  assign n35835 = n34675 & n35805;
  assign n35836 = n6221 & n35809;
  assign n35837 = ~n6221 & n35813;
  assign n35838 = pi224 & ~n35836;
  assign n35839 = ~n35837 & n35838;
  assign n35840 = pi215 & ~n35835;
  assign n35841 = ~n35839 & n35840;
  assign n35842 = pi299 & ~n35841;
  assign n35843 = ~n35834 & n35842;
  assign n35844 = pi39 & ~n35820;
  assign n35845 = ~n35843 & n35844;
  assign n35846 = ~n35785 & ~n35845;
  assign n35847 = ~pi38 & ~n35846;
  assign n35848 = n9829 & ~n35770;
  assign n35849 = ~n35847 & n35848;
  assign n35850 = ~n35613 & ~n35849;
  assign n35851 = ~pi778 & ~n35850;
  assign n35852 = pi625 & n35850;
  assign n35853 = ~pi625 & ~n35610;
  assign n35854 = pi1153 & ~n35853;
  assign n35855 = ~n35852 & n35854;
  assign n35856 = ~pi625 & n35850;
  assign n35857 = pi625 & ~n35610;
  assign n35858 = ~pi1153 & ~n35857;
  assign n35859 = ~n35856 & n35858;
  assign n35860 = ~n35855 & ~n35859;
  assign n35861 = pi778 & ~n35860;
  assign n35862 = ~n35851 & ~n35861;
  assign n35863 = ~n15741 & n35862;
  assign n35864 = ~n35768 & ~n35863;
  assign n35865 = ~n15747 & ~n35864;
  assign n35866 = n15747 & ~n35610;
  assign n35867 = ~n35865 & ~n35866;
  assign n35868 = ~n15753 & ~n35867;
  assign n35869 = ~n15759 & n35868;
  assign n35870 = ~n35767 & ~n35869;
  assign n35871 = ~n15765 & ~n35870;
  assign n35872 = ~n35766 & ~n35871;
  assign n35873 = ~pi787 & n35872;
  assign n35874 = n19394 & n35872;
  assign n35875 = ~n19394 & n35610;
  assign n35876 = ~n35874 & ~n35875;
  assign n35877 = pi787 & ~n35876;
  assign n35878 = ~n35873 & ~n35877;
  assign n35879 = pi644 & n35878;
  assign n35880 = n15832 & ~n35610;
  assign n35881 = ~n35759 & ~n35880;
  assign n35882 = ~n15925 & ~n35881;
  assign n35883 = n15925 & ~n35610;
  assign n35884 = n19478 & ~n35883;
  assign n35885 = ~n35882 & n35884;
  assign n35886 = ~n15959 & ~n35766;
  assign n35887 = ~n35876 & n35886;
  assign n35888 = ~n35885 & ~n35887;
  assign n35889 = pi787 & ~n35888;
  assign n35890 = pi628 & ~n35610;
  assign n35891 = ~pi628 & ~n35870;
  assign n35892 = n15923 & ~n35890;
  assign n35893 = ~n35891 & n35892;
  assign n35894 = ~n16633 & n35881;
  assign n35895 = ~pi628 & ~n35610;
  assign n35896 = pi628 & ~n35870;
  assign n35897 = n15922 & ~n35895;
  assign n35898 = ~n35896 & n35897;
  assign n35899 = ~n35893 & ~n35898;
  assign n35900 = ~n35894 & n35899;
  assign n35901 = pi792 & ~n35900;
  assign n35902 = n15753 & ~n35610;
  assign n35903 = ~n35868 & ~n35902;
  assign n35904 = n15828 & ~n35903;
  assign n35905 = ~pi626 & n35610;
  assign n35906 = pi626 & ~n35758;
  assign n35907 = n15756 & ~n35905;
  assign n35908 = ~n35906 & n35907;
  assign n35909 = pi626 & n35610;
  assign n35910 = ~pi626 & ~n35758;
  assign n35911 = n15757 & ~n35909;
  assign n35912 = ~n35910 & n35911;
  assign n35913 = ~n35904 & ~n35908;
  assign n35914 = ~n35912 & n35913;
  assign n35915 = pi788 & ~n35914;
  assign n35916 = pi618 & ~n35864;
  assign n35917 = pi609 & n35862;
  assign n35918 = pi662 & n16664;
  assign n35919 = n16228 & n35918;
  assign n35920 = n35617 & ~n35919;
  assign n35921 = n18059 & n35771;
  assign n35922 = ~n35621 & ~n35921;
  assign n35923 = ~pi224 & ~n35922;
  assign n35924 = n18059 & ~n35771;
  assign n35925 = ~n34931 & n35619;
  assign n35926 = ~n35924 & n35925;
  assign n35927 = ~n35923 & ~n35926;
  assign n35928 = ~pi299 & ~n35927;
  assign n35929 = n35629 & ~n35771;
  assign n35930 = ~pi614 & n16524;
  assign n35931 = ~n34944 & ~n35930;
  assign n35932 = pi224 & ~n35931;
  assign n35933 = ~pi224 & ~n35625;
  assign n35934 = ~n34940 & n35933;
  assign n35935 = ~n35932 & ~n35934;
  assign n35936 = n35771 & ~n35935;
  assign n35937 = pi299 & ~n35929;
  assign n35938 = ~n35936 & n35937;
  assign n35939 = ~n35928 & ~n35938;
  assign n35940 = ~pi39 & ~n35939;
  assign n35941 = ~pi662 & n35633;
  assign n35942 = ~pi614 & n16751;
  assign n35943 = ~n34865 & ~n35942;
  assign n35944 = pi680 & ~n35943;
  assign n35945 = pi680 & ~n16787;
  assign n35946 = ~n16715 & ~n35945;
  assign n35947 = pi662 & ~n35944;
  assign n35948 = ~n35946 & n35947;
  assign n35949 = ~pi224 & ~n35941;
  assign n35950 = ~n35948 & n35949;
  assign n35951 = ~pi614 & ~n22848;
  assign n35952 = pi614 & ~n34772;
  assign n35953 = ~n35951 & ~n35952;
  assign n35954 = ~n16060 & n35953;
  assign n35955 = pi616 & ~n35954;
  assign n35956 = ~n16723 & ~n35955;
  assign n35957 = pi680 & ~n35956;
  assign n35958 = ~n35653 & ~n35957;
  assign n35959 = pi662 & ~n35958;
  assign n35960 = ~pi662 & ~n6162;
  assign n35961 = ~n35650 & n35960;
  assign n35962 = pi224 & ~n35961;
  assign n35963 = ~n35656 & n35962;
  assign n35964 = ~n35959 & n35963;
  assign n35965 = ~n35950 & ~n35964;
  assign n35966 = n6194 & n35965;
  assign n35967 = pi680 & ~n16709;
  assign n35968 = ~n35652 & ~n35967;
  assign n35969 = ~n35639 & n35968;
  assign n35970 = pi662 & ~n35969;
  assign n35971 = ~n35638 & n35960;
  assign n35972 = pi224 & ~n35971;
  assign n35973 = ~n35643 & n35972;
  assign n35974 = ~n35970 & n35973;
  assign n35975 = pi614 & n16530;
  assign n35976 = ~n34507 & n35975;
  assign n35977 = pi614 & ~n16808;
  assign n35978 = ~n16081 & n35977;
  assign n35979 = n16177 & n16797;
  assign n35980 = ~n35978 & ~n35979;
  assign n35981 = pi662 & ~n35980;
  assign n35982 = ~pi224 & ~n35976;
  assign n35983 = ~n35981 & n35982;
  assign n35984 = ~n35974 & ~n35983;
  assign n35985 = ~n6194 & n35984;
  assign n35986 = pi223 & ~n35985;
  assign n35987 = ~n35966 & n35986;
  assign n35988 = ~n15780 & n35821;
  assign n35989 = ~n16715 & ~n35988;
  assign n35990 = ~pi224 & ~n35989;
  assign n35991 = ~pi222 & n35990;
  assign n35992 = n16775 & n35771;
  assign n35993 = ~n35702 & ~n35992;
  assign n35994 = ~n6194 & n35993;
  assign n35995 = ~n16715 & ~n34885;
  assign n35996 = ~n35944 & ~n35995;
  assign n35997 = pi662 & ~n35996;
  assign n35998 = ~pi662 & ~n35704;
  assign n35999 = ~n35997 & ~n35998;
  assign n36000 = n6194 & ~n35999;
  assign n36001 = n5754 & ~n35994;
  assign n36002 = ~n36000 & n36001;
  assign n36003 = ~n35674 & n35960;
  assign n36004 = ~n16689 & ~n16717;
  assign n36005 = ~pi616 & ~n36004;
  assign n36006 = ~n35955 & ~n36005;
  assign n36007 = pi680 & ~n36006;
  assign n36008 = ~n35676 & ~n36007;
  assign n36009 = pi662 & ~n36008;
  assign n36010 = ~n35679 & ~n36003;
  assign n36011 = ~n36009 & n36010;
  assign n36012 = n6194 & n36011;
  assign n36013 = ~n35666 & n35960;
  assign n36014 = n34846 & ~n34874;
  assign n36015 = ~n35652 & ~n35668;
  assign n36016 = ~n36014 & n36015;
  assign n36017 = pi662 & ~n36016;
  assign n36018 = ~n35671 & ~n36013;
  assign n36019 = ~n36017 & n36018;
  assign n36020 = ~n6194 & n36019;
  assign n36021 = pi224 & ~n36020;
  assign n36022 = ~n36012 & n36021;
  assign n36023 = ~pi223 & ~n35991;
  assign n36024 = ~n36002 & n36023;
  assign n36025 = ~n36022 & n36024;
  assign n36026 = ~n35987 & ~n36025;
  assign n36027 = ~pi299 & ~n36026;
  assign n36028 = ~n6221 & ~n35984;
  assign n36029 = n6221 & ~n35965;
  assign n36030 = pi215 & ~n36028;
  assign n36031 = ~n36029 & n36030;
  assign n36032 = ~n35647 & ~n35771;
  assign n36033 = n16065 & n36032;
  assign n36034 = n35771 & n35953;
  assign n36035 = pi224 & ~n36033;
  assign n36036 = ~n36034 & n36035;
  assign n36037 = n35696 & ~n36036;
  assign n36038 = ~n35990 & n36037;
  assign n36039 = n6221 & ~n36011;
  assign n36040 = ~n6221 & ~n36019;
  assign n36041 = pi224 & ~n36040;
  assign n36042 = ~n36039 & n36041;
  assign n36043 = ~n6221 & ~n35993;
  assign n36044 = n6221 & n35999;
  assign n36045 = ~pi224 & ~n36043;
  assign n36046 = ~n36044 & n36045;
  assign n36047 = ~n36042 & ~n36046;
  assign n36048 = ~n3302 & ~n36047;
  assign n36049 = ~pi215 & ~n36038;
  assign n36050 = ~n36048 & n36049;
  assign n36051 = pi299 & ~n36031;
  assign n36052 = ~n36050 & n36051;
  assign n36053 = pi39 & ~n36027;
  assign n36054 = ~n36052 & n36053;
  assign n36055 = ~pi38 & ~n35940;
  assign n36056 = ~n36054 & n36055;
  assign n36057 = n9829 & ~n35920;
  assign n36058 = ~n36056 & n36057;
  assign n36059 = ~n35613 & ~n36058;
  assign n36060 = ~pi625 & n36059;
  assign n36061 = pi625 & n35720;
  assign n36062 = ~pi1153 & ~n36061;
  assign n36063 = ~n36060 & n36062;
  assign n36064 = ~pi608 & ~n35855;
  assign n36065 = ~n36063 & n36064;
  assign n36066 = ~pi625 & n35720;
  assign n36067 = pi625 & n36059;
  assign n36068 = pi1153 & ~n36066;
  assign n36069 = ~n36067 & n36068;
  assign n36070 = pi608 & ~n35859;
  assign n36071 = ~n36069 & n36070;
  assign n36072 = ~n36065 & ~n36071;
  assign n36073 = pi778 & ~n36072;
  assign n36074 = ~pi778 & n36059;
  assign n36075 = ~n36073 & ~n36074;
  assign n36076 = ~pi609 & ~n36075;
  assign n36077 = ~pi1155 & ~n35917;
  assign n36078 = ~n36076 & n36077;
  assign n36079 = ~pi660 & ~n35727;
  assign n36080 = ~n36078 & n36079;
  assign n36081 = ~pi609 & n35862;
  assign n36082 = pi609 & ~n36075;
  assign n36083 = pi1155 & ~n36081;
  assign n36084 = ~n36082 & n36083;
  assign n36085 = pi660 & ~n35731;
  assign n36086 = ~n36084 & n36085;
  assign n36087 = ~n36080 & ~n36086;
  assign n36088 = pi785 & ~n36087;
  assign n36089 = ~pi785 & ~n36075;
  assign n36090 = ~n36088 & ~n36089;
  assign n36091 = ~pi618 & ~n36090;
  assign n36092 = ~pi1154 & ~n35916;
  assign n36093 = ~n36091 & n36092;
  assign n36094 = ~pi627 & ~n35739;
  assign n36095 = ~n36093 & n36094;
  assign n36096 = ~pi618 & ~n35864;
  assign n36097 = pi618 & ~n36090;
  assign n36098 = pi1154 & ~n36096;
  assign n36099 = ~n36097 & n36098;
  assign n36100 = pi627 & ~n35743;
  assign n36101 = ~n36099 & n36100;
  assign n36102 = ~n36095 & ~n36101;
  assign n36103 = pi781 & ~n36102;
  assign n36104 = ~pi781 & ~n36090;
  assign n36105 = ~n36103 & ~n36104;
  assign n36106 = ~pi789 & n36105;
  assign n36107 = ~pi619 & ~n35867;
  assign n36108 = pi619 & ~n36105;
  assign n36109 = pi1159 & ~n36107;
  assign n36110 = ~n36108 & n36109;
  assign n36111 = pi648 & ~n35755;
  assign n36112 = ~n36110 & n36111;
  assign n36113 = pi619 & ~n35867;
  assign n36114 = ~pi619 & ~n36105;
  assign n36115 = ~pi1159 & ~n36113;
  assign n36116 = ~n36114 & n36115;
  assign n36117 = ~pi648 & ~n35751;
  assign n36118 = ~n36116 & n36117;
  assign n36119 = pi789 & ~n36112;
  assign n36120 = ~n36118 & n36119;
  assign n36121 = n15833 & ~n36106;
  assign n36122 = ~n36120 & n36121;
  assign n36123 = ~n16644 & ~n35915;
  assign n36124 = ~n36122 & n36123;
  assign n36125 = ~n35901 & ~n36124;
  assign n36126 = n18841 & ~n36125;
  assign n36127 = ~n35889 & ~n36126;
  assign n36128 = ~pi644 & n36127;
  assign n36129 = ~pi715 & ~n35879;
  assign n36130 = ~n36128 & n36129;
  assign n36131 = ~pi1160 & ~n35765;
  assign n36132 = ~n36130 & n36131;
  assign n36133 = ~pi644 & n35878;
  assign n36134 = pi644 & n36127;
  assign n36135 = pi715 & ~n36133;
  assign n36136 = ~n36134 & n36135;
  assign n36137 = pi644 & ~n35761;
  assign n36138 = ~pi644 & ~n35610;
  assign n36139 = ~pi715 & ~n36138;
  assign n36140 = ~n36137 & n36139;
  assign n36141 = pi1160 & ~n36140;
  assign n36142 = ~n36136 & n36141;
  assign n36143 = ~n36132 & ~n36142;
  assign n36144 = pi790 & ~n36143;
  assign n36145 = ~pi790 & n36127;
  assign n36146 = ~n36144 & ~n36145;
  assign n36147 = ~po1038 & ~n36146;
  assign n36148 = ~pi224 & po1038;
  assign po381 = ~n36147 & ~n36148;
  assign n36150 = n2554 & n2628;
  assign n36151 = n3316 & n36150;
  assign n36152 = ~pi62 & n36151;
  assign n36153 = ~n3291 & ~n36152;
  assign n36154 = pi62 & n36151;
  assign n36155 = n2535 & n36150;
  assign n36156 = pi54 & ~n36155;
  assign n36157 = pi92 & n2534;
  assign n36158 = n36150 & n36157;
  assign n36159 = ~n6090 & n6150;
  assign n36160 = ~pi137 & ~n36159;
  assign n36161 = n7228 & ~n36160;
  assign n36162 = pi75 & ~n36161;
  assign n36163 = pi87 & n36150;
  assign n36164 = n6083 & ~n36160;
  assign n36165 = pi38 & ~pi137;
  assign n36166 = pi39 & n2554;
  assign n36167 = ~n2740 & ~n2971;
  assign n36168 = pi137 & ~n36167;
  assign n36169 = ~n2739 & ~n36168;
  assign n36170 = ~pi332 & ~n36169;
  assign n36171 = n2737 & ~n11004;
  assign n36172 = ~pi137 & n2716;
  assign n36173 = ~n36171 & n36172;
  assign n36174 = n3149 & ~n11003;
  assign n36175 = ~n2904 & n36174;
  assign n36176 = n2745 & ~n36175;
  assign n36177 = n2743 & ~n36176;
  assign n36178 = ~n2715 & ~n36177;
  assign n36179 = ~pi95 & ~n36178;
  assign n36180 = n3069 & ~n36179;
  assign n36181 = pi332 & ~n36173;
  assign n36182 = ~n36180 & n36181;
  assign n36183 = ~n36170 & ~n36182;
  assign n36184 = pi210 & ~n36183;
  assign n36185 = n2920 & ~n36171;
  assign n36186 = pi1093 & ~n36185;
  assign n36187 = n2920 & n11104;
  assign n36188 = n2701 & ~n7387;
  assign n36189 = ~n2953 & n36188;
  assign n36190 = ~pi32 & ~n36189;
  assign n36191 = n36187 & ~n36190;
  assign n36192 = ~pi1093 & ~n36191;
  assign n36193 = ~n11104 & n36185;
  assign n36194 = n11002 & n36188;
  assign n36195 = n36187 & n36194;
  assign n36196 = ~n36193 & ~n36195;
  assign n36197 = n36192 & n36196;
  assign n36198 = ~n36186 & ~n36197;
  assign n36199 = n11140 & ~n36198;
  assign n36200 = ~n2919 & ~n36177;
  assign n36201 = ~pi95 & ~n36200;
  assign n36202 = ~n2740 & ~n36201;
  assign n36203 = pi137 & ~n36202;
  assign n36204 = n3010 & ~n11104;
  assign n36205 = n36192 & ~n36204;
  assign n36206 = ~n2982 & n36188;
  assign n36207 = ~pi32 & ~n36206;
  assign n36208 = n36187 & ~n36207;
  assign n36209 = pi1093 & ~n36204;
  assign n36210 = ~n36208 & n36209;
  assign n36211 = ~n36205 & ~n36210;
  assign n36212 = n11108 & ~n36211;
  assign n36213 = n36196 & n36212;
  assign n36214 = ~n36199 & ~n36213;
  assign n36215 = ~n36203 & n36214;
  assign n36216 = pi332 & ~n36215;
  assign n36217 = ~n2740 & ~n2978;
  assign n36218 = pi137 & ~n36217;
  assign n36219 = pi1093 & ~n3010;
  assign n36220 = ~n36205 & ~n36219;
  assign n36221 = n11140 & ~n36220;
  assign n36222 = ~n36212 & ~n36221;
  assign n36223 = ~n36218 & n36222;
  assign n36224 = ~pi332 & ~n36223;
  assign n36225 = ~n36216 & ~n36224;
  assign n36226 = ~n2666 & n36225;
  assign n36227 = ~pi137 & ~n36185;
  assign n36228 = ~n36203 & ~n36227;
  assign n36229 = pi332 & ~n36228;
  assign n36230 = ~n3011 & ~n36218;
  assign n36231 = ~pi332 & ~n36230;
  assign n36232 = ~n36229 & ~n36231;
  assign n36233 = n2666 & n36232;
  assign n36234 = ~pi210 & ~n36226;
  assign n36235 = ~n36233 & n36234;
  assign n36236 = pi299 & ~n36184;
  assign n36237 = ~n36235 & n36236;
  assign n36238 = pi198 & ~n36183;
  assign n36239 = ~n6320 & n36225;
  assign n36240 = n6320 & n36232;
  assign n36241 = ~pi198 & ~n36239;
  assign n36242 = ~n36240 & n36241;
  assign n36243 = ~pi299 & ~n36238;
  assign n36244 = ~n36242 & n36243;
  assign n36245 = ~n36237 & ~n36244;
  assign n36246 = ~pi39 & ~n36245;
  assign n36247 = ~pi38 & ~n36166;
  assign n36248 = ~n36246 & n36247;
  assign n36249 = n6118 & ~n36165;
  assign n36250 = ~n36248 & n36249;
  assign n36251 = ~n36164 & ~n36250;
  assign n36252 = ~pi87 & ~n36251;
  assign n36253 = ~pi75 & ~n36163;
  assign n36254 = ~n36252 & n36253;
  assign n36255 = ~pi92 & ~n36162;
  assign n36256 = ~n36254 & n36255;
  assign n36257 = ~pi54 & ~n36158;
  assign n36258 = ~n36256 & n36257;
  assign n36259 = ~pi74 & ~n36156;
  assign n36260 = ~n36258 & n36259;
  assign n36261 = pi74 & n6074;
  assign n36262 = n36150 & n36261;
  assign n36263 = ~pi55 & ~n36262;
  assign n36264 = ~n36260 & n36263;
  assign n36265 = n7278 & ~n36264;
  assign n36266 = pi56 & n2537;
  assign n36267 = n36150 & n36266;
  assign n36268 = ~n36265 & ~n36267;
  assign n36269 = ~pi62 & ~n36268;
  assign n36270 = n3291 & ~n36154;
  assign n36271 = ~n36269 & n36270;
  assign n36272 = ~n6068 & ~n36153;
  assign po382 = ~n36271 & n36272;
  assign n36274 = pi228 & pi231;
  assign n36275 = ~n7290 & ~n36274;
  assign n36276 = pi56 & ~n36275;
  assign n36277 = pi55 & ~n36274;
  assign n36278 = ~n7295 & ~n36274;
  assign n36279 = ~n6276 & ~n36274;
  assign n36280 = pi74 & ~n36279;
  assign n36281 = ~n36278 & n36280;
  assign n36282 = pi54 & ~n36274;
  assign n36283 = pi75 & ~n36278;
  assign n36284 = pi87 & ~n36274;
  assign n36285 = ~n7289 & n36284;
  assign n36286 = ~n7294 & ~n36274;
  assign n36287 = pi100 & ~n36286;
  assign n36288 = ~n2729 & ~n3105;
  assign n36289 = ~pi70 & ~n36288;
  assign n36290 = ~pi51 & ~n36289;
  assign n36291 = n2748 & ~n36290;
  assign n36292 = n3149 & ~n36291;
  assign n36293 = n2745 & ~n36292;
  assign n36294 = n2743 & ~n36293;
  assign n36295 = ~n6154 & ~n36294;
  assign n36296 = ~pi95 & ~n36295;
  assign n36297 = n2741 & ~n36296;
  assign n36298 = ~pi39 & ~n36297;
  assign n36299 = ~pi38 & ~n3378;
  assign n36300 = ~n36298 & n36299;
  assign n36301 = ~pi228 & n36300;
  assign n36302 = ~n36274 & ~n36301;
  assign n36303 = ~pi100 & ~n36302;
  assign n36304 = ~pi87 & ~n36287;
  assign n36305 = ~n36303 & n36304;
  assign n36306 = ~pi75 & ~n36285;
  assign n36307 = ~n36305 & n36306;
  assign n36308 = ~pi92 & ~n36283;
  assign n36309 = ~n36307 & n36308;
  assign n36310 = pi92 & ~n36274;
  assign n36311 = ~n7300 & n36310;
  assign n36312 = ~n36309 & ~n36311;
  assign n36313 = ~pi54 & ~n36312;
  assign n36314 = ~pi74 & ~n36282;
  assign n36315 = ~n36313 & n36314;
  assign n36316 = ~pi55 & ~n36281;
  assign n36317 = ~n36315 & n36316;
  assign n36318 = ~pi56 & ~n36277;
  assign n36319 = ~n36317 & n36318;
  assign n36320 = ~pi62 & ~n36276;
  assign n36321 = ~n36319 & n36320;
  assign n36322 = pi62 & ~n36274;
  assign n36323 = ~n7286 & n36322;
  assign n36324 = ~n36321 & ~n36323;
  assign n36325 = n3291 & ~n36324;
  assign n36326 = ~n3291 & ~n36274;
  assign po383 = ~n36325 & ~n36326;
  assign n36328 = n2711 & ~n6419;
  assign n36329 = ~pi91 & ~n2761;
  assign n36330 = ~n6102 & n10622;
  assign n36331 = n2754 & n10631;
  assign n36332 = n10629 & n36331;
  assign n36333 = n36329 & ~n36330;
  assign n36334 = ~n36332 & n36333;
  assign n36335 = n36328 & ~n36334;
  assign n36336 = ~pi72 & ~n36335;
  assign n36337 = n6432 & ~n36336;
  assign n36338 = n6176 & ~n36337;
  assign n36339 = n10643 & ~n12392;
  assign n36340 = n6432 & n36339;
  assign n36341 = ~n6340 & ~n36340;
  assign n36342 = pi1093 & ~n36341;
  assign n36343 = n36328 & ~n36329;
  assign n36344 = ~pi72 & ~n36343;
  assign n36345 = n10622 & n36328;
  assign n36346 = ~n7348 & n36345;
  assign n36347 = ~n8617 & n36344;
  assign n36348 = ~n36346 & n36347;
  assign n36349 = n6432 & ~n36348;
  assign n36350 = ~n36342 & ~n36349;
  assign n36351 = n36344 & ~n36345;
  assign n36352 = n6432 & ~n36351;
  assign n36353 = n6179 & ~n36352;
  assign n36354 = ~n36338 & ~n36353;
  assign n36355 = ~n36350 & n36354;
  assign n36356 = ~pi39 & ~n36355;
  assign po384 = ~n11061 | n36356;
  assign n36358 = ~pi39 & pi228;
  assign n36359 = n6348 & n12465;
  assign n36360 = ~n6178 & ~n8618;
  assign n36361 = n9824 & ~n36360;
  assign n36362 = n2958 & n36361;
  assign n36363 = ~n11076 & n36362;
  assign n36364 = ~n36359 & ~n36363;
  assign n36365 = n9833 & ~n36364;
  assign po385 = n36358 | n36365;
  assign n36367 = ~n6117 & n9830;
  assign n36368 = pi120 & n6181;
  assign n36369 = n16062 & ~n36368;
  assign n36370 = ~n33895 & ~n36369;
  assign n36371 = ~n6194 & ~n36370;
  assign n36372 = ~n6205 & n16062;
  assign n36373 = ~n36369 & ~n36372;
  assign n36374 = n6194 & ~n36373;
  assign n36375 = pi223 & ~n36371;
  assign n36376 = ~n36374 & n36375;
  assign n36377 = ~n6103 & n7453;
  assign n36378 = n16128 & n36377;
  assign n36379 = n16059 & ~n36377;
  assign n36380 = pi1091 & ~n36378;
  assign n36381 = ~n36379 & n36380;
  assign n36382 = n6336 & n16128;
  assign n36383 = ~n6336 & n16059;
  assign n36384 = ~pi1091 & ~n36382;
  assign n36385 = ~n36383 & n36384;
  assign n36386 = ~n36381 & ~n36385;
  assign n36387 = ~pi120 & ~n36386;
  assign n36388 = ~n16061 & ~n36387;
  assign n36389 = ~n6197 & n36388;
  assign n36390 = ~n33895 & ~n36389;
  assign n36391 = ~n6194 & n36390;
  assign n36392 = n6205 & n36388;
  assign n36393 = ~n36372 & ~n36392;
  assign n36394 = n6194 & n36393;
  assign n36395 = ~n2608 & ~n36391;
  assign n36396 = ~n36394 & n36395;
  assign n36397 = ~pi223 & ~n16231;
  assign n36398 = ~n36396 & n36397;
  assign n36399 = ~pi299 & ~n36376;
  assign n36400 = ~n36398 & n36399;
  assign n36401 = ~n6221 & ~n36370;
  assign n36402 = n6221 & ~n36373;
  assign n36403 = pi215 & ~n36401;
  assign n36404 = ~n36402 & n36403;
  assign n36405 = ~n6221 & n36390;
  assign n36406 = n6221 & n36393;
  assign n36407 = ~n3302 & ~n36405;
  assign n36408 = ~n36406 & n36407;
  assign n36409 = ~pi215 & ~n16316;
  assign n36410 = ~n36408 & n36409;
  assign n36411 = pi299 & ~n36404;
  assign n36412 = ~n36410 & n36411;
  assign n36413 = ~n36400 & ~n36412;
  assign n36414 = pi39 & ~n36413;
  assign n36415 = ~n6344 & n7348;
  assign n36416 = n16007 & ~n36415;
  assign n36417 = n6150 & ~n16024;
  assign n36418 = ~n6344 & ~n36417;
  assign n36419 = ~n36416 & ~n36418;
  assign n36420 = pi1091 & n16044;
  assign n36421 = pi1091 & ~n6344;
  assign n36422 = n11104 & n36421;
  assign n36423 = n36416 & ~n36422;
  assign n36424 = ~n6150 & ~n16038;
  assign n36425 = ~n36420 & n36424;
  assign n36426 = ~n36423 & n36425;
  assign n36427 = ~n36419 & ~n36426;
  assign n36428 = pi1093 & ~n36427;
  assign n36429 = n6130 & n8623;
  assign n36430 = ~n15997 & n36429;
  assign n36431 = ~pi40 & ~n36430;
  assign n36432 = n9914 & ~n36431;
  assign n36433 = pi252 & ~n36432;
  assign n36434 = n6104 & ~n15994;
  assign n36435 = ~n36433 & n36434;
  assign n36436 = ~n6104 & n16007;
  assign n36437 = ~pi1093 & ~n36435;
  assign n36438 = ~n36436 & n36437;
  assign n36439 = ~pi39 & ~n36438;
  assign n36440 = ~n36428 & n36439;
  assign n36441 = ~pi38 & ~n36440;
  assign n36442 = ~n36414 & n36441;
  assign po387 = n36367 & ~n36442;
  assign n36444 = ~pi81 & ~n2865;
  assign n36445 = n6392 & ~n36444;
  assign n36446 = n2464 & ~n36445;
  assign n36447 = n2873 & ~n36446;
  assign n36448 = n2783 & ~n36447;
  assign n36449 = n2877 & ~n36448;
  assign n36450 = n2719 & ~n36449;
  assign n36451 = ~n2722 & ~n36450;
  assign n36452 = ~pi86 & ~n36451;
  assign n36453 = n2780 & ~n36452;
  assign n36454 = n2778 & ~n36453;
  assign n36455 = ~n2775 & ~n36454;
  assign n36456 = ~pi108 & ~n36455;
  assign n36457 = n2774 & ~n36456;
  assign n36458 = n2890 & ~n36457;
  assign n36459 = ~n2766 & ~n36458;
  assign n36460 = n2765 & ~n36459;
  assign n36461 = n2764 & ~n36460;
  assign n36462 = n2757 & ~n36461;
  assign n36463 = n3090 & ~n36462;
  assign n36464 = n2516 & ~n36463;
  assign n36465 = n14767 & ~n36464;
  assign n36466 = ~pi70 & ~n36465;
  assign n36467 = ~n3081 & ~n36466;
  assign n36468 = ~pi51 & ~n36467;
  assign n36469 = n2748 & ~n36468;
  assign n36470 = n3149 & ~n36469;
  assign n36471 = n2745 & ~n36470;
  assign n36472 = ~pi1082 & n2742;
  assign n36473 = ~pi32 & ~n36472;
  assign n36474 = ~n36471 & n36473;
  assign n36475 = ~n3388 & ~n36474;
  assign n36476 = ~pi95 & ~n36475;
  assign n36477 = ~n2740 & ~n36476;
  assign n36478 = ~pi39 & ~n36477;
  assign po950 = ~n6102 | ~n6180;
  assign n36480 = n6334 & ~po950;
  assign n36481 = ~n11007 & n36480;
  assign n36482 = pi39 & n9857;
  assign n36483 = n6171 & n36482;
  assign n36484 = ~n36481 & n36483;
  assign n36485 = ~n3378 & ~n36484;
  assign n36486 = ~n36478 & n36485;
  assign n36487 = ~pi38 & ~n36486;
  assign n36488 = n6118 & ~n36487;
  assign n36489 = ~pi87 & ~n6083;
  assign n36490 = ~n36488 & n36489;
  assign n36491 = ~n6079 & ~n36490;
  assign n36492 = n2572 & ~n36491;
  assign n36493 = n7235 & ~n36492;
  assign n36494 = ~pi54 & ~n36493;
  assign n36495 = ~n7271 & ~n36494;
  assign n36496 = n6246 & ~n36495;
  assign n36497 = n14831 & ~n36496;
  assign n36498 = ~pi56 & ~n36497;
  assign n36499 = ~n6248 & ~n36498;
  assign n36500 = ~pi62 & ~n36499;
  assign n36501 = ~n6252 & ~n36500;
  assign n36502 = n3291 & ~n36501;
  assign po389 = n6071 & ~n36502;
  assign n36504 = ~pi230 & ~pi233;
  assign n36505 = pi199 & pi1142;
  assign n36506 = ~pi200 & ~n36505;
  assign n36507 = ~pi199 & pi1144;
  assign n36508 = n36506 & ~n36507;
  assign n36509 = ~pi199 & pi1143;
  assign n36510 = pi200 & ~n36509;
  assign n36511 = ~n36508 & ~n36510;
  assign n36512 = ~pi299 & ~n36511;
  assign n36513 = ~pi207 & ~n36512;
  assign n36514 = pi207 & ~pi299;
  assign n36515 = n36506 & ~n36509;
  assign n36516 = ~pi199 & pi1142;
  assign n36517 = pi200 & ~n36516;
  assign n36518 = n36514 & ~n36517;
  assign n36519 = ~n36515 & n36518;
  assign n36520 = ~n36513 & ~n36519;
  assign n36521 = pi208 & ~n36520;
  assign n36522 = pi207 & ~pi208;
  assign n36523 = n36511 & n36522;
  assign n36524 = ~n36521 & ~n36523;
  assign n36525 = n15574 & n36524;
  assign n36526 = pi211 & pi1143;
  assign n36527 = ~pi211 & pi1144;
  assign n36528 = ~n36526 & ~n36527;
  assign n36529 = ~n10332 & n36528;
  assign n36530 = ~pi211 & pi1143;
  assign n36531 = pi211 & pi1142;
  assign n36532 = n10332 & ~n36530;
  assign n36533 = ~n36531 & n36532;
  assign n36534 = ~n36529 & ~n36533;
  assign n36535 = ~pi219 & ~n36534;
  assign n36536 = ~pi212 & ~pi214;
  assign n36537 = ~pi211 & pi1142;
  assign n36538 = pi219 & ~n36537;
  assign n36539 = ~n36536 & ~n36538;
  assign n36540 = ~n36535 & n36539;
  assign n36541 = ~n15574 & ~n36540;
  assign n36542 = ~n36525 & ~n36541;
  assign n36543 = pi213 & ~n36542;
  assign n36544 = ~pi212 & pi214;
  assign n36545 = pi299 & pi1155;
  assign n36546 = n36544 & n36545;
  assign n36547 = pi299 & pi1153;
  assign n36548 = pi214 & ~n36547;
  assign n36549 = pi299 & pi1154;
  assign n36550 = ~pi214 & ~n36549;
  assign n36551 = pi212 & ~n36548;
  assign n36552 = ~n36550 & n36551;
  assign n36553 = ~n36546 & ~n36552;
  assign n36554 = ~pi211 & pi219;
  assign n36555 = ~n36553 & n36554;
  assign n36556 = ~pi299 & ~n36524;
  assign n36557 = ~pi211 & pi1157;
  assign n36558 = pi211 & pi1156;
  assign n36559 = ~n36557 & ~n36558;
  assign n36560 = n36544 & ~n36559;
  assign n36561 = ~pi211 & pi1155;
  assign n36562 = pi211 & pi1154;
  assign n36563 = ~n36561 & ~n36562;
  assign n36564 = pi214 & n36563;
  assign n36565 = ~pi211 & pi1156;
  assign n36566 = pi211 & pi1155;
  assign n36567 = ~n36565 & ~n36566;
  assign n36568 = ~pi214 & n36567;
  assign n36569 = pi212 & ~n36564;
  assign n36570 = ~n36568 & n36569;
  assign n36571 = ~n36560 & ~n36570;
  assign n36572 = ~pi219 & pi299;
  assign n36573 = ~n36571 & n36572;
  assign n36574 = ~n36555 & ~n36573;
  assign n36575 = ~n36556 & n36574;
  assign n36576 = ~po1038 & ~n36575;
  assign n36577 = ~pi219 & ~n36560;
  assign n36578 = ~n36570 & n36577;
  assign n36579 = ~pi211 & pi1154;
  assign n36580 = ~pi214 & ~n36579;
  assign n36581 = ~pi211 & pi1153;
  assign n36582 = n10332 & ~n36581;
  assign n36583 = ~pi211 & pi214;
  assign n36584 = pi1155 & n36583;
  assign n36585 = ~pi212 & ~n36584;
  assign n36586 = ~n36580 & ~n36582;
  assign n36587 = ~n36585 & n36586;
  assign n36588 = pi219 & ~n36587;
  assign n36589 = po1038 & ~n36588;
  assign n36590 = ~n36578 & n36589;
  assign n36591 = ~pi213 & ~n36590;
  assign n36592 = ~n36576 & n36591;
  assign n36593 = pi209 & ~n36543;
  assign n36594 = ~n36592 & n36593;
  assign n36595 = po1038 & n36540;
  assign n36596 = pi299 & pi1143;
  assign n36597 = pi199 & pi200;
  assign n36598 = ~pi299 & ~n36597;
  assign n36599 = pi1153 & ~n36598;
  assign n36600 = pi1154 & ~n36599;
  assign n36601 = ~pi200 & pi1155;
  assign n36602 = n10970 & n36601;
  assign n36603 = ~n10421 & ~n36597;
  assign n36604 = ~pi1153 & ~n10970;
  assign n36605 = pi1154 & n36603;
  assign n36606 = ~n36604 & n36605;
  assign n36607 = ~n36602 & ~n36606;
  assign n36608 = n36600 & ~n36607;
  assign n36609 = ~pi199 & ~pi1155;
  assign n36610 = ~pi200 & ~pi299;
  assign n36611 = pi199 & ~pi1153;
  assign n36612 = n36610 & ~n36611;
  assign n36613 = ~pi1154 & ~n36609;
  assign n36614 = n36612 & n36613;
  assign n36615 = ~n36608 & ~n36614;
  assign n36616 = pi207 & n36615;
  assign n36617 = ~n36596 & n36616;
  assign n36618 = ~pi199 & pi1155;
  assign n36619 = pi200 & ~pi299;
  assign n36620 = n36618 & n36619;
  assign n36621 = ~pi1154 & ~n36620;
  assign n36622 = ~n36596 & n36621;
  assign n36623 = ~pi1155 & n36596;
  assign n36624 = ~pi299 & ~n36603;
  assign n36625 = pi1155 & ~n36624;
  assign n36626 = pi299 & ~pi1143;
  assign n36627 = n36625 & ~n36626;
  assign n36628 = pi199 & ~pi200;
  assign n36629 = ~pi299 & n36628;
  assign n36630 = ~pi1155 & n36629;
  assign n36631 = pi1154 & ~n36630;
  assign n36632 = ~n36623 & n36631;
  assign n36633 = ~n36627 & n36632;
  assign n36634 = ~pi1156 & ~n36622;
  assign n36635 = ~n36633 & n36634;
  assign n36636 = pi200 & ~n36618;
  assign n36637 = ~pi299 & ~n36636;
  assign n36638 = pi1154 & ~n36637;
  assign n36639 = ~n36596 & n36638;
  assign n36640 = pi1155 & ~n10957;
  assign n36641 = ~pi1155 & ~n10422;
  assign n36642 = ~n36640 & ~n36641;
  assign n36643 = ~n36626 & ~n36642;
  assign n36644 = ~pi1154 & ~n36643;
  assign n36645 = pi1156 & ~n36639;
  assign n36646 = ~n36644 & n36645;
  assign n36647 = ~n36635 & ~n36646;
  assign n36648 = ~pi207 & n36647;
  assign n36649 = pi208 & ~n36617;
  assign n36650 = ~n36648 & n36649;
  assign n36651 = pi1155 & n36629;
  assign n36652 = ~pi1156 & ~n36651;
  assign n36653 = pi1155 & n36628;
  assign n36654 = ~pi299 & ~n11035;
  assign n36655 = pi1156 & ~n36653;
  assign n36656 = n36654 & n36655;
  assign n36657 = ~n36652 & ~n36656;
  assign n36658 = ~pi299 & ~n36657;
  assign n36659 = ~pi207 & ~pi299;
  assign n36660 = ~pi208 & ~n36659;
  assign n36661 = ~n36658 & n36660;
  assign n36662 = ~pi1157 & n36661;
  assign n36663 = ~pi208 & pi1157;
  assign n36664 = pi1155 & ~n36619;
  assign n36665 = ~n36641 & ~n36664;
  assign n36666 = pi199 & ~pi1155;
  assign n36667 = pi1156 & ~n36666;
  assign n36668 = n36598 & n36667;
  assign n36669 = n36665 & ~n36668;
  assign n36670 = ~n36659 & n36663;
  assign n36671 = ~n36669 & n36670;
  assign n36672 = ~n36662 & ~n36671;
  assign n36673 = ~pi208 & ~n36626;
  assign n36674 = ~n36672 & n36673;
  assign n36675 = ~n10332 & ~n36536;
  assign n36676 = pi211 & ~n36675;
  assign n36677 = ~n10335 & ~n36676;
  assign n36678 = ~n36674 & n36677;
  assign n36679 = ~n36650 & n36678;
  assign n36680 = pi299 & ~pi1144;
  assign n36681 = ~n36672 & ~n36680;
  assign n36682 = pi207 & ~n36615;
  assign n36683 = pi299 & pi1144;
  assign n36684 = n36621 & ~n36683;
  assign n36685 = ~pi1155 & n36683;
  assign n36686 = n36625 & ~n36680;
  assign n36687 = n36631 & ~n36685;
  assign n36688 = ~n36686 & n36687;
  assign n36689 = ~pi1156 & ~n36684;
  assign n36690 = ~n36688 & n36689;
  assign n36691 = n36638 & ~n36683;
  assign n36692 = ~n36642 & ~n36680;
  assign n36693 = ~pi1154 & ~n36692;
  assign n36694 = pi1156 & ~n36691;
  assign n36695 = ~n36693 & n36694;
  assign n36696 = ~n36690 & ~n36695;
  assign n36697 = ~pi207 & ~n36696;
  assign n36698 = pi207 & n36683;
  assign n36699 = ~n36682 & ~n36698;
  assign n36700 = ~n36697 & n36699;
  assign n36701 = pi208 & ~n36700;
  assign n36702 = n10335 & ~n36536;
  assign n36703 = ~n36681 & n36702;
  assign n36704 = ~n36701 & n36703;
  assign n36705 = ~n36679 & ~n36704;
  assign n36706 = ~pi219 & ~n36705;
  assign n36707 = ~pi299 & n36603;
  assign n36708 = ~n36666 & n36707;
  assign n36709 = ~n36652 & n36708;
  assign n36710 = pi207 & n36709;
  assign n36711 = ~pi208 & ~n36710;
  assign n36712 = n10422 & ~n36636;
  assign n36713 = ~n36621 & n36712;
  assign n36714 = pi200 & ~pi1155;
  assign n36715 = n10970 & ~n36714;
  assign n36716 = pi1156 & n36715;
  assign n36717 = ~n36713 & ~n36716;
  assign n36718 = ~n10101 & n36717;
  assign n36719 = ~n36616 & ~n36718;
  assign n36720 = pi208 & ~n36719;
  assign n36721 = ~n36711 & ~n36720;
  assign n36722 = ~pi1157 & ~n36721;
  assign n36723 = ~pi1156 & n36610;
  assign n36724 = ~n36666 & n36723;
  assign n36725 = ~n36668 & ~n36724;
  assign n36726 = pi207 & ~n36725;
  assign n36727 = ~pi208 & ~n36726;
  assign n36728 = ~n36720 & ~n36727;
  assign n36729 = pi1157 & ~n36728;
  assign n36730 = ~n36722 & ~n36729;
  assign n36731 = ~pi211 & ~n36536;
  assign n36732 = ~pi219 & ~n36536;
  assign n36733 = ~n36731 & ~n36732;
  assign n36734 = ~n36730 & n36733;
  assign n36735 = pi299 & ~pi1142;
  assign n36736 = ~n36611 & n36707;
  assign n36737 = ~n36640 & ~n36736;
  assign n36738 = ~pi1154 & n36619;
  assign n36739 = ~n36737 & ~n36738;
  assign n36740 = ~pi299 & ~n36739;
  assign n36741 = ~n36735 & ~n36740;
  assign n36742 = pi207 & ~n36741;
  assign n36743 = ~pi299 & ~n36628;
  assign n36744 = ~pi1155 & ~n36743;
  assign n36745 = ~n36625 & ~n36744;
  assign n36746 = pi1154 & ~n36745;
  assign n36747 = pi1156 & ~n36642;
  assign n36748 = ~n36746 & ~n36747;
  assign n36749 = ~n36735 & ~n36748;
  assign n36750 = pi299 & pi1142;
  assign n36751 = ~n36620 & ~n36750;
  assign n36752 = ~pi1154 & ~pi1156;
  assign n36753 = ~n36751 & n36752;
  assign n36754 = ~pi207 & ~n36753;
  assign n36755 = ~n36749 & n36754;
  assign n36756 = pi208 & ~n36742;
  assign n36757 = ~n36755 & n36756;
  assign n36758 = ~pi1157 & ~n36661;
  assign n36759 = n10957 & ~n36601;
  assign n36760 = pi1156 & ~n36759;
  assign n36761 = n36665 & ~n36760;
  assign n36762 = n36660 & ~n36761;
  assign n36763 = pi1157 & ~n36762;
  assign n36764 = ~n36735 & ~n36763;
  assign n36765 = ~n36758 & n36764;
  assign n36766 = ~n10100 & ~n36733;
  assign n36767 = ~n36765 & n36766;
  assign n36768 = ~n36757 & n36767;
  assign n36769 = ~po1038 & ~n36768;
  assign n36770 = ~n36706 & n36769;
  assign n36771 = ~n36734 & n36770;
  assign n36772 = pi213 & ~n36595;
  assign n36773 = ~n36771 & n36772;
  assign n36774 = ~pi207 & ~n36545;
  assign n36775 = ~pi208 & ~n36774;
  assign n36776 = ~pi1155 & ~n10970;
  assign n36777 = ~pi299 & n36652;
  assign n36778 = ~n36624 & ~n36776;
  assign n36779 = ~n36777 & n36778;
  assign n36780 = pi1157 & n12341;
  assign n36781 = ~n36779 & ~n36780;
  assign n36782 = n36775 & ~n36781;
  assign n36783 = pi207 & ~n36739;
  assign n36784 = ~n36545 & n36717;
  assign n36785 = ~pi207 & n36784;
  assign n36786 = pi208 & ~n36783;
  assign n36787 = ~n36785 & n36786;
  assign n36788 = ~n36782 & ~n36787;
  assign n36789 = ~pi211 & ~pi214;
  assign n36790 = ~n10098 & ~n36789;
  assign n36791 = ~n36788 & n36790;
  assign n36792 = n36717 & ~n36746;
  assign n36793 = ~pi207 & ~n36792;
  assign n36794 = ~pi299 & n36737;
  assign n36795 = pi1154 & ~n36794;
  assign n36796 = ~n36614 & ~n36795;
  assign n36797 = pi207 & ~n36796;
  assign n36798 = ~n36793 & ~n36797;
  assign n36799 = pi208 & ~n36798;
  assign n36800 = ~n36549 & ~n36710;
  assign n36801 = ~pi208 & ~n36800;
  assign n36802 = pi299 & ~pi1154;
  assign n36803 = pi1157 & ~n36802;
  assign n36804 = ~n36801 & ~n36803;
  assign n36805 = ~n36763 & ~n36804;
  assign n36806 = ~n36799 & ~n36805;
  assign n36807 = n10098 & ~n36806;
  assign n36808 = ~n36652 & n36661;
  assign n36809 = ~n36713 & ~n36747;
  assign n36810 = ~n36514 & ~n36809;
  assign n36811 = ~n36682 & ~n36810;
  assign n36812 = pi208 & ~n36811;
  assign n36813 = pi299 & pi1156;
  assign n36814 = ~n36726 & ~n36813;
  assign n36815 = n36663 & ~n36814;
  assign n36816 = ~n36808 & ~n36815;
  assign n36817 = ~n36812 & n36816;
  assign n36818 = n36789 & ~n36817;
  assign n36819 = ~n36791 & ~n36818;
  assign n36820 = ~n36807 & n36819;
  assign n36821 = pi212 & ~n36820;
  assign n36822 = ~pi214 & ~n36730;
  assign n36823 = ~pi212 & ~n36822;
  assign n36824 = pi211 & ~n36817;
  assign n36825 = pi299 & ~pi1155;
  assign n36826 = pi1155 & ~n36654;
  assign n36827 = ~n36825 & ~n36826;
  assign n36828 = n36748 & n36827;
  assign n36829 = ~pi207 & n36828;
  assign n36830 = pi1153 & ~n36743;
  assign n36831 = n36607 & ~n36830;
  assign n36832 = n36514 & n36831;
  assign n36833 = pi208 & ~n36832;
  assign n36834 = ~n36829 & n36833;
  assign n36835 = n36763 & ~n36834;
  assign n36836 = ~pi211 & ~n36835;
  assign n36837 = ~n36722 & n36836;
  assign n36838 = pi214 & ~n36824;
  assign n36839 = ~n36837 & n36838;
  assign n36840 = n36823 & ~n36839;
  assign n36841 = ~n36821 & ~n36840;
  assign n36842 = ~pi219 & ~n36841;
  assign n36843 = pi211 & ~n36730;
  assign n36844 = n36583 & n36788;
  assign n36845 = n36823 & ~n36844;
  assign n36846 = pi207 & ~n36831;
  assign n36847 = pi299 & ~pi1153;
  assign n36848 = ~pi207 & ~n36847;
  assign n36849 = ~n36828 & n36848;
  assign n36850 = ~n36846 & ~n36849;
  assign n36851 = pi208 & ~n36850;
  assign n36852 = ~n36763 & ~n36847;
  assign n36853 = ~n36758 & n36852;
  assign n36854 = n36583 & ~n36853;
  assign n36855 = ~n36851 & n36854;
  assign n36856 = n36789 & n36806;
  assign n36857 = pi212 & ~n36855;
  assign n36858 = ~n36856 & n36857;
  assign n36859 = ~n36845 & ~n36858;
  assign n36860 = pi219 & ~n36843;
  assign n36861 = ~n36859 & n36860;
  assign n36862 = ~n36842 & ~n36861;
  assign n36863 = ~po1038 & ~n36862;
  assign n36864 = n36591 & ~n36863;
  assign n36865 = ~pi209 & ~n36773;
  assign n36866 = ~n36864 & n36865;
  assign n36867 = ~n36594 & ~n36866;
  assign n36868 = pi230 & ~n36867;
  assign po390 = n36504 | n36868;
  assign n36870 = ~pi230 & pi234;
  assign n36871 = pi211 & pi1153;
  assign n36872 = ~n36579 & ~n36871;
  assign n36873 = ~n10332 & n36872;
  assign n36874 = n36732 & ~n36873;
  assign n36875 = ~n36582 & n36874;
  assign n36876 = po1038 & n36875;
  assign n36877 = ~pi1152 & ~n36876;
  assign n36878 = ~pi207 & ~pi208;
  assign n36879 = ~n10101 & ~n36878;
  assign n36880 = pi1154 & ~n36624;
  assign n36881 = ~n36602 & ~n36880;
  assign n36882 = pi207 & ~n36881;
  assign n36883 = ~pi299 & n36882;
  assign n36884 = ~n36879 & ~n36883;
  assign n36885 = ~n36718 & ~n36884;
  assign n36886 = ~pi214 & ~n36885;
  assign n36887 = ~pi212 & ~n36886;
  assign n36888 = pi207 & ~n36792;
  assign n36889 = ~n36549 & ~n36888;
  assign n36890 = ~pi208 & ~n36889;
  assign n36891 = ~n36793 & ~n36882;
  assign n36892 = pi208 & ~n36891;
  assign n36893 = ~n36890 & ~n36892;
  assign n36894 = ~pi211 & ~n36893;
  assign n36895 = pi208 & pi299;
  assign n36896 = pi207 & n36828;
  assign n36897 = n36660 & ~n36896;
  assign n36898 = ~n36810 & ~n36883;
  assign n36899 = pi208 & ~n36898;
  assign n36900 = ~n36895 & ~n36899;
  assign n36901 = ~n36897 & n36900;
  assign n36902 = ~n36847 & ~n36901;
  assign n36903 = pi211 & n36902;
  assign n36904 = ~n36894 & ~n36903;
  assign n36905 = pi214 & n36904;
  assign n36906 = n36887 & ~n36905;
  assign n36907 = ~pi219 & ~n36906;
  assign n36908 = ~pi214 & ~n36904;
  assign n36909 = ~pi211 & ~n36902;
  assign n36910 = pi214 & ~n36909;
  assign n36911 = pi211 & ~n36885;
  assign n36912 = n36910 & ~n36911;
  assign n36913 = ~n36908 & ~n36912;
  assign n36914 = pi212 & ~n36913;
  assign n36915 = n36907 & ~n36914;
  assign n36916 = pi219 & ~n36885;
  assign n36917 = ~po1038 & ~n36916;
  assign n36918 = ~n36915 & n36917;
  assign n36919 = n36877 & ~n36918;
  assign n36920 = pi219 & ~n36731;
  assign n36921 = po1038 & ~n36920;
  assign n36922 = pi1153 & ~n36789;
  assign n36923 = ~n36580 & ~n36583;
  assign n36924 = ~n36922 & ~n36923;
  assign n36925 = pi212 & ~n36924;
  assign n36926 = n36544 & ~n36872;
  assign n36927 = ~pi219 & ~n36926;
  assign n36928 = ~n36925 & n36927;
  assign n36929 = n36921 & ~n36928;
  assign n36930 = pi1152 & ~n36929;
  assign n36931 = ~n36901 & n36910;
  assign n36932 = ~n36908 & ~n36931;
  assign n36933 = pi212 & ~n36932;
  assign n36934 = n36907 & ~n36933;
  assign n36935 = ~n36731 & n36885;
  assign n36936 = pi219 & ~n36935;
  assign n36937 = n36731 & ~n36901;
  assign n36938 = n36936 & ~n36937;
  assign n36939 = ~po1038 & ~n36938;
  assign n36940 = ~n36934 & n36939;
  assign n36941 = n36930 & ~n36940;
  assign n36942 = ~pi213 & ~n36919;
  assign n36943 = ~n36941 & n36942;
  assign n36944 = ~n36536 & n36894;
  assign n36945 = n36936 & ~n36944;
  assign n36946 = n36660 & ~n36809;
  assign n36947 = ~n36899 & ~n36946;
  assign n36948 = ~pi211 & ~n36947;
  assign n36949 = ~n36545 & ~n36885;
  assign n36950 = pi211 & ~n36949;
  assign n36951 = ~n36948 & ~n36950;
  assign n36952 = pi214 & n36951;
  assign n36953 = n36887 & ~n36952;
  assign n36954 = pi211 & ~n36893;
  assign n36955 = ~pi211 & ~n36949;
  assign n36956 = pi214 & ~n36955;
  assign n36957 = ~n36954 & n36956;
  assign n36958 = ~pi214 & n36951;
  assign n36959 = pi212 & ~n36957;
  assign n36960 = ~n36958 & n36959;
  assign n36961 = ~pi219 & ~n36953;
  assign n36962 = ~n36960 & n36961;
  assign n36963 = n34036 & ~n36945;
  assign n36964 = ~n36962 & n36963;
  assign n36965 = ~n36943 & ~n36964;
  assign n36966 = pi209 & ~n36965;
  assign n36967 = ~pi1153 & ~n12341;
  assign n36968 = n36600 & ~n36967;
  assign n36969 = ~pi199 & ~pi1153;
  assign n36970 = n36707 & ~n36969;
  assign n36971 = ~n36968 & ~n36970;
  assign n36972 = pi208 & n36514;
  assign n36973 = n36971 & ~n36972;
  assign n36974 = ~pi299 & n36597;
  assign n36975 = ~pi1153 & ~n10422;
  assign n36976 = n10101 & ~n36974;
  assign n36977 = ~n36975 & n36976;
  assign n36978 = ~n36660 & ~n36879;
  assign n36979 = ~n36977 & n36978;
  assign n36980 = ~n36973 & ~n36979;
  assign n36981 = pi211 & ~n36980;
  assign n36982 = ~pi200 & ~pi1153;
  assign n36983 = ~pi199 & ~n36982;
  assign n36984 = ~pi299 & ~n36983;
  assign n36985 = ~n36628 & n36984;
  assign n36986 = pi207 & ~n36985;
  assign n36987 = pi1153 & n11036;
  assign n36988 = pi1154 & ~n36619;
  assign n36989 = ~n36987 & ~n36988;
  assign n36990 = n36743 & n36989;
  assign n36991 = ~pi207 & ~n36990;
  assign n36992 = ~n36986 & ~n36991;
  assign n36993 = pi208 & ~n36992;
  assign n36994 = n36660 & ~n36990;
  assign n36995 = ~n36993 & ~n36994;
  assign n36996 = ~pi211 & n36995;
  assign n36997 = ~n36981 & ~n36996;
  assign n36998 = ~n36536 & n36997;
  assign n36999 = pi219 & ~n36536;
  assign n37000 = pi219 & ~n36980;
  assign n37001 = ~n36999 & ~n37000;
  assign n37002 = ~n36998 & ~n37001;
  assign n37003 = ~po1038 & ~n37002;
  assign n37004 = pi211 & ~n36995;
  assign n37005 = ~pi1153 & ~n36610;
  assign n37006 = pi1154 & ~n10957;
  assign n37007 = n36624 & ~n37006;
  assign n37008 = ~n37005 & ~n37007;
  assign n37009 = ~n36979 & n37008;
  assign n37010 = ~n36977 & ~n37009;
  assign n37011 = ~pi211 & ~n37010;
  assign n37012 = pi214 & ~n37011;
  assign n37013 = ~n37004 & n37012;
  assign n37014 = ~n36549 & ~n36980;
  assign n37015 = ~pi211 & ~n37014;
  assign n37016 = pi211 & ~n37010;
  assign n37017 = ~n37015 & ~n37016;
  assign n37018 = ~pi214 & n37017;
  assign n37019 = pi212 & ~n37013;
  assign n37020 = ~n37018 & n37019;
  assign n37021 = ~pi214 & ~n36980;
  assign n37022 = ~pi212 & ~n37021;
  assign n37023 = pi214 & n37017;
  assign n37024 = n37022 & ~n37023;
  assign n37025 = ~pi219 & ~n37020;
  assign n37026 = ~n37024 & n37025;
  assign n37027 = n37003 & ~n37026;
  assign n37028 = n36930 & ~n37027;
  assign n37029 = pi1154 & ~n10422;
  assign n37030 = ~n36987 & ~n37029;
  assign n37031 = n36514 & n37030;
  assign n37032 = n36660 & ~n37031;
  assign n37033 = n36659 & n37030;
  assign n37034 = pi1153 & ~n10422;
  assign n37035 = n36514 & ~n37034;
  assign n37036 = pi208 & ~n37035;
  assign n37037 = ~n37033 & n37036;
  assign n37038 = ~n37032 & ~n37037;
  assign n37039 = pi200 & pi207;
  assign n37040 = ~pi199 & ~n37039;
  assign n37041 = ~pi299 & ~n37040;
  assign n37042 = pi208 & ~n37041;
  assign n37043 = ~pi299 & n37042;
  assign n37044 = n10970 & n36522;
  assign n37045 = ~n37043 & ~n37044;
  assign n37046 = ~n37038 & ~n37045;
  assign n37047 = pi219 & ~n37046;
  assign n37048 = ~po1038 & ~n37047;
  assign n37049 = ~pi211 & n10332;
  assign n37050 = ~n37005 & ~n37038;
  assign n37051 = n37049 & ~n37050;
  assign n37052 = ~n36802 & ~n37038;
  assign n37053 = ~pi211 & ~n37052;
  assign n37054 = pi211 & ~n37050;
  assign n37055 = ~n37053 & ~n37054;
  assign n37056 = n36675 & ~n37055;
  assign n37057 = ~n37051 & ~n37056;
  assign n37058 = ~pi219 & ~n37057;
  assign n37059 = ~n36583 & ~n36675;
  assign n37060 = ~n37046 & n37059;
  assign n37061 = n37048 & ~n37060;
  assign n37062 = ~n37058 & n37061;
  assign n37063 = n36877 & ~n37062;
  assign n37064 = ~n37028 & ~n37063;
  assign n37065 = ~pi213 & ~n37064;
  assign n37066 = ~pi1152 & ~po1038;
  assign n37067 = n36536 & n37046;
  assign n37068 = pi299 & ~n36567;
  assign n37069 = ~n37046 & ~n37068;
  assign n37070 = n36675 & ~n37069;
  assign n37071 = ~pi211 & ~n36545;
  assign n37072 = ~n37046 & n37071;
  assign n37073 = pi211 & ~n37052;
  assign n37074 = n10332 & ~n37072;
  assign n37075 = ~n37073 & n37074;
  assign n37076 = ~n37070 & ~n37075;
  assign n37077 = ~pi219 & ~n37076;
  assign n37078 = pi211 & ~n37046;
  assign n37079 = n36999 & ~n37053;
  assign n37080 = ~n37078 & n37079;
  assign n37081 = ~n37067 & ~n37080;
  assign n37082 = ~n37077 & n37081;
  assign n37083 = n37066 & ~n37082;
  assign n37084 = ~n36536 & n37015;
  assign n37085 = ~n36980 & ~n37084;
  assign n37086 = pi219 & ~n37085;
  assign n37087 = ~pi212 & n37021;
  assign n37088 = ~n36825 & ~n36995;
  assign n37089 = ~pi211 & n37088;
  assign n37090 = pi211 & ~n37014;
  assign n37091 = n10332 & ~n37090;
  assign n37092 = ~n37089 & n37091;
  assign n37093 = pi211 & n37088;
  assign n37094 = ~pi208 & ~n36813;
  assign n37095 = ~n36980 & n37094;
  assign n37096 = pi299 & ~pi1156;
  assign n37097 = n36986 & ~n37096;
  assign n37098 = ~n36813 & n36971;
  assign n37099 = ~pi207 & ~n37098;
  assign n37100 = pi208 & ~n37097;
  assign n37101 = ~n37099 & n37100;
  assign n37102 = ~pi211 & ~n37095;
  assign n37103 = ~n37101 & n37102;
  assign n37104 = n36675 & ~n37093;
  assign n37105 = ~n37103 & n37104;
  assign n37106 = ~pi219 & ~n37087;
  assign n37107 = ~n37092 & n37106;
  assign n37108 = ~n37105 & n37107;
  assign n37109 = ~n37086 & ~n37108;
  assign n37110 = pi1152 & ~po1038;
  assign n37111 = ~n37109 & n37110;
  assign n37112 = pi213 & ~n37083;
  assign n37113 = ~n37111 & n37112;
  assign n37114 = ~pi209 & ~n37113;
  assign n37115 = ~n37065 & n37114;
  assign n37116 = pi219 & ~n36579;
  assign n37117 = n36544 & ~n36567;
  assign n37118 = ~pi219 & ~n37117;
  assign n37119 = ~n36570 & n37118;
  assign n37120 = pi213 & ~n37116;
  assign n37121 = n36921 & n37120;
  assign n37122 = ~n37119 & n37121;
  assign n37123 = ~n37115 & ~n37122;
  assign n37124 = ~n36966 & n37123;
  assign n37125 = pi230 & ~n37124;
  assign po391 = n36870 | n37125;
  assign n37127 = pi214 & n36567;
  assign n37128 = ~pi214 & n36559;
  assign n37129 = pi212 & ~n37127;
  assign n37130 = ~n37128 & n37129;
  assign n37131 = n36577 & ~n37130;
  assign n37132 = pi219 & ~n36675;
  assign n37133 = pi219 & ~n36561;
  assign n37134 = ~n37132 & ~n37133;
  assign n37135 = po1038 & n37134;
  assign n37136 = ~n37131 & n37135;
  assign n37137 = ~pi1156 & n36620;
  assign n37138 = ~n36747 & ~n37137;
  assign n37139 = pi207 & ~n37138;
  assign n37140 = ~pi207 & n36657;
  assign n37141 = ~n37139 & ~n37140;
  assign n37142 = pi208 & ~n37141;
  assign n37143 = ~n36808 & ~n37142;
  assign n37144 = n36780 & n36879;
  assign n37145 = n37143 & ~n37144;
  assign n37146 = ~pi299 & ~n37145;
  assign n37147 = ~n36545 & ~n37146;
  assign n37148 = ~pi211 & n37147;
  assign n37149 = ~pi299 & ~n36878;
  assign n37150 = ~n36597 & n37149;
  assign n37151 = ~n37143 & n37150;
  assign n37152 = ~pi1157 & ~n37151;
  assign n37153 = ~pi207 & n36725;
  assign n37154 = n10101 & ~n36716;
  assign n37155 = ~n37137 & n37154;
  assign n37156 = ~n37153 & ~n37155;
  assign n37157 = ~n36727 & n37156;
  assign n37158 = pi1157 & ~n37157;
  assign n37159 = ~n37152 & ~n37158;
  assign n37160 = pi211 & ~n37159;
  assign n37161 = n36675 & ~n37160;
  assign n37162 = ~n37148 & n37161;
  assign n37163 = ~n36675 & n37159;
  assign n37164 = pi219 & ~n37163;
  assign n37165 = ~n37162 & n37164;
  assign n37166 = pi211 & ~n37147;
  assign n37167 = ~pi211 & ~n37145;
  assign n37168 = n10332 & ~n37167;
  assign n37169 = ~n37166 & n37168;
  assign n37170 = n36536 & ~n37159;
  assign n37171 = pi211 & ~n37145;
  assign n37172 = ~pi299 & n37145;
  assign n37173 = pi1157 & n37172;
  assign n37174 = ~pi211 & ~n37152;
  assign n37175 = ~n37173 & n37174;
  assign n37176 = n36675 & ~n37171;
  assign n37177 = ~n37175 & n37176;
  assign n37178 = ~n37169 & ~n37170;
  assign n37179 = ~n37177 & n37178;
  assign n37180 = ~pi219 & ~n37179;
  assign n37181 = pi209 & ~n37165;
  assign n37182 = ~n37180 & n37181;
  assign n37183 = n36739 & n36775;
  assign n37184 = pi208 & ~n37031;
  assign n37185 = ~n36514 & ~n36739;
  assign n37186 = n37184 & ~n37185;
  assign n37187 = ~n37183 & ~n37186;
  assign n37188 = ~pi211 & n37187;
  assign n37189 = ~pi1154 & ~n36987;
  assign n37190 = pi200 & ~pi1153;
  assign n37191 = n10970 & ~n37190;
  assign n37192 = ~n37189 & n37191;
  assign n37193 = n10101 & ~n37192;
  assign n37194 = ~n36615 & ~n36878;
  assign n37195 = ~n10101 & ~n37194;
  assign n37196 = ~n37193 & ~n37195;
  assign n37197 = pi211 & ~n37196;
  assign n37198 = n36675 & ~n37197;
  assign n37199 = ~n37188 & n37198;
  assign n37200 = ~n36675 & n37196;
  assign n37201 = pi219 & ~n37200;
  assign n37202 = ~n37199 & n37201;
  assign n37203 = n36536 & ~n37196;
  assign n37204 = n36660 & ~n36832;
  assign n37205 = n36659 & n36831;
  assign n37206 = n37184 & ~n37205;
  assign n37207 = ~n37204 & ~n37206;
  assign n37208 = pi1157 & ~n37207;
  assign n37209 = ~pi1157 & n37196;
  assign n37210 = ~pi211 & ~n37208;
  assign n37211 = ~n37209 & n37210;
  assign n37212 = ~n36813 & ~n37196;
  assign n37213 = pi211 & n37212;
  assign n37214 = ~n37211 & ~n37213;
  assign n37215 = n36675 & ~n37214;
  assign n37216 = ~pi211 & ~n37212;
  assign n37217 = pi211 & ~n37187;
  assign n37218 = n10332 & ~n37217;
  assign n37219 = ~n37216 & n37218;
  assign n37220 = ~n37203 & ~n37219;
  assign n37221 = ~n37215 & n37220;
  assign n37222 = ~pi219 & ~n37221;
  assign n37223 = ~pi209 & ~n37202;
  assign n37224 = ~n37222 & n37223;
  assign n37225 = ~n37182 & ~n37224;
  assign n37226 = ~po1038 & ~n37225;
  assign n37227 = pi213 & ~n37136;
  assign n37228 = ~n37226 & n37227;
  assign n37229 = ~pi219 & po1038;
  assign n37230 = po1038 & n36581;
  assign n37231 = ~n37229 & ~n37230;
  assign n37232 = ~n36563 & n36675;
  assign n37233 = n10332 & ~n36872;
  assign n37234 = ~pi219 & ~n37232;
  assign n37235 = ~n37233 & n37234;
  assign n37236 = ~n37132 & ~n37235;
  assign n37237 = ~n37231 & n37236;
  assign n37238 = ~n36621 & ~n36827;
  assign n37239 = ~n36716 & ~n37238;
  assign n37240 = pi207 & ~n37239;
  assign n37241 = pi1154 & ~n36656;
  assign n37242 = ~n36708 & ~n37241;
  assign n37243 = ~pi207 & ~n36777;
  assign n37244 = ~n37242 & n37243;
  assign n37245 = ~n37240 & ~n37244;
  assign n37246 = pi208 & ~n37245;
  assign n37247 = ~n36801 & ~n37246;
  assign n37248 = ~pi1157 & ~n37247;
  assign n37249 = n36803 & ~n37172;
  assign n37250 = ~n37248 & ~n37249;
  assign n37251 = pi211 & n37250;
  assign n37252 = ~n37148 & ~n37251;
  assign n37253 = n36675 & ~n37252;
  assign n37254 = ~pi211 & ~n37250;
  assign n37255 = pi211 & ~n36847;
  assign n37256 = ~n37172 & n37255;
  assign n37257 = n10332 & ~n37256;
  assign n37258 = ~n37254 & n37257;
  assign n37259 = ~n37170 & ~n37258;
  assign n37260 = ~n37253 & n37259;
  assign n37261 = ~pi219 & ~n37260;
  assign n37262 = ~pi211 & ~n36547;
  assign n37263 = ~n37146 & n37262;
  assign n37264 = n37161 & ~n37263;
  assign n37265 = n37164 & ~n37264;
  assign n37266 = pi209 & ~n37265;
  assign n37267 = ~n37261 & n37266;
  assign n37268 = n36660 & ~n36796;
  assign n37269 = ~n36514 & n36796;
  assign n37270 = n37184 & ~n37269;
  assign n37271 = ~n37268 & ~n37270;
  assign n37272 = pi211 & n37271;
  assign n37273 = ~n37188 & ~n37272;
  assign n37274 = n36675 & ~n37273;
  assign n37275 = ~pi211 & ~n37271;
  assign n37276 = n36660 & ~n36831;
  assign n37277 = ~n36604 & n37206;
  assign n37278 = ~n37276 & ~n37277;
  assign n37279 = pi211 & ~n37278;
  assign n37280 = n10332 & ~n37279;
  assign n37281 = ~n37275 & n37280;
  assign n37282 = ~n37203 & ~n37281;
  assign n37283 = ~n37274 & n37282;
  assign n37284 = ~pi219 & ~n37283;
  assign n37285 = ~pi211 & n37278;
  assign n37286 = n37198 & ~n37285;
  assign n37287 = n37201 & ~n37286;
  assign n37288 = ~pi209 & ~n37287;
  assign n37289 = ~n37284 & n37288;
  assign n37290 = ~n37267 & ~n37289;
  assign n37291 = ~po1038 & ~n37290;
  assign n37292 = ~pi213 & ~n37237;
  assign n37293 = ~n37291 & n37292;
  assign n37294 = ~n37228 & ~n37293;
  assign n37295 = pi230 & ~n37294;
  assign n37296 = ~pi230 & ~pi235;
  assign po392 = ~n37295 & ~n37296;
  assign n37298 = ~pi100 & n36300;
  assign n37299 = n36489 & ~n37298;
  assign n37300 = ~n6079 & ~n37299;
  assign n37301 = ~pi75 & ~n37300;
  assign n37302 = ~n7229 & ~n37301;
  assign n37303 = ~pi92 & ~n37302;
  assign n37304 = n12909 & ~n37303;
  assign n37305 = ~pi74 & ~n37304;
  assign n37306 = n6077 & ~n37305;
  assign n37307 = ~pi56 & ~n37306;
  assign n37308 = ~n6248 & ~n37307;
  assign n37309 = ~pi62 & ~n37308;
  assign po393 = n12917 & ~n37309;
  assign n37311 = pi211 & pi1157;
  assign n37312 = ~pi211 & pi1158;
  assign n37313 = ~n37311 & ~n37312;
  assign n37314 = n36544 & ~n37313;
  assign n37315 = ~pi219 & ~n37314;
  assign n37316 = ~n37130 & n37315;
  assign n37317 = n36544 & n36565;
  assign n37318 = po1038 & n37317;
  assign n37319 = ~n37229 & ~n37318;
  assign n37320 = ~pi214 & n36561;
  assign n37321 = pi1154 & n36583;
  assign n37322 = ~n37320 & ~n37321;
  assign n37323 = pi212 & ~n37322;
  assign n37324 = po1038 & n37323;
  assign n37325 = n37319 & ~n37324;
  assign n37326 = ~n37316 & ~n37325;
  assign n37327 = ~pi213 & ~n37326;
  assign n37328 = n36572 & ~n37316;
  assign n37329 = pi199 & pi1143;
  assign n37330 = ~pi200 & ~n37329;
  assign n37331 = ~n36507 & n37330;
  assign n37332 = ~n36510 & n36972;
  assign n37333 = ~n37331 & n37332;
  assign n37334 = pi200 & ~n36507;
  assign n37335 = ~pi199 & pi1145;
  assign n37336 = n37330 & ~n37335;
  assign n37337 = n36879 & ~n37334;
  assign n37338 = ~n37336 & n37337;
  assign n37339 = ~n37333 & ~n37338;
  assign n37340 = ~pi299 & ~n37339;
  assign n37341 = n36544 & n36813;
  assign n37342 = pi214 & ~n36549;
  assign n37343 = ~pi214 & ~n36545;
  assign n37344 = pi212 & ~n37342;
  assign n37345 = ~n37343 & n37344;
  assign n37346 = ~n37341 & ~n37345;
  assign n37347 = n36554 & ~n37346;
  assign n37348 = ~n37340 & ~n37347;
  assign n37349 = ~n37328 & n37348;
  assign n37350 = ~po1038 & ~n37349;
  assign n37351 = n37327 & ~n37350;
  assign n37352 = pi299 & ~n36536;
  assign n37353 = pi219 & ~n36530;
  assign n37354 = ~pi211 & pi1145;
  assign n37355 = pi211 & pi1144;
  assign n37356 = ~n37354 & ~n37355;
  assign n37357 = ~n10332 & n37356;
  assign n37358 = n10332 & n36528;
  assign n37359 = ~n36536 & ~n37357;
  assign n37360 = ~n37358 & n37359;
  assign n37361 = ~pi219 & ~n37360;
  assign n37362 = n37352 & ~n37353;
  assign n37363 = ~n37361 & n37362;
  assign n37364 = ~n37340 & ~n37363;
  assign n37365 = ~po1038 & ~n37364;
  assign n37366 = n36921 & ~n37353;
  assign n37367 = ~n37361 & n37366;
  assign n37368 = ~n37365 & ~n37367;
  assign n37369 = pi213 & n37368;
  assign n37370 = pi209 & ~n37351;
  assign n37371 = ~n37369 & n37370;
  assign n37372 = ~pi200 & pi207;
  assign n37373 = ~pi200 & ~pi1158;
  assign n37374 = ~pi199 & ~n37373;
  assign n37375 = ~pi1156 & ~n12341;
  assign n37376 = pi1158 & ~n37375;
  assign n37377 = pi199 & pi1156;
  assign n37378 = ~n37376 & ~n37377;
  assign n37379 = n37372 & ~n37378;
  assign n37380 = ~n37374 & ~n37379;
  assign n37381 = n36514 & ~n37380;
  assign n37382 = ~pi208 & n37381;
  assign n37383 = n37372 & n37382;
  assign n37384 = pi207 & n36717;
  assign n37385 = ~pi207 & ~n36709;
  assign n37386 = pi208 & ~n37384;
  assign n37387 = ~n37385 & n37386;
  assign n37388 = ~n37383 & ~n37387;
  assign n37389 = ~pi1157 & ~n37388;
  assign n37390 = ~pi200 & n37377;
  assign n37391 = ~n37374 & ~n37390;
  assign n37392 = n36514 & ~n37391;
  assign n37393 = ~pi208 & ~n37392;
  assign n37394 = ~n37153 & ~n37384;
  assign n37395 = pi208 & ~n37394;
  assign n37396 = pi1157 & ~n37393;
  assign n37397 = ~n37395 & n37396;
  assign n37398 = ~n37389 & ~n37397;
  assign n37399 = ~n36731 & n37398;
  assign n37400 = ~pi1157 & ~n37383;
  assign n37401 = n37382 & ~n37400;
  assign n37402 = ~pi208 & ~n37401;
  assign n37403 = ~n36596 & n37402;
  assign n37404 = n36658 & ~n36780;
  assign n37405 = ~pi207 & ~n36626;
  assign n37406 = ~n37404 & n37405;
  assign n37407 = pi207 & ~n36647;
  assign n37408 = pi208 & ~n37406;
  assign n37409 = ~n37407 & n37408;
  assign n37410 = ~n37403 & ~n37409;
  assign n37411 = n36731 & ~n37410;
  assign n37412 = ~n37399 & ~n37411;
  assign n37413 = pi219 & ~n37412;
  assign n37414 = ~pi214 & n37398;
  assign n37415 = ~pi212 & ~n37414;
  assign n37416 = ~n36683 & n37402;
  assign n37417 = ~pi207 & ~n36680;
  assign n37418 = ~n37404 & n37417;
  assign n37419 = pi207 & ~n36696;
  assign n37420 = pi208 & ~n37418;
  assign n37421 = ~n37419 & n37420;
  assign n37422 = ~n37416 & ~n37421;
  assign n37423 = pi211 & ~n37422;
  assign n37424 = pi299 & pi1145;
  assign n37425 = n37402 & ~n37424;
  assign n37426 = ~pi299 & ~n36809;
  assign n37427 = ~n37424 & ~n37426;
  assign n37428 = pi207 & ~n37427;
  assign n37429 = pi299 & ~pi1145;
  assign n37430 = ~pi207 & ~n37429;
  assign n37431 = ~n37404 & n37430;
  assign n37432 = pi208 & ~n37431;
  assign n37433 = ~n37428 & n37432;
  assign n37434 = ~n37425 & ~n37433;
  assign n37435 = ~pi211 & ~n37434;
  assign n37436 = ~n37423 & ~n37435;
  assign n37437 = pi214 & ~n37436;
  assign n37438 = n37415 & ~n37437;
  assign n37439 = ~pi211 & n37422;
  assign n37440 = pi211 & n37410;
  assign n37441 = pi214 & ~n37439;
  assign n37442 = ~n37440 & n37441;
  assign n37443 = ~pi214 & ~n37436;
  assign n37444 = pi212 & ~n37442;
  assign n37445 = ~n37443 & n37444;
  assign n37446 = ~pi219 & ~n37438;
  assign n37447 = ~n37445 & n37446;
  assign n37448 = ~po1038 & ~n37413;
  assign n37449 = ~n37447 & n37448;
  assign n37450 = pi213 & ~n37367;
  assign n37451 = ~n37449 & n37450;
  assign n37452 = pi208 & pi1157;
  assign n37453 = pi207 & ~n36809;
  assign n37454 = ~n36724 & ~n36760;
  assign n37455 = ~pi207 & ~n37454;
  assign n37456 = ~n37453 & ~n37455;
  assign n37457 = n37452 & ~n37456;
  assign n37458 = ~n36813 & ~n37392;
  assign n37459 = n36663 & ~n37458;
  assign n37460 = n37094 & ~n37379;
  assign n37461 = pi208 & ~n37140;
  assign n37462 = ~n37453 & n37461;
  assign n37463 = ~pi1157 & ~n37460;
  assign n37464 = ~n37462 & n37463;
  assign n37465 = ~n37457 & ~n37459;
  assign n37466 = ~n37464 & n37465;
  assign n37467 = n36544 & n37466;
  assign n37468 = ~n36545 & ~n37381;
  assign n37469 = n36663 & ~n37468;
  assign n37470 = ~pi207 & n36779;
  assign n37471 = pi207 & ~n36784;
  assign n37472 = ~n37470 & ~n37471;
  assign n37473 = pi208 & ~n37472;
  assign n37474 = ~pi299 & ~n37372;
  assign n37475 = ~pi208 & ~n37474;
  assign n37476 = ~n37468 & n37475;
  assign n37477 = ~n37473 & ~n37476;
  assign n37478 = ~pi1157 & ~n37477;
  assign n37479 = ~n10970 & ~n36664;
  assign n37480 = pi1156 & ~n37479;
  assign n37481 = ~pi1156 & ~n36619;
  assign n37482 = ~n36744 & n37481;
  assign n37483 = ~n37480 & ~n37482;
  assign n37484 = ~pi207 & ~n37483;
  assign n37485 = ~n37471 & ~n37484;
  assign n37486 = n37452 & ~n37485;
  assign n37487 = ~n37469 & ~n37486;
  assign n37488 = ~n37478 & n37487;
  assign n37489 = ~pi214 & ~n37488;
  assign n37490 = ~n36549 & n37402;
  assign n37491 = ~pi207 & ~n36761;
  assign n37492 = ~n36802 & n37491;
  assign n37493 = pi1157 & ~n37492;
  assign n37494 = ~n37244 & n37400;
  assign n37495 = ~n37493 & ~n37494;
  assign n37496 = pi208 & ~n36888;
  assign n37497 = ~n37495 & n37496;
  assign n37498 = pi214 & ~n37490;
  assign n37499 = ~n37497 & n37498;
  assign n37500 = pi212 & ~n37489;
  assign n37501 = ~n37499 & n37500;
  assign n37502 = ~n37467 & ~n37501;
  assign n37503 = ~pi211 & ~n37502;
  assign n37504 = ~n37399 & ~n37503;
  assign n37505 = pi219 & ~n37504;
  assign n37506 = n36790 & ~n37466;
  assign n37507 = n10098 & ~n37488;
  assign n37508 = ~pi299 & n37391;
  assign n37509 = n36660 & ~n37508;
  assign n37510 = ~pi207 & n36761;
  assign n37511 = pi208 & ~n37510;
  assign n37512 = ~n36896 & n37511;
  assign n37513 = ~n37509 & ~n37512;
  assign n37514 = pi1157 & ~n37513;
  assign n37515 = ~n37389 & ~n37514;
  assign n37516 = n36789 & ~n37515;
  assign n37517 = ~n37506 & ~n37507;
  assign n37518 = ~n37516 & n37517;
  assign n37519 = pi212 & ~n37518;
  assign n37520 = pi211 & n37515;
  assign n37521 = ~pi1158 & n36717;
  assign n37522 = pi1158 & n36828;
  assign n37523 = pi207 & ~n37521;
  assign n37524 = ~n37522 & n37523;
  assign n37525 = pi299 & ~pi1158;
  assign n37526 = n37491 & ~n37525;
  assign n37527 = ~n37524 & ~n37526;
  assign n37528 = n37452 & ~n37527;
  assign n37529 = pi207 & ~n10422;
  assign n37530 = ~pi299 & ~n37529;
  assign n37531 = pi1158 & ~n37530;
  assign n37532 = pi1157 & n37381;
  assign n37533 = ~n37531 & ~n37532;
  assign n37534 = ~pi208 & ~n37533;
  assign n37535 = ~pi207 & ~n37525;
  assign n37536 = ~n36658 & n37535;
  assign n37537 = ~n37524 & ~n37536;
  assign n37538 = pi208 & ~n37537;
  assign n37539 = ~n37383 & ~n37538;
  assign n37540 = ~pi1157 & ~n37539;
  assign n37541 = ~pi211 & ~n37534;
  assign n37542 = ~n37528 & n37541;
  assign n37543 = ~n37540 & n37542;
  assign n37544 = ~n37520 & ~n37543;
  assign n37545 = pi214 & ~n37544;
  assign n37546 = n37415 & ~n37545;
  assign n37547 = ~pi219 & ~n37519;
  assign n37548 = ~n37546 & n37547;
  assign n37549 = ~po1038 & ~n37548;
  assign n37550 = ~n37505 & n37549;
  assign n37551 = n37327 & ~n37550;
  assign n37552 = ~pi209 & ~n37451;
  assign n37553 = ~n37551 & n37552;
  assign n37554 = ~n37371 & ~n37553;
  assign n37555 = pi230 & ~n37554;
  assign n37556 = ~pi230 & ~pi237;
  assign po394 = n37555 | n37556;
  assign n37558 = ~pi230 & pi238;
  assign n37559 = n36522 & n36983;
  assign n37560 = ~n10101 & n36982;
  assign n37561 = n37043 & ~n37560;
  assign n37562 = ~pi299 & ~n37559;
  assign n37563 = ~n37561 & n37562;
  assign n37564 = ~pi211 & ~n36802;
  assign n37565 = ~n37563 & n37564;
  assign n37566 = n10421 & n36879;
  assign n37567 = ~pi299 & ~n37566;
  assign n37568 = pi1153 & ~n37567;
  assign n37569 = ~n36879 & ~n37529;
  assign n37570 = ~n10101 & n36654;
  assign n37571 = ~n37569 & ~n37570;
  assign n37572 = n37567 & n37571;
  assign n37573 = ~n37568 & ~n37572;
  assign n37574 = pi211 & ~n37573;
  assign n37575 = ~n37565 & ~n37574;
  assign n37576 = n10332 & ~n37575;
  assign n37577 = n36675 & ~n37563;
  assign n37578 = pi299 & n36563;
  assign n37579 = n37577 & ~n37578;
  assign n37580 = ~n37576 & ~n37579;
  assign n37581 = ~pi219 & ~n37580;
  assign n37582 = ~n37045 & ~n37560;
  assign n37583 = n36581 & n37352;
  assign n37584 = ~n37582 & ~n37583;
  assign n37585 = ~n36732 & ~n37584;
  assign n37586 = ~n37581 & ~n37585;
  assign n37587 = ~pi1151 & ~po1038;
  assign n37588 = ~n37586 & n37587;
  assign n37589 = ~n36878 & ~n36985;
  assign n37590 = n37563 & ~n37589;
  assign n37591 = ~pi211 & ~n37590;
  assign n37592 = ~n36825 & n37591;
  assign n37593 = pi211 & ~n37590;
  assign n37594 = ~n36802 & n37593;
  assign n37595 = ~n37592 & ~n37594;
  assign n37596 = n36675 & ~n37595;
  assign n37597 = n37150 & ~n37566;
  assign n37598 = n12341 & n36879;
  assign n37599 = pi1153 & n37598;
  assign n37600 = ~n37597 & ~n37599;
  assign n37601 = n36536 & ~n37600;
  assign n37602 = n36871 & ~n37567;
  assign n37603 = ~n37597 & ~n37602;
  assign n37604 = ~n37565 & n37603;
  assign n37605 = n10332 & ~n37604;
  assign n37606 = ~pi219 & ~n37601;
  assign n37607 = ~n37605 & n37606;
  assign n37608 = ~n37596 & n37607;
  assign n37609 = pi211 & pi299;
  assign n37610 = ~pi214 & ~n37598;
  assign n37611 = ~pi212 & n37610;
  assign n37612 = ~n37567 & ~n37609;
  assign n37613 = ~n37611 & n37612;
  assign n37614 = pi1153 & n37613;
  assign n37615 = pi219 & ~n37597;
  assign n37616 = ~n37614 & n37615;
  assign n37617 = pi1151 & ~po1038;
  assign n37618 = ~n37616 & n37617;
  assign n37619 = ~n37608 & n37618;
  assign n37620 = pi1152 & ~n37588;
  assign n37621 = ~n37619 & n37620;
  assign n37622 = ~n36732 & ~n37614;
  assign n37623 = ~n36549 & ~n37599;
  assign n37624 = ~pi211 & ~n37623;
  assign n37625 = n10332 & ~n37602;
  assign n37626 = ~n37624 & n37625;
  assign n37627 = pi299 & ~n36563;
  assign n37628 = n36675 & ~n37627;
  assign n37629 = ~n37599 & n37628;
  assign n37630 = ~n37626 & ~n37629;
  assign n37631 = ~pi219 & ~n37630;
  assign n37632 = n37587 & ~n37622;
  assign n37633 = ~n37631 & n37632;
  assign n37634 = n36610 & n36879;
  assign n37635 = n36603 & n36972;
  assign n37636 = ~n37634 & ~n37635;
  assign n37637 = ~pi214 & n37636;
  assign n37638 = ~pi212 & ~n37637;
  assign n37639 = ~pi1153 & n10421;
  assign n37640 = ~n37636 & ~n37639;
  assign n37641 = ~n37627 & ~n37640;
  assign n37642 = n37638 & ~n37641;
  assign n37643 = pi207 & n36624;
  assign n37644 = pi200 & n36659;
  assign n37645 = pi208 & ~n37644;
  assign n37646 = ~n37643 & n37645;
  assign n37647 = ~n37475 & ~n37646;
  assign n37648 = ~n36975 & ~n37647;
  assign n37649 = n10098 & ~n37648;
  assign n37650 = ~n36549 & n36790;
  assign n37651 = ~n36545 & n36789;
  assign n37652 = ~n37650 & ~n37651;
  assign n37653 = ~n37640 & ~n37652;
  assign n37654 = pi212 & ~n37653;
  assign n37655 = ~n37649 & n37654;
  assign n37656 = ~pi219 & ~n37642;
  assign n37657 = ~n37655 & n37656;
  assign n37658 = ~n37583 & ~n37640;
  assign n37659 = pi219 & n37658;
  assign n37660 = n37617 & ~n37659;
  assign n37661 = ~n37657 & n37660;
  assign n37662 = ~pi1152 & ~n37633;
  assign n37663 = ~n37661 & n37662;
  assign n37664 = ~pi209 & ~n37663;
  assign n37665 = ~n37621 & n37664;
  assign n37666 = ~pi1153 & n36554;
  assign n37667 = n36921 & ~n37666;
  assign n37668 = ~n37235 & n37667;
  assign n37669 = pi1153 & ~pi1154;
  assign n37670 = n36707 & n37669;
  assign n37671 = n10101 & ~n37670;
  assign n37672 = ~n36968 & n37671;
  assign n37673 = ~n37195 & ~n37672;
  assign n37674 = n36536 & ~n37673;
  assign n37675 = pi211 & n37673;
  assign n37676 = pi1153 & ~n36624;
  assign n37677 = n36514 & ~n37676;
  assign n37678 = ~n36968 & n37677;
  assign n37679 = pi208 & ~n37678;
  assign n37680 = ~n36604 & ~n37205;
  assign n37681 = n37679 & n37680;
  assign n37682 = ~n37276 & ~n37681;
  assign n37683 = ~pi211 & ~n37682;
  assign n37684 = ~n37675 & ~n37683;
  assign n37685 = n36999 & n37684;
  assign n37686 = ~po1038 & ~n37674;
  assign n37687 = ~n37685 & n37686;
  assign n37688 = ~n37185 & n37679;
  assign n37689 = ~n37183 & ~n37688;
  assign n37690 = ~pi211 & ~n37689;
  assign n37691 = ~n37269 & n37679;
  assign n37692 = ~n37268 & ~n37691;
  assign n37693 = pi211 & ~n37692;
  assign n37694 = n36544 & ~n37690;
  assign n37695 = ~n37693 & n37694;
  assign n37696 = n36789 & ~n37689;
  assign n37697 = pi211 & ~pi214;
  assign n37698 = ~n36583 & ~n37697;
  assign n37699 = ~n37692 & ~n37698;
  assign n37700 = n10098 & ~n37682;
  assign n37701 = pi212 & ~n37696;
  assign n37702 = ~n37700 & n37701;
  assign n37703 = ~n37699 & n37702;
  assign n37704 = ~n37695 & ~n37703;
  assign n37705 = ~pi219 & ~n37704;
  assign n37706 = pi209 & n37687;
  assign n37707 = ~n37705 & n37706;
  assign n37708 = ~n37668 & ~n37707;
  assign n37709 = ~n37665 & n37708;
  assign n37710 = pi213 & ~n37709;
  assign n37711 = ~n10099 & n36732;
  assign n37712 = po1038 & n37711;
  assign n37713 = ~pi211 & ~pi1153;
  assign n37714 = ~n10332 & ~n37713;
  assign n37715 = ~n37049 & ~n37714;
  assign n37716 = n37712 & ~n37715;
  assign n37717 = ~pi1151 & ~n37716;
  assign n37718 = pi219 & ~n37582;
  assign n37719 = ~po1038 & ~n37718;
  assign n37720 = pi299 & n37049;
  assign n37721 = ~pi211 & n37573;
  assign n37722 = n37577 & ~n37721;
  assign n37723 = ~n36675 & n37582;
  assign n37724 = ~pi219 & ~n37720;
  assign n37725 = ~n37723 & n37724;
  assign n37726 = ~n37722 & n37725;
  assign n37727 = n37719 & ~n37726;
  assign n37728 = n37717 & ~n37727;
  assign n37729 = ~n10100 & n36921;
  assign n37730 = pi1151 & ~n37729;
  assign n37731 = ~n37716 & n37730;
  assign n37732 = ~n37591 & n37600;
  assign n37733 = pi214 & n37732;
  assign n37734 = ~pi214 & ~n37597;
  assign n37735 = ~n37599 & n37734;
  assign n37736 = ~n37733 & ~n37735;
  assign n37737 = ~pi212 & ~n37736;
  assign n37738 = ~n37732 & ~n37737;
  assign n37739 = pi219 & ~n37738;
  assign n37740 = ~po1038 & ~n37739;
  assign n37741 = ~pi212 & ~n37735;
  assign n37742 = ~n37568 & ~n37593;
  assign n37743 = pi214 & ~n37597;
  assign n37744 = n37742 & n37743;
  assign n37745 = n37741 & ~n37744;
  assign n37746 = n37734 & n37742;
  assign n37747 = pi214 & n37590;
  assign n37748 = pi212 & ~n37747;
  assign n37749 = ~n37746 & n37748;
  assign n37750 = ~pi219 & ~n37745;
  assign n37751 = ~n37749 & n37750;
  assign n37752 = n37740 & ~n37751;
  assign n37753 = n37731 & ~n37752;
  assign n37754 = ~n37728 & ~n37753;
  assign n37755 = pi1152 & ~n37754;
  assign n37756 = ~pi219 & n36675;
  assign n37757 = n37230 & n37756;
  assign n37758 = n37730 & ~n37757;
  assign n37759 = n12342 & ~n36536;
  assign n37760 = ~pi212 & ~n37759;
  assign n37761 = ~n37640 & n37760;
  assign n37762 = ~pi214 & ~n12342;
  assign n37763 = ~n37599 & ~n37609;
  assign n37764 = pi214 & n37763;
  assign n37765 = ~n37762 & ~n37764;
  assign n37766 = pi212 & ~n37640;
  assign n37767 = ~n37765 & n37766;
  assign n37768 = ~n37761 & ~n37767;
  assign n37769 = ~n10422 & n37713;
  assign n37770 = n37768 & ~n37769;
  assign n37771 = ~pi219 & ~n37770;
  assign n37772 = pi219 & ~n37759;
  assign n37773 = ~n37640 & n37772;
  assign n37774 = ~po1038 & ~n37773;
  assign n37775 = ~n37771 & n37774;
  assign n37776 = n37758 & ~n37775;
  assign n37777 = ~pi1151 & ~n37757;
  assign n37778 = pi219 & ~n37598;
  assign n37779 = ~po1038 & ~n37778;
  assign n37780 = n37613 & n37779;
  assign n37781 = ~pi211 & n37610;
  assign n37782 = pi212 & ~n37567;
  assign n37783 = ~n37781 & n37782;
  assign n37784 = n37583 & ~n37783;
  assign n37785 = ~pi214 & n37609;
  assign n37786 = pi212 & ~n37785;
  assign n37787 = ~n37763 & n37786;
  assign n37788 = ~pi219 & ~n37787;
  assign n37789 = ~n37598 & ~n37784;
  assign n37790 = n37788 & n37789;
  assign n37791 = pi1153 & n37780;
  assign n37792 = ~n37790 & n37791;
  assign n37793 = n37777 & ~n37792;
  assign n37794 = ~n37776 & ~n37793;
  assign n37795 = ~pi1152 & ~n37794;
  assign n37796 = ~n37755 & ~n37795;
  assign n37797 = ~pi209 & ~n37796;
  assign n37798 = ~pi214 & ~n37673;
  assign n37799 = pi214 & n37684;
  assign n37800 = ~n37798 & ~n37799;
  assign n37801 = ~pi212 & ~n37800;
  assign n37802 = ~pi214 & ~n37684;
  assign n37803 = ~pi299 & n37682;
  assign n37804 = pi211 & ~n37803;
  assign n37805 = ~pi211 & n37673;
  assign n37806 = ~n37804 & ~n37805;
  assign n37807 = pi214 & ~n37806;
  assign n37808 = pi212 & ~n37802;
  assign n37809 = ~n37807 & n37808;
  assign n37810 = ~n37801 & ~n37809;
  assign n37811 = ~pi219 & ~n37810;
  assign n37812 = ~po1038 & ~n37772;
  assign n37813 = ~n37687 & ~n37812;
  assign n37814 = ~n37811 & ~n37813;
  assign n37815 = n37758 & ~n37814;
  assign n37816 = ~n37673 & ~n37756;
  assign n37817 = n37684 & n37756;
  assign n37818 = ~po1038 & ~n37816;
  assign n37819 = ~n37817 & n37818;
  assign n37820 = n37777 & ~n37819;
  assign n37821 = ~n37815 & ~n37820;
  assign n37822 = ~pi1152 & ~n37821;
  assign n37823 = ~n37609 & n37682;
  assign n37824 = pi214 & n37823;
  assign n37825 = ~pi212 & ~n37798;
  assign n37826 = ~n37824 & n37825;
  assign n37827 = ~pi219 & ~n37826;
  assign n37828 = pi214 & pi299;
  assign n37829 = ~n37785 & ~n37828;
  assign n37830 = n37682 & n37829;
  assign n37831 = pi212 & ~n37830;
  assign n37832 = n37827 & ~n37831;
  assign n37833 = ~n37813 & ~n37832;
  assign n37834 = n37731 & ~n37833;
  assign n37835 = pi219 & ~n37673;
  assign n37836 = ~pi214 & n37823;
  assign n37837 = ~n12342 & n37799;
  assign n37838 = pi212 & ~n37836;
  assign n37839 = ~n37837 & n37838;
  assign n37840 = n37827 & ~n37839;
  assign n37841 = ~po1038 & ~n37835;
  assign n37842 = ~n37840 & n37841;
  assign n37843 = n37717 & ~n37842;
  assign n37844 = ~n37834 & ~n37843;
  assign n37845 = pi1152 & ~n37844;
  assign n37846 = ~n37822 & ~n37845;
  assign n37847 = pi209 & ~n37846;
  assign n37848 = ~pi213 & ~n37797;
  assign n37849 = ~n37847 & n37848;
  assign n37850 = ~n37710 & ~n37849;
  assign n37851 = pi230 & ~n37850;
  assign po395 = n37558 | n37851;
  assign n37853 = po1038 & ~n37116;
  assign n37854 = n36544 & ~n37118;
  assign n37855 = n37853 & n37854;
  assign n37856 = n36522 & ~n36717;
  assign n37857 = pi212 & ~n37856;
  assign n37858 = ~po1038 & ~n37857;
  assign n37859 = ~pi214 & n37856;
  assign n37860 = ~pi212 & ~n37859;
  assign n37861 = pi219 & n37860;
  assign n37862 = pi211 & ~n37856;
  assign n37863 = pi214 & ~n37862;
  assign n37864 = ~n36549 & ~n36890;
  assign n37865 = n37863 & ~n37864;
  assign n37866 = n37861 & ~n37865;
  assign n37867 = ~pi219 & n37860;
  assign n37868 = ~pi211 & ~n36813;
  assign n37869 = ~n36946 & n37868;
  assign n37870 = ~n36545 & n37862;
  assign n37871 = pi214 & ~n37869;
  assign n37872 = ~n37870 & n37871;
  assign n37873 = n37867 & ~n37872;
  assign n37874 = n37858 & ~n37873;
  assign n37875 = ~n37866 & n37874;
  assign n37876 = ~pi209 & ~n37875;
  assign n37877 = pi212 & ~n37401;
  assign n37878 = ~po1038 & ~n37877;
  assign n37879 = ~pi214 & n37401;
  assign n37880 = ~pi212 & ~n37879;
  assign n37881 = ~pi219 & n37880;
  assign n37882 = ~n37068 & ~n37401;
  assign n37883 = pi214 & ~n37882;
  assign n37884 = n37881 & ~n37883;
  assign n37885 = ~pi211 & n37828;
  assign n37886 = pi1154 & n37885;
  assign n37887 = ~pi212 & pi219;
  assign n37888 = ~n37886 & n37887;
  assign n37889 = ~n37401 & n37888;
  assign n37890 = n37878 & ~n37889;
  assign n37891 = ~n37884 & n37890;
  assign n37892 = pi209 & ~n37891;
  assign n37893 = ~n37876 & ~n37892;
  assign n37894 = ~pi213 & ~n37855;
  assign n37895 = ~n37893 & n37894;
  assign n37896 = ~n37315 & ~n37319;
  assign n37897 = pi1157 & ~n36895;
  assign n37898 = ~n37509 & n37897;
  assign n37899 = ~n37400 & ~n37898;
  assign n37900 = pi211 & ~n37899;
  assign n37901 = pi299 & pi1158;
  assign n37902 = ~pi211 & ~n37901;
  assign n37903 = ~n37401 & n37902;
  assign n37904 = pi214 & ~n37900;
  assign n37905 = ~n37903 & n37904;
  assign n37906 = n37881 & ~n37905;
  assign n37907 = ~pi211 & ~n37868;
  assign n37908 = ~n37401 & ~n37907;
  assign n37909 = pi214 & ~n37908;
  assign n37910 = pi219 & n37880;
  assign n37911 = ~n37909 & n37910;
  assign n37912 = pi209 & n37878;
  assign n37913 = ~n37906 & n37912;
  assign n37914 = ~n37911 & n37913;
  assign n37915 = n37863 & ~n37869;
  assign n37916 = n37861 & ~n37915;
  assign n37917 = ~n36522 & n37901;
  assign n37918 = ~pi208 & n37524;
  assign n37919 = ~n37917 & ~n37918;
  assign n37920 = ~pi211 & ~n37919;
  assign n37921 = ~pi1157 & ~n37856;
  assign n37922 = ~n36897 & n37897;
  assign n37923 = pi211 & ~n37921;
  assign n37924 = ~n37922 & n37923;
  assign n37925 = ~n37920 & ~n37924;
  assign n37926 = pi214 & ~n37925;
  assign n37927 = n37867 & ~n37926;
  assign n37928 = ~pi209 & n37858;
  assign n37929 = ~n37916 & n37928;
  assign n37930 = ~n37927 & n37929;
  assign n37931 = pi213 & ~n37896;
  assign n37932 = ~n37930 & n37931;
  assign n37933 = ~n37914 & n37932;
  assign n37934 = ~n37895 & ~n37933;
  assign n37935 = pi230 & ~n37934;
  assign n37936 = ~pi230 & ~pi239;
  assign po396 = ~n37935 & ~n37936;
  assign n37938 = ~pi211 & pi1146;
  assign n37939 = pi211 & pi1145;
  assign n37940 = ~n37938 & ~n37939;
  assign n37941 = pi214 & ~n37940;
  assign n37942 = pi1146 & n37697;
  assign n37943 = ~n37941 & ~n37942;
  assign n37944 = pi212 & ~n37943;
  assign n37945 = pi211 & pi1146;
  assign n37946 = n36544 & n37945;
  assign n37947 = ~n37944 & ~n37946;
  assign n37948 = ~n36999 & n37947;
  assign n37949 = po1038 & n37354;
  assign n37950 = ~n37229 & ~n37949;
  assign n37951 = ~n37948 & ~n37950;
  assign n37952 = ~pi1147 & ~n37951;
  assign n37953 = ~pi199 & pi1146;
  assign n37954 = pi200 & ~n37953;
  assign n37955 = ~pi299 & ~n37954;
  assign n37956 = pi199 & pi1145;
  assign n37957 = n36628 & ~n37956;
  assign n37958 = n37955 & ~n37957;
  assign n37959 = ~n10101 & ~n37958;
  assign n37960 = ~pi200 & ~n37956;
  assign n37961 = ~n37953 & n37960;
  assign n37962 = pi200 & ~n37335;
  assign n37963 = n36514 & ~n37962;
  assign n37964 = ~n37961 & n37963;
  assign n37965 = ~n36879 & ~n37964;
  assign n37966 = ~n37959 & ~n37965;
  assign n37967 = pi299 & pi1146;
  assign n37968 = ~n37966 & ~n37967;
  assign n37969 = n36659 & n37960;
  assign n37970 = pi208 & ~n37969;
  assign n37971 = ~n37968 & n37970;
  assign n37972 = n36522 & ~n37960;
  assign n37973 = n37955 & n37972;
  assign n37974 = ~n37971 & ~n37973;
  assign n37975 = n37966 & ~n37974;
  assign n37976 = ~n36732 & ~n37975;
  assign n37977 = ~po1038 & ~n37976;
  assign n37978 = ~pi211 & n37424;
  assign n37979 = n36999 & n37978;
  assign n37980 = pi219 & ~n37979;
  assign n37981 = ~po1038 & ~n37980;
  assign n37982 = ~n37977 & ~n37981;
  assign n37983 = pi211 & n37967;
  assign n37984 = ~n37975 & ~n37983;
  assign n37985 = ~pi214 & ~n37975;
  assign n37986 = ~pi212 & ~n37985;
  assign n37987 = ~n37984 & n37986;
  assign n37988 = pi299 & ~n37943;
  assign n37989 = ~n37975 & ~n37988;
  assign n37990 = pi212 & ~n37989;
  assign n37991 = ~pi219 & ~n37990;
  assign n37992 = ~n37987 & n37991;
  assign n37993 = ~n37982 & ~n37992;
  assign n37994 = n37952 & ~n37993;
  assign n37995 = ~n37966 & n37980;
  assign n37996 = ~po1038 & ~n37995;
  assign n37997 = ~n12342 & ~n37966;
  assign n37998 = ~pi214 & ~n37966;
  assign n37999 = ~pi212 & ~n37998;
  assign n38000 = ~n37997 & n37999;
  assign n38001 = pi214 & ~n37983;
  assign n38002 = ~n37762 & ~n38001;
  assign n38003 = ~pi299 & ~n37966;
  assign n38004 = pi211 & ~n38003;
  assign n38005 = pi214 & n38004;
  assign n38006 = ~n37966 & ~n38002;
  assign n38007 = ~n38005 & n38006;
  assign n38008 = pi212 & ~n38007;
  assign n38009 = ~pi219 & ~n38000;
  assign n38010 = ~n38008 & n38009;
  assign n38011 = ~n37997 & ~n38010;
  assign n38012 = n37992 & ~n38011;
  assign n38013 = n37996 & ~n38012;
  assign n38014 = ~pi211 & n37229;
  assign n38015 = n36675 & n38014;
  assign n38016 = pi1147 & ~n38015;
  assign n38017 = ~n37951 & n38016;
  assign n38018 = ~n38013 & n38017;
  assign n38019 = ~n37994 & ~n38018;
  assign n38020 = ~pi213 & n38019;
  assign n38021 = ~n37812 & ~n37996;
  assign n38022 = pi299 & n10098;
  assign n38023 = ~pi299 & n37974;
  assign n38024 = pi214 & ~n38023;
  assign n38025 = ~n38004 & ~n38024;
  assign n38026 = pi212 & ~n38025;
  assign n38027 = ~pi219 & ~n37966;
  assign n38028 = ~n38022 & n38027;
  assign n38029 = ~n38026 & n38028;
  assign n38030 = ~n38021 & ~n38029;
  assign n38031 = pi211 & n36544;
  assign n38032 = pi212 & ~n36789;
  assign n38033 = ~n38031 & ~n38032;
  assign n38034 = ~pi219 & n38033;
  assign n38035 = n36921 & ~n38034;
  assign n38036 = pi1147 & ~n38035;
  assign n38037 = ~n38030 & n38036;
  assign n38038 = ~n36536 & n38023;
  assign n38039 = n10332 & n37997;
  assign n38040 = ~n38038 & ~n38039;
  assign n38041 = ~pi219 & ~n38040;
  assign n38042 = n37977 & ~n38041;
  assign n38043 = ~n38029 & n38042;
  assign n38044 = ~n10099 & ~n38033;
  assign n38045 = n37229 & n38044;
  assign n38046 = ~pi1147 & ~n38045;
  assign n38047 = ~n38043 & n38046;
  assign n38048 = ~pi1149 & ~n38037;
  assign n38049 = ~n38047 & n38048;
  assign n38050 = ~n36536 & n36921;
  assign n38051 = ~n37352 & n38027;
  assign n38052 = ~n38021 & ~n38051;
  assign n38053 = pi1147 & ~n38050;
  assign n38054 = ~n38052 & n38053;
  assign n38055 = ~pi1147 & ~n37712;
  assign n38056 = ~n38042 & n38055;
  assign n38057 = pi1149 & ~n38054;
  assign n38058 = ~n38056 & n38057;
  assign n38059 = pi1148 & ~n38058;
  assign n38060 = ~n38049 & n38059;
  assign n38061 = ~pi1147 & ~po1038;
  assign n38062 = n37975 & n38061;
  assign n38063 = ~pi1149 & n38062;
  assign n38064 = n10335 & n36732;
  assign n38065 = n15574 & n38064;
  assign n38066 = n37974 & n38065;
  assign n38067 = ~pi1147 & n38064;
  assign n38068 = ~n38062 & ~n38067;
  assign n38069 = pi1149 & ~n38066;
  assign n38070 = ~n38068 & n38069;
  assign n38071 = n10335 & n37712;
  assign n38072 = ~n38010 & ~n38021;
  assign n38073 = ~n38071 & ~n38072;
  assign n38074 = pi1149 & ~n38073;
  assign n38075 = ~n38010 & n38030;
  assign n38076 = ~n37729 & ~n38074;
  assign n38077 = ~n38075 & n38076;
  assign n38078 = pi1147 & ~n38077;
  assign n38079 = ~pi1148 & ~n38063;
  assign n38080 = ~n38070 & n38079;
  assign n38081 = ~n38078 & n38080;
  assign n38082 = pi213 & ~n38060;
  assign n38083 = ~n38081 & n38082;
  assign n38084 = ~pi209 & ~n38020;
  assign n38085 = ~n38083 & n38084;
  assign n38086 = ~pi211 & ~n15574;
  assign n38087 = n37756 & n38086;
  assign n38088 = n15574 & n37566;
  assign n38089 = ~n38087 & ~n38088;
  assign n38090 = ~pi1147 & n38089;
  assign n38091 = ~pi211 & ~n37636;
  assign n38092 = pi211 & ~n37647;
  assign n38093 = pi214 & ~n38092;
  assign n38094 = ~n38091 & n38093;
  assign n38095 = n10332 & ~n38094;
  assign n38096 = ~n12342 & n37636;
  assign n38097 = pi214 & n38096;
  assign n38098 = n37638 & ~n38097;
  assign n38099 = ~pi219 & ~n38098;
  assign n38100 = pi212 & ~n38096;
  assign n38101 = ~n38094 & n38100;
  assign n38102 = n38099 & ~n38101;
  assign n38103 = ~n38095 & n38102;
  assign n38104 = pi219 & n37636;
  assign n38105 = ~po1038 & ~n38104;
  assign n38106 = ~n37812 & ~n38105;
  assign n38107 = ~n38103 & ~n38106;
  assign n38108 = ~n37729 & ~n38071;
  assign n38109 = ~n38107 & n38108;
  assign n38110 = pi1147 & n38109;
  assign n38111 = pi1149 & ~n38090;
  assign n38112 = ~n38110 & n38111;
  assign n38113 = n37786 & ~n37885;
  assign n38114 = ~pi212 & ~n38022;
  assign n38115 = ~n38113 & ~n38114;
  assign n38116 = ~n37597 & ~n38115;
  assign n38117 = ~pi219 & n38116;
  assign n38118 = n36743 & ~n37039;
  assign n38119 = pi208 & ~n38118;
  assign n38120 = ~pi199 & ~n38119;
  assign n38121 = n37597 & ~n38120;
  assign n38122 = ~pi299 & ~n38121;
  assign n38123 = ~pi219 & n38122;
  assign n38124 = ~n38117 & ~n38123;
  assign n38125 = ~pi211 & ~n38124;
  assign n38126 = ~n37597 & ~n37885;
  assign n38127 = ~pi212 & ~n38126;
  assign n38128 = ~pi219 & ~n38127;
  assign n38129 = ~pi299 & ~n37150;
  assign n38130 = pi212 & ~n38129;
  assign n38131 = n37783 & ~n38022;
  assign n38132 = n38130 & ~n38131;
  assign n38133 = n38128 & ~n38132;
  assign n38134 = ~po1038 & n37597;
  assign n38135 = ~n37812 & ~n38134;
  assign n38136 = ~n38133 & ~n38135;
  assign n38137 = ~n38122 & n38136;
  assign n38138 = ~n38125 & n38137;
  assign n38139 = ~n37729 & ~n38138;
  assign n38140 = pi1147 & ~pi1149;
  assign n38141 = ~n38139 & n38140;
  assign n38142 = ~n38112 & ~n38141;
  assign n38143 = ~pi1148 & ~n38142;
  assign n38144 = ~po1038 & ~n37045;
  assign n38145 = ~n37779 & ~n38144;
  assign n38146 = n10100 & n37352;
  assign n38147 = ~pi219 & ~n38146;
  assign n38148 = n37045 & n38147;
  assign n38149 = ~n38145 & ~n38148;
  assign n38150 = ~n37712 & ~n38149;
  assign n38151 = ~pi1147 & n38150;
  assign n38152 = ~po1038 & ~n36920;
  assign n38153 = n37352 & n38152;
  assign n38154 = ~po1038 & n37150;
  assign n38155 = ~n38153 & ~n38154;
  assign n38156 = ~n38050 & n38155;
  assign n38157 = pi1147 & n38156;
  assign n38158 = pi1149 & ~n38157;
  assign n38159 = ~n38151 & n38158;
  assign n38160 = ~pi299 & ~n37571;
  assign n38161 = n10098 & ~n37567;
  assign n38162 = ~n38160 & ~n38161;
  assign n38163 = pi212 & ~n38162;
  assign n38164 = pi214 & ~n38160;
  assign n38165 = ~pi214 & n37572;
  assign n38166 = ~pi212 & ~n38164;
  assign n38167 = ~n38165 & n38166;
  assign n38168 = ~n38163 & ~n38167;
  assign n38169 = ~n37572 & ~n37609;
  assign n38170 = ~n38164 & n38169;
  assign n38171 = pi212 & ~n38170;
  assign n38172 = n38168 & n38171;
  assign n38173 = ~pi212 & n37572;
  assign n38174 = pi299 & n38031;
  assign n38175 = ~pi219 & ~n38174;
  assign n38176 = ~n38173 & n38175;
  assign n38177 = ~n38172 & n38176;
  assign n38178 = pi219 & ~n37572;
  assign n38179 = ~po1038 & ~n38178;
  assign n38180 = ~n38177 & n38179;
  assign n38181 = ~n38045 & ~n38180;
  assign n38182 = ~pi1147 & n38181;
  assign n38183 = ~n38050 & ~n38153;
  assign n38184 = ~n38034 & ~n38183;
  assign n38185 = ~n38134 & ~n38184;
  assign n38186 = pi1147 & n38185;
  assign n38187 = ~pi1149 & ~n38186;
  assign n38188 = ~n38182 & n38187;
  assign n38189 = ~n38159 & ~n38188;
  assign n38190 = pi1148 & ~n38189;
  assign n38191 = ~n38143 & ~n38190;
  assign n38192 = pi213 & ~n38191;
  assign n38193 = ~po1038 & n37979;
  assign n38194 = pi299 & ~n37947;
  assign n38195 = n34315 & n38194;
  assign n38196 = pi219 & ~n37150;
  assign n38197 = ~po1038 & ~n38196;
  assign n38198 = pi299 & n38032;
  assign n38199 = n38130 & ~n38198;
  assign n38200 = ~n37150 & ~n37885;
  assign n38201 = ~pi212 & ~n38200;
  assign n38202 = ~pi219 & ~n38201;
  assign n38203 = ~n38199 & n38202;
  assign n38204 = n38197 & ~n38203;
  assign n38205 = ~n38193 & ~n38195;
  assign n38206 = ~n38204 & n38205;
  assign n38207 = n38017 & n38206;
  assign n38208 = n37045 & n37772;
  assign n38209 = ~po1038 & ~n38208;
  assign n38210 = n10970 & n38209;
  assign n38211 = ~n37981 & ~n38210;
  assign n38212 = pi214 & n37609;
  assign n38213 = n37045 & ~n38212;
  assign n38214 = ~pi212 & ~n38213;
  assign n38215 = n37045 & ~n37967;
  assign n38216 = n38214 & ~n38215;
  assign n38217 = n37045 & ~n37988;
  assign n38218 = pi212 & ~n38217;
  assign n38219 = ~pi219 & ~n38218;
  assign n38220 = ~n38216 & n38219;
  assign n38221 = ~n38211 & ~n38220;
  assign n38222 = n37952 & ~n38221;
  assign n38223 = pi1148 & ~n38207;
  assign n38224 = ~n38222 & n38223;
  assign n38225 = n37952 & ~n38195;
  assign n38226 = ~n38193 & n38225;
  assign n38227 = ~n38088 & n38226;
  assign n38228 = ~n37981 & ~n38105;
  assign n38229 = ~n12342 & ~n37983;
  assign n38230 = ~n10332 & n38229;
  assign n38231 = pi299 & ~n37940;
  assign n38232 = n10332 & ~n38231;
  assign n38233 = ~n36536 & ~n38230;
  assign n38234 = ~n38232 & n38233;
  assign n38235 = ~pi219 & n37636;
  assign n38236 = ~n38234 & n38235;
  assign n38237 = ~n38228 & ~n38236;
  assign n38238 = n38017 & ~n38237;
  assign n38239 = ~pi1148 & ~n38238;
  assign n38240 = ~n38227 & n38239;
  assign n38241 = ~n38224 & ~n38240;
  assign n38242 = pi1149 & ~n38241;
  assign n38243 = ~n37981 & ~n38134;
  assign n38244 = n36536 & n37597;
  assign n38245 = ~pi219 & ~n38244;
  assign n38246 = ~n37597 & ~n38231;
  assign n38247 = n10332 & ~n38246;
  assign n38248 = ~n37597 & n38229;
  assign n38249 = n36675 & ~n38248;
  assign n38250 = n38245 & ~n38247;
  assign n38251 = ~n38249 & n38250;
  assign n38252 = ~n38243 & ~n38251;
  assign n38253 = n38017 & ~n38252;
  assign n38254 = ~po1038 & n37572;
  assign n38255 = n38226 & ~n38254;
  assign n38256 = pi1148 & ~n38253;
  assign n38257 = ~n38255 & n38256;
  assign n38258 = pi219 & ~n38121;
  assign n38259 = ~n36732 & n38121;
  assign n38260 = ~pi1146 & n37609;
  assign n38261 = n36675 & ~n38260;
  assign n38262 = ~n38247 & ~n38261;
  assign n38263 = ~n38259 & n38262;
  assign n38264 = ~n38122 & ~n38258;
  assign n38265 = ~n38263 & n38264;
  assign n38266 = ~n37979 & ~n38265;
  assign n38267 = ~po1038 & ~n38266;
  assign n38268 = n38017 & ~n38267;
  assign n38269 = ~pi1148 & ~n38226;
  assign n38270 = ~n38268 & n38269;
  assign n38271 = ~n38257 & ~n38270;
  assign n38272 = ~pi1149 & ~n38271;
  assign n38273 = ~n38242 & ~n38272;
  assign n38274 = ~pi213 & ~n38273;
  assign n38275 = pi209 & ~n38274;
  assign n38276 = ~n38192 & n38275;
  assign n38277 = ~n38085 & ~n38276;
  assign n38278 = pi230 & ~n38277;
  assign n38279 = ~pi230 & ~pi240;
  assign po397 = ~n38278 & ~n38279;
  assign n38281 = pi209 & ~n37796;
  assign n38282 = ~pi299 & n37045;
  assign n38283 = pi212 & ~n38282;
  assign n38284 = pi211 & ~n38282;
  assign n38285 = ~pi211 & ~n36847;
  assign n38286 = ~n10957 & n36660;
  assign n38287 = ~n37042 & ~n38286;
  assign n38288 = n38285 & ~n38287;
  assign n38289 = ~n38284 & ~n38288;
  assign n38290 = ~pi214 & n38289;
  assign n38291 = n38283 & ~n38290;
  assign n38292 = ~pi214 & n37045;
  assign n38293 = ~pi212 & ~n38292;
  assign n38294 = pi214 & n38289;
  assign n38295 = n38293 & ~n38294;
  assign n38296 = ~pi219 & ~n38291;
  assign n38297 = ~n38295 & n38296;
  assign n38298 = n38209 & ~n38297;
  assign n38299 = n37731 & ~n38298;
  assign n38300 = n38168 & n38179;
  assign n38301 = n37721 & ~n37783;
  assign n38302 = n38300 & ~n38301;
  assign n38303 = n37717 & ~n38302;
  assign n38304 = pi1152 & ~n38303;
  assign n38305 = ~n38299 & n38304;
  assign n38306 = pi214 & ~n12342;
  assign n38307 = n37045 & n38306;
  assign n38308 = n38293 & ~n38307;
  assign n38309 = pi299 & ~n37698;
  assign n38310 = n38283 & ~n38309;
  assign n38311 = ~pi219 & ~n38308;
  assign n38312 = ~n38310 & n38311;
  assign n38313 = n38209 & ~n38312;
  assign n38314 = ~n38297 & n38313;
  assign n38315 = n37758 & ~n38314;
  assign n38316 = ~n36847 & ~n38160;
  assign n38317 = ~n37567 & ~n38064;
  assign n38318 = ~po1038 & ~n38317;
  assign n38319 = n38316 & n38318;
  assign n38320 = n37777 & ~n38319;
  assign n38321 = ~pi1152 & ~n38320;
  assign n38322 = ~n38315 & n38321;
  assign n38323 = pi1150 & ~n38305;
  assign n38324 = ~n38322 & n38323;
  assign n38325 = n12343 & n36675;
  assign n38326 = pi1153 & n38325;
  assign n38327 = n37777 & ~n38326;
  assign n38328 = ~pi1152 & ~n38327;
  assign n38329 = ~n37779 & ~n38153;
  assign n38330 = ~n37790 & ~n38329;
  assign n38331 = n37758 & ~n38330;
  assign n38332 = n38328 & ~n38331;
  assign n38333 = ~n37715 & n38146;
  assign n38334 = n37717 & ~n38333;
  assign n38335 = ~pi212 & ~n37567;
  assign n38336 = ~n37610 & n38335;
  assign n38337 = ~n12342 & n38336;
  assign n38338 = ~pi219 & ~n38337;
  assign n38339 = ~n37783 & n38338;
  assign n38340 = ~n38329 & ~n38339;
  assign n38341 = n37731 & ~n38330;
  assign n38342 = ~n38340 & n38341;
  assign n38343 = pi1152 & ~n38334;
  assign n38344 = ~n38342 & n38343;
  assign n38345 = ~pi1150 & ~n38332;
  assign n38346 = ~n38344 & n38345;
  assign n38347 = ~pi1149 & ~n38346;
  assign n38348 = ~n38324 & n38347;
  assign n38349 = ~n37352 & ~n38121;
  assign n38350 = ~n36707 & n37715;
  assign n38351 = ~n38349 & ~n38350;
  assign n38352 = ~pi219 & ~n38351;
  assign n38353 = ~po1038 & ~n38258;
  assign n38354 = ~n38352 & n38353;
  assign n38355 = n37717 & ~n38354;
  assign n38356 = ~n37637 & ~n38094;
  assign n38357 = ~pi219 & ~n38356;
  assign n38358 = n37658 & ~n38198;
  assign n38359 = n38357 & n38358;
  assign n38360 = ~n38106 & ~n38359;
  assign n38361 = n37731 & ~n38360;
  assign n38362 = pi1152 & ~n38355;
  assign n38363 = ~n38361 & n38362;
  assign n38364 = pi299 & n37713;
  assign n38365 = ~n38121 & ~n38325;
  assign n38366 = ~po1038 & ~n38365;
  assign n38367 = ~n38364 & n38366;
  assign n38368 = n37777 & ~n38367;
  assign n38369 = ~n37647 & n38285;
  assign n38370 = n10719 & ~n38369;
  assign n38371 = n38107 & ~n38370;
  assign n38372 = n37758 & ~n38371;
  assign n38373 = ~pi1152 & ~n38368;
  assign n38374 = ~n38372 & n38373;
  assign n38375 = ~pi1150 & ~n38363;
  assign n38376 = ~n38374 & n38375;
  assign n38377 = ~pi219 & ~n37150;
  assign n38378 = ~n38198 & n38377;
  assign n38379 = ~pi1153 & n38378;
  assign n38380 = n10332 & n37609;
  assign n38381 = ~pi219 & ~n38380;
  assign n38382 = n37812 & ~n38381;
  assign n38383 = ~n38204 & ~n38382;
  assign n38384 = ~n38379 & ~n38383;
  assign n38385 = n37758 & ~n38384;
  assign n38386 = ~pi1151 & ~n38134;
  assign n38387 = ~pi1152 & ~n38386;
  assign n38388 = ~n38328 & ~n38387;
  assign n38389 = ~n38385 & ~n38388;
  assign n38390 = ~po1038 & ~n37615;
  assign n38391 = ~n12342 & ~n37597;
  assign n38392 = n10332 & ~n38391;
  assign n38393 = ~pi299 & ~n37597;
  assign n38394 = n36675 & ~n38364;
  assign n38395 = ~n38393 & n38394;
  assign n38396 = n38245 & ~n38392;
  assign n38397 = ~n38395 & n38396;
  assign n38398 = n38390 & ~n38397;
  assign n38399 = n37717 & ~n38398;
  assign n38400 = ~pi211 & n38378;
  assign n38401 = ~n38155 & ~n38400;
  assign n38402 = n37731 & ~n38401;
  assign n38403 = ~n38384 & n38402;
  assign n38404 = pi1152 & ~n38399;
  assign n38405 = ~n38403 & n38404;
  assign n38406 = pi1150 & ~n38389;
  assign n38407 = ~n38405 & n38406;
  assign n38408 = pi1149 & ~n38407;
  assign n38409 = ~n38376 & n38408;
  assign n38410 = ~pi209 & ~n38409;
  assign n38411 = ~n38348 & n38410;
  assign n38412 = pi213 & ~n38411;
  assign n38413 = ~n38281 & n38412;
  assign n38414 = ~pi1150 & pi1151;
  assign n38415 = ~n38089 & n38414;
  assign n38416 = ~pi1151 & ~n38045;
  assign n38417 = ~n38180 & n38416;
  assign n38418 = pi1151 & ~n37712;
  assign n38419 = ~n38149 & n38418;
  assign n38420 = pi1150 & ~n38419;
  assign n38421 = ~n38417 & n38420;
  assign n38422 = ~pi1149 & ~n38415;
  assign n38423 = ~n38421 & n38422;
  assign n38424 = n37730 & ~n38071;
  assign n38425 = ~n38107 & n38424;
  assign n38426 = ~pi1151 & ~n37729;
  assign n38427 = ~n38138 & n38426;
  assign n38428 = ~pi1150 & ~n38427;
  assign n38429 = ~n38425 & n38428;
  assign n38430 = pi1151 & ~n38050;
  assign n38431 = n38155 & n38430;
  assign n38432 = ~n38184 & n38386;
  assign n38433 = pi1150 & ~n38431;
  assign n38434 = ~n38432 & n38433;
  assign n38435 = pi1149 & ~n38434;
  assign n38436 = ~n38429 & n38435;
  assign n38437 = ~n38423 & ~n38436;
  assign n38438 = ~pi209 & ~n38437;
  assign n38439 = pi1152 & n37587;
  assign n38440 = n37582 & n38439;
  assign n38441 = ~pi1151 & n37599;
  assign n38442 = n37066 & n38441;
  assign n38443 = po1038 & ~n38064;
  assign n38444 = n37591 & n37756;
  assign n38445 = n37600 & ~n38444;
  assign n38446 = pi1152 & ~n38445;
  assign n38447 = ~n37640 & ~n38325;
  assign n38448 = ~pi1152 & ~n38447;
  assign n38449 = ~po1038 & ~n38448;
  assign n38450 = ~n38446 & n38449;
  assign n38451 = pi1151 & ~n38443;
  assign n38452 = ~n38450 & n38451;
  assign n38453 = ~n38440 & ~n38442;
  assign n38454 = ~n38452 & n38453;
  assign n38455 = ~pi1150 & ~n38454;
  assign n38456 = pi219 & ~n37599;
  assign n38457 = ~po1038 & ~n38456;
  assign n38458 = ~n38131 & n38338;
  assign n38459 = ~n37599 & n37788;
  assign n38460 = ~pi299 & n38459;
  assign n38461 = ~n38458 & ~n38460;
  assign n38462 = n38457 & n38461;
  assign n38463 = ~pi1152 & ~n38462;
  assign n38464 = ~n37582 & ~n38461;
  assign n38465 = n37719 & ~n38464;
  assign n38466 = pi1152 & ~n38465;
  assign n38467 = ~n38463 & ~n38466;
  assign n38468 = n38416 & ~n38467;
  assign n38469 = ~n38134 & ~n38457;
  assign n38470 = n37741 & ~n37747;
  assign n38471 = ~pi219 & ~n38470;
  assign n38472 = ~pi214 & n37590;
  assign n38473 = pi212 & ~n38472;
  assign n38474 = ~n37733 & n38473;
  assign n38475 = n38471 & ~n38474;
  assign n38476 = pi1152 & ~n38475;
  assign n38477 = ~pi299 & ~n37648;
  assign n38478 = ~pi214 & n37647;
  assign n38479 = pi212 & ~n38478;
  assign n38480 = ~n38097 & n38479;
  assign n38481 = n37638 & ~n37735;
  assign n38482 = ~n38480 & ~n38481;
  assign n38483 = ~n38477 & ~n38482;
  assign n38484 = ~pi219 & ~n38483;
  assign n38485 = ~pi1152 & ~n38104;
  assign n38486 = ~n38484 & n38485;
  assign n38487 = ~n38476 & ~n38486;
  assign n38488 = ~n38469 & ~n38487;
  assign n38489 = n38418 & ~n38488;
  assign n38490 = pi1150 & ~n38468;
  assign n38491 = ~n38489 & n38490;
  assign n38492 = ~pi1149 & ~n38455;
  assign n38493 = ~n38491 & n38492;
  assign n38494 = ~n37812 & ~n38457;
  assign n38495 = ~n37719 & n38494;
  assign n38496 = ~n38459 & ~n38494;
  assign n38497 = ~pi1152 & ~n38496;
  assign n38498 = pi1152 & ~n37582;
  assign n38499 = n37788 & n38498;
  assign n38500 = ~n38495 & ~n38499;
  assign n38501 = ~n38497 & n38500;
  assign n38502 = n38426 & ~n38501;
  assign n38503 = ~pi219 & ~n37768;
  assign n38504 = n37066 & ~n37773;
  assign n38505 = ~n38503 & n38504;
  assign n38506 = ~n37590 & n37698;
  assign n38507 = pi212 & n37600;
  assign n38508 = ~n38506 & n38507;
  assign n38509 = ~n37737 & ~n38508;
  assign n38510 = ~pi219 & ~n38509;
  assign n38511 = pi1152 & ~n38510;
  assign n38512 = n37740 & n38511;
  assign n38513 = n38424 & ~n38505;
  assign n38514 = ~n38512 & n38513;
  assign n38515 = ~pi1150 & ~n38502;
  assign n38516 = ~n38514 & n38515;
  assign n38517 = ~pi1151 & ~n38035;
  assign n38518 = n10332 & n37563;
  assign n38519 = ~n37611 & ~n37763;
  assign n38520 = ~n10332 & ~n38519;
  assign n38521 = ~n37582 & n38520;
  assign n38522 = ~n38518 & ~n38521;
  assign n38523 = ~pi219 & ~n38522;
  assign n38524 = ~n38495 & ~n38523;
  assign n38525 = pi1152 & ~n38524;
  assign n38526 = n38463 & ~n38496;
  assign n38527 = ~n38525 & ~n38526;
  assign n38528 = n38517 & ~n38527;
  assign n38529 = pi211 & pi219;
  assign n38530 = n37352 & ~n38529;
  assign n38531 = ~n37640 & ~n38530;
  assign n38532 = n37066 & ~n38531;
  assign n38533 = pi212 & ~n37590;
  assign n38534 = n38471 & ~n38533;
  assign n38535 = pi1152 & ~n38534;
  assign n38536 = n37740 & n38535;
  assign n38537 = n38430 & ~n38532;
  assign n38538 = ~n38536 & n38537;
  assign n38539 = pi1150 & ~n38528;
  assign n38540 = ~n38538 & n38539;
  assign n38541 = pi1149 & ~n38516;
  assign n38542 = ~n38540 & n38541;
  assign n38543 = ~n38493 & ~n38542;
  assign n38544 = pi209 & ~n38543;
  assign n38545 = ~pi213 & ~n38438;
  assign n38546 = ~n38544 & n38545;
  assign n38547 = ~n38413 & ~n38546;
  assign n38548 = pi230 & ~n38547;
  assign n38549 = ~pi230 & pi241;
  assign po398 = n38548 | n38549;
  assign n38551 = ~pi230 & ~pi242;
  assign n38552 = pi219 & ~n36527;
  assign n38553 = ~pi212 & n37941;
  assign n38554 = pi214 & ~n37356;
  assign n38555 = ~pi214 & ~n37940;
  assign n38556 = ~n38554 & ~n38555;
  assign n38557 = pi212 & ~n38556;
  assign n38558 = ~pi219 & ~n38553;
  assign n38559 = ~n38557 & n38558;
  assign n38560 = ~n36920 & ~n38552;
  assign n38561 = ~n38559 & n38560;
  assign n38562 = po1038 & n38561;
  assign n38563 = pi199 & pi1144;
  assign n38564 = ~pi200 & ~n38563;
  assign n38565 = ~n37953 & n38564;
  assign n38566 = ~pi299 & ~n37962;
  assign n38567 = ~n38565 & n38566;
  assign n38568 = n36879 & n38567;
  assign n38569 = ~pi207 & ~n38567;
  assign n38570 = ~pi299 & ~n37334;
  assign n38571 = ~n37335 & n38564;
  assign n38572 = n38570 & ~n38571;
  assign n38573 = pi207 & ~n38572;
  assign n38574 = pi208 & ~n38569;
  assign n38575 = ~n38573 & n38574;
  assign n38576 = ~n38568 & ~n38575;
  assign n38577 = n36527 & n37352;
  assign n38578 = pi219 & ~n38577;
  assign n38579 = n38576 & n38578;
  assign n38580 = ~n10332 & ~n38231;
  assign n38581 = pi299 & n38554;
  assign n38582 = ~n36675 & ~n38581;
  assign n38583 = ~n38580 & ~n38582;
  assign n38584 = ~pi219 & ~n38583;
  assign n38585 = n38576 & n38584;
  assign n38586 = ~po1038 & ~n38579;
  assign n38587 = ~n38585 & n38586;
  assign n38588 = ~n38562 & ~n38587;
  assign n38589 = pi213 & n38588;
  assign n38590 = n36536 & ~n38568;
  assign n38591 = pi211 & ~n38568;
  assign n38592 = n36522 & n38567;
  assign n38593 = n36731 & ~n36750;
  assign n38594 = pi219 & ~n38593;
  assign n38595 = ~n38592 & ~n38594;
  assign n38596 = ~n38591 & ~n38595;
  assign n38597 = pi299 & n36534;
  assign n38598 = ~n36536 & ~n38592;
  assign n38599 = ~n38597 & n38598;
  assign n38600 = ~pi219 & ~n38599;
  assign n38601 = ~n38596 & ~n38600;
  assign n38602 = ~n38590 & ~n38601;
  assign n38603 = ~n38575 & ~n38602;
  assign n38604 = ~po1038 & ~n38603;
  assign n38605 = ~pi213 & ~n36595;
  assign n38606 = ~n38604 & n38605;
  assign n38607 = ~n38589 & ~n38606;
  assign n38608 = pi209 & ~n38607;
  assign n38609 = ~n15574 & ~n38561;
  assign n38610 = pi213 & ~n38609;
  assign n38611 = ~n36525 & n38610;
  assign n38612 = ~pi213 & n36542;
  assign n38613 = ~pi209 & ~n38611;
  assign n38614 = ~n38612 & n38613;
  assign n38615 = ~n38608 & ~n38614;
  assign n38616 = pi230 & ~n38615;
  assign po399 = ~n38551 & ~n38616;
  assign n38618 = pi243 & ~pi1091;
  assign n38619 = pi1155 & ~n38618;
  assign n38620 = pi200 & pi1091;
  assign n38621 = ~pi299 & n38620;
  assign n38622 = n38619 & ~n38621;
  assign n38623 = pi1091 & ~n36629;
  assign n38624 = ~n38618 & ~n38623;
  assign n38625 = ~pi243 & ~pi1091;
  assign n38626 = ~pi1155 & n10421;
  assign n38627 = pi1091 & n36598;
  assign n38628 = ~n38626 & n38627;
  assign n38629 = ~n38625 & ~n38628;
  assign n38630 = pi1156 & ~n38629;
  assign n38631 = pi1157 & ~n38630;
  assign n38632 = ~n38622 & ~n38624;
  assign n38633 = n38631 & n38632;
  assign n38634 = pi199 & pi1091;
  assign n38635 = ~pi299 & n38634;
  assign n38636 = n38619 & ~n38635;
  assign n38637 = ~pi1155 & ~n38618;
  assign n38638 = pi1091 & ~n11036;
  assign n38639 = n38637 & ~n38638;
  assign n38640 = ~n38636 & ~n38639;
  assign n38641 = ~pi299 & pi1091;
  assign n38642 = pi200 & ~pi1156;
  assign n38643 = n38641 & n38642;
  assign n38644 = ~n38640 & ~n38643;
  assign n38645 = ~pi1157 & ~n38644;
  assign n38646 = ~pi211 & ~n38645;
  assign n38647 = ~n38633 & n38646;
  assign n38648 = pi1091 & ~n12341;
  assign n38649 = pi1156 & ~n36974;
  assign n38650 = n38648 & n38649;
  assign n38651 = ~n38619 & ~n38625;
  assign n38652 = n36610 & ~n38651;
  assign n38653 = ~n38624 & ~n38652;
  assign n38654 = ~pi1156 & ~n38653;
  assign n38655 = n38631 & ~n38654;
  assign n38656 = ~n38650 & n38655;
  assign n38657 = ~pi1156 & ~n38648;
  assign n38658 = ~n38651 & n38657;
  assign n38659 = pi1091 & n36654;
  assign n38660 = n38637 & ~n38659;
  assign n38661 = ~n38636 & ~n38660;
  assign n38662 = pi1156 & ~n38661;
  assign n38663 = ~pi1157 & ~n38658;
  assign n38664 = ~n38662 & n38663;
  assign n38665 = pi211 & ~n38664;
  assign n38666 = ~n38656 & n38665;
  assign n38667 = ~n38647 & ~n38666;
  assign n38668 = ~pi219 & ~n38667;
  assign n38669 = pi211 & n38655;
  assign n38670 = pi299 & pi1091;
  assign n38671 = n38644 & ~n38670;
  assign n38672 = ~pi1157 & ~n38671;
  assign n38673 = pi1091 & n36743;
  assign n38674 = n38637 & ~n38673;
  assign n38675 = ~n38622 & ~n38674;
  assign n38676 = ~pi1156 & ~n38675;
  assign n38677 = n36557 & ~n38650;
  assign n38678 = ~n38630 & n38677;
  assign n38679 = ~n38676 & n38678;
  assign n38680 = pi219 & ~n38672;
  assign n38681 = ~n38679 & n38680;
  assign n38682 = ~n38669 & n38681;
  assign n38683 = ~n38668 & ~n38682;
  assign n38684 = ~po1038 & n38683;
  assign n38685 = pi272 & pi283;
  assign n38686 = pi275 & n38685;
  assign n38687 = pi268 & n38686;
  assign n38688 = ~n36558 & ~n36561;
  assign n38689 = ~pi219 & ~n38688;
  assign n38690 = pi219 & n36557;
  assign n38691 = ~n38689 & ~n38690;
  assign n38692 = pi1091 & ~n38691;
  assign n38693 = ~n38625 & ~n38692;
  assign n38694 = po1038 & n38693;
  assign n38695 = ~n38687 & ~n38694;
  assign n38696 = ~n38684 & n38695;
  assign n38697 = pi253 & pi254;
  assign n38698 = pi267 & n38697;
  assign n38699 = ~pi263 & n38698;
  assign n38700 = ~n38683 & ~n38699;
  assign n38701 = ~pi83 & ~pi85;
  assign n38702 = pi314 & ~n38701;
  assign n38703 = pi802 & n38702;
  assign n38704 = pi276 & n38703;
  assign n38705 = ~pi1091 & n38704;
  assign n38706 = pi271 & n38705;
  assign n38707 = pi273 & n38706;
  assign n38708 = pi299 & ~n38707;
  assign n38709 = ~pi81 & n38701;
  assign n38710 = pi314 & ~n38709;
  assign n38711 = pi802 & n38710;
  assign n38712 = pi276 & n38711;
  assign n38713 = ~pi1091 & n38712;
  assign n38714 = ~pi1091 & ~n38704;
  assign n38715 = pi271 & ~n38714;
  assign n38716 = ~pi1091 & ~n38715;
  assign n38717 = pi273 & ~n38716;
  assign n38718 = ~pi1091 & ~n38717;
  assign n38719 = pi199 & ~n38718;
  assign n38720 = pi271 & n38713;
  assign n38721 = pi273 & n38720;
  assign n38722 = n38718 & ~n38721;
  assign n38723 = ~pi199 & ~n38722;
  assign n38724 = ~n38719 & ~n38723;
  assign n38725 = n38713 & ~n38724;
  assign n38726 = ~pi299 & ~n38725;
  assign n38727 = ~n38708 & ~n38726;
  assign n38728 = n38625 & ~n38727;
  assign n38729 = ~pi1155 & ~n38728;
  assign n38730 = pi243 & n38727;
  assign n38731 = n38729 & ~n38730;
  assign n38732 = ~n38723 & n38726;
  assign n38733 = ~pi200 & ~n38718;
  assign n38734 = n38726 & ~n38733;
  assign n38735 = ~n38708 & ~n38734;
  assign n38736 = pi243 & n38735;
  assign n38737 = ~n38732 & n38736;
  assign n38738 = ~pi200 & ~n38713;
  assign n38739 = ~n38724 & ~n38738;
  assign n38740 = ~pi299 & ~n38739;
  assign n38741 = ~n38719 & n38740;
  assign n38742 = pi299 & n38718;
  assign n38743 = ~n38741 & ~n38742;
  assign n38744 = ~pi243 & ~n38743;
  assign n38745 = pi1155 & ~n38744;
  assign n38746 = ~n38737 & n38745;
  assign n38747 = ~n38731 & ~n38746;
  assign n38748 = ~pi1156 & ~n38747;
  assign n38749 = ~n38721 & n38742;
  assign n38750 = ~n38732 & ~n38749;
  assign n38751 = ~n38740 & n38750;
  assign n38752 = ~pi1155 & ~n38751;
  assign n38753 = n38733 & n38752;
  assign n38754 = ~n38719 & n38726;
  assign n38755 = ~n38742 & ~n38754;
  assign n38756 = ~pi243 & ~n38755;
  assign n38757 = ~n38753 & n38756;
  assign n38758 = ~n38708 & ~n38732;
  assign n38759 = pi1155 & n38758;
  assign n38760 = ~n38740 & n38758;
  assign n38761 = ~n38759 & ~n38760;
  assign n38762 = pi243 & ~n38761;
  assign n38763 = pi1156 & ~n38762;
  assign n38764 = ~n38757 & n38763;
  assign n38765 = ~n38748 & ~n38764;
  assign n38766 = ~pi1157 & ~n38765;
  assign n38767 = ~n38740 & ~n38749;
  assign n38768 = ~pi243 & ~n38767;
  assign n38769 = ~n38736 & ~n38768;
  assign n38770 = pi1155 & ~n38769;
  assign n38771 = ~n38723 & n38740;
  assign n38772 = ~n38742 & ~n38771;
  assign n38773 = ~pi243 & ~n38772;
  assign n38774 = n38735 & ~n38754;
  assign n38775 = pi243 & n38774;
  assign n38776 = ~n38773 & ~n38775;
  assign n38777 = ~n38770 & n38776;
  assign n38778 = ~pi1156 & ~n38777;
  assign n38779 = ~n38733 & n38754;
  assign n38780 = ~n38742 & ~n38779;
  assign n38781 = ~pi243 & n38780;
  assign n38782 = ~n38723 & n38734;
  assign n38783 = ~n38708 & ~n38782;
  assign n38784 = ~n38741 & n38783;
  assign n38785 = pi243 & ~n38784;
  assign n38786 = ~n38781 & ~n38785;
  assign n38787 = ~pi1155 & ~n38773;
  assign n38788 = pi1155 & ~n38768;
  assign n38789 = pi243 & n38783;
  assign n38790 = n38788 & ~n38789;
  assign n38791 = ~n38787 & ~n38790;
  assign n38792 = ~n38786 & ~n38791;
  assign n38793 = pi1156 & ~n38792;
  assign n38794 = n37311 & ~n38778;
  assign n38795 = ~n38793 & n38794;
  assign n38796 = ~n38734 & ~n38742;
  assign n38797 = pi243 & ~n38796;
  assign n38798 = pi243 & n38754;
  assign n38799 = ~n38708 & ~n38771;
  assign n38800 = ~pi243 & n38799;
  assign n38801 = ~n38798 & ~n38800;
  assign n38802 = ~pi1155 & ~n38801;
  assign n38803 = n38788 & n38800;
  assign n38804 = ~pi1156 & ~n38797;
  assign n38805 = ~n38803 & n38804;
  assign n38806 = ~n38802 & n38805;
  assign n38807 = ~n38708 & ~n38740;
  assign n38808 = n38781 & n38807;
  assign n38809 = ~n38784 & n38797;
  assign n38810 = pi1155 & ~n38809;
  assign n38811 = ~n38808 & n38810;
  assign n38812 = pi299 & ~n38721;
  assign n38813 = ~n38779 & ~n38812;
  assign n38814 = ~n38618 & ~n38813;
  assign n38815 = n38776 & ~n38814;
  assign n38816 = ~pi1155 & ~n38815;
  assign n38817 = ~n38811 & ~n38816;
  assign n38818 = pi1156 & ~n38817;
  assign n38819 = n36557 & ~n38806;
  assign n38820 = ~n38818 & n38819;
  assign n38821 = ~n38766 & ~n38795;
  assign n38822 = ~n38820 & n38821;
  assign n38823 = pi219 & ~n38822;
  assign n38824 = ~n38740 & ~n38812;
  assign n38825 = ~pi243 & n38824;
  assign n38826 = ~n38734 & ~n38749;
  assign n38827 = pi243 & ~n38826;
  assign n38828 = ~n38825 & ~n38827;
  assign n38829 = ~n38741 & ~n38812;
  assign n38830 = ~n38782 & n38829;
  assign n38831 = pi243 & ~n38830;
  assign n38832 = ~n38771 & ~n38779;
  assign n38833 = ~pi243 & ~n38749;
  assign n38834 = n38832 & n38833;
  assign n38835 = ~n38831 & ~n38834;
  assign n38836 = n38828 & n38835;
  assign n38837 = ~pi1155 & ~n38836;
  assign n38838 = ~pi1156 & ~n38837;
  assign n38839 = n38828 & n38838;
  assign n38840 = ~n38749 & ~n38782;
  assign n38841 = pi1155 & n38840;
  assign n38842 = ~n38810 & ~n38841;
  assign n38843 = ~n38779 & n38825;
  assign n38844 = ~n38842 & ~n38843;
  assign n38845 = ~pi1155 & n38835;
  assign n38846 = ~n38844 & ~n38845;
  assign n38847 = pi1156 & ~n38846;
  assign n38848 = pi1157 & ~n38839;
  assign n38849 = ~n38847 & n38848;
  assign n38850 = ~pi1155 & n38826;
  assign n38851 = ~n38824 & n38850;
  assign n38852 = ~n38726 & ~n38812;
  assign n38853 = pi243 & n38852;
  assign n38854 = ~n38754 & ~n38812;
  assign n38855 = ~n38618 & ~n38854;
  assign n38856 = ~n38853 & ~n38855;
  assign n38857 = pi1156 & ~n38856;
  assign n38858 = ~n38753 & n38857;
  assign n38859 = ~n38851 & n38858;
  assign n38860 = ~pi1155 & n38852;
  assign n38861 = ~n38729 & ~n38860;
  assign n38862 = ~n38853 & ~n38861;
  assign n38863 = ~pi1156 & ~n38862;
  assign n38864 = n38828 & ~n38856;
  assign n38865 = pi1155 & ~n38864;
  assign n38866 = n38863 & ~n38865;
  assign n38867 = ~pi1157 & ~n38859;
  assign n38868 = ~n38866 & n38867;
  assign n38869 = ~pi211 & ~n38868;
  assign n38870 = ~n38849 & n38869;
  assign n38871 = ~n38734 & ~n38812;
  assign n38872 = pi243 & n38871;
  assign n38873 = n38788 & ~n38872;
  assign n38874 = n38619 & n38719;
  assign n38875 = ~n38873 & ~n38874;
  assign n38876 = n38863 & n38875;
  assign n38877 = ~pi1157 & ~n38858;
  assign n38878 = ~n38876 & n38877;
  assign n38879 = n38838 & ~n38873;
  assign n38880 = ~n38814 & n38846;
  assign n38881 = pi1156 & ~n38880;
  assign n38882 = pi1157 & ~n38879;
  assign n38883 = ~n38881 & n38882;
  assign n38884 = pi211 & ~n38878;
  assign n38885 = ~n38883 & n38884;
  assign n38886 = ~pi219 & ~n38870;
  assign n38887 = ~n38885 & n38886;
  assign n38888 = n38699 & ~n38823;
  assign n38889 = ~n38887 & n38888;
  assign n38890 = ~po1038 & ~n38700;
  assign n38891 = ~n38889 & n38890;
  assign n38892 = pi1091 & n38688;
  assign n38893 = pi243 & n38722;
  assign n38894 = ~pi243 & n38721;
  assign n38895 = ~n38892 & ~n38894;
  assign n38896 = ~n38893 & n38895;
  assign n38897 = ~pi219 & ~n38896;
  assign n38898 = ~pi243 & n38718;
  assign n38899 = n36557 & ~n38618;
  assign n38900 = ~n38705 & n38899;
  assign n38901 = pi243 & n38707;
  assign n38902 = pi219 & ~n38900;
  assign n38903 = ~n38901 & n38902;
  assign n38904 = ~n38898 & n38903;
  assign n38905 = n38699 & ~n38904;
  assign n38906 = ~n38897 & n38905;
  assign n38907 = ~n38693 & ~n38699;
  assign n38908 = po1038 & ~n38907;
  assign n38909 = ~n38906 & n38908;
  assign n38910 = n38687 & ~n38909;
  assign n38911 = ~n38891 & n38910;
  assign n38912 = ~pi230 & ~n38696;
  assign n38913 = ~n38911 & n38912;
  assign n38914 = ~n15574 & ~n38691;
  assign n38915 = ~pi200 & pi1157;
  assign n38916 = pi199 & ~n38915;
  assign n38917 = ~n38626 & ~n38642;
  assign n38918 = ~n38916 & n38917;
  assign n38919 = n15574 & n38918;
  assign n38920 = pi230 & ~n38914;
  assign n38921 = ~n38919 & n38920;
  assign po400 = ~n38913 & ~n38921;
  assign n38923 = ~pi230 & ~pi244;
  assign n38924 = pi213 & ~n38019;
  assign n38925 = pi299 & n37356;
  assign n38926 = ~n38003 & ~n38925;
  assign n38927 = pi214 & ~n38926;
  assign n38928 = n37999 & ~n38927;
  assign n38929 = n36528 & n37828;
  assign n38930 = ~pi214 & ~n38926;
  assign n38931 = pi212 & ~n38929;
  assign n38932 = ~n38930 & n38931;
  assign n38933 = ~n38003 & n38932;
  assign n38934 = ~pi219 & ~n38928;
  assign n38935 = ~n38933 & n38934;
  assign n38936 = pi299 & n37353;
  assign n38937 = pi1147 & ~n38936;
  assign n38938 = ~n38021 & n38937;
  assign n38939 = ~n38935 & n38938;
  assign n38940 = n37986 & ~n38927;
  assign n38941 = ~n38932 & ~n38940;
  assign n38942 = ~n38023 & ~n38941;
  assign n38943 = ~pi219 & ~n38942;
  assign n38944 = ~n37353 & ~n37772;
  assign n38945 = ~n37975 & ~n38944;
  assign n38946 = n38061 & ~n38945;
  assign n38947 = ~n38943 & n38946;
  assign n38948 = ~pi213 & ~n37367;
  assign n38949 = ~n38939 & n38948;
  assign n38950 = ~n38947 & n38949;
  assign n38951 = ~n38924 & ~n38950;
  assign n38952 = pi209 & ~n38951;
  assign n38953 = ~pi213 & ~n37368;
  assign n38954 = ~n38017 & ~n38225;
  assign n38955 = n37952 & ~n38194;
  assign n38956 = n36732 & ~n38230;
  assign n38957 = ~n38232 & n38956;
  assign n38958 = ~n38955 & n38957;
  assign n38959 = ~n37340 & ~n37979;
  assign n38960 = ~n38958 & n38959;
  assign n38961 = ~po1038 & ~n38960;
  assign n38962 = ~n38954 & ~n38961;
  assign n38963 = pi213 & ~n38962;
  assign n38964 = ~pi209 & ~n38953;
  assign n38965 = ~n38963 & n38964;
  assign n38966 = ~n38952 & ~n38965;
  assign n38967 = pi230 & ~n38966;
  assign po401 = ~n38923 & ~n38967;
  assign n38969 = ~pi213 & n38588;
  assign n38970 = pi1146 & n37729;
  assign n38971 = ~pi1147 & ~n38970;
  assign n38972 = ~n38015 & n38971;
  assign n38973 = n37352 & n37938;
  assign n38974 = pi219 & ~n38973;
  assign n38975 = n38576 & n38974;
  assign n38976 = ~po1038 & ~n38975;
  assign n38977 = n38001 & n38576;
  assign n38978 = pi212 & ~n38977;
  assign n38979 = ~pi214 & n38576;
  assign n38980 = ~n12342 & n38979;
  assign n38981 = n38978 & ~n38980;
  assign n38982 = ~n12342 & n38576;
  assign n38983 = ~pi212 & ~n38979;
  assign n38984 = ~n38982 & n38983;
  assign n38985 = ~pi219 & ~n38981;
  assign n38986 = ~n38984 & n38985;
  assign n38987 = n38976 & ~n38986;
  assign n38988 = n38972 & ~n38987;
  assign n38989 = pi299 & n38983;
  assign n38990 = n10098 & ~n37967;
  assign n38991 = pi299 & ~n38990;
  assign n38992 = n38576 & ~n38991;
  assign n38993 = pi212 & ~n38992;
  assign n38994 = ~pi212 & ~n38576;
  assign n38995 = ~pi219 & ~n38994;
  assign n38996 = ~n38993 & n38995;
  assign n38997 = ~n38989 & n38996;
  assign n38998 = n38976 & ~n38997;
  assign n38999 = pi1147 & ~n37712;
  assign n39000 = ~n38970 & n38999;
  assign n39001 = ~n38998 & n39000;
  assign n39002 = ~n38988 & ~n39001;
  assign n39003 = pi1148 & ~n39002;
  assign n39004 = n38978 & ~n38979;
  assign n39005 = n38995 & ~n39004;
  assign n39006 = n38976 & ~n39005;
  assign n39007 = n38971 & ~n39006;
  assign n39008 = ~n38036 & ~n39000;
  assign n39009 = ~n37609 & n38576;
  assign n39010 = ~n38983 & ~n38993;
  assign n39011 = ~n39009 & ~n39010;
  assign n39012 = pi214 & n38993;
  assign n39013 = ~pi219 & ~n39012;
  assign n39014 = ~n39011 & n39013;
  assign n39015 = n38976 & ~n39014;
  assign n39016 = ~n39008 & ~n39015;
  assign n39017 = ~n39007 & ~n39016;
  assign n39018 = ~pi1148 & ~n39017;
  assign n39019 = ~n39003 & ~n39018;
  assign n39020 = pi213 & ~n39019;
  assign n39021 = ~pi209 & ~n38969;
  assign n39022 = ~n39020 & n39021;
  assign n39023 = pi199 & pi1146;
  assign n39024 = n36628 & ~n39023;
  assign n39025 = pi208 & ~n39024;
  assign n39026 = n37955 & n39025;
  assign n39027 = ~n36879 & ~n39026;
  assign n39028 = n36598 & ~n39027;
  assign n39029 = ~n39024 & n39028;
  assign n39030 = ~n37828 & ~n39029;
  assign n39031 = ~pi212 & ~n39030;
  assign n39032 = ~n38991 & ~n39029;
  assign n39033 = pi212 & ~n39032;
  assign n39034 = ~pi219 & ~n39031;
  assign n39035 = ~n39033 & n39034;
  assign n39036 = n38974 & ~n39029;
  assign n39037 = ~po1038 & ~n39036;
  assign n39038 = ~n39035 & n39037;
  assign n39039 = n39000 & ~n39038;
  assign n39040 = ~pi208 & n37967;
  assign n39041 = n37634 & ~n39024;
  assign n39042 = ~pi200 & ~n39023;
  assign n39043 = n37955 & ~n39042;
  assign n39044 = ~pi299 & ~n39043;
  assign n39045 = pi1146 & n38119;
  assign n39046 = ~n39044 & n39045;
  assign n39047 = ~n39040 & ~n39041;
  assign n39048 = ~n39046 & n39047;
  assign n39049 = ~pi299 & ~n39048;
  assign n39050 = ~n36731 & n39049;
  assign n39051 = pi219 & ~n39050;
  assign n39052 = n36731 & ~n39048;
  assign n39053 = n39051 & ~n39052;
  assign n39054 = ~pi214 & ~n39049;
  assign n39055 = ~pi212 & ~n39054;
  assign n39056 = ~n10101 & ~n37634;
  assign n39057 = n39043 & ~n39056;
  assign n39058 = pi211 & ~n39057;
  assign n39059 = ~n39044 & ~n39048;
  assign n39060 = ~pi299 & ~n39059;
  assign n39061 = ~pi211 & n39060;
  assign n39062 = ~n39058 & ~n39061;
  assign n39063 = ~n39049 & ~n39062;
  assign n39064 = n39055 & ~n39063;
  assign n39065 = ~pi214 & n39063;
  assign n39066 = n38001 & ~n39049;
  assign n39067 = pi212 & ~n39066;
  assign n39068 = ~n39065 & n39067;
  assign n39069 = ~pi219 & ~n39064;
  assign n39070 = ~n39068 & n39069;
  assign n39071 = ~po1038 & ~n39053;
  assign n39072 = ~n39070 & n39071;
  assign n39073 = n38972 & ~n39072;
  assign n39074 = pi1148 & ~n39039;
  assign n39075 = ~n39073 & n39074;
  assign n39076 = ~pi219 & ~n37945;
  assign n39077 = ~n38381 & ~n39076;
  assign n39078 = ~n39057 & ~n39077;
  assign n39079 = pi219 & ~n39057;
  assign n39080 = ~n36999 & ~n39079;
  assign n39081 = ~n36536 & ~n39058;
  assign n39082 = n39059 & n39081;
  assign n39083 = ~n39080 & ~n39082;
  assign n39084 = ~po1038 & ~n39078;
  assign n39085 = ~n39083 & n39084;
  assign n39086 = n38971 & ~n39085;
  assign n39087 = ~n10101 & n39042;
  assign n39088 = n39028 & ~n39087;
  assign n39089 = n38114 & ~n39088;
  assign n39090 = ~pi299 & ~n39088;
  assign n39091 = pi214 & ~n39090;
  assign n39092 = ~n12342 & ~n39029;
  assign n39093 = n39091 & ~n39092;
  assign n39094 = pi212 & ~n39093;
  assign n39095 = ~pi214 & n39088;
  assign n39096 = ~n37785 & ~n39095;
  assign n39097 = n39094 & n39096;
  assign n39098 = ~n39089 & ~n39097;
  assign n39099 = ~pi219 & ~n39098;
  assign n39100 = n38198 & ~n38990;
  assign n39101 = n39099 & ~n39100;
  assign n39102 = pi219 & ~n39088;
  assign n39103 = ~n38973 & n39102;
  assign n39104 = ~po1038 & ~n39103;
  assign n39105 = ~n39101 & n39104;
  assign n39106 = ~n39008 & ~n39105;
  assign n39107 = ~pi1148 & ~n39086;
  assign n39108 = ~n39106 & n39107;
  assign n39109 = ~n39075 & ~n39108;
  assign n39110 = pi213 & n39109;
  assign n39111 = ~pi214 & n39057;
  assign n39112 = ~n38231 & ~n39049;
  assign n39113 = pi214 & ~n39060;
  assign n39114 = ~n39112 & n39113;
  assign n39115 = ~n39111 & ~n39114;
  assign n39116 = ~pi212 & ~n39115;
  assign n39117 = pi299 & ~n38556;
  assign n39118 = ~n39049 & ~n39117;
  assign n39119 = pi212 & ~n39118;
  assign n39120 = ~n39044 & n39119;
  assign n39121 = ~pi219 & ~n39120;
  assign n39122 = ~n39116 & n39121;
  assign n39123 = ~n36536 & ~n36680;
  assign n39124 = n39062 & n39123;
  assign n39125 = ~n39080 & ~n39124;
  assign n39126 = n38061 & ~n39125;
  assign n39127 = ~n39122 & n39126;
  assign n39128 = ~n38577 & n39102;
  assign n39129 = ~pi212 & n39095;
  assign n39130 = ~pi214 & ~n39029;
  assign n39131 = ~pi212 & ~n39130;
  assign n39132 = ~n38231 & ~n39029;
  assign n39133 = n39131 & ~n39132;
  assign n39134 = n39091 & n39133;
  assign n39135 = ~n39029 & ~n39117;
  assign n39136 = pi212 & ~n39135;
  assign n39137 = ~n39090 & n39136;
  assign n39138 = ~pi219 & ~n39129;
  assign n39139 = ~n39137 & n39138;
  assign n39140 = ~n39134 & n39139;
  assign n39141 = pi1147 & ~po1038;
  assign n39142 = ~n39128 & n39141;
  assign n39143 = ~n39140 & n39142;
  assign n39144 = ~pi1148 & ~n38562;
  assign n39145 = ~n39143 & n39144;
  assign n39146 = ~n39127 & n39145;
  assign n39147 = n39055 & ~n39112;
  assign n39148 = ~pi219 & ~n39119;
  assign n39149 = ~n39147 & n39148;
  assign n39150 = ~pi299 & n39048;
  assign n39151 = n36731 & ~n39150;
  assign n39152 = ~n36680 & n39151;
  assign n39153 = n39051 & ~n39152;
  assign n39154 = n38061 & ~n39153;
  assign n39155 = ~n39149 & n39154;
  assign n39156 = n38578 & ~n39029;
  assign n39157 = ~pi219 & ~n39136;
  assign n39158 = ~n39133 & n39157;
  assign n39159 = n39141 & ~n39156;
  assign n39160 = ~n39158 & n39159;
  assign n39161 = pi1148 & ~n38562;
  assign n39162 = ~n39160 & n39161;
  assign n39163 = ~n39155 & n39162;
  assign n39164 = ~n39146 & ~n39163;
  assign n39165 = ~pi213 & ~n39164;
  assign n39166 = pi209 & ~n39165;
  assign n39167 = ~n39110 & n39166;
  assign n39168 = ~n39022 & ~n39167;
  assign n39169 = pi230 & ~n39168;
  assign n39170 = ~pi230 & pi245;
  assign po402 = n39169 | n39170;
  assign n39172 = ~pi209 & n39109;
  assign n39173 = ~n38972 & ~n39000;
  assign n39174 = ~po1038 & ~n38974;
  assign n39175 = ~n38134 & ~n39174;
  assign n39176 = ~n37597 & ~n38002;
  assign n39177 = pi212 & ~n39176;
  assign n39178 = n38132 & ~n38391;
  assign n39179 = n38116 & ~n39178;
  assign n39180 = ~n38972 & ~n39179;
  assign n39181 = n38128 & ~n39177;
  assign n39182 = ~n39180 & n39181;
  assign n39183 = ~n39175 & ~n39182;
  assign n39184 = ~n39173 & ~n39183;
  assign n39185 = ~pi1150 & ~n39184;
  assign n39186 = n39077 & n39174;
  assign n39187 = ~n38204 & ~n39186;
  assign n39188 = n38972 & n39187;
  assign n39189 = pi1146 & n38153;
  assign n39190 = ~n38146 & n38377;
  assign n39191 = n38197 & ~n39190;
  assign n39192 = ~n39189 & ~n39191;
  assign n39193 = n39000 & n39192;
  assign n39194 = pi1150 & ~n39193;
  assign n39195 = ~n39188 & n39194;
  assign n39196 = pi1148 & ~n39195;
  assign n39197 = ~n39185 & n39196;
  assign n39198 = ~n38179 & ~n39189;
  assign n39199 = n38177 & ~n39077;
  assign n39200 = ~n39198 & ~n39199;
  assign n39201 = ~n39008 & ~n39200;
  assign n39202 = ~pi1146 & ~n37572;
  assign n39203 = ~n38254 & ~n38382;
  assign n39204 = ~n39202 & ~n39203;
  assign n39205 = n38971 & ~n39204;
  assign n39206 = ~n39201 & ~n39205;
  assign n39207 = ~pi1150 & ~n39206;
  assign n39208 = ~n38971 & n39008;
  assign n39209 = ~n38210 & ~n39174;
  assign n39210 = ~n37609 & n38292;
  assign n39211 = pi212 & ~n38307;
  assign n39212 = ~n39210 & n39211;
  assign n39213 = ~pi219 & ~n39212;
  assign n39214 = ~n38214 & n39213;
  assign n39215 = n38215 & n39214;
  assign n39216 = n38213 & n39213;
  assign n39217 = ~n38313 & n38971;
  assign n39218 = ~n39209 & ~n39216;
  assign n39219 = ~n39215 & n39218;
  assign n39220 = ~n39217 & n39219;
  assign n39221 = pi1150 & ~n39208;
  assign n39222 = ~n39220 & n39221;
  assign n39223 = ~n39207 & ~n39222;
  assign n39224 = ~pi1148 & ~n39223;
  assign n39225 = pi1149 & ~n39197;
  assign n39226 = ~n39224 & n39225;
  assign n39227 = pi1150 & n38088;
  assign n39228 = pi299 & n38044;
  assign n39229 = n39174 & n39228;
  assign n39230 = ~n38971 & n39229;
  assign n39231 = ~pi1148 & ~n39186;
  assign n39232 = ~n39227 & n39231;
  assign n39233 = ~n39230 & n39232;
  assign n39234 = ~n39208 & n39233;
  assign n39235 = ~n38105 & ~n39174;
  assign n39236 = n37636 & ~n38002;
  assign n39237 = pi212 & ~n39236;
  assign n39238 = n38099 & ~n39237;
  assign n39239 = ~n39235 & ~n39238;
  assign n39240 = n38972 & ~n39239;
  assign n39241 = ~pi212 & ~n37636;
  assign n39242 = ~pi219 & ~n39241;
  assign n39243 = ~n38336 & n39242;
  assign n39244 = ~n38480 & n39243;
  assign n39245 = ~n39237 & n39244;
  assign n39246 = ~n39235 & ~n39245;
  assign n39247 = n39000 & ~n39246;
  assign n39248 = ~n39240 & ~n39247;
  assign n39249 = pi1150 & ~n39248;
  assign n39250 = ~n38123 & ~n38133;
  assign n39251 = n38972 & ~n39250;
  assign n39252 = ~po1038 & n38121;
  assign n39253 = ~n39174 & ~n39252;
  assign n39254 = ~n36675 & n38260;
  assign n39255 = ~n38349 & ~n39254;
  assign n39256 = ~pi219 & ~n39255;
  assign n39257 = ~n39253 & ~n39256;
  assign n39258 = ~n39251 & n39257;
  assign n39259 = ~pi1150 & ~n39173;
  assign n39260 = ~n39258 & n39259;
  assign n39261 = ~n39249 & ~n39260;
  assign n39262 = pi1148 & ~n39261;
  assign n39263 = ~pi1149 & ~n39234;
  assign n39264 = ~n39262 & n39263;
  assign n39265 = pi209 & ~n39264;
  assign n39266 = ~n39226 & n39265;
  assign n39267 = ~pi213 & ~n39172;
  assign n39268 = ~n39266 & n39267;
  assign n39269 = n37772 & ~n39029;
  assign n39270 = n39141 & ~n39269;
  assign n39271 = pi214 & ~n37609;
  assign n39272 = ~n39029 & n39271;
  assign n39273 = ~n12342 & n39130;
  assign n39274 = pi212 & ~n39272;
  assign n39275 = ~n39273 & n39274;
  assign n39276 = ~n39092 & n39131;
  assign n39277 = ~pi219 & ~n39275;
  assign n39278 = ~n39276 & n39277;
  assign n39279 = n39270 & ~n39278;
  assign n39280 = n39051 & ~n39151;
  assign n39281 = n38061 & ~n39280;
  assign n39282 = ~n38380 & n39070;
  assign n39283 = n39281 & ~n39282;
  assign n39284 = pi1150 & n38108;
  assign n39285 = ~n39279 & n39284;
  assign n39286 = ~n39283 & n39285;
  assign n39287 = ~pi219 & ~n39029;
  assign n39288 = ~n38380 & n39287;
  assign n39289 = n39270 & ~n39288;
  assign n39290 = n38381 & ~n39049;
  assign n39291 = n39281 & ~n39290;
  assign n39292 = ~pi1150 & ~n37729;
  assign n39293 = ~n39289 & n39292;
  assign n39294 = ~n39291 & n39293;
  assign n39295 = ~pi1149 & ~n39294;
  assign n39296 = ~n39286 & n39295;
  assign n39297 = pi57 & n36733;
  assign n39298 = ~n36733 & ~n39150;
  assign n39299 = ~n6258 & ~n36733;
  assign n39300 = ~pi57 & ~n39299;
  assign n39301 = n6258 & ~n36732;
  assign n39302 = n39050 & n39301;
  assign n39303 = ~pi1147 & n39300;
  assign n39304 = ~n39298 & n39303;
  assign n39305 = ~n39302 & n39304;
  assign n39306 = ~n38530 & ~n39029;
  assign n39307 = n6258 & ~n39306;
  assign n39308 = pi1147 & n39300;
  assign n39309 = ~n39307 & n39308;
  assign n39310 = ~n39297 & ~n39309;
  assign n39311 = ~n39305 & n39310;
  assign n39312 = pi1150 & ~n39311;
  assign n39313 = ~n37609 & ~n39057;
  assign n39314 = ~n36536 & ~n39313;
  assign n39315 = pi212 & n39113;
  assign n39316 = ~pi219 & ~n39314;
  assign n39317 = ~n39049 & n39316;
  assign n39318 = ~n39315 & n39317;
  assign n39319 = n39281 & ~n39318;
  assign n39320 = ~n38400 & n39141;
  assign n39321 = ~n39306 & n39320;
  assign n39322 = ~pi1150 & ~n38035;
  assign n39323 = ~n39321 & n39322;
  assign n39324 = ~n39319 & n39323;
  assign n39325 = pi1149 & ~n39312;
  assign n39326 = ~n39324 & n39325;
  assign n39327 = ~n39296 & ~n39326;
  assign n39328 = pi1148 & ~n39327;
  assign n39329 = ~n39102 & n39141;
  assign n39330 = ~n39099 & n39329;
  assign n39331 = ~pi1150 & ~n38045;
  assign n39332 = ~pi214 & ~n39313;
  assign n39333 = pi214 & n39062;
  assign n39334 = pi212 & ~n39333;
  assign n39335 = ~pi219 & ~n39332;
  assign n39336 = n39334 & n39335;
  assign n39337 = ~pi219 & ~n38114;
  assign n39338 = ~n39057 & ~n39337;
  assign n39339 = n38061 & ~n39338;
  assign n39340 = ~n39336 & n39339;
  assign n39341 = ~n39330 & n39331;
  assign n39342 = ~n39340 & n39341;
  assign n39343 = ~pi214 & ~n39060;
  assign n39344 = n39334 & ~n39343;
  assign n39345 = ~pi212 & ~n39111;
  assign n39346 = ~n39113 & n39345;
  assign n39347 = ~n39344 & ~n39346;
  assign n39348 = ~pi219 & ~n39347;
  assign n39349 = ~n39079 & ~n39348;
  assign n39350 = ~pi1147 & ~n39349;
  assign n39351 = pi299 & n36732;
  assign n39352 = ~n39088 & ~n39351;
  assign n39353 = pi214 & n39287;
  assign n39354 = n39094 & n39353;
  assign n39355 = ~n39352 & ~n39354;
  assign n39356 = pi1147 & ~n39355;
  assign n39357 = ~po1038 & ~n39356;
  assign n39358 = ~n39350 & n39357;
  assign n39359 = pi1150 & ~n37712;
  assign n39360 = ~n39358 & n39359;
  assign n39361 = ~n39342 & ~n39360;
  assign n39362 = pi1149 & ~n39361;
  assign n39363 = pi1150 & n38064;
  assign n39364 = n39057 & ~n39363;
  assign n39365 = ~pi1147 & ~n39364;
  assign n39366 = pi1147 & ~n39088;
  assign n39367 = ~po1038 & ~n39365;
  assign n39368 = ~n39366 & n39367;
  assign n39369 = ~pi1147 & n39059;
  assign n39370 = n15574 & ~n39369;
  assign n39371 = n39363 & ~n39370;
  assign n39372 = ~pi1149 & ~n39368;
  assign n39373 = ~n39371 & n39372;
  assign n39374 = ~pi1148 & ~n39373;
  assign n39375 = ~n39362 & n39374;
  assign n39376 = ~pi209 & ~n39328;
  assign n39377 = ~n39375 & n39376;
  assign n39378 = pi1150 & n38150;
  assign n39379 = ~n38180 & n39331;
  assign n39380 = pi1149 & ~n39378;
  assign n39381 = ~n39379 & n39380;
  assign n39382 = ~pi1149 & pi1150;
  assign n39383 = ~n38089 & n39382;
  assign n39384 = ~n39381 & ~n39383;
  assign n39385 = ~pi1148 & ~n39384;
  assign n39386 = ~pi1150 & ~n38185;
  assign n39387 = pi1150 & ~n38156;
  assign n39388 = pi1149 & ~n39387;
  assign n39389 = ~n39386 & n39388;
  assign n39390 = pi1150 & ~n38109;
  assign n39391 = ~pi1150 & ~n38139;
  assign n39392 = ~pi1149 & ~n39391;
  assign n39393 = ~n39390 & n39392;
  assign n39394 = pi1148 & ~n39389;
  assign n39395 = ~n39393 & n39394;
  assign n39396 = ~n39385 & ~n39395;
  assign n39397 = pi209 & n39396;
  assign n39398 = pi213 & ~n39397;
  assign n39399 = ~n39377 & n39398;
  assign n39400 = ~n39268 & ~n39399;
  assign n39401 = pi230 & ~n39400;
  assign n39402 = ~pi230 & pi246;
  assign po403 = n39401 | n39402;
  assign n39404 = pi213 & ~n38437;
  assign n39405 = ~pi1151 & ~n37712;
  assign n39406 = ~n36675 & n38126;
  assign n39407 = ~n38122 & ~n39406;
  assign n39408 = n38353 & n39407;
  assign n39409 = n39405 & ~n39408;
  assign n39410 = n38105 & ~n39244;
  assign n39411 = ~n37712 & ~n39410;
  assign n39412 = pi1151 & n39411;
  assign n39413 = ~pi1147 & ~n39409;
  assign n39414 = ~n39412 & n39413;
  assign n39415 = pi212 & ~n37647;
  assign n39416 = n39243 & ~n39415;
  assign n39417 = ~n38106 & ~n39416;
  assign n39418 = n38430 & ~n39417;
  assign n39419 = pi1147 & ~n39418;
  assign n39420 = ~pi1151 & ~n38050;
  assign n39421 = ~n39408 & n39420;
  assign n39422 = ~n38137 & n39421;
  assign n39423 = n39419 & ~n39422;
  assign n39424 = pi1149 & ~n39423;
  assign n39425 = ~n39414 & n39424;
  assign n39426 = ~pi219 & ~n15574;
  assign n39427 = n38044 & n39426;
  assign n39428 = ~pi1151 & ~n39427;
  assign n39429 = ~pi1147 & ~n39428;
  assign n39430 = pi1151 & ~n38045;
  assign n39431 = n37779 & ~n38458;
  assign n39432 = n39430 & ~n39431;
  assign n39433 = n39429 & ~n39432;
  assign n39434 = pi1151 & ~n38035;
  assign n39435 = ~n38340 & n39434;
  assign n39436 = ~pi1151 & ~n38184;
  assign n39437 = pi1147 & ~n39436;
  assign n39438 = ~n39435 & n39437;
  assign n39439 = ~pi1149 & ~n39433;
  assign n39440 = ~n39438 & n39439;
  assign n39441 = ~pi1150 & ~n39440;
  assign n39442 = ~n39425 & n39441;
  assign n39443 = pi1147 & ~n38431;
  assign n39444 = n38183 & n38386;
  assign n39445 = n39443 & ~n39444;
  assign n39446 = n38128 & ~n39178;
  assign n39447 = n38390 & ~n39446;
  assign n39448 = ~n38117 & n38390;
  assign n39449 = ~n39447 & ~n39448;
  assign n39450 = n39405 & n39449;
  assign n39451 = n38418 & ~n39191;
  assign n39452 = ~pi1147 & ~n39451;
  assign n39453 = ~n39450 & n39452;
  assign n39454 = pi1149 & ~n39445;
  assign n39455 = ~n39453 & n39454;
  assign n39456 = n38209 & ~n39216;
  assign n39457 = n39434 & ~n39456;
  assign n39458 = ~n38171 & n38176;
  assign n39459 = ~n38153 & ~n38179;
  assign n39460 = ~n39458 & ~n39459;
  assign n39461 = ~n38035 & ~n39460;
  assign n39462 = ~pi1151 & n39461;
  assign n39463 = pi1147 & ~n39457;
  assign n39464 = ~n39462 & n39463;
  assign n39465 = ~pi1147 & ~n38417;
  assign n39466 = ~n38145 & ~n39214;
  assign n39467 = n39430 & ~n39466;
  assign n39468 = n39465 & ~n39467;
  assign n39469 = ~pi1149 & ~n39464;
  assign n39470 = ~n39468 & n39469;
  assign n39471 = pi1150 & ~n39455;
  assign n39472 = ~n39470 & n39471;
  assign n39473 = pi1148 & ~n39442;
  assign n39474 = ~n39472 & n39473;
  assign n39475 = pi1151 & n38088;
  assign n39476 = ~n37729 & ~n38382;
  assign n39477 = pi1147 & ~n39476;
  assign n39478 = ~pi1150 & ~n39475;
  assign n39479 = ~n39477 & n39478;
  assign n39480 = ~pi1151 & ~n38254;
  assign n39481 = ~pi1147 & ~n39480;
  assign n39482 = pi1151 & ~n38144;
  assign n39483 = n39481 & ~n39482;
  assign n39484 = ~n38312 & n39456;
  assign n39485 = n37730 & ~n39484;
  assign n39486 = n38426 & n39203;
  assign n39487 = pi1147 & ~n39486;
  assign n39488 = ~n39485 & n39487;
  assign n39489 = pi1150 & ~n39483;
  assign n39490 = ~n39488 & n39489;
  assign n39491 = ~pi1149 & ~n39479;
  assign n39492 = ~n39490 & n39491;
  assign n39493 = ~n38102 & n38105;
  assign n39494 = pi1151 & ~n38015;
  assign n39495 = ~n39493 & n39494;
  assign n39496 = ~pi1151 & ~n38015;
  assign n39497 = ~n38366 & n39496;
  assign n39498 = ~pi1147 & ~n39497;
  assign n39499 = ~n39495 & n39498;
  assign n39500 = pi1147 & ~n38425;
  assign n39501 = ~n38071 & n38426;
  assign n39502 = ~n38137 & n39501;
  assign n39503 = n39500 & ~n39502;
  assign n39504 = ~pi1150 & ~n39499;
  assign n39505 = ~n39503 & n39504;
  assign n39506 = n38383 & n38424;
  assign n39507 = pi1147 & ~n39506;
  assign n39508 = ~n38136 & n39501;
  assign n39509 = n39507 & ~n39508;
  assign n39510 = ~n39447 & n39496;
  assign n39511 = ~n38204 & n39494;
  assign n39512 = ~pi1147 & ~n39511;
  assign n39513 = ~n39510 & n39512;
  assign n39514 = pi1150 & ~n39509;
  assign n39515 = ~n39513 & n39514;
  assign n39516 = pi1149 & ~n39515;
  assign n39517 = ~n39505 & n39516;
  assign n39518 = ~pi1148 & ~n39492;
  assign n39519 = ~n39517 & n39518;
  assign n39520 = ~n39474 & ~n39519;
  assign n39521 = ~pi213 & ~n39520;
  assign n39522 = pi209 & ~n39404;
  assign n39523 = ~n39521 & n39522;
  assign n39524 = ~pi213 & n38191;
  assign n39525 = ~n38160 & ~n38317;
  assign n39526 = ~po1038 & ~n39525;
  assign n39527 = ~n38443 & ~n39526;
  assign n39528 = n39481 & n39527;
  assign n39529 = ~n39447 & n39494;
  assign n39530 = pi1147 & ~n38386;
  assign n39531 = ~n39529 & n39530;
  assign n39532 = ~pi1150 & ~n39528;
  assign n39533 = ~n39531 & n39532;
  assign n39534 = n38416 & ~n39448;
  assign n39535 = n38418 & n39449;
  assign n39536 = pi1147 & ~n39534;
  assign n39537 = ~n39535 & n39536;
  assign n39538 = ~n38300 & n38418;
  assign n39539 = n39465 & ~n39538;
  assign n39540 = pi1150 & ~n39537;
  assign n39541 = ~n39539 & n39540;
  assign n39542 = ~n39533 & ~n39541;
  assign n39543 = ~pi1149 & ~n39542;
  assign n39544 = ~pi1151 & n39476;
  assign n39545 = ~n38154 & n39544;
  assign n39546 = n39507 & ~n39545;
  assign n39547 = n38426 & ~n39484;
  assign n39548 = n38108 & ~n38313;
  assign n39549 = ~pi1147 & ~n39548;
  assign n39550 = ~n39547 & n39549;
  assign n39551 = ~pi1150 & ~n39546;
  assign n39552 = ~n39550 & n39551;
  assign n39553 = ~n38035 & ~n38401;
  assign n39554 = ~pi1151 & n39553;
  assign n39555 = n39443 & ~n39554;
  assign n39556 = n38517 & ~n39456;
  assign n39557 = ~n38153 & n38430;
  assign n39558 = ~n38144 & n39557;
  assign n39559 = ~pi1147 & ~n39558;
  assign n39560 = ~n39556 & n39559;
  assign n39561 = pi1150 & ~n39555;
  assign n39562 = ~n39560 & n39561;
  assign n39563 = ~n39552 & ~n39562;
  assign n39564 = pi1149 & ~n39563;
  assign n39565 = pi1148 & ~n39564;
  assign n39566 = ~n39543 & n39565;
  assign n39567 = ~n38088 & ~n38382;
  assign n39568 = ~n10332 & n37780;
  assign n39569 = n39567 & ~n39568;
  assign n39570 = n38424 & n39569;
  assign n39571 = ~pi1151 & ~n38088;
  assign n39572 = n39476 & n39571;
  assign n39573 = ~pi1147 & ~n39572;
  assign n39574 = ~n39570 & n39573;
  assign n39575 = ~n37783 & n38357;
  assign n39576 = ~n38106 & ~n39575;
  assign n39577 = ~n38103 & n39576;
  assign n39578 = n38426 & ~n39577;
  assign n39579 = n39500 & ~n39578;
  assign n39580 = ~pi1150 & ~n39574;
  assign n39581 = ~n39579 & n39580;
  assign n39582 = ~n38340 & n38517;
  assign n39583 = ~n39431 & n39557;
  assign n39584 = ~pi1147 & ~n39582;
  assign n39585 = ~n39583 & n39584;
  assign n39586 = ~n38035 & ~n39576;
  assign n39587 = ~pi1151 & n39586;
  assign n39588 = n39419 & ~n39587;
  assign n39589 = pi1150 & ~n39585;
  assign n39590 = ~n39588 & n39589;
  assign n39591 = ~n39581 & ~n39590;
  assign n39592 = pi1149 & ~n39591;
  assign n39593 = n38124 & n38353;
  assign n39594 = ~n38045 & ~n39593;
  assign n39595 = ~pi1151 & n39594;
  assign n39596 = n38418 & ~n39408;
  assign n39597 = pi1150 & ~n39596;
  assign n39598 = ~n39595 & n39597;
  assign n39599 = ~n38015 & ~n38366;
  assign n39600 = ~pi1151 & ~n39252;
  assign n39601 = ~pi1150 & ~n39600;
  assign n39602 = ~n39599 & n39601;
  assign n39603 = ~n39598 & ~n39602;
  assign n39604 = pi1147 & ~n39603;
  assign n39605 = ~n15574 & n37711;
  assign n39606 = pi1151 & ~n39605;
  assign n39607 = pi1150 & ~n39606;
  assign n39608 = n39429 & n39607;
  assign n39609 = ~pi1147 & n38414;
  assign n39610 = n38087 & n39609;
  assign n39611 = ~pi1149 & ~n39610;
  assign n39612 = ~n39608 & n39611;
  assign n39613 = ~n39604 & n39612;
  assign n39614 = ~pi1148 & ~n39613;
  assign n39615 = ~n39592 & n39614;
  assign n39616 = pi213 & ~n39566;
  assign n39617 = ~n39615 & n39616;
  assign n39618 = ~pi209 & ~n39524;
  assign n39619 = ~n39617 & n39618;
  assign n39620 = ~n39523 & ~n39619;
  assign n39621 = pi230 & ~n39620;
  assign n39622 = ~pi230 & pi247;
  assign po404 = n39621 | n39622;
  assign n39624 = ~pi213 & n39396;
  assign n39625 = pi1151 & ~pi1152;
  assign n39626 = n39427 & n39625;
  assign n39627 = ~pi1151 & ~n38087;
  assign n39628 = pi1152 & ~n39606;
  assign n39629 = ~n39627 & n39628;
  assign n39630 = ~pi1150 & ~n39626;
  assign n39631 = ~n39629 & n39630;
  assign n39632 = ~pi1152 & ~n39572;
  assign n39633 = ~n39435 & n39632;
  assign n39634 = n39501 & n39569;
  assign n39635 = pi1152 & ~n39634;
  assign n39636 = ~n39583 & n39635;
  assign n39637 = pi1150 & ~n39633;
  assign n39638 = ~n39636 & n39637;
  assign n39639 = ~n39631 & ~n39638;
  assign n39640 = ~pi1149 & ~n39639;
  assign n39641 = ~n38180 & n39430;
  assign n39642 = ~pi1152 & ~n39641;
  assign n39643 = ~n39480 & n39642;
  assign n39644 = ~pi1151 & ~n39527;
  assign n39645 = pi1152 & ~n39644;
  assign n39646 = ~n39538 & n39645;
  assign n39647 = ~n39643 & ~n39646;
  assign n39648 = ~pi1150 & ~n39647;
  assign n39649 = ~n38313 & n39501;
  assign n39650 = pi1152 & ~n39558;
  assign n39651 = ~n39649 & n39650;
  assign n39652 = ~pi1152 & ~n39457;
  assign n39653 = ~n39547 & n39652;
  assign n39654 = ~n39651 & ~n39653;
  assign n39655 = pi1150 & ~n39654;
  assign n39656 = pi1149 & ~n39655;
  assign n39657 = ~n39648 & n39656;
  assign n39658 = ~n39640 & ~n39657;
  assign n39659 = ~pi1148 & ~n39658;
  assign n39660 = pi1152 & ~n39497;
  assign n39661 = ~n39596 & n39660;
  assign n39662 = pi1151 & n39594;
  assign n39663 = ~pi1152 & ~n39600;
  assign n39664 = ~n39662 & n39663;
  assign n39665 = ~pi1150 & ~n39661;
  assign n39666 = ~n39664 & n39665;
  assign n39667 = pi1151 & n39586;
  assign n39668 = ~pi1152 & ~n39578;
  assign n39669 = ~n39667 & n39668;
  assign n39670 = ~n38107 & n39501;
  assign n39671 = pi1152 & ~n39670;
  assign n39672 = ~n39418 & n39671;
  assign n39673 = pi1150 & ~n39672;
  assign n39674 = ~n39669 & n39673;
  assign n39675 = ~pi1149 & ~n39666;
  assign n39676 = ~n39674 & n39675;
  assign n39677 = pi1151 & n39553;
  assign n39678 = ~pi1152 & ~n39545;
  assign n39679 = ~n39677 & n39678;
  assign n39680 = pi1152 & ~n38431;
  assign n39681 = n38383 & n39501;
  assign n39682 = n39680 & ~n39681;
  assign n39683 = pi1150 & ~n39679;
  assign n39684 = ~n39682 & n39683;
  assign n39685 = pi1152 & ~n39510;
  assign n39686 = ~n39535 & n39685;
  assign n39687 = n39430 & ~n39448;
  assign n39688 = n38387 & ~n39687;
  assign n39689 = ~pi1150 & ~n39688;
  assign n39690 = ~n39686 & n39689;
  assign n39691 = pi1149 & ~n39684;
  assign n39692 = ~n39690 & n39691;
  assign n39693 = pi1148 & ~n39692;
  assign n39694 = ~n39676 & n39693;
  assign n39695 = ~n39659 & ~n39694;
  assign n39696 = pi213 & ~n39695;
  assign n39697 = ~pi209 & ~n39624;
  assign n39698 = ~n39696 & n39697;
  assign n39699 = ~n38087 & n39571;
  assign n39700 = pi1152 & ~n39699;
  assign n39701 = ~n38419 & n39700;
  assign n39702 = ~n38181 & n39625;
  assign n39703 = ~pi1150 & ~n39701;
  assign n39704 = ~n39702 & n39703;
  assign n39705 = pi1151 & n38185;
  assign n39706 = ~pi1152 & ~n39705;
  assign n39707 = ~n38427 & n39706;
  assign n39708 = ~n39670 & n39680;
  assign n39709 = pi1150 & ~n39707;
  assign n39710 = ~n39708 & n39709;
  assign n39711 = ~n39704 & ~n39710;
  assign n39712 = pi213 & ~n39711;
  assign n39713 = n38254 & n39625;
  assign n39714 = pi1152 & ~n39571;
  assign n39715 = ~n39482 & n39714;
  assign n39716 = ~pi1150 & ~n39713;
  assign n39717 = ~n39715 & n39716;
  assign n39718 = ~pi1152 & ~n39497;
  assign n39719 = ~n39529 & n39718;
  assign n39720 = ~n39493 & n39496;
  assign n39721 = pi1152 & ~n39511;
  assign n39722 = ~n39720 & n39721;
  assign n39723 = pi1150 & ~n39719;
  assign n39724 = ~n39722 & n39723;
  assign n39725 = ~pi1148 & ~n39717;
  assign n39726 = ~n39724 & n39725;
  assign n39727 = ~n37729 & n39203;
  assign n39728 = ~pi1152 & ~n39544;
  assign n39729 = ~n39727 & n39728;
  assign n39730 = pi1152 & ~n39572;
  assign n39731 = ~n39485 & n39730;
  assign n39732 = ~pi1150 & ~n39729;
  assign n39733 = ~n39731 & n39732;
  assign n39734 = ~n39506 & n39671;
  assign n39735 = n38108 & ~n38136;
  assign n39736 = ~pi1152 & ~n39735;
  assign n39737 = ~n39502 & n39736;
  assign n39738 = pi1150 & ~n39737;
  assign n39739 = ~n39734 & n39738;
  assign n39740 = pi1148 & ~n39733;
  assign n39741 = ~n39739 & n39740;
  assign n39742 = ~pi1149 & ~n39726;
  assign n39743 = ~n39741 & n39742;
  assign n39744 = n38416 & ~n39431;
  assign n39745 = pi1152 & ~n39744;
  assign n39746 = ~n39467 & n39745;
  assign n39747 = ~n39428 & n39642;
  assign n39748 = ~pi1150 & ~n39746;
  assign n39749 = ~n39747 & n39748;
  assign n39750 = ~pi1151 & n39411;
  assign n39751 = pi1152 & ~n39451;
  assign n39752 = ~n39750 & n39751;
  assign n39753 = ~pi1152 & ~n39409;
  assign n39754 = ~n39535 & n39753;
  assign n39755 = pi1150 & ~n39752;
  assign n39756 = ~n39754 & n39755;
  assign n39757 = ~pi1148 & ~n39756;
  assign n39758 = ~n39749 & n39757;
  assign n39759 = pi1152 & ~n39582;
  assign n39760 = ~n39457 & n39759;
  assign n39761 = pi1151 & n39461;
  assign n39762 = ~pi1152 & ~n39436;
  assign n39763 = ~n39761 & n39762;
  assign n39764 = ~pi1150 & ~n39760;
  assign n39765 = ~n39763 & n39764;
  assign n39766 = ~n39417 & n39420;
  assign n39767 = n39680 & ~n39766;
  assign n39768 = ~n38134 & n39557;
  assign n39769 = ~pi1152 & ~n39768;
  assign n39770 = ~n39422 & n39769;
  assign n39771 = pi1150 & ~n39767;
  assign n39772 = ~n39770 & n39771;
  assign n39773 = pi1148 & ~n39772;
  assign n39774 = ~n39765 & n39773;
  assign n39775 = pi1149 & ~n39774;
  assign n39776 = ~n39758 & n39775;
  assign n39777 = ~n39743 & ~n39776;
  assign n39778 = ~pi213 & ~n39777;
  assign n39779 = pi209 & ~n39712;
  assign n39780 = ~n39778 & n39779;
  assign n39781 = ~n39698 & ~n39780;
  assign n39782 = pi230 & ~n39781;
  assign n39783 = ~pi230 & pi248;
  assign po405 = n39782 | n39783;
  assign n39785 = ~pi213 & ~n39711;
  assign n39786 = pi57 & ~n36875;
  assign n39787 = ~n6258 & n36875;
  assign n39788 = pi299 & n36872;
  assign n39789 = ~n38393 & ~n39788;
  assign n39790 = n37741 & n39789;
  assign n39791 = ~pi211 & n36547;
  assign n39792 = n37743 & ~n39791;
  assign n39793 = ~pi214 & ~n39789;
  assign n39794 = pi212 & ~n39792;
  assign n39795 = ~n39793 & n39794;
  assign n39796 = ~pi219 & ~n39790;
  assign n39797 = ~n39795 & n39796;
  assign n39798 = n6258 & ~n37615;
  assign n39799 = ~n39797 & n39798;
  assign n39800 = ~pi57 & pi1151;
  assign n39801 = ~n39787 & n39800;
  assign n39802 = ~n39799 & n39801;
  assign n39803 = ~n37734 & ~n39788;
  assign n39804 = ~pi212 & ~n39803;
  assign n39805 = n36580 & ~n36871;
  assign n39806 = n10332 & n37713;
  assign n39807 = ~n39805 & ~n39806;
  assign n39808 = pi299 & ~n39807;
  assign n39809 = ~n38380 & ~n39808;
  assign n39810 = ~n38122 & n39809;
  assign n39811 = ~n39804 & n39810;
  assign n39812 = ~pi219 & ~n39811;
  assign n39813 = n6258 & ~n38258;
  assign n39814 = ~n39812 & n39813;
  assign n39815 = ~pi57 & ~pi1151;
  assign n39816 = ~n39787 & n39815;
  assign n39817 = ~n39814 & n39816;
  assign n39818 = ~n39786 & ~n39802;
  assign n39819 = ~n39817 & n39818;
  assign n39820 = ~pi1152 & ~n39819;
  assign n39821 = pi299 & ~n36872;
  assign n39822 = ~n10332 & n39821;
  assign n39823 = ~n36925 & ~n39822;
  assign n39824 = n37352 & ~n39823;
  assign n39825 = n38377 & ~n39824;
  assign n39826 = ~n37812 & ~n38197;
  assign n39827 = pi1151 & ~n39826;
  assign n39828 = ~n39825 & n39827;
  assign n39829 = n38336 & ~n39788;
  assign n39830 = ~n37150 & n39805;
  assign n39831 = n38093 & ~n38369;
  assign n39832 = n38479 & ~n39830;
  assign n39833 = ~n39831 & n39832;
  assign n39834 = n39242 & ~n39829;
  assign n39835 = ~n39833 & n39834;
  assign n39836 = ~pi1151 & ~n38106;
  assign n39837 = ~n39835 & n39836;
  assign n39838 = n36930 & ~n39828;
  assign n39839 = ~n39837 & n39838;
  assign n39840 = ~n39820 & ~n39839;
  assign n39841 = pi1150 & ~n39840;
  assign n39842 = ~n39791 & ~n39822;
  assign n39843 = n36874 & n37587;
  assign n39844 = ~n39842 & n39843;
  assign n39845 = n38292 & ~n39821;
  assign n39846 = pi212 & ~n39845;
  assign n39847 = ~n38294 & n39846;
  assign n39848 = ~pi212 & ~n37045;
  assign n39849 = ~pi219 & ~n39829;
  assign n39850 = ~n39848 & n39849;
  assign n39851 = ~n39847 & n39850;
  assign n39852 = pi1151 & n38209;
  assign n39853 = ~n39851 & n39852;
  assign n39854 = ~pi1151 & ~n39567;
  assign n39855 = n36930 & ~n39854;
  assign n39856 = ~n39853 & n39855;
  assign n39857 = n37059 & ~n37572;
  assign n39858 = n37049 & ~n38316;
  assign n39859 = ~n38160 & ~n39788;
  assign n39860 = n36675 & ~n39859;
  assign n39861 = ~n39857 & ~n39858;
  assign n39862 = ~n39860 & n39861;
  assign n39863 = ~pi219 & ~n39862;
  assign n39864 = pi1151 & n38179;
  assign n39865 = ~n39863 & n39864;
  assign n39866 = n36877 & ~n39865;
  assign n39867 = ~n39856 & ~n39866;
  assign n39868 = ~pi1150 & ~n39844;
  assign n39869 = ~n39867 & n39868;
  assign n39870 = ~n39841 & ~n39869;
  assign n39871 = pi213 & ~n39870;
  assign n39872 = ~pi209 & ~n39785;
  assign n39873 = ~n39871 & n39872;
  assign n39874 = pi213 & ~n37064;
  assign n39875 = pi212 & n36790;
  assign n39876 = n37045 & ~n39875;
  assign n39877 = ~n37038 & ~n39876;
  assign n39878 = n38175 & ~n39877;
  assign n39879 = n37048 & ~n39878;
  assign n39880 = n39430 & ~n39879;
  assign n39881 = n37046 & n37066;
  assign n39882 = ~n39625 & ~n39881;
  assign n39883 = ~n39880 & ~n39882;
  assign n39884 = ~n36997 & n37756;
  assign n39885 = ~n36980 & ~n37756;
  assign n39886 = ~po1038 & ~n39885;
  assign n39887 = ~n39884 & n39886;
  assign n39888 = n39496 & ~n39887;
  assign n39889 = pi214 & n36995;
  assign n39890 = n37022 & ~n39889;
  assign n39891 = ~pi219 & ~n39890;
  assign n39892 = pi214 & ~n36997;
  assign n39893 = ~pi214 & n36995;
  assign n39894 = pi212 & ~n39893;
  assign n39895 = ~n39892 & n39894;
  assign n39896 = n39891 & ~n39895;
  assign n39897 = ~po1038 & ~n37000;
  assign n39898 = ~n39896 & n39897;
  assign n39899 = n38418 & ~n39898;
  assign n39900 = pi1152 & ~n39888;
  assign n39901 = ~n39899 & n39900;
  assign n39902 = ~pi1150 & ~n39883;
  assign n39903 = ~n39901 & n39902;
  assign n39904 = n39434 & ~n39879;
  assign n39905 = ~n38426 & ~n39904;
  assign n39906 = ~n37038 & n38152;
  assign n39907 = ~n37048 & ~n39906;
  assign n39908 = ~n37046 & n38381;
  assign n39909 = ~n39907 & ~n39908;
  assign n39910 = ~n39905 & ~n39909;
  assign n39911 = ~pi1152 & ~n39910;
  assign n39912 = pi212 & ~n36995;
  assign n39913 = n39891 & ~n39912;
  assign n39914 = n37003 & ~n39913;
  assign n39915 = n38430 & ~n39914;
  assign n39916 = ~n37021 & ~n39892;
  assign n39917 = ~pi212 & ~n39916;
  assign n39918 = ~pi211 & n36980;
  assign n39919 = ~n37004 & ~n39918;
  assign n39920 = pi214 & ~n39919;
  assign n39921 = ~pi214 & n36997;
  assign n39922 = pi212 & ~n39920;
  assign n39923 = ~n39921 & n39922;
  assign n39924 = ~n39917 & ~n39923;
  assign n39925 = ~pi219 & ~n39924;
  assign n39926 = n37003 & ~n39925;
  assign n39927 = n39501 & ~n39926;
  assign n39928 = pi1152 & ~n39915;
  assign n39929 = ~n39927 & n39928;
  assign n39930 = pi1150 & ~n39911;
  assign n39931 = ~n39929 & n39930;
  assign n39932 = ~n39903 & ~n39931;
  assign n39933 = ~pi213 & ~n39932;
  assign n39934 = pi209 & ~n39874;
  assign n39935 = ~n39933 & n39934;
  assign n39936 = ~n39873 & ~n39935;
  assign n39937 = pi230 & ~n39936;
  assign n39938 = ~pi230 & pi249;
  assign po406 = n39937 | n39938;
  assign n39940 = n2532 & n11103;
  assign n39941 = ~n6083 & ~n39940;
  assign n39942 = ~pi75 & ~n39941;
  assign n39943 = n7236 & n8670;
  assign n39944 = ~n39942 & ~n39943;
  assign n39945 = ~pi87 & ~pi250;
  assign n39946 = n8598 & n39945;
  assign po407 = ~n39944 & n39946;
  assign n39948 = pi897 & n10421;
  assign n39949 = ~pi476 & n11035;
  assign n39950 = ~n39948 & ~n39949;
  assign n39951 = ~pi200 & pi1053;
  assign n39952 = pi200 & pi1039;
  assign n39953 = ~pi199 & ~n39951;
  assign n39954 = ~n39952 & n39953;
  assign n39955 = ~n39950 & ~n39954;
  assign n39956 = pi251 & n39950;
  assign po408 = n39955 | n39956;
  assign n39958 = ~n10585 & n11143;
  assign n39959 = ~n6205 & n11143;
  assign n39960 = ~pi979 & ~pi984;
  assign n39961 = pi1001 & n39960;
  assign n39962 = n6172 & n39961;
  assign n39963 = ~n6103 & n39962;
  assign n39964 = n6333 & n39963;
  assign n39965 = ~pi252 & ~n39964;
  assign n39966 = pi1092 & ~pi1093;
  assign n39967 = ~n39965 & n39966;
  assign n39968 = n6349 & ~n39967;
  assign n39969 = n6348 & n39967;
  assign n39970 = ~n39968 & ~n39969;
  assign n39971 = n6205 & n39970;
  assign n39972 = ~n39959 & ~n39971;
  assign n39973 = n6221 & ~n39972;
  assign n39974 = ~n6197 & n39970;
  assign n39975 = n6197 & n11143;
  assign n39976 = ~n39974 & ~n39975;
  assign n39977 = ~n6221 & ~n39976;
  assign n39978 = pi299 & ~n39973;
  assign n39979 = ~n39977 & n39978;
  assign n39980 = n6194 & ~n39972;
  assign n39981 = ~n6194 & ~n39976;
  assign n39982 = ~pi299 & ~n39980;
  assign n39983 = ~n39981 & n39982;
  assign n39984 = n10585 & ~n39979;
  assign n39985 = ~n39983 & n39984;
  assign n39986 = ~n7578 & ~n39958;
  assign n39987 = ~n39985 & n39986;
  assign n39988 = pi57 & n11142;
  assign n39989 = n10584 & n39962;
  assign n39990 = n20005 & n39989;
  assign n39991 = n6180 & n39990;
  assign n39992 = ~n11007 & n39991;
  assign n39993 = n6333 & n39992;
  assign n39994 = ~pi252 & ~n39993;
  assign n39995 = ~pi57 & pi1092;
  assign n39996 = ~n39994 & n39995;
  assign n39997 = n7578 & ~n39988;
  assign n39998 = ~n39996 & n39997;
  assign po409 = ~n39987 & ~n39998;
  assign n40000 = ~pi1151 & n10333;
  assign n40001 = ~n37231 & ~n40000;
  assign n40002 = pi1153 & ~n36619;
  assign n40003 = ~n37609 & n40002;
  assign n40004 = ~n10970 & ~n36572;
  assign n40005 = pi1151 & n40004;
  assign n40006 = ~n40003 & n40005;
  assign n40007 = n36554 & n37676;
  assign n40008 = ~pi1151 & ~n11038;
  assign n40009 = ~n36736 & n40008;
  assign n40010 = ~n40007 & n40009;
  assign n40011 = ~po1038 & ~n40006;
  assign n40012 = ~n40010 & n40011;
  assign n40013 = pi1152 & ~n40001;
  assign n40014 = ~n40012 & n40013;
  assign n40015 = ~n36572 & ~n37609;
  assign n40016 = ~n36743 & n40015;
  assign n40017 = ~po1038 & n40016;
  assign n40018 = po1038 & n36554;
  assign n40019 = ~n40017 & ~n40018;
  assign n40020 = ~pi1151 & pi1153;
  assign n40021 = ~n40019 & n40020;
  assign n40022 = ~n11037 & ~n37231;
  assign n40023 = pi211 & ~n36612;
  assign n40024 = n10333 & ~n40002;
  assign n40025 = ~n36975 & n40024;
  assign n40026 = ~n40023 & ~n40025;
  assign n40027 = ~n36604 & ~n36619;
  assign n40028 = n36554 & ~n40027;
  assign n40029 = ~po1038 & ~n40028;
  assign n40030 = n40026 & n40029;
  assign n40031 = ~n40022 & ~n40030;
  assign n40032 = pi1151 & ~n40031;
  assign n40033 = ~pi1152 & ~n40021;
  assign n40034 = ~n40032 & n40033;
  assign n40035 = ~n40014 & ~n40034;
  assign n40036 = pi230 & ~n40035;
  assign n40037 = pi253 & po1038;
  assign n40038 = pi219 & pi1091;
  assign n40039 = ~n36581 & n40038;
  assign n40040 = ~pi219 & ~n38721;
  assign n40041 = ~pi211 & ~n38718;
  assign n40042 = pi219 & ~n38707;
  assign n40043 = ~n40041 & n40042;
  assign n40044 = po1038 & ~n40043;
  assign n40045 = ~n40040 & n40044;
  assign n40046 = ~n40039 & n40045;
  assign n40047 = ~n40037 & ~n40046;
  assign n40048 = ~pi219 & ~n38722;
  assign n40049 = ~n38707 & ~n40039;
  assign n40050 = ~n40048 & n40049;
  assign n40051 = pi253 & ~n40050;
  assign n40052 = ~n40047 & ~n40051;
  assign n40053 = ~pi211 & ~n38721;
  assign n40054 = n40048 & ~n40053;
  assign n40055 = ~pi219 & ~n40054;
  assign n40056 = po1038 & n40055;
  assign n40057 = ~n38718 & n40056;
  assign n40058 = pi1151 & ~n40057;
  assign n40059 = ~n40052 & n40058;
  assign n40060 = ~n38734 & n38755;
  assign n40061 = ~pi211 & n40060;
  assign n40062 = ~n38783 & ~n40061;
  assign n40063 = pi1153 & ~n40062;
  assign n40064 = ~n38758 & ~n40063;
  assign n40065 = pi219 & ~n40064;
  assign n40066 = ~n38813 & ~n40061;
  assign n40067 = n40048 & ~n40066;
  assign n40068 = pi1153 & n38796;
  assign n40069 = ~pi219 & ~n38750;
  assign n40070 = ~n40068 & n40069;
  assign n40071 = n40067 & ~n40070;
  assign n40072 = ~n40065 & ~n40071;
  assign n40073 = ~n38734 & ~n40072;
  assign n40074 = ~pi253 & ~n40073;
  assign n40075 = ~n38741 & ~n38749;
  assign n40076 = ~pi211 & n38812;
  assign n40077 = n40075 & ~n40076;
  assign n40078 = n40048 & n40077;
  assign n40079 = pi1153 & ~n38767;
  assign n40080 = n40078 & ~n40079;
  assign n40081 = n38772 & ~n38779;
  assign n40082 = n40077 & n40081;
  assign n40083 = ~n38799 & ~n40082;
  assign n40084 = pi1153 & n40083;
  assign n40085 = pi219 & n38743;
  assign n40086 = ~n40084 & n40085;
  assign n40087 = ~n40080 & ~n40086;
  assign n40088 = pi253 & ~n40087;
  assign n40089 = ~po1038 & ~n40088;
  assign n40090 = ~n40074 & n40089;
  assign n40091 = ~pi1152 & n40059;
  assign n40092 = ~n40090 & n40091;
  assign n40093 = n40040 & ~n40041;
  assign n40094 = n40048 & ~n40093;
  assign n40095 = pi219 & ~n38718;
  assign n40096 = po1038 & ~n40095;
  assign n40097 = ~n40094 & n40096;
  assign n40098 = pi1091 & n40097;
  assign n40099 = pi219 & n40064;
  assign n40100 = ~pi253 & ~n40070;
  assign n40101 = ~n40099 & n40100;
  assign n40102 = ~n38812 & n38832;
  assign n40103 = ~n38772 & ~n40102;
  assign n40104 = ~pi1153 & n40103;
  assign n40105 = ~n38832 & ~n40104;
  assign n40106 = ~pi219 & n38854;
  assign n40107 = ~n40105 & n40106;
  assign n40108 = pi1153 & ~n40082;
  assign n40109 = ~pi1153 & ~n38755;
  assign n40110 = pi219 & ~n40109;
  assign n40111 = ~n40108 & n40110;
  assign n40112 = pi253 & ~n40111;
  assign n40113 = ~n40107 & n40112;
  assign n40114 = ~n40101 & ~n40113;
  assign n40115 = ~po1038 & ~n40114;
  assign n40116 = n40059 & ~n40115;
  assign n40117 = ~n38782 & n40078;
  assign n40118 = ~n40104 & n40117;
  assign n40119 = ~n38741 & n40065;
  assign n40120 = ~n40118 & ~n40119;
  assign n40121 = ~pi253 & ~n40120;
  assign n40122 = pi219 & n38780;
  assign n40123 = ~n40084 & n40122;
  assign n40124 = n40067 & ~n40105;
  assign n40125 = pi253 & ~n40123;
  assign n40126 = ~n40124 & n40125;
  assign n40127 = ~n40121 & ~n40126;
  assign n40128 = ~po1038 & ~n40127;
  assign n40129 = ~pi1151 & ~n40128;
  assign n40130 = ~n40116 & ~n40129;
  assign n40131 = pi1152 & ~n40098;
  assign n40132 = ~n40130 & n40131;
  assign n40133 = pi219 & ~n38754;
  assign n40134 = ~n38734 & n38854;
  assign n40135 = ~n40133 & ~n40134;
  assign n40136 = n40101 & ~n40135;
  assign n40137 = ~pi1091 & ~n38758;
  assign n40138 = ~pi1153 & ~n40137;
  assign n40139 = ~pi219 & ~n40103;
  assign n40140 = pi253 & ~n40138;
  assign n40141 = n40083 & n40140;
  assign n40142 = ~n40139 & n40141;
  assign n40143 = ~n40136 & ~n40142;
  assign n40144 = ~po1038 & ~n40143;
  assign n40145 = ~pi1151 & ~pi1152;
  assign n40146 = ~n40144 & n40145;
  assign n40147 = ~n40132 & ~n40146;
  assign n40148 = ~n40052 & ~n40147;
  assign n40149 = n38687 & ~n40092;
  assign n40150 = ~n40148 & n40149;
  assign n40151 = ~pi253 & ~pi1091;
  assign n40152 = po1038 & ~n40151;
  assign n40153 = ~n40039 & n40152;
  assign n40154 = pi1091 & n40000;
  assign n40155 = n40153 & ~n40154;
  assign n40156 = pi1091 & n36736;
  assign n40157 = pi253 & ~pi1091;
  assign n40158 = ~n11037 & ~n36554;
  assign n40159 = ~n40157 & n40158;
  assign n40160 = pi211 & ~pi253;
  assign n40161 = ~n38670 & n40160;
  assign n40162 = ~n40159 & ~n40161;
  assign n40163 = ~n40156 & ~n40162;
  assign n40164 = n11037 & n38641;
  assign n40165 = ~n36736 & n40164;
  assign n40166 = pi1091 & n36554;
  assign n40167 = n36624 & n40166;
  assign n40168 = ~n37666 & ~n40167;
  assign n40169 = n38638 & ~n40168;
  assign n40170 = pi253 & ~n40165;
  assign n40171 = ~n40169 & n40170;
  assign n40172 = n36969 & n38621;
  assign n40173 = pi1091 & pi1153;
  assign n40174 = ~n36624 & n40173;
  assign n40175 = n36554 & ~n40172;
  assign n40176 = ~n40174 & n40175;
  assign n40177 = ~pi253 & ~n40176;
  assign n40178 = ~n40171 & ~n40177;
  assign n40179 = n37587 & ~n40163;
  assign n40180 = ~n40178 & n40179;
  assign n40181 = pi1091 & ~pi1153;
  assign n40182 = ~n12342 & ~n36610;
  assign n40183 = ~n40157 & n40182;
  assign n40184 = ~n40181 & ~n40183;
  assign n40185 = n40004 & ~n40184;
  assign n40186 = n37617 & ~n40151;
  assign n40187 = ~n40185 & n40186;
  assign n40188 = pi1152 & ~n40155;
  assign n40189 = ~n40187 & n40188;
  assign n40190 = ~n40180 & n40189;
  assign n40191 = n40017 & n40173;
  assign n40192 = pi219 & n40153;
  assign n40193 = ~pi1151 & ~n40157;
  assign n40194 = ~n40191 & n40193;
  assign n40195 = ~n40192 & n40194;
  assign n40196 = n12344 & ~n40003;
  assign n40197 = pi1091 & ~n40196;
  assign n40198 = ~pi253 & ~n40197;
  assign n40199 = ~n36967 & ~n38621;
  assign n40200 = n36554 & ~n40199;
  assign n40201 = n40026 & ~n40200;
  assign n40202 = pi253 & pi1091;
  assign n40203 = ~n40201 & n40202;
  assign n40204 = ~po1038 & ~n40198;
  assign n40205 = ~n40203 & n40204;
  assign n40206 = pi219 & n40181;
  assign n40207 = pi211 & pi1091;
  assign n40208 = ~n40206 & ~n40207;
  assign n40209 = n40152 & n40208;
  assign n40210 = pi1151 & ~n40209;
  assign n40211 = ~n40205 & n40210;
  assign n40212 = ~n40195 & ~n40211;
  assign n40213 = ~pi1152 & ~n40212;
  assign n40214 = ~n38687 & ~n40190;
  assign n40215 = ~n40213 & n40214;
  assign n40216 = ~pi230 & ~n40215;
  assign n40217 = ~n40150 & n40216;
  assign po410 = ~n40036 & ~n40217;
  assign n40219 = ~pi219 & ~n36871;
  assign n40220 = ~n37116 & ~n40219;
  assign n40221 = po1038 & n40220;
  assign n40222 = pi299 & n36554;
  assign n40223 = ~n11037 & n36970;
  assign n40224 = ~n40222 & ~n40223;
  assign n40225 = ~n37189 & ~n40224;
  assign n40226 = n36654 & ~n36880;
  assign n40227 = n11037 & ~n37005;
  assign n40228 = ~n40226 & n40227;
  assign n40229 = ~n40225 & ~n40228;
  assign n40230 = ~po1038 & ~n40229;
  assign n40231 = ~pi1152 & ~n40221;
  assign n40232 = ~n40230 & n40231;
  assign n40233 = n11037 & ~n36871;
  assign n40234 = n37853 & ~n40233;
  assign n40235 = ~pi200 & pi1154;
  assign n40236 = n10957 & ~n40235;
  assign n40237 = ~n12342 & n37005;
  assign n40238 = ~n40236 & ~n40237;
  assign n40239 = ~pi219 & ~n40238;
  assign n40240 = ~n36599 & ~n37005;
  assign n40241 = n36562 & ~n40240;
  assign n40242 = n36989 & ~n37191;
  assign n40243 = ~n40241 & ~n40242;
  assign n40244 = pi219 & ~n40243;
  assign n40245 = ~po1038 & ~n40239;
  assign n40246 = ~n40244 & n40245;
  assign n40247 = pi1152 & ~n40234;
  assign n40248 = ~n40246 & n40247;
  assign n40249 = ~n40232 & ~n40248;
  assign n40250 = pi230 & ~n40249;
  assign n40251 = pi1091 & ~n40220;
  assign n40252 = ~pi254 & ~pi1091;
  assign n40253 = po1038 & ~n40252;
  assign n40254 = ~n40251 & n40253;
  assign n40255 = pi1091 & n38014;
  assign n40256 = ~n40254 & ~n40255;
  assign n40257 = ~pi1153 & ~n38648;
  assign n40258 = pi1153 & ~n38635;
  assign n40259 = ~pi1154 & ~n40258;
  assign n40260 = ~n37769 & ~n40257;
  assign n40261 = n40259 & n40260;
  assign n40262 = pi1153 & ~n10957;
  assign n40263 = pi1091 & n36562;
  assign n40264 = ~n36610 & n40263;
  assign n40265 = ~n40262 & n40264;
  assign n40266 = ~n40261 & ~n40265;
  assign n40267 = ~pi219 & ~n40266;
  assign n40268 = ~pi211 & pi1091;
  assign n40269 = pi1154 & n40268;
  assign n40270 = ~n40038 & ~n40269;
  assign n40271 = ~n40243 & ~n40270;
  assign n40272 = ~n40267 & ~n40271;
  assign n40273 = pi254 & ~n40272;
  assign n40274 = n36988 & ~n37609;
  assign n40275 = pi219 & ~n37191;
  assign n40276 = ~n40274 & n40275;
  assign n40277 = ~n40239 & ~n40276;
  assign n40278 = ~pi254 & ~n40277;
  assign n40279 = ~n40252 & ~n40278;
  assign n40280 = ~n40273 & n40279;
  assign n40281 = ~po1038 & n40280;
  assign n40282 = pi1152 & n40256;
  assign n40283 = ~n40281 & n40282;
  assign n40284 = ~n37676 & n38623;
  assign n40285 = n40207 & ~n40259;
  assign n40286 = ~n40284 & n40285;
  assign n40287 = pi1091 & n36970;
  assign n40288 = n11036 & n40173;
  assign n40289 = ~pi1154 & ~n40288;
  assign n40290 = ~pi211 & ~n40289;
  assign n40291 = n40287 & n40290;
  assign n40292 = ~n40286 & ~n40291;
  assign n40293 = ~pi219 & ~n40292;
  assign n40294 = ~pi1153 & ~n36743;
  assign n40295 = ~n37676 & ~n40294;
  assign n40296 = pi1091 & ~n40295;
  assign n40297 = n36579 & ~n40296;
  assign n40298 = n36562 & ~n40287;
  assign n40299 = pi219 & ~n40289;
  assign n40300 = ~n40298 & n40299;
  assign n40301 = ~n40297 & n40300;
  assign n40302 = ~n40293 & ~n40301;
  assign n40303 = ~pi254 & ~n40302;
  assign n40304 = ~pi1154 & n38659;
  assign n40305 = ~n40284 & ~n40304;
  assign n40306 = n11037 & ~n40305;
  assign n40307 = pi1091 & ~n11037;
  assign n40308 = ~n36987 & n40307;
  assign n40309 = ~pi1154 & ~n40308;
  assign n40310 = n38673 & ~n40168;
  assign n40311 = pi1091 & ~n36707;
  assign n40312 = ~n40284 & ~n40311;
  assign n40313 = n40158 & ~n40312;
  assign n40314 = pi1154 & ~n40310;
  assign n40315 = ~n40313 & n40314;
  assign n40316 = ~n40309 & ~n40315;
  assign n40317 = pi254 & ~n40306;
  assign n40318 = ~n40316 & n40317;
  assign n40319 = ~n40303 & ~n40318;
  assign n40320 = ~po1038 & ~n40319;
  assign n40321 = ~pi1152 & ~n40254;
  assign n40322 = ~n40320 & n40321;
  assign n40323 = ~n38687 & ~n40283;
  assign n40324 = ~n40322 & n40323;
  assign n40325 = pi1091 & n37116;
  assign n40326 = ~pi211 & ~n38705;
  assign n40327 = n40095 & ~n40326;
  assign n40328 = ~pi219 & n38721;
  assign n40329 = ~n40327 & ~n40328;
  assign n40330 = n11037 & n40181;
  assign n40331 = pi254 & ~n40330;
  assign n40332 = ~n40325 & n40331;
  assign n40333 = n40329 & n40332;
  assign n40334 = n40093 & ~n40173;
  assign n40335 = ~pi254 & ~n40325;
  assign n40336 = ~n40043 & n40335;
  assign n40337 = ~n40334 & n40336;
  assign n40338 = pi253 & ~n40333;
  assign n40339 = ~n40337 & n40338;
  assign n40340 = ~n40037 & n40256;
  assign n40341 = ~n40339 & ~n40340;
  assign n40342 = ~pi253 & ~n40280;
  assign n40343 = n38743 & ~n38782;
  assign n40344 = pi1154 & n40343;
  assign n40345 = ~n38750 & ~n40344;
  assign n40346 = ~n38871 & ~n40076;
  assign n40347 = ~pi1153 & n40346;
  assign n40348 = ~n40345 & ~n40347;
  assign n40349 = ~pi254 & ~n40348;
  assign n40350 = pi1153 & ~n38813;
  assign n40351 = ~n38740 & ~n40350;
  assign n40352 = pi1154 & ~n40351;
  assign n40353 = ~pi1153 & n38772;
  assign n40354 = n40066 & ~n40353;
  assign n40355 = ~pi1154 & n40354;
  assign n40356 = pi254 & n40077;
  assign n40357 = ~n40352 & n40356;
  assign n40358 = ~n40355 & n40357;
  assign n40359 = ~pi219 & ~n40349;
  assign n40360 = ~n40358 & n40359;
  assign n40361 = ~n38807 & ~n40082;
  assign n40362 = pi1154 & ~n40108;
  assign n40363 = ~n40361 & n40362;
  assign n40364 = pi1153 & ~n38755;
  assign n40365 = ~pi1154 & n38743;
  assign n40366 = ~n40364 & n40365;
  assign n40367 = ~n40363 & ~n40366;
  assign n40368 = pi254 & ~n40367;
  assign n40369 = ~n40109 & n40343;
  assign n40370 = n36579 & ~n40369;
  assign n40371 = ~pi1153 & ~n38727;
  assign n40372 = n38760 & ~n40371;
  assign n40373 = ~pi1154 & ~n40372;
  assign n40374 = n38784 & ~n40109;
  assign n40375 = n36562 & ~n40374;
  assign n40376 = ~n40370 & ~n40373;
  assign n40377 = ~n40375 & n40376;
  assign n40378 = ~n38734 & n38758;
  assign n40379 = ~pi254 & ~n40378;
  assign n40380 = ~n40377 & n40379;
  assign n40381 = pi219 & ~n40380;
  assign n40382 = ~n40368 & n40381;
  assign n40383 = pi253 & ~n40360;
  assign n40384 = ~n40382 & n40383;
  assign n40385 = ~po1038 & ~n40342;
  assign n40386 = ~n40384 & n40385;
  assign n40387 = pi1152 & ~n40341;
  assign n40388 = ~n40386 & n40387;
  assign n40389 = ~n40037 & ~n40254;
  assign n40390 = ~n40094 & n40333;
  assign n40391 = ~n40055 & n40337;
  assign n40392 = pi253 & ~n40390;
  assign n40393 = ~n40391 & n40392;
  assign n40394 = ~n40389 & ~n40393;
  assign n40395 = ~pi253 & n40319;
  assign n40396 = pi219 & ~n40377;
  assign n40397 = pi1154 & n38771;
  assign n40398 = ~n40354 & ~n40397;
  assign n40399 = ~n38718 & ~n40398;
  assign n40400 = ~pi219 & ~n38852;
  assign n40401 = ~n40399 & n40400;
  assign n40402 = ~n40396 & ~n40401;
  assign n40403 = ~pi254 & ~n40402;
  assign n40404 = ~pi219 & ~n40398;
  assign n40405 = ~n38780 & ~n40138;
  assign n40406 = n36579 & ~n38799;
  assign n40407 = ~n40397 & ~n40406;
  assign n40408 = ~n40405 & n40407;
  assign n40409 = pi219 & ~n40408;
  assign n40410 = pi254 & ~n40409;
  assign n40411 = ~n40404 & n40410;
  assign n40412 = ~n40403 & ~n40411;
  assign n40413 = pi253 & ~n40412;
  assign n40414 = ~po1038 & ~n40395;
  assign n40415 = ~n40413 & n40414;
  assign n40416 = ~pi1152 & ~n40394;
  assign n40417 = ~n40415 & n40416;
  assign n40418 = n38687 & ~n40388;
  assign n40419 = ~n40417 & n40418;
  assign n40420 = ~pi230 & ~n40324;
  assign n40421 = ~n40419 & n40420;
  assign po411 = ~n40250 & ~n40421;
  assign n40423 = pi200 & ~pi1036;
  assign n40424 = ~pi200 & ~pi1049;
  assign n40425 = ~n40423 & ~n40424;
  assign n40426 = ~n39950 & n40425;
  assign n40427 = pi255 & n39950;
  assign po412 = n40426 | n40427;
  assign n40429 = pi200 & ~pi1070;
  assign n40430 = ~pi200 & ~pi1048;
  assign n40431 = ~n40429 & ~n40430;
  assign n40432 = ~n39950 & n40431;
  assign n40433 = pi256 & n39950;
  assign po413 = n40432 | n40433;
  assign n40435 = pi200 & ~pi1065;
  assign n40436 = ~pi200 & ~pi1084;
  assign n40437 = ~n40435 & ~n40436;
  assign n40438 = ~n39950 & n40437;
  assign n40439 = pi257 & n39950;
  assign po414 = n40438 | n40439;
  assign n40441 = pi200 & ~pi1062;
  assign n40442 = ~pi200 & ~pi1072;
  assign n40443 = ~n40441 & ~n40442;
  assign n40444 = ~n39950 & n40443;
  assign n40445 = pi258 & n39950;
  assign po415 = n40444 | n40445;
  assign n40447 = pi200 & ~pi1069;
  assign n40448 = ~pi200 & ~pi1059;
  assign n40449 = ~n40447 & ~n40448;
  assign n40450 = ~n39950 & n40449;
  assign n40451 = pi259 & n39950;
  assign po416 = n40450 | n40451;
  assign n40453 = ~pi200 & pi1044;
  assign n40454 = pi200 & pi1067;
  assign n40455 = ~pi199 & ~n40453;
  assign n40456 = ~n40454 & n40455;
  assign n40457 = ~n39950 & ~n40456;
  assign n40458 = pi260 & n39950;
  assign po417 = n40457 | n40458;
  assign n40460 = ~pi200 & pi1037;
  assign n40461 = pi200 & pi1040;
  assign n40462 = ~pi199 & ~n40460;
  assign n40463 = ~n40461 & n40462;
  assign n40464 = ~n39950 & ~n40463;
  assign n40465 = pi261 & n39950;
  assign po418 = n40464 | n40465;
  assign n40467 = ~pi123 & pi228;
  assign n40468 = ~pi228 & pi1093;
  assign n40469 = ~n40467 & ~n40468;
  assign n40470 = pi199 & ~n40469;
  assign n40471 = pi1093 & pi1142;
  assign n40472 = ~pi262 & ~pi1093;
  assign n40473 = ~n40471 & ~n40472;
  assign n40474 = ~pi228 & ~n40473;
  assign n40475 = ~pi123 & ~pi1142;
  assign n40476 = pi123 & pi262;
  assign n40477 = pi228 & ~n40475;
  assign n40478 = ~n40476 & n40477;
  assign n40479 = ~n40474 & ~n40478;
  assign n40480 = n37039 & ~n40469;
  assign n40481 = ~n40479 & ~n40480;
  assign n40482 = pi208 & ~n40481;
  assign n40483 = ~n40470 & ~n40482;
  assign n40484 = ~pi299 & ~n40483;
  assign n40485 = ~pi262 & n40469;
  assign n40486 = ~n37149 & ~n40485;
  assign n40487 = ~n38146 & n40486;
  assign n40488 = ~n36522 & ~n38146;
  assign n40489 = n40479 & ~n40488;
  assign n40490 = ~po1038 & ~n40487;
  assign n40491 = ~n40489 & n40490;
  assign n40492 = ~n40484 & n40491;
  assign n40493 = ~n37711 & ~n40469;
  assign n40494 = po1038 & ~n40479;
  assign n40495 = ~n40493 & n40494;
  assign po419 = n40492 | n40495;
  assign n40497 = ~pi199 & ~pi1154;
  assign n40498 = n36610 & ~n40497;
  assign n40499 = n40207 & ~n40498;
  assign n40500 = ~n36826 & n40499;
  assign n40501 = pi1155 & ~n36974;
  assign n40502 = n38621 & ~n40501;
  assign n40503 = ~pi1154 & n40311;
  assign n40504 = ~n40502 & ~n40503;
  assign n40505 = ~pi211 & ~n40504;
  assign n40506 = pi1156 & ~n40500;
  assign n40507 = ~n40505 & n40506;
  assign n40508 = ~n36620 & ~n37029;
  assign n40509 = n40268 & n40508;
  assign n40510 = pi1091 & ~pi1154;
  assign n40511 = ~n38648 & ~n40510;
  assign n40512 = ~n36826 & ~n40511;
  assign n40513 = pi211 & n40512;
  assign n40514 = ~pi1156 & ~n40509;
  assign n40515 = ~n40513 & n40514;
  assign n40516 = ~n40507 & ~n40515;
  assign n40517 = ~pi219 & ~n40516;
  assign n40518 = pi1154 & ~n36636;
  assign n40519 = pi1156 & ~n40518;
  assign n40520 = n40268 & n40519;
  assign n40521 = n36745 & n40520;
  assign n40522 = ~n38670 & n40504;
  assign n40523 = n36558 & ~n40522;
  assign n40524 = ~pi1156 & ~n36620;
  assign n40525 = ~n40511 & n40524;
  assign n40526 = pi219 & ~n40525;
  assign n40527 = ~n40521 & n40526;
  assign n40528 = ~n40523 & n40527;
  assign n40529 = ~n40517 & ~n40528;
  assign n40530 = ~pi263 & ~n40529;
  assign n40531 = ~pi299 & ~n40519;
  assign n40532 = ~n40508 & n40531;
  assign n40533 = ~n12342 & ~n36712;
  assign n40534 = ~n40531 & n40533;
  assign n40535 = pi1156 & ~n40534;
  assign n40536 = pi219 & ~n40532;
  assign n40537 = ~n40535 & n40536;
  assign n40538 = ~n36714 & ~n37481;
  assign n40539 = n36707 & n40538;
  assign n40540 = ~n37029 & ~n40539;
  assign n40541 = ~pi211 & ~n40540;
  assign n40542 = ~pi219 & ~n40541;
  assign n40543 = ~pi1156 & n40512;
  assign n40544 = ~n36610 & ~n36640;
  assign n40545 = pi1154 & ~n40544;
  assign n40546 = ~pi1154 & ~n36641;
  assign n40547 = ~n36745 & n40546;
  assign n40548 = pi1156 & ~n40545;
  assign n40549 = ~n40547 & n40548;
  assign n40550 = pi211 & ~n40543;
  assign n40551 = ~n40549 & n40550;
  assign n40552 = n40542 & ~n40551;
  assign n40553 = pi263 & pi1091;
  assign n40554 = ~n40537 & n40553;
  assign n40555 = ~n40552 & n40554;
  assign n40556 = ~n40530 & ~n40555;
  assign n40557 = ~po1038 & n40556;
  assign n40558 = pi219 & ~n36565;
  assign n40559 = ~pi219 & ~n36566;
  assign n40560 = ~n36579 & n40559;
  assign n40561 = ~n40558 & ~n40560;
  assign n40562 = pi1091 & ~n40561;
  assign n40563 = pi263 & ~pi1091;
  assign n40564 = ~n40562 & ~n40563;
  assign n40565 = po1038 & ~n40564;
  assign n40566 = ~n38687 & ~n40565;
  assign n40567 = ~n40557 & n40566;
  assign n40568 = pi1091 & n40558;
  assign n40569 = pi211 & n38718;
  assign n40570 = ~pi211 & ~n40510;
  assign n40571 = ~n36566 & ~n40570;
  assign n40572 = ~n40569 & n40571;
  assign n40573 = ~n38721 & ~n40572;
  assign n40574 = ~pi219 & ~n40573;
  assign n40575 = ~pi263 & ~n40327;
  assign n40576 = ~n40574 & n40575;
  assign n40577 = ~n36566 & ~n40269;
  assign n40578 = ~n40569 & ~n40577;
  assign n40579 = n40040 & ~n40578;
  assign n40580 = pi263 & ~n40043;
  assign n40581 = ~n40579 & n40580;
  assign n40582 = ~n40576 & ~n40581;
  assign n40583 = n38698 & ~n40568;
  assign n40584 = ~n40582 & n40583;
  assign n40585 = ~n38698 & n40564;
  assign n40586 = po1038 & ~n40585;
  assign n40587 = ~n40584 & n40586;
  assign n40588 = ~n38698 & ~n40556;
  assign n40589 = ~pi1155 & n40137;
  assign n40590 = pi1155 & ~n38780;
  assign n40591 = ~pi1154 & ~n40590;
  assign n40592 = ~n40589 & n40591;
  assign n40593 = pi1155 & n38779;
  assign n40594 = pi1154 & n38743;
  assign n40595 = ~n40593 & n40594;
  assign n40596 = ~n40592 & ~n40595;
  assign n40597 = ~pi1156 & ~n40596;
  assign n40598 = pi299 & n36558;
  assign n40599 = ~n38718 & n40598;
  assign n40600 = ~pi1154 & n38758;
  assign n40601 = ~n38807 & ~n40600;
  assign n40602 = pi1156 & ~n40593;
  assign n40603 = ~n40601 & n40602;
  assign n40604 = pi219 & ~n40599;
  assign n40605 = ~n40603 & n40604;
  assign n40606 = ~n40597 & n40605;
  assign n40607 = n38772 & n40591;
  assign n40608 = pi1155 & ~n38813;
  assign n40609 = ~pi1154 & ~n40608;
  assign n40610 = ~n40103 & n40609;
  assign n40611 = pi1156 & ~n40610;
  assign n40612 = pi1155 & ~n38854;
  assign n40613 = pi1154 & ~n40612;
  assign n40614 = n38829 & n40613;
  assign n40615 = ~n38738 & n40614;
  assign n40616 = ~n40607 & ~n40615;
  assign n40617 = n40611 & n40616;
  assign n40618 = ~n38750 & n40589;
  assign n40619 = n40609 & ~n40618;
  assign n40620 = ~pi1156 & ~n40619;
  assign n40621 = ~n40592 & ~n40614;
  assign n40622 = n40620 & n40621;
  assign n40623 = ~pi211 & ~n40617;
  assign n40624 = ~n40622 & n40623;
  assign n40625 = n40075 & n40613;
  assign n40626 = n40620 & ~n40625;
  assign n40627 = n38767 & n40613;
  assign n40628 = n40611 & ~n40627;
  assign n40629 = pi211 & ~n40626;
  assign n40630 = ~n40628 & n40629;
  assign n40631 = ~pi219 & ~n40624;
  assign n40632 = ~n40630 & n40631;
  assign n40633 = ~pi263 & ~n40606;
  assign n40634 = ~n40632 & n40633;
  assign n40635 = ~n38759 & ~n38796;
  assign n40636 = pi1154 & n38741;
  assign n40637 = ~n38784 & ~n40636;
  assign n40638 = ~pi1156 & n38732;
  assign n40639 = ~n40635 & ~n40638;
  assign n40640 = ~n40637 & n40639;
  assign n40641 = n36813 & n40041;
  assign n40642 = ~n40640 & ~n40641;
  assign n40643 = pi219 & ~n40642;
  assign n40644 = n38850 & ~n40346;
  assign n40645 = pi1154 & ~n38841;
  assign n40646 = ~n40644 & n40645;
  assign n40647 = ~n38732 & n38824;
  assign n40648 = n36561 & n40647;
  assign n40649 = n36566 & n38751;
  assign n40650 = ~pi1154 & ~n38860;
  assign n40651 = ~n40648 & n40650;
  assign n40652 = ~n40649 & n40651;
  assign n40653 = ~pi1156 & n40397;
  assign n40654 = ~n40652 & ~n40653;
  assign n40655 = pi1156 & n40134;
  assign n40656 = ~n40654 & ~n40655;
  assign n40657 = ~pi219 & ~n40646;
  assign n40658 = ~n40656 & n40657;
  assign n40659 = pi263 & ~n40643;
  assign n40660 = ~n40658 & n40659;
  assign n40661 = n38698 & ~n40660;
  assign n40662 = ~n40634 & n40661;
  assign n40663 = ~po1038 & ~n40588;
  assign n40664 = ~n40662 & n40663;
  assign n40665 = n38687 & ~n40587;
  assign n40666 = ~n40664 & n40665;
  assign n40667 = ~pi230 & ~n40567;
  assign n40668 = ~n40666 & n40667;
  assign n40669 = po1038 & n40561;
  assign n40670 = ~pi1154 & n10421;
  assign n40671 = ~n36621 & n36715;
  assign n40672 = ~pi1156 & ~n40671;
  assign n40673 = n36637 & ~n40670;
  assign n40674 = ~n40672 & n40673;
  assign n40675 = pi1156 & n12342;
  assign n40676 = pi219 & ~n40675;
  assign n40677 = ~n40674 & n40676;
  assign n40678 = ~n36545 & ~n40674;
  assign n40679 = pi211 & ~n40678;
  assign n40680 = n40542 & ~n40679;
  assign n40681 = ~po1038 & ~n40677;
  assign n40682 = ~n40680 & n40681;
  assign n40683 = pi230 & ~n40669;
  assign n40684 = ~n40682 & n40683;
  assign po420 = ~n40668 & ~n40684;
  assign n40686 = pi1091 & pi1143;
  assign n40687 = ~pi200 & n40686;
  assign n40688 = ~pi796 & n38702;
  assign n40689 = pi264 & ~n38702;
  assign n40690 = ~pi1091 & ~n40688;
  assign n40691 = ~n40689 & n40690;
  assign n40692 = pi199 & ~n40687;
  assign n40693 = ~n40691 & n40692;
  assign n40694 = pi1091 & pi1141;
  assign n40695 = ~pi796 & n38710;
  assign n40696 = pi264 & ~n38710;
  assign n40697 = ~pi1091 & ~n40695;
  assign n40698 = ~n40696 & n40697;
  assign n40699 = ~n40694 & ~n40698;
  assign n40700 = ~pi200 & ~n40699;
  assign n40701 = pi1091 & pi1142;
  assign n40702 = ~n40698 & ~n40701;
  assign n40703 = pi200 & ~n40702;
  assign n40704 = ~pi199 & ~n40700;
  assign n40705 = ~n40703 & n40704;
  assign n40706 = n15574 & ~n40693;
  assign n40707 = ~n40705 & n40706;
  assign n40708 = pi219 & ~n40268;
  assign n40709 = ~n37353 & ~n40708;
  assign n40710 = ~n40691 & ~n40709;
  assign n40711 = ~pi211 & ~n40699;
  assign n40712 = pi211 & ~n40702;
  assign n40713 = ~pi219 & ~n40711;
  assign n40714 = ~n40712 & n40713;
  assign n40715 = ~n15574 & ~n40710;
  assign n40716 = ~n40714 & n40715;
  assign n40717 = ~n40707 & ~n40716;
  assign n40718 = ~pi230 & ~n40717;
  assign n40719 = ~pi211 & pi1141;
  assign n40720 = ~pi219 & ~n36531;
  assign n40721 = ~n40719 & n40720;
  assign n40722 = ~n37353 & ~n40721;
  assign n40723 = ~n15574 & ~n40722;
  assign n40724 = ~pi199 & pi1141;
  assign n40725 = n37330 & ~n40724;
  assign n40726 = ~n36517 & ~n40725;
  assign n40727 = n15574 & ~n40726;
  assign n40728 = pi230 & ~n40723;
  assign n40729 = ~n40727 & n40728;
  assign po421 = n40718 | n40729;
  assign n40731 = pi1091 & pi1144;
  assign n40732 = ~pi200 & n40731;
  assign n40733 = ~pi819 & n38702;
  assign n40734 = pi265 & ~n38702;
  assign n40735 = ~pi1091 & ~n40733;
  assign n40736 = ~n40734 & n40735;
  assign n40737 = pi199 & ~n40732;
  assign n40738 = ~n40736 & n40737;
  assign n40739 = ~pi819 & n38710;
  assign n40740 = pi265 & ~n38710;
  assign n40741 = ~pi1091 & ~n40739;
  assign n40742 = ~n40740 & n40741;
  assign n40743 = ~n40701 & ~n40742;
  assign n40744 = ~pi200 & ~n40743;
  assign n40745 = ~n40686 & ~n40742;
  assign n40746 = pi200 & ~n40745;
  assign n40747 = ~pi199 & ~n40744;
  assign n40748 = ~n40746 & n40747;
  assign n40749 = n15574 & ~n40738;
  assign n40750 = ~n40748 & n40749;
  assign n40751 = ~n38552 & ~n40708;
  assign n40752 = ~n40736 & ~n40751;
  assign n40753 = ~pi211 & ~n40743;
  assign n40754 = pi211 & ~n40745;
  assign n40755 = ~pi219 & ~n40753;
  assign n40756 = ~n40754 & n40755;
  assign n40757 = ~n15574 & ~n40752;
  assign n40758 = ~n40756 & n40757;
  assign n40759 = ~n40750 & ~n40758;
  assign n40760 = ~pi230 & ~n40759;
  assign n40761 = ~pi219 & ~n36526;
  assign n40762 = ~n36537 & n40761;
  assign n40763 = ~n38552 & ~n40762;
  assign n40764 = ~n15574 & ~n40763;
  assign n40765 = ~n36516 & n38564;
  assign n40766 = ~n36510 & ~n40765;
  assign n40767 = n15574 & ~n40766;
  assign n40768 = pi230 & ~n40764;
  assign n40769 = ~n40767 & n40768;
  assign po422 = n40760 | n40769;
  assign n40771 = ~pi211 & pi1136;
  assign n40772 = pi219 & ~n40771;
  assign n40773 = pi211 & ~pi1135;
  assign n40774 = ~n40772 & ~n40773;
  assign n40775 = ~n10333 & n40774;
  assign n40776 = po1038 & n40775;
  assign n40777 = pi299 & n40775;
  assign n40778 = ~pi199 & pi1135;
  assign n40779 = pi200 & ~n40778;
  assign n40780 = pi199 & pi1136;
  assign n40781 = ~pi200 & ~n40780;
  assign n40782 = ~pi299 & ~n40779;
  assign n40783 = ~n40781 & n40782;
  assign n40784 = ~n40777 & ~n40783;
  assign n40785 = ~po1038 & ~n40784;
  assign n40786 = pi230 & ~n40776;
  assign n40787 = ~n40785 & n40786;
  assign n40788 = ~n40708 & ~n40772;
  assign n40789 = ~pi266 & ~n38702;
  assign n40790 = ~pi948 & n38702;
  assign n40791 = ~pi1091 & ~n40789;
  assign n40792 = ~n40790 & n40791;
  assign n40793 = ~n40788 & ~n40792;
  assign n40794 = ~n15574 & ~n40793;
  assign n40795 = ~pi266 & ~n38710;
  assign n40796 = ~pi948 & n38710;
  assign n40797 = ~pi1091 & ~n40795;
  assign n40798 = ~n40796 & n40797;
  assign n40799 = ~pi219 & ~n40798;
  assign n40800 = pi1135 & n40207;
  assign n40801 = n40799 & ~n40800;
  assign n40802 = n40794 & ~n40801;
  assign n40803 = ~pi199 & ~n40798;
  assign n40804 = pi1091 & pi1136;
  assign n40805 = pi199 & ~n40792;
  assign n40806 = ~n40804 & n40805;
  assign n40807 = ~n40803 & ~n40806;
  assign n40808 = ~pi200 & n40807;
  assign n40809 = pi1091 & pi1135;
  assign n40810 = n40803 & ~n40809;
  assign n40811 = pi200 & ~n40805;
  assign n40812 = ~n40810 & n40811;
  assign n40813 = ~n40808 & ~n40812;
  assign n40814 = n15574 & ~n40813;
  assign n40815 = ~pi230 & ~n40802;
  assign n40816 = ~n40814 & n40815;
  assign n40817 = ~n40787 & ~n40816;
  assign n40818 = ~pi1134 & ~n40817;
  assign n40819 = n36628 & ~n40780;
  assign n40820 = ~n40779 & ~n40819;
  assign n40821 = n15574 & n40820;
  assign n40822 = ~n15574 & n40774;
  assign n40823 = pi230 & ~n40821;
  assign n40824 = ~n40822 & n40823;
  assign n40825 = pi1091 & ~n40773;
  assign n40826 = n40799 & ~n40825;
  assign n40827 = n40794 & ~n40826;
  assign n40828 = ~pi199 & pi1091;
  assign n40829 = ~n40807 & ~n40828;
  assign n40830 = ~pi200 & ~n40829;
  assign n40831 = ~n40812 & ~n40830;
  assign n40832 = n15574 & ~n40831;
  assign n40833 = ~pi230 & ~n40827;
  assign n40834 = ~n40832 & n40833;
  assign n40835 = ~n40824 & ~n40834;
  assign n40836 = pi1134 & ~n40835;
  assign po423 = ~n40818 & ~n40836;
  assign n40838 = ~n36744 & ~n38623;
  assign n40839 = pi1153 & n12341;
  assign n40840 = n40510 & ~n40839;
  assign n40841 = ~n40838 & n40840;
  assign n40842 = n36598 & ~n37639;
  assign n40843 = pi1155 & n40842;
  assign n40844 = pi1154 & ~n40843;
  assign n40845 = pi1091 & n40844;
  assign n40846 = pi219 & pi299;
  assign n40847 = ~pi1155 & ~n36984;
  assign n40848 = ~n36625 & ~n40847;
  assign n40849 = ~n40846 & ~n40848;
  assign n40850 = n40845 & ~n40849;
  assign n40851 = pi211 & ~n40841;
  assign n40852 = ~n40850 & n40851;
  assign n40853 = ~n40002 & ~n40294;
  assign n40854 = ~n36744 & ~n40853;
  assign n40855 = n40510 & ~n40854;
  assign n40856 = pi1091 & n40501;
  assign n40857 = ~n40257 & n40856;
  assign n40858 = pi1154 & ~n40857;
  assign n40859 = ~pi299 & n36983;
  assign n40860 = pi1091 & ~n40859;
  assign n40861 = n40858 & n40860;
  assign n40862 = ~n40855 & ~n40861;
  assign n40863 = pi219 & ~n40862;
  assign n40864 = pi1091 & ~n37034;
  assign n40865 = ~n40838 & n40864;
  assign n40866 = ~pi1154 & n40865;
  assign n40867 = ~n11036 & ~n40258;
  assign n40868 = n40845 & n40867;
  assign n40869 = ~n40866 & ~n40868;
  assign n40870 = ~pi219 & ~n40869;
  assign n40871 = ~pi211 & ~n40863;
  assign n40872 = ~n40870 & n40871;
  assign n40873 = ~n40852 & ~n40872;
  assign n40874 = pi267 & ~n40873;
  assign n40875 = n38641 & ~n40865;
  assign n40876 = pi211 & ~pi1154;
  assign n40877 = ~n40875 & n40876;
  assign n40878 = n40268 & n40862;
  assign n40879 = n40501 & n40844;
  assign n40880 = pi1091 & ~pi1155;
  assign n40881 = n40859 & n40880;
  assign n40882 = n40858 & ~n40881;
  assign n40883 = pi211 & ~n40879;
  assign n40884 = ~n40882 & n40883;
  assign n40885 = ~n40878 & ~n40884;
  assign n40886 = pi219 & ~n40885;
  assign n40887 = ~n36984 & n40880;
  assign n40888 = n36562 & ~n40887;
  assign n40889 = ~n40857 & n40888;
  assign n40890 = ~n36738 & ~n36759;
  assign n40891 = ~n36975 & n40890;
  assign n40892 = pi1091 & n40891;
  assign n40893 = ~pi211 & ~n40892;
  assign n40894 = ~pi219 & ~n40889;
  assign n40895 = ~n40893 & n40894;
  assign n40896 = ~n40886 & ~n40895;
  assign n40897 = ~pi267 & ~n40877;
  assign n40898 = ~n40896 & n40897;
  assign n40899 = ~n40874 & ~n40898;
  assign n40900 = ~po1038 & n40899;
  assign n40901 = ~pi219 & ~n36562;
  assign n40902 = ~n36581 & n40901;
  assign n40903 = ~n37133 & ~n40902;
  assign n40904 = pi1091 & ~n40903;
  assign n40905 = ~pi267 & ~pi1091;
  assign n40906 = ~n40904 & ~n40905;
  assign n40907 = po1038 & ~n40906;
  assign n40908 = ~n38687 & ~n40907;
  assign n40909 = ~n40900 & n40908;
  assign n40910 = ~pi267 & ~n38722;
  assign n40911 = ~n40043 & n40910;
  assign n40912 = pi267 & n40329;
  assign n40913 = n38697 & ~n40911;
  assign n40914 = ~n40912 & n40913;
  assign n40915 = ~n38697 & n40905;
  assign n40916 = ~n40904 & ~n40915;
  assign n40917 = ~n40914 & n40916;
  assign n40918 = po1038 & ~n40917;
  assign n40919 = ~n38697 & ~n40899;
  assign n40920 = ~n40371 & n40378;
  assign n40921 = ~pi1154 & ~n38774;
  assign n40922 = ~n40920 & n40921;
  assign n40923 = pi1153 & n38783;
  assign n40924 = pi1154 & pi1155;
  assign n40925 = ~n38784 & n40924;
  assign n40926 = ~n40923 & n40925;
  assign n40927 = ~n40922 & ~n40926;
  assign n40928 = pi211 & ~n40927;
  assign n40929 = n36561 & ~n40060;
  assign n40930 = ~n40068 & n40929;
  assign n40931 = ~n40344 & n40930;
  assign n40932 = pi1154 & n38760;
  assign n40933 = ~pi1155 & ~n40920;
  assign n40934 = ~n40932 & n40933;
  assign n40935 = ~pi267 & ~n40931;
  assign n40936 = ~n40934 & n40935;
  assign n40937 = ~n40928 & n40936;
  assign n40938 = pi1155 & ~n40079;
  assign n40939 = n38779 & ~n40600;
  assign n40940 = n40938 & ~n40939;
  assign n40941 = ~n40083 & n40940;
  assign n40942 = ~pi1154 & ~n38743;
  assign n40943 = ~n40138 & n40942;
  assign n40944 = n38780 & ~n40364;
  assign n40945 = pi1154 & ~n40944;
  assign n40946 = ~pi1155 & ~n40943;
  assign n40947 = ~n40945 & n40946;
  assign n40948 = pi267 & ~n40941;
  assign n40949 = ~n40947 & n40948;
  assign n40950 = pi219 & ~n40949;
  assign n40951 = ~n40937 & n40950;
  assign n40952 = ~pi1153 & n38826;
  assign n40953 = ~n38854 & ~n40952;
  assign n40954 = pi1154 & n40953;
  assign n40955 = ~pi1153 & n38750;
  assign n40956 = ~pi1154 & ~n40955;
  assign n40957 = ~n38829 & n40956;
  assign n40958 = ~pi1155 & ~n40957;
  assign n40959 = ~n38824 & ~n40955;
  assign n40960 = ~n40958 & n40959;
  assign n40961 = ~pi211 & ~n40954;
  assign n40962 = ~n40960 & n40961;
  assign n40963 = ~pi1155 & n38813;
  assign n40964 = ~n40953 & n40963;
  assign n40965 = n40102 & n40938;
  assign n40966 = pi1154 & ~n40964;
  assign n40967 = ~n40965 & n40966;
  assign n40968 = ~n38767 & n40956;
  assign n40969 = ~n40958 & n40968;
  assign n40970 = pi211 & ~n40967;
  assign n40971 = ~n40969 & n40970;
  assign n40972 = pi267 & ~n40962;
  assign n40973 = ~n40971 & n40972;
  assign n40974 = pi1154 & n40647;
  assign n40975 = ~n40068 & ~n40134;
  assign n40976 = ~pi1155 & n38732;
  assign n40977 = ~n40975 & ~n40976;
  assign n40978 = ~n40974 & ~n40977;
  assign n40979 = ~pi211 & ~n40978;
  assign n40980 = n38752 & ~n40920;
  assign n40981 = ~pi1153 & ~n38854;
  assign n40982 = ~pi1154 & ~n40981;
  assign n40983 = pi1155 & ~n40982;
  assign n40984 = n38871 & ~n40983;
  assign n40985 = pi1155 & ~n40343;
  assign n40986 = n40975 & n40985;
  assign n40987 = pi1154 & ~n40986;
  assign n40988 = ~n40984 & ~n40987;
  assign n40989 = pi211 & ~n40980;
  assign n40990 = ~n40988 & n40989;
  assign n40991 = ~n40979 & ~n40990;
  assign n40992 = ~pi267 & ~n40991;
  assign n40993 = ~pi219 & ~n40973;
  assign n40994 = ~n40992 & n40993;
  assign n40995 = n38697 & ~n40951;
  assign n40996 = ~n40994 & n40995;
  assign n40997 = ~po1038 & ~n40919;
  assign n40998 = ~n40996 & n40997;
  assign n40999 = n38687 & ~n40918;
  assign n41000 = ~n40998 & n40999;
  assign n41001 = ~pi230 & ~n40909;
  assign n41002 = ~n41000 & n41001;
  assign n41003 = po1038 & n40903;
  assign n41004 = pi219 & ~n40842;
  assign n41005 = ~pi1155 & n40839;
  assign n41006 = ~pi1154 & ~n41005;
  assign n41007 = ~n36984 & ~n41006;
  assign n41008 = pi1155 & n36610;
  assign n41009 = ~n36969 & n41008;
  assign n41010 = ~n41007 & ~n41009;
  assign n41011 = ~n41004 & ~n41010;
  assign n41012 = pi211 & ~n41011;
  assign n41013 = ~pi199 & pi1154;
  assign n41014 = pi200 & ~n41013;
  assign n41015 = ~n36776 & ~n37639;
  assign n41016 = ~n41014 & n41015;
  assign n41017 = ~n36545 & ~n41016;
  assign n41018 = pi219 & ~n41017;
  assign n41019 = ~pi219 & n40891;
  assign n41020 = ~pi211 & ~n41019;
  assign n41021 = ~n41018 & n41020;
  assign n41022 = ~po1038 & ~n41021;
  assign n41023 = ~n41012 & n41022;
  assign n41024 = pi230 & ~n41003;
  assign n41025 = ~n41023 & n41024;
  assign po424 = ~n41002 & ~n41025;
  assign n41027 = ~po1038 & n36610;
  assign n41028 = ~n38086 & ~n41027;
  assign n41029 = ~pi199 & n15574;
  assign n41030 = ~n39426 & ~n41029;
  assign n41031 = pi1151 & ~n41030;
  assign n41032 = n41028 & ~n41031;
  assign n41033 = pi1150 & ~n41032;
  assign n41034 = pi1152 & n41033;
  assign n41035 = pi1091 & ~n41034;
  assign n41036 = pi268 & ~n41035;
  assign n41037 = ~pi1152 & n41030;
  assign n41038 = n41033 & ~n41037;
  assign n41039 = ~pi1151 & n40019;
  assign n41040 = ~po1038 & ~n11039;
  assign n41041 = po1038 & n11037;
  assign n41042 = ~n41040 & ~n41041;
  assign n41043 = pi1151 & ~n41042;
  assign n41044 = ~pi1152 & ~n41043;
  assign n41045 = ~n15574 & ~n40158;
  assign n41046 = ~po1038 & n36707;
  assign n41047 = ~n41045 & ~n41046;
  assign n41048 = pi1151 & n41047;
  assign n41049 = pi1152 & n41048;
  assign n41050 = ~pi1150 & ~n41039;
  assign n41051 = ~n41044 & n41050;
  assign n41052 = ~n41049 & n41051;
  assign n41053 = ~n41038 & ~n41052;
  assign n41054 = pi1091 & ~n41053;
  assign n41055 = ~n41036 & ~n41054;
  assign n41056 = ~n38686 & ~n41055;
  assign n41057 = po1038 & n40042;
  assign n41058 = ~po1038 & ~n40106;
  assign n41059 = ~n38727 & n41058;
  assign n41060 = ~n40040 & ~n41057;
  assign n41061 = ~n41059 & n41060;
  assign n41062 = ~pi1151 & n41061;
  assign n41063 = pi219 & ~n40062;
  assign n41064 = ~n38741 & n41063;
  assign n41065 = ~n40117 & ~n41064;
  assign n41066 = ~n38807 & ~n40139;
  assign n41067 = ~n41065 & ~n41066;
  assign n41068 = ~po1038 & ~n41067;
  assign n41069 = ~n40056 & ~n41057;
  assign n41070 = ~n41068 & n41069;
  assign n41071 = pi1151 & n41070;
  assign n41072 = ~pi268 & ~n41062;
  assign n41073 = ~n41071 & n41072;
  assign n41074 = n40096 & ~n40328;
  assign n41075 = pi219 & n38755;
  assign n41076 = n41058 & ~n41075;
  assign n41077 = ~n41074 & ~n41076;
  assign n41078 = n38718 & ~n41077;
  assign n41079 = ~pi1151 & n41078;
  assign n41080 = ~po1038 & ~n40122;
  assign n41081 = ~n40067 & n41080;
  assign n41082 = ~n40097 & ~n41081;
  assign n41083 = pi1151 & ~n41082;
  assign n41084 = pi268 & ~n41079;
  assign n41085 = ~n41083 & n41084;
  assign n41086 = ~pi1150 & ~n41085;
  assign n41087 = ~n41073 & n41086;
  assign n41088 = ~n38718 & ~n41077;
  assign n41089 = ~n41061 & ~n41088;
  assign n41090 = pi1151 & ~n41089;
  assign n41091 = po1038 & ~n40327;
  assign n41092 = ~n40048 & n41091;
  assign n41093 = n40044 & ~n40093;
  assign n41094 = ~n41092 & n41093;
  assign n41095 = pi219 & ~n38708;
  assign n41096 = ~n40067 & ~n41095;
  assign n41097 = ~n38734 & ~n41096;
  assign n41098 = ~po1038 & ~n38732;
  assign n41099 = n41097 & n41098;
  assign n41100 = ~n41094 & ~n41099;
  assign n41101 = ~pi1151 & ~n41100;
  assign n41102 = ~pi268 & ~n41090;
  assign n41103 = ~n41101 & n41102;
  assign n41104 = ~n40054 & n40096;
  assign n41105 = ~po1038 & ~n40082;
  assign n41106 = n41065 & n41105;
  assign n41107 = ~n41104 & ~n41106;
  assign n41108 = ~pi1151 & ~n41107;
  assign n41109 = pi1151 & ~n41077;
  assign n41110 = pi268 & ~n41109;
  assign n41111 = ~n41108 & n41110;
  assign n41112 = pi1150 & ~n41103;
  assign n41113 = ~n41111 & n41112;
  assign n41114 = ~pi1152 & ~n41087;
  assign n41115 = ~n41113 & n41114;
  assign n41116 = ~pi219 & n38840;
  assign n41117 = ~n41063 & ~n41116;
  assign n41118 = ~po1038 & ~n41117;
  assign n41119 = ~n40135 & n41118;
  assign n41120 = ~n40045 & ~n41119;
  assign n41121 = ~pi1151 & ~n41120;
  assign n41122 = n40044 & ~n40055;
  assign n41123 = ~po1038 & ~n41065;
  assign n41124 = ~n41122 & ~n41123;
  assign n41125 = pi1151 & ~n41124;
  assign n41126 = ~pi268 & ~n41121;
  assign n41127 = ~n41125 & n41126;
  assign n41128 = pi219 & ~n40083;
  assign n41129 = ~po1038 & ~n40139;
  assign n41130 = ~n41128 & n41129;
  assign n41131 = ~n41092 & ~n41130;
  assign n41132 = ~pi1151 & ~n41131;
  assign n41133 = ~n40094 & n41091;
  assign n41134 = ~n40067 & ~n41128;
  assign n41135 = n38832 & ~n41134;
  assign n41136 = ~po1038 & ~n41135;
  assign n41137 = ~n41133 & ~n41136;
  assign n41138 = pi1151 & ~n41137;
  assign n41139 = pi268 & ~n41132;
  assign n41140 = ~n41138 & n41139;
  assign n41141 = ~pi1150 & ~n41140;
  assign n41142 = ~n41127 & n41141;
  assign n41143 = ~n40054 & n41091;
  assign n41144 = ~n38707 & ~n40361;
  assign n41145 = n41068 & ~n41144;
  assign n41146 = ~n41143 & ~n41145;
  assign n41147 = ~pi1151 & ~n41146;
  assign n41148 = ~n38714 & n41105;
  assign n41149 = n41077 & ~n41092;
  assign n41150 = ~n41148 & n41149;
  assign n41151 = pi1151 & ~n41150;
  assign n41152 = pi268 & ~n41151;
  assign n41153 = ~n41147 & n41152;
  assign n41154 = ~n40061 & ~n41097;
  assign n41155 = ~po1038 & ~n41154;
  assign n41156 = ~n41093 & ~n41155;
  assign n41157 = ~pi1151 & ~n41156;
  assign n41158 = ~n41094 & ~n41122;
  assign n41159 = ~n41118 & n41158;
  assign n41160 = pi1151 & ~n41159;
  assign n41161 = ~pi268 & ~n41160;
  assign n41162 = ~n41157 & n41161;
  assign n41163 = pi1150 & ~n41162;
  assign n41164 = ~n41153 & n41163;
  assign n41165 = pi1152 & ~n41142;
  assign n41166 = ~n41164 & n41165;
  assign n41167 = n38686 & ~n41115;
  assign n41168 = ~n41166 & n41167;
  assign n41169 = ~n41056 & ~n41168;
  assign n41170 = ~pi230 & ~n41169;
  assign n41171 = pi230 & ~n41053;
  assign po425 = n41170 | n41171;
  assign n41173 = pi211 & pi1137;
  assign n41174 = ~n40771 & ~n41173;
  assign n41175 = pi1091 & ~n41174;
  assign n41176 = n39426 & ~n41175;
  assign n41177 = ~pi200 & n40804;
  assign n41178 = pi1137 & n38620;
  assign n41179 = ~n41177 & ~n41178;
  assign n41180 = n41029 & n41179;
  assign n41181 = ~n41176 & ~n41180;
  assign n41182 = ~pi817 & n38710;
  assign n41183 = pi269 & ~n38710;
  assign n41184 = ~pi1091 & ~n41182;
  assign n41185 = ~n41183 & n41184;
  assign n41186 = ~n41181 & ~n41185;
  assign n41187 = pi219 & ~n15574;
  assign n41188 = pi1138 & n40268;
  assign n41189 = n41187 & ~n41188;
  assign n41190 = ~pi200 & pi1091;
  assign n41191 = pi1138 & n41190;
  assign n41192 = pi199 & ~n41191;
  assign n41193 = n15574 & n41192;
  assign n41194 = ~n41189 & ~n41193;
  assign n41195 = ~pi817 & n38702;
  assign n41196 = pi269 & ~n38702;
  assign n41197 = ~pi1091 & ~n41195;
  assign n41198 = ~n41196 & n41197;
  assign n41199 = ~n41194 & ~n41198;
  assign n41200 = ~n41186 & ~n41199;
  assign n41201 = ~pi230 & ~n41200;
  assign n41202 = ~pi199 & pi1137;
  assign n41203 = pi200 & ~n41202;
  assign n41204 = pi199 & pi1138;
  assign n41205 = ~pi199 & pi1136;
  assign n41206 = ~pi200 & ~n41204;
  assign n41207 = ~n41205 & n41206;
  assign n41208 = ~n41203 & ~n41207;
  assign n41209 = n15574 & ~n41208;
  assign n41210 = ~pi219 & ~n41174;
  assign n41211 = ~pi211 & pi1138;
  assign n41212 = pi219 & n41211;
  assign n41213 = ~n41210 & ~n41212;
  assign n41214 = ~n15574 & n41213;
  assign n41215 = ~n41209 & ~n41214;
  assign n41216 = pi230 & ~n41215;
  assign po426 = ~n41201 & ~n41216;
  assign n41218 = pi1091 & n40719;
  assign n41219 = n41187 & ~n41218;
  assign n41220 = ~pi200 & n40694;
  assign n41221 = pi199 & ~n41220;
  assign n41222 = n15574 & n41221;
  assign n41223 = ~n41219 & ~n41222;
  assign n41224 = ~pi805 & n38702;
  assign n41225 = pi270 & ~n38702;
  assign n41226 = ~pi1091 & ~n41224;
  assign n41227 = ~n41225 & n41226;
  assign n41228 = ~n41223 & ~n41227;
  assign n41229 = ~pi211 & pi1139;
  assign n41230 = pi211 & pi1140;
  assign n41231 = ~n41229 & ~n41230;
  assign n41232 = pi1091 & ~n41231;
  assign n41233 = n39426 & ~n41232;
  assign n41234 = pi1140 & n38620;
  assign n41235 = pi1139 & n41190;
  assign n41236 = ~n41234 & ~n41235;
  assign n41237 = n41029 & n41236;
  assign n41238 = ~n41233 & ~n41237;
  assign n41239 = ~pi805 & n38710;
  assign n41240 = pi270 & ~n38710;
  assign n41241 = ~pi1091 & ~n41239;
  assign n41242 = ~n41240 & n41241;
  assign n41243 = ~n41238 & ~n41242;
  assign n41244 = ~pi230 & ~n41228;
  assign n41245 = ~n41243 & n41244;
  assign n41246 = ~pi219 & ~n41231;
  assign n41247 = pi219 & n40719;
  assign n41248 = ~n41246 & ~n41247;
  assign n41249 = ~n15574 & n41248;
  assign n41250 = ~pi199 & pi1140;
  assign n41251 = pi200 & ~n41250;
  assign n41252 = pi199 & pi1141;
  assign n41253 = ~pi199 & pi1139;
  assign n41254 = ~pi200 & ~n41252;
  assign n41255 = ~n41253 & n41254;
  assign n41256 = ~n41251 & ~n41255;
  assign n41257 = n15574 & ~n41256;
  assign n41258 = pi230 & ~n41249;
  assign n41259 = ~n41257 & n41258;
  assign po427 = n41245 | n41259;
  assign n41261 = ~pi271 & ~n38705;
  assign n41262 = ~n38715 & ~n41261;
  assign n41263 = pi199 & ~n41262;
  assign n41264 = pi1091 & pi1146;
  assign n41265 = ~n38713 & ~n41262;
  assign n41266 = ~n38720 & ~n41265;
  assign n41267 = ~n41264 & ~n41266;
  assign n41268 = ~pi199 & n41267;
  assign n41269 = ~n41263 & ~n41268;
  assign n41270 = pi200 & ~n41269;
  assign n41271 = pi1147 & n38634;
  assign n41272 = pi1091 & pi1145;
  assign n41273 = ~pi199 & ~n41272;
  assign n41274 = ~n41266 & n41273;
  assign n41275 = ~n41263 & ~n41274;
  assign n41276 = ~pi200 & ~n41271;
  assign n41277 = ~n41275 & n41276;
  assign n41278 = ~n41270 & ~n41277;
  assign n41279 = n15574 & ~n41278;
  assign n41280 = ~pi211 & pi1147;
  assign n41281 = n40038 & n41280;
  assign n41282 = pi219 & ~n41262;
  assign n41283 = ~pi211 & n41264;
  assign n41284 = ~n41267 & ~n41283;
  assign n41285 = pi1091 & n37354;
  assign n41286 = ~pi219 & ~n41285;
  assign n41287 = ~n41284 & n41286;
  assign n41288 = ~n41282 & ~n41287;
  assign n41289 = ~n15574 & ~n41281;
  assign n41290 = ~n41288 & n41289;
  assign n41291 = ~n41279 & ~n41290;
  assign n41292 = ~pi230 & ~n41291;
  assign n41293 = ~pi200 & ~n37335;
  assign n41294 = n37955 & ~n41293;
  assign n41295 = pi1147 & n40016;
  assign n41296 = ~n37978 & ~n37983;
  assign n41297 = ~pi219 & ~n41296;
  assign n41298 = ~n41294 & ~n41295;
  assign n41299 = ~n41297 & n41298;
  assign n41300 = ~po1038 & ~n41299;
  assign n41301 = pi219 & ~n41280;
  assign n41302 = ~n37354 & n39076;
  assign n41303 = ~n41301 & ~n41302;
  assign n41304 = po1038 & n41303;
  assign n41305 = pi230 & ~n41304;
  assign n41306 = ~n41300 & n41305;
  assign po428 = ~n41292 & ~n41306;
  assign n41308 = ~n12345 & ~n38014;
  assign n41309 = ~pi1149 & ~n41308;
  assign n41310 = ~pi1150 & ~n41309;
  assign n41311 = ~n41028 & ~n41310;
  assign n41312 = pi1149 & ~n41030;
  assign n41313 = ~n41311 & ~n41312;
  assign n41314 = pi1148 & ~n41313;
  assign n41315 = pi1150 & ~n40019;
  assign n41316 = ~pi1149 & ~n41315;
  assign n41317 = ~pi1150 & ~n41042;
  assign n41318 = pi1149 & ~pi1150;
  assign n41319 = pi1149 & n41047;
  assign n41320 = ~n41318 & ~n41319;
  assign n41321 = ~n41317 & ~n41320;
  assign n41322 = ~pi1148 & ~n41316;
  assign n41323 = ~n41321 & n41322;
  assign n41324 = ~n41314 & ~n41323;
  assign n41325 = pi1091 & ~n41324;
  assign n41326 = ~pi283 & ~n41325;
  assign n41327 = pi1150 & n41124;
  assign n41328 = ~pi1150 & ~n41070;
  assign n41329 = pi1149 & ~n41327;
  assign n41330 = ~n41328 & n41329;
  assign n41331 = pi1150 & n41120;
  assign n41332 = ~pi1150 & ~n41061;
  assign n41333 = ~pi1149 & ~n41332;
  assign n41334 = ~n41331 & n41333;
  assign n41335 = ~n41330 & ~n41334;
  assign n41336 = ~pi1148 & ~n41335;
  assign n41337 = ~pi1150 & ~n41089;
  assign n41338 = pi1150 & ~n41159;
  assign n41339 = pi1149 & ~n41337;
  assign n41340 = ~n41338 & n41339;
  assign n41341 = ~pi1150 & ~n41100;
  assign n41342 = pi1150 & ~n41156;
  assign n41343 = ~pi1149 & ~n41341;
  assign n41344 = ~n41342 & n41343;
  assign n41345 = pi1148 & ~n41340;
  assign n41346 = ~n41344 & n41345;
  assign n41347 = pi283 & ~n41346;
  assign n41348 = ~n41336 & n41347;
  assign n41349 = ~pi272 & ~n41326;
  assign n41350 = ~n41348 & n41349;
  assign n41351 = pi1091 & n41326;
  assign n41352 = pi1150 & ~n41146;
  assign n41353 = ~pi1150 & ~n41107;
  assign n41354 = ~pi1149 & ~n41353;
  assign n41355 = ~n41352 & n41354;
  assign n41356 = ~n41092 & ~n41148;
  assign n41357 = pi1150 & ~n41356;
  assign n41358 = pi1149 & n41077;
  assign n41359 = ~n41357 & n41358;
  assign n41360 = ~n41355 & ~n41359;
  assign n41361 = pi1148 & ~n41360;
  assign n41362 = pi1150 & n41137;
  assign n41363 = ~pi1150 & n41082;
  assign n41364 = pi1149 & ~n41363;
  assign n41365 = ~n41362 & n41364;
  assign n41366 = ~pi1150 & ~n41078;
  assign n41367 = pi1150 & n41131;
  assign n41368 = ~pi1149 & ~n41366;
  assign n41369 = ~n41367 & n41368;
  assign n41370 = ~pi1148 & ~n41369;
  assign n41371 = ~n41365 & n41370;
  assign n41372 = ~n41361 & ~n41371;
  assign n41373 = pi283 & ~n41372;
  assign n41374 = pi272 & ~n41351;
  assign n41375 = ~n41373 & n41374;
  assign n41376 = ~n41350 & ~n41375;
  assign n41377 = ~pi230 & ~n41376;
  assign n41378 = pi230 & ~n41324;
  assign po429 = n41377 | n41378;
  assign n41380 = ~pi273 & ~n38706;
  assign n41381 = ~n38717 & ~n41380;
  assign n41382 = pi219 & ~n41381;
  assign n41383 = ~n38720 & ~n41381;
  assign n41384 = ~n38721 & ~n41383;
  assign n41385 = ~pi219 & ~n41283;
  assign n41386 = ~n41384 & n41385;
  assign n41387 = ~n41382 & ~n41386;
  assign n41388 = po1038 & n41387;
  assign n41389 = ~n11038 & ~n38760;
  assign n41390 = pi1091 & ~n41389;
  assign n41391 = pi199 & ~n41381;
  assign n41392 = ~pi200 & n41264;
  assign n41393 = ~pi199 & ~n41392;
  assign n41394 = ~n41384 & n41393;
  assign n41395 = ~n41391 & ~n41394;
  assign n41396 = ~pi299 & ~n41395;
  assign n41397 = pi299 & ~n41387;
  assign n41398 = ~n41396 & ~n41397;
  assign n41399 = ~n41390 & ~n41398;
  assign n41400 = ~po1038 & ~n41399;
  assign n41401 = ~n40098 & ~n41400;
  assign n41402 = pi1147 & ~n41401;
  assign n41403 = n38061 & n41398;
  assign n41404 = ~pi1148 & ~n41403;
  assign n41405 = pi1091 & n40018;
  assign n41406 = n38635 & ~n41270;
  assign n41407 = n40268 & n40846;
  assign n41408 = ~n41406 & ~n41407;
  assign n41409 = ~n41398 & n41408;
  assign n41410 = ~po1038 & ~n41409;
  assign n41411 = pi1148 & ~n41405;
  assign n41412 = ~n41410 & n41411;
  assign n41413 = ~n41404 & ~n41412;
  assign n41414 = ~n41388 & ~n41413;
  assign n41415 = ~n41402 & n41414;
  assign n41416 = ~pi230 & ~n41415;
  assign n41417 = ~pi1148 & n41030;
  assign n41418 = ~pi1146 & n10333;
  assign n41419 = pi1147 & n39426;
  assign n41420 = ~n38086 & ~n41419;
  assign n41421 = ~n41418 & ~n41420;
  assign n41422 = ~pi199 & pi1147;
  assign n41423 = pi200 & ~n41422;
  assign n41424 = ~pi1146 & n10421;
  assign n41425 = ~n41423 & ~n41424;
  assign n41426 = n15574 & n41425;
  assign n41427 = ~n41421 & ~n41426;
  assign n41428 = pi230 & ~n41417;
  assign n41429 = ~n41427 & n41428;
  assign po430 = n41416 | n41429;
  assign n41431 = ~pi200 & n41272;
  assign n41432 = ~pi659 & n38702;
  assign n41433 = pi274 & ~n38702;
  assign n41434 = ~pi1091 & ~n41432;
  assign n41435 = ~n41433 & n41434;
  assign n41436 = pi199 & ~n41431;
  assign n41437 = ~n41435 & n41436;
  assign n41438 = ~pi659 & n38710;
  assign n41439 = pi274 & ~n38710;
  assign n41440 = ~pi1091 & ~n41438;
  assign n41441 = ~n41439 & n41440;
  assign n41442 = ~n40731 & ~n41441;
  assign n41443 = pi200 & ~n41442;
  assign n41444 = ~n40686 & ~n41441;
  assign n41445 = ~pi200 & ~n41444;
  assign n41446 = ~pi199 & ~n41443;
  assign n41447 = ~n41445 & n41446;
  assign n41448 = n15574 & ~n41437;
  assign n41449 = ~n41447 & n41448;
  assign n41450 = pi211 & ~n41442;
  assign n41451 = ~pi211 & ~n41444;
  assign n41452 = ~pi219 & ~n41450;
  assign n41453 = ~n41451 & n41452;
  assign n41454 = pi219 & ~n41285;
  assign n41455 = ~n41435 & n41454;
  assign n41456 = ~n15574 & ~n41455;
  assign n41457 = ~n41453 & n41456;
  assign n41458 = ~pi230 & ~n41449;
  assign n41459 = ~n41457 & n41458;
  assign n41460 = ~n36572 & ~n37978;
  assign n41461 = ~pi219 & ~n36530;
  assign n41462 = ~n37355 & n41461;
  assign n41463 = ~n41460 & ~n41462;
  assign n41464 = ~n36509 & n37960;
  assign n41465 = n38570 & ~n41464;
  assign n41466 = ~n41463 & ~n41465;
  assign n41467 = ~po1038 & ~n41466;
  assign n41468 = ~n37950 & ~n41462;
  assign n41469 = pi230 & ~n41467;
  assign n41470 = ~n41468 & n41469;
  assign po431 = ~n41459 & ~n41470;
  assign n41472 = pi1150 & ~n41070;
  assign n41473 = ~pi1151 & ~n41332;
  assign n41474 = ~n41472 & n41473;
  assign n41475 = ~pi1150 & n41120;
  assign n41476 = pi1151 & ~n41327;
  assign n41477 = ~n41475 & n41476;
  assign n41478 = ~pi275 & ~n41474;
  assign n41479 = ~n41477 & n41478;
  assign n41480 = pi1150 & n41082;
  assign n41481 = ~pi1151 & ~n41366;
  assign n41482 = ~n41480 & n41481;
  assign n41483 = ~pi1150 & n41131;
  assign n41484 = pi1151 & ~n41483;
  assign n41485 = ~n41362 & n41484;
  assign n41486 = pi275 & ~n41482;
  assign n41487 = ~n41485 & n41486;
  assign n41488 = ~pi1149 & ~n41487;
  assign n41489 = ~n41479 & n41488;
  assign n41490 = pi1151 & ~n41146;
  assign n41491 = ~pi1150 & ~n41108;
  assign n41492 = ~n41490 & n41491;
  assign n41493 = pi1150 & n41077;
  assign n41494 = ~n41151 & n41493;
  assign n41495 = ~n41492 & ~n41494;
  assign n41496 = pi275 & ~n41495;
  assign n41497 = pi1151 & ~n41156;
  assign n41498 = ~n41101 & ~n41497;
  assign n41499 = ~pi1150 & ~n41498;
  assign n41500 = ~pi1151 & ~n41089;
  assign n41501 = ~n41160 & ~n41500;
  assign n41502 = pi1150 & ~n41501;
  assign n41503 = ~pi275 & ~n41502;
  assign n41504 = ~n41499 & n41503;
  assign n41505 = pi1149 & ~n41504;
  assign n41506 = ~n41496 & n41505;
  assign n41507 = n38685 & ~n41489;
  assign n41508 = ~n41506 & n41507;
  assign n41509 = ~pi1151 & n41042;
  assign n41510 = ~pi1149 & n41509;
  assign n41511 = pi1149 & n41028;
  assign n41512 = pi1151 & ~n40019;
  assign n41513 = ~pi1149 & ~n41512;
  assign n41514 = ~pi1151 & n41308;
  assign n41515 = ~pi1150 & ~n41511;
  assign n41516 = ~n41513 & ~n41514;
  assign n41517 = n41515 & n41516;
  assign n41518 = ~pi1149 & n41048;
  assign n41519 = pi1151 & ~n41028;
  assign n41520 = pi1149 & n41030;
  assign n41521 = ~n41519 & n41520;
  assign n41522 = pi1150 & ~n41518;
  assign n41523 = ~n41521 & n41522;
  assign n41524 = ~n41517 & ~n41523;
  assign n41525 = ~n41510 & ~n41524;
  assign n41526 = pi1091 & ~n41525;
  assign n41527 = pi275 & ~n41526;
  assign n41528 = n41028 & n41318;
  assign n41529 = n38414 & ~n40019;
  assign n41530 = pi1150 & ~n41509;
  assign n41531 = ~n41048 & n41530;
  assign n41532 = ~pi1149 & ~n41529;
  assign n41533 = ~n41531 & n41532;
  assign n41534 = ~n41521 & ~n41528;
  assign n41535 = ~n41533 & n41534;
  assign n41536 = ~pi275 & pi1091;
  assign n41537 = n41535 & n41536;
  assign n41538 = ~n38685 & ~n41537;
  assign n41539 = ~n41527 & n41538;
  assign n41540 = ~n41508 & ~n41539;
  assign n41541 = ~pi230 & ~n41540;
  assign n41542 = pi230 & ~n41535;
  assign po432 = ~n41541 & ~n41542;
  assign n41544 = ~pi276 & ~n38703;
  assign n41545 = n38714 & ~n41544;
  assign n41546 = n41187 & ~n41283;
  assign n41547 = pi199 & ~n41392;
  assign n41548 = n15574 & n41547;
  assign n41549 = ~n41546 & ~n41548;
  assign n41550 = ~n41545 & ~n41549;
  assign n41551 = ~n36527 & ~n37939;
  assign n41552 = pi1091 & ~n41551;
  assign n41553 = n39426 & ~n41552;
  assign n41554 = pi1145 & n38620;
  assign n41555 = ~n40732 & ~n41554;
  assign n41556 = n41029 & n41555;
  assign n41557 = ~n41553 & ~n41556;
  assign n41558 = ~pi276 & ~n38711;
  assign n41559 = ~pi1091 & ~n38712;
  assign n41560 = ~n41558 & n41559;
  assign n41561 = ~n41557 & ~n41560;
  assign n41562 = ~pi230 & ~n41550;
  assign n41563 = ~n41561 & n41562;
  assign n41564 = ~n36507 & n39042;
  assign n41565 = ~n37962 & ~n41564;
  assign n41566 = n15574 & ~n41565;
  assign n41567 = pi219 & n37938;
  assign n41568 = ~pi219 & ~n41551;
  assign n41569 = ~n41567 & ~n41568;
  assign n41570 = ~n15574 & n41569;
  assign n41571 = pi230 & ~n41566;
  assign n41572 = ~n41570 & n41571;
  assign po433 = n41563 | n41572;
  assign n41574 = ~pi200 & n40701;
  assign n41575 = ~pi820 & n38702;
  assign n41576 = pi277 & ~n38702;
  assign n41577 = ~pi1091 & ~n41575;
  assign n41578 = ~n41576 & n41577;
  assign n41579 = pi199 & ~n41574;
  assign n41580 = ~n41578 & n41579;
  assign n41581 = pi1091 & pi1140;
  assign n41582 = ~pi820 & n38710;
  assign n41583 = pi277 & ~n38710;
  assign n41584 = ~pi1091 & ~n41582;
  assign n41585 = ~n41583 & n41584;
  assign n41586 = ~n41581 & ~n41585;
  assign n41587 = ~pi200 & ~n41586;
  assign n41588 = ~n40694 & ~n41585;
  assign n41589 = pi200 & ~n41588;
  assign n41590 = ~pi199 & ~n41587;
  assign n41591 = ~n41589 & n41590;
  assign n41592 = n15574 & ~n41580;
  assign n41593 = ~n41591 & n41592;
  assign n41594 = ~n36538 & ~n40708;
  assign n41595 = ~n41578 & ~n41594;
  assign n41596 = ~pi211 & ~n41586;
  assign n41597 = pi211 & ~n41588;
  assign n41598 = ~pi219 & ~n41596;
  assign n41599 = ~n41597 & n41598;
  assign n41600 = ~n15574 & ~n41595;
  assign n41601 = ~n41599 & n41600;
  assign n41602 = ~n41593 & ~n41601;
  assign n41603 = ~pi230 & ~n41602;
  assign n41604 = pi211 & pi1141;
  assign n41605 = ~pi211 & pi1140;
  assign n41606 = ~pi219 & ~n41604;
  assign n41607 = ~n41605 & n41606;
  assign n41608 = ~n36538 & ~n41607;
  assign n41609 = ~n15574 & ~n41608;
  assign n41610 = n36506 & ~n41250;
  assign n41611 = pi200 & ~n40724;
  assign n41612 = ~n41610 & ~n41611;
  assign n41613 = n15574 & ~n41612;
  assign n41614 = pi230 & ~n41609;
  assign n41615 = ~n41613 & n41614;
  assign po434 = n41603 | n41615;
  assign n41617 = ~pi278 & ~n38702;
  assign n41618 = ~pi976 & n38702;
  assign n41619 = ~pi1091 & ~n41617;
  assign n41620 = ~n41618 & n41619;
  assign n41621 = pi199 & ~n41620;
  assign n41622 = pi1091 & ~pi1132;
  assign n41623 = pi976 & n38710;
  assign n41624 = pi278 & ~n38710;
  assign n41625 = ~pi1091 & ~n41623;
  assign n41626 = ~n41624 & n41625;
  assign n41627 = ~n41622 & ~n41626;
  assign n41628 = ~pi199 & ~n41627;
  assign n41629 = ~n41621 & ~n41628;
  assign n41630 = ~pi200 & ~n41629;
  assign n41631 = pi1091 & ~pi1133;
  assign n41632 = ~n41626 & ~n41631;
  assign n41633 = ~pi199 & ~n41632;
  assign n41634 = ~n41621 & ~n41633;
  assign n41635 = pi200 & ~n41634;
  assign n41636 = ~pi299 & ~n41635;
  assign n41637 = ~n41630 & n41636;
  assign n41638 = pi219 & ~n41620;
  assign n41639 = ~pi211 & pi1132;
  assign n41640 = pi211 & pi1133;
  assign n41641 = ~n41639 & ~n41640;
  assign n41642 = pi1091 & n41641;
  assign n41643 = ~n41626 & ~n41642;
  assign n41644 = ~pi219 & ~n41643;
  assign n41645 = ~n41638 & ~n41644;
  assign n41646 = pi299 & n41645;
  assign n41647 = ~n41637 & ~n41646;
  assign n41648 = ~po1038 & ~n41647;
  assign n41649 = po1038 & n41645;
  assign n41650 = ~pi230 & ~n41649;
  assign n41651 = ~n41648 & n41650;
  assign n41652 = ~pi199 & pi1132;
  assign n41653 = ~pi200 & ~n41652;
  assign n41654 = ~pi199 & pi1133;
  assign n41655 = pi200 & ~n41654;
  assign n41656 = ~pi299 & ~n41655;
  assign n41657 = ~n41653 & n41656;
  assign n41658 = n36572 & ~n41641;
  assign n41659 = ~n41657 & ~n41658;
  assign n41660 = ~po1038 & ~n41659;
  assign n41661 = n37229 & ~n41641;
  assign n41662 = pi230 & ~n41661;
  assign n41663 = ~n41660 & n41662;
  assign n41664 = ~n41651 & ~n41663;
  assign n41665 = ~pi1134 & ~n41664;
  assign n41666 = n10421 & ~n41652;
  assign n41667 = n41656 & ~n41666;
  assign n41668 = ~n40222 & ~n41658;
  assign n41669 = ~n41667 & n41668;
  assign n41670 = ~po1038 & ~n41669;
  assign n41671 = ~n40018 & ~n41670;
  assign n41672 = n41662 & n41671;
  assign n41673 = ~n38634 & n41630;
  assign n41674 = n41636 & ~n41673;
  assign n41675 = ~n41407 & ~n41646;
  assign n41676 = ~n41674 & n41675;
  assign n41677 = ~po1038 & ~n41676;
  assign n41678 = ~n41405 & n41650;
  assign n41679 = ~n41677 & n41678;
  assign n41680 = ~n41672 & ~n41679;
  assign n41681 = pi1134 & ~n41680;
  assign po435 = ~n41665 & ~n41681;
  assign n41683 = ~pi279 & ~n38702;
  assign n41684 = ~pi958 & n38702;
  assign n41685 = ~pi1091 & ~n41683;
  assign n41686 = ~n41684 & n41685;
  assign n41687 = pi1135 & n41190;
  assign n41688 = ~n41686 & ~n41687;
  assign n41689 = pi199 & ~n41688;
  assign n41690 = pi958 & n38710;
  assign n41691 = pi279 & ~n38710;
  assign n41692 = ~pi1091 & ~n41690;
  assign n41693 = ~n41691 & n41692;
  assign n41694 = ~pi1133 & n41190;
  assign n41695 = ~pi199 & ~n41694;
  assign n41696 = ~n41693 & n41695;
  assign n41697 = ~n41689 & ~n41696;
  assign n41698 = n15574 & ~n41697;
  assign n41699 = ~n38620 & n41698;
  assign n41700 = ~n40207 & ~n41631;
  assign n41701 = ~n41693 & n41700;
  assign n41702 = ~pi219 & ~n41701;
  assign n41703 = pi1135 & n40268;
  assign n41704 = pi219 & ~n41703;
  assign n41705 = ~n41686 & n41704;
  assign n41706 = ~n15574 & ~n41705;
  assign n41707 = ~n41702 & n41706;
  assign n41708 = ~pi230 & ~n41707;
  assign n41709 = ~n41699 & n41708;
  assign n41710 = pi1135 & n36554;
  assign n41711 = ~pi211 & ~pi1133;
  assign n41712 = ~pi219 & ~n41711;
  assign n41713 = ~pi211 & n41712;
  assign n41714 = ~n41710 & ~n41713;
  assign n41715 = po1038 & ~n41714;
  assign n41716 = pi199 & pi1135;
  assign n41717 = ~n41654 & ~n41716;
  assign n41718 = n36610 & ~n41717;
  assign n41719 = pi299 & ~n41714;
  assign n41720 = ~n41718 & ~n41719;
  assign n41721 = ~po1038 & ~n41720;
  assign n41722 = pi230 & ~n41715;
  assign n41723 = ~n41721 & n41722;
  assign n41724 = ~n41709 & ~n41723;
  assign n41725 = ~pi1134 & ~n41724;
  assign n41726 = ~pi1133 & n10421;
  assign n41727 = ~pi200 & pi1135;
  assign n41728 = pi199 & ~n41727;
  assign n41729 = ~n41726 & ~n41728;
  assign n41730 = n15574 & ~n41729;
  assign n41731 = ~n41710 & ~n41712;
  assign n41732 = ~n15574 & n41731;
  assign n41733 = ~n41730 & ~n41732;
  assign n41734 = pi230 & ~n41733;
  assign n41735 = pi1091 & ~n41711;
  assign n41736 = n39426 & n41735;
  assign n41737 = ~n41698 & ~n41736;
  assign n41738 = n41708 & n41737;
  assign n41739 = ~n41734 & ~n41738;
  assign n41740 = pi1134 & ~n41739;
  assign po436 = ~n41725 & ~n41740;
  assign n41742 = pi1137 & n41190;
  assign n41743 = ~pi914 & n38702;
  assign n41744 = pi280 & ~n38702;
  assign n41745 = ~pi1091 & ~n41743;
  assign n41746 = ~n41744 & n41745;
  assign n41747 = ~n41742 & ~n41746;
  assign n41748 = pi199 & ~n41747;
  assign n41749 = ~pi280 & ~n38710;
  assign n41750 = pi914 & n38710;
  assign n41751 = ~pi1091 & ~n41749;
  assign n41752 = ~n41750 & n41751;
  assign n41753 = pi200 & pi1136;
  assign n41754 = pi1091 & ~n41727;
  assign n41755 = ~n41753 & n41754;
  assign n41756 = ~pi199 & ~n41755;
  assign n41757 = ~n41752 & n41756;
  assign n41758 = ~n41748 & ~n41757;
  assign n41759 = n15574 & ~n41758;
  assign n41760 = ~pi211 & pi1137;
  assign n41761 = pi219 & ~n41760;
  assign n41762 = ~n40708 & ~n41761;
  assign n41763 = ~n41746 & ~n41762;
  assign n41764 = ~pi211 & pi1135;
  assign n41765 = pi211 & pi1136;
  assign n41766 = ~n41764 & ~n41765;
  assign n41767 = pi1091 & n41766;
  assign n41768 = ~n41752 & ~n41767;
  assign n41769 = ~pi219 & ~n41768;
  assign n41770 = ~n15574 & ~n41763;
  assign n41771 = ~n41769 & n41770;
  assign n41772 = ~n41759 & ~n41771;
  assign n41773 = ~pi230 & ~n41772;
  assign n41774 = ~pi219 & n41766;
  assign n41775 = ~n41761 & ~n41774;
  assign n41776 = ~n15574 & ~n41775;
  assign n41777 = pi200 & ~n41205;
  assign n41778 = pi199 & pi1137;
  assign n41779 = ~pi200 & ~n40778;
  assign n41780 = ~n41778 & n41779;
  assign n41781 = ~n41777 & ~n41780;
  assign n41782 = n15574 & ~n41781;
  assign n41783 = pi230 & ~n41776;
  assign n41784 = ~n41782 & n41783;
  assign po437 = n41773 | n41784;
  assign n41786 = pi211 & pi1138;
  assign n41787 = ~n41760 & ~n41786;
  assign n41788 = pi1091 & ~n41787;
  assign n41789 = n39426 & ~n41788;
  assign n41790 = pi1138 & n38620;
  assign n41791 = ~n41742 & ~n41790;
  assign n41792 = n41029 & n41791;
  assign n41793 = ~n41789 & ~n41792;
  assign n41794 = ~pi830 & n38710;
  assign n41795 = pi281 & ~n38710;
  assign n41796 = ~pi1091 & ~n41794;
  assign n41797 = ~n41795 & n41796;
  assign n41798 = ~n41793 & ~n41797;
  assign n41799 = pi1139 & n40268;
  assign n41800 = n41187 & ~n41799;
  assign n41801 = pi199 & ~n41235;
  assign n41802 = n15574 & n41801;
  assign n41803 = ~n41800 & ~n41802;
  assign n41804 = ~pi830 & n38702;
  assign n41805 = pi281 & ~n38702;
  assign n41806 = ~pi1091 & ~n41804;
  assign n41807 = ~n41805 & n41806;
  assign n41808 = ~n41803 & ~n41807;
  assign n41809 = ~n41798 & ~n41808;
  assign n41810 = ~pi230 & ~n41809;
  assign n41811 = ~pi199 & pi1138;
  assign n41812 = pi200 & ~n41811;
  assign n41813 = pi199 & pi1139;
  assign n41814 = ~pi200 & ~n41202;
  assign n41815 = ~n41813 & n41814;
  assign n41816 = ~n41812 & ~n41815;
  assign n41817 = n15574 & ~n41816;
  assign n41818 = pi219 & n41229;
  assign n41819 = ~pi219 & ~n41787;
  assign n41820 = ~n41818 & ~n41819;
  assign n41821 = ~n15574 & n41820;
  assign n41822 = ~n41817 & ~n41821;
  assign n41823 = pi230 & ~n41822;
  assign po438 = ~n41810 & ~n41823;
  assign n41825 = pi211 & pi1139;
  assign n41826 = ~n41211 & ~n41825;
  assign n41827 = pi1091 & ~n41826;
  assign n41828 = n39426 & ~n41827;
  assign n41829 = pi1139 & n38620;
  assign n41830 = ~n41191 & ~n41829;
  assign n41831 = n41029 & n41830;
  assign n41832 = ~n41828 & ~n41831;
  assign n41833 = ~pi836 & n38710;
  assign n41834 = pi282 & ~n38710;
  assign n41835 = ~pi1091 & ~n41833;
  assign n41836 = ~n41834 & n41835;
  assign n41837 = ~n41832 & ~n41836;
  assign n41838 = pi1140 & n40268;
  assign n41839 = n41187 & ~n41838;
  assign n41840 = ~pi200 & n41581;
  assign n41841 = pi199 & ~n41840;
  assign n41842 = n15574 & n41841;
  assign n41843 = ~n41839 & ~n41842;
  assign n41844 = ~pi836 & n38702;
  assign n41845 = pi282 & ~n38702;
  assign n41846 = ~pi1091 & ~n41844;
  assign n41847 = ~n41845 & n41846;
  assign n41848 = ~n41843 & ~n41847;
  assign n41849 = ~n41837 & ~n41848;
  assign n41850 = ~pi230 & ~n41849;
  assign n41851 = pi200 & ~n41253;
  assign n41852 = pi199 & pi1140;
  assign n41853 = ~pi200 & ~n41811;
  assign n41854 = ~n41852 & n41853;
  assign n41855 = ~n41851 & ~n41854;
  assign n41856 = n15574 & ~n41855;
  assign n41857 = pi219 & n41605;
  assign n41858 = ~pi219 & ~n41826;
  assign n41859 = ~n41857 & ~n41858;
  assign n41860 = ~n15574 & n41859;
  assign n41861 = ~n41856 & ~n41860;
  assign n41862 = pi230 & ~n41861;
  assign po439 = ~n41850 & ~n41862;
  assign n41864 = ~pi1147 & n41120;
  assign n41865 = pi1147 & n41156;
  assign n41866 = pi1149 & ~n41864;
  assign n41867 = ~n41865 & n41866;
  assign n41868 = ~pi1147 & ~n41061;
  assign n41869 = pi1147 & n41100;
  assign n41870 = ~pi1149 & ~n41868;
  assign n41871 = ~n41869 & n41870;
  assign n41872 = ~n41867 & ~n41871;
  assign n41873 = ~pi1148 & ~n41872;
  assign n41874 = ~pi1147 & n41124;
  assign n41875 = pi1147 & n41159;
  assign n41876 = pi1149 & ~n41875;
  assign n41877 = ~n41874 & n41876;
  assign n41878 = ~pi1147 & ~n41070;
  assign n41879 = pi1147 & n41089;
  assign n41880 = ~pi1149 & ~n41879;
  assign n41881 = ~n41878 & n41880;
  assign n41882 = ~n41877 & ~n41881;
  assign n41883 = pi1148 & ~n41882;
  assign n41884 = ~pi283 & ~n41873;
  assign n41885 = ~n41883 & n41884;
  assign n41886 = ~pi1147 & ~n41082;
  assign n41887 = pi1147 & ~n41077;
  assign n41888 = pi1148 & ~n41887;
  assign n41889 = ~n41886 & n41888;
  assign n41890 = pi1147 & ~n41107;
  assign n41891 = ~pi1147 & n41078;
  assign n41892 = ~pi1148 & ~n41891;
  assign n41893 = ~n41890 & n41892;
  assign n41894 = ~pi1149 & ~n41889;
  assign n41895 = ~n41893 & n41894;
  assign n41896 = ~pi1147 & ~n41137;
  assign n41897 = pi1147 & ~n41150;
  assign n41898 = pi1148 & ~n41897;
  assign n41899 = ~n41896 & n41898;
  assign n41900 = pi1147 & ~n41146;
  assign n41901 = ~pi1147 & ~n41131;
  assign n41902 = ~pi1148 & ~n41901;
  assign n41903 = ~n41900 & n41902;
  assign n41904 = pi1149 & ~n41899;
  assign n41905 = ~n41903 & n41904;
  assign n41906 = pi283 & ~n41895;
  assign n41907 = ~n41905 & n41906;
  assign n41908 = ~n41885 & ~n41907;
  assign n41909 = ~pi230 & ~n41908;
  assign n41910 = pi1147 & ~n41308;
  assign n41911 = pi1149 & ~n40019;
  assign n41912 = ~n41910 & ~n41911;
  assign n41913 = ~pi1148 & ~n41912;
  assign n41914 = n41319 & ~n41910;
  assign n41915 = pi1147 & ~n41030;
  assign n41916 = ~pi1149 & n41042;
  assign n41917 = ~n41915 & n41916;
  assign n41918 = pi1148 & ~n41914;
  assign n41919 = ~n41917 & n41918;
  assign n41920 = pi230 & ~n41913;
  assign n41921 = ~n41919 & n41920;
  assign po440 = ~n41909 & ~n41921;
  assign n41923 = ~pi284 & n40469;
  assign n41924 = pi1143 & ~n40469;
  assign n41925 = ~n38089 & n41924;
  assign po441 = n41923 | n41925;
  assign n41927 = n2577 & ~n10031;
  assign po637 = ~po1038 & n41927;
  assign n41929 = ~n7351 & n41927;
  assign n41930 = pi286 & n41929;
  assign n41931 = pi288 & pi289;
  assign n41932 = n41930 & n41931;
  assign n41933 = ~pi285 & ~n41932;
  assign n41934 = pi285 & n41932;
  assign n41935 = po637 & ~n41933;
  assign n41936 = ~n41934 & n41935;
  assign n41937 = ~po1038 & n41932;
  assign n41938 = pi285 & ~pi289;
  assign n41939 = ~pi286 & n7351;
  assign n41940 = ~pi288 & n41939;
  assign n41941 = n41938 & n41940;
  assign n41942 = pi285 & ~n41941;
  assign n41943 = ~n41937 & n41942;
  assign n41944 = ~n41936 & ~n41943;
  assign po442 = ~pi793 & ~n41944;
  assign n41946 = ~pi288 & ~n7355;
  assign n41947 = n7351 & n41946;
  assign n41948 = pi286 & ~n41947;
  assign n41949 = ~pi286 & n41947;
  assign n41950 = po1038 & ~n41948;
  assign n41951 = ~n41949 & n41950;
  assign n41952 = n7351 & ~n41927;
  assign n41953 = pi286 & ~n41952;
  assign n41954 = ~n41927 & n41939;
  assign n41955 = ~n41953 & ~n41954;
  assign n41956 = n41946 & ~n41955;
  assign n41957 = ~pi286 & ~n41929;
  assign n41958 = pi288 & ~n41930;
  assign n41959 = ~n41957 & n41958;
  assign n41960 = ~po1038 & ~n41956;
  assign n41961 = ~n41959 & n41960;
  assign n41962 = ~pi793 & ~n41951;
  assign po443 = ~n41961 & n41962;
  assign n41964 = ~pi287 & pi457;
  assign po444 = ~pi332 & ~n41964;
  assign n41966 = pi288 & ~n7351;
  assign n41967 = ~n41947 & ~n41966;
  assign n41968 = po637 & ~n41967;
  assign n41969 = ~po637 & n41967;
  assign n41970 = ~pi793 & ~n41968;
  assign po445 = ~n41969 & n41970;
  assign n41972 = pi289 & ~n41940;
  assign n41973 = po1038 & ~n41941;
  assign n41974 = ~n41972 & n41973;
  assign n41975 = ~pi289 & n41958;
  assign n41976 = n41938 & n41954;
  assign n41977 = pi289 & ~n41954;
  assign n41978 = ~pi288 & ~n41976;
  assign n41979 = ~n41977 & n41978;
  assign n41980 = ~n41932 & ~n41975;
  assign n41981 = ~n41979 & n41980;
  assign n41982 = ~po1038 & ~n41981;
  assign n41983 = ~pi793 & ~n41974;
  assign po446 = ~n41982 & n41983;
  assign n41985 = ~pi476 & pi1048;
  assign n41986 = pi290 & pi476;
  assign po447 = n41985 | n41986;
  assign n41988 = ~pi476 & pi1049;
  assign n41989 = pi291 & pi476;
  assign po448 = n41988 | n41989;
  assign n41991 = ~pi476 & pi1084;
  assign n41992 = pi292 & pi476;
  assign po449 = n41991 | n41992;
  assign n41994 = ~pi476 & pi1059;
  assign n41995 = pi293 & pi476;
  assign po450 = n41994 | n41995;
  assign n41997 = ~pi476 & pi1072;
  assign n41998 = pi294 & pi476;
  assign po451 = n41997 | n41998;
  assign n42000 = ~pi476 & pi1053;
  assign n42001 = pi295 & pi476;
  assign po452 = n42000 | n42001;
  assign n42003 = ~pi476 & pi1037;
  assign n42004 = pi296 & pi476;
  assign po453 = n42003 | n42004;
  assign n42006 = ~pi476 & pi1044;
  assign n42007 = pi297 & pi476;
  assign po454 = n42006 | n42007;
  assign n42009 = ~pi298 & pi478;
  assign n42010 = ~pi478 & ~pi1044;
  assign po455 = ~n42009 & ~n42010;
  assign n42012 = pi54 & n2523;
  assign n42013 = ~pi54 & n12429;
  assign n42014 = n12670 & n42013;
  assign n42015 = ~n42012 & ~n42014;
  assign n42016 = n2575 & n8597;
  assign n42017 = ~n42015 & n42016;
  assign n42018 = ~pi39 & ~n42017;
  assign po456 = ~n10850 & ~n42018;
  assign n42020 = pi57 & ~pi59;
  assign n42021 = n9705 & n42020;
  assign n42022 = ~pi312 & n42021;
  assign n42023 = pi300 & ~n42022;
  assign n42024 = ~pi300 & n42022;
  assign n42025 = ~pi55 & ~n42024;
  assign po457 = n42023 | ~n42025;
  assign n42027 = ~pi301 & n42025;
  assign n42028 = ~pi300 & pi301;
  assign n42029 = ~pi55 & n42028;
  assign n42030 = n42022 & n42029;
  assign po458 = n42027 | n42030;
  assign n42032 = n5784 & ~po1038;
  assign n42033 = ~pi222 & ~pi223;
  assign n42034 = pi937 & ~n42033;
  assign n42035 = pi273 & n3328;
  assign n42036 = ~n42034 & ~n42035;
  assign n42037 = n42032 & n42036;
  assign n42038 = ~n2608 & n42037;
  assign n42039 = n3303 & ~n15574;
  assign n42040 = ~n42037 & ~n42039;
  assign n42041 = pi237 & ~n42040;
  assign n42042 = ~n5729 & ~n15574;
  assign n42043 = ~n42032 & ~n42042;
  assign n42044 = ~pi1148 & n42043;
  assign n42045 = ~pi215 & n3293;
  assign n42046 = ~pi273 & n42045;
  assign n42047 = ~pi937 & n5728;
  assign n42048 = ~n42046 & ~n42047;
  assign n42049 = ~n15574 & ~n42048;
  assign n42050 = ~n42038 & ~n42049;
  assign n42051 = ~n42041 & n42050;
  assign po459 = ~n42044 & n42051;
  assign n42053 = ~pi303 & pi478;
  assign n42054 = ~pi478 & ~pi1049;
  assign po460 = ~n42053 & ~n42054;
  assign n42056 = ~pi304 & pi478;
  assign n42057 = ~pi478 & ~pi1048;
  assign po461 = ~n42056 & ~n42057;
  assign n42059 = ~pi305 & pi478;
  assign n42060 = ~pi478 & ~pi1084;
  assign po462 = ~n42059 & ~n42060;
  assign n42062 = ~pi306 & pi478;
  assign n42063 = ~pi478 & ~pi1059;
  assign po463 = ~n42062 & ~n42063;
  assign n42065 = ~pi307 & pi478;
  assign n42066 = ~pi478 & ~pi1053;
  assign po464 = ~n42065 & ~n42066;
  assign n42068 = ~pi308 & pi478;
  assign n42069 = ~pi478 & ~pi1037;
  assign po465 = ~n42068 & ~n42069;
  assign n42071 = ~pi309 & pi478;
  assign n42072 = ~pi478 & ~pi1072;
  assign po466 = ~n42071 & ~n42072;
  assign n42074 = pi271 & n3293;
  assign n42075 = pi934 & ~n2461;
  assign n42076 = ~pi233 & n3303;
  assign n42077 = ~n42074 & ~n42075;
  assign n42078 = ~n42076 & n42077;
  assign n42079 = ~n5729 & n42078;
  assign n42080 = ~pi1147 & ~n3303;
  assign n42081 = n5729 & n42080;
  assign n42082 = ~n15574 & ~n42079;
  assign n42083 = ~n42081 & n42082;
  assign n42084 = pi233 & n2609;
  assign n42085 = pi222 & ~pi934;
  assign n42086 = ~pi271 & n3328;
  assign n42087 = ~n42085 & ~n42086;
  assign n42088 = n2598 & ~n42087;
  assign n42089 = ~pi1147 & ~n2598;
  assign n42090 = ~n42084 & ~n42088;
  assign n42091 = ~n42089 & n42090;
  assign n42092 = n15574 & n42091;
  assign po467 = n42083 | n42092;
  assign n42094 = pi311 & ~n42030;
  assign n42095 = ~pi55 & ~n42030;
  assign n42096 = ~pi311 & ~n42095;
  assign po468 = ~n42094 & ~n42096;
  assign n42098 = pi312 & ~n42021;
  assign n42099 = ~n42022 & ~n42098;
  assign po469 = ~pi55 & ~n42099;
  assign n42101 = ~n10010 & ~n12703;
  assign n42102 = po740 & ~n12710;
  assign n42103 = n9782 & ~n42102;
  assign po634 = n42101 | ~n42103;
  assign n42105 = ~pi954 & po634;
  assign n42106 = pi313 & pi954;
  assign po470 = ~n42105 & ~n42106;
  assign n42108 = n2572 & n12403;
  assign n42109 = n13616 & ~n42108;
  assign n42110 = ~pi39 & ~n13692;
  assign n42111 = pi39 & ~n14187;
  assign n42112 = n2613 & ~n42111;
  assign n42113 = ~n42110 & n42112;
  assign n42114 = ~n14480 & ~n42113;
  assign n42115 = n2535 & n12403;
  assign n42116 = ~n42114 & n42115;
  assign n42117 = ~n42109 & ~n42116;
  assign n42118 = n13608 & n13609;
  assign po471 = ~n42117 & n42118;
  assign n42120 = ~pi340 & n41927;
  assign n42121 = ~po1038 & n42120;
  assign n42122 = pi315 & ~n42121;
  assign n42123 = pi1080 & n42121;
  assign po472 = n42122 | n42123;
  assign n42125 = pi316 & ~n42121;
  assign n42126 = pi1047 & n42121;
  assign po473 = n42125 | n42126;
  assign n42128 = ~pi330 & po637;
  assign n42129 = pi317 & ~n42128;
  assign n42130 = pi1078 & n42128;
  assign po474 = n42129 | n42130;
  assign n42132 = ~pi341 & n41927;
  assign n42133 = ~po1038 & n42132;
  assign n42134 = pi318 & ~n42133;
  assign n42135 = pi1074 & n42133;
  assign po475 = n42134 | n42135;
  assign n42137 = pi319 & ~n42133;
  assign n42138 = pi1072 & n42133;
  assign po476 = n42137 | n42138;
  assign n42140 = pi320 & ~n42121;
  assign n42141 = pi1048 & n42121;
  assign po477 = n42140 | n42141;
  assign n42143 = pi321 & ~n42121;
  assign n42144 = pi1058 & n42121;
  assign po478 = n42143 | n42144;
  assign n42146 = pi322 & ~n42121;
  assign n42147 = pi1051 & n42121;
  assign po479 = n42146 | n42147;
  assign n42149 = pi323 & ~n42121;
  assign n42150 = pi1065 & n42121;
  assign po480 = n42149 | n42150;
  assign n42152 = pi324 & ~n42133;
  assign n42153 = pi1086 & n42133;
  assign po481 = n42152 | n42153;
  assign n42155 = pi325 & ~n42133;
  assign n42156 = pi1063 & n42133;
  assign po482 = n42155 | n42156;
  assign n42158 = pi326 & ~n42133;
  assign n42159 = pi1057 & n42133;
  assign po483 = n42158 | n42159;
  assign n42161 = pi327 & ~n42121;
  assign n42162 = pi1040 & n42121;
  assign po484 = n42161 | n42162;
  assign n42164 = pi328 & ~n42133;
  assign n42165 = pi1058 & n42133;
  assign po485 = n42164 | n42165;
  assign n42167 = pi329 & ~n42133;
  assign n42168 = pi1043 & n42133;
  assign po486 = n42167 | n42168;
  assign n42170 = pi1092 & ~n6178;
  assign n42171 = po1038 & n42170;
  assign n42172 = ~pi330 & n42171;
  assign n42173 = ~po1038 & n42170;
  assign n42174 = ~pi330 & ~n41927;
  assign n42175 = ~n42120 & ~n42174;
  assign n42176 = n42173 & ~n42175;
  assign po487 = n42172 | n42176;
  assign n42178 = ~pi331 & n42171;
  assign n42179 = ~pi331 & ~n41927;
  assign n42180 = ~n42132 & ~n42179;
  assign n42181 = n42173 & ~n42180;
  assign po488 = n42178 | n42181;
  assign n42183 = n10603 & n12445;
  assign n42184 = ~n10603 & ~n12379;
  assign n42185 = n7376 & ~n42184;
  assign n42186 = ~pi70 & ~n42185;
  assign n42187 = pi332 & n8798;
  assign n42188 = ~n42186 & n42187;
  assign n42189 = ~n42183 & ~n42188;
  assign n42190 = ~pi39 & ~n42189;
  assign n42191 = pi39 & n10001;
  assign n42192 = ~pi38 & ~n42191;
  assign n42193 = ~n42190 & n42192;
  assign po489 = n36367 & ~n42193;
  assign n42195 = pi333 & ~n42133;
  assign n42196 = pi1040 & n42133;
  assign po490 = n42195 | n42196;
  assign n42198 = pi334 & ~n42133;
  assign n42199 = pi1065 & n42133;
  assign po491 = n42198 | n42199;
  assign n42201 = pi335 & ~n42133;
  assign n42202 = pi1069 & n42133;
  assign po492 = n42201 | n42202;
  assign n42204 = pi336 & ~n42128;
  assign n42205 = pi1070 & n42128;
  assign po493 = n42204 | n42205;
  assign n42207 = pi337 & ~n42128;
  assign n42208 = pi1044 & n42128;
  assign po494 = n42207 | n42208;
  assign n42210 = pi338 & ~n42128;
  assign n42211 = pi1072 & n42128;
  assign po495 = n42210 | n42211;
  assign n42213 = pi339 & ~n42128;
  assign n42214 = pi1086 & n42128;
  assign po496 = n42213 | n42214;
  assign n42216 = pi340 & n42171;
  assign n42217 = ~pi340 & ~n41927;
  assign n42218 = ~pi331 & n41927;
  assign n42219 = n42173 & ~n42217;
  assign n42220 = ~n42218 & n42219;
  assign po497 = ~n42216 & ~n42220;
  assign n42222 = ~pi341 & ~po637;
  assign n42223 = ~n42128 & ~n42222;
  assign po498 = n42170 & ~n42223;
  assign n42225 = pi342 & ~n42121;
  assign n42226 = pi1049 & n42121;
  assign po499 = n42225 | n42226;
  assign n42228 = pi343 & ~n42121;
  assign n42229 = pi1062 & n42121;
  assign po500 = n42228 | n42229;
  assign n42231 = pi344 & ~n42121;
  assign n42232 = pi1069 & n42121;
  assign po501 = n42231 | n42232;
  assign n42234 = pi345 & ~n42121;
  assign n42235 = pi1039 & n42121;
  assign po502 = n42234 | n42235;
  assign n42237 = pi346 & ~n42121;
  assign n42238 = pi1067 & n42121;
  assign po503 = n42237 | n42238;
  assign n42240 = pi347 & ~n42121;
  assign n42241 = pi1055 & n42121;
  assign po504 = n42240 | n42241;
  assign n42243 = pi348 & ~n42121;
  assign n42244 = pi1087 & n42121;
  assign po505 = n42243 | n42244;
  assign n42246 = pi349 & ~n42121;
  assign n42247 = pi1043 & n42121;
  assign po506 = n42246 | n42247;
  assign n42249 = pi350 & ~n42121;
  assign n42250 = pi1035 & n42121;
  assign po507 = n42249 | n42250;
  assign n42252 = pi351 & ~n42121;
  assign n42253 = pi1079 & n42121;
  assign po508 = n42252 | n42253;
  assign n42255 = pi352 & ~n42121;
  assign n42256 = pi1078 & n42121;
  assign po509 = n42255 | n42256;
  assign n42258 = pi353 & ~n42121;
  assign n42259 = pi1063 & n42121;
  assign po510 = n42258 | n42259;
  assign n42261 = pi354 & ~n42121;
  assign n42262 = pi1045 & n42121;
  assign po511 = n42261 | n42262;
  assign n42264 = pi355 & ~n42121;
  assign n42265 = pi1084 & n42121;
  assign po512 = n42264 | n42265;
  assign n42267 = pi356 & ~n42121;
  assign n42268 = pi1081 & n42121;
  assign po513 = n42267 | n42268;
  assign n42270 = pi357 & ~n42121;
  assign n42271 = pi1076 & n42121;
  assign po514 = n42270 | n42271;
  assign n42273 = pi358 & ~n42121;
  assign n42274 = pi1071 & n42121;
  assign po515 = n42273 | n42274;
  assign n42276 = pi359 & ~n42121;
  assign n42277 = pi1068 & n42121;
  assign po516 = n42276 | n42277;
  assign n42279 = pi360 & ~n42121;
  assign n42280 = pi1042 & n42121;
  assign po517 = n42279 | n42280;
  assign n42282 = pi361 & ~n42121;
  assign n42283 = pi1059 & n42121;
  assign po518 = n42282 | n42283;
  assign n42285 = pi362 & ~n42121;
  assign n42286 = pi1070 & n42121;
  assign po519 = n42285 | n42286;
  assign n42288 = pi363 & ~n42128;
  assign n42289 = pi1049 & n42128;
  assign po520 = n42288 | n42289;
  assign n42291 = pi364 & ~n42128;
  assign n42292 = pi1062 & n42128;
  assign po521 = n42291 | n42292;
  assign n42294 = pi365 & ~n42128;
  assign n42295 = pi1065 & n42128;
  assign po522 = n42294 | n42295;
  assign n42297 = pi366 & ~n42128;
  assign n42298 = pi1069 & n42128;
  assign po523 = n42297 | n42298;
  assign n42300 = pi367 & ~n42128;
  assign n42301 = pi1039 & n42128;
  assign po524 = n42300 | n42301;
  assign n42303 = pi368 & ~n42128;
  assign n42304 = pi1067 & n42128;
  assign po525 = n42303 | n42304;
  assign n42306 = pi369 & ~n42128;
  assign n42307 = pi1080 & n42128;
  assign po526 = n42306 | n42307;
  assign n42309 = pi370 & ~n42128;
  assign n42310 = pi1055 & n42128;
  assign po527 = n42309 | n42310;
  assign n42312 = pi371 & ~n42128;
  assign n42313 = pi1051 & n42128;
  assign po528 = n42312 | n42313;
  assign n42315 = pi372 & ~n42128;
  assign n42316 = pi1048 & n42128;
  assign po529 = n42315 | n42316;
  assign n42318 = pi373 & ~n42128;
  assign n42319 = pi1087 & n42128;
  assign po530 = n42318 | n42319;
  assign n42321 = pi374 & ~n42128;
  assign n42322 = pi1035 & n42128;
  assign po531 = n42321 | n42322;
  assign n42324 = pi375 & ~n42128;
  assign n42325 = pi1047 & n42128;
  assign po532 = n42324 | n42325;
  assign n42327 = pi376 & ~n42128;
  assign n42328 = pi1079 & n42128;
  assign po533 = n42327 | n42328;
  assign n42330 = pi377 & ~n42128;
  assign n42331 = pi1074 & n42128;
  assign po534 = n42330 | n42331;
  assign n42333 = pi378 & ~n42128;
  assign n42334 = pi1063 & n42128;
  assign po535 = n42333 | n42334;
  assign n42336 = pi379 & ~n42128;
  assign n42337 = pi1045 & n42128;
  assign po536 = n42336 | n42337;
  assign n42339 = pi380 & ~n42128;
  assign n42340 = pi1084 & n42128;
  assign po537 = n42339 | n42340;
  assign n42342 = pi381 & ~n42128;
  assign n42343 = pi1081 & n42128;
  assign po538 = n42342 | n42343;
  assign n42345 = pi382 & ~n42128;
  assign n42346 = pi1076 & n42128;
  assign po539 = n42345 | n42346;
  assign n42348 = pi383 & ~n42128;
  assign n42349 = pi1071 & n42128;
  assign po540 = n42348 | n42349;
  assign n42351 = pi384 & ~n42128;
  assign n42352 = pi1068 & n42128;
  assign po541 = n42351 | n42352;
  assign n42354 = pi385 & ~n42128;
  assign n42355 = pi1042 & n42128;
  assign po542 = n42354 | n42355;
  assign n42357 = pi386 & ~n42128;
  assign n42358 = pi1059 & n42128;
  assign po543 = n42357 | n42358;
  assign n42360 = pi387 & ~n42128;
  assign n42361 = pi1053 & n42128;
  assign po544 = n42360 | n42361;
  assign n42363 = pi388 & ~n42128;
  assign n42364 = pi1037 & n42128;
  assign po545 = n42363 | n42364;
  assign n42366 = pi389 & ~n42128;
  assign n42367 = pi1036 & n42128;
  assign po546 = n42366 | n42367;
  assign n42369 = pi390 & ~n42133;
  assign n42370 = pi1049 & n42133;
  assign po547 = n42369 | n42370;
  assign n42372 = pi391 & ~n42133;
  assign n42373 = pi1062 & n42133;
  assign po548 = n42372 | n42373;
  assign n42375 = pi392 & ~n42133;
  assign n42376 = pi1039 & n42133;
  assign po549 = n42375 | n42376;
  assign n42378 = pi393 & ~n42133;
  assign n42379 = pi1067 & n42133;
  assign po550 = n42378 | n42379;
  assign n42381 = pi394 & ~n42133;
  assign n42382 = pi1080 & n42133;
  assign po551 = n42381 | n42382;
  assign n42384 = pi395 & ~n42133;
  assign n42385 = pi1055 & n42133;
  assign po552 = n42384 | n42385;
  assign n42387 = pi396 & ~n42133;
  assign n42388 = pi1051 & n42133;
  assign po553 = n42387 | n42388;
  assign n42390 = pi397 & ~n42133;
  assign n42391 = pi1048 & n42133;
  assign po554 = n42390 | n42391;
  assign n42393 = pi398 & ~n42133;
  assign n42394 = pi1087 & n42133;
  assign po555 = n42393 | n42394;
  assign n42396 = pi399 & ~n42133;
  assign n42397 = pi1047 & n42133;
  assign po556 = n42396 | n42397;
  assign n42399 = pi400 & ~n42133;
  assign n42400 = pi1035 & n42133;
  assign po557 = n42399 | n42400;
  assign n42402 = pi401 & ~n42133;
  assign n42403 = pi1079 & n42133;
  assign po558 = n42402 | n42403;
  assign n42405 = pi402 & ~n42133;
  assign n42406 = pi1078 & n42133;
  assign po559 = n42405 | n42406;
  assign n42408 = pi403 & ~n42133;
  assign n42409 = pi1045 & n42133;
  assign po560 = n42408 | n42409;
  assign n42411 = pi404 & ~n42133;
  assign n42412 = pi1084 & n42133;
  assign po561 = n42411 | n42412;
  assign n42414 = pi405 & ~n42133;
  assign n42415 = pi1081 & n42133;
  assign po562 = n42414 | n42415;
  assign n42417 = pi406 & ~n42133;
  assign n42418 = pi1076 & n42133;
  assign po563 = n42417 | n42418;
  assign n42420 = pi407 & ~n42133;
  assign n42421 = pi1071 & n42133;
  assign po564 = n42420 | n42421;
  assign n42423 = pi408 & ~n42133;
  assign n42424 = pi1068 & n42133;
  assign po565 = n42423 | n42424;
  assign n42426 = pi409 & ~n42133;
  assign n42427 = pi1042 & n42133;
  assign po566 = n42426 | n42427;
  assign n42429 = pi410 & ~n42133;
  assign n42430 = pi1059 & n42133;
  assign po567 = n42429 | n42430;
  assign n42432 = pi411 & ~n42133;
  assign n42433 = pi1053 & n42133;
  assign po568 = n42432 | n42433;
  assign n42435 = pi412 & ~n42133;
  assign n42436 = pi1037 & n42133;
  assign po569 = n42435 | n42436;
  assign n42438 = pi413 & ~n42133;
  assign n42439 = pi1036 & n42133;
  assign po570 = n42438 | n42439;
  assign n42441 = ~po1038 & n42218;
  assign n42442 = pi414 & ~n42441;
  assign n42443 = pi1049 & n42441;
  assign po571 = n42442 | n42443;
  assign n42445 = pi415 & ~n42441;
  assign n42446 = pi1062 & n42441;
  assign po572 = n42445 | n42446;
  assign n42448 = pi416 & ~n42441;
  assign n42449 = pi1069 & n42441;
  assign po573 = n42448 | n42449;
  assign n42451 = pi417 & ~n42441;
  assign n42452 = pi1039 & n42441;
  assign po574 = n42451 | n42452;
  assign n42454 = pi418 & ~n42441;
  assign n42455 = pi1067 & n42441;
  assign po575 = n42454 | n42455;
  assign n42457 = pi419 & ~n42441;
  assign n42458 = pi1080 & n42441;
  assign po576 = n42457 | n42458;
  assign n42460 = pi420 & ~n42441;
  assign n42461 = pi1055 & n42441;
  assign po577 = n42460 | n42461;
  assign n42463 = pi421 & ~n42441;
  assign n42464 = pi1051 & n42441;
  assign po578 = n42463 | n42464;
  assign n42466 = pi422 & ~n42441;
  assign n42467 = pi1048 & n42441;
  assign po579 = n42466 | n42467;
  assign n42469 = pi423 & ~n42441;
  assign n42470 = pi1087 & n42441;
  assign po580 = n42469 | n42470;
  assign n42472 = pi424 & ~n42441;
  assign n42473 = pi1047 & n42441;
  assign po581 = n42472 | n42473;
  assign n42475 = pi425 & ~n42441;
  assign n42476 = pi1035 & n42441;
  assign po582 = n42475 | n42476;
  assign n42478 = pi426 & ~n42441;
  assign n42479 = pi1079 & n42441;
  assign po583 = n42478 | n42479;
  assign n42481 = pi427 & ~n42441;
  assign n42482 = pi1078 & n42441;
  assign po584 = n42481 | n42482;
  assign n42484 = pi428 & ~n42441;
  assign n42485 = pi1045 & n42441;
  assign po585 = n42484 | n42485;
  assign n42487 = pi429 & ~n42441;
  assign n42488 = pi1084 & n42441;
  assign po586 = n42487 | n42488;
  assign n42490 = pi430 & ~n42441;
  assign n42491 = pi1076 & n42441;
  assign po587 = n42490 | n42491;
  assign n42493 = pi431 & ~n42441;
  assign n42494 = pi1071 & n42441;
  assign po588 = n42493 | n42494;
  assign n42496 = pi432 & ~n42441;
  assign n42497 = pi1068 & n42441;
  assign po589 = n42496 | n42497;
  assign n42499 = pi433 & ~n42441;
  assign n42500 = pi1042 & n42441;
  assign po590 = n42499 | n42500;
  assign n42502 = pi434 & ~n42441;
  assign n42503 = pi1059 & n42441;
  assign po591 = n42502 | n42503;
  assign n42505 = pi435 & ~n42441;
  assign n42506 = pi1053 & n42441;
  assign po592 = n42505 | n42506;
  assign n42508 = pi436 & ~n42441;
  assign n42509 = pi1037 & n42441;
  assign po593 = n42508 | n42509;
  assign n42511 = pi437 & ~n42441;
  assign n42512 = pi1070 & n42441;
  assign po594 = n42511 | n42512;
  assign n42514 = pi438 & ~n42441;
  assign n42515 = pi1036 & n42441;
  assign po595 = n42514 | n42515;
  assign n42517 = pi439 & ~n42128;
  assign n42518 = pi1057 & n42128;
  assign po596 = n42517 | n42518;
  assign n42520 = pi440 & ~n42128;
  assign n42521 = pi1043 & n42128;
  assign po597 = n42520 | n42521;
  assign n42523 = pi441 & ~n42121;
  assign n42524 = pi1044 & n42121;
  assign po598 = n42523 | n42524;
  assign n42526 = pi442 & ~n42128;
  assign n42527 = pi1058 & n42128;
  assign po599 = n42526 | n42527;
  assign n42529 = pi443 & ~n42441;
  assign n42530 = pi1044 & n42441;
  assign po600 = n42529 | n42530;
  assign n42532 = pi444 & ~n42441;
  assign n42533 = pi1072 & n42441;
  assign po601 = n42532 | n42533;
  assign n42535 = pi445 & ~n42441;
  assign n42536 = pi1081 & n42441;
  assign po602 = n42535 | n42536;
  assign n42538 = pi446 & ~n42441;
  assign n42539 = pi1086 & n42441;
  assign po603 = n42538 | n42539;
  assign n42541 = pi447 & ~n42128;
  assign n42542 = pi1040 & n42128;
  assign po604 = n42541 | n42542;
  assign n42544 = pi448 & ~n42441;
  assign n42545 = pi1074 & n42441;
  assign po605 = n42544 | n42545;
  assign n42547 = pi449 & ~n42441;
  assign n42548 = pi1057 & n42441;
  assign po606 = n42547 | n42548;
  assign n42550 = pi450 & ~n42121;
  assign n42551 = pi1036 & n42121;
  assign po607 = n42550 | n42551;
  assign n42553 = pi451 & ~n42441;
  assign n42554 = pi1063 & n42441;
  assign po608 = n42553 | n42554;
  assign n42556 = pi452 & ~n42121;
  assign n42557 = pi1053 & n42121;
  assign po609 = n42556 | n42557;
  assign n42559 = pi453 & ~n42441;
  assign n42560 = pi1040 & n42441;
  assign po610 = n42559 | n42560;
  assign n42562 = pi454 & ~n42441;
  assign n42563 = pi1043 & n42441;
  assign po611 = n42562 | n42563;
  assign n42565 = pi455 & ~n42121;
  assign n42566 = pi1037 & n42121;
  assign po612 = n42565 | n42566;
  assign n42568 = pi456 & ~n42133;
  assign n42569 = pi1044 & n42133;
  assign po613 = n42568 | n42569;
  assign n42571 = ~pi804 & ~pi810;
  assign n42572 = ~pi595 & ~n42571;
  assign n42573 = ~pi599 & pi810;
  assign n42574 = pi596 & ~n42573;
  assign n42575 = pi804 & ~n42574;
  assign n42576 = pi815 & ~n42575;
  assign n42577 = pi595 & ~n42576;
  assign n42578 = pi594 & pi600;
  assign n42579 = pi597 & n42578;
  assign n42580 = pi601 & n42579;
  assign n42581 = ~n42572 & n42580;
  assign n42582 = ~n42577 & n42581;
  assign n42583 = pi600 & ~pi810;
  assign n42584 = pi804 & ~n42583;
  assign n42585 = ~pi601 & ~n42571;
  assign n42586 = ~pi815 & ~n42584;
  assign n42587 = ~n42585 & n42586;
  assign n42588 = ~n42582 & ~n42587;
  assign n42589 = pi605 & ~n42588;
  assign n42590 = pi990 & n42578;
  assign n42591 = ~pi815 & n42584;
  assign n42592 = n42590 & n42591;
  assign n42593 = ~n42589 & ~n42592;
  assign po614 = pi821 & ~n42593;
  assign n42595 = pi458 & ~n42121;
  assign n42596 = pi1072 & n42121;
  assign po615 = n42595 | n42596;
  assign n42598 = pi459 & ~n42441;
  assign n42599 = pi1058 & n42441;
  assign po616 = n42598 | n42599;
  assign n42601 = pi460 & ~n42121;
  assign n42602 = pi1086 & n42121;
  assign po617 = n42601 | n42602;
  assign n42604 = pi461 & ~n42121;
  assign n42605 = pi1057 & n42121;
  assign po618 = n42604 | n42605;
  assign n42607 = pi462 & ~n42121;
  assign n42608 = pi1074 & n42121;
  assign po619 = n42607 | n42608;
  assign n42610 = pi463 & ~n42133;
  assign n42611 = pi1070 & n42133;
  assign po620 = n42610 | n42611;
  assign n42613 = pi464 & ~n42441;
  assign n42614 = pi1065 & n42441;
  assign po621 = n42613 | n42614;
  assign n42616 = pi926 & n5728;
  assign n42617 = pi1157 & n5729;
  assign n42618 = ~pi243 & n42045;
  assign n42619 = ~n42616 & ~n42618;
  assign n42620 = ~n42617 & n42619;
  assign n42621 = po1038 & ~n42620;
  assign n42622 = ~pi243 & pi1157;
  assign n42623 = pi926 & n42622;
  assign n42624 = ~n11010 & n42623;
  assign n42625 = ~n10982 & ~n10985;
  assign n42626 = ~pi243 & ~n42625;
  assign n42627 = ~n5784 & ~n5802;
  assign n42628 = ~pi926 & ~n42627;
  assign n42629 = ~pi1157 & n42627;
  assign n42630 = ~pi299 & n42033;
  assign n42631 = pi299 & n2461;
  assign n42632 = ~n42630 & ~n42631;
  assign n42633 = ~n42622 & ~n42632;
  assign n42634 = ~n42628 & ~n42633;
  assign n42635 = ~n42629 & n42634;
  assign n42636 = ~n42626 & ~n42635;
  assign n42637 = ~po1038 & ~n42624;
  assign n42638 = ~n42636 & n42637;
  assign po622 = n42621 | n42638;
  assign n42640 = ~po1038 & n11008;
  assign n42641 = ~n42039 & ~n42640;
  assign n42642 = pi943 & ~n42641;
  assign n42643 = ~po1038 & ~n42625;
  assign n42644 = po1038 & n42045;
  assign n42645 = ~n42643 & ~n42644;
  assign n42646 = ~pi943 & ~n42645;
  assign n42647 = ~pi1151 & n42043;
  assign n42648 = ~n42646 & n42647;
  assign n42649 = ~n2461 & po1038;
  assign n42650 = ~po1038 & n42632;
  assign n42651 = ~n42649 & ~n42650;
  assign n42652 = ~pi275 & n42651;
  assign n42653 = ~pi943 & n42645;
  assign n42654 = ~n42043 & n42653;
  assign n42655 = ~n42642 & ~n42652;
  assign n42656 = ~n42654 & n42655;
  assign po623 = ~n42648 & n42656;
  assign n42658 = pi40 & ~pi287;
  assign n42659 = n39961 & n42658;
  assign n42660 = po950 & n42659;
  assign n42661 = ~n9781 & ~n42660;
  assign n42662 = ~pi102 & ~n12645;
  assign n42663 = n10960 & n15988;
  assign n42664 = ~n42662 & n42663;
  assign n42665 = n15986 & n42664;
  assign n42666 = ~n42659 & ~n42665;
  assign n42667 = n42659 & n42665;
  assign n42668 = ~n42666 & ~n42667;
  assign n42669 = n7425 & n42668;
  assign n42670 = ~n6104 & ~n42668;
  assign n42671 = n6104 & ~n42665;
  assign n42672 = ~n42670 & ~n42671;
  assign n42673 = ~n7425 & n42672;
  assign n42674 = pi1091 & ~n42669;
  assign n42675 = ~n42673 & n42674;
  assign n42676 = ~n7348 & ~n42668;
  assign n42677 = n7348 & ~n42665;
  assign n42678 = pi1093 & ~n42677;
  assign n42679 = ~n42676 & n42678;
  assign n42680 = ~pi1093 & n42672;
  assign n42681 = ~pi1091 & ~n42679;
  assign n42682 = ~n42680 & n42681;
  assign n42683 = ~n42675 & ~n42682;
  assign n42684 = n2616 & n12403;
  assign n42685 = ~n42683 & n42684;
  assign po624 = ~n42661 & ~n42685;
  assign n42687 = n9833 & n10924;
  assign n42688 = n9830 & n18596;
  assign n42689 = n7413 & n42688;
  assign n42690 = pi468 & ~n42689;
  assign po625 = n42687 | n42690;
  assign n42692 = pi942 & n5728;
  assign n42693 = pi1156 & n5729;
  assign n42694 = ~pi263 & n42045;
  assign n42695 = ~n42692 & ~n42694;
  assign n42696 = ~n42693 & n42695;
  assign n42697 = po1038 & ~n42696;
  assign n42698 = ~pi263 & pi1156;
  assign n42699 = pi942 & n42698;
  assign n42700 = ~n11010 & n42699;
  assign n42701 = ~pi263 & ~n42625;
  assign n42702 = ~pi942 & ~n42627;
  assign n42703 = ~pi1156 & n42627;
  assign n42704 = ~n42632 & ~n42698;
  assign n42705 = ~n42702 & ~n42704;
  assign n42706 = ~n42703 & n42705;
  assign n42707 = ~n42701 & ~n42706;
  assign n42708 = ~po1038 & ~n42700;
  assign n42709 = ~n42707 & n42708;
  assign po626 = n42697 | n42709;
  assign n42711 = pi925 & n5728;
  assign n42712 = pi1155 & n5729;
  assign n42713 = pi267 & n42045;
  assign n42714 = ~n42711 & ~n42713;
  assign n42715 = ~n42712 & n42714;
  assign n42716 = po1038 & ~n42715;
  assign n42717 = pi267 & pi1155;
  assign n42718 = pi925 & n42717;
  assign n42719 = ~n11010 & n42718;
  assign n42720 = pi267 & ~n42625;
  assign n42721 = ~pi925 & ~n42627;
  assign n42722 = ~pi1155 & n42627;
  assign n42723 = ~n42632 & ~n42717;
  assign n42724 = ~n42721 & ~n42723;
  assign n42725 = ~n42722 & n42724;
  assign n42726 = ~n42720 & ~n42725;
  assign n42727 = ~po1038 & ~n42719;
  assign n42728 = ~n42726 & n42727;
  assign po627 = n42716 | n42728;
  assign n42730 = pi941 & n5728;
  assign n42731 = pi1153 & n5729;
  assign n42732 = pi253 & n42045;
  assign n42733 = ~n42730 & ~n42732;
  assign n42734 = ~n42731 & n42733;
  assign n42735 = po1038 & ~n42734;
  assign n42736 = pi253 & pi1153;
  assign n42737 = pi941 & n42736;
  assign n42738 = ~n11010 & n42737;
  assign n42739 = pi253 & ~n42625;
  assign n42740 = ~pi941 & ~n42627;
  assign n42741 = ~pi1153 & n42627;
  assign n42742 = ~n42632 & ~n42736;
  assign n42743 = ~n42740 & ~n42742;
  assign n42744 = ~n42741 & n42743;
  assign n42745 = ~n42739 & ~n42744;
  assign n42746 = ~po1038 & ~n42738;
  assign n42747 = ~n42745 & n42746;
  assign po628 = n42735 | n42747;
  assign n42749 = pi923 & n5728;
  assign n42750 = pi1154 & n5729;
  assign n42751 = pi254 & n42045;
  assign n42752 = ~n42749 & ~n42751;
  assign n42753 = ~n42750 & n42752;
  assign n42754 = po1038 & ~n42753;
  assign n42755 = pi254 & pi1154;
  assign n42756 = pi923 & n42755;
  assign n42757 = ~n11010 & n42756;
  assign n42758 = pi254 & ~n42625;
  assign n42759 = ~pi923 & ~n42627;
  assign n42760 = ~pi1154 & n42627;
  assign n42761 = ~n42632 & ~n42755;
  assign n42762 = ~n42759 & ~n42761;
  assign n42763 = ~n42760 & n42762;
  assign n42764 = ~n42758 & ~n42763;
  assign n42765 = ~po1038 & ~n42757;
  assign n42766 = ~n42764 & n42765;
  assign po629 = n42754 | n42766;
  assign n42768 = pi922 & ~n42641;
  assign n42769 = ~pi922 & ~n42645;
  assign n42770 = ~pi1152 & n42043;
  assign n42771 = ~n42769 & n42770;
  assign n42772 = ~pi268 & n42651;
  assign n42773 = ~pi922 & n42645;
  assign n42774 = ~n42043 & n42773;
  assign n42775 = ~n42768 & ~n42772;
  assign n42776 = ~n42774 & n42775;
  assign po630 = ~n42771 & n42776;
  assign n42778 = pi931 & ~n42641;
  assign n42779 = ~pi931 & ~n42645;
  assign n42780 = ~pi1150 & n42043;
  assign n42781 = ~n42779 & n42780;
  assign n42782 = ~pi272 & n42651;
  assign n42783 = ~pi931 & n42645;
  assign n42784 = ~n42043 & n42783;
  assign n42785 = ~n42778 & ~n42782;
  assign n42786 = ~n42784 & n42785;
  assign po631 = ~n42781 & n42786;
  assign n42788 = pi936 & ~n42641;
  assign n42789 = ~pi936 & ~n42645;
  assign n42790 = ~pi1149 & n42043;
  assign n42791 = ~n42789 & n42790;
  assign n42792 = ~pi283 & n42651;
  assign n42793 = ~pi936 & n42645;
  assign n42794 = ~n42043 & n42793;
  assign n42795 = ~n42788 & ~n42792;
  assign n42796 = ~n42794 & n42795;
  assign po632 = ~n42791 & n42796;
  assign n42798 = pi71 & n41041;
  assign n42799 = pi71 & ~n11039;
  assign n42800 = n11039 & n12327;
  assign n42801 = n9788 & ~n11039;
  assign n42802 = n9785 & n42801;
  assign n42803 = ~n42800 & ~n42802;
  assign n42804 = n10880 & ~n42803;
  assign n42805 = n12332 & n42804;
  assign n42806 = ~n42799 & ~n42805;
  assign n42807 = ~po1038 & ~n42806;
  assign po633 = n42798 | n42807;
  assign po635 = pi71 & ~n41308;
  assign n42810 = pi481 & ~n33034;
  assign n42811 = pi248 & n33034;
  assign po638 = n42810 | n42811;
  assign n42813 = pi482 & ~n33050;
  assign n42814 = pi249 & n33050;
  assign po639 = n42813 | n42814;
  assign n42816 = pi483 & ~n33169;
  assign n42817 = pi242 & n33169;
  assign po640 = n42816 | n42817;
  assign n42819 = pi484 & ~n33169;
  assign n42820 = pi249 & n33169;
  assign po641 = n42819 | n42820;
  assign n42822 = pi485 & ~n34312;
  assign n42823 = pi234 & n34312;
  assign po642 = n42822 | n42823;
  assign n42825 = pi486 & ~n34312;
  assign n42826 = pi244 & n34312;
  assign po643 = n42825 | n42826;
  assign n42828 = pi487 & ~n33034;
  assign n42829 = pi246 & n33034;
  assign po644 = n42828 | n42829;
  assign n42831 = pi488 & ~n33034;
  assign n42832 = ~pi239 & n33034;
  assign po645 = ~n42831 & ~n42832;
  assign n42834 = pi489 & ~n34312;
  assign n42835 = pi242 & n34312;
  assign po646 = n42834 | n42835;
  assign n42837 = pi490 & ~n33169;
  assign n42838 = pi241 & n33169;
  assign po647 = n42837 | n42838;
  assign n42840 = pi491 & ~n33169;
  assign n42841 = pi238 & n33169;
  assign po648 = n42840 | n42841;
  assign n42843 = pi492 & ~n33169;
  assign n42844 = pi240 & n33169;
  assign po649 = n42843 | n42844;
  assign n42846 = pi493 & ~n33169;
  assign n42847 = pi244 & n33169;
  assign po650 = n42846 | n42847;
  assign n42849 = pi494 & ~n33169;
  assign n42850 = ~pi239 & n33169;
  assign po651 = ~n42849 & ~n42850;
  assign n42852 = pi495 & ~n33169;
  assign n42853 = pi235 & n33169;
  assign po652 = n42852 | n42853;
  assign n42855 = pi496 & ~n33161;
  assign n42856 = pi249 & n33161;
  assign po653 = n42855 | n42856;
  assign n42858 = pi497 & ~n33161;
  assign n42859 = ~pi239 & n33161;
  assign po654 = ~n42858 & ~n42859;
  assign n42861 = pi498 & ~n33050;
  assign n42862 = pi238 & n33050;
  assign po655 = n42861 | n42862;
  assign n42864 = pi499 & ~n33161;
  assign n42865 = pi246 & n33161;
  assign po656 = n42864 | n42865;
  assign n42867 = pi500 & ~n33161;
  assign n42868 = pi241 & n33161;
  assign po657 = n42867 | n42868;
  assign n42870 = pi501 & ~n33161;
  assign n42871 = pi248 & n33161;
  assign po658 = n42870 | n42871;
  assign n42873 = pi502 & ~n33161;
  assign n42874 = pi247 & n33161;
  assign po659 = n42873 | n42874;
  assign n42876 = pi503 & ~n33161;
  assign n42877 = pi245 & n33161;
  assign po660 = n42876 | n42877;
  assign n42879 = pi504 & ~n33154;
  assign n42880 = pi242 & n33154;
  assign po661 = n42879 | n42880;
  assign n42882 = pi505 & ~n33161;
  assign n42883 = pi234 & n33153;
  assign n42884 = n33037 & n42883;
  assign po662 = n42882 | n42884;
  assign n42886 = pi506 & ~n33154;
  assign n42887 = pi241 & n33154;
  assign po663 = n42886 | n42887;
  assign n42889 = pi507 & ~n33154;
  assign n42890 = pi238 & n33154;
  assign po664 = n42889 | n42890;
  assign n42892 = pi508 & ~n33154;
  assign n42893 = pi247 & n33154;
  assign po665 = n42892 | n42893;
  assign n42895 = pi509 & ~n33154;
  assign n42896 = pi245 & n33154;
  assign po666 = n42895 | n42896;
  assign n42898 = pi510 & ~n33034;
  assign n42899 = pi242 & n33034;
  assign po667 = n42898 | n42899;
  assign n42901 = n6536 & ~po1038;
  assign n42902 = ~n33028 & ~n42901;
  assign n42903 = ~pi234 & n42902;
  assign n42904 = n33034 & ~n42903;
  assign n42905 = pi511 & ~n33034;
  assign po668 = n42904 | n42905;
  assign n42907 = pi512 & ~n33034;
  assign n42908 = pi235 & n33034;
  assign po669 = n42907 | n42908;
  assign n42910 = pi513 & ~n33034;
  assign n42911 = pi244 & n33034;
  assign po670 = n42910 | n42911;
  assign n42913 = pi514 & ~n33034;
  assign n42914 = pi245 & n33034;
  assign po671 = n42913 | n42914;
  assign n42916 = pi515 & ~n33034;
  assign n42917 = pi240 & n33034;
  assign po672 = n42916 | n42917;
  assign n42919 = pi516 & ~n33034;
  assign n42920 = pi247 & n33034;
  assign po673 = n42919 | n42920;
  assign n42922 = pi517 & ~n33034;
  assign n42923 = pi238 & n33034;
  assign po674 = n42922 | n42923;
  assign n42925 = pi518 & ~n33042;
  assign n42926 = pi234 & n33033;
  assign n42927 = n33037 & n42926;
  assign po675 = n42925 | n42927;
  assign n42929 = pi519 & ~n33042;
  assign n42930 = ~pi239 & n33042;
  assign po676 = ~n42929 & ~n42930;
  assign n42932 = pi520 & ~n33042;
  assign n42933 = pi246 & n33042;
  assign po677 = n42932 | n42933;
  assign n42935 = pi521 & ~n33042;
  assign n42936 = pi248 & n33042;
  assign po678 = n42935 | n42936;
  assign n42938 = pi522 & ~n33042;
  assign n42939 = pi238 & n33042;
  assign po679 = n42938 | n42939;
  assign n42941 = pi523 & ~n34340;
  assign n42942 = n33164 & n42926;
  assign po680 = n42941 | n42942;
  assign n42944 = pi524 & ~n34340;
  assign n42945 = ~pi239 & n34340;
  assign po681 = ~n42944 & ~n42945;
  assign n42947 = pi525 & ~n34340;
  assign n42948 = pi245 & n34340;
  assign po682 = n42947 | n42948;
  assign n42950 = pi526 & ~n34340;
  assign n42951 = pi246 & n34340;
  assign po683 = n42950 | n42951;
  assign n42953 = pi527 & ~n34340;
  assign n42954 = pi247 & n34340;
  assign po684 = n42953 | n42954;
  assign n42956 = pi528 & ~n34340;
  assign n42957 = pi249 & n34340;
  assign po685 = n42956 | n42957;
  assign n42959 = pi529 & ~n34340;
  assign n42960 = pi238 & n34340;
  assign po686 = n42959 | n42960;
  assign n42962 = pi530 & ~n34340;
  assign n42963 = pi240 & n34340;
  assign po687 = n42962 | n42963;
  assign n42965 = pi531 & ~n33050;
  assign n42966 = pi235 & n33050;
  assign po688 = n42965 | n42966;
  assign n42968 = pi532 & ~n33050;
  assign n42969 = pi247 & n33050;
  assign po689 = n42968 | n42969;
  assign n42971 = pi533 & ~n33154;
  assign n42972 = pi235 & n33154;
  assign po690 = n42971 | n42972;
  assign n42974 = pi534 & ~n33154;
  assign n42975 = ~pi239 & n33154;
  assign po691 = ~n42974 & ~n42975;
  assign n42977 = pi535 & ~n33154;
  assign n42978 = pi240 & n33154;
  assign po692 = n42977 | n42978;
  assign n42980 = pi536 & ~n33154;
  assign n42981 = pi246 & n33154;
  assign po693 = n42980 | n42981;
  assign n42983 = pi537 & ~n33154;
  assign n42984 = pi248 & n33154;
  assign po694 = n42983 | n42984;
  assign n42986 = pi538 & ~n33154;
  assign n42987 = pi249 & n33154;
  assign po695 = n42986 | n42987;
  assign n42989 = pi539 & ~n33161;
  assign n42990 = pi242 & n33161;
  assign po696 = n42989 | n42990;
  assign n42992 = pi540 & ~n33161;
  assign n42993 = pi235 & n33161;
  assign po697 = n42992 | n42993;
  assign n42995 = pi541 & ~n33161;
  assign n42996 = pi244 & n33161;
  assign po698 = n42995 | n42996;
  assign n42998 = pi542 & ~n33161;
  assign n42999 = pi240 & n33161;
  assign po699 = n42998 | n42999;
  assign n43001 = pi543 & ~n33161;
  assign n43002 = pi238 & n33161;
  assign po700 = n43001 | n43002;
  assign n43004 = pi544 & ~n33169;
  assign n43005 = n33164 & n42883;
  assign po701 = n43004 | n43005;
  assign n43007 = pi545 & ~n33169;
  assign n43008 = pi245 & n33169;
  assign po702 = n43007 | n43008;
  assign n43010 = pi546 & ~n33169;
  assign n43011 = pi246 & n33169;
  assign po703 = n43010 | n43011;
  assign n43013 = pi547 & ~n33169;
  assign n43014 = pi247 & n33169;
  assign po704 = n43013 | n43014;
  assign n43016 = pi548 & ~n33169;
  assign n43017 = pi248 & n33169;
  assign po705 = n43016 | n43017;
  assign n43019 = pi549 & ~n34312;
  assign n43020 = pi235 & n34312;
  assign po706 = n43019 | n43020;
  assign n43022 = pi550 & ~n34312;
  assign n43023 = ~pi239 & n34312;
  assign po707 = ~n43022 & ~n43023;
  assign n43025 = pi551 & ~n34312;
  assign n43026 = pi240 & n34312;
  assign po708 = n43025 | n43026;
  assign n43028 = pi552 & ~n34312;
  assign n43029 = pi247 & n34312;
  assign po709 = n43028 | n43029;
  assign n43031 = pi553 & ~n34312;
  assign n43032 = pi241 & n34312;
  assign po710 = n43031 | n43032;
  assign n43034 = pi554 & ~n34312;
  assign n43035 = pi248 & n34312;
  assign po711 = n43034 | n43035;
  assign n43037 = pi555 & ~n34312;
  assign n43038 = pi249 & n34312;
  assign po712 = n43037 | n43038;
  assign n43040 = pi556 & ~n33050;
  assign n43041 = pi242 & n33050;
  assign po713 = n43040 | n43041;
  assign n43043 = pi557 & ~n33154;
  assign n43044 = n32850 & n42883;
  assign po714 = n43043 | n43044;
  assign n43046 = pi558 & ~n33154;
  assign n43047 = pi244 & n33154;
  assign po715 = n43046 | n43047;
  assign n43049 = pi559 & ~n33034;
  assign n43050 = pi241 & n33034;
  assign po716 = n43049 | n43050;
  assign n43052 = pi560 & ~n33050;
  assign n43053 = pi240 & n33050;
  assign po717 = n43052 | n43053;
  assign n43055 = pi561 & ~n33042;
  assign n43056 = pi247 & n33042;
  assign po718 = n43055 | n43056;
  assign n43058 = pi562 & ~n33050;
  assign n43059 = pi241 & n33050;
  assign po719 = n43058 | n43059;
  assign n43061 = pi563 & ~n34312;
  assign n43062 = pi246 & n34312;
  assign po720 = n43061 | n43062;
  assign n43064 = pi564 & ~n33050;
  assign n43065 = pi246 & n33050;
  assign po721 = n43064 | n43065;
  assign n43067 = pi565 & ~n33050;
  assign n43068 = pi248 & n33050;
  assign po722 = n43067 | n43068;
  assign n43070 = pi566 & ~n33050;
  assign n43071 = pi244 & n33050;
  assign po723 = n43070 | n43071;
  assign n43073 = ~pi567 & pi1092;
  assign n43074 = ~pi1093 & n43073;
  assign n43075 = pi680 & n16232;
  assign n43076 = ~n17581 & n43075;
  assign n43077 = ~n43074 & ~n43076;
  assign n43078 = n17586 & ~n43077;
  assign n43079 = ~n15765 & n43078;
  assign n43080 = ~n17768 & n43079;
  assign n43081 = ~n43074 & ~n43080;
  assign n43082 = pi644 & ~n43081;
  assign n43083 = pi647 & n43079;
  assign n43084 = pi1157 & ~n43074;
  assign n43085 = ~n43083 & n43084;
  assign n43086 = pi603 & n16486;
  assign n43087 = n18872 & n43086;
  assign n43088 = ~n15832 & n43087;
  assign n43089 = ~n15925 & n43088;
  assign n43090 = ~n43074 & ~n43089;
  assign n43091 = pi647 & ~n43090;
  assign n43092 = n22052 & ~n43077;
  assign n43093 = ~n43074 & ~n43087;
  assign n43094 = ~n43092 & n43093;
  assign n43095 = n15833 & ~n43094;
  assign n43096 = n22348 & ~n43093;
  assign n43097 = pi641 & n43092;
  assign n43098 = ~n43074 & ~n43097;
  assign n43099 = n15818 & ~n43098;
  assign n43100 = ~pi641 & n43092;
  assign n43101 = ~n43074 & ~n43100;
  assign n43102 = n15819 & ~n43101;
  assign n43103 = ~n43096 & ~n43099;
  assign n43104 = ~n43102 & n43103;
  assign n43105 = pi788 & ~n43104;
  assign n43106 = ~n43095 & ~n43105;
  assign n43107 = ~n16644 & ~n43106;
  assign n43108 = ~n43074 & ~n43088;
  assign n43109 = n15763 & ~n43108;
  assign n43110 = pi628 & n43078;
  assign n43111 = ~n43074 & ~n43110;
  assign n43112 = pi1156 & ~n43111;
  assign n43113 = ~pi629 & ~n43109;
  assign n43114 = ~n43112 & n43113;
  assign n43115 = n15762 & ~n43108;
  assign n43116 = ~pi628 & n43078;
  assign n43117 = ~n43074 & ~n43116;
  assign n43118 = ~pi1156 & ~n43117;
  assign n43119 = pi629 & ~n43115;
  assign n43120 = ~n43118 & n43119;
  assign n43121 = pi792 & ~n43114;
  assign n43122 = ~n43120 & n43121;
  assign n43123 = ~n43107 & ~n43122;
  assign n43124 = ~pi647 & ~n43123;
  assign n43125 = ~pi1157 & ~n43091;
  assign n43126 = ~n43124 & n43125;
  assign n43127 = ~pi630 & ~n43085;
  assign n43128 = ~n43126 & n43127;
  assign n43129 = ~pi647 & n43079;
  assign n43130 = ~pi1157 & ~n43074;
  assign n43131 = ~n43129 & n43130;
  assign n43132 = ~pi647 & ~n43090;
  assign n43133 = pi647 & ~n43123;
  assign n43134 = pi1157 & ~n43132;
  assign n43135 = ~n43133 & n43134;
  assign n43136 = pi630 & ~n43131;
  assign n43137 = ~n43135 & n43136;
  assign n43138 = ~n43128 & ~n43137;
  assign n43139 = pi787 & ~n43138;
  assign n43140 = ~pi787 & ~n43123;
  assign n43141 = ~n43139 & ~n43140;
  assign n43142 = ~pi644 & ~n43141;
  assign n43143 = ~pi715 & ~n43082;
  assign n43144 = ~n43142 & n43143;
  assign n43145 = n19771 & ~n43108;
  assign n43146 = ~pi644 & n43145;
  assign n43147 = pi715 & ~n43074;
  assign n43148 = ~n43146 & n43147;
  assign n43149 = ~pi1160 & ~n43148;
  assign n43150 = ~n43144 & n43149;
  assign n43151 = pi644 & ~n43141;
  assign n43152 = ~pi644 & ~n43081;
  assign n43153 = pi715 & ~n43152;
  assign n43154 = ~n43151 & n43153;
  assign n43155 = pi644 & n43145;
  assign n43156 = ~pi715 & ~n43074;
  assign n43157 = ~n43155 & n43156;
  assign n43158 = pi1160 & ~n43157;
  assign n43159 = ~n43154 & n43158;
  assign n43160 = ~n43150 & ~n43159;
  assign n43161 = pi790 & ~n43160;
  assign n43162 = ~pi790 & ~n43141;
  assign n43163 = ~n43161 & ~n43162;
  assign n43164 = pi230 & ~n43163;
  assign n43165 = ~pi230 & n43073;
  assign po724 = n43164 | n43165;
  assign n43167 = pi568 & ~n33050;
  assign n43168 = pi245 & n33050;
  assign po725 = n43167 | n43168;
  assign n43170 = pi569 & ~n33050;
  assign n43171 = ~pi239 & n33050;
  assign po726 = ~n43170 & ~n43171;
  assign n43173 = pi570 & ~n33050;
  assign n43174 = n33045 & n42926;
  assign po727 = n43173 | n43174;
  assign n43176 = pi571 & ~n34340;
  assign n43177 = pi241 & n34340;
  assign po728 = n43176 | n43177;
  assign n43179 = pi572 & ~n34340;
  assign n43180 = pi244 & n34340;
  assign po729 = n43179 | n43180;
  assign n43182 = pi573 & ~n34340;
  assign n43183 = pi242 & n34340;
  assign po730 = n43182 | n43183;
  assign n43185 = pi574 & ~n33042;
  assign n43186 = pi241 & n33042;
  assign po731 = n43185 | n43186;
  assign n43188 = pi575 & ~n34340;
  assign n43189 = pi235 & n34340;
  assign po732 = n43188 | n43189;
  assign n43191 = pi576 & ~n34340;
  assign n43192 = pi248 & n34340;
  assign po733 = n43191 | n43192;
  assign n43194 = pi577 & ~n34312;
  assign n43195 = pi238 & n34312;
  assign po734 = n43194 | n43195;
  assign n43197 = pi578 & ~n33042;
  assign n43198 = pi249 & n33042;
  assign po735 = n43197 | n43198;
  assign n43200 = pi579 & ~n33034;
  assign n43201 = pi249 & n33034;
  assign po736 = n43200 | n43201;
  assign n43203 = pi580 & ~n34312;
  assign n43204 = pi245 & n34312;
  assign po737 = n43203 | n43204;
  assign n43206 = pi581 & ~n33042;
  assign n43207 = pi235 & n33042;
  assign po738 = n43206 | n43207;
  assign n43209 = pi582 & ~n33042;
  assign n43210 = pi240 & n33042;
  assign po739 = n43209 | n43210;
  assign n43212 = pi584 & ~n33042;
  assign n43213 = pi245 & n33042;
  assign po741 = n43212 | n43213;
  assign n43215 = pi585 & ~n33042;
  assign n43216 = pi244 & n33042;
  assign po742 = n43215 | n43216;
  assign n43218 = pi586 & ~n33042;
  assign n43219 = pi242 & n33042;
  assign po743 = n43218 | n43219;
  assign n43221 = ~pi230 & pi587;
  assign n43222 = pi230 & n15780;
  assign n43223 = ~n33800 & n43222;
  assign n43224 = n18872 & n43223;
  assign n43225 = n28954 & n43224;
  assign po744 = n43221 | n43225;
  assign n43227 = ~pi123 & n11855;
  assign n43228 = ~pi588 & ~n43227;
  assign n43229 = ~pi591 & n43227;
  assign n43230 = n42170 & ~n43228;
  assign po745 = ~n43229 & n43230;
  assign n43232 = ~n6279 & n15574;
  assign n43233 = ~n33149 & ~n43232;
  assign n43234 = ~pi205 & n43233;
  assign n43235 = ~pi202 & n42902;
  assign n43236 = ~pi233 & ~n43234;
  assign n43237 = ~n43235 & n43236;
  assign n43238 = ~pi204 & n43233;
  assign n43239 = ~pi201 & n42902;
  assign n43240 = pi233 & ~n43238;
  assign n43241 = ~n43239 & n43240;
  assign n43242 = ~n43237 & ~n43241;
  assign n43243 = pi237 & ~n43242;
  assign n43244 = ~pi218 & n43233;
  assign n43245 = ~pi203 & n42902;
  assign n43246 = ~pi233 & ~n43244;
  assign n43247 = ~n43245 & n43246;
  assign n43248 = ~pi206 & n43233;
  assign n43249 = ~pi220 & n42902;
  assign n43250 = pi233 & ~n43248;
  assign n43251 = ~n43249 & n43250;
  assign n43252 = ~n43247 & ~n43251;
  assign n43253 = ~pi237 & ~n43252;
  assign po746 = ~n43243 & ~n43253;
  assign n43255 = pi588 & n43227;
  assign n43256 = pi590 & ~n43227;
  assign n43257 = n42170 & ~n43255;
  assign po747 = n43256 | ~n43257;
  assign n43259 = ~pi591 & ~n43227;
  assign n43260 = ~pi592 & n43227;
  assign n43261 = n42170 & ~n43259;
  assign po748 = ~n43260 & n43261;
  assign n43263 = ~pi592 & ~n43227;
  assign n43264 = ~pi590 & n43227;
  assign n43265 = n42170 & ~n43263;
  assign po749 = ~n43264 & n43265;
  assign n43267 = ~pi248 & pi521;
  assign n43268 = ~pi240 & pi582;
  assign n43269 = ~pi239 & ~pi519;
  assign n43270 = pi240 & ~pi582;
  assign n43271 = pi247 & ~pi561;
  assign n43272 = ~pi247 & pi561;
  assign n43273 = ~pi245 & ~pi584;
  assign n43274 = pi245 & pi584;
  assign n43275 = ~n43273 & ~n43274;
  assign n43276 = pi241 & ~pi574;
  assign n43277 = ~pi241 & pi574;
  assign n43278 = pi246 & ~pi520;
  assign n43279 = ~pi246 & pi520;
  assign n43280 = ~pi249 & pi578;
  assign n43281 = pi244 & ~pi585;
  assign n43282 = pi249 & ~pi578;
  assign n43283 = ~pi235 & pi581;
  assign n43284 = ~pi244 & pi585;
  assign n43285 = pi235 & ~pi581;
  assign n43286 = pi242 & ~pi586;
  assign n43287 = pi239 & pi519;
  assign n43288 = ~pi518 & n42903;
  assign n43289 = pi234 & n42902;
  assign n43290 = pi518 & n43289;
  assign n43291 = ~n43288 & ~n43290;
  assign n43292 = pi248 & ~pi521;
  assign n43293 = ~pi242 & pi586;
  assign n43294 = ~n43267 & ~n43268;
  assign n43295 = ~n43269 & ~n43270;
  assign n43296 = ~n43271 & ~n43272;
  assign n43297 = ~n43276 & ~n43277;
  assign n43298 = ~n43278 & ~n43279;
  assign n43299 = ~n43280 & ~n43281;
  assign n43300 = ~n43282 & ~n43283;
  assign n43301 = ~n43284 & ~n43285;
  assign n43302 = ~n43286 & ~n43287;
  assign n43303 = ~n43292 & ~n43293;
  assign n43304 = n43302 & n43303;
  assign n43305 = n43300 & n43301;
  assign n43306 = n43298 & n43299;
  assign n43307 = n43296 & n43297;
  assign n43308 = n43294 & n43295;
  assign n43309 = ~n43275 & n43308;
  assign n43310 = n43306 & n43307;
  assign n43311 = n43304 & n43305;
  assign n43312 = n43310 & n43311;
  assign n43313 = n43309 & n43312;
  assign n43314 = ~n43291 & n43313;
  assign n43315 = ~pi522 & n43314;
  assign n43316 = ~pi249 & pi496;
  assign n43317 = pi246 & ~pi499;
  assign n43318 = ~pi246 & pi499;
  assign n43319 = pi241 & ~pi500;
  assign n43320 = pi249 & ~pi496;
  assign n43321 = ~n43316 & ~n43317;
  assign n43322 = ~n43318 & ~n43319;
  assign n43323 = ~n43320 & n43322;
  assign n43324 = n43321 & n43323;
  assign n43325 = ~pi245 & ~pi503;
  assign n43326 = pi245 & pi503;
  assign n43327 = ~n43325 & ~n43326;
  assign n43328 = ~pi248 & pi501;
  assign n43329 = ~pi235 & pi540;
  assign n43330 = ~pi242 & pi539;
  assign n43331 = pi235 & ~pi540;
  assign n43332 = pi240 & ~pi542;
  assign n43333 = ~pi241 & pi500;
  assign n43334 = ~pi234 & n43233;
  assign n43335 = ~pi505 & n43334;
  assign n43336 = pi234 & n43233;
  assign n43337 = pi505 & n43336;
  assign n43338 = ~n43335 & ~n43337;
  assign n43339 = pi248 & ~pi501;
  assign n43340 = ~pi240 & pi542;
  assign n43341 = pi239 & pi497;
  assign n43342 = pi242 & ~pi539;
  assign n43343 = ~pi239 & ~pi497;
  assign n43344 = pi244 & ~pi541;
  assign n43345 = ~pi244 & pi541;
  assign n43346 = pi247 & ~pi502;
  assign n43347 = ~pi247 & pi502;
  assign n43348 = ~n43328 & ~n43329;
  assign n43349 = ~n43330 & ~n43331;
  assign n43350 = ~n43332 & ~n43333;
  assign n43351 = ~n43339 & ~n43340;
  assign n43352 = ~n43341 & ~n43342;
  assign n43353 = ~n43343 & ~n43344;
  assign n43354 = ~n43345 & ~n43346;
  assign n43355 = ~n43347 & n43354;
  assign n43356 = n43352 & n43353;
  assign n43357 = n43350 & n43351;
  assign n43358 = n43348 & n43349;
  assign n43359 = ~n43327 & n43358;
  assign n43360 = n43356 & n43357;
  assign n43361 = n43355 & n43360;
  assign n43362 = n43359 & n43361;
  assign n43363 = ~n43338 & n43362;
  assign n43364 = ~pi543 & n43324;
  assign n43365 = n43363 & n43364;
  assign n43366 = ~pi238 & ~n43315;
  assign n43367 = ~n43365 & n43366;
  assign n43368 = pi522 & n43314;
  assign n43369 = pi543 & n43324;
  assign n43370 = n43363 & n43369;
  assign n43371 = pi238 & ~n43368;
  assign n43372 = ~n43370 & n43371;
  assign n43373 = ~pi233 & ~n43367;
  assign n43374 = ~n43372 & n43373;
  assign n43375 = ~pi240 & ~pi535;
  assign n43376 = pi240 & pi535;
  assign n43377 = ~n43375 & ~n43376;
  assign n43378 = pi557 & ~n43336;
  assign n43379 = pi246 & ~pi536;
  assign n43380 = ~pi246 & pi536;
  assign n43381 = ~pi248 & ~pi537;
  assign n43382 = pi248 & pi537;
  assign n43383 = ~n43381 & ~n43382;
  assign n43384 = pi249 & ~pi538;
  assign n43385 = ~pi249 & pi538;
  assign n43386 = ~pi557 & ~n43334;
  assign n43387 = ~n43379 & ~n43380;
  assign n43388 = ~n43384 & ~n43385;
  assign n43389 = n43387 & n43388;
  assign n43390 = ~n43383 & n43389;
  assign n43391 = ~n43378 & n43390;
  assign n43392 = ~n43386 & n43391;
  assign n43393 = ~pi241 & ~pi506;
  assign n43394 = pi241 & pi506;
  assign n43395 = ~n43393 & ~n43394;
  assign n43396 = n43392 & ~n43395;
  assign n43397 = ~n43377 & n43396;
  assign n43398 = pi534 & n43397;
  assign n43399 = ~pi239 & ~n43398;
  assign n43400 = ~pi534 & n43397;
  assign n43401 = pi239 & ~n43400;
  assign n43402 = ~n43399 & ~n43401;
  assign n43403 = pi504 & n43402;
  assign n43404 = pi242 & ~n43403;
  assign n43405 = ~pi504 & n43402;
  assign n43406 = ~pi242 & ~n43405;
  assign n43407 = ~n43404 & ~n43406;
  assign n43408 = pi533 & n43407;
  assign n43409 = pi235 & ~n43408;
  assign n43410 = ~pi533 & n43407;
  assign n43411 = ~pi235 & ~n43410;
  assign n43412 = ~n43409 & ~n43411;
  assign n43413 = pi558 & n43412;
  assign n43414 = pi244 & ~n43413;
  assign n43415 = ~pi558 & n43412;
  assign n43416 = ~pi244 & ~n43415;
  assign n43417 = ~n43414 & ~n43416;
  assign n43418 = pi509 & n43417;
  assign n43419 = pi245 & ~n43418;
  assign n43420 = ~pi509 & n43417;
  assign n43421 = ~pi245 & ~n43420;
  assign n43422 = ~n43419 & ~n43421;
  assign n43423 = pi508 & n43422;
  assign n43424 = pi247 & ~n43423;
  assign n43425 = ~pi508 & n43422;
  assign n43426 = ~pi247 & ~n43425;
  assign n43427 = ~n43424 & ~n43426;
  assign n43428 = ~pi238 & n43427;
  assign n43429 = pi511 & ~n43289;
  assign n43430 = pi246 & ~pi487;
  assign n43431 = ~pi246 & pi487;
  assign n43432 = ~pi248 & ~pi481;
  assign n43433 = pi248 & pi481;
  assign n43434 = ~n43432 & ~n43433;
  assign n43435 = pi249 & ~pi579;
  assign n43436 = ~pi249 & pi579;
  assign n43437 = ~pi511 & ~n42903;
  assign n43438 = ~n43430 & ~n43431;
  assign n43439 = ~n43435 & ~n43436;
  assign n43440 = n43438 & n43439;
  assign n43441 = ~n43434 & n43440;
  assign n43442 = ~n43429 & n43441;
  assign n43443 = ~n43437 & n43442;
  assign n43444 = pi559 & n43443;
  assign n43445 = pi241 & ~n43444;
  assign n43446 = ~pi559 & n43443;
  assign n43447 = ~pi241 & ~n43446;
  assign n43448 = ~n43445 & ~n43447;
  assign n43449 = pi515 & n43448;
  assign n43450 = pi240 & ~n43449;
  assign n43451 = ~pi515 & n43448;
  assign n43452 = ~pi240 & ~n43451;
  assign n43453 = ~n43450 & ~n43452;
  assign n43454 = pi239 & ~pi488;
  assign n43455 = ~pi239 & pi488;
  assign n43456 = ~n43454 & ~n43455;
  assign n43457 = n43453 & ~n43456;
  assign n43458 = ~pi242 & ~pi510;
  assign n43459 = pi242 & pi510;
  assign n43460 = ~n43458 & ~n43459;
  assign n43461 = n43457 & ~n43460;
  assign n43462 = ~pi235 & ~pi512;
  assign n43463 = pi235 & pi512;
  assign n43464 = ~n43462 & ~n43463;
  assign n43465 = n43461 & ~n43464;
  assign n43466 = ~pi244 & ~pi513;
  assign n43467 = pi244 & pi513;
  assign n43468 = ~n43466 & ~n43467;
  assign n43469 = n43465 & ~n43468;
  assign n43470 = ~pi245 & ~pi514;
  assign n43471 = pi245 & pi514;
  assign n43472 = ~n43470 & ~n43471;
  assign n43473 = n43469 & ~n43472;
  assign n43474 = ~pi247 & ~pi516;
  assign n43475 = pi247 & pi516;
  assign n43476 = ~n43474 & ~n43475;
  assign n43477 = n43473 & ~n43476;
  assign n43478 = pi238 & n43477;
  assign n43479 = pi517 & ~n43478;
  assign n43480 = ~n43428 & n43479;
  assign n43481 = ~n43396 & n43447;
  assign n43482 = ~n43445 & ~n43481;
  assign n43483 = pi506 & n43392;
  assign n43484 = ~n43447 & n43483;
  assign n43485 = ~n43482 & ~n43484;
  assign n43486 = ~pi515 & ~n43485;
  assign n43487 = pi515 & n43396;
  assign n43488 = ~pi240 & ~n43487;
  assign n43489 = ~n43486 & n43488;
  assign n43490 = ~n43450 & ~n43489;
  assign n43491 = ~pi535 & ~n43490;
  assign n43492 = pi515 & ~n43485;
  assign n43493 = ~pi515 & n43396;
  assign n43494 = pi240 & ~n43493;
  assign n43495 = ~n43492 & n43494;
  assign n43496 = ~n43452 & ~n43495;
  assign n43497 = pi535 & ~n43496;
  assign n43498 = ~n43491 & ~n43497;
  assign n43499 = ~pi534 & n43498;
  assign n43500 = pi534 & n43453;
  assign n43501 = pi239 & ~n43500;
  assign n43502 = ~n43499 & n43501;
  assign n43503 = ~n43399 & ~n43502;
  assign n43504 = ~pi488 & ~n43503;
  assign n43505 = pi534 & n43498;
  assign n43506 = ~pi534 & n43453;
  assign n43507 = ~pi239 & ~n43506;
  assign n43508 = ~n43505 & n43507;
  assign n43509 = ~n43401 & ~n43508;
  assign n43510 = pi488 & ~n43509;
  assign n43511 = ~n43504 & ~n43510;
  assign n43512 = ~pi504 & n43511;
  assign n43513 = pi504 & n43457;
  assign n43514 = ~pi242 & ~n43513;
  assign n43515 = ~n43512 & n43514;
  assign n43516 = ~n43404 & ~n43515;
  assign n43517 = ~pi510 & ~n43516;
  assign n43518 = pi504 & n43511;
  assign n43519 = ~pi504 & n43457;
  assign n43520 = pi242 & ~n43519;
  assign n43521 = ~n43518 & n43520;
  assign n43522 = ~n43406 & ~n43521;
  assign n43523 = pi510 & ~n43522;
  assign n43524 = ~n43517 & ~n43523;
  assign n43525 = ~pi533 & n43524;
  assign n43526 = pi533 & n43461;
  assign n43527 = ~pi235 & ~n43526;
  assign n43528 = ~n43525 & n43527;
  assign n43529 = ~n43409 & ~n43528;
  assign n43530 = ~pi512 & ~n43529;
  assign n43531 = pi533 & n43524;
  assign n43532 = ~pi533 & n43461;
  assign n43533 = pi235 & ~n43532;
  assign n43534 = ~n43531 & n43533;
  assign n43535 = ~n43411 & ~n43534;
  assign n43536 = pi512 & ~n43535;
  assign n43537 = ~n43530 & ~n43536;
  assign n43538 = ~pi558 & n43537;
  assign n43539 = pi558 & n43465;
  assign n43540 = ~pi244 & ~n43539;
  assign n43541 = ~n43538 & n43540;
  assign n43542 = ~n43414 & ~n43541;
  assign n43543 = ~pi513 & ~n43542;
  assign n43544 = pi558 & n43537;
  assign n43545 = ~pi558 & n43465;
  assign n43546 = pi244 & ~n43545;
  assign n43547 = ~n43544 & n43546;
  assign n43548 = ~n43416 & ~n43547;
  assign n43549 = pi513 & ~n43548;
  assign n43550 = ~n43543 & ~n43549;
  assign n43551 = ~pi509 & n43550;
  assign n43552 = pi509 & n43469;
  assign n43553 = ~pi245 & ~n43552;
  assign n43554 = ~n43551 & n43553;
  assign n43555 = ~n43419 & ~n43554;
  assign n43556 = ~pi514 & ~n43555;
  assign n43557 = pi509 & n43550;
  assign n43558 = ~pi509 & n43469;
  assign n43559 = pi245 & ~n43558;
  assign n43560 = ~n43557 & n43559;
  assign n43561 = ~n43421 & ~n43560;
  assign n43562 = pi514 & ~n43561;
  assign n43563 = ~n43556 & ~n43562;
  assign n43564 = ~pi508 & n43563;
  assign n43565 = pi508 & n43473;
  assign n43566 = ~pi247 & ~n43565;
  assign n43567 = ~n43564 & n43566;
  assign n43568 = ~n43424 & ~n43567;
  assign n43569 = ~pi516 & ~n43568;
  assign n43570 = pi508 & n43563;
  assign n43571 = ~pi508 & n43473;
  assign n43572 = pi247 & ~n43571;
  assign n43573 = ~n43570 & n43572;
  assign n43574 = ~n43426 & ~n43573;
  assign n43575 = pi516 & ~n43574;
  assign n43576 = ~n43569 & ~n43575;
  assign n43577 = ~pi238 & n43576;
  assign n43578 = ~pi517 & ~n43577;
  assign n43579 = ~pi507 & ~n43480;
  assign n43580 = ~n43578 & n43579;
  assign n43581 = pi238 & n43427;
  assign n43582 = ~pi238 & n43477;
  assign n43583 = ~pi517 & ~n43582;
  assign n43584 = ~n43581 & n43583;
  assign n43585 = pi238 & n43576;
  assign n43586 = pi517 & ~n43585;
  assign n43587 = pi507 & ~n43584;
  assign n43588 = ~n43586 & n43587;
  assign n43589 = ~n43580 & ~n43588;
  assign n43590 = pi233 & ~n43589;
  assign n43591 = pi237 & ~n43374;
  assign n43592 = ~n43590 & n43591;
  assign n43593 = pi485 & ~n43336;
  assign n43594 = ~pi235 & ~pi549;
  assign n43595 = pi235 & pi549;
  assign n43596 = ~n43594 & ~n43595;
  assign n43597 = ~pi241 & pi553;
  assign n43598 = ~pi245 & pi580;
  assign n43599 = pi241 & ~pi553;
  assign n43600 = ~pi239 & ~pi550;
  assign n43601 = pi239 & pi550;
  assign n43602 = pi242 & ~pi489;
  assign n43603 = ~pi242 & pi489;
  assign n43604 = pi244 & ~pi486;
  assign n43605 = ~pi244 & pi486;
  assign n43606 = ~pi248 & pi554;
  assign n43607 = pi245 & ~pi580;
  assign n43608 = pi246 & ~pi563;
  assign n43609 = ~pi246 & pi563;
  assign n43610 = ~pi247 & ~pi552;
  assign n43611 = pi247 & pi552;
  assign n43612 = ~n43610 & ~n43611;
  assign n43613 = ~pi485 & ~n43334;
  assign n43614 = ~n43597 & ~n43598;
  assign n43615 = ~n43599 & ~n43600;
  assign n43616 = ~n43601 & ~n43602;
  assign n43617 = ~n43603 & ~n43604;
  assign n43618 = ~n43605 & ~n43606;
  assign n43619 = ~n43607 & ~n43608;
  assign n43620 = ~n43609 & n43619;
  assign n43621 = n43617 & n43618;
  assign n43622 = n43615 & n43616;
  assign n43623 = ~n43596 & n43614;
  assign n43624 = ~n43612 & n43623;
  assign n43625 = n43621 & n43622;
  assign n43626 = n43620 & n43625;
  assign n43627 = n43624 & n43626;
  assign n43628 = ~n43593 & n43627;
  assign n43629 = ~n43613 & n43628;
  assign n43630 = pi240 & ~pi551;
  assign n43631 = ~pi240 & pi551;
  assign n43632 = pi248 & ~pi554;
  assign n43633 = ~pi249 & ~pi555;
  assign n43634 = pi249 & pi555;
  assign n43635 = ~n43633 & ~n43634;
  assign n43636 = ~n43630 & ~n43631;
  assign n43637 = ~n43632 & n43636;
  assign n43638 = ~n43635 & n43637;
  assign n43639 = ~pi577 & n43638;
  assign n43640 = n43629 & n43639;
  assign n43641 = ~pi245 & ~pi568;
  assign n43642 = pi245 & pi568;
  assign n43643 = ~n43641 & ~n43642;
  assign n43644 = ~pi246 & ~pi564;
  assign n43645 = pi246 & pi564;
  assign n43646 = ~n43644 & ~n43645;
  assign n43647 = ~pi235 & pi531;
  assign n43648 = pi242 & ~pi556;
  assign n43649 = ~pi248 & pi565;
  assign n43650 = ~pi249 & pi482;
  assign n43651 = ~pi241 & ~pi562;
  assign n43652 = pi241 & pi562;
  assign n43653 = ~n43651 & ~n43652;
  assign n43654 = pi244 & ~pi566;
  assign n43655 = ~pi244 & pi566;
  assign n43656 = pi240 & ~pi560;
  assign n43657 = ~pi240 & pi560;
  assign n43658 = ~pi239 & ~pi569;
  assign n43659 = pi249 & ~pi482;
  assign n43660 = pi248 & ~pi565;
  assign n43661 = pi570 & ~n43289;
  assign n43662 = pi239 & pi569;
  assign n43663 = pi235 & ~pi531;
  assign n43664 = ~pi570 & ~n42903;
  assign n43665 = ~pi242 & pi556;
  assign n43666 = ~n43647 & ~n43648;
  assign n43667 = ~n43649 & ~n43650;
  assign n43668 = ~n43654 & ~n43655;
  assign n43669 = ~n43656 & ~n43657;
  assign n43670 = ~n43658 & ~n43659;
  assign n43671 = ~n43660 & ~n43662;
  assign n43672 = ~n43663 & ~n43665;
  assign n43673 = n43671 & n43672;
  assign n43674 = n43669 & n43670;
  assign n43675 = n43667 & n43668;
  assign n43676 = ~n43643 & n43666;
  assign n43677 = ~n43646 & ~n43653;
  assign n43678 = n43676 & n43677;
  assign n43679 = n43674 & n43675;
  assign n43680 = n43673 & n43679;
  assign n43681 = n43678 & n43680;
  assign n43682 = ~n43661 & n43681;
  assign n43683 = ~n43664 & n43682;
  assign n43684 = pi247 & ~pi532;
  assign n43685 = ~pi247 & pi532;
  assign n43686 = ~n43684 & ~n43685;
  assign n43687 = ~pi498 & n43686;
  assign n43688 = n43683 & n43687;
  assign n43689 = ~pi238 & ~n43640;
  assign n43690 = ~n43688 & n43689;
  assign n43691 = pi577 & n43638;
  assign n43692 = n43629 & n43691;
  assign n43693 = pi498 & n43686;
  assign n43694 = n43683 & n43693;
  assign n43695 = pi238 & ~n43692;
  assign n43696 = ~n43694 & n43695;
  assign n43697 = ~pi233 & ~n43690;
  assign n43698 = ~n43696 & n43697;
  assign n43699 = ~pi246 & pi526;
  assign n43700 = ~pi241 & ~pi571;
  assign n43701 = pi241 & pi571;
  assign n43702 = ~n43700 & ~n43701;
  assign n43703 = ~pi240 & pi530;
  assign n43704 = pi523 & ~n43289;
  assign n43705 = pi240 & ~pi530;
  assign n43706 = pi248 & ~pi576;
  assign n43707 = ~pi248 & pi576;
  assign n43708 = pi235 & ~pi575;
  assign n43709 = ~pi235 & pi575;
  assign n43710 = ~pi249 & ~pi528;
  assign n43711 = pi249 & pi528;
  assign n43712 = ~n43710 & ~n43711;
  assign n43713 = pi239 & pi524;
  assign n43714 = ~pi242 & pi573;
  assign n43715 = ~pi523 & ~n42903;
  assign n43716 = ~pi239 & ~pi524;
  assign n43717 = pi242 & ~pi573;
  assign n43718 = pi246 & ~pi526;
  assign n43719 = ~n43699 & ~n43703;
  assign n43720 = ~n43705 & ~n43706;
  assign n43721 = ~n43707 & ~n43708;
  assign n43722 = ~n43709 & ~n43713;
  assign n43723 = ~n43714 & ~n43716;
  assign n43724 = ~n43717 & ~n43718;
  assign n43725 = n43723 & n43724;
  assign n43726 = n43721 & n43722;
  assign n43727 = n43719 & n43720;
  assign n43728 = ~n43702 & ~n43712;
  assign n43729 = n43727 & n43728;
  assign n43730 = n43725 & n43726;
  assign n43731 = n43729 & n43730;
  assign n43732 = ~n43704 & n43731;
  assign n43733 = ~n43715 & n43732;
  assign n43734 = ~pi572 & n43733;
  assign n43735 = ~pi244 & ~n43734;
  assign n43736 = pi572 & n43733;
  assign n43737 = pi244 & ~n43736;
  assign n43738 = ~n43735 & ~n43737;
  assign n43739 = ~pi245 & ~pi525;
  assign n43740 = pi245 & pi525;
  assign n43741 = ~n43739 & ~n43740;
  assign n43742 = n43738 & ~n43741;
  assign n43743 = ~pi247 & ~pi527;
  assign n43744 = pi247 & pi527;
  assign n43745 = ~n43743 & ~n43744;
  assign n43746 = n43742 & ~n43745;
  assign n43747 = pi238 & n43746;
  assign n43748 = pi544 & ~n43336;
  assign n43749 = ~pi240 & pi492;
  assign n43750 = ~pi242 & pi483;
  assign n43751 = pi240 & ~pi492;
  assign n43752 = pi246 & ~pi546;
  assign n43753 = ~pi246 & pi546;
  assign n43754 = pi235 & ~pi495;
  assign n43755 = ~pi235 & pi495;
  assign n43756 = ~pi248 & ~pi548;
  assign n43757 = pi248 & pi548;
  assign n43758 = ~n43756 & ~n43757;
  assign n43759 = pi241 & ~pi490;
  assign n43760 = ~pi241 & pi490;
  assign n43761 = pi249 & ~pi484;
  assign n43762 = ~pi249 & pi484;
  assign n43763 = pi242 & ~pi483;
  assign n43764 = ~pi239 & ~pi494;
  assign n43765 = pi239 & pi494;
  assign n43766 = ~pi544 & ~n43334;
  assign n43767 = ~n43749 & ~n43750;
  assign n43768 = ~n43751 & ~n43752;
  assign n43769 = ~n43753 & ~n43754;
  assign n43770 = ~n43755 & ~n43759;
  assign n43771 = ~n43760 & ~n43761;
  assign n43772 = ~n43762 & ~n43763;
  assign n43773 = ~n43764 & ~n43765;
  assign n43774 = n43772 & n43773;
  assign n43775 = n43770 & n43771;
  assign n43776 = n43768 & n43769;
  assign n43777 = ~n43758 & n43767;
  assign n43778 = n43776 & n43777;
  assign n43779 = n43774 & n43775;
  assign n43780 = n43778 & n43779;
  assign n43781 = ~n43748 & n43780;
  assign n43782 = ~n43766 & n43781;
  assign n43783 = ~pi244 & ~pi493;
  assign n43784 = pi244 & pi493;
  assign n43785 = ~n43783 & ~n43784;
  assign n43786 = n43782 & ~n43785;
  assign n43787 = pi545 & n43786;
  assign n43788 = pi245 & ~n43787;
  assign n43789 = ~pi545 & n43786;
  assign n43790 = ~pi245 & ~n43789;
  assign n43791 = ~n43788 & ~n43790;
  assign n43792 = pi547 & n43791;
  assign n43793 = pi247 & ~n43792;
  assign n43794 = ~pi547 & n43791;
  assign n43795 = ~pi247 & ~n43794;
  assign n43796 = ~n43793 & ~n43795;
  assign n43797 = ~pi238 & n43796;
  assign n43798 = pi529 & ~n43747;
  assign n43799 = ~n43797 & n43798;
  assign n43800 = n43735 & ~n43786;
  assign n43801 = ~n43737 & ~n43800;
  assign n43802 = pi493 & n43782;
  assign n43803 = ~n43735 & n43802;
  assign n43804 = ~n43801 & ~n43803;
  assign n43805 = ~pi545 & ~n43804;
  assign n43806 = pi545 & n43738;
  assign n43807 = ~pi245 & ~n43806;
  assign n43808 = ~n43805 & n43807;
  assign n43809 = ~n43788 & ~n43808;
  assign n43810 = ~pi525 & ~n43809;
  assign n43811 = pi545 & ~n43804;
  assign n43812 = ~pi545 & n43738;
  assign n43813 = pi245 & ~n43812;
  assign n43814 = ~n43811 & n43813;
  assign n43815 = ~n43790 & ~n43814;
  assign n43816 = pi525 & ~n43815;
  assign n43817 = ~n43810 & ~n43816;
  assign n43818 = ~pi547 & n43817;
  assign n43819 = pi547 & n43742;
  assign n43820 = ~pi247 & ~n43819;
  assign n43821 = ~n43818 & n43820;
  assign n43822 = ~n43793 & ~n43821;
  assign n43823 = ~pi527 & ~n43822;
  assign n43824 = ~pi547 & n43742;
  assign n43825 = pi547 & n43817;
  assign n43826 = pi247 & ~n43824;
  assign n43827 = ~n43825 & n43826;
  assign n43828 = ~n43795 & ~n43827;
  assign n43829 = pi527 & ~n43828;
  assign n43830 = ~n43823 & ~n43829;
  assign n43831 = ~pi238 & n43830;
  assign n43832 = ~pi529 & ~n43831;
  assign n43833 = ~pi491 & ~n43799;
  assign n43834 = ~n43832 & n43833;
  assign n43835 = ~pi238 & n43746;
  assign n43836 = pi238 & n43796;
  assign n43837 = ~pi529 & ~n43835;
  assign n43838 = ~n43836 & n43837;
  assign n43839 = pi238 & n43830;
  assign n43840 = pi529 & ~n43839;
  assign n43841 = pi491 & ~n43838;
  assign n43842 = ~n43840 & n43841;
  assign n43843 = ~n43834 & ~n43842;
  assign n43844 = pi233 & ~n43843;
  assign n43845 = ~pi237 & ~n43698;
  assign n43846 = ~n43844 & n43845;
  assign po750 = ~n43592 & ~n43846;
  assign n43848 = ~pi806 & n42590;
  assign n43849 = ~pi332 & ~pi806;
  assign n43850 = pi990 & n43849;
  assign n43851 = pi600 & n43850;
  assign n43852 = ~pi332 & pi594;
  assign n43853 = ~n43851 & ~n43852;
  assign po751 = ~n43848 & ~n43853;
  assign n43855 = pi605 & ~pi806;
  assign n43856 = n42580 & n43855;
  assign n43857 = ~pi595 & ~n43856;
  assign n43858 = pi595 & n43856;
  assign n43859 = ~pi332 & ~n43857;
  assign po752 = ~n43858 & n43859;
  assign n43861 = ~pi332 & pi596;
  assign n43862 = pi595 & n42579;
  assign n43863 = n43850 & n43862;
  assign n43864 = ~n43861 & ~n43863;
  assign n43865 = pi596 & n43863;
  assign po753 = ~n43864 & ~n43865;
  assign n43867 = ~pi597 & ~n43848;
  assign n43868 = pi597 & n43848;
  assign n43869 = ~pi332 & ~n43867;
  assign po754 = ~n43868 & n43869;
  assign n43871 = ~pi882 & ~po1038;
  assign n43872 = pi947 & n43871;
  assign n43873 = pi598 & ~n43872;
  assign n43874 = pi740 & pi780;
  assign n43875 = n6161 & n43874;
  assign po755 = n43873 | n43875;
  assign n43877 = ~pi332 & pi599;
  assign n43878 = ~n43865 & ~n43877;
  assign n43879 = pi599 & n43865;
  assign po756 = ~n43878 & ~n43879;
  assign n43881 = ~pi332 & pi600;
  assign n43882 = ~n43850 & ~n43881;
  assign po757 = ~n43851 & ~n43882;
  assign n43884 = ~pi806 & ~pi989;
  assign n43885 = ~pi601 & pi806;
  assign n43886 = ~pi332 & ~n43884;
  assign po758 = ~n43885 & n43886;
  assign n43888 = ~pi230 & pi602;
  assign n43889 = pi715 & pi1160;
  assign n43890 = ~pi715 & ~pi1160;
  assign n43891 = pi790 & ~n43889;
  assign n43892 = ~n43890 & n43891;
  assign n43893 = pi230 & n15725;
  assign n43894 = ~n15765 & n43893;
  assign n43895 = ~n17581 & ~n17768;
  assign n43896 = ~n43892 & n43895;
  assign n43897 = n43894 & n43896;
  assign n43898 = n17586 & n43897;
  assign po759 = n43888 | n43898;
  assign n43900 = pi871 & pi966;
  assign n43901 = pi872 & pi966;
  assign n43902 = pi832 & ~pi1100;
  assign n43903 = ~pi980 & pi1038;
  assign n43904 = pi1060 & n43903;
  assign n43905 = pi952 & ~pi1061;
  assign n43906 = n43904 & n43905;
  assign n43907 = n43902 & n43906;
  assign po897 = pi832 & n43906;
  assign n43909 = ~pi603 & ~po897;
  assign n43910 = ~pi966 & ~n43907;
  assign n43911 = ~n43909 & n43910;
  assign n43912 = ~n43900 & ~n43901;
  assign po760 = n43911 | ~n43912;
  assign n43914 = pi823 & n16108;
  assign n43915 = ~pi779 & n43914;
  assign n43916 = ~pi299 & pi983;
  assign n43917 = pi907 & n43916;
  assign n43918 = pi604 & ~n43917;
  assign n43919 = ~n43914 & n43918;
  assign po761 = n43915 | n43919;
  assign n43921 = ~pi605 & ~n43849;
  assign n43922 = ~pi332 & ~n43855;
  assign po762 = ~n43921 & n43922;
  assign n43924 = pi606 & ~po897;
  assign n43925 = pi1104 & po897;
  assign n43926 = ~n43924 & ~n43925;
  assign n43927 = ~pi966 & ~n43926;
  assign n43928 = pi837 & pi966;
  assign po763 = n43927 | n43928;
  assign n43930 = ~pi607 & ~po897;
  assign n43931 = ~pi1107 & po897;
  assign n43932 = ~pi966 & ~n43930;
  assign po764 = ~n43931 & n43932;
  assign n43934 = ~pi608 & ~po897;
  assign n43935 = ~pi1116 & po897;
  assign n43936 = ~pi966 & ~n43934;
  assign po765 = ~n43935 & n43936;
  assign n43938 = ~pi609 & ~po897;
  assign n43939 = ~pi1118 & po897;
  assign n43940 = ~pi966 & ~n43938;
  assign po766 = ~n43939 & n43940;
  assign n43942 = ~pi610 & ~po897;
  assign n43943 = ~pi1113 & po897;
  assign n43944 = ~pi966 & ~n43942;
  assign po767 = ~n43943 & n43944;
  assign n43946 = ~pi611 & ~po897;
  assign n43947 = ~pi1114 & po897;
  assign n43948 = ~pi966 & ~n43946;
  assign po768 = ~n43947 & n43948;
  assign n43950 = ~pi612 & ~po897;
  assign n43951 = ~pi1111 & po897;
  assign n43952 = ~pi966 & ~n43950;
  assign po769 = ~n43951 & n43952;
  assign n43954 = ~pi613 & ~po897;
  assign n43955 = ~pi1115 & po897;
  assign n43956 = ~pi966 & ~n43954;
  assign po770 = ~n43955 & n43956;
  assign n43958 = ~pi614 & ~po897;
  assign n43959 = ~pi1102 & po897;
  assign n43960 = ~pi966 & ~n43958;
  assign n43961 = ~n43959 & n43960;
  assign po771 = n43900 | n43961;
  assign n43963 = pi907 & n43871;
  assign n43964 = ~pi615 & ~n43963;
  assign n43965 = pi779 & pi797;
  assign n43966 = n6164 & n43965;
  assign po772 = n43964 | n43966;
  assign n43968 = ~pi616 & ~po897;
  assign n43969 = ~pi1101 & po897;
  assign n43970 = ~pi966 & ~n43968;
  assign n43971 = ~n43969 & n43970;
  assign po773 = n43901 | n43971;
  assign n43973 = pi617 & ~po897;
  assign n43974 = pi1105 & po897;
  assign n43975 = ~n43973 & ~n43974;
  assign n43976 = ~pi966 & ~n43975;
  assign n43977 = pi850 & pi966;
  assign po774 = n43976 | n43977;
  assign n43979 = ~pi618 & ~po897;
  assign n43980 = ~pi1117 & po897;
  assign n43981 = ~pi966 & ~n43979;
  assign po775 = ~n43980 & n43981;
  assign n43983 = ~pi619 & ~po897;
  assign n43984 = ~pi1122 & po897;
  assign n43985 = ~pi966 & ~n43983;
  assign po776 = ~n43984 & n43985;
  assign n43987 = ~pi620 & ~po897;
  assign n43988 = ~pi1112 & po897;
  assign n43989 = ~pi966 & ~n43987;
  assign po777 = ~n43988 & n43989;
  assign n43991 = ~pi621 & ~po897;
  assign n43992 = ~pi1108 & po897;
  assign n43993 = ~pi966 & ~n43991;
  assign po778 = ~n43992 & n43993;
  assign n43995 = ~pi622 & ~po897;
  assign n43996 = ~pi1109 & po897;
  assign n43997 = ~pi966 & ~n43995;
  assign po779 = ~n43996 & n43997;
  assign n43999 = ~pi623 & ~po897;
  assign n44000 = ~pi1106 & po897;
  assign n44001 = ~pi966 & ~n43999;
  assign po780 = ~n44000 & n44001;
  assign n44003 = pi831 & n16452;
  assign n44004 = ~pi780 & n44003;
  assign n44005 = pi947 & n43916;
  assign n44006 = pi624 & ~n44005;
  assign n44007 = ~n44003 & n44006;
  assign po781 = n44004 | n44007;
  assign n44009 = pi832 & ~pi973;
  assign n44010 = ~pi1054 & pi1066;
  assign n44011 = pi1088 & n44010;
  assign n44012 = n44009 & n44011;
  assign po954 = ~pi953 & n44012;
  assign n44014 = ~pi625 & ~po954;
  assign n44015 = ~pi1116 & po954;
  assign n44016 = ~pi962 & ~n44014;
  assign po782 = ~n44015 & n44016;
  assign n44018 = ~pi626 & ~po897;
  assign n44019 = ~pi1121 & po897;
  assign n44020 = ~pi966 & ~n44018;
  assign po783 = ~n44019 & n44020;
  assign n44022 = ~pi627 & ~po954;
  assign n44023 = ~pi1117 & po954;
  assign n44024 = ~pi962 & ~n44022;
  assign po784 = ~n44023 & n44024;
  assign n44026 = ~pi628 & ~po954;
  assign n44027 = ~pi1119 & po954;
  assign n44028 = ~pi962 & ~n44026;
  assign po785 = ~n44027 & n44028;
  assign n44030 = ~pi629 & ~po897;
  assign n44031 = ~pi1119 & po897;
  assign n44032 = ~pi966 & ~n44030;
  assign po786 = ~n44031 & n44032;
  assign n44034 = ~pi630 & ~po897;
  assign n44035 = ~pi1120 & po897;
  assign n44036 = ~pi966 & ~n44034;
  assign po787 = ~n44035 & n44036;
  assign n44038 = ~pi1113 & po954;
  assign n44039 = pi631 & ~po954;
  assign n44040 = ~pi962 & ~n44038;
  assign po788 = ~n44039 & n44040;
  assign n44042 = ~pi1115 & po954;
  assign n44043 = pi632 & ~po954;
  assign n44044 = ~pi962 & ~n44042;
  assign po789 = ~n44043 & n44044;
  assign n44046 = ~pi633 & ~po897;
  assign n44047 = ~pi1110 & po897;
  assign n44048 = ~pi966 & ~n44046;
  assign po790 = ~n44047 & n44048;
  assign n44050 = ~pi634 & ~po954;
  assign n44051 = ~pi1110 & po954;
  assign n44052 = ~pi962 & ~n44050;
  assign po791 = ~n44051 & n44052;
  assign n44054 = ~pi1112 & po954;
  assign n44055 = pi635 & ~po954;
  assign n44056 = ~pi962 & ~n44054;
  assign po792 = ~n44055 & n44056;
  assign n44058 = ~pi636 & ~po897;
  assign n44059 = ~pi1127 & po897;
  assign n44060 = ~pi966 & ~n44058;
  assign po793 = ~n44059 & n44060;
  assign n44062 = ~pi637 & ~po954;
  assign n44063 = ~pi1105 & po954;
  assign n44064 = ~pi962 & ~n44062;
  assign po794 = ~n44063 & n44064;
  assign n44066 = ~pi638 & ~po954;
  assign n44067 = ~pi1107 & po954;
  assign n44068 = ~pi962 & ~n44066;
  assign po795 = ~n44067 & n44068;
  assign n44070 = ~pi639 & ~po954;
  assign n44071 = ~pi1109 & po954;
  assign n44072 = ~pi962 & ~n44070;
  assign po796 = ~n44071 & n44072;
  assign n44074 = ~pi640 & ~po897;
  assign n44075 = ~pi1128 & po897;
  assign n44076 = ~pi966 & ~n44074;
  assign po797 = ~n44075 & n44076;
  assign n44078 = ~pi641 & ~po954;
  assign n44079 = ~pi1121 & po954;
  assign n44080 = ~pi962 & ~n44078;
  assign po798 = ~n44079 & n44080;
  assign n44082 = ~pi642 & ~po897;
  assign n44083 = ~pi1103 & po897;
  assign n44084 = ~pi966 & ~n44082;
  assign po799 = ~n44083 & n44084;
  assign n44086 = ~pi643 & ~po954;
  assign n44087 = ~pi1104 & po954;
  assign n44088 = ~pi962 & ~n44086;
  assign po800 = ~n44087 & n44088;
  assign n44090 = ~pi644 & ~po897;
  assign n44091 = ~pi1123 & po897;
  assign n44092 = ~pi966 & ~n44090;
  assign po801 = ~n44091 & n44092;
  assign n44094 = ~pi645 & ~po897;
  assign n44095 = ~pi1125 & po897;
  assign n44096 = ~pi966 & ~n44094;
  assign po802 = ~n44095 & n44096;
  assign n44098 = ~pi1114 & po954;
  assign n44099 = pi646 & ~po954;
  assign n44100 = ~pi962 & ~n44098;
  assign po803 = ~n44099 & n44100;
  assign n44102 = ~pi647 & ~po954;
  assign n44103 = ~pi1120 & po954;
  assign n44104 = ~pi962 & ~n44102;
  assign po804 = ~n44103 & n44104;
  assign n44106 = ~pi648 & ~po954;
  assign n44107 = ~pi1122 & po954;
  assign n44108 = ~pi962 & ~n44106;
  assign po805 = ~n44107 & n44108;
  assign n44110 = ~pi1126 & po954;
  assign n44111 = pi649 & ~po954;
  assign n44112 = ~pi962 & ~n44110;
  assign po806 = ~n44111 & n44112;
  assign n44114 = ~pi1127 & po954;
  assign n44115 = pi650 & ~po954;
  assign n44116 = ~pi962 & ~n44114;
  assign po807 = ~n44115 & n44116;
  assign n44118 = ~pi651 & ~po897;
  assign n44119 = ~pi1130 & po897;
  assign n44120 = ~pi966 & ~n44118;
  assign po808 = ~n44119 & n44120;
  assign n44122 = ~pi652 & ~po897;
  assign n44123 = ~pi1131 & po897;
  assign n44124 = ~pi966 & ~n44122;
  assign po809 = ~n44123 & n44124;
  assign n44126 = ~pi653 & ~po897;
  assign n44127 = ~pi1129 & po897;
  assign n44128 = ~pi966 & ~n44126;
  assign po810 = ~n44127 & n44128;
  assign n44130 = ~pi1130 & po954;
  assign n44131 = pi654 & ~po954;
  assign n44132 = ~pi962 & ~n44130;
  assign po811 = ~n44131 & n44132;
  assign n44134 = ~pi1124 & po954;
  assign n44135 = pi655 & ~po954;
  assign n44136 = ~pi962 & ~n44134;
  assign po812 = ~n44135 & n44136;
  assign n44138 = ~pi656 & ~po897;
  assign n44139 = ~pi1126 & po897;
  assign n44140 = ~pi966 & ~n44138;
  assign po813 = ~n44139 & n44140;
  assign n44142 = ~pi1131 & po954;
  assign n44143 = pi657 & ~po954;
  assign n44144 = ~pi962 & ~n44142;
  assign po814 = ~n44143 & n44144;
  assign n44146 = ~pi658 & ~po897;
  assign n44147 = ~pi1124 & po897;
  assign n44148 = ~pi966 & ~n44146;
  assign po815 = ~n44147 & n44148;
  assign n44150 = pi266 & pi992;
  assign n44151 = ~pi280 & n44150;
  assign n44152 = ~pi269 & n44151;
  assign n44153 = ~pi281 & n44152;
  assign n44154 = ~pi270 & ~pi277;
  assign n44155 = ~pi282 & n44154;
  assign n44156 = n44153 & n44155;
  assign n44157 = ~pi264 & n44156;
  assign n44158 = ~pi265 & n44157;
  assign po959 = ~pi274 & n44158;
  assign n44160 = pi274 & ~n44158;
  assign po816 = ~po959 & ~n44160;
  assign n44162 = ~pi660 & ~po954;
  assign n44163 = ~pi1118 & po954;
  assign n44164 = ~pi962 & ~n44162;
  assign po817 = ~n44163 & n44164;
  assign n44166 = ~pi661 & ~po954;
  assign n44167 = ~pi1101 & po954;
  assign n44168 = ~pi962 & ~n44166;
  assign po818 = ~n44167 & n44168;
  assign n44170 = ~pi662 & ~po954;
  assign n44171 = ~pi1102 & po954;
  assign n44172 = ~pi962 & ~n44170;
  assign po819 = ~n44171 & n44172;
  assign n44174 = pi464 & n7580;
  assign n44175 = pi588 & ~n44174;
  assign n44176 = ~pi223 & ~pi224;
  assign n44177 = ~pi591 & ~pi592;
  assign n44178 = pi590 & n44177;
  assign n44179 = pi323 & n44178;
  assign n44180 = ~pi591 & pi592;
  assign n44181 = pi365 & n44180;
  assign n44182 = pi334 & pi591;
  assign n44183 = ~pi592 & n44182;
  assign n44184 = ~n44181 & ~n44183;
  assign n44185 = ~pi590 & ~n44184;
  assign n44186 = ~pi588 & ~n44179;
  assign n44187 = ~n44185 & n44186;
  assign n44188 = ~n44175 & n44176;
  assign n44189 = ~n44187 & n44188;
  assign n44190 = ~pi199 & ~pi257;
  assign n44191 = pi199 & ~pi1065;
  assign n44192 = ~n44176 & ~n44190;
  assign n44193 = ~n44191 & n44192;
  assign n44194 = ~n44189 & ~n44193;
  assign n44195 = n7578 & ~n44194;
  assign n44196 = ~pi1137 & ~pi1138;
  assign n44197 = ~pi1134 & n44196;
  assign n44198 = ~pi784 & ~pi1136;
  assign n44199 = ~pi634 & pi1136;
  assign n44200 = pi1135 & ~n44198;
  assign n44201 = ~n44199 & n44200;
  assign n44202 = ~pi815 & ~pi1136;
  assign n44203 = ~pi633 & pi1136;
  assign n44204 = ~pi1135 & ~n44202;
  assign n44205 = ~n44203 & n44204;
  assign n44206 = ~n44201 & ~n44205;
  assign n44207 = n44197 & ~n44206;
  assign n44208 = ~pi700 & pi1135;
  assign n44209 = pi1135 & ~pi1136;
  assign n44210 = pi1134 & n44196;
  assign n44211 = ~n44209 & n44210;
  assign n44212 = ~pi855 & ~pi1136;
  assign n44213 = pi1135 & n44196;
  assign n44214 = pi1136 & ~n44213;
  assign n44215 = ~pi766 & n44214;
  assign n44216 = ~n44208 & ~n44212;
  assign n44217 = n44211 & n44216;
  assign n44218 = ~n44215 & n44217;
  assign n44219 = ~n44207 & ~n44218;
  assign n44220 = ~n7578 & ~n44219;
  assign po820 = n44195 | n44220;
  assign n44222 = pi429 & n7580;
  assign n44223 = pi588 & ~n44222;
  assign n44224 = ~pi590 & pi591;
  assign n44225 = pi404 & n44224;
  assign n44226 = ~pi590 & pi592;
  assign n44227 = ~pi588 & ~n44226;
  assign n44228 = ~n44225 & n44227;
  assign n44229 = pi380 & ~pi591;
  assign n44230 = pi592 & ~n44229;
  assign n44231 = ~n44228 & ~n44230;
  assign n44232 = pi355 & n44178;
  assign n44233 = ~n44231 & ~n44232;
  assign n44234 = n44176 & ~n44223;
  assign n44235 = ~n44233 & n44234;
  assign n44236 = ~pi199 & ~pi292;
  assign n44237 = pi199 & ~pi1084;
  assign n44238 = ~n44176 & ~n44236;
  assign n44239 = ~n44237 & n44238;
  assign n44240 = ~n44235 & ~n44239;
  assign n44241 = n7578 & ~n44240;
  assign n44242 = ~pi1135 & ~pi1136;
  assign n44243 = pi872 & n44242;
  assign n44244 = ~pi772 & ~pi1135;
  assign n44245 = ~pi727 & pi1135;
  assign n44246 = pi1136 & ~n44244;
  assign n44247 = ~n44245 & n44246;
  assign n44248 = pi1134 & ~n44243;
  assign n44249 = ~n44247 & n44248;
  assign n44250 = ~n7578 & n44196;
  assign n44251 = pi614 & ~pi1135;
  assign n44252 = pi662 & pi1135;
  assign n44253 = pi1136 & ~n44251;
  assign n44254 = ~n44252 & n44253;
  assign n44255 = pi811 & ~pi1135;
  assign n44256 = pi785 & pi1135;
  assign n44257 = ~pi1136 & ~n44255;
  assign n44258 = ~n44256 & n44257;
  assign n44259 = ~n44254 & ~n44258;
  assign n44260 = ~pi1134 & ~n44259;
  assign n44261 = ~n44249 & n44250;
  assign n44262 = ~n44260 & n44261;
  assign po821 = n44241 | n44262;
  assign n44264 = ~pi665 & ~po954;
  assign n44265 = ~pi1108 & po954;
  assign n44266 = ~pi962 & ~n44264;
  assign po822 = ~n44265 & n44266;
  assign n44268 = ~pi607 & ~pi1135;
  assign n44269 = ~pi638 & pi1135;
  assign n44270 = pi1136 & ~n44268;
  assign n44271 = ~n44269 & n44270;
  assign n44272 = ~pi790 & pi1135;
  assign n44273 = pi799 & ~pi1135;
  assign n44274 = ~pi1136 & ~n44272;
  assign n44275 = ~n44273 & n44274;
  assign n44276 = ~n44271 & ~n44275;
  assign n44277 = n44197 & ~n44276;
  assign n44278 = ~pi691 & pi1135;
  assign n44279 = ~pi764 & n44214;
  assign n44280 = ~pi873 & ~pi1136;
  assign n44281 = ~n44278 & ~n44280;
  assign n44282 = n44211 & n44281;
  assign n44283 = ~n44279 & n44282;
  assign n44284 = ~n44277 & ~n44283;
  assign n44285 = ~n7578 & ~n44284;
  assign n44286 = ~pi199 & ~pi297;
  assign n44287 = pi199 & ~pi1044;
  assign n44288 = ~n44176 & ~n44286;
  assign n44289 = ~n44287 & n44288;
  assign n44290 = pi443 & n7580;
  assign n44291 = pi588 & ~n44290;
  assign n44292 = pi456 & n44224;
  assign n44293 = n44227 & ~n44292;
  assign n44294 = pi337 & ~pi591;
  assign n44295 = pi592 & ~n44294;
  assign n44296 = ~n44293 & ~n44295;
  assign n44297 = pi441 & n44178;
  assign n44298 = ~n44296 & ~n44297;
  assign n44299 = n44176 & ~n44291;
  assign n44300 = ~n44298 & n44299;
  assign n44301 = ~n44289 & ~n44300;
  assign n44302 = n7578 & ~n44301;
  assign po823 = n44285 | n44302;
  assign n44304 = pi444 & n7580;
  assign n44305 = pi588 & ~n44304;
  assign n44306 = pi319 & n44224;
  assign n44307 = n44227 & ~n44306;
  assign n44308 = pi338 & ~pi591;
  assign n44309 = pi592 & ~n44308;
  assign n44310 = ~n44307 & ~n44309;
  assign n44311 = pi458 & n44178;
  assign n44312 = ~n44310 & ~n44311;
  assign n44313 = n44176 & ~n44305;
  assign n44314 = ~n44312 & n44313;
  assign n44315 = ~pi199 & ~pi294;
  assign n44316 = pi199 & ~pi1072;
  assign n44317 = ~n44176 & ~n44315;
  assign n44318 = ~n44316 & n44317;
  assign n44319 = ~n44314 & ~n44318;
  assign n44320 = n7578 & ~n44319;
  assign n44321 = pi871 & n44242;
  assign n44322 = ~pi763 & ~pi1135;
  assign n44323 = ~pi699 & pi1135;
  assign n44324 = pi1136 & ~n44322;
  assign n44325 = ~n44323 & n44324;
  assign n44326 = pi1134 & ~n44321;
  assign n44327 = ~n44325 & n44326;
  assign n44328 = pi792 & ~pi1136;
  assign n44329 = pi681 & pi1136;
  assign n44330 = pi1135 & ~n44328;
  assign n44331 = ~n44329 & n44330;
  assign n44332 = ~pi809 & ~pi1136;
  assign n44333 = pi642 & pi1136;
  assign n44334 = ~pi1135 & ~n44332;
  assign n44335 = ~n44333 & n44334;
  assign n44336 = ~n44331 & ~n44335;
  assign n44337 = ~pi1134 & ~n44336;
  assign n44338 = n44250 & ~n44327;
  assign n44339 = ~n44337 & n44338;
  assign po824 = n44320 | n44339;
  assign n44341 = ~pi603 & ~pi1135;
  assign n44342 = ~pi680 & pi1135;
  assign n44343 = pi1136 & ~n44341;
  assign n44344 = ~n44342 & n44343;
  assign n44345 = ~pi981 & ~pi1135;
  assign n44346 = ~pi778 & pi1135;
  assign n44347 = ~pi1136 & ~n44345;
  assign n44348 = ~n44346 & n44347;
  assign n44349 = ~n44344 & ~n44348;
  assign n44350 = n44197 & ~n44349;
  assign n44351 = ~pi696 & pi1135;
  assign n44352 = ~pi759 & n44214;
  assign n44353 = ~pi837 & ~pi1136;
  assign n44354 = ~n44351 & ~n44353;
  assign n44355 = n44211 & n44354;
  assign n44356 = ~n44352 & n44355;
  assign n44357 = ~n44350 & ~n44356;
  assign n44358 = ~n7578 & ~n44357;
  assign n44359 = ~pi199 & ~pi291;
  assign n44360 = pi199 & ~pi1049;
  assign n44361 = ~n44176 & ~n44359;
  assign n44362 = ~n44360 & n44361;
  assign n44363 = pi414 & n7580;
  assign n44364 = pi588 & ~n44363;
  assign n44365 = pi390 & n44224;
  assign n44366 = n44227 & ~n44365;
  assign n44367 = pi363 & ~pi591;
  assign n44368 = pi592 & ~n44367;
  assign n44369 = ~n44366 & ~n44368;
  assign n44370 = pi342 & n44178;
  assign n44371 = ~n44369 & ~n44370;
  assign n44372 = n44176 & ~n44364;
  assign n44373 = ~n44371 & n44372;
  assign n44374 = ~n44362 & ~n44373;
  assign n44375 = n7578 & ~n44374;
  assign po825 = n44358 | n44375;
  assign n44377 = ~pi1125 & po954;
  assign n44378 = pi669 & ~po954;
  assign n44379 = ~pi962 & ~n44377;
  assign po826 = ~n44378 & n44379;
  assign n44381 = pi695 & pi1135;
  assign n44382 = pi1136 & n44196;
  assign n44383 = ~pi612 & ~pi1135;
  assign n44384 = ~pi1134 & ~n44381;
  assign n44385 = ~n44383 & n44384;
  assign n44386 = n44382 & n44385;
  assign n44387 = pi723 & pi1135;
  assign n44388 = ~pi852 & ~pi1136;
  assign n44389 = pi745 & n44214;
  assign n44390 = ~n44387 & ~n44388;
  assign n44391 = n44211 & n44390;
  assign n44392 = ~n44389 & n44391;
  assign n44393 = ~n44386 & ~n44392;
  assign n44394 = ~n7578 & ~n44393;
  assign n44395 = ~pi199 & ~pi258;
  assign n44396 = pi199 & ~pi1062;
  assign n44397 = ~n44176 & ~n44395;
  assign n44398 = ~n44396 & n44397;
  assign n44399 = pi415 & n7580;
  assign n44400 = pi588 & ~n44399;
  assign n44401 = pi343 & n44178;
  assign n44402 = pi364 & n44180;
  assign n44403 = pi391 & pi591;
  assign n44404 = ~pi592 & n44403;
  assign n44405 = ~n44402 & ~n44404;
  assign n44406 = ~pi590 & ~n44405;
  assign n44407 = ~pi588 & ~n44401;
  assign n44408 = ~n44406 & n44407;
  assign n44409 = n44176 & ~n44400;
  assign n44410 = ~n44408 & n44409;
  assign n44411 = ~n44398 & ~n44410;
  assign n44412 = n7578 & ~n44411;
  assign po827 = n44394 | n44412;
  assign n44414 = pi646 & pi1135;
  assign n44415 = ~pi611 & ~pi1135;
  assign n44416 = ~pi1134 & ~n44414;
  assign n44417 = ~n44415 & n44416;
  assign n44418 = n44382 & n44417;
  assign n44419 = pi724 & pi1135;
  assign n44420 = ~pi865 & ~pi1136;
  assign n44421 = pi741 & n44214;
  assign n44422 = ~n44419 & ~n44420;
  assign n44423 = n44211 & n44422;
  assign n44424 = ~n44421 & n44423;
  assign n44425 = ~n44418 & ~n44424;
  assign n44426 = ~n7578 & ~n44425;
  assign n44427 = ~pi199 & ~pi261;
  assign n44428 = pi199 & ~pi1040;
  assign n44429 = ~n44176 & ~n44427;
  assign n44430 = ~n44428 & n44429;
  assign n44431 = pi453 & n7580;
  assign n44432 = pi588 & ~n44431;
  assign n44433 = pi327 & n44178;
  assign n44434 = pi447 & n44180;
  assign n44435 = pi333 & pi591;
  assign n44436 = ~pi592 & n44435;
  assign n44437 = ~n44434 & ~n44436;
  assign n44438 = ~pi590 & ~n44437;
  assign n44439 = ~pi588 & ~n44433;
  assign n44440 = ~n44438 & n44439;
  assign n44441 = n44176 & ~n44432;
  assign n44442 = ~n44440 & n44441;
  assign n44443 = ~n44430 & ~n44442;
  assign n44444 = n7578 & ~n44443;
  assign po828 = n44426 | n44444;
  assign n44446 = ~pi616 & ~pi1135;
  assign n44447 = ~pi661 & pi1135;
  assign n44448 = pi1136 & ~n44446;
  assign n44449 = ~n44447 & n44448;
  assign n44450 = ~pi808 & ~pi1135;
  assign n44451 = ~pi781 & pi1135;
  assign n44452 = ~pi1136 & ~n44450;
  assign n44453 = ~n44451 & n44452;
  assign n44454 = ~n44449 & ~n44453;
  assign n44455 = n44197 & ~n44454;
  assign n44456 = ~pi736 & pi1135;
  assign n44457 = ~pi758 & n44214;
  assign n44458 = ~pi850 & ~pi1136;
  assign n44459 = ~n44456 & ~n44458;
  assign n44460 = n44211 & n44459;
  assign n44461 = ~n44457 & n44460;
  assign n44462 = ~n44455 & ~n44461;
  assign n44463 = ~n7578 & ~n44462;
  assign n44464 = ~pi199 & ~pi290;
  assign n44465 = pi199 & ~pi1048;
  assign n44466 = ~n44176 & ~n44464;
  assign n44467 = ~n44465 & n44466;
  assign n44468 = pi422 & n7580;
  assign n44469 = pi588 & ~n44468;
  assign n44470 = pi397 & n44224;
  assign n44471 = n44227 & ~n44470;
  assign n44472 = pi372 & ~pi591;
  assign n44473 = pi592 & ~n44472;
  assign n44474 = ~n44471 & ~n44473;
  assign n44475 = pi320 & n44178;
  assign n44476 = ~n44474 & ~n44475;
  assign n44477 = n44176 & ~n44469;
  assign n44478 = ~n44476 & n44477;
  assign n44479 = ~n44467 & ~n44478;
  assign n44480 = n7578 & ~n44479;
  assign po829 = n44463 | n44480;
  assign n44482 = ~pi617 & ~pi1135;
  assign n44483 = ~pi637 & pi1135;
  assign n44484 = pi1136 & ~n44482;
  assign n44485 = ~n44483 & n44484;
  assign n44486 = ~pi788 & pi1135;
  assign n44487 = pi814 & ~pi1135;
  assign n44488 = ~pi1136 & ~n44486;
  assign n44489 = ~n44487 & n44488;
  assign n44490 = ~n44485 & ~n44489;
  assign n44491 = n44197 & ~n44490;
  assign n44492 = ~pi706 & pi1135;
  assign n44493 = ~pi749 & n44214;
  assign n44494 = ~pi866 & ~pi1136;
  assign n44495 = ~n44492 & ~n44494;
  assign n44496 = n44211 & n44495;
  assign n44497 = ~n44493 & n44496;
  assign n44498 = ~n44491 & ~n44497;
  assign n44499 = ~n7578 & ~n44498;
  assign n44500 = ~pi199 & ~pi295;
  assign n44501 = pi199 & ~pi1053;
  assign n44502 = ~n44176 & ~n44500;
  assign n44503 = ~n44501 & n44502;
  assign n44504 = pi435 & n7580;
  assign n44505 = pi588 & ~n44504;
  assign n44506 = pi411 & n44224;
  assign n44507 = n44227 & ~n44506;
  assign n44508 = pi387 & ~pi591;
  assign n44509 = pi592 & ~n44508;
  assign n44510 = ~n44507 & ~n44509;
  assign n44511 = pi452 & n44178;
  assign n44512 = ~n44510 & ~n44511;
  assign n44513 = n44176 & ~n44505;
  assign n44514 = ~n44512 & n44513;
  assign n44515 = ~n44503 & ~n44514;
  assign n44516 = n7578 & ~n44515;
  assign po830 = n44499 | n44516;
  assign n44518 = pi437 & n7580;
  assign n44519 = pi588 & ~n44518;
  assign n44520 = pi362 & n44178;
  assign n44521 = pi336 & n44180;
  assign n44522 = pi463 & pi591;
  assign n44523 = ~pi592 & n44522;
  assign n44524 = ~n44521 & ~n44523;
  assign n44525 = ~pi590 & ~n44524;
  assign n44526 = ~pi588 & ~n44520;
  assign n44527 = ~n44525 & n44526;
  assign n44528 = n44176 & ~n44519;
  assign n44529 = ~n44527 & n44528;
  assign n44530 = ~pi199 & ~pi256;
  assign n44531 = pi199 & ~pi1070;
  assign n44532 = ~n44176 & ~n44530;
  assign n44533 = ~n44531 & n44532;
  assign n44534 = ~n44529 & ~n44533;
  assign n44535 = n7578 & ~n44534;
  assign n44536 = pi859 & n44242;
  assign n44537 = ~pi743 & ~pi1135;
  assign n44538 = ~pi735 & pi1135;
  assign n44539 = pi1136 & ~n44537;
  assign n44540 = ~n44538 & n44539;
  assign n44541 = pi1134 & ~n44536;
  assign n44542 = ~n44540 & n44541;
  assign n44543 = pi622 & ~pi1135;
  assign n44544 = pi639 & pi1135;
  assign n44545 = pi1136 & ~n44543;
  assign n44546 = ~n44544 & n44545;
  assign n44547 = pi804 & ~pi1135;
  assign n44548 = pi783 & pi1135;
  assign n44549 = ~pi1136 & ~n44547;
  assign n44550 = ~n44548 & n44549;
  assign n44551 = ~n44546 & ~n44550;
  assign n44552 = ~pi1134 & ~n44551;
  assign n44553 = n44250 & ~n44542;
  assign n44554 = ~n44552 & n44553;
  assign po831 = n44535 | n44554;
  assign n44556 = pi876 & n44242;
  assign n44557 = ~pi748 & ~pi1135;
  assign n44558 = ~pi730 & pi1135;
  assign n44559 = pi1136 & ~n44557;
  assign n44560 = ~n44558 & n44559;
  assign n44561 = ~n44556 & ~n44560;
  assign n44562 = n44210 & ~n44561;
  assign n44563 = ~pi623 & n44214;
  assign n44564 = ~pi803 & ~pi1135;
  assign n44565 = pi789 & n44209;
  assign n44566 = ~pi710 & pi1135;
  assign n44567 = pi1136 & ~n44566;
  assign n44568 = ~n44564 & ~n44565;
  assign n44569 = ~n44567 & n44568;
  assign n44570 = n44197 & ~n44563;
  assign n44571 = ~n44569 & n44570;
  assign n44572 = ~n44562 & ~n44571;
  assign n44573 = ~n7578 & ~n44572;
  assign n44574 = ~pi199 & ~pi296;
  assign n44575 = pi199 & ~pi1037;
  assign n44576 = ~n44176 & ~n44574;
  assign n44577 = ~n44575 & n44576;
  assign n44578 = pi436 & n7580;
  assign n44579 = pi588 & ~n44578;
  assign n44580 = pi412 & n44224;
  assign n44581 = n44227 & ~n44580;
  assign n44582 = pi388 & ~pi591;
  assign n44583 = pi592 & ~n44582;
  assign n44584 = ~n44581 & ~n44583;
  assign n44585 = pi455 & n44178;
  assign n44586 = ~n44584 & ~n44585;
  assign n44587 = n44176 & ~n44579;
  assign n44588 = ~n44586 & n44587;
  assign n44589 = ~n44577 & ~n44588;
  assign n44590 = n7578 & ~n44589;
  assign po832 = n44573 | n44590;
  assign n44592 = ~pi606 & ~pi1135;
  assign n44593 = ~pi643 & pi1135;
  assign n44594 = pi1136 & ~n44592;
  assign n44595 = ~n44593 & n44594;
  assign n44596 = ~pi787 & pi1135;
  assign n44597 = pi812 & ~pi1135;
  assign n44598 = ~pi1136 & ~n44596;
  assign n44599 = ~n44597 & n44598;
  assign n44600 = ~n44595 & ~n44599;
  assign n44601 = n44197 & ~n44600;
  assign n44602 = ~pi729 & pi1135;
  assign n44603 = ~pi746 & n44214;
  assign n44604 = ~pi881 & ~pi1136;
  assign n44605 = ~n44602 & ~n44604;
  assign n44606 = n44211 & n44605;
  assign n44607 = ~n44603 & n44606;
  assign n44608 = ~n44601 & ~n44607;
  assign n44609 = ~n7578 & ~n44608;
  assign n44610 = ~pi199 & ~pi293;
  assign n44611 = pi199 & ~pi1059;
  assign n44612 = ~n44176 & ~n44610;
  assign n44613 = ~n44611 & n44612;
  assign n44614 = pi434 & n7580;
  assign n44615 = pi588 & ~n44614;
  assign n44616 = pi410 & n44224;
  assign n44617 = n44227 & ~n44616;
  assign n44618 = pi386 & ~pi591;
  assign n44619 = pi592 & ~n44618;
  assign n44620 = ~n44617 & ~n44619;
  assign n44621 = pi361 & n44178;
  assign n44622 = ~n44620 & ~n44621;
  assign n44623 = n44176 & ~n44615;
  assign n44624 = ~n44622 & n44623;
  assign n44625 = ~n44613 & ~n44624;
  assign n44626 = n7578 & ~n44625;
  assign po833 = n44609 | n44626;
  assign n44628 = pi635 & pi1135;
  assign n44629 = ~pi620 & ~pi1135;
  assign n44630 = ~pi1134 & ~n44628;
  assign n44631 = ~n44629 & n44630;
  assign n44632 = n44382 & n44631;
  assign n44633 = pi704 & pi1135;
  assign n44634 = ~pi870 & ~pi1136;
  assign n44635 = pi742 & n44214;
  assign n44636 = ~n44633 & ~n44634;
  assign n44637 = n44211 & n44636;
  assign n44638 = ~n44635 & n44637;
  assign n44639 = ~n44632 & ~n44638;
  assign n44640 = ~n7578 & ~n44639;
  assign n44641 = ~pi199 & ~pi259;
  assign n44642 = pi199 & ~pi1069;
  assign n44643 = ~n44176 & ~n44641;
  assign n44644 = ~n44642 & n44643;
  assign n44645 = pi416 & n7580;
  assign n44646 = pi588 & ~n44645;
  assign n44647 = pi344 & n44178;
  assign n44648 = pi366 & n44180;
  assign n44649 = pi335 & pi591;
  assign n44650 = ~pi592 & n44649;
  assign n44651 = ~n44648 & ~n44650;
  assign n44652 = ~pi590 & ~n44651;
  assign n44653 = ~pi588 & ~n44647;
  assign n44654 = ~n44652 & n44653;
  assign n44655 = n44176 & ~n44646;
  assign n44656 = ~n44654 & n44655;
  assign n44657 = ~n44644 & ~n44656;
  assign n44658 = n7578 & ~n44657;
  assign po834 = n44640 | n44658;
  assign n44660 = pi632 & pi1135;
  assign n44661 = ~pi613 & ~pi1135;
  assign n44662 = ~pi1134 & ~n44660;
  assign n44663 = ~n44661 & n44662;
  assign n44664 = n44382 & n44663;
  assign n44665 = pi688 & pi1135;
  assign n44666 = ~pi856 & ~pi1136;
  assign n44667 = pi760 & n44214;
  assign n44668 = ~n44665 & ~n44666;
  assign n44669 = n44211 & n44668;
  assign n44670 = ~n44667 & n44669;
  assign n44671 = ~n44664 & ~n44670;
  assign n44672 = ~n7578 & ~n44671;
  assign n44673 = ~pi199 & ~pi260;
  assign n44674 = pi199 & ~pi1067;
  assign n44675 = ~n44176 & ~n44673;
  assign n44676 = ~n44674 & n44675;
  assign n44677 = pi418 & n7580;
  assign n44678 = pi588 & ~n44677;
  assign n44679 = pi346 & n44178;
  assign n44680 = pi368 & n44180;
  assign n44681 = pi393 & pi591;
  assign n44682 = ~pi592 & n44681;
  assign n44683 = ~n44680 & ~n44682;
  assign n44684 = ~pi590 & ~n44683;
  assign n44685 = ~pi588 & ~n44679;
  assign n44686 = ~n44684 & n44685;
  assign n44687 = n44176 & ~n44678;
  assign n44688 = ~n44686 & n44687;
  assign n44689 = ~n44676 & ~n44688;
  assign n44690 = n7578 & ~n44689;
  assign po835 = n44672 | n44690;
  assign n44692 = pi438 & n7580;
  assign n44693 = pi588 & ~n44692;
  assign n44694 = pi450 & n44178;
  assign n44695 = pi389 & n44180;
  assign n44696 = pi413 & pi591;
  assign n44697 = ~pi592 & n44696;
  assign n44698 = ~n44695 & ~n44697;
  assign n44699 = ~pi590 & ~n44698;
  assign n44700 = ~pi588 & ~n44694;
  assign n44701 = ~n44699 & n44700;
  assign n44702 = n44176 & ~n44693;
  assign n44703 = ~n44701 & n44702;
  assign n44704 = ~pi199 & ~pi255;
  assign n44705 = pi199 & ~pi1036;
  assign n44706 = ~n44176 & ~n44704;
  assign n44707 = ~n44705 & n44706;
  assign n44708 = ~n44703 & ~n44707;
  assign n44709 = n7578 & ~n44708;
  assign n44710 = ~pi791 & ~pi1136;
  assign n44711 = ~pi665 & pi1136;
  assign n44712 = pi1135 & ~n44710;
  assign n44713 = ~n44711 & n44712;
  assign n44714 = ~pi810 & ~pi1136;
  assign n44715 = ~pi621 & pi1136;
  assign n44716 = ~pi1135 & ~n44714;
  assign n44717 = ~n44715 & n44716;
  assign n44718 = ~n44713 & ~n44717;
  assign n44719 = n44197 & ~n44718;
  assign n44720 = ~pi690 & pi1135;
  assign n44721 = ~pi874 & ~pi1136;
  assign n44722 = ~pi739 & n44214;
  assign n44723 = ~n44720 & ~n44721;
  assign n44724 = n44211 & n44723;
  assign n44725 = ~n44722 & n44724;
  assign n44726 = ~n44719 & ~n44725;
  assign n44727 = ~n7578 & ~n44726;
  assign po836 = n44709 | n44727;
  assign n44729 = ~pi680 & ~po954;
  assign n44730 = ~pi1100 & po954;
  assign n44731 = ~pi962 & ~n44729;
  assign po837 = ~n44730 & n44731;
  assign n44733 = ~pi681 & ~po954;
  assign n44734 = ~pi1103 & po954;
  assign n44735 = ~pi962 & ~n44733;
  assign po838 = ~n44734 & n44735;
  assign n44737 = pi631 & pi1135;
  assign n44738 = ~pi610 & ~pi1135;
  assign n44739 = ~pi1134 & ~n44737;
  assign n44740 = ~n44738 & n44739;
  assign n44741 = n44382 & n44740;
  assign n44742 = pi686 & pi1135;
  assign n44743 = ~pi848 & ~pi1136;
  assign n44744 = pi757 & n44214;
  assign n44745 = ~n44742 & ~n44743;
  assign n44746 = n44211 & n44745;
  assign n44747 = ~n44744 & n44746;
  assign n44748 = ~n44741 & ~n44747;
  assign n44749 = ~n7578 & ~n44748;
  assign n44750 = ~pi199 & ~pi251;
  assign n44751 = pi199 & ~pi1039;
  assign n44752 = ~n44176 & ~n44750;
  assign n44753 = ~n44751 & n44752;
  assign n44754 = pi417 & n7580;
  assign n44755 = pi588 & ~n44754;
  assign n44756 = pi345 & n44178;
  assign n44757 = pi367 & n44180;
  assign n44758 = pi392 & pi591;
  assign n44759 = ~pi592 & n44758;
  assign n44760 = ~n44757 & ~n44759;
  assign n44761 = ~pi590 & ~n44760;
  assign n44762 = ~pi588 & ~n44756;
  assign n44763 = ~n44761 & n44762;
  assign n44764 = n44176 & ~n44755;
  assign n44765 = ~n44763 & n44764;
  assign n44766 = ~n44753 & ~n44765;
  assign n44767 = n7578 & ~n44766;
  assign po839 = n44749 | n44767;
  assign po980 = pi953 & n44012;
  assign n44770 = ~pi1130 & po980;
  assign n44771 = pi684 & ~po980;
  assign n44772 = ~pi962 & ~n44770;
  assign po841 = ~n44771 & n44772;
  assign n44774 = pi590 & ~pi592;
  assign n44775 = pi357 & n44774;
  assign n44776 = pi382 & n44226;
  assign n44777 = ~n44775 & ~n44776;
  assign n44778 = ~pi591 & ~n44777;
  assign n44779 = pi406 & ~pi592;
  assign n44780 = n44224 & n44779;
  assign n44781 = ~n44778 & ~n44780;
  assign n44782 = ~pi588 & ~n44781;
  assign n44783 = pi588 & ~pi590;
  assign n44784 = pi430 & n44177;
  assign n44785 = n44783 & n44784;
  assign n44786 = ~n44782 & ~n44785;
  assign n44787 = n44176 & ~n44786;
  assign n44788 = pi199 & ~pi1076;
  assign n44789 = ~n44176 & ~n44788;
  assign n44790 = ~n40456 & n44789;
  assign n44791 = ~n44787 & ~n44790;
  assign n44792 = n7578 & ~n44791;
  assign n44793 = pi860 & n44242;
  assign n44794 = pi744 & ~pi1135;
  assign n44795 = pi728 & pi1135;
  assign n44796 = pi1136 & ~n44794;
  assign n44797 = ~n44795 & n44796;
  assign n44798 = ~n44793 & ~n44797;
  assign n44799 = n44210 & ~n44798;
  assign n44800 = pi1136 & ~n44196;
  assign n44801 = ~pi1134 & ~n44800;
  assign n44802 = ~pi652 & ~pi1135;
  assign n44803 = pi657 & pi1135;
  assign n44804 = pi1136 & ~n44802;
  assign n44805 = ~n44803 & n44804;
  assign n44806 = pi813 & n44196;
  assign n44807 = n44242 & n44806;
  assign n44808 = ~n44805 & ~n44807;
  assign n44809 = n44801 & ~n44808;
  assign n44810 = ~n44799 & ~n44809;
  assign n44811 = ~n7578 & ~n44810;
  assign po842 = n44792 | n44811;
  assign n44813 = ~pi1113 & po980;
  assign n44814 = pi686 & ~po980;
  assign n44815 = ~pi962 & ~n44813;
  assign po843 = ~n44814 & n44815;
  assign n44817 = ~pi687 & ~po980;
  assign n44818 = ~pi1127 & po980;
  assign n44819 = ~pi962 & ~n44817;
  assign po844 = ~n44818 & n44819;
  assign n44821 = ~pi1115 & po980;
  assign n44822 = pi688 & ~po980;
  assign n44823 = ~pi962 & ~n44821;
  assign po845 = ~n44822 & n44823;
  assign n44825 = pi351 & n44774;
  assign n44826 = pi376 & n44226;
  assign n44827 = ~n44825 & ~n44826;
  assign n44828 = ~pi591 & ~n44827;
  assign n44829 = pi401 & ~pi592;
  assign n44830 = n44224 & n44829;
  assign n44831 = ~n44828 & ~n44830;
  assign n44832 = ~pi588 & ~n44831;
  assign n44833 = pi426 & n44177;
  assign n44834 = n44783 & n44833;
  assign n44835 = ~n44832 & ~n44834;
  assign n44836 = n44176 & ~n44835;
  assign n44837 = pi199 & ~pi1079;
  assign n44838 = ~pi199 & ~n40425;
  assign n44839 = ~n44176 & ~n44837;
  assign n44840 = ~n44838 & n44839;
  assign n44841 = ~n44836 & ~n44840;
  assign n44842 = n7578 & ~n44841;
  assign n44843 = pi798 & n44242;
  assign n44844 = ~pi658 & ~pi1135;
  assign n44845 = pi655 & pi1135;
  assign n44846 = pi1136 & ~n44844;
  assign n44847 = ~n44845 & n44846;
  assign n44848 = ~n44843 & ~n44847;
  assign n44849 = n44197 & ~n44848;
  assign n44850 = ~pi703 & pi1135;
  assign n44851 = pi752 & n44214;
  assign n44852 = ~pi843 & ~pi1136;
  assign n44853 = ~n44850 & ~n44852;
  assign n44854 = n44211 & n44853;
  assign n44855 = ~n44851 & n44854;
  assign n44856 = ~n44849 & ~n44855;
  assign n44857 = ~n7578 & ~n44856;
  assign po846 = n44842 | n44857;
  assign n44859 = ~pi690 & ~po980;
  assign n44860 = ~pi1108 & po980;
  assign n44861 = ~pi962 & ~n44859;
  assign po847 = ~n44860 & n44861;
  assign n44863 = ~pi691 & ~po980;
  assign n44864 = ~pi1107 & po980;
  assign n44865 = ~pi962 & ~n44863;
  assign po848 = ~n44864 & n44865;
  assign n44867 = pi352 & n44774;
  assign n44868 = pi317 & n44226;
  assign n44869 = ~n44867 & ~n44868;
  assign n44870 = ~pi591 & ~n44869;
  assign n44871 = pi402 & ~pi592;
  assign n44872 = n44224 & n44871;
  assign n44873 = ~n44870 & ~n44872;
  assign n44874 = ~pi588 & ~n44873;
  assign n44875 = pi427 & n44177;
  assign n44876 = n44783 & n44875;
  assign n44877 = ~n44874 & ~n44876;
  assign n44878 = n44176 & ~n44877;
  assign n44879 = pi199 & ~pi1078;
  assign n44880 = ~pi199 & ~n40437;
  assign n44881 = ~n44176 & ~n44879;
  assign n44882 = ~n44880 & n44881;
  assign n44883 = ~n44878 & ~n44882;
  assign n44884 = n7578 & ~n44883;
  assign n44885 = pi844 & n44242;
  assign n44886 = ~pi726 & pi1135;
  assign n44887 = pi770 & ~pi1135;
  assign n44888 = pi1136 & ~n44886;
  assign n44889 = ~n44887 & n44888;
  assign n44890 = pi1134 & ~n44885;
  assign n44891 = ~n44889 & n44890;
  assign n44892 = pi801 & n44242;
  assign n44893 = ~pi656 & ~pi1135;
  assign n44894 = pi649 & pi1135;
  assign n44895 = pi1136 & ~n44893;
  assign n44896 = ~n44894 & n44895;
  assign n44897 = ~pi1134 & ~n44892;
  assign n44898 = ~n44896 & n44897;
  assign n44899 = n44250 & ~n44891;
  assign n44900 = ~n44898 & n44899;
  assign po849 = n44884 | n44900;
  assign n44902 = ~pi1129 & po954;
  assign n44903 = pi693 & ~po954;
  assign n44904 = ~pi962 & ~n44902;
  assign po850 = ~n44903 & n44904;
  assign n44906 = ~pi1128 & po980;
  assign n44907 = pi694 & ~po980;
  assign n44908 = ~pi962 & ~n44906;
  assign po851 = ~n44907 & n44908;
  assign n44910 = ~pi1111 & po954;
  assign n44911 = pi695 & ~po954;
  assign n44912 = ~pi962 & ~n44910;
  assign po852 = ~n44911 & n44912;
  assign n44914 = ~pi696 & ~po980;
  assign n44915 = ~pi1100 & po980;
  assign n44916 = ~pi962 & ~n44914;
  assign po853 = ~n44915 & n44916;
  assign n44918 = ~pi1129 & po980;
  assign n44919 = pi697 & ~po980;
  assign n44920 = ~pi962 & ~n44918;
  assign po854 = ~n44919 & n44920;
  assign n44922 = ~pi1116 & po980;
  assign n44923 = pi698 & ~po980;
  assign n44924 = ~pi962 & ~n44922;
  assign po855 = ~n44923 & n44924;
  assign n44926 = ~pi699 & ~po980;
  assign n44927 = ~pi1103 & po980;
  assign n44928 = ~pi962 & ~n44926;
  assign po856 = ~n44927 & n44928;
  assign n44930 = ~pi700 & ~po980;
  assign n44931 = ~pi1110 & po980;
  assign n44932 = ~pi962 & ~n44930;
  assign po857 = ~n44931 & n44932;
  assign n44934 = ~pi1123 & po980;
  assign n44935 = pi701 & ~po980;
  assign n44936 = ~pi962 & ~n44934;
  assign po858 = ~n44935 & n44936;
  assign n44938 = ~pi1117 & po980;
  assign n44939 = pi702 & ~po980;
  assign n44940 = ~pi962 & ~n44938;
  assign po859 = ~n44939 & n44940;
  assign n44942 = ~pi703 & ~po980;
  assign n44943 = ~pi1124 & po980;
  assign n44944 = ~pi962 & ~n44942;
  assign po860 = ~n44943 & n44944;
  assign n44946 = ~pi1112 & po980;
  assign n44947 = pi704 & ~po980;
  assign n44948 = ~pi962 & ~n44946;
  assign po861 = ~n44947 & n44948;
  assign n44950 = ~pi705 & ~po980;
  assign n44951 = ~pi1125 & po980;
  assign n44952 = ~pi962 & ~n44950;
  assign po862 = ~n44951 & n44952;
  assign n44954 = ~pi706 & ~po980;
  assign n44955 = ~pi1105 & po980;
  assign n44956 = ~pi962 & ~n44954;
  assign po863 = ~n44955 & n44956;
  assign n44958 = ~pi627 & pi1135;
  assign n44959 = ~pi618 & ~pi1135;
  assign n44960 = ~pi1134 & ~n44958;
  assign n44961 = ~n44959 & n44960;
  assign n44962 = n44382 & n44961;
  assign n44963 = ~pi847 & ~pi1136;
  assign n44964 = pi753 & n44214;
  assign n44965 = pi702 & pi1135;
  assign n44966 = ~n44963 & ~n44965;
  assign n44967 = n44211 & n44966;
  assign n44968 = ~n44964 & n44967;
  assign n44969 = ~n7578 & ~n44962;
  assign n44970 = ~n44968 & n44969;
  assign n44971 = n7580 & n44176;
  assign n44972 = pi420 & pi588;
  assign n44973 = n44971 & n44972;
  assign n44974 = pi370 & n44180;
  assign n44975 = pi395 & pi591;
  assign n44976 = ~pi592 & n44975;
  assign n44977 = ~n44974 & ~n44976;
  assign n44978 = ~pi590 & ~n44977;
  assign n44979 = pi347 & n44178;
  assign n44980 = ~n44978 & ~n44979;
  assign n44981 = ~pi588 & n44176;
  assign n44982 = ~n44980 & n44981;
  assign n44983 = pi199 & ~pi1055;
  assign n44984 = ~pi200 & ~pi304;
  assign n44985 = pi200 & ~pi1048;
  assign n44986 = ~n44984 & ~n44985;
  assign n44987 = ~pi199 & ~n44986;
  assign n44988 = ~n44176 & ~n44983;
  assign n44989 = ~n44987 & n44988;
  assign n44990 = n7578 & ~n44973;
  assign n44991 = ~n44989 & n44990;
  assign n44992 = ~n44982 & n44991;
  assign po864 = ~n44970 & ~n44992;
  assign n44994 = pi199 & ~pi1058;
  assign n44995 = ~pi200 & ~pi305;
  assign n44996 = pi200 & ~pi1084;
  assign n44997 = ~n44995 & ~n44996;
  assign n44998 = ~pi199 & ~n44997;
  assign n44999 = ~n44176 & ~n44994;
  assign n45000 = ~n44998 & n44999;
  assign n45001 = n44176 & n44177;
  assign n45002 = pi459 & n44783;
  assign n45003 = n45001 & n45002;
  assign n45004 = n44176 & n44180;
  assign n45005 = pi442 & n45004;
  assign n45006 = ~pi592 & n44176;
  assign n45007 = pi328 & pi591;
  assign n45008 = n45006 & n45007;
  assign n45009 = ~n45005 & ~n45008;
  assign n45010 = ~pi590 & ~n45009;
  assign n45011 = pi321 & n44176;
  assign n45012 = n44178 & n45011;
  assign n45013 = ~n45010 & ~n45012;
  assign n45014 = ~pi588 & ~n45013;
  assign n45015 = n7578 & ~n45003;
  assign n45016 = ~n45000 & n45015;
  assign n45017 = ~n45014 & n45016;
  assign n45018 = ~pi660 & pi1135;
  assign n45019 = ~pi609 & ~pi1135;
  assign n45020 = ~pi1134 & ~n45018;
  assign n45021 = ~n45019 & n45020;
  assign n45022 = n44382 & n45021;
  assign n45023 = ~pi857 & ~pi1136;
  assign n45024 = pi754 & n44214;
  assign n45025 = pi709 & pi1135;
  assign n45026 = ~n45023 & ~n45025;
  assign n45027 = n44211 & n45026;
  assign n45028 = ~n45024 & n45027;
  assign n45029 = ~n7578 & ~n45022;
  assign n45030 = ~n45028 & n45029;
  assign po865 = ~n45017 & ~n45030;
  assign n45032 = ~pi1118 & po980;
  assign n45033 = pi709 & ~po980;
  assign n45034 = ~pi962 & ~n45032;
  assign po866 = ~n45033 & n45034;
  assign n45036 = ~pi710 & ~po954;
  assign n45037 = ~pi1106 & po954;
  assign n45038 = ~pi962 & ~n45036;
  assign po867 = ~n45037 & n45038;
  assign n45040 = ~pi647 & pi1135;
  assign n45041 = ~pi630 & ~pi1135;
  assign n45042 = ~pi1134 & ~n45040;
  assign n45043 = ~n45041 & n45042;
  assign n45044 = n44382 & n45043;
  assign n45045 = ~pi858 & ~pi1136;
  assign n45046 = pi755 & n44214;
  assign n45047 = pi725 & pi1135;
  assign n45048 = ~n45045 & ~n45047;
  assign n45049 = n44211 & n45048;
  assign n45050 = ~n45046 & n45049;
  assign n45051 = ~n7578 & ~n45044;
  assign n45052 = ~n45050 & n45051;
  assign n45053 = pi423 & pi588;
  assign n45054 = n44971 & n45053;
  assign n45055 = pi373 & n44180;
  assign n45056 = pi398 & pi591;
  assign n45057 = ~pi592 & n45056;
  assign n45058 = ~n45055 & ~n45057;
  assign n45059 = ~pi590 & ~n45058;
  assign n45060 = pi348 & n44178;
  assign n45061 = ~n45059 & ~n45060;
  assign n45062 = n44981 & ~n45061;
  assign n45063 = pi199 & ~pi1087;
  assign n45064 = ~pi200 & ~pi306;
  assign n45065 = pi200 & ~pi1059;
  assign n45066 = ~n45064 & ~n45065;
  assign n45067 = ~pi199 & ~n45066;
  assign n45068 = ~n44176 & ~n45063;
  assign n45069 = ~n45067 & n45068;
  assign n45070 = n7578 & ~n45054;
  assign n45071 = ~n45069 & n45070;
  assign n45072 = ~n45062 & n45071;
  assign po868 = ~n45052 & ~n45072;
  assign n45074 = ~pi715 & pi1135;
  assign n45075 = ~pi644 & ~pi1135;
  assign n45076 = ~pi1134 & ~n45074;
  assign n45077 = ~n45075 & n45076;
  assign n45078 = n44382 & n45077;
  assign n45079 = pi701 & pi1135;
  assign n45080 = ~pi842 & ~pi1136;
  assign n45081 = pi751 & n44214;
  assign n45082 = ~n45079 & ~n45080;
  assign n45083 = n44211 & n45082;
  assign n45084 = ~n45081 & n45083;
  assign n45085 = ~n45078 & ~n45084;
  assign n45086 = ~n7578 & ~n45085;
  assign n45087 = pi425 & n44177;
  assign n45088 = n44783 & n45087;
  assign n45089 = pi374 & n44180;
  assign n45090 = pi400 & pi591;
  assign n45091 = ~pi592 & n45090;
  assign n45092 = ~n45089 & ~n45091;
  assign n45093 = ~pi590 & ~n45092;
  assign n45094 = pi350 & n44178;
  assign n45095 = ~n45093 & ~n45094;
  assign n45096 = ~pi588 & ~n45095;
  assign n45097 = n44176 & ~n45088;
  assign n45098 = ~n45096 & n45097;
  assign n45099 = pi199 & pi1035;
  assign n45100 = pi298 & n10421;
  assign n45101 = pi1044 & n11035;
  assign n45102 = ~n44176 & ~n45099;
  assign n45103 = ~n45100 & n45102;
  assign n45104 = ~n45101 & n45103;
  assign n45105 = n7578 & ~n45104;
  assign n45106 = ~n45098 & n45105;
  assign po869 = n45086 | n45106;
  assign n45108 = ~pi628 & pi1135;
  assign n45109 = ~pi629 & ~pi1135;
  assign n45110 = ~pi1134 & ~n45108;
  assign n45111 = ~n45109 & n45110;
  assign n45112 = n44382 & n45111;
  assign n45113 = ~pi854 & ~pi1136;
  assign n45114 = pi756 & n44214;
  assign n45115 = pi734 & pi1135;
  assign n45116 = ~n45113 & ~n45115;
  assign n45117 = n44211 & n45116;
  assign n45118 = ~n45114 & n45117;
  assign n45119 = ~n7578 & ~n45112;
  assign n45120 = ~n45118 & n45119;
  assign n45121 = pi421 & pi588;
  assign n45122 = n44971 & n45121;
  assign n45123 = pi371 & n44180;
  assign n45124 = pi396 & pi591;
  assign n45125 = ~pi592 & n45124;
  assign n45126 = ~n45123 & ~n45125;
  assign n45127 = ~pi590 & ~n45126;
  assign n45128 = pi322 & n44178;
  assign n45129 = ~n45127 & ~n45128;
  assign n45130 = n44981 & ~n45129;
  assign n45131 = pi199 & ~pi1051;
  assign n45132 = ~pi200 & ~pi309;
  assign n45133 = pi200 & ~pi1072;
  assign n45134 = ~n45132 & ~n45133;
  assign n45135 = ~pi199 & ~n45134;
  assign n45136 = ~n44176 & ~n45131;
  assign n45137 = ~n45135 & n45136;
  assign n45138 = n7578 & ~n45122;
  assign n45139 = ~n45137 & n45138;
  assign n45140 = ~n45130 & n45139;
  assign po870 = ~n45120 & ~n45140;
  assign n45142 = pi461 & n44774;
  assign n45143 = pi439 & n44226;
  assign n45144 = ~n45142 & ~n45143;
  assign n45145 = ~pi591 & ~n45144;
  assign n45146 = pi326 & ~pi592;
  assign n45147 = n44224 & n45146;
  assign n45148 = ~n45145 & ~n45147;
  assign n45149 = ~pi588 & ~n45148;
  assign n45150 = pi449 & n44177;
  assign n45151 = n44783 & n45150;
  assign n45152 = ~n45149 & ~n45151;
  assign n45153 = n44176 & ~n45152;
  assign n45154 = pi199 & ~pi1057;
  assign n45155 = ~n44176 & ~n45154;
  assign n45156 = ~n39954 & n45155;
  assign n45157 = ~n45153 & ~n45156;
  assign n45158 = n7578 & ~n45157;
  assign n45159 = pi867 & n44242;
  assign n45160 = pi762 & ~pi1135;
  assign n45161 = pi697 & pi1135;
  assign n45162 = pi1136 & ~n45160;
  assign n45163 = ~n45161 & n45162;
  assign n45164 = ~n45159 & ~n45163;
  assign n45165 = n44210 & ~n45164;
  assign n45166 = ~pi653 & ~pi1135;
  assign n45167 = pi693 & pi1135;
  assign n45168 = pi1136 & ~n45166;
  assign n45169 = ~n45167 & n45168;
  assign n45170 = pi816 & n44196;
  assign n45171 = n44242 & n45170;
  assign n45172 = ~n45169 & ~n45171;
  assign n45173 = n44801 & ~n45172;
  assign n45174 = ~n45165 & ~n45173;
  assign n45175 = ~n7578 & ~n45174;
  assign po871 = n45158 | n45175;
  assign n45177 = ~pi715 & ~po954;
  assign n45178 = ~pi1123 & po954;
  assign n45179 = ~pi962 & ~n45177;
  assign po872 = ~n45178 & n45179;
  assign n45181 = pi199 & ~pi1043;
  assign n45182 = ~pi200 & ~pi307;
  assign n45183 = pi200 & ~pi1053;
  assign n45184 = ~n45182 & ~n45183;
  assign n45185 = ~pi199 & ~n45184;
  assign n45186 = ~n44176 & ~n45181;
  assign n45187 = ~n45185 & n45186;
  assign n45188 = pi454 & n44783;
  assign n45189 = n45001 & n45188;
  assign n45190 = pi440 & n45004;
  assign n45191 = pi329 & pi591;
  assign n45192 = n45006 & n45191;
  assign n45193 = ~n45190 & ~n45192;
  assign n45194 = ~pi590 & ~n45193;
  assign n45195 = pi349 & n44176;
  assign n45196 = n44178 & n45195;
  assign n45197 = ~n45194 & ~n45196;
  assign n45198 = ~pi588 & ~n45197;
  assign n45199 = n7578 & ~n45189;
  assign n45200 = ~n45187 & n45199;
  assign n45201 = ~n45198 & n45200;
  assign n45202 = ~pi641 & pi1135;
  assign n45203 = ~pi626 & ~pi1135;
  assign n45204 = ~pi1134 & ~n45202;
  assign n45205 = ~n45203 & n45204;
  assign n45206 = n44382 & n45205;
  assign n45207 = ~pi845 & ~pi1136;
  assign n45208 = pi761 & n44214;
  assign n45209 = pi738 & pi1135;
  assign n45210 = ~n45207 & ~n45209;
  assign n45211 = n44211 & n45210;
  assign n45212 = ~n45208 & n45211;
  assign n45213 = ~n7578 & ~n45206;
  assign n45214 = ~n45212 & n45213;
  assign po873 = ~n45201 & ~n45214;
  assign n45216 = pi377 & n44180;
  assign n45217 = pi318 & pi591;
  assign n45218 = ~pi592 & n45217;
  assign n45219 = ~n45216 & ~n45218;
  assign n45220 = ~pi590 & ~n45219;
  assign n45221 = pi462 & n44178;
  assign n45222 = ~n45220 & ~n45221;
  assign n45223 = n44981 & ~n45222;
  assign n45224 = pi199 & ~pi1074;
  assign n45225 = ~pi199 & ~n40431;
  assign n45226 = ~n44176 & ~n45224;
  assign n45227 = ~n45225 & n45226;
  assign n45228 = pi448 & pi588;
  assign n45229 = n44971 & n45228;
  assign n45230 = ~n45227 & ~n45229;
  assign n45231 = ~n45223 & n45230;
  assign n45232 = n7578 & ~n45231;
  assign n45233 = pi800 & n44242;
  assign n45234 = ~pi645 & ~pi1135;
  assign n45235 = pi669 & pi1135;
  assign n45236 = pi1136 & ~n45234;
  assign n45237 = ~n45235 & n45236;
  assign n45238 = ~n45233 & ~n45237;
  assign n45239 = n44197 & ~n45238;
  assign n45240 = ~pi705 & pi1135;
  assign n45241 = pi768 & n44214;
  assign n45242 = ~pi839 & ~pi1136;
  assign n45243 = ~n45240 & ~n45242;
  assign n45244 = n44211 & n45243;
  assign n45245 = ~n45241 & n45244;
  assign n45246 = ~n45239 & ~n45245;
  assign n45247 = ~n7578 & ~n45246;
  assign po874 = n45232 | n45247;
  assign n45249 = pi199 & ~pi1080;
  assign n45250 = ~pi200 & ~pi303;
  assign n45251 = pi200 & ~pi1049;
  assign n45252 = ~n45250 & ~n45251;
  assign n45253 = ~pi199 & ~n45252;
  assign n45254 = ~n44176 & ~n45249;
  assign n45255 = ~n45253 & n45254;
  assign n45256 = pi419 & n44783;
  assign n45257 = n45001 & n45256;
  assign n45258 = pi369 & n45004;
  assign n45259 = pi394 & pi591;
  assign n45260 = n45006 & n45259;
  assign n45261 = ~n45258 & ~n45260;
  assign n45262 = ~pi590 & ~n45261;
  assign n45263 = pi315 & n44176;
  assign n45264 = n44178 & n45263;
  assign n45265 = ~n45262 & ~n45264;
  assign n45266 = ~pi588 & ~n45265;
  assign n45267 = n7578 & ~n45257;
  assign n45268 = ~n45255 & n45267;
  assign n45269 = ~n45266 & n45268;
  assign n45270 = ~pi625 & pi1135;
  assign n45271 = ~pi608 & ~pi1135;
  assign n45272 = ~pi1134 & ~n45270;
  assign n45273 = ~n45271 & n45272;
  assign n45274 = n44382 & n45273;
  assign n45275 = ~pi853 & ~pi1136;
  assign n45276 = pi767 & n44214;
  assign n45277 = pi698 & pi1135;
  assign n45278 = ~n45275 & ~n45277;
  assign n45279 = n44211 & n45278;
  assign n45280 = ~n45276 & n45279;
  assign n45281 = ~n7578 & ~n45274;
  assign n45282 = ~n45280 & n45281;
  assign po875 = ~n45269 & ~n45282;
  assign n45284 = pi378 & n44180;
  assign n45285 = pi325 & pi591;
  assign n45286 = ~pi592 & n45285;
  assign n45287 = ~n45284 & ~n45286;
  assign n45288 = ~pi590 & ~n45287;
  assign n45289 = pi353 & n44178;
  assign n45290 = ~n45288 & ~n45289;
  assign n45291 = n44981 & ~n45290;
  assign n45292 = pi199 & ~pi1063;
  assign n45293 = ~pi199 & ~n40443;
  assign n45294 = ~n44176 & ~n45292;
  assign n45295 = ~n45293 & n45294;
  assign n45296 = pi451 & pi588;
  assign n45297 = n44971 & n45296;
  assign n45298 = ~n45295 & ~n45297;
  assign n45299 = ~n45291 & n45298;
  assign n45300 = n7578 & ~n45299;
  assign n45301 = pi807 & n44242;
  assign n45302 = ~pi636 & ~pi1135;
  assign n45303 = pi650 & pi1135;
  assign n45304 = pi1136 & ~n45302;
  assign n45305 = ~n45303 & n45304;
  assign n45306 = ~n45301 & ~n45305;
  assign n45307 = n44197 & ~n45306;
  assign n45308 = ~pi687 & pi1135;
  assign n45309 = pi774 & n44214;
  assign n45310 = ~pi868 & ~pi1136;
  assign n45311 = ~n45308 & ~n45310;
  assign n45312 = n44211 & n45311;
  assign n45313 = ~n45309 & n45312;
  assign n45314 = ~n45307 & ~n45313;
  assign n45315 = ~n7578 & ~n45314;
  assign po876 = n45300 | n45315;
  assign n45317 = pi356 & n44774;
  assign n45318 = pi381 & n44226;
  assign n45319 = ~n45317 & ~n45318;
  assign n45320 = ~pi591 & ~n45319;
  assign n45321 = pi405 & ~pi592;
  assign n45322 = n44224 & n45321;
  assign n45323 = ~n45320 & ~n45322;
  assign n45324 = ~pi588 & ~n45323;
  assign n45325 = pi445 & n44177;
  assign n45326 = n44783 & n45325;
  assign n45327 = ~n45324 & ~n45326;
  assign n45328 = n44176 & ~n45327;
  assign n45329 = pi199 & ~pi1081;
  assign n45330 = ~n44176 & ~n45329;
  assign n45331 = ~n40463 & n45330;
  assign n45332 = ~n45328 & ~n45331;
  assign n45333 = n7578 & ~n45332;
  assign n45334 = pi880 & n44242;
  assign n45335 = pi750 & ~pi1135;
  assign n45336 = pi684 & pi1135;
  assign n45337 = pi1136 & ~n45335;
  assign n45338 = ~n45336 & n45337;
  assign n45339 = ~n45334 & ~n45338;
  assign n45340 = n44210 & ~n45339;
  assign n45341 = ~pi651 & ~pi1135;
  assign n45342 = pi654 & pi1135;
  assign n45343 = pi1136 & ~n45341;
  assign n45344 = ~n45342 & n45343;
  assign n45345 = pi794 & n44196;
  assign n45346 = n44242 & n45345;
  assign n45347 = ~n45344 & ~n45346;
  assign n45348 = n44801 & ~n45347;
  assign n45349 = ~n45340 & ~n45348;
  assign n45350 = ~n7578 & ~n45349;
  assign po877 = n45333 | n45350;
  assign n45352 = ~pi945 & pi988;
  assign n45353 = pi731 & n45352;
  assign n45354 = pi721 & pi813;
  assign n45355 = pi765 & ~pi798;
  assign n45356 = ~pi765 & pi798;
  assign n45357 = ~n45355 & ~n45356;
  assign n45358 = pi807 & n45357;
  assign n45359 = pi747 & n45358;
  assign n45360 = ~pi747 & ~pi807;
  assign n45361 = n45357 & n45360;
  assign n45362 = ~n45359 & ~n45361;
  assign n45363 = ~pi771 & ~pi800;
  assign n45364 = pi771 & pi800;
  assign n45365 = ~n45363 & ~n45364;
  assign n45366 = ~pi769 & ~pi794;
  assign n45367 = pi769 & pi794;
  assign n45368 = ~n45366 & ~n45367;
  assign n45369 = ~n45365 & ~n45368;
  assign n45370 = ~n45362 & n45369;
  assign n45371 = pi773 & ~pi801;
  assign n45372 = ~pi773 & pi801;
  assign n45373 = ~n45371 & ~n45372;
  assign n45374 = n45370 & n45373;
  assign n45375 = n45354 & n45374;
  assign n45376 = ~pi721 & ~pi813;
  assign n45377 = pi794 & ~n45365;
  assign n45378 = pi801 & n45376;
  assign n45379 = n45358 & n45378;
  assign n45380 = n45377 & n45379;
  assign n45381 = ~n45375 & ~n45380;
  assign n45382 = pi816 & ~n45381;
  assign n45383 = pi747 & pi773;
  assign n45384 = pi769 & n45383;
  assign n45385 = pi721 & n45384;
  assign n45386 = ~pi721 & ~n45384;
  assign n45387 = pi775 & ~n45385;
  assign n45388 = ~n45386 & n45387;
  assign n45389 = ~n45382 & n45388;
  assign n45390 = pi795 & ~n45389;
  assign n45391 = pi721 & ~pi775;
  assign n45392 = ~n45388 & ~n45391;
  assign n45393 = n45353 & ~n45392;
  assign n45394 = ~n45390 & n45393;
  assign n45395 = ~pi816 & n45375;
  assign n45396 = n45391 & ~n45395;
  assign n45397 = ~pi731 & ~pi795;
  assign n45398 = pi731 & pi795;
  assign n45399 = ~n45397 & ~n45398;
  assign n45400 = ~pi775 & ~pi816;
  assign n45401 = pi775 & pi816;
  assign n45402 = ~n45400 & ~n45401;
  assign n45403 = ~n45354 & ~n45376;
  assign n45404 = ~n45402 & ~n45403;
  assign n45405 = n45374 & n45404;
  assign po978 = ~n45399 & n45405;
  assign n45407 = ~n45353 & ~po978;
  assign n45408 = pi721 & n45407;
  assign n45409 = ~n45396 & ~n45408;
  assign po878 = n45394 | ~n45409;
  assign n45411 = pi379 & n44180;
  assign n45412 = pi403 & pi591;
  assign n45413 = ~pi592 & n45412;
  assign n45414 = ~n45411 & ~n45413;
  assign n45415 = ~pi590 & ~n45414;
  assign n45416 = pi354 & n44178;
  assign n45417 = ~n45415 & ~n45416;
  assign n45418 = n44981 & ~n45417;
  assign n45419 = pi199 & ~pi1045;
  assign n45420 = ~pi199 & ~n40449;
  assign n45421 = ~n44176 & ~n45419;
  assign n45422 = ~n45420 & n45421;
  assign n45423 = pi428 & pi588;
  assign n45424 = n44971 & n45423;
  assign n45425 = ~n45422 & ~n45424;
  assign n45426 = ~n45418 & n45425;
  assign n45427 = n7578 & ~n45426;
  assign n45428 = ~pi795 & ~pi1134;
  assign n45429 = ~pi851 & pi1134;
  assign n45430 = ~pi1136 & ~n45428;
  assign n45431 = ~n45429 & n45430;
  assign n45432 = ~pi640 & ~pi1134;
  assign n45433 = pi776 & pi1134;
  assign n45434 = pi1136 & ~n45432;
  assign n45435 = ~n45433 & n45434;
  assign n45436 = ~n45431 & ~n45435;
  assign n45437 = ~pi1135 & ~n45436;
  assign n45438 = pi694 & pi1134;
  assign n45439 = pi732 & ~pi1134;
  assign n45440 = pi1135 & pi1136;
  assign n45441 = ~n45438 & n45440;
  assign n45442 = ~n45439 & n45441;
  assign n45443 = ~n45437 & ~n45442;
  assign n45444 = n44250 & ~n45443;
  assign po879 = n45427 | n45444;
  assign n45446 = ~pi1111 & po980;
  assign n45447 = pi723 & ~po980;
  assign n45448 = ~pi962 & ~n45446;
  assign po880 = ~n45447 & n45448;
  assign n45450 = ~pi1114 & po980;
  assign n45451 = pi724 & ~po980;
  assign n45452 = ~pi962 & ~n45450;
  assign po881 = ~n45451 & n45452;
  assign n45454 = ~pi1120 & po980;
  assign n45455 = pi725 & ~po980;
  assign n45456 = ~pi962 & ~n45454;
  assign po882 = ~n45455 & n45456;
  assign n45458 = ~pi726 & ~po980;
  assign n45459 = ~pi1126 & po980;
  assign n45460 = ~pi962 & ~n45458;
  assign po883 = ~n45459 & n45460;
  assign n45462 = ~pi727 & ~po980;
  assign n45463 = ~pi1102 & po980;
  assign n45464 = ~pi962 & ~n45462;
  assign po884 = ~n45463 & n45464;
  assign n45466 = ~pi1131 & po980;
  assign n45467 = pi728 & ~po980;
  assign n45468 = ~pi962 & ~n45466;
  assign po885 = ~n45467 & n45468;
  assign n45470 = ~pi729 & ~po980;
  assign n45471 = ~pi1104 & po980;
  assign n45472 = ~pi962 & ~n45470;
  assign po886 = ~n45471 & n45472;
  assign n45474 = ~pi730 & ~po980;
  assign n45475 = ~pi1106 & po980;
  assign n45476 = ~pi962 & ~n45474;
  assign po887 = ~n45475 & n45476;
  assign n45478 = pi795 & n45405;
  assign n45479 = n45352 & n45383;
  assign n45480 = pi731 & ~n45479;
  assign n45481 = ~n45478 & n45480;
  assign n45482 = ~n45399 & n45404;
  assign n45483 = pi801 & n45370;
  assign n45484 = n45482 & n45483;
  assign n45485 = ~pi731 & n45479;
  assign n45486 = ~n45484 & n45485;
  assign po888 = n45481 | n45486;
  assign n45488 = ~pi1128 & po954;
  assign n45489 = pi732 & ~po954;
  assign n45490 = ~pi962 & ~n45488;
  assign po889 = ~n45489 & n45490;
  assign n45492 = pi199 & ~pi1047;
  assign n45493 = ~pi200 & ~pi308;
  assign n45494 = pi200 & ~pi1037;
  assign n45495 = ~n45493 & ~n45494;
  assign n45496 = ~pi199 & ~n45495;
  assign n45497 = ~n44176 & ~n45492;
  assign n45498 = ~n45496 & n45497;
  assign n45499 = pi424 & n44783;
  assign n45500 = n45001 & n45499;
  assign n45501 = pi375 & n45004;
  assign n45502 = pi399 & pi591;
  assign n45503 = n45006 & n45502;
  assign n45504 = ~n45501 & ~n45503;
  assign n45505 = ~pi590 & ~n45504;
  assign n45506 = pi316 & n44176;
  assign n45507 = n44178 & n45506;
  assign n45508 = ~n45505 & ~n45507;
  assign n45509 = ~pi588 & ~n45508;
  assign n45510 = n7578 & ~n45500;
  assign n45511 = ~n45498 & n45510;
  assign n45512 = ~n45509 & n45511;
  assign n45513 = ~pi648 & pi1135;
  assign n45514 = ~pi619 & ~pi1135;
  assign n45515 = ~pi1134 & ~n45513;
  assign n45516 = ~n45514 & n45515;
  assign n45517 = n44382 & n45516;
  assign n45518 = ~pi838 & ~pi1136;
  assign n45519 = pi777 & n44214;
  assign n45520 = pi737 & pi1135;
  assign n45521 = ~n45518 & ~n45520;
  assign n45522 = n44211 & n45521;
  assign n45523 = ~n45519 & n45522;
  assign n45524 = ~n7578 & ~n45517;
  assign n45525 = ~n45523 & n45524;
  assign po890 = ~n45512 & ~n45525;
  assign n45527 = ~pi1119 & po980;
  assign n45528 = pi734 & ~po980;
  assign n45529 = ~pi962 & ~n45527;
  assign po891 = ~n45528 & n45529;
  assign n45531 = ~pi735 & ~po980;
  assign n45532 = ~pi1109 & po980;
  assign n45533 = ~pi962 & ~n45531;
  assign po892 = ~n45532 & n45533;
  assign n45535 = ~pi736 & ~po980;
  assign n45536 = ~pi1101 & po980;
  assign n45537 = ~pi962 & ~n45535;
  assign po893 = ~n45536 & n45537;
  assign n45539 = ~pi1122 & po980;
  assign n45540 = pi737 & ~po980;
  assign n45541 = ~pi962 & ~n45539;
  assign po894 = ~n45540 & n45541;
  assign n45543 = ~pi1121 & po980;
  assign n45544 = pi738 & ~po980;
  assign n45545 = ~pi962 & ~n45543;
  assign po895 = ~n45544 & n45545;
  assign n45547 = ~pi952 & ~pi1061;
  assign n45548 = n43904 & n45547;
  assign po988 = pi832 & n45548;
  assign n45550 = pi1108 & po988;
  assign n45551 = pi739 & ~po988;
  assign n45552 = ~pi966 & ~n45550;
  assign po896 = n45551 | ~n45552;
  assign n45554 = ~pi741 & ~po988;
  assign n45555 = pi1114 & po988;
  assign n45556 = ~pi966 & ~n45554;
  assign po898 = n45555 | ~n45556;
  assign n45558 = ~pi742 & ~po988;
  assign n45559 = pi1112 & po988;
  assign n45560 = ~pi966 & ~n45558;
  assign po899 = n45559 | ~n45560;
  assign n45562 = pi1109 & po988;
  assign n45563 = pi743 & ~po988;
  assign n45564 = ~pi966 & ~n45562;
  assign po900 = n45563 | ~n45564;
  assign n45566 = ~pi744 & ~po988;
  assign n45567 = pi1131 & po988;
  assign n45568 = ~pi966 & ~n45566;
  assign po901 = n45567 | ~n45568;
  assign n45570 = ~pi745 & ~po988;
  assign n45571 = pi1111 & po988;
  assign n45572 = ~pi966 & ~n45570;
  assign po902 = n45571 | ~n45572;
  assign n45574 = pi1104 & po988;
  assign n45575 = pi746 & ~po988;
  assign n45576 = ~pi966 & ~n45574;
  assign po903 = n45575 | ~n45576;
  assign n45578 = pi773 & n45352;
  assign n45579 = ~pi747 & ~n45578;
  assign n45580 = pi801 & n45361;
  assign n45581 = n45373 & ~n45578;
  assign n45582 = n45358 & n45581;
  assign n45583 = ~n45580 & ~n45582;
  assign n45584 = n45369 & n45482;
  assign n45585 = ~n45583 & n45584;
  assign n45586 = ~n45479 & ~n45579;
  assign po904 = ~n45585 & n45586;
  assign n45588 = pi1106 & po988;
  assign n45589 = pi748 & ~po988;
  assign n45590 = ~pi966 & ~n45588;
  assign po905 = n45589 | ~n45590;
  assign n45592 = pi1105 & po988;
  assign n45593 = pi749 & ~po988;
  assign n45594 = ~pi966 & ~n45592;
  assign po906 = n45593 | ~n45594;
  assign n45596 = ~pi750 & ~po988;
  assign n45597 = pi1130 & po988;
  assign n45598 = ~pi966 & ~n45596;
  assign po907 = n45597 | ~n45598;
  assign n45600 = ~pi751 & ~po988;
  assign n45601 = pi1123 & po988;
  assign n45602 = ~pi966 & ~n45600;
  assign po908 = n45601 | ~n45602;
  assign n45604 = ~pi752 & ~po988;
  assign n45605 = pi1124 & po988;
  assign n45606 = ~pi966 & ~n45604;
  assign po909 = n45605 | ~n45606;
  assign n45608 = ~pi753 & ~po988;
  assign n45609 = pi1117 & po988;
  assign n45610 = ~pi966 & ~n45608;
  assign po910 = n45609 | ~n45610;
  assign n45612 = ~pi754 & ~po988;
  assign n45613 = pi1118 & po988;
  assign n45614 = ~pi966 & ~n45612;
  assign po911 = n45613 | ~n45614;
  assign n45616 = ~pi755 & ~po988;
  assign n45617 = pi1120 & po988;
  assign n45618 = ~pi966 & ~n45616;
  assign po912 = n45617 | ~n45618;
  assign n45620 = ~pi756 & ~po988;
  assign n45621 = pi1119 & po988;
  assign n45622 = ~pi966 & ~n45620;
  assign po913 = n45621 | ~n45622;
  assign n45624 = ~pi757 & ~po988;
  assign n45625 = pi1113 & po988;
  assign n45626 = ~pi966 & ~n45624;
  assign po914 = n45625 | ~n45626;
  assign n45628 = pi1101 & po988;
  assign n45629 = pi758 & ~po988;
  assign n45630 = ~pi966 & ~n45628;
  assign po915 = n45629 | ~n45630;
  assign n45632 = ~pi759 & ~po988;
  assign n45633 = n43902 & n45548;
  assign n45634 = ~n45632 & ~n45633;
  assign po916 = pi966 | n45634;
  assign n45636 = ~pi760 & ~po988;
  assign n45637 = pi1115 & po988;
  assign n45638 = ~pi966 & ~n45636;
  assign po917 = n45637 | ~n45638;
  assign n45640 = ~pi761 & ~po988;
  assign n45641 = pi1121 & po988;
  assign n45642 = ~pi966 & ~n45640;
  assign po918 = n45641 | ~n45642;
  assign n45644 = ~pi762 & ~po988;
  assign n45645 = pi1129 & po988;
  assign n45646 = ~pi966 & ~n45644;
  assign po919 = n45645 | ~n45646;
  assign n45648 = pi1103 & po988;
  assign n45649 = pi763 & ~po988;
  assign n45650 = ~pi966 & ~n45648;
  assign po920 = n45649 | ~n45650;
  assign n45652 = pi1107 & po988;
  assign n45653 = pi764 & ~po988;
  assign n45654 = ~pi966 & ~n45652;
  assign po921 = n45653 | ~n45654;
  assign n45656 = pi945 & ~po978;
  assign n45657 = pi765 & ~n45656;
  assign n45658 = ~pi765 & ~pi773;
  assign n45659 = ~n45364 & n45658;
  assign n45660 = ~n45367 & n45659;
  assign n45661 = ~n45359 & n45660;
  assign n45662 = n45374 & ~n45661;
  assign n45663 = ~pi721 & ~pi731;
  assign n45664 = ~pi775 & n45663;
  assign n45665 = ~n45662 & n45664;
  assign po963 = po978 & ~n45665;
  assign n45667 = ~pi945 & ~po963;
  assign n45668 = ~pi765 & ~n45667;
  assign po922 = ~n45657 & ~n45668;
  assign n45670 = pi1110 & po988;
  assign n45671 = pi766 & ~po988;
  assign n45672 = ~pi966 & ~n45670;
  assign po923 = n45671 | ~n45672;
  assign n45674 = ~pi767 & ~po988;
  assign n45675 = pi1116 & po988;
  assign n45676 = ~pi966 & ~n45674;
  assign po924 = n45675 | ~n45676;
  assign n45678 = ~pi768 & ~po988;
  assign n45679 = pi1125 & po988;
  assign n45680 = ~pi966 & ~n45678;
  assign po925 = n45679 | ~n45680;
  assign n45682 = pi769 & n45407;
  assign n45683 = n45401 & ~n45403;
  assign n45684 = n45374 & n45683;
  assign n45685 = ~pi775 & n45373;
  assign n45686 = n45377 & n45685;
  assign n45687 = n45404 & n45686;
  assign n45688 = ~n45362 & n45687;
  assign n45689 = ~n45684 & ~n45688;
  assign n45690 = pi795 & ~n45689;
  assign n45691 = pi775 & n45383;
  assign n45692 = ~pi769 & ~n45691;
  assign n45693 = pi769 & n45691;
  assign n45694 = n45353 & ~n45692;
  assign n45695 = ~n45693 & n45694;
  assign n45696 = ~n45690 & n45695;
  assign po926 = n45682 | n45696;
  assign n45698 = ~pi770 & ~po988;
  assign n45699 = pi1126 & po988;
  assign n45700 = ~pi966 & ~n45698;
  assign po927 = n45699 | ~n45700;
  assign n45702 = pi987 & n45667;
  assign n45703 = pi771 & n45656;
  assign po928 = n45702 | n45703;
  assign n45705 = pi1102 & po988;
  assign n45706 = pi772 & ~po988;
  assign n45707 = ~pi966 & ~n45705;
  assign po929 = n45706 | ~n45707;
  assign n45709 = ~n45483 & po963;
  assign n45710 = n45352 & ~n45709;
  assign n45711 = pi773 & ~n45484;
  assign n45712 = ~n45710 & ~n45711;
  assign po930 = ~n45578 & ~n45712;
  assign n45714 = ~pi774 & ~po988;
  assign n45715 = pi1127 & po988;
  assign n45716 = ~pi966 & ~n45714;
  assign po931 = n45715 | ~n45716;
  assign n45718 = pi775 & ~po978;
  assign n45719 = pi731 & ~pi945;
  assign n45720 = pi765 & pi771;
  assign n45721 = n45383 & n45720;
  assign n45722 = pi795 & pi800;
  assign n45723 = pi801 & ~pi816;
  assign n45724 = n45722 & n45723;
  assign n45725 = ~n45368 & n45724;
  assign n45726 = ~n45403 & n45725;
  assign n45727 = ~n45362 & n45726;
  assign n45728 = n45721 & ~n45727;
  assign n45729 = ~pi775 & ~n45728;
  assign n45730 = n45719 & ~n45729;
  assign n45731 = ~n45718 & ~n45730;
  assign n45732 = ~n45478 & ~n45721;
  assign n45733 = pi775 & n45719;
  assign n45734 = ~n45732 & n45733;
  assign po932 = ~n45731 & ~n45734;
  assign n45736 = ~pi776 & ~po988;
  assign n45737 = pi1128 & po988;
  assign n45738 = ~pi966 & ~n45736;
  assign po933 = n45737 | ~n45738;
  assign n45740 = ~pi777 & ~po988;
  assign n45741 = pi1122 & po988;
  assign n45742 = ~pi966 & ~n45740;
  assign po934 = n45741 | ~n45742;
  assign n45744 = pi832 & pi956;
  assign n45745 = ~pi1046 & ~pi1083;
  assign n45746 = pi1085 & n45745;
  assign n45747 = n45744 & n45746;
  assign n45748 = ~pi968 & n45747;
  assign n45749 = pi778 & ~n45748;
  assign n45750 = pi1100 & n45748;
  assign po935 = n45749 | n45750;
  assign po936 = ~pi779 | n43963;
  assign po937 = ~pi780 | n43872;
  assign n45754 = pi781 & ~n45748;
  assign n45755 = pi1101 & n45748;
  assign po938 = n45754 | n45755;
  assign n45757 = ~n39960 & ~n43916;
  assign po939 = n43871 | ~n45757;
  assign n45759 = pi783 & ~n45748;
  assign n45760 = pi1109 & n45748;
  assign po940 = n45759 | n45760;
  assign n45762 = pi784 & ~n45748;
  assign n45763 = pi1110 & n45748;
  assign po941 = n45762 | n45763;
  assign n45765 = pi785 & ~n45748;
  assign n45766 = pi1102 & n45748;
  assign po942 = n45765 | n45766;
  assign n45768 = ~pi786 & pi954;
  assign n45769 = ~pi24 & ~pi954;
  assign po943 = n45768 | n45769;
  assign n45771 = pi787 & ~n45748;
  assign n45772 = pi1104 & n45748;
  assign po944 = n45771 | n45772;
  assign n45774 = pi788 & ~n45748;
  assign n45775 = pi1105 & n45748;
  assign po945 = n45774 | n45775;
  assign n45777 = pi789 & ~n45748;
  assign n45778 = pi1106 & n45748;
  assign po946 = n45777 | n45778;
  assign n45780 = pi790 & ~n45748;
  assign n45781 = pi1107 & n45748;
  assign po947 = n45780 | n45781;
  assign n45783 = pi791 & ~n45748;
  assign n45784 = pi1108 & n45748;
  assign po948 = n45783 | n45784;
  assign n45786 = pi792 & ~n45748;
  assign n45787 = pi1103 & n45748;
  assign po949 = n45786 | n45787;
  assign n45789 = pi968 & n45747;
  assign n45790 = pi794 & ~n45789;
  assign n45791 = pi1130 & n45789;
  assign po951 = n45790 | n45791;
  assign n45793 = pi795 & ~n45789;
  assign n45794 = pi1128 & n45789;
  assign po952 = n45793 | n45794;
  assign n45796 = pi266 & ~pi269;
  assign n45797 = pi278 & pi279;
  assign n45798 = ~pi280 & n45797;
  assign n45799 = n45796 & n45798;
  assign n45800 = ~pi281 & n45799;
  assign n45801 = n44155 & n45800;
  assign n45802 = pi264 & ~n45801;
  assign n45803 = ~pi264 & n45801;
  assign po953 = ~n45802 & ~n45803;
  assign n45805 = pi798 & ~n45789;
  assign n45806 = pi1124 & n45789;
  assign po955 = n45805 | n45806;
  assign n45808 = pi799 & ~n45789;
  assign n45809 = ~pi1107 & n45789;
  assign po956 = ~n45808 & ~n45809;
  assign n45811 = pi800 & ~n45789;
  assign n45812 = pi1125 & n45789;
  assign po957 = n45811 | n45812;
  assign n45814 = pi801 & ~n45789;
  assign n45815 = pi1126 & n45789;
  assign po958 = n45814 | n45815;
  assign n45817 = pi803 & ~n45789;
  assign n45818 = ~pi1106 & n45789;
  assign po960 = ~n45817 & ~n45818;
  assign n45820 = pi804 & ~n45789;
  assign n45821 = pi1109 & n45789;
  assign po961 = n45820 | n45821;
  assign n45823 = ~pi282 & n44153;
  assign n45824 = ~pi270 & n45823;
  assign n45825 = pi270 & ~n45823;
  assign po962 = ~n45824 & ~n45825;
  assign n45827 = pi807 & ~n45789;
  assign n45828 = pi1127 & n45789;
  assign po964 = n45827 | n45828;
  assign n45830 = pi808 & ~n45789;
  assign n45831 = pi1101 & n45789;
  assign po965 = n45830 | n45831;
  assign n45833 = pi809 & ~n45789;
  assign n45834 = ~pi1103 & n45789;
  assign po966 = ~n45833 & ~n45834;
  assign n45836 = pi810 & ~n45789;
  assign n45837 = pi1108 & n45789;
  assign po967 = n45836 | n45837;
  assign n45839 = pi811 & ~n45789;
  assign n45840 = pi1102 & n45789;
  assign po968 = n45839 | n45840;
  assign n45842 = pi812 & ~n45789;
  assign n45843 = ~pi1104 & n45789;
  assign po969 = ~n45842 & ~n45843;
  assign n45845 = pi813 & ~n45789;
  assign n45846 = pi1131 & n45789;
  assign po970 = n45845 | n45846;
  assign n45848 = pi814 & ~n45789;
  assign n45849 = ~pi1105 & n45789;
  assign po971 = ~n45848 & ~n45849;
  assign n45851 = pi815 & ~n45789;
  assign n45852 = pi1110 & n45789;
  assign po972 = n45851 | n45852;
  assign n45854 = pi816 & ~n45789;
  assign n45855 = pi1129 & n45789;
  assign po973 = n45854 | n45855;
  assign n45857 = pi269 & ~n44151;
  assign po974 = ~n44152 & ~n45857;
  assign n45859 = n7578 & n13384;
  assign po975 = n13261 | n45859;
  assign n45861 = pi265 & ~n44157;
  assign po976 = ~n44158 & ~n45861;
  assign n45863 = pi277 & ~n45824;
  assign po977 = ~n44156 & ~n45863;
  assign po979 = ~pi811 & ~pi893;
  assign n45866 = ~pi982 & ~n6179;
  assign n45867 = n7561 & n7578;
  assign n45868 = ~n45866 & ~n45867;
  assign po981 = n6102 & ~n45868;
  assign n45870 = pi123 & n2609;
  assign n45871 = pi1131 & ~n45870;
  assign n45872 = pi1127 & ~n45870;
  assign n45873 = ~n45871 & ~n45872;
  assign n45874 = ~pi825 & n45870;
  assign n45875 = n45873 & ~n45874;
  assign n45876 = pi1131 & n45872;
  assign n45877 = ~n45875 & ~n45876;
  assign n45878 = pi1128 & ~pi1129;
  assign n45879 = ~pi1128 & pi1129;
  assign n45880 = ~n45878 & ~n45879;
  assign n45881 = ~pi1124 & ~pi1130;
  assign n45882 = pi1124 & pi1130;
  assign n45883 = ~n45881 & ~n45882;
  assign n45884 = ~pi1125 & ~pi1126;
  assign n45885 = pi1125 & pi1126;
  assign n45886 = ~n45884 & ~n45885;
  assign n45887 = n45883 & ~n45886;
  assign n45888 = ~n45883 & n45886;
  assign n45889 = ~n45887 & ~n45888;
  assign n45890 = n45880 & n45889;
  assign n45891 = ~n45880 & ~n45889;
  assign n45892 = ~n45890 & ~n45891;
  assign n45893 = ~n45877 & ~n45892;
  assign n45894 = pi825 & n45870;
  assign n45895 = n45873 & ~n45894;
  assign n45896 = ~n45876 & n45892;
  assign n45897 = ~n45895 & n45896;
  assign po982 = ~n45893 & ~n45897;
  assign n45899 = pi1123 & ~n45870;
  assign n45900 = pi1122 & ~n45870;
  assign n45901 = ~n45899 & ~n45900;
  assign n45902 = ~pi826 & n45870;
  assign n45903 = n45901 & ~n45902;
  assign n45904 = pi1123 & n45900;
  assign n45905 = ~n45903 & ~n45904;
  assign n45906 = pi1120 & ~pi1121;
  assign n45907 = ~pi1120 & pi1121;
  assign n45908 = ~n45906 & ~n45907;
  assign n45909 = ~pi1118 & ~pi1119;
  assign n45910 = pi1118 & pi1119;
  assign n45911 = ~n45909 & ~n45910;
  assign n45912 = ~pi1116 & ~pi1117;
  assign n45913 = pi1116 & pi1117;
  assign n45914 = ~n45912 & ~n45913;
  assign n45915 = n45911 & ~n45914;
  assign n45916 = ~n45911 & n45914;
  assign n45917 = ~n45915 & ~n45916;
  assign n45918 = n45908 & n45917;
  assign n45919 = ~n45908 & ~n45917;
  assign n45920 = ~n45918 & ~n45919;
  assign n45921 = ~n45905 & ~n45920;
  assign n45922 = pi826 & n45870;
  assign n45923 = n45901 & ~n45922;
  assign n45924 = ~n45904 & n45920;
  assign n45925 = ~n45923 & n45924;
  assign po983 = ~n45921 & ~n45925;
  assign n45927 = pi1100 & ~n45870;
  assign n45928 = pi1107 & ~n45870;
  assign n45929 = ~n45927 & ~n45928;
  assign n45930 = ~pi827 & n45870;
  assign n45931 = n45929 & ~n45930;
  assign n45932 = pi1100 & n45928;
  assign n45933 = ~n45931 & ~n45932;
  assign n45934 = pi1101 & ~pi1102;
  assign n45935 = ~pi1101 & pi1102;
  assign n45936 = ~n45934 & ~n45935;
  assign n45937 = ~pi1103 & ~pi1105;
  assign n45938 = pi1103 & pi1105;
  assign n45939 = ~n45937 & ~n45938;
  assign n45940 = ~pi1104 & ~pi1106;
  assign n45941 = pi1104 & pi1106;
  assign n45942 = ~n45940 & ~n45941;
  assign n45943 = n45939 & ~n45942;
  assign n45944 = ~n45939 & n45942;
  assign n45945 = ~n45943 & ~n45944;
  assign n45946 = n45936 & n45945;
  assign n45947 = ~n45936 & ~n45945;
  assign n45948 = ~n45946 & ~n45947;
  assign n45949 = ~n45933 & ~n45948;
  assign n45950 = pi827 & n45870;
  assign n45951 = n45929 & ~n45950;
  assign n45952 = ~n45932 & n45948;
  assign n45953 = ~n45951 & n45952;
  assign po984 = ~n45949 & ~n45953;
  assign n45955 = pi1115 & ~n45870;
  assign n45956 = pi1114 & ~n45870;
  assign n45957 = ~n45955 & ~n45956;
  assign n45958 = ~pi828 & n45870;
  assign n45959 = n45957 & ~n45958;
  assign n45960 = pi1115 & n45956;
  assign n45961 = ~n45959 & ~n45960;
  assign n45962 = pi1112 & ~pi1113;
  assign n45963 = ~pi1112 & pi1113;
  assign n45964 = ~n45962 & ~n45963;
  assign n45965 = ~pi1110 & ~pi1111;
  assign n45966 = pi1110 & pi1111;
  assign n45967 = ~n45965 & ~n45966;
  assign n45968 = ~pi1108 & ~pi1109;
  assign n45969 = pi1108 & pi1109;
  assign n45970 = ~n45968 & ~n45969;
  assign n45971 = n45967 & ~n45970;
  assign n45972 = ~n45967 & n45970;
  assign n45973 = ~n45971 & ~n45972;
  assign n45974 = n45964 & n45973;
  assign n45975 = ~n45964 & ~n45973;
  assign n45976 = ~n45974 & ~n45975;
  assign n45977 = ~n45961 & ~n45976;
  assign n45978 = pi828 & n45870;
  assign n45979 = n45957 & ~n45978;
  assign n45980 = ~n45960 & n45976;
  assign n45981 = ~n45979 & n45980;
  assign po985 = ~n45977 & ~n45981;
  assign n45983 = n6178 & n7578;
  assign n45984 = pi951 & ~n45983;
  assign po986 = pi1092 & ~n45984;
  assign n45986 = pi281 & ~n45799;
  assign po987 = ~n45800 & ~n45986;
  assign n45988 = ~pi832 & pi1091;
  assign n45989 = pi1162 & n45988;
  assign po989 = n8593 & n45989;
  assign n45991 = pi1092 & n6178;
  assign n45992 = pi833 & ~n2923;
  assign po990 = n45991 | n45992;
  assign po991 = pi946 & n2923;
  assign n45995 = pi282 & ~n44153;
  assign po992 = ~n45823 & ~n45995;
  assign n45997 = ~pi837 & pi955;
  assign n45998 = ~pi955 & ~pi1049;
  assign po993 = ~n45997 & ~n45998;
  assign n46000 = ~pi838 & pi955;
  assign n46001 = ~pi955 & ~pi1047;
  assign po994 = ~n46000 & ~n46001;
  assign n46003 = ~pi839 & pi955;
  assign n46004 = ~pi955 & ~pi1074;
  assign po995 = ~n46003 & ~n46004;
  assign n46006 = pi840 & ~n2923;
  assign n46007 = pi1196 & n2923;
  assign po996 = n46006 | n46007;
  assign po997 = ~pi33 & n8684;
  assign n46010 = ~pi842 & pi955;
  assign n46011 = ~pi955 & ~pi1035;
  assign po998 = ~n46010 & ~n46011;
  assign n46013 = ~pi843 & pi955;
  assign n46014 = ~pi955 & ~pi1079;
  assign po999 = ~n46013 & ~n46014;
  assign n46016 = ~pi844 & pi955;
  assign n46017 = ~pi955 & ~pi1078;
  assign po1000 = ~n46016 & ~n46017;
  assign n46019 = ~pi845 & pi955;
  assign n46020 = ~pi955 & ~pi1043;
  assign po1001 = ~n46019 & ~n46020;
  assign n46022 = pi1134 & ~n40469;
  assign n46023 = pi846 & n40469;
  assign po1002 = n46022 | n46023;
  assign n46025 = ~pi847 & pi955;
  assign n46026 = ~pi955 & ~pi1055;
  assign po1003 = ~n46025 & ~n46026;
  assign n46028 = ~pi848 & pi955;
  assign n46029 = ~pi955 & ~pi1039;
  assign po1004 = ~n46028 & ~n46029;
  assign n46031 = pi849 & ~n2923;
  assign n46032 = pi1198 & n2923;
  assign po1005 = n46031 | n46032;
  assign n46034 = ~pi850 & pi955;
  assign n46035 = ~pi955 & ~pi1048;
  assign po1006 = ~n46034 & ~n46035;
  assign n46037 = ~pi851 & pi955;
  assign n46038 = ~pi955 & ~pi1045;
  assign po1007 = ~n46037 & ~n46038;
  assign n46040 = ~pi852 & pi955;
  assign n46041 = ~pi955 & ~pi1062;
  assign po1008 = ~n46040 & ~n46041;
  assign n46043 = ~pi853 & pi955;
  assign n46044 = ~pi955 & ~pi1080;
  assign po1009 = ~n46043 & ~n46044;
  assign n46046 = ~pi854 & pi955;
  assign n46047 = ~pi955 & ~pi1051;
  assign po1010 = ~n46046 & ~n46047;
  assign n46049 = ~pi855 & pi955;
  assign n46050 = ~pi955 & ~pi1065;
  assign po1011 = ~n46049 & ~n46050;
  assign n46052 = ~pi856 & pi955;
  assign n46053 = ~pi955 & ~pi1067;
  assign po1012 = ~n46052 & ~n46053;
  assign n46055 = ~pi857 & pi955;
  assign n46056 = ~pi955 & ~pi1058;
  assign po1013 = ~n46055 & ~n46056;
  assign n46058 = ~pi858 & pi955;
  assign n46059 = ~pi955 & ~pi1087;
  assign po1014 = ~n46058 & ~n46059;
  assign n46061 = ~pi859 & pi955;
  assign n46062 = ~pi955 & ~pi1070;
  assign po1015 = ~n46061 & ~n46062;
  assign n46064 = ~pi860 & pi955;
  assign n46065 = ~pi955 & ~pi1076;
  assign po1016 = ~n46064 & ~n46065;
  assign n46067 = pi1093 & pi1141;
  assign n46068 = pi861 & ~pi1093;
  assign n46069 = ~n46067 & ~n46068;
  assign n46070 = ~pi228 & ~n46069;
  assign n46071 = ~pi123 & ~pi1141;
  assign n46072 = pi123 & ~pi861;
  assign n46073 = pi228 & ~n46071;
  assign n46074 = ~n46072 & n46073;
  assign po1017 = n46070 | n46074;
  assign n46076 = pi1139 & ~n40469;
  assign n46077 = pi862 & n40469;
  assign po1018 = n46076 | n46077;
  assign n46079 = pi863 & ~n2923;
  assign n46080 = pi1199 & n2923;
  assign po1019 = n46079 | n46080;
  assign n46082 = pi864 & ~n2923;
  assign n46083 = pi1197 & n2923;
  assign po1020 = n46082 | n46083;
  assign n46085 = ~pi865 & pi955;
  assign n46086 = ~pi955 & ~pi1040;
  assign po1021 = ~n46085 & ~n46086;
  assign n46088 = ~pi866 & pi955;
  assign n46089 = ~pi955 & ~pi1053;
  assign po1022 = ~n46088 & ~n46089;
  assign n46091 = ~pi867 & pi955;
  assign n46092 = ~pi955 & ~pi1057;
  assign po1023 = ~n46091 & ~n46092;
  assign n46094 = ~pi868 & pi955;
  assign n46095 = ~pi955 & ~pi1063;
  assign po1024 = ~n46094 & ~n46095;
  assign n46097 = pi1093 & pi1140;
  assign n46098 = pi869 & ~pi1093;
  assign n46099 = ~n46097 & ~n46098;
  assign n46100 = ~pi228 & ~n46099;
  assign n46101 = ~pi123 & ~pi1140;
  assign n46102 = pi123 & ~pi869;
  assign n46103 = pi228 & ~n46101;
  assign n46104 = ~n46102 & n46103;
  assign po1025 = n46100 | n46104;
  assign n46106 = ~pi870 & pi955;
  assign n46107 = ~pi955 & ~pi1069;
  assign po1026 = ~n46106 & ~n46107;
  assign n46109 = ~pi871 & pi955;
  assign n46110 = ~pi955 & ~pi1072;
  assign po1027 = ~n46109 & ~n46110;
  assign n46112 = ~pi872 & pi955;
  assign n46113 = ~pi955 & ~pi1084;
  assign po1028 = ~n46112 & ~n46113;
  assign n46115 = ~pi873 & pi955;
  assign n46116 = ~pi955 & ~pi1044;
  assign po1029 = ~n46115 & ~n46116;
  assign n46118 = ~pi874 & pi955;
  assign n46119 = ~pi955 & ~pi1036;
  assign po1030 = ~n46118 & ~n46119;
  assign n46121 = pi1093 & ~pi1136;
  assign n46122 = ~pi875 & ~pi1093;
  assign n46123 = ~n46121 & ~n46122;
  assign n46124 = ~pi228 & ~n46123;
  assign n46125 = ~pi123 & pi1136;
  assign n46126 = pi123 & pi875;
  assign n46127 = pi228 & ~n46125;
  assign n46128 = ~n46126 & n46127;
  assign po1031 = ~n46124 & ~n46128;
  assign n46130 = ~pi876 & pi955;
  assign n46131 = ~pi955 & ~pi1037;
  assign po1032 = ~n46130 & ~n46131;
  assign n46133 = pi1093 & pi1138;
  assign n46134 = pi877 & ~pi1093;
  assign n46135 = ~n46133 & ~n46134;
  assign n46136 = ~pi228 & ~n46135;
  assign n46137 = ~pi123 & ~pi1138;
  assign n46138 = pi123 & ~pi877;
  assign n46139 = pi228 & ~n46137;
  assign n46140 = ~n46138 & n46139;
  assign po1033 = n46136 | n46140;
  assign n46142 = pi1093 & pi1137;
  assign n46143 = pi878 & ~pi1093;
  assign n46144 = ~n46142 & ~n46143;
  assign n46145 = ~pi228 & ~n46144;
  assign n46146 = ~pi123 & ~pi1137;
  assign n46147 = pi123 & ~pi878;
  assign n46148 = pi228 & ~n46146;
  assign n46149 = ~n46147 & n46148;
  assign po1034 = n46145 | n46149;
  assign n46151 = pi1093 & pi1135;
  assign n46152 = pi879 & ~pi1093;
  assign n46153 = ~n46151 & ~n46152;
  assign n46154 = ~pi228 & ~n46153;
  assign n46155 = ~pi123 & ~pi1135;
  assign n46156 = pi123 & ~pi879;
  assign n46157 = pi228 & ~n46155;
  assign n46158 = ~n46156 & n46157;
  assign po1035 = n46154 | n46158;
  assign n46160 = ~pi880 & pi955;
  assign n46161 = ~pi955 & ~pi1081;
  assign po1036 = ~n46160 & ~n46161;
  assign n46163 = ~pi881 & pi955;
  assign n46164 = ~pi955 & ~pi1059;
  assign po1037 = ~n46163 & ~n46164;
  assign n46166 = ~pi883 & n45870;
  assign po1039 = n45928 | n46166;
  assign n46168 = pi1124 & ~n45870;
  assign n46169 = ~pi884 & n45870;
  assign po1040 = n46168 | n46169;
  assign n46171 = pi1125 & ~n45870;
  assign n46172 = ~pi885 & n45870;
  assign po1041 = n46171 | n46172;
  assign n46174 = pi1109 & ~n45870;
  assign n46175 = ~pi886 & n45870;
  assign po1042 = n46174 | n46175;
  assign n46177 = ~pi887 & n45870;
  assign po1043 = n45927 | n46177;
  assign n46179 = pi1120 & ~n45870;
  assign n46180 = ~pi888 & n45870;
  assign po1044 = n46179 | n46180;
  assign n46182 = pi1103 & ~n45870;
  assign n46183 = ~pi889 & n45870;
  assign po1045 = n46182 | n46183;
  assign n46185 = pi1126 & ~n45870;
  assign n46186 = ~pi890 & n45870;
  assign po1046 = n46185 | n46186;
  assign n46188 = pi1116 & ~n45870;
  assign n46189 = ~pi891 & n45870;
  assign po1047 = n46188 | n46189;
  assign n46191 = pi1101 & ~n45870;
  assign n46192 = ~pi892 & n45870;
  assign po1048 = n46191 | n46192;
  assign n46194 = pi1119 & ~n45870;
  assign n46195 = ~pi894 & n45870;
  assign po1050 = n46194 | n46195;
  assign n46197 = pi1113 & ~n45870;
  assign n46198 = ~pi895 & n45870;
  assign po1051 = n46197 | n46198;
  assign n46200 = pi1118 & ~n45870;
  assign n46201 = ~pi896 & n45870;
  assign po1052 = n46200 | n46201;
  assign n46203 = pi1129 & ~n45870;
  assign n46204 = ~pi898 & n45870;
  assign po1054 = n46203 | n46204;
  assign n46206 = ~pi899 & n45870;
  assign po1055 = n45955 | n46206;
  assign n46208 = pi1110 & ~n45870;
  assign n46209 = ~pi900 & n45870;
  assign po1056 = n46208 | n46209;
  assign n46211 = pi1111 & ~n45870;
  assign n46212 = ~pi902 & n45870;
  assign po1058 = n46211 | n46212;
  assign n46214 = pi1121 & ~n45870;
  assign n46215 = ~pi903 & n45870;
  assign po1059 = n46214 | n46215;
  assign n46217 = ~pi904 & n45870;
  assign po1060 = n45872 | n46217;
  assign n46219 = ~pi905 & n45870;
  assign po1061 = n45871 | n46219;
  assign n46221 = pi1128 & ~n45870;
  assign n46222 = ~pi906 & n45870;
  assign po1062 = n46221 | n46222;
  assign n46224 = ~pi782 & ~pi907;
  assign n46225 = ~pi624 & ~pi979;
  assign n46226 = ~pi598 & pi979;
  assign n46227 = pi782 & ~n46225;
  assign n46228 = ~n46226 & n46227;
  assign n46229 = ~pi604 & ~pi979;
  assign n46230 = pi615 & pi979;
  assign n46231 = ~n46229 & ~n46230;
  assign n46232 = pi782 & ~n46231;
  assign n46233 = ~n46224 & ~n46228;
  assign po1063 = ~n46232 & n46233;
  assign n46235 = ~pi908 & n45870;
  assign po1064 = n45900 | n46235;
  assign n46237 = pi1105 & ~n45870;
  assign n46238 = ~pi909 & n45870;
  assign po1065 = n46237 | n46238;
  assign n46240 = pi1117 & ~n45870;
  assign n46241 = ~pi910 & n45870;
  assign po1066 = n46240 | n46241;
  assign n46243 = pi1130 & ~n45870;
  assign n46244 = ~pi911 & n45870;
  assign po1067 = n46243 | n46244;
  assign n46246 = ~pi912 & n45870;
  assign po1068 = n45956 | n46246;
  assign n46248 = pi1106 & ~n45870;
  assign n46249 = ~pi913 & n45870;
  assign po1069 = n46248 | n46249;
  assign n46251 = pi280 & ~n44150;
  assign po1070 = ~n44151 & ~n46251;
  assign n46253 = pi1108 & ~n45870;
  assign n46254 = ~pi915 & n45870;
  assign po1071 = n46253 | n46254;
  assign n46256 = ~pi916 & n45870;
  assign po1072 = n45899 | n46256;
  assign n46258 = pi1112 & ~n45870;
  assign n46259 = ~pi917 & n45870;
  assign po1073 = n46258 | n46259;
  assign n46261 = pi1104 & ~n45870;
  assign n46262 = ~pi918 & n45870;
  assign po1074 = n46261 | n46262;
  assign n46264 = pi1102 & ~n45870;
  assign n46265 = ~pi919 & n45870;
  assign po1075 = n46264 | n46265;
  assign n46267 = ~pi920 & ~pi1093;
  assign n46268 = pi1093 & ~pi1139;
  assign po1076 = ~n46267 & ~n46268;
  assign n46270 = pi921 & ~pi1093;
  assign po1077 = n46097 | n46270;
  assign n46272 = pi1093 & pi1152;
  assign n46273 = pi922 & ~pi1093;
  assign po1078 = n46272 | n46273;
  assign n46275 = pi1093 & pi1154;
  assign n46276 = pi923 & ~pi1093;
  assign po1079 = n46275 | n46276;
  assign n46278 = pi311 & ~pi312;
  assign po1080 = n42028 & n46278;
  assign n46280 = pi1093 & pi1155;
  assign n46281 = pi925 & ~pi1093;
  assign po1081 = n46280 | n46281;
  assign n46283 = pi1093 & pi1157;
  assign n46284 = pi926 & ~pi1093;
  assign po1082 = n46283 | n46284;
  assign n46286 = pi1093 & pi1145;
  assign n46287 = pi927 & ~pi1093;
  assign po1083 = n46286 | n46287;
  assign n46289 = ~pi928 & ~pi1093;
  assign po1084 = ~n46121 & ~n46289;
  assign n46291 = pi1093 & pi1144;
  assign n46292 = pi929 & ~pi1093;
  assign po1085 = n46291 | n46292;
  assign n46294 = pi1093 & pi1134;
  assign n46295 = pi930 & ~pi1093;
  assign po1086 = n46294 | n46295;
  assign n46297 = pi1093 & pi1150;
  assign n46298 = pi931 & ~pi1093;
  assign po1087 = n46297 | n46298;
  assign n46300 = pi932 & ~pi1093;
  assign po1088 = n40471 | n46300;
  assign n46302 = pi933 & ~pi1093;
  assign po1089 = n46142 | n46302;
  assign n46304 = pi1093 & pi1147;
  assign n46305 = pi934 & ~pi1093;
  assign po1090 = n46304 | n46305;
  assign n46307 = pi935 & ~pi1093;
  assign po1091 = n46067 | n46307;
  assign n46309 = pi1093 & pi1149;
  assign n46310 = pi936 & ~pi1093;
  assign po1092 = n46309 | n46310;
  assign n46312 = pi1093 & pi1148;
  assign n46313 = pi937 & ~pi1093;
  assign po1093 = n46312 | n46313;
  assign n46315 = pi938 & ~pi1093;
  assign po1094 = n46151 | n46315;
  assign n46317 = pi1093 & pi1146;
  assign n46318 = pi939 & ~pi1093;
  assign po1095 = n46317 | n46318;
  assign n46320 = pi940 & ~pi1093;
  assign po1096 = n46133 | n46320;
  assign n46322 = pi1093 & pi1153;
  assign n46323 = pi941 & ~pi1093;
  assign po1097 = n46322 | n46323;
  assign n46325 = pi1093 & pi1156;
  assign n46326 = pi942 & ~pi1093;
  assign po1098 = n46325 | n46326;
  assign n46328 = pi1093 & pi1151;
  assign n46329 = pi943 & ~pi1093;
  assign po1099 = n46328 | n46329;
  assign n46331 = ~pi944 & ~pi1093;
  assign n46332 = pi1093 & ~pi1143;
  assign po1100 = ~n46331 & ~n46332;
  assign po1102 = pi230 & n2923;
  assign n46335 = ~pi782 & pi947;
  assign po1103 = n46228 | n46335;
  assign n46337 = ~pi266 & ~pi992;
  assign po1104 = ~n44150 & ~n46337;
  assign n46339 = ~pi949 & pi954;
  assign n46340 = pi313 & ~pi954;
  assign po1105 = ~n46339 & ~n46340;
  assign po1106 = n2921 & n45991;
  assign po1107 = n7470 & ~n7561;
  assign n46344 = pi957 & pi1092;
  assign po1112 = pi31 | n46344;
  assign po1115 = ~pi782 & pi960;
  assign po1116 = ~pi230 & pi961;
  assign po1118 = ~pi782 & pi963;
  assign po1122 = ~pi230 & pi967;
  assign po1124 = ~pi230 & pi969;
  assign po1125 = ~pi782 & pi970;
  assign po1126 = ~pi230 & pi971;
  assign po1127 = ~pi782 & pi972;
  assign po1128 = ~pi230 & pi974;
  assign po1129 = ~pi782 & pi975;
  assign po1131 = ~pi230 & pi977;
  assign po1132 = ~pi782 & pi978;
  assign po1133 = pi598 | ~pi615;
  assign po1135 = pi824 & pi1092;
  assign po1137 = pi604 | pi624;
  assign po166 = 1'b1;
  assign po170 = ~pi1090;
  assign po1110 = ~pi954;
  assign po1130 = ~pi278;
  assign po1146 = ~pi915;
  assign po1147 = ~pi825;
  assign po1148 = ~pi826;
  assign po1149 = ~pi913;
  assign po1150 = ~pi894;
  assign po1151 = ~pi905;
  assign po1153 = ~pi890;
  assign po1155 = ~pi906;
  assign po1156 = ~pi896;
  assign po1157 = ~pi909;
  assign po1158 = ~pi911;
  assign po1159 = ~pi908;
  assign po1160 = ~pi891;
  assign po1161 = ~pi902;
  assign po1162 = ~pi903;
  assign po1163 = ~pi883;
  assign po1164 = ~pi888;
  assign po1165 = ~pi919;
  assign po1166 = ~pi886;
  assign po1167 = ~pi912;
  assign po1168 = ~pi895;
  assign po1169 = ~pi916;
  assign po1170 = ~pi889;
  assign po1171 = ~pi900;
  assign po1172 = ~pi885;
  assign po1173 = ~pi904;
  assign po1174 = ~pi899;
  assign po1175 = ~pi918;
  assign po1176 = ~pi898;
  assign po1177 = ~pi917;
  assign po1178 = ~pi827;
  assign po1179 = ~pi887;
  assign po1180 = ~pi884;
  assign po1181 = ~pi910;
  assign po1182 = ~pi828;
  assign po1183 = ~pi892;
  assign po0 = pi668;
  assign po1 = pi672;
  assign po2 = pi664;
  assign po3 = pi667;
  assign po4 = pi676;
  assign po5 = pi673;
  assign po6 = pi675;
  assign po7 = pi666;
  assign po8 = pi679;
  assign po9 = pi674;
  assign po10 = pi663;
  assign po11 = pi670;
  assign po12 = pi677;
  assign po13 = pi682;
  assign po14 = pi671;
  assign po15 = pi678;
  assign po16 = pi718;
  assign po17 = pi707;
  assign po18 = pi708;
  assign po19 = pi713;
  assign po20 = pi711;
  assign po21 = pi716;
  assign po22 = pi733;
  assign po23 = pi712;
  assign po24 = pi689;
  assign po25 = pi717;
  assign po26 = pi692;
  assign po27 = pi719;
  assign po28 = pi722;
  assign po29 = pi714;
  assign po30 = pi720;
  assign po31 = pi685;
  assign po32 = pi837;
  assign po33 = pi850;
  assign po34 = pi872;
  assign po35 = pi871;
  assign po36 = pi881;
  assign po37 = pi866;
  assign po38 = pi876;
  assign po39 = pi873;
  assign po40 = pi874;
  assign po41 = pi859;
  assign po42 = pi855;
  assign po43 = pi852;
  assign po44 = pi870;
  assign po45 = pi848;
  assign po46 = pi865;
  assign po47 = pi856;
  assign po48 = pi853;
  assign po49 = pi847;
  assign po50 = pi857;
  assign po51 = pi854;
  assign po52 = pi858;
  assign po53 = pi845;
  assign po54 = pi838;
  assign po55 = pi842;
  assign po56 = pi843;
  assign po57 = pi839;
  assign po58 = pi844;
  assign po59 = pi868;
  assign po60 = pi851;
  assign po61 = pi867;
  assign po62 = pi880;
  assign po63 = pi860;
  assign po64 = pi1030;
  assign po65 = pi1034;
  assign po66 = pi1015;
  assign po67 = pi1020;
  assign po68 = pi1025;
  assign po69 = pi1005;
  assign po70 = pi996;
  assign po71 = pi1012;
  assign po72 = pi993;
  assign po73 = pi1016;
  assign po74 = pi1021;
  assign po75 = pi1010;
  assign po76 = pi1027;
  assign po77 = pi1018;
  assign po78 = pi1017;
  assign po79 = pi1024;
  assign po80 = pi1009;
  assign po81 = pi1032;
  assign po82 = pi1003;
  assign po83 = pi997;
  assign po84 = pi1013;
  assign po85 = pi1011;
  assign po86 = pi1008;
  assign po87 = pi1019;
  assign po88 = pi1031;
  assign po89 = pi1022;
  assign po90 = pi1000;
  assign po91 = pi1023;
  assign po92 = pi1002;
  assign po93 = pi1026;
  assign po94 = pi1006;
  assign po95 = pi998;
  assign po96 = pi31;
  assign po97 = pi80;
  assign po98 = pi893;
  assign po99 = pi467;
  assign po100 = pi78;
  assign po101 = pi112;
  assign po102 = pi13;
  assign po103 = pi25;
  assign po104 = pi226;
  assign po105 = pi127;
  assign po106 = pi822;
  assign po107 = pi808;
  assign po108 = pi227;
  assign po109 = pi477;
  assign po110 = pi834;
  assign po111 = pi229;
  assign po112 = pi12;
  assign po113 = pi11;
  assign po114 = pi10;
  assign po115 = pi9;
  assign po116 = pi8;
  assign po117 = pi7;
  assign po118 = pi6;
  assign po119 = pi5;
  assign po120 = pi4;
  assign po121 = pi3;
  assign po122 = pi0;
  assign po123 = pi2;
  assign po124 = pi1;
  assign po125 = pi310;
  assign po126 = pi302;
  assign po127 = pi475;
  assign po128 = pi474;
  assign po129 = pi466;
  assign po130 = pi473;
  assign po131 = pi471;
  assign po132 = pi472;
  assign po133 = pi470;
  assign po134 = pi469;
  assign po135 = pi465;
  assign po136 = pi1028;
  assign po137 = pi1033;
  assign po138 = pi995;
  assign po139 = pi994;
  assign po140 = pi28;
  assign po141 = pi27;
  assign po142 = pi26;
  assign po143 = pi29;
  assign po144 = pi15;
  assign po145 = pi14;
  assign po146 = pi21;
  assign po147 = pi20;
  assign po148 = pi19;
  assign po149 = pi18;
  assign po150 = pi17;
  assign po151 = pi16;
  assign po152 = pi1096;
  assign po168 = pi228;
  assign po169 = pi22;
  assign po179 = pi1089;
  assign po180 = pi23;
  assign po181 = po167;
  assign po188 = pi37;
  assign po263 = pi117;
  assign po285 = pi131;
  assign po386 = pi232;
  assign po388 = pi236;
  assign po636 = pi583;
  assign po1053 = pi67;
  assign po1108 = pi1134;
  assign po1109 = pi964;
  assign po1111 = pi965;
  assign po1113 = pi991;
  assign po1114 = pi985;
  assign po1117 = pi1014;
  assign po1119 = pi1029;
  assign po1120 = pi1004;
  assign po1121 = pi1007;
  assign po1123 = pi1135;
  assign po1134 = pi1064;
  assign po1136 = pi299;
  assign po1138 = pi1075;
  assign po1139 = pi1052;
  assign po1140 = pi771;
  assign po1141 = pi765;
  assign po1142 = pi605;
  assign po1143 = pi601;
  assign po1144 = pi278;
  assign po1145 = pi279;
  assign po1152 = pi1095;
  assign po1154 = pi1094;
  assign po1184 = pi1187;
  assign po1185 = pi1172;
  assign po1186 = pi1170;
  assign po1187 = pi1138;
  assign po1188 = pi1177;
  assign po1189 = pi1178;
  assign po1190 = pi863;
  assign po1191 = pi1203;
  assign po1192 = pi1185;
  assign po1193 = pi1171;
  assign po1194 = pi1192;
  assign po1195 = pi1137;
  assign po1196 = pi1186;
  assign po1197 = pi1165;
  assign po1198 = pi1164;
  assign po1199 = pi1098;
  assign po1200 = pi1183;
  assign po1201 = pi230;
  assign po1202 = pi1169;
  assign po1203 = pi1136;
  assign po1204 = pi1181;
  assign po1205 = pi849;
  assign po1206 = pi1193;
  assign po1207 = pi1182;
  assign po1208 = pi1168;
  assign po1209 = pi1175;
  assign po1210 = pi1191;
  assign po1211 = pi1099;
  assign po1212 = pi1174;
  assign po1213 = pi1179;
  assign po1214 = pi1202;
  assign po1215 = pi1176;
  assign po1216 = pi1173;
  assign po1217 = pi1201;
  assign po1218 = pi1167;
  assign po1219 = pi840;
  assign po1220 = pi1189;
  assign po1221 = pi1195;
  assign po1222 = pi864;
  assign po1223 = pi1190;
  assign po1224 = pi1188;
  assign po1225 = pi1180;
  assign po1226 = pi1194;
  assign po1227 = pi1097;
  assign po1228 = pi1166;
  assign po1229 = pi1200;
  assign po1230 = pi1184;
endmodule
