module alu4_cl ( 
    pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09, pi10, pi11,
    pi12, pi13,
    po0, po1, po2, po3, po4, po5, po6, po7  );
  input  pi00, pi01, pi02, pi03, pi04, pi05, pi06, pi07, pi08, pi09,
    pi10, pi11, pi12, pi13;
  output po0, po1, po2, po3, po4, po5, po6, po7;
  wire n23, n24, n25, n26, n27, n28, n29,
    n30, n31, n32, n33, n34, n35, n36, n37,
    n38, n39, n40, n41, n42, n43, n44, n45,
    n46, n47, n48, n49, n50, n51, n52, n53,
    n54, n55, n56, n57, n58, n59, n60, n61,
    n62, n63, n64, n65, n66, n67, n68, n69,
    n70, n71, n72, n73, n74, n75, n76, n77,
    n78, n79, n80, n81, n82, n83, n84, n85,
    n86, n87, n88, n89, n90, n91, n92, n93,
    n94, n95, n96, n97, n98, n99, n100,
    n101, n102, n103, n104, n105, n106, n107,
    n108, n109, n110, n111, n112, n113, n114,
    n115, n116, n117, n118, n119, n120, n121,
    n122, n123, n124, n125, n126, n127, n128,
    n129, n130, n131, n132, n133, n134, n135,
    n136, n137, n138, n139, n140, n141, n142,
    n143, n144, n145, n146, n147, n148, n149,
    n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163,
    n164, n165, n166, n167, n168, n169, n170,
    n171, n172, n173, n174, n175, n176, n177,
    n178, n179, n180, n182, n183, n184, n185,
    n186, n187, n188, n189, n190, n191, n192,
    n193, n194, n195, n196, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n215, n216, n217, n218, n219, n220,
    n221, n222, n223, n224, n225, n226, n227,
    n228, n229, n230, n231, n232, n233, n234,
    n235, n236, n237, n238, n239, n240, n241,
    n242, n243, n244, n245, n246, n247, n248,
    n249, n250, n251, n252, n253, n254, n255,
    n256, n257, n258, n259, n260, n261, n262,
    n263, n264, n265, n266, n267, n268, n269,
    n270, n271, n272, n273, n274, n275, n276,
    n277, n278, n279, n280, n281, n282, n283,
    n284, n285, n286, n287, n288, n289, n290,
    n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n332, n333,
    n334, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n372, n373, n374, n375,
    n376, n377, n378, n379, n380, n381, n382,
    n383, n384, n385, n386, n387, n388, n389,
    n390, n391, n392, n393, n394, n395, n396,
    n397, n398, n399, n400, n401, n402, n403,
    n404, n405, n406, n407, n408, n409, n410,
    n411, n412, n413, n414, n415, n416, n417,
    n418, n419, n420, n421, n422, n423, n424,
    n425, n426, n427, n428, n429, n430, n431,
    n432, n433, n434, n435, n436, n437, n438,
    n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n448, n449, n450, n451, n452,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n464, n465, n466,
    n467, n468, n469, n470, n471, n472, n473,
    n474, n475, n476, n477, n478, n479, n480,
    n481, n482, n483, n485, n486, n488, n489,
    n490, n491, n492, n493, n494, n495, n496,
    n497, n498, n499, n500, n501, n502, n503,
    n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517,
    n518, n519, n520, n521, n522, n523, n524,
    n525, n526, n527, n528, n529, n530, n531,
    n532, n533, n534, n535, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n545,
    n546, n547, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566,
    n567, n568, n569, n570, n571, n572, n573,
    n574, n575, n576, n577, n578, n579, n580,
    n581, n582, n583, n584, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n600, n601,
    n602, n603, n604, n605, n606, n607, n608,
    n609, n610, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n629,
    n630, n631, n632, n633, n634, n635, n636,
    n637, n638, n639, n640, n641, n644, n645,
    n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659,
    n660, n661, n662, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n672, n673,
    n674, n675, n677, n678;
  assign n23 = pi00 & pi11;
  assign n24 = ~pi08 & ~pi09;
  assign n25 = ~pi10 & ~n24;
  assign n26 = n23 & ~n25;
  assign n27 = ~pi00 & pi04;
  assign n28 = pi08 & ~pi10;
  assign n29 = pi11 & n28;
  assign n30 = n27 & n29;
  assign n31 = ~pi08 & pi10;
  assign n32 = ~pi10 & ~pi11;
  assign n33 = pi08 & n32;
  assign n34 = ~n31 & ~n33;
  assign n35 = pi09 & pi11;
  assign n36 = ~pi10 & ~pi13;
  assign n37 = ~n35 & n36;
  assign n38 = ~pi08 & n37;
  assign n39 = ~pi00 & n38;
  assign n40 = ~pi00 & ~pi04;
  assign n41 = ~pi10 & pi13;
  assign n42 = pi08 & ~pi09;
  assign n43 = ~pi13 & ~n32;
  assign n44 = ~n41 & n42;
  assign n45 = ~n43 & n44;
  assign n46 = ~n40 & n45;
  assign n47 = ~pi09 & pi11;
  assign n48 = pi08 & pi10;
  assign n49 = ~pi13 & n47;
  assign n50 = n48 & n49;
  assign n51 = pi10 & ~pi11;
  assign n52 = ~pi08 & pi09;
  assign n53 = pi13 & n52;
  assign n54 = ~n51 & n53;
  assign n55 = pi08 & pi09;
  assign n56 = n51 & n55;
  assign n57 = ~n50 & ~n56;
  assign n58 = ~n54 & n57;
  assign n59 = ~pi04 & ~n58;
  assign n60 = ~n24 & ~n55;
  assign n61 = ~pi10 & pi11;
  assign n62 = ~n60 & n61;
  assign n63 = pi13 & n62;
  assign n64 = ~pi09 & ~pi11;
  assign n65 = n31 & n64;
  assign n66 = ~n63 & ~n65;
  assign n67 = pi00 & pi04;
  assign n68 = ~n66 & n67;
  assign n69 = ~n40 & ~n67;
  assign n70 = ~pi00 & ~n51;
  assign n71 = n53 & n69;
  assign n72 = ~n70 & n71;
  assign n73 = ~n46 & ~n72;
  assign n74 = ~n59 & n73;
  assign n75 = ~n68 & n74;
  assign n76 = ~n39 & n75;
  assign n77 = ~n34 & n76;
  assign n78 = pi08 & n51;
  assign n79 = ~n23 & ~n78;
  assign n80 = ~pi04 & ~n79;
  assign n81 = ~n30 & ~n80;
  assign n82 = ~n77 & n81;
  assign n83 = ~pi09 & ~n82;
  assign n84 = ~pi08 & n51;
  assign n85 = n40 & n84;
  assign n86 = pi00 & ~n75;
  assign n87 = n48 & n86;
  assign n88 = ~pi11 & ~n31;
  assign n89 = ~pi08 & pi11;
  assign n90 = ~pi00 & ~n89;
  assign n91 = pi04 & ~n88;
  assign n92 = ~n90 & n91;
  assign n93 = ~n85 & ~n92;
  assign n94 = ~n87 & n93;
  assign n95 = pi09 & ~n94;
  assign n96 = ~pi08 & ~pi10;
  assign n97 = pi04 & n96;
  assign n98 = ~pi09 & ~n28;
  assign n99 = ~n51 & n98;
  assign n100 = ~n97 & ~n99;
  assign n101 = ~n76 & ~n100;
  assign n102 = ~n26 & ~n101;
  assign n103 = ~n83 & n102;
  assign n104 = ~n95 & n103;
  assign n105 = ~pi13 & ~n104;
  assign n106 = pi09 & pi13;
  assign n107 = n33 & n106;
  assign n108 = ~pi09 & pi10;
  assign n109 = ~pi13 & n89;
  assign n110 = n108 & n109;
  assign n111 = ~n107 & ~n110;
  assign n112 = pi10 & n55;
  assign n113 = ~pi00 & pi11;
  assign n114 = n112 & n113;
  assign n115 = n55 & n61;
  assign n116 = n51 & n52;
  assign n117 = ~n115 & ~n116;
  assign n118 = n23 & ~n55;
  assign n119 = ~pi08 & pi13;
  assign n120 = n35 & n119;
  assign n121 = ~pi10 & n120;
  assign n122 = n67 & n121;
  assign n123 = ~pi00 & n76;
  assign n124 = n120 & ~n123;
  assign n125 = pi13 & n51;
  assign n126 = n24 & n76;
  assign n127 = n55 & n86;
  assign n128 = n42 & n67;
  assign n129 = ~n126 & ~n128;
  assign n130 = ~n127 & n129;
  assign n131 = n125 & ~n130;
  assign n132 = ~n124 & ~n131;
  assign n133 = n42 & n125;
  assign n134 = n132 & n133;
  assign n135 = ~n122 & ~n134;
  assign n136 = pi08 & n64;
  assign n137 = ~n135 & n136;
  assign n138 = ~n118 & ~n137;
  assign n139 = pi10 & ~n138;
  assign n140 = n117 & ~n139;
  assign n141 = n76 & ~n140;
  assign n142 = n52 & n61;
  assign n143 = ~n135 & n142;
  assign n144 = ~n56 & ~n143;
  assign n145 = n132 & ~n144;
  assign n146 = n135 & n142;
  assign n147 = ~pi00 & n65;
  assign n148 = ~n146 & ~n147;
  assign n149 = ~n132 & ~n148;
  assign n150 = n42 & n51;
  assign n151 = n135 & n150;
  assign n152 = ~n25 & n113;
  assign n153 = ~n151 & ~n152;
  assign n154 = ~n76 & ~n153;
  assign n155 = pi04 & n28;
  assign n156 = pi00 & ~pi08;
  assign n157 = n132 & n156;
  assign n158 = ~n155 & ~n157;
  assign n159 = n64 & ~n158;
  assign n160 = ~pi09 & n28;
  assign n161 = n69 & n160;
  assign n162 = pi09 & ~n76;
  assign n163 = ~pi00 & ~n162;
  assign n164 = ~pi09 & n76;
  assign n165 = pi11 & ~n164;
  assign n166 = n96 & ~n163;
  assign n167 = ~n165 & n166;
  assign n168 = ~n114 & ~n161;
  assign n169 = ~n167 & n168;
  assign n170 = ~n159 & n169;
  assign n171 = ~n145 & n170;
  assign n172 = ~n149 & ~n154;
  assign n173 = n171 & n172;
  assign n174 = ~n141 & n173;
  assign n175 = ~pi12 & pi13;
  assign n176 = ~n174 & n175;
  assign n177 = pi12 & n174;
  assign n178 = pi13 & ~n176;
  assign n179 = ~n177 & n178;
  assign n180 = ~n105 & n111;
  assign po0 = n179 | ~n180;
  assign n182 = ~pi01 & pi05;
  assign n183 = n29 & n182;
  assign n184 = pi01 & pi05;
  assign n185 = ~pi09 & n51;
  assign n186 = pi13 & n185;
  assign n187 = n66 & ~n186;
  assign n188 = ~pi08 & n27;
  assign n189 = n125 & n188;
  assign n190 = n187 & ~n189;
  assign n191 = n184 & ~n190;
  assign n192 = n23 & n108;
  assign n193 = ~pi01 & ~pi05;
  assign n194 = n27 & n193;
  assign n195 = ~pi01 & ~n51;
  assign n196 = ~n184 & ~n193;
  assign n197 = ~n27 & ~n195;
  assign n198 = n196 & n197;
  assign n199 = ~n194 & ~n198;
  assign n200 = pi09 & ~n199;
  assign n201 = ~n192 & ~n200;
  assign n202 = n119 & ~n201;
  assign n203 = n45 & ~n193;
  assign n204 = ~pi01 & n38;
  assign n205 = ~pi05 & ~n58;
  assign n206 = ~n203 & ~n204;
  assign n207 = ~n205 & n206;
  assign n208 = ~n202 & n207;
  assign n209 = ~n191 & n208;
  assign n210 = ~n34 & n209;
  assign n211 = pi01 & pi11;
  assign n212 = ~n78 & ~n211;
  assign n213 = ~pi05 & ~n212;
  assign n214 = ~n183 & ~n213;
  assign n215 = ~n210 & n214;
  assign n216 = ~pi09 & ~n215;
  assign n217 = pi11 & ~n25;
  assign n218 = pi09 & ~n209;
  assign n219 = n48 & n218;
  assign n220 = ~n217 & ~n219;
  assign n221 = pi01 & ~n220;
  assign n222 = pi05 & n96;
  assign n223 = ~n99 & ~n222;
  assign n224 = ~n209 & ~n223;
  assign n225 = n84 & n193;
  assign n226 = pi01 & ~n88;
  assign n227 = ~n89 & ~n226;
  assign n228 = pi05 & ~n227;
  assign n229 = ~n225 & ~n228;
  assign n230 = pi09 & ~n229;
  assign n231 = ~n224 & ~n230;
  assign n232 = ~n216 & n231;
  assign n233 = ~n221 & n232;
  assign n234 = ~pi13 & ~n233;
  assign n235 = pi05 & n28;
  assign n236 = ~n76 & ~n135;
  assign n237 = n121 & n184;
  assign n238 = ~pi01 & n208;
  assign n239 = n120 & ~n238;
  assign n240 = n24 & n209;
  assign n241 = pi05 & ~pi09;
  assign n242 = ~n218 & ~n241;
  assign n243 = pi01 & pi08;
  assign n244 = ~n242 & n243;
  assign n245 = ~n240 & ~n244;
  assign n246 = n125 & ~n245;
  assign n247 = ~n239 & ~n246;
  assign n248 = n133 & n247;
  assign n249 = ~n237 & ~n248;
  assign n250 = n236 & ~n249;
  assign n251 = ~n236 & n249;
  assign n252 = ~n250 & ~n251;
  assign n253 = n209 & ~n252;
  assign n254 = ~n209 & n252;
  assign n255 = n48 & ~n253;
  assign n256 = ~n254 & n255;
  assign n257 = pi00 & ~n132;
  assign n258 = n247 & ~n257;
  assign n259 = ~n132 & ~n247;
  assign n260 = pi00 & n259;
  assign n261 = ~n258 & ~n260;
  assign n262 = pi01 & ~pi08;
  assign n263 = ~n261 & n262;
  assign n264 = ~n235 & ~n263;
  assign n265 = ~n256 & n264;
  assign n266 = n64 & ~n265;
  assign n267 = n132 & n247;
  assign n268 = ~n259 & ~n267;
  assign n269 = n112 & ~n268;
  assign n270 = pi09 & n96;
  assign n271 = ~n209 & n270;
  assign n272 = ~n269 & ~n271;
  assign n273 = ~pi11 & ~n272;
  assign n274 = pi10 & ~n55;
  assign n275 = ~n24 & ~n274;
  assign n276 = pi11 & ~n275;
  assign n277 = n86 & ~n209;
  assign n278 = ~n86 & n209;
  assign n279 = ~n277 & ~n278;
  assign n280 = n276 & n279;
  assign n281 = n65 & n261;
  assign n282 = ~n280 & ~n281;
  assign n283 = ~pi01 & ~n282;
  assign n284 = ~pi05 & ~n67;
  assign n285 = n160 & n284;
  assign n286 = ~n51 & ~n275;
  assign n287 = ~n279 & n286;
  assign n288 = n23 & n112;
  assign n289 = n32 & ~n55;
  assign n290 = ~n285 & ~n289;
  assign n291 = ~n288 & n290;
  assign n292 = ~n287 & n291;
  assign n293 = pi01 & ~n292;
  assign n294 = ~pi11 & n52;
  assign n295 = ~n115 & ~n294;
  assign n296 = ~n76 & ~n295;
  assign n297 = ~n209 & n296;
  assign n298 = n76 & n209;
  assign n299 = ~n117 & n298;
  assign n300 = ~pi00 & ~pi01;
  assign n301 = n112 & n300;
  assign n302 = n67 & n193;
  assign n303 = n160 & n302;
  assign n304 = ~n301 & ~n303;
  assign n305 = pi11 & ~n304;
  assign n306 = ~n67 & ~n182;
  assign n307 = n67 & ~n184;
  assign n308 = n160 & ~n306;
  assign n309 = ~n307 & n308;
  assign n310 = n122 & ~n132;
  assign n311 = ~n249 & n310;
  assign n312 = n249 & ~n310;
  assign n313 = ~n311 & ~n312;
  assign n314 = n247 & ~n313;
  assign n315 = ~n247 & n313;
  assign n316 = n142 & ~n314;
  assign n317 = ~n315 & n316;
  assign n318 = ~n305 & ~n309;
  assign n319 = ~n297 & n318;
  assign n320 = ~n299 & n319;
  assign n321 = ~n293 & n320;
  assign n322 = ~n273 & n321;
  assign n323 = ~n283 & n322;
  assign n324 = ~n317 & n323;
  assign n325 = ~n266 & n324;
  assign n326 = ~n176 & n325;
  assign n327 = n176 & ~n325;
  assign n328 = pi13 & ~n326;
  assign n329 = ~n327 & n328;
  assign n330 = n111 & ~n234;
  assign po1 = n329 | ~n330;
  assign n332 = ~pi02 & n38;
  assign n333 = n108 & n211;
  assign n334 = pi01 & ~pi05;
  assign n335 = ~n27 & ~n182;
  assign n336 = ~n334 & ~n335;
  assign n337 = ~pi06 & ~n336;
  assign n338 = pi09 & n337;
  assign n339 = pi06 & n51;
  assign n340 = n336 & n339;
  assign n341 = ~n338 & ~n340;
  assign n342 = pi02 & ~n341;
  assign n343 = pi06 & n336;
  assign n344 = ~n336 & ~n339;
  assign n345 = ~pi02 & pi09;
  assign n346 = ~n343 & n345;
  assign n347 = ~n344 & n346;
  assign n348 = ~n333 & ~n347;
  assign n349 = ~n342 & n348;
  assign n350 = n119 & ~n349;
  assign n351 = pi02 & pi06;
  assign n352 = ~n187 & n351;
  assign n353 = ~pi02 & ~pi06;
  assign n354 = n45 & ~n353;
  assign n355 = ~pi06 & ~n58;
  assign n356 = ~n354 & ~n355;
  assign n357 = ~n352 & n356;
  assign n358 = ~n350 & n357;
  assign n359 = ~n332 & n358;
  assign n360 = ~n34 & n359;
  assign n361 = ~pi06 & n78;
  assign n362 = ~n360 & ~n361;
  assign n363 = ~pi09 & ~n362;
  assign n364 = ~n88 & n351;
  assign n365 = n84 & n353;
  assign n366 = ~n364 & ~n365;
  assign n367 = pi09 & ~n366;
  assign n368 = pi09 & n89;
  assign n369 = ~pi02 & n28;
  assign n370 = n47 & n369;
  assign n371 = ~n368 & ~n370;
  assign n372 = pi06 & ~n371;
  assign n373 = pi02 & pi11;
  assign n374 = ~pi06 & ~pi09;
  assign n375 = n25 & ~n374;
  assign n376 = n373 & ~n375;
  assign n377 = pi02 & n112;
  assign n378 = pi06 & n96;
  assign n379 = ~n99 & ~n378;
  assign n380 = ~n377 & n379;
  assign n381 = ~n359 & ~n380;
  assign n382 = ~n367 & ~n376;
  assign n383 = ~n372 & n382;
  assign n384 = ~n381 & n383;
  assign n385 = ~n363 & n384;
  assign n386 = ~pi13 & ~n385;
  assign n387 = n121 & n351;
  assign n388 = ~pi02 & n359;
  assign n389 = n120 & ~n388;
  assign n390 = n24 & n359;
  assign n391 = pi09 & n359;
  assign n392 = pi02 & pi08;
  assign n393 = ~n374 & n392;
  assign n394 = ~n391 & n393;
  assign n395 = ~n390 & ~n394;
  assign n396 = n125 & ~n395;
  assign n397 = ~n389 & ~n396;
  assign n398 = n133 & n397;
  assign n399 = ~n387 & ~n398;
  assign n400 = n359 & n399;
  assign n401 = ~n359 & ~n399;
  assign n402 = ~n400 & ~n401;
  assign n403 = ~n209 & ~n251;
  assign n404 = ~n250 & ~n403;
  assign n405 = ~n402 & n404;
  assign n406 = n402 & ~n404;
  assign n407 = n48 & ~n405;
  assign n408 = ~n406 & n407;
  assign n409 = pi06 & n28;
  assign n410 = pi01 & ~n258;
  assign n411 = ~n260 & ~n410;
  assign n412 = ~n397 & n411;
  assign n413 = n397 & ~n411;
  assign n414 = ~n412 & ~n413;
  assign n415 = pi02 & ~pi08;
  assign n416 = n414 & n415;
  assign n417 = ~n409 & ~n416;
  assign n418 = ~n408 & n417;
  assign n419 = n64 & ~n418;
  assign n420 = n65 & ~n414;
  assign n421 = pi01 & ~n278;
  assign n422 = ~n277 & ~n421;
  assign n423 = n276 & ~n359;
  assign n424 = n422 & n423;
  assign n425 = ~n420 & ~n424;
  assign n426 = ~pi02 & ~n425;
  assign n427 = ~pi02 & n300;
  assign n428 = pi11 & n427;
  assign n429 = ~n300 & n373;
  assign n430 = n267 & n397;
  assign n431 = ~n267 & ~n397;
  assign n432 = ~n430 & ~n431;
  assign n433 = ~pi11 & ~n432;
  assign n434 = ~n428 & ~n429;
  assign n435 = ~n433 & n434;
  assign n436 = n112 & ~n435;
  assign n437 = ~n359 & ~n422;
  assign n438 = n286 & n437;
  assign n439 = ~n289 & ~n438;
  assign n440 = pi02 & ~n439;
  assign n441 = pi02 & ~n422;
  assign n442 = pi02 & n286;
  assign n443 = n276 & ~n422;
  assign n444 = ~n442 & ~n443;
  assign n445 = n359 & ~n441;
  assign n446 = ~n444 & n445;
  assign n447 = ~n67 & ~n184;
  assign n448 = ~n193 & ~n447;
  assign n449 = ~n351 & ~n353;
  assign n450 = ~n448 & ~n449;
  assign n451 = pi11 & n353;
  assign n452 = ~n351 & ~n451;
  assign n453 = n448 & n452;
  assign n454 = n160 & ~n450;
  assign n455 = ~n453 & n454;
  assign n456 = n299 & n359;
  assign n457 = ~pi10 & n294;
  assign n458 = n298 & ~n457;
  assign n459 = ~n295 & ~n359;
  assign n460 = ~n458 & n459;
  assign n461 = ~n247 & ~n312;
  assign n462 = ~n311 & ~n461;
  assign n463 = n399 & n462;
  assign n464 = ~n399 & ~n462;
  assign n465 = ~n463 & ~n464;
  assign n466 = n397 & ~n465;
  assign n467 = ~n397 & n465;
  assign n468 = n142 & ~n466;
  assign n469 = ~n467 & n468;
  assign n470 = ~n455 & ~n456;
  assign n471 = ~n460 & n470;
  assign n472 = ~n446 & n471;
  assign n473 = ~n440 & n472;
  assign n474 = ~n436 & n473;
  assign n475 = ~n426 & n474;
  assign n476 = ~n419 & n475;
  assign n477 = ~n469 & n476;
  assign n478 = pi13 & n327;
  assign n479 = ~n477 & n478;
  assign n480 = ~n327 & n477;
  assign n481 = pi13 & ~n479;
  assign n482 = ~n480 & n481;
  assign n483 = n111 & ~n386;
  assign po2 = n482 | ~n483;
  assign n485 = ~pi03 & ~pi07;
  assign n486 = n84 & n485;
  assign po5 = pi03 & pi07;
  assign n488 = ~n88 & po5;
  assign n489 = n45 & ~n485;
  assign n490 = pi02 & ~n343;
  assign n491 = ~n337 & ~n490;
  assign n492 = n125 & n491;
  assign n493 = ~n185 & ~n492;
  assign n494 = po5 & ~n493;
  assign n495 = pi07 & n51;
  assign n496 = n106 & n495;
  assign n497 = ~n491 & n496;
  assign n498 = ~n37 & ~n497;
  assign n499 = ~pi03 & ~n498;
  assign n500 = n108 & n373;
  assign n501 = pi09 & n485;
  assign n502 = n491 & n501;
  assign n503 = ~n500 & ~n502;
  assign n504 = pi13 & ~n503;
  assign n505 = ~n494 & ~n499;
  assign n506 = ~n504 & n505;
  assign n507 = ~pi08 & ~n506;
  assign n508 = pi03 & n53;
  assign n509 = ~n491 & n508;
  assign n510 = n58 & ~n509;
  assign n511 = ~pi07 & ~n510;
  assign n512 = ~n62 & ~n185;
  assign n513 = pi13 & po5;
  assign n514 = ~n512 & n513;
  assign n515 = ~n489 & ~n514;
  assign n516 = ~n511 & n515;
  assign n517 = ~n507 & n516;
  assign n518 = pi03 & ~n517;
  assign n519 = n48 & n518;
  assign n520 = ~n486 & ~n488;
  assign n521 = ~n519 & n520;
  assign n522 = pi09 & ~n521;
  assign n523 = ~n34 & n517;
  assign n524 = ~pi07 & n78;
  assign n525 = ~n523 & ~n524;
  assign n526 = ~pi09 & ~n525;
  assign n527 = pi07 & n96;
  assign n528 = ~n99 & ~n527;
  assign n529 = ~n517 & ~n528;
  assign n530 = pi03 & pi11;
  assign n531 = ~pi07 & ~pi09;
  assign n532 = n25 & ~n531;
  assign n533 = n530 & ~n532;
  assign n534 = ~pi03 & n28;
  assign n535 = n47 & n534;
  assign n536 = ~n368 & ~n535;
  assign n537 = pi07 & ~n536;
  assign n538 = ~n533 & ~n537;
  assign n539 = ~n529 & n538;
  assign n540 = ~n526 & n539;
  assign n541 = ~n522 & n540;
  assign n542 = ~pi13 & ~n541;
  assign n543 = ~pi03 & n517;
  assign n544 = n120 & ~n543;
  assign n545 = n55 & n518;
  assign n546 = n42 & po5;
  assign n547 = n24 & n517;
  assign n548 = ~n546 & ~n547;
  assign n549 = ~n545 & n548;
  assign n550 = n125 & ~n549;
  assign n551 = ~n544 & ~n550;
  assign n552 = n121 & po5;
  assign n553 = n133 & n551;
  assign n554 = ~n552 & ~n553;
  assign n555 = ~n397 & ~n463;
  assign n556 = ~n464 & ~n555;
  assign n557 = n554 & n556;
  assign n558 = ~n554 & ~n556;
  assign n559 = ~n557 & ~n558;
  assign n560 = n551 & ~n559;
  assign n561 = ~n551 & n559;
  assign n562 = n270 & ~n560;
  assign n563 = ~n561 & n562;
  assign n564 = ~pi03 & n112;
  assign n565 = n427 & n564;
  assign n566 = ~n351 & ~n448;
  assign n567 = ~n353 & ~n566;
  assign n568 = ~pi07 & n567;
  assign n569 = ~pi03 & n160;
  assign n570 = n568 & n569;
  assign n571 = ~n565 & ~n570;
  assign n572 = ~n563 & n571;
  assign n573 = pi11 & ~n572;
  assign n574 = ~n517 & n554;
  assign n575 = n517 & ~n554;
  assign n576 = ~n574 & ~n575;
  assign n577 = ~n400 & ~n404;
  assign n578 = ~n401 & ~n577;
  assign n579 = n576 & n578;
  assign n580 = ~n576 & ~n578;
  assign n581 = pi08 & ~n579;
  assign n582 = ~n580 & n581;
  assign n583 = ~pi02 & n397;
  assign n584 = ~n411 & ~n583;
  assign n585 = pi02 & ~n397;
  assign n586 = ~n584 & ~n585;
  assign n587 = ~n551 & ~n586;
  assign n588 = ~pi03 & ~n587;
  assign n589 = n551 & n586;
  assign n590 = ~pi08 & ~n589;
  assign n591 = n588 & n590;
  assign n592 = ~n582 & ~n591;
  assign n593 = n185 & ~n592;
  assign n594 = pi02 & ~n358;
  assign n595 = ~n437 & ~n594;
  assign n596 = ~n441 & n595;
  assign n597 = ~n517 & n596;
  assign n598 = n517 & ~n596;
  assign n599 = ~n597 & ~n598;
  assign n600 = n286 & n599;
  assign n601 = ~n289 & ~n600;
  assign n602 = pi03 & ~n601;
  assign n603 = n276 & ~n599;
  assign n604 = pi07 & n160;
  assign n605 = ~n567 & n604;
  assign n606 = ~n603 & ~n605;
  assign n607 = ~pi03 & ~n606;
  assign n608 = pi07 & ~n567;
  assign n609 = pi03 & n160;
  assign n610 = ~n568 & n609;
  assign n611 = ~n608 & n610;
  assign n612 = n456 & n517;
  assign n613 = n112 & n530;
  assign n614 = ~n427 & n613;
  assign n615 = n298 & n359;
  assign n616 = ~n457 & n615;
  assign n617 = ~n295 & ~n517;
  assign n618 = ~n616 & n617;
  assign n619 = n430 & n551;
  assign n620 = ~n430 & ~n551;
  assign n621 = ~n619 & ~n620;
  assign n622 = n112 & ~n621;
  assign n623 = ~n587 & ~n589;
  assign n624 = pi03 & n24;
  assign n625 = ~n623 & n624;
  assign n626 = ~n604 & ~n622;
  assign n627 = ~n625 & n626;
  assign n628 = ~pi11 & ~n627;
  assign n629 = ~n611 & ~n614;
  assign n630 = ~n612 & n629;
  assign n631 = ~n618 & n630;
  assign n632 = ~n602 & n631;
  assign n633 = ~n607 & n632;
  assign n634 = ~n628 & n633;
  assign n635 = ~n593 & n634;
  assign n636 = ~n573 & n635;
  assign n637 = ~n479 & n636;
  assign n638 = n479 & ~n636;
  assign n639 = pi13 & ~n637;
  assign n640 = ~n638 & n639;
  assign n641 = n111 & ~n542;
  assign po3 = n640 | ~n641;
  assign po4 = n485 | po5;
  assign n644 = ~po5 & ~n567;
  assign n645 = n160 & ~n485;
  assign n646 = ~n644 & n645;
  assign n647 = ~n518 & n596;
  assign n648 = ~n275 & ~n543;
  assign n649 = ~n647 & n648;
  assign n650 = n551 & ~n558;
  assign n651 = n270 & ~n557;
  assign n652 = ~n650 & n651;
  assign n653 = ~n565 & ~n646;
  assign n654 = ~n649 & n653;
  assign n655 = ~n652 & n654;
  assign n656 = pi11 & ~n655;
  assign n657 = ~n28 & ~n84;
  assign n658 = pi09 & ~n657;
  assign n659 = n615 & n658;
  assign n660 = n517 & n659;
  assign n661 = ~n588 & n590;
  assign n662 = n554 & n578;
  assign n663 = ~n554 & ~n578;
  assign n664 = n517 & ~n663;
  assign n665 = pi08 & ~n662;
  assign n666 = ~n664 & n665;
  assign n667 = ~n661 & ~n666;
  assign n668 = n108 & ~n667;
  assign n669 = pi10 & ~n619;
  assign n670 = n55 & ~n669;
  assign n671 = ~n668 & ~n670;
  assign n672 = ~pi11 & ~n671;
  assign n673 = ~n656 & ~n660;
  assign n674 = ~n672 & n673;
  assign n675 = ~n638 & n674;
  assign po6 = pi13 & ~n675;
  assign n677 = ~n69 & ~n196;
  assign n678 = ~n449 & po4;
  assign po7 = n677 & n678;
endmodule
