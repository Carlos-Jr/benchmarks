module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 , pi16 ,
    pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 , pi11 , pi12 , pi13 , pi14 , pi15 ,
    pi16 , pi17 , pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ,
    po7 , po8 , po9 , po10 , po11 , po12 ,
    po13 , po14 , po15 , po16 , po17 , po18 ,
    po19 , po20 , po21 , po22 , po23 , po24 ;
  wire n50, n51, n52, n53, n54, n55, n56,
    n57, n58, n59, n60, n61, n62, n63, n64,
    n65, n66, n67, n68, n69, n70, n71, n72,
    n73, n74, n75, n76, n77, n78, n79, n80,
    n81, n82, n83, n84, n85, n86, n87, n88,
    n89, n90, n91, n92, n93, n94, n95, n96,
    n97, n98, n99, n100, n101, n102, n103,
    n104, n105, n106, n107, n108, n109, n110,
    n111, n112, n113, n114, n115, n116, n117,
    n118, n119, n120, n121, n122, n123, n124,
    n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138,
    n139, n140, n141, n142, n143, n144, n145,
    n146, n147, n148, n149, n150, n151, n152,
    n153, n154, n155, n156, n157, n158, n159,
    n160, n161, n162, n163, n164, n165, n166,
    n167, n168, n169, n170, n171, n172, n173,
    n174, n175, n176, n177, n178, n179, n180,
    n181, n182, n183, n184, n185, n186, n187,
    n188, n189, n190, n191, n192, n193, n194,
    n195, n196, n197, n198, n199, n200, n201,
    n202, n203, n204, n205, n206, n207, n208,
    n209, n210, n211, n212, n213, n214, n215,
    n216, n217, n218, n219, n220, n221, n222,
    n223, n224, n225, n226, n227, n228, n229,
    n230, n231, n232, n233, n234, n235, n236,
    n237, n238, n239, n240, n241, n242, n243,
    n244, n245, n246, n247, n248, n249, n250,
    n251, n252, n253, n254, n255, n256, n257,
    n258, n259, n260, n261, n262, n263, n264,
    n265, n266, n267, n268, n269, n270, n271,
    n272, n273, n274, n275, n276, n277, n278,
    n279, n280, n281, n282, n283, n284, n285,
    n286, n287, n288, n289, n290, n291, n292,
    n293, n294, n295, n296, n297, n298, n299,
    n300, n301, n302, n303, n304, n305, n306,
    n307, n308, n309, n310, n311, n312, n313,
    n314, n315, n316, n317, n318, n319, n320,
    n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n334,
    n335, n336, n337, n338, n339, n340, n341,
    n342, n343, n344, n345, n346, n347, n348,
    n349, n350, n351, n352, n353, n354, n355,
    n356, n357, n358, n359, n360, n361, n362,
    n363, n364, n365, n366, n367, n368, n369,
    n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n405, n406, n407, n408, n409, n410, n411,
    n412, n413, n414, n415, n416, n417, n418,
    n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432,
    n433, n434, n435, n436, n437, n438, n439,
    n440, n441, n442, n443, n444, n445, n446,
    n447, n448, n449, n450, n451, n452, n453,
    n454, n455, n456, n457, n458, n459, n460,
    n461, n462, n463, n464, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481,
    n482, n483, n484, n485, n486, n487, n488,
    n489, n490, n491, n492, n493, n494, n495,
    n496, n497, n498, n499, n500, n501, n502,
    n503, n504, n505, n506, n507, n508, n509,
    n510, n511, n512, n513, n514, n515, n516,
    n517, n518, n519, n520, n521, n522, n523,
    n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537,
    n538, n539, n540, n541, n542, n543, n544,
    n545, n546, n547, n548, n549, n550, n551,
    n552, n553, n554, n555, n556, n557, n558,
    n559, n560, n561, n562, n563, n564, n565,
    n566, n567, n568, n569, n570, n571, n572,
    n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586,
    n587, n588, n589, n590, n591, n592, n593,
    n594, n595, n596, n597, n598, n599, n600,
    n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614,
    n615, n616, n617, n618, n619, n620, n621,
    n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635,
    n636, n637, n638, n639, n640, n641, n642,
    n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591,
    n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3626, n3627,
    n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651,
    n3652, n3653, n3654, n3655, n3656, n3657,
    n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681,
    n3682, n3683, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3693, n3694,
    n3695, n3696, n3697, n3698, n3699, n3700,
    n3701, n3702, n3703, n3704, n3705, n3706,
    n3707, n3708, n3709, n3710, n3711, n3712,
    n3713, n3714, n3715, n3716, n3717, n3718,
    n3719, n3720, n3721, n3722, n3723, n3724,
    n3725, n3726, n3727, n3728, n3729, n3730,
    n3731, n3732, n3733, n3734, n3735, n3736,
    n3737, n3738, n3739, n3740, n3741, n3742,
    n3743, n3744, n3745, n3746, n3747, n3748,
    n3749, n3750, n3751, n3752, n3753, n3754,
    n3755, n3756, n3757, n3758, n3759, n3760,
    n3761, n3762, n3763, n3764, n3765, n3766,
    n3767, n3768, n3769, n3770, n3771, n3772,
    n3773, n3774, n3775, n3776, n3777, n3778,
    n3779, n3780, n3781, n3782, n3783, n3784,
    n3785, n3786, n3787, n3788, n3789, n3790,
    n3791, n3792, n3793, n3794, n3795, n3796,
    n3797, n3798, n3799, n3800, n3801, n3802,
    n3803, n3804, n3805, n3806, n3807, n3808,
    n3809, n3810, n3811, n3812, n3813, n3814,
    n3815, n3816, n3817, n3818, n3819, n3820,
    n3821, n3822, n3823, n3824, n3825, n3826,
    n3827, n3828, n3829, n3830, n3831, n3832,
    n3833, n3834, n3835, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845,
    n3846, n3847, n3848, n3849, n3850, n3851,
    n3852, n3853, n3854, n3855, n3856, n3857,
    n3858, n3859, n3860, n3861, n3862, n3863,
    n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875,
    n3876, n3877, n3878, n3879, n3880, n3881,
    n3882, n3883, n3884, n3885, n3886, n3887,
    n3888, n3889, n3890, n3891, n3892, n3893,
    n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3901, n3902, n3903, n3904, n3905,
    n3906, n3907, n3908, n3909, n3910, n3911,
    n3912, n3913, n3914, n3915, n3916, n3917,
    n3918, n3919, n3920, n3921, n3922, n3923,
    n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3934, n3935,
    n3936, n3937, n3938, n3939, n3940, n3941,
    n3942, n3943, n3944, n3945, n3946, n3947,
    n3948, n3949, n3950, n3951, n3952, n3953,
    n3954, n3956, n3957, n3958, n3959, n3960,
    n3961, n3962, n3963, n3964, n3965, n3966,
    n3967, n3968, n3969, n3970, n3971, n3972,
    n3973, n3974, n3975, n3976, n3977, n3978,
    n3979, n3980, n3981, n3982, n3983, n3984,
    n3985, n3986, n3987, n3988, n3989, n3990,
    n3991, n3992, n3993, n3994, n3995, n3996,
    n3997, n3998, n3999, n4000, n4001, n4002,
    n4003, n4004, n4005, n4006, n4007, n4008,
    n4009, n4010, n4011, n4012, n4013, n4014,
    n4015, n4016, n4017, n4018, n4019, n4020,
    n4021, n4022, n4023, n4024, n4025, n4026,
    n4027, n4028, n4029, n4030, n4031, n4032,
    n4033, n4034, n4035, n4036, n4037, n4038,
    n4039, n4040, n4041, n4042, n4043, n4044,
    n4045, n4046, n4047, n4048, n4049, n4050,
    n4051, n4052, n4053, n4054, n4055, n4056,
    n4057, n4058, n4059, n4060, n4061, n4062,
    n4063, n4064, n4065, n4066, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075,
    n4076, n4077, n4078, n4079, n4080, n4081,
    n4082, n4083, n4084, n4085, n4086, n4087,
    n4088, n4089, n4090, n4091, n4092, n4093,
    n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105,
    n4106, n4107, n4108, n4109, n4110, n4111,
    n4112, n4113, n4114, n4115, n4116, n4117,
    n4118, n4119, n4120, n4121, n4122, n4123,
    n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135,
    n4136, n4137, n4138, n4139, n4140, n4141,
    n4142, n4143, n4144, n4145, n4146, n4147,
    n4148, n4149, n4150, n4151, n4152, n4153,
    n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165,
    n4166, n4167, n4168, n4169, n4170, n4172,
    n4173, n4174, n4175, n4176, n4177, n4178,
    n4179, n4180, n4181, n4182, n4183, n4184,
    n4185, n4186, n4187, n4188, n4189, n4190,
    n4191, n4192, n4193, n4194, n4195, n4196,
    n4197, n4198, n4199, n4200, n4201, n4202,
    n4203, n4204, n4205, n4206, n4207, n4208,
    n4209, n4210, n4211, n4212, n4213, n4214,
    n4215, n4216, n4217, n4218, n4219, n4220,
    n4221, n4222, n4223, n4224, n4225, n4226,
    n4227, n4228, n4229, n4230, n4231, n4232,
    n4233, n4234, n4235, n4236, n4237, n4238,
    n4239, n4240, n4241, n4242, n4243, n4244,
    n4245, n4246, n4247, n4248, n4249, n4250,
    n4251, n4252, n4253, n4254, n4255, n4256,
    n4257, n4258, n4259, n4260, n4261, n4262,
    n4263, n4264, n4265, n4266, n4267, n4268,
    n4269, n4270, n4271, n4272, n4273, n4274,
    n4275, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317,
    n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341,
    n4342, n4343, n4344, n4345, n4346, n4347,
    n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4375, n4376, n4377,
    n4378, n4379, n4381, n4382, n4383, n4384,
    n4385, n4386, n4387, n4388, n4389, n4390,
    n4391, n4392, n4393, n4394, n4395, n4396,
    n4397, n4398, n4399, n4400, n4401, n4402,
    n4403, n4404, n4405, n4406, n4407, n4408,
    n4409, n4410, n4411, n4412, n4413, n4414,
    n4415, n4416, n4417, n4418, n4419, n4420,
    n4421, n4422, n4423, n4424, n4425, n4426,
    n4427, n4428, n4429, n4430, n4431, n4432,
    n4433, n4434, n4435, n4436, n4437, n4438,
    n4439, n4440, n4441, n4442, n4443, n4444,
    n4445, n4446, n4447, n4448, n4449, n4450,
    n4451, n4452, n4453, n4454, n4455, n4456,
    n4457, n4458, n4459, n4460, n4461, n4462,
    n4463, n4464, n4465, n4466, n4467, n4468,
    n4469, n4470, n4471, n4473, n4474, n4475,
    n4476, n4477, n4478, n4479, n4480, n4481,
    n4482, n4483, n4484, n4485, n4486, n4487,
    n4488, n4489, n4490, n4491, n4492, n4493,
    n4494, n4495, n4496, n4497, n4498, n4499,
    n4500, n4501, n4502, n4503, n4504, n4505,
    n4506, n4507, n4508, n4509, n4510, n4511,
    n4512, n4513, n4514, n4515, n4516, n4517,
    n4518, n4519, n4520, n4521, n4522, n4523,
    n4524, n4525, n4526, n4527, n4528, n4529,
    n4530, n4531, n4532, n4533, n4534, n4535,
    n4536, n4537, n4538, n4539, n4540, n4541,
    n4542, n4543, n4544, n4545, n4546, n4547,
    n4548, n4549, n4550, n4551, n4552, n4553,
    n4554, n4555, n4556, n4557, n4558, n4559,
    n4560, n4561, n4562, n4564, n4565, n4566,
    n4567, n4568, n4569, n4570, n4571, n4572,
    n4573, n4574, n4575, n4576, n4577, n4578,
    n4579, n4580, n4581, n4582, n4583, n4584,
    n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596,
    n4597, n4598, n4599, n4600, n4601, n4602,
    n4603, n4604, n4605, n4606, n4607, n4608,
    n4609, n4610, n4611, n4612, n4613, n4614,
    n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626,
    n4627, n4628, n4629, n4630, n4631, n4632,
    n4633, n4634, n4635, n4636, n4637, n4638,
    n4639, n4640, n4641, n4642, n4644, n4645,
    n4646, n4647, n4648, n4649, n4650, n4651,
    n4652, n4653, n4654, n4655, n4656, n4657,
    n4658, n4659, n4660, n4661, n4662, n4663,
    n4664, n4665, n4666, n4667, n4668, n4669,
    n4670, n4671, n4672, n4673, n4674, n4675,
    n4676, n4677, n4678, n4679, n4680, n4681,
    n4682, n4683, n4684, n4685, n4686, n4687,
    n4688, n4689, n4690, n4691, n4692, n4693,
    n4694, n4695, n4696, n4697, n4698, n4699,
    n4700, n4701, n4702, n4703, n4704, n4705,
    n4706, n4707, n4708, n4709, n4710, n4711,
    n4712, n4713, n4714, n4715, n4716, n4717,
    n4718, n4719, n4721, n4722, n4723, n4724,
    n4725, n4726, n4727, n4728, n4729, n4730,
    n4731, n4732, n4733, n4734, n4735, n4736,
    n4737, n4738, n4739, n4740, n4741, n4742,
    n4743, n4744, n4745, n4746, n4747, n4748,
    n4749, n4750, n4751, n4752, n4753, n4754,
    n4755, n4756, n4757, n4758, n4759, n4760,
    n4761, n4762, n4763, n4764, n4765, n4766,
    n4767, n4768, n4769, n4770, n4771, n4772,
    n4773, n4774, n4775, n4776, n4777, n4778,
    n4779, n4780, n4781, n4782, n4783, n4785,
    n4786, n4787, n4788, n4789, n4790, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797,
    n4798, n4799, n4800, n4801, n4802, n4803,
    n4804, n4805, n4806, n4807, n4808, n4809,
    n4810, n4811, n4812, n4813, n4814, n4815,
    n4816, n4817, n4818, n4819, n4820, n4821,
    n4822, n4823, n4824, n4825, n4826, n4827,
    n4828, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845,
    n4846, n4847, n4849, n4850, n4851, n4852,
    n4853, n4854, n4855, n4856, n4857, n4858,
    n4859, n4860, n4861, n4862, n4863, n4864,
    n4865, n4866, n4867, n4868, n4869, n4870,
    n4871, n4872, n4873, n4874, n4875, n4876,
    n4877, n4878, n4879, n4880, n4881, n4882,
    n4883, n4884, n4885, n4886, n4887, n4888,
    n4889, n4890, n4891, n4892, n4893, n4894,
    n4895, n4896, n4897, n4898, n4899, n4900,
    n4901, n4902, n4903, n4904, n4905, n4906,
    n4907, n4908, n4909, n4910, n4912, n4913,
    n4914, n4915, n4916, n4917, n4918, n4919,
    n4920, n4921, n4922, n4923, n4924, n4925,
    n4926, n4927, n4928, n4929, n4930, n4931,
    n4932, n4933, n4934, n4935, n4936, n4937,
    n4938, n4939, n4940, n4941, n4942, n4943,
    n4944, n4945, n4946, n4947, n4948, n4949,
    n4950, n4951, n4952, n4953, n4954, n4955,
    n4956, n4957, n4958, n4959, n4960, n4961,
    n4962, n4963, n4965, n4966, n4967, n4968,
    n4969, n4970, n4971, n4972, n4973, n4974,
    n4975, n4976, n4977, n4978, n4979, n4980,
    n4981, n4982, n4983, n4984, n4985, n4986,
    n4987, n4988, n4989, n4990, n4991, n4992,
    n4993, n4994, n4995, n4996, n4997, n4998,
    n4999, n5000, n5001, n5002, n5003, n5004,
    n5005, n5006, n5007, n5008, n5009, n5010,
    n5012, n5013, n5014, n5015, n5016, n5017,
    n5018, n5019, n5020, n5021, n5022, n5023,
    n5024, n5025, n5026, n5027, n5028, n5029,
    n5030, n5031, n5032, n5033, n5034, n5035,
    n5036, n5037, n5038, n5039, n5040, n5041,
    n5042, n5043, n5044, n5045, n5046, n5047,
    n5048, n5049, n5051, n5052, n5053, n5054,
    n5055, n5056, n5057, n5058, n5059, n5060,
    n5061, n5062, n5063, n5064, n5065, n5066,
    n5067, n5068, n5069, n5070, n5071, n5072,
    n5073, n5075, n5076, n5077, n5078, n5079,
    n5080, n5081, n5082, n5083, n5084, n5085,
    n5086, n5087, n5088, n5089, n5090, n5091,
    n5092, n5093, n5095, n5096, n5097, n5098,
    n5099, n5100, n5101, n5102, n5103, n5104,
    n5105, n5106, n5107, n5108, n5109, n5110,
    n5111, n5112, n5113, n5114, n5115, n5116,
    n5118, n5119, n5120, n5121, n5122, n5123,
    n5124, n5125, n5126, n5127, n5128, n5129,
    n5130, n5131, n5132, n5133, n5135, n5136,
    n5137, n5138, n5139, n5140, n5141, n5142,
    n5143, n5144, n5145, n5146, n5147, n5148,
    n5149, n5151, n5152, n5153, n5154, n5155,
    n5156, n5157, n5158, n5159, n5161, n5162,
    n5163, n5164, n5165, n5166, n5167, n5168,
    n5169, n5171, n5172, n5173, n5174, n5175;
  assign n50 = ~pi0  & ~pi1 ;
  assign n51 = ~pi2  & n50;
  assign n52 = ~pi3  & n51;
  assign n53 = ~pi4  & n52;
  assign n54 = ~pi22  & ~n53;
  assign n55 = pi5  & ~n54;
  assign n56 = ~pi5  & n54;
  assign n57 = ~n55 & ~n56;
  assign n58 = ~pi22  & ~n51;
  assign n59 = pi3  & ~n58;
  assign n60 = ~pi3  & n58;
  assign n61 = ~n59 & ~n60;
  assign n62 = pi2  & pi22 ;
  assign n63 = pi2  & ~n50;
  assign n64 = n58 & ~n63;
  assign n65 = ~n62 & ~n64;
  assign n66 = n61 & n65;
  assign n67 = ~n61 & ~n65;
  assign n68 = ~n66 & ~n67;
  assign n69 = pi4  & pi22 ;
  assign n70 = pi4  & ~n52;
  assign n71 = n54 & ~n70;
  assign n72 = ~n69 & ~n71;
  assign n73 = n61 & n72;
  assign n74 = ~n61 & ~n72;
  assign n75 = ~n73 & ~n74;
  assign n76 = ~n68 & n75;
  assign n77 = ~pi5  & n53;
  assign n78 = ~pi6  & n77;
  assign n79 = ~pi7  & n78;
  assign n80 = ~pi8  & n79;
  assign n81 = ~pi9  & n80;
  assign n82 = ~pi10  & n81;
  assign n83 = ~pi11  & n82;
  assign n84 = ~pi12  & n83;
  assign n85 = ~pi13  & n84;
  assign n86 = ~pi14  & n85;
  assign n87 = ~pi15  & n86;
  assign n88 = ~pi16  & n87;
  assign n89 = ~pi22  & ~n88;
  assign n90 = pi17  & ~n89;
  assign n91 = ~pi17  & n89;
  assign n92 = ~n90 & ~n91;
  assign n93 = ~pi22  & ~n87;
  assign n94 = pi16  & ~n93;
  assign n95 = ~pi16  & n93;
  assign n96 = ~n94 & ~n95;
  assign n97 = n92 & n96;
  assign n98 = ~pi17  & n88;
  assign n99 = ~pi18  & n98;
  assign n100 = ~pi22  & ~n99;
  assign n101 = pi19  & ~n100;
  assign n102 = ~pi19  & n100;
  assign n103 = ~n101 & ~n102;
  assign n104 = pi18  & pi22 ;
  assign n105 = pi18  & ~n98;
  assign n106 = n100 & ~n105;
  assign n107 = ~n104 & ~n106;
  assign n108 = ~n103 & ~n107;
  assign n109 = n97 & n108;
  assign n110 = pi15  & pi22 ;
  assign n111 = pi15  & ~n86;
  assign n112 = n93 & ~n111;
  assign n113 = ~n110 & ~n112;
  assign n114 = pi21  & pi22 ;
  assign n115 = ~pi19  & n99;
  assign n116 = ~pi20  & n115;
  assign n117 = pi21  & ~n116;
  assign n118 = ~pi21  & n116;
  assign n119 = ~pi22  & ~n117;
  assign n120 = ~n118 & n119;
  assign n121 = ~n114 & ~n120;
  assign n122 = pi20  & pi22 ;
  assign n123 = pi20  & ~n115;
  assign n124 = ~pi22  & ~n116;
  assign n125 = ~n123 & n124;
  assign n126 = ~n122 & ~n125;
  assign n127 = n121 & ~n126;
  assign n128 = ~n113 & n127;
  assign n129 = n109 & n128;
  assign n130 = ~n92 & n96;
  assign n131 = n103 & n107;
  assign n132 = n130 & n131;
  assign n133 = n128 & n132;
  assign n134 = ~n129 & ~n133;
  assign n135 = n103 & ~n107;
  assign n136 = ~n92 & ~n96;
  assign n137 = n135 & n136;
  assign n138 = n128 & n137;
  assign n139 = n108 & n130;
  assign n140 = n121 & n126;
  assign n141 = n113 & n140;
  assign n142 = n139 & n141;
  assign n143 = ~n113 & n140;
  assign n144 = n132 & n143;
  assign n145 = ~n121 & ~n126;
  assign n146 = ~n103 & n107;
  assign n147 = n92 & ~n96;
  assign n148 = n146 & n147;
  assign n149 = n145 & n148;
  assign n150 = n113 & n149;
  assign n151 = n97 & n131;
  assign n152 = n128 & n151;
  assign n153 = ~n121 & n126;
  assign n154 = ~n113 & n153;
  assign n155 = n97 & n135;
  assign n156 = n154 & n155;
  assign n157 = n135 & n147;
  assign n158 = n154 & n157;
  assign n159 = ~n156 & ~n158;
  assign n160 = ~n152 & n159;
  assign n161 = n131 & n147;
  assign n162 = n143 & n161;
  assign n163 = n130 & n146;
  assign n164 = n113 & n127;
  assign n165 = n163 & n164;
  assign n166 = n136 & n146;
  assign n167 = n154 & n166;
  assign n168 = n148 & n154;
  assign n169 = ~n162 & ~n165;
  assign n170 = ~n167 & ~n168;
  assign n171 = n169 & n170;
  assign n172 = n139 & n143;
  assign n173 = n97 & n146;
  assign n174 = n141 & n173;
  assign n175 = n128 & n161;
  assign n176 = n130 & n135;
  assign n177 = n164 & n176;
  assign n178 = n113 & n145;
  assign n179 = n173 & n178;
  assign n180 = n148 & n164;
  assign n181 = ~n172 & ~n174;
  assign n182 = ~n175 & ~n177;
  assign n183 = ~n179 & ~n180;
  assign n184 = n182 & n183;
  assign n185 = n181 & n184;
  assign n186 = ~n138 & ~n142;
  assign n187 = ~n144 & ~n150;
  assign n188 = n186 & n187;
  assign n189 = n134 & n188;
  assign n190 = n160 & n171;
  assign n191 = n189 & n190;
  assign n192 = n185 & n191;
  assign n193 = n151 & n178;
  assign n194 = n161 & n178;
  assign n195 = n143 & n151;
  assign n196 = ~n194 & ~n195;
  assign n197 = n131 & n136;
  assign n198 = n145 & n197;
  assign n199 = ~n113 & n198;
  assign n200 = n141 & n163;
  assign n201 = n155 & n164;
  assign n202 = n109 & n141;
  assign n203 = n108 & n147;
  assign n204 = n164 & n203;
  assign n205 = ~n193 & ~n199;
  assign n206 = ~n200 & ~n201;
  assign n207 = ~n202 & ~n204;
  assign n208 = n206 & n207;
  assign n209 = n196 & n205;
  assign n210 = n208 & n209;
  assign n211 = ~n113 & n145;
  assign n212 = n137 & n211;
  assign n213 = n108 & n136;
  assign n214 = n143 & n213;
  assign n215 = n127 & n166;
  assign n216 = ~n113 & n215;
  assign n217 = n137 & n154;
  assign n218 = n164 & n197;
  assign n219 = n140 & n166;
  assign n220 = n113 & n219;
  assign n221 = ~n212 & ~n214;
  assign n222 = ~n216 & ~n217;
  assign n223 = ~n218 & ~n220;
  assign n224 = n222 & n223;
  assign n225 = n221 & n224;
  assign n226 = n139 & n153;
  assign n227 = n155 & n178;
  assign n228 = n143 & n197;
  assign n229 = n141 & n148;
  assign n230 = n137 & n141;
  assign n231 = n113 & n153;
  assign n232 = n173 & n231;
  assign n233 = n143 & n176;
  assign n234 = n128 & n173;
  assign n235 = ~n233 & ~n234;
  assign n236 = n128 & n213;
  assign n237 = n141 & n203;
  assign n238 = ~n236 & ~n237;
  assign n239 = n113 & n198;
  assign n240 = n109 & n231;
  assign n241 = n157 & n164;
  assign n242 = n153 & n163;
  assign n243 = n113 & n242;
  assign n244 = n176 & n231;
  assign n245 = n173 & n211;
  assign n246 = n137 & n178;
  assign n247 = ~n245 & ~n246;
  assign n248 = ~n240 & ~n241;
  assign n249 = ~n243 & ~n244;
  assign n250 = n248 & n249;
  assign n251 = n247 & n250;
  assign n252 = n139 & n164;
  assign n253 = n143 & n157;
  assign n254 = n155 & n231;
  assign n255 = n143 & n155;
  assign n256 = ~n254 & ~n255;
  assign n257 = ~n253 & n256;
  assign n258 = ~n229 & ~n230;
  assign n259 = ~n232 & ~n239;
  assign n260 = ~n252 & n259;
  assign n261 = n235 & n258;
  assign n262 = n238 & n261;
  assign n263 = n257 & n260;
  assign n264 = n262 & n263;
  assign n265 = n251 & n264;
  assign n266 = n132 & n154;
  assign n267 = n154 & n203;
  assign n268 = n161 & n231;
  assign n269 = ~n266 & ~n267;
  assign n270 = ~n268 & n269;
  assign n271 = n151 & n211;
  assign n272 = n155 & n211;
  assign n273 = n128 & n176;
  assign n274 = ~n271 & ~n272;
  assign n275 = ~n273 & n274;
  assign n276 = ~n226 & ~n227;
  assign n277 = ~n228 & n276;
  assign n278 = n270 & n277;
  assign n279 = n275 & n278;
  assign n280 = n210 & n225;
  assign n281 = n279 & n280;
  assign n282 = n192 & n281;
  assign n283 = n265 & n282;
  assign n284 = n132 & n178;
  assign n285 = n163 & n211;
  assign n286 = n132 & n231;
  assign n287 = ~n285 & ~n286;
  assign n288 = ~n284 & n287;
  assign n289 = n143 & n148;
  assign n290 = n128 & n148;
  assign n291 = n109 & n154;
  assign n292 = n164 & n213;
  assign n293 = ~n289 & ~n290;
  assign n294 = ~n291 & ~n292;
  assign n295 = n293 & n294;
  assign n296 = n203 & n231;
  assign n297 = ~n113 & n226;
  assign n298 = ~n142 & ~n297;
  assign n299 = ~n113 & n149;
  assign n300 = n109 & n178;
  assign n301 = ~n236 & ~n299;
  assign n302 = ~n300 & n301;
  assign n303 = n203 & n211;
  assign n304 = n109 & n164;
  assign n305 = ~n202 & ~n303;
  assign n306 = ~n304 & n305;
  assign n307 = ~n199 & ~n218;
  assign n308 = ~n243 & ~n296;
  assign n309 = n307 & n308;
  assign n310 = n298 & n309;
  assign n311 = n288 & n295;
  assign n312 = n302 & n306;
  assign n313 = n311 & n312;
  assign n314 = n310 & n313;
  assign n315 = n128 & n139;
  assign n316 = ~n241 & ~n315;
  assign n317 = n141 & n161;
  assign n318 = ~n253 & ~n266;
  assign n319 = n141 & n197;
  assign n320 = n154 & n161;
  assign n321 = ~n319 & ~n320;
  assign n322 = ~n200 & ~n317;
  assign n323 = n316 & n322;
  assign n324 = n318 & n321;
  assign n325 = n323 & n324;
  assign n326 = n134 & n325;
  assign n327 = n143 & n203;
  assign n328 = n113 & n226;
  assign n329 = ~n204 & ~n328;
  assign n330 = ~n228 & ~n327;
  assign n331 = n329 & n330;
  assign n332 = n148 & n231;
  assign n333 = ~n267 & ~n332;
  assign n334 = n109 & n211;
  assign n335 = ~n168 & ~n334;
  assign n336 = n178 & n213;
  assign n337 = n128 & n155;
  assign n338 = ~n336 & ~n337;
  assign n339 = n154 & n173;
  assign n340 = n178 & n203;
  assign n341 = ~n339 & ~n340;
  assign n342 = n211 & n213;
  assign n343 = n139 & n178;
  assign n344 = ~n239 & ~n343;
  assign n345 = ~n138 & ~n165;
  assign n346 = n141 & n157;
  assign n347 = n137 & n164;
  assign n348 = n163 & n178;
  assign n349 = n145 & n166;
  assign n350 = n113 & n349;
  assign n351 = ~n348 & ~n350;
  assign n352 = n139 & n211;
  assign n353 = n161 & n211;
  assign n354 = ~n352 & ~n353;
  assign n355 = n137 & n143;
  assign n356 = n157 & n231;
  assign n357 = ~n244 & ~n356;
  assign n358 = n151 & n164;
  assign n359 = ~n172 & ~n358;
  assign n360 = n132 & n211;
  assign n361 = ~n272 & ~n360;
  assign n362 = ~n113 & n349;
  assign n363 = ~n355 & ~n362;
  assign n364 = n357 & n363;
  assign n365 = n359 & n361;
  assign n366 = n364 & n365;
  assign n367 = ~n158 & ~n227;
  assign n368 = ~n346 & ~n347;
  assign n369 = n367 & n368;
  assign n370 = n344 & n345;
  assign n371 = n351 & n354;
  assign n372 = n370 & n371;
  assign n373 = n369 & n372;
  assign n374 = n366 & n373;
  assign n375 = ~n174 & ~n342;
  assign n376 = n374 & n375;
  assign n377 = n132 & n164;
  assign n378 = ~n113 & n219;
  assign n379 = ~n152 & ~n162;
  assign n380 = ~n377 & ~n378;
  assign n381 = n379 & n380;
  assign n382 = n333 & n335;
  assign n383 = n338 & n341;
  assign n384 = n382 & n383;
  assign n385 = n331 & n381;
  assign n386 = n384 & n385;
  assign n387 = n326 & n386;
  assign n388 = n314 & n387;
  assign n389 = n376 & n388;
  assign n390 = ~n283 & ~n389;
  assign n391 = n132 & n141;
  assign n392 = n128 & n197;
  assign n393 = ~n214 & ~n228;
  assign n394 = ~n392 & n393;
  assign n395 = ~n152 & ~n303;
  assign n396 = n166 & n231;
  assign n397 = ~n254 & ~n300;
  assign n398 = ~n220 & ~n290;
  assign n399 = ~n334 & ~n396;
  assign n400 = n395 & n399;
  assign n401 = n397 & n398;
  assign n402 = n400 & n401;
  assign n403 = n145 & n157;
  assign n404 = n141 & n213;
  assign n405 = n141 & n176;
  assign n406 = ~n144 & ~n405;
  assign n407 = ~n403 & ~n404;
  assign n408 = n406 & n407;
  assign n409 = n153 & n203;
  assign n410 = ~n378 & ~n409;
  assign n411 = ~n285 & ~n342;
  assign n412 = ~n362 & n411;
  assign n413 = ~n244 & ~n343;
  assign n414 = ~n391 & n413;
  assign n415 = n410 & n414;
  assign n416 = n394 & n408;
  assign n417 = n412 & n416;
  assign n418 = n402 & n415;
  assign n419 = n417 & n418;
  assign n420 = n176 & n211;
  assign n421 = ~n156 & ~n167;
  assign n422 = ~n420 & n421;
  assign n423 = n153 & n197;
  assign n424 = ~n113 & n423;
  assign n425 = ~n179 & ~n202;
  assign n426 = ~n236 & ~n424;
  assign n427 = n425 & n426;
  assign n428 = n422 & n427;
  assign n429 = n143 & n163;
  assign n430 = n164 & n173;
  assign n431 = ~n180 & ~n429;
  assign n432 = ~n430 & n431;
  assign n433 = n338 & n432;
  assign n434 = n176 & n178;
  assign n435 = ~n150 & ~n434;
  assign n436 = ~n352 & ~n355;
  assign n437 = n316 & n351;
  assign n438 = n436 & n437;
  assign n439 = ~n252 & ~n340;
  assign n440 = ~n212 & ~n233;
  assign n441 = ~n246 & ~n297;
  assign n442 = ~n299 & n441;
  assign n443 = n435 & n440;
  assign n444 = n439 & n443;
  assign n445 = n442 & n444;
  assign n446 = n438 & n445;
  assign n447 = ~n201 & ~n245;
  assign n448 = n446 & n447;
  assign n449 = ~n158 & ~n165;
  assign n450 = ~n113 & n242;
  assign n451 = ~n174 & ~n328;
  assign n452 = ~n450 & n451;
  assign n453 = n449 & n452;
  assign n454 = ~n291 & ~n319;
  assign n455 = n113 & n423;
  assign n456 = n128 & n203;
  assign n457 = ~n240 & ~n356;
  assign n458 = ~n455 & ~n456;
  assign n459 = n457 & n458;
  assign n460 = ~n234 & ~n292;
  assign n461 = ~n358 & n460;
  assign n462 = ~n230 & n454;
  assign n463 = n459 & n462;
  assign n464 = n461 & n463;
  assign n465 = n428 & n433;
  assign n466 = n453 & n465;
  assign n467 = n464 & n466;
  assign n468 = n419 & n467;
  assign n469 = n448 & n468;
  assign n470 = ~n390 & ~n469;
  assign n471 = ~pi22  & ~n80;
  assign n472 = pi9  & ~n471;
  assign n473 = ~pi9  & n471;
  assign n474 = ~n472 & ~n473;
  assign n475 = ~n113 & n403;
  assign n476 = ~n217 & ~n475;
  assign n477 = ~n434 & n476;
  assign n478 = n113 & n403;
  assign n479 = n154 & n176;
  assign n480 = n137 & n231;
  assign n481 = ~n479 & ~n480;
  assign n482 = ~n179 & ~n396;
  assign n483 = ~n150 & n482;
  assign n484 = ~n167 & ~n242;
  assign n485 = ~n245 & ~n478;
  assign n486 = n484 & n485;
  assign n487 = n481 & n486;
  assign n488 = n477 & n483;
  assign n489 = n487 & n488;
  assign n490 = ~n132 & ~n213;
  assign n491 = n145 & ~n490;
  assign n492 = n213 & n231;
  assign n493 = ~n362 & ~n492;
  assign n494 = ~n226 & ~n300;
  assign n495 = ~n334 & n494;
  assign n496 = n493 & n495;
  assign n497 = n154 & n213;
  assign n498 = ~n193 & ~n497;
  assign n499 = ~n271 & ~n303;
  assign n500 = ~n212 & ~n232;
  assign n501 = ~n339 & n500;
  assign n502 = ~n227 & ~n246;
  assign n503 = ~n332 & ~n420;
  assign n504 = n502 & n503;
  assign n505 = ~n168 & ~n272;
  assign n506 = n501 & n505;
  assign n507 = n504 & n506;
  assign n508 = ~n239 & ~n291;
  assign n509 = ~n199 & ~n267;
  assign n510 = ~n285 & n509;
  assign n511 = n351 & n508;
  assign n512 = n510 & n511;
  assign n513 = ~n240 & ~n296;
  assign n514 = n512 & n513;
  assign n515 = ~n194 & ~n299;
  assign n516 = ~n340 & ~n343;
  assign n517 = n515 & n516;
  assign n518 = n498 & n499;
  assign n519 = n517 & n518;
  assign n520 = n507 & n519;
  assign n521 = n514 & n520;
  assign n522 = n354 & ~n491;
  assign n523 = n496 & n522;
  assign n524 = n489 & n523;
  assign n525 = n521 & n524;
  assign n526 = ~n474 & ~n525;
  assign n527 = ~n470 & n526;
  assign n528 = pi10  & pi22 ;
  assign n529 = ~pi22  & ~n82;
  assign n530 = pi10  & ~n81;
  assign n531 = n529 & ~n530;
  assign n532 = ~n528 & ~n531;
  assign n533 = ~n525 & ~n532;
  assign n534 = n470 & ~n526;
  assign n535 = ~n527 & ~n534;
  assign n536 = n533 & n535;
  assign n537 = ~n527 & ~n536;
  assign n538 = ~n268 & ~n497;
  assign n539 = ~n214 & ~n233;
  assign n540 = ~n340 & ~n475;
  assign n541 = n539 & n540;
  assign n542 = n538 & n541;
  assign n543 = n288 & n542;
  assign n544 = ~n199 & ~n320;
  assign n545 = n543 & n544;
  assign n546 = n128 & n157;
  assign n547 = ~n424 & ~n546;
  assign n548 = n151 & n231;
  assign n549 = ~n237 & ~n548;
  assign n550 = n247 & ~n327;
  assign n551 = ~n180 & ~n303;
  assign n552 = ~n193 & ~n492;
  assign n553 = ~n266 & ~n273;
  assign n554 = ~n334 & ~n336;
  assign n555 = n553 & n554;
  assign n556 = n551 & n552;
  assign n557 = n555 & n556;
  assign n558 = ~n179 & ~n194;
  assign n559 = ~n430 & n558;
  assign n560 = ~n271 & ~n478;
  assign n561 = ~n212 & ~n290;
  assign n562 = n560 & n561;
  assign n563 = n109 & n143;
  assign n564 = ~n455 & ~n563;
  assign n565 = n141 & n155;
  assign n566 = n151 & n154;
  assign n567 = ~n142 & ~n255;
  assign n568 = ~n177 & ~n234;
  assign n569 = ~n152 & ~n299;
  assign n570 = ~n405 & ~n420;
  assign n571 = n569 & n570;
  assign n572 = n435 & n567;
  assign n573 = n568 & n572;
  assign n574 = n571 & n573;
  assign n575 = ~n156 & ~n253;
  assign n576 = ~n565 & ~n566;
  assign n577 = n575 & n576;
  assign n578 = n564 & n577;
  assign n579 = n559 & n562;
  assign n580 = n578 & n579;
  assign n581 = n574 & n580;
  assign n582 = n376 & n581;
  assign n583 = ~n230 & ~n404;
  assign n584 = n397 & n583;
  assign n585 = n547 & n549;
  assign n586 = n584 & n585;
  assign n587 = n550 & n586;
  assign n588 = n557 & n587;
  assign n589 = n545 & n588;
  assign n590 = n582 & n589;
  assign n591 = n469 & ~n590;
  assign n592 = ~n469 & n590;
  assign n593 = ~n591 & ~n592;
  assign n594 = n143 & n173;
  assign n595 = ~n229 & ~n594;
  assign n596 = ~n254 & ~n356;
  assign n597 = ~n327 & ~n563;
  assign n598 = n140 & n213;
  assign n599 = ~n142 & ~n598;
  assign n600 = ~n237 & n599;
  assign n601 = n359 & n596;
  assign n602 = n597 & n601;
  assign n603 = n160 & n600;
  assign n604 = n602 & n603;
  assign n605 = ~n202 & ~n219;
  assign n606 = ~n429 & n605;
  assign n607 = n604 & n606;
  assign n608 = ~n286 & ~n424;
  assign n609 = ~n244 & ~n292;
  assign n610 = ~n304 & ~n566;
  assign n611 = ~n266 & ~n320;
  assign n612 = ~n129 & ~n456;
  assign n613 = ~n204 & n612;
  assign n614 = ~n215 & ~n315;
  assign n615 = n613 & n614;
  assign n616 = n128 & n163;
  assign n617 = ~n236 & ~n252;
  assign n618 = ~n268 & ~n455;
  assign n619 = ~n616 & n618;
  assign n620 = n617 & n619;
  assign n621 = ~n548 & n608;
  assign n622 = n609 & n610;
  assign n623 = n611 & n622;
  assign n624 = n621 & n623;
  assign n625 = n615 & n620;
  assign n626 = n624 & n625;
  assign n627 = ~n200 & ~n289;
  assign n628 = n595 & n627;
  assign n629 = n607 & n628;
  assign n630 = n626 & n629;
  assign n631 = ~n593 & ~n630;
  assign n632 = pi14  & pi22 ;
  assign n633 = pi14  & ~n85;
  assign n634 = ~pi22  & ~n86;
  assign n635 = ~n633 & n634;
  assign n636 = ~n632 & ~n635;
  assign n637 = n631 & ~n636;
  assign n638 = ~n593 & n630;
  assign n639 = n636 & n638;
  assign n640 = ~pi22  & ~n84;
  assign n641 = pi13  & ~n640;
  assign n642 = ~pi13  & n640;
  assign n643 = ~n641 & ~n642;
  assign n644 = ~n590 & n630;
  assign n645 = n593 & ~n644;
  assign n646 = ~n643 & n645;
  assign n647 = ~n469 & ~n590;
  assign n648 = ~n630 & ~n647;
  assign n649 = n593 & ~n648;
  assign n650 = n643 & n649;
  assign n651 = ~n637 & ~n639;
  assign n652 = ~n646 & ~n650;
  assign n653 = n651 & n652;
  assign n654 = pi11  & ~n529;
  assign n655 = ~pi11  & n529;
  assign n656 = ~n654 & ~n655;
  assign n657 = n161 & n164;
  assign n658 = ~n337 & ~n657;
  assign n659 = ~n175 & ~n218;
  assign n660 = ~n377 & n659;
  assign n661 = n658 & n660;
  assign n662 = ~n133 & ~n201;
  assign n663 = ~n392 & n662;
  assign n664 = n661 & n663;
  assign n665 = ~n241 & n664;
  assign n666 = ~n177 & ~n347;
  assign n667 = ~n546 & n666;
  assign n668 = ~n290 & ~n430;
  assign n669 = ~n180 & ~n234;
  assign n670 = ~n273 & n669;
  assign n671 = n345 & n668;
  assign n672 = n670 & n671;
  assign n673 = n667 & n672;
  assign n674 = n159 & n596;
  assign n675 = n673 & n674;
  assign n676 = n626 & n675;
  assign n677 = n665 & n676;
  assign n678 = n630 & ~n677;
  assign n679 = ~n630 & n677;
  assign n680 = ~n678 & ~n679;
  assign n681 = n525 & ~n630;
  assign n682 = n680 & ~n681;
  assign n683 = ~n656 & n682;
  assign n684 = pi12  & pi22 ;
  assign n685 = pi12  & ~n83;
  assign n686 = n640 & ~n685;
  assign n687 = ~n684 & ~n686;
  assign n688 = ~n525 & ~n687;
  assign n689 = n525 & n687;
  assign n690 = ~n688 & ~n689;
  assign n691 = ~n680 & ~n690;
  assign n692 = ~n630 & ~n677;
  assign n693 = ~n525 & ~n692;
  assign n694 = n680 & ~n693;
  assign n695 = n656 & n694;
  assign n696 = ~n683 & ~n691;
  assign n697 = ~n695 & n696;
  assign n698 = n653 & n697;
  assign n699 = n283 & ~n389;
  assign n700 = ~n283 & n389;
  assign n701 = ~n699 & ~n700;
  assign n702 = ~n636 & n701;
  assign n703 = ~n470 & ~n702;
  assign n704 = ~n389 & n469;
  assign n705 = n701 & ~n704;
  assign n706 = ~n636 & n705;
  assign n707 = ~n703 & ~n706;
  assign n708 = ~n526 & n707;
  assign n709 = n526 & ~n707;
  assign n710 = ~n708 & ~n709;
  assign n711 = n631 & ~n643;
  assign n712 = n638 & n643;
  assign n713 = n645 & ~n687;
  assign n714 = n649 & n687;
  assign n715 = ~n711 & ~n712;
  assign n716 = ~n713 & ~n714;
  assign n717 = n715 & n716;
  assign n718 = n710 & n717;
  assign n719 = ~n708 & ~n718;
  assign n720 = ~n653 & ~n697;
  assign n721 = ~n698 & ~n720;
  assign n722 = ~n719 & n721;
  assign n723 = ~n698 & ~n722;
  assign n724 = ~n537 & ~n723;
  assign n725 = ~n537 & n723;
  assign n726 = n537 & ~n723;
  assign n727 = ~n725 & ~n726;
  assign n728 = ~n525 & ~n656;
  assign n729 = n593 & ~n636;
  assign n730 = ~n648 & ~n729;
  assign n731 = ~n636 & n645;
  assign n732 = ~n730 & ~n731;
  assign n733 = ~n728 & n732;
  assign n734 = n728 & ~n732;
  assign n735 = ~n733 & ~n734;
  assign n736 = n682 & ~n687;
  assign n737 = ~n525 & ~n643;
  assign n738 = n525 & n643;
  assign n739 = ~n737 & ~n738;
  assign n740 = ~n680 & ~n739;
  assign n741 = n687 & n694;
  assign n742 = ~n736 & ~n740;
  assign n743 = ~n741 & n742;
  assign n744 = n735 & n743;
  assign n745 = ~n735 & ~n743;
  assign n746 = ~n744 & ~n745;
  assign n747 = ~n727 & n746;
  assign n748 = ~n724 & ~n747;
  assign n749 = ~n733 & ~n744;
  assign n750 = ~n643 & n682;
  assign n751 = n643 & n694;
  assign n752 = n525 & ~n636;
  assign n753 = ~n525 & n636;
  assign n754 = ~n752 & ~n753;
  assign n755 = ~n680 & n754;
  assign n756 = ~n750 & ~n755;
  assign n757 = ~n751 & n756;
  assign n758 = ~n749 & n757;
  assign n759 = n749 & ~n757;
  assign n760 = ~n758 & ~n759;
  assign n761 = ~n648 & n728;
  assign n762 = n648 & ~n728;
  assign n763 = ~n761 & ~n762;
  assign n764 = n688 & n763;
  assign n765 = ~n688 & ~n763;
  assign n766 = ~n764 & ~n765;
  assign n767 = n760 & n766;
  assign n768 = ~n760 & ~n766;
  assign n769 = ~n767 & ~n768;
  assign n770 = ~n748 & n769;
  assign n771 = ~pi22  & ~n78;
  assign n772 = pi7  & ~n771;
  assign n773 = ~pi7  & n771;
  assign n774 = ~n772 & ~n773;
  assign n775 = ~n525 & ~n774;
  assign n776 = ~n286 & ~n292;
  assign n777 = n595 & n776;
  assign n778 = ~n165 & ~n285;
  assign n779 = ~n319 & ~n404;
  assign n780 = n778 & n779;
  assign n781 = n501 & n780;
  assign n782 = ~n150 & ~n480;
  assign n783 = ~n199 & ~n241;
  assign n784 = ~n332 & n783;
  assign n785 = n551 & n782;
  assign n786 = n784 & n785;
  assign n787 = n394 & n777;
  assign n788 = n786 & n787;
  assign n789 = n781 & n788;
  assign n790 = ~n174 & ~n272;
  assign n791 = ~n352 & n790;
  assign n792 = ~n204 & ~n566;
  assign n793 = ~n144 & ~n230;
  assign n794 = ~n378 & n793;
  assign n795 = n439 & n792;
  assign n796 = n794 & n795;
  assign n797 = ~n218 & ~n430;
  assign n798 = ~n343 & ~n360;
  assign n799 = ~n479 & n798;
  assign n800 = ~n236 & ~n475;
  assign n801 = ~n217 & ~n492;
  assign n802 = n797 & n800;
  assign n803 = n801 & n802;
  assign n804 = n799 & n803;
  assign n805 = ~n202 & ~n396;
  assign n806 = n196 & ~n243;
  assign n807 = n805 & n806;
  assign n808 = ~n273 & ~n304;
  assign n809 = ~n138 & ~n175;
  assign n810 = ~n291 & ~n336;
  assign n811 = ~n350 & ~n355;
  assign n812 = n810 & n811;
  assign n813 = n808 & n809;
  assign n814 = n812 & n813;
  assign n815 = n796 & n814;
  assign n816 = n807 & n815;
  assign n817 = n804 & n816;
  assign n818 = n113 & n215;
  assign n819 = ~n342 & ~n818;
  assign n820 = ~n172 & n819;
  assign n821 = ~n266 & ~n391;
  assign n822 = n141 & n151;
  assign n823 = ~n168 & ~n822;
  assign n824 = ~n162 & ~n240;
  assign n825 = ~n254 & ~n271;
  assign n826 = ~n297 & ~n450;
  assign n827 = ~n563 & n826;
  assign n828 = n824 & n825;
  assign n829 = n827 & n828;
  assign n830 = ~n317 & ~n497;
  assign n831 = n658 & n830;
  assign n832 = n821 & n823;
  assign n833 = n831 & n832;
  assign n834 = n422 & n791;
  assign n835 = n820 & n834;
  assign n836 = n829 & n833;
  assign n837 = n835 & n836;
  assign n838 = n789 & n837;
  assign n839 = n817 & n838;
  assign n840 = ~n480 & ~n566;
  assign n841 = ~n232 & ~n297;
  assign n842 = ~n200 & n841;
  assign n843 = ~n214 & ~n429;
  assign n844 = ~n218 & ~n340;
  assign n845 = n840 & n844;
  assign n846 = n843 & n845;
  assign n847 = n842 & n846;
  assign n848 = ~n347 & ~n392;
  assign n849 = ~n216 & ~n290;
  assign n850 = ~n424 & n849;
  assign n851 = ~n201 & ~n240;
  assign n852 = ~n243 & ~n352;
  assign n853 = n851 & n852;
  assign n854 = n848 & n853;
  assign n855 = n850 & n854;
  assign n856 = ~n273 & ~n818;
  assign n857 = ~n396 & n856;
  assign n858 = ~n156 & ~n220;
  assign n859 = n857 & n858;
  assign n860 = ~n179 & ~n334;
  assign n861 = ~n194 & ~n227;
  assign n862 = ~n245 & ~n296;
  assign n863 = ~n342 & n862;
  assign n864 = n861 & n863;
  assign n865 = ~n300 & ~n336;
  assign n866 = ~n343 & ~n456;
  assign n867 = n865 & n866;
  assign n868 = ~n284 & ~n289;
  assign n869 = ~n420 & n868;
  assign n870 = n329 & n395;
  assign n871 = n538 & n870;
  assign n872 = n777 & n869;
  assign n873 = n867 & n872;
  assign n874 = n864 & n871;
  assign n875 = n873 & n874;
  assign n876 = ~n174 & ~n230;
  assign n877 = n860 & n876;
  assign n878 = n875 & n877;
  assign n879 = ~n180 & ~n332;
  assign n880 = ~n404 & n879;
  assign n881 = n435 & n880;
  assign n882 = n366 & n881;
  assign n883 = n859 & n882;
  assign n884 = n847 & n855;
  assign n885 = n883 & n884;
  assign n886 = n878 & n885;
  assign n887 = ~n839 & ~n886;
  assign n888 = ~n283 & ~n887;
  assign n889 = n775 & ~n888;
  assign n890 = ~n775 & n888;
  assign n891 = ~n889 & ~n890;
  assign n892 = pi8  & pi22 ;
  assign n893 = pi8  & ~n79;
  assign n894 = n471 & ~n893;
  assign n895 = ~n892 & ~n894;
  assign n896 = ~n525 & ~n895;
  assign n897 = n891 & n896;
  assign n898 = ~n889 & ~n897;
  assign n899 = ~n532 & n682;
  assign n900 = n525 & n656;
  assign n901 = ~n728 & ~n900;
  assign n902 = ~n680 & ~n901;
  assign n903 = n532 & n694;
  assign n904 = ~n899 & ~n902;
  assign n905 = ~n903 & n904;
  assign n906 = ~n898 & n905;
  assign n907 = n469 & ~n701;
  assign n908 = n636 & n907;
  assign n909 = ~n643 & n705;
  assign n910 = ~n469 & ~n701;
  assign n911 = ~n636 & n910;
  assign n912 = ~n470 & n701;
  assign n913 = n643 & n912;
  assign n914 = ~n908 & ~n909;
  assign n915 = ~n911 & ~n913;
  assign n916 = n914 & n915;
  assign n917 = n631 & ~n687;
  assign n918 = n638 & n687;
  assign n919 = n645 & ~n656;
  assign n920 = n649 & n656;
  assign n921 = ~n917 & ~n918;
  assign n922 = ~n919 & ~n920;
  assign n923 = n921 & n922;
  assign n924 = n916 & ~n923;
  assign n925 = ~n916 & n923;
  assign n926 = ~n924 & ~n925;
  assign n927 = ~n474 & n682;
  assign n928 = n525 & n532;
  assign n929 = ~n533 & ~n928;
  assign n930 = ~n680 & ~n929;
  assign n931 = n474 & n694;
  assign n932 = ~n927 & ~n930;
  assign n933 = ~n931 & n932;
  assign n934 = ~n926 & n933;
  assign n935 = n916 & n923;
  assign n936 = ~n934 & ~n935;
  assign n937 = n898 & ~n905;
  assign n938 = ~n906 & ~n937;
  assign n939 = ~n936 & n938;
  assign n940 = ~n906 & ~n939;
  assign n941 = ~n533 & ~n535;
  assign n942 = ~n536 & ~n941;
  assign n943 = ~n940 & n942;
  assign n944 = n940 & ~n942;
  assign n945 = ~n943 & ~n944;
  assign n946 = n719 & ~n721;
  assign n947 = ~n722 & ~n946;
  assign n948 = n945 & n947;
  assign n949 = ~n943 & ~n948;
  assign n950 = ~n727 & ~n746;
  assign n951 = n727 & n746;
  assign n952 = ~n950 & ~n951;
  assign n953 = ~n949 & ~n952;
  assign n954 = n631 & ~n656;
  assign n955 = n638 & n656;
  assign n956 = ~n532 & n645;
  assign n957 = n532 & n649;
  assign n958 = ~n954 & ~n955;
  assign n959 = ~n956 & ~n957;
  assign n960 = n958 & n959;
  assign n961 = n682 & ~n895;
  assign n962 = n474 & n525;
  assign n963 = ~n526 & ~n962;
  assign n964 = ~n680 & ~n963;
  assign n965 = n694 & n895;
  assign n966 = ~n961 & ~n964;
  assign n967 = ~n965 & n966;
  assign n968 = n960 & n967;
  assign n969 = ~n960 & ~n967;
  assign n970 = ~n968 & ~n969;
  assign n971 = ~n240 & ~n594;
  assign n972 = ~n138 & ~n195;
  assign n973 = ~n377 & n972;
  assign n974 = n499 & n608;
  assign n975 = n971 & n974;
  assign n976 = n973 & n975;
  assign n977 = ~n289 & ~n565;
  assign n978 = ~n337 & ~n616;
  assign n979 = ~n172 & ~n242;
  assign n980 = ~n215 & n978;
  assign n981 = n979 & n980;
  assign n982 = ~n180 & ~n237;
  assign n983 = ~n334 & ~n455;
  assign n984 = n982 & n983;
  assign n985 = ~n175 & ~n244;
  assign n986 = ~n657 & n985;
  assign n987 = ~n328 & ~n391;
  assign n988 = ~n566 & n987;
  assign n989 = ~n236 & ~n336;
  assign n990 = ~n429 & ~n480;
  assign n991 = n989 & n990;
  assign n992 = n316 & n991;
  assign n993 = n984 & n986;
  assign n994 = n988 & n993;
  assign n995 = n864 & n992;
  assign n996 = n994 & n995;
  assign n997 = ~n129 & ~n156;
  assign n998 = ~n212 & ~n234;
  assign n999 = ~n332 & ~n378;
  assign n1000 = n998 & n999;
  assign n1001 = n318 & n997;
  assign n1002 = n397 & n808;
  assign n1003 = n1001 & n1002;
  assign n1004 = n1000 & n1003;
  assign n1005 = ~n339 & ~n434;
  assign n1006 = ~n133 & ~n204;
  assign n1007 = ~n230 & ~n239;
  assign n1008 = ~n297 & n1007;
  assign n1009 = n361 & n1006;
  assign n1010 = n823 & n977;
  assign n1011 = n1005 & n1010;
  assign n1012 = n1008 & n1009;
  assign n1013 = n408 & n1012;
  assign n1014 = n981 & n1011;
  assign n1015 = n1013 & n1014;
  assign n1016 = n976 & n1004;
  assign n1017 = n1015 & n1016;
  assign n1018 = n996 & n1017;
  assign n1019 = n839 & n1018;
  assign n1020 = pi6  & pi22 ;
  assign n1021 = pi6  & ~n77;
  assign n1022 = n771 & ~n1021;
  assign n1023 = ~n1020 & ~n1022;
  assign n1024 = ~n525 & ~n1023;
  assign n1025 = ~n290 & ~n336;
  assign n1026 = ~n342 & ~n420;
  assign n1027 = n335 & n1026;
  assign n1028 = n611 & n977;
  assign n1029 = n1027 & n1028;
  assign n1030 = ~n218 & ~n343;
  assign n1031 = ~n346 & ~n348;
  assign n1032 = ~n548 & n1031;
  assign n1033 = n476 & n1030;
  assign n1034 = n1025 & n1033;
  assign n1035 = n550 & n1032;
  assign n1036 = n791 & n1035;
  assign n1037 = n981 & n1034;
  assign n1038 = n1029 & n1037;
  assign n1039 = n1036 & n1038;
  assign n1040 = ~n201 & ~n347;
  assign n1041 = ~n358 & ~n377;
  assign n1042 = n1040 & n1041;
  assign n1043 = n547 & n1042;
  assign n1044 = ~n162 & ~n230;
  assign n1045 = ~n244 & ~n271;
  assign n1046 = ~n332 & ~n353;
  assign n1047 = n1045 & n1046;
  assign n1048 = n552 & n1044;
  assign n1049 = n805 & n1048;
  assign n1050 = n1047 & n1049;
  assign n1051 = ~n167 & ~n195;
  assign n1052 = ~n255 & ~n317;
  assign n1053 = ~n339 & ~n355;
  assign n1054 = ~n822 & n1053;
  assign n1055 = n1051 & n1052;
  assign n1056 = n159 & n410;
  assign n1057 = n1055 & n1056;
  assign n1058 = n842 & n1054;
  assign n1059 = n1057 & n1058;
  assign n1060 = n1050 & n1059;
  assign n1061 = ~n227 & ~n252;
  assign n1062 = ~n304 & ~n478;
  assign n1063 = n1061 & n1062;
  assign n1064 = ~n199 & ~n350;
  assign n1065 = ~n657 & n1064;
  assign n1066 = n238 & n345;
  assign n1067 = n435 & n1066;
  assign n1068 = n613 & n1065;
  assign n1069 = n1063 & n1068;
  assign n1070 = n1043 & n1067;
  assign n1071 = n1069 & n1070;
  assign n1072 = n1060 & n1071;
  assign n1073 = n1039 & n1072;
  assign n1074 = ~n1018 & n1073;
  assign n1075 = ~n839 & n1074;
  assign n1076 = n1024 & ~n1075;
  assign n1077 = ~n1019 & ~n1076;
  assign n1078 = n970 & ~n1077;
  assign n1079 = ~n968 & ~n1078;
  assign n1080 = n839 & ~n886;
  assign n1081 = ~n839 & n886;
  assign n1082 = ~n1080 & ~n1081;
  assign n1083 = ~n636 & n1082;
  assign n1084 = ~n888 & ~n1083;
  assign n1085 = n839 & n886;
  assign n1086 = n283 & ~n1085;
  assign n1087 = n1083 & ~n1086;
  assign n1088 = ~n1084 & ~n1087;
  assign n1089 = ~n775 & n1088;
  assign n1090 = n775 & ~n1088;
  assign n1091 = ~n1089 & ~n1090;
  assign n1092 = n643 & n907;
  assign n1093 = ~n687 & n705;
  assign n1094 = ~n643 & n910;
  assign n1095 = n687 & n912;
  assign n1096 = ~n1092 & ~n1093;
  assign n1097 = ~n1094 & ~n1095;
  assign n1098 = n1096 & n1097;
  assign n1099 = n1091 & n1098;
  assign n1100 = ~n1089 & ~n1099;
  assign n1101 = ~n1079 & ~n1100;
  assign n1102 = ~n1079 & n1100;
  assign n1103 = n1079 & ~n1100;
  assign n1104 = ~n1102 & ~n1103;
  assign n1105 = ~n891 & ~n896;
  assign n1106 = ~n897 & ~n1105;
  assign n1107 = ~n1104 & n1106;
  assign n1108 = ~n1101 & ~n1107;
  assign n1109 = ~n710 & ~n717;
  assign n1110 = ~n718 & ~n1109;
  assign n1111 = ~n1108 & n1110;
  assign n1112 = n1108 & ~n1110;
  assign n1113 = ~n1111 & ~n1112;
  assign n1114 = n936 & ~n938;
  assign n1115 = ~n939 & ~n1114;
  assign n1116 = n1113 & n1115;
  assign n1117 = ~n1111 & ~n1116;
  assign n1118 = ~n945 & ~n947;
  assign n1119 = ~n948 & ~n1118;
  assign n1120 = ~n1117 & n1119;
  assign n1121 = ~n1113 & ~n1115;
  assign n1122 = ~n1116 & ~n1121;
  assign n1123 = ~n532 & n631;
  assign n1124 = n532 & n638;
  assign n1125 = ~n474 & n645;
  assign n1126 = n474 & n649;
  assign n1127 = ~n1123 & ~n1124;
  assign n1128 = ~n1125 & ~n1126;
  assign n1129 = n1127 & n1128;
  assign n1130 = n682 & ~n774;
  assign n1131 = n525 & n895;
  assign n1132 = ~n896 & ~n1131;
  assign n1133 = ~n680 & ~n1132;
  assign n1134 = n694 & n774;
  assign n1135 = ~n1130 & ~n1133;
  assign n1136 = ~n1134 & n1135;
  assign n1137 = n1129 & ~n1136;
  assign n1138 = ~n1129 & n1136;
  assign n1139 = ~n1137 & ~n1138;
  assign n1140 = ~n283 & ~n1082;
  assign n1141 = ~n636 & n1140;
  assign n1142 = n283 & ~n1082;
  assign n1143 = n636 & n1142;
  assign n1144 = n1082 & ~n1086;
  assign n1145 = ~n643 & n1144;
  assign n1146 = ~n888 & n1082;
  assign n1147 = n643 & n1146;
  assign n1148 = ~n1141 & ~n1143;
  assign n1149 = ~n1145 & ~n1147;
  assign n1150 = n1148 & n1149;
  assign n1151 = ~n1139 & n1150;
  assign n1152 = n1129 & n1136;
  assign n1153 = ~n1151 & ~n1152;
  assign n1154 = ~n1091 & ~n1098;
  assign n1155 = ~n1099 & ~n1154;
  assign n1156 = ~n1153 & n1155;
  assign n1157 = ~n970 & n1077;
  assign n1158 = ~n1078 & ~n1157;
  assign n1159 = n1153 & ~n1155;
  assign n1160 = ~n1156 & ~n1159;
  assign n1161 = n1158 & n1160;
  assign n1162 = ~n1156 & ~n1161;
  assign n1163 = n926 & n933;
  assign n1164 = ~n926 & ~n933;
  assign n1165 = ~n1163 & ~n1164;
  assign n1166 = n1162 & n1165;
  assign n1167 = ~n1162 & ~n1165;
  assign n1168 = ~n1104 & ~n1106;
  assign n1169 = n1104 & n1106;
  assign n1170 = ~n1168 & ~n1169;
  assign n1171 = ~n1167 & n1170;
  assign n1172 = ~n1166 & ~n1171;
  assign n1173 = n1122 & n1172;
  assign n1174 = n687 & n907;
  assign n1175 = ~n656 & n705;
  assign n1176 = ~n687 & n910;
  assign n1177 = n656 & n912;
  assign n1178 = ~n1174 & ~n1175;
  assign n1179 = ~n1176 & ~n1177;
  assign n1180 = n1178 & n1179;
  assign n1181 = ~n1019 & ~n1075;
  assign n1182 = n1024 & ~n1181;
  assign n1183 = ~n1076 & n1181;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = n1180 & ~n1184;
  assign n1186 = ~n57 & ~n525;
  assign n1187 = ~n1018 & n1186;
  assign n1188 = n1018 & ~n1186;
  assign n1189 = ~n1187 & ~n1188;
  assign n1190 = ~n1018 & ~n1073;
  assign n1191 = ~n839 & ~n1190;
  assign n1192 = n1018 & ~n1073;
  assign n1193 = ~n1074 & ~n1192;
  assign n1194 = ~n636 & n1193;
  assign n1195 = ~n1191 & ~n1194;
  assign n1196 = n1018 & n1073;
  assign n1197 = n839 & ~n1196;
  assign n1198 = n1194 & ~n1197;
  assign n1199 = ~n1195 & ~n1198;
  assign n1200 = n1189 & n1199;
  assign n1201 = ~n1187 & ~n1200;
  assign n1202 = ~n1180 & n1184;
  assign n1203 = ~n1185 & ~n1202;
  assign n1204 = ~n1201 & n1203;
  assign n1205 = ~n1185 & ~n1204;
  assign n1206 = ~n643 & n1140;
  assign n1207 = n643 & n1142;
  assign n1208 = ~n687 & n1144;
  assign n1209 = n687 & n1146;
  assign n1210 = ~n1206 & ~n1207;
  assign n1211 = ~n1208 & ~n1209;
  assign n1212 = n1210 & n1211;
  assign n1213 = n656 & n907;
  assign n1214 = ~n532 & n705;
  assign n1215 = ~n656 & n910;
  assign n1216 = n532 & n912;
  assign n1217 = ~n1213 & ~n1214;
  assign n1218 = ~n1215 & ~n1216;
  assign n1219 = n1217 & n1218;
  assign n1220 = n1212 & n1219;
  assign n1221 = n1212 & ~n1219;
  assign n1222 = ~n1212 & n1219;
  assign n1223 = ~n1221 & ~n1222;
  assign n1224 = ~n474 & n631;
  assign n1225 = n474 & n638;
  assign n1226 = n645 & ~n895;
  assign n1227 = n649 & n895;
  assign n1228 = ~n1224 & ~n1225;
  assign n1229 = ~n1226 & ~n1227;
  assign n1230 = n1228 & n1229;
  assign n1231 = ~n1223 & n1230;
  assign n1232 = ~n1220 & ~n1231;
  assign n1233 = n1139 & ~n1150;
  assign n1234 = ~n1151 & ~n1233;
  assign n1235 = ~n1232 & n1234;
  assign n1236 = ~n72 & ~n525;
  assign n1237 = ~n1018 & n1236;
  assign n1238 = n1018 & ~n1236;
  assign n1239 = ~n1237 & ~n1238;
  assign n1240 = ~n839 & ~n1193;
  assign n1241 = ~n636 & n1240;
  assign n1242 = n839 & ~n1193;
  assign n1243 = n636 & n1242;
  assign n1244 = n1193 & ~n1197;
  assign n1245 = ~n643 & n1244;
  assign n1246 = ~n1191 & n1193;
  assign n1247 = n643 & n1246;
  assign n1248 = ~n1241 & ~n1243;
  assign n1249 = ~n1245 & ~n1247;
  assign n1250 = n1248 & n1249;
  assign n1251 = n1239 & n1250;
  assign n1252 = ~n1237 & ~n1251;
  assign n1253 = n682 & ~n1023;
  assign n1254 = n525 & n774;
  assign n1255 = ~n775 & ~n1254;
  assign n1256 = ~n680 & ~n1255;
  assign n1257 = n694 & n1023;
  assign n1258 = ~n1253 & ~n1256;
  assign n1259 = ~n1257 & n1258;
  assign n1260 = ~n1252 & n1259;
  assign n1261 = n1252 & ~n1259;
  assign n1262 = ~n1260 & ~n1261;
  assign n1263 = n532 & n907;
  assign n1264 = ~n474 & n705;
  assign n1265 = ~n532 & n910;
  assign n1266 = n474 & n912;
  assign n1267 = ~n1263 & ~n1264;
  assign n1268 = ~n1265 & ~n1266;
  assign n1269 = n1267 & n1268;
  assign n1270 = ~n687 & n1140;
  assign n1271 = n687 & n1142;
  assign n1272 = ~n656 & n1144;
  assign n1273 = n656 & n1146;
  assign n1274 = ~n1270 & ~n1271;
  assign n1275 = ~n1272 & ~n1273;
  assign n1276 = n1274 & n1275;
  assign n1277 = n1269 & n1276;
  assign n1278 = ~n1269 & n1276;
  assign n1279 = n1269 & ~n1276;
  assign n1280 = ~n1278 & ~n1279;
  assign n1281 = n631 & ~n895;
  assign n1282 = n638 & n895;
  assign n1283 = n645 & ~n774;
  assign n1284 = n649 & n774;
  assign n1285 = ~n1281 & ~n1282;
  assign n1286 = ~n1283 & ~n1284;
  assign n1287 = n1285 & n1286;
  assign n1288 = ~n1280 & n1287;
  assign n1289 = ~n1277 & ~n1288;
  assign n1290 = n1262 & ~n1289;
  assign n1291 = ~n1260 & ~n1290;
  assign n1292 = n1232 & ~n1234;
  assign n1293 = ~n1235 & ~n1292;
  assign n1294 = ~n1291 & n1293;
  assign n1295 = ~n1235 & ~n1294;
  assign n1296 = ~n1205 & ~n1295;
  assign n1297 = ~n1205 & n1295;
  assign n1298 = n1205 & ~n1295;
  assign n1299 = ~n1297 & ~n1298;
  assign n1300 = ~n1158 & ~n1160;
  assign n1301 = ~n1161 & ~n1300;
  assign n1302 = ~n1299 & n1301;
  assign n1303 = ~n1296 & ~n1302;
  assign n1304 = ~n1166 & ~n1167;
  assign n1305 = n1170 & n1304;
  assign n1306 = ~n1170 & ~n1304;
  assign n1307 = ~n1305 & ~n1306;
  assign n1308 = ~n1303 & ~n1307;
  assign n1309 = ~n1299 & ~n1301;
  assign n1310 = n1299 & n1301;
  assign n1311 = ~n1309 & ~n1310;
  assign n1312 = n1223 & n1230;
  assign n1313 = ~n1223 & ~n1230;
  assign n1314 = ~n1312 & ~n1313;
  assign n1315 = ~n1189 & ~n1199;
  assign n1316 = ~n1200 & ~n1315;
  assign n1317 = ~n1314 & n1316;
  assign n1318 = n1314 & n1316;
  assign n1319 = ~n1314 & ~n1316;
  assign n1320 = ~n1318 & ~n1319;
  assign n1321 = ~n61 & ~n525;
  assign n1322 = ~n317 & ~n546;
  assign n1323 = ~n218 & ~n243;
  assign n1324 = ~n420 & n1323;
  assign n1325 = ~n179 & ~n271;
  assign n1326 = ~n296 & ~n392;
  assign n1327 = ~n404 & n1326;
  assign n1328 = n354 & n1325;
  assign n1329 = n549 & n841;
  assign n1330 = n1328 & n1329;
  assign n1331 = n459 & n1327;
  assign n1332 = n1324 & n1331;
  assign n1333 = n1330 & n1332;
  assign n1334 = ~n168 & ~n230;
  assign n1335 = ~n292 & ~n396;
  assign n1336 = n1334 & n1335;
  assign n1337 = n321 & n800;
  assign n1338 = n821 & n1337;
  assign n1339 = n1336 & n1338;
  assign n1340 = ~n152 & ~n165;
  assign n1341 = ~n180 & ~n355;
  assign n1342 = ~n358 & ~n424;
  assign n1343 = ~n563 & ~n566;
  assign n1344 = ~n822 & n1343;
  assign n1345 = n1341 & n1342;
  assign n1346 = n1340 & n1345;
  assign n1347 = n1344 & n1346;
  assign n1348 = ~n253 & ~n300;
  assign n1349 = ~n337 & ~n478;
  assign n1350 = ~n565 & n1349;
  assign n1351 = n567 & n1348;
  assign n1352 = n1322 & n1351;
  assign n1353 = n1350 & n1352;
  assign n1354 = n512 & n1353;
  assign n1355 = n1339 & n1347;
  assign n1356 = n1354 & n1355;
  assign n1357 = n1333 & n1356;
  assign n1358 = ~n1018 & ~n1357;
  assign n1359 = n636 & ~n1018;
  assign n1360 = ~n1358 & ~n1359;
  assign n1361 = n1321 & ~n1360;
  assign n1362 = ~n1321 & n1360;
  assign n1363 = ~n1361 & ~n1362;
  assign n1364 = ~n643 & n1240;
  assign n1365 = n643 & n1242;
  assign n1366 = ~n687 & n1244;
  assign n1367 = n687 & n1246;
  assign n1368 = ~n1364 & ~n1365;
  assign n1369 = ~n1366 & ~n1367;
  assign n1370 = n1368 & n1369;
  assign n1371 = n1363 & n1370;
  assign n1372 = ~n1361 & ~n1371;
  assign n1373 = ~n57 & n682;
  assign n1374 = n525 & n1023;
  assign n1375 = ~n1024 & ~n1374;
  assign n1376 = ~n680 & ~n1375;
  assign n1377 = n57 & n694;
  assign n1378 = ~n1373 & ~n1376;
  assign n1379 = ~n1377 & n1378;
  assign n1380 = ~n1372 & n1379;
  assign n1381 = n1372 & ~n1379;
  assign n1382 = ~n1380 & ~n1381;
  assign n1383 = n474 & n907;
  assign n1384 = n705 & ~n895;
  assign n1385 = ~n474 & n910;
  assign n1386 = n895 & n912;
  assign n1387 = ~n1383 & ~n1384;
  assign n1388 = ~n1385 & ~n1386;
  assign n1389 = n1387 & n1388;
  assign n1390 = ~n656 & n1140;
  assign n1391 = n656 & n1142;
  assign n1392 = ~n532 & n1144;
  assign n1393 = n532 & n1146;
  assign n1394 = ~n1390 & ~n1391;
  assign n1395 = ~n1392 & ~n1393;
  assign n1396 = n1394 & n1395;
  assign n1397 = n1389 & n1396;
  assign n1398 = ~n1389 & n1396;
  assign n1399 = n1389 & ~n1396;
  assign n1400 = ~n1398 & ~n1399;
  assign n1401 = n631 & ~n774;
  assign n1402 = n638 & n774;
  assign n1403 = n645 & ~n1023;
  assign n1404 = n649 & n1023;
  assign n1405 = ~n1401 & ~n1402;
  assign n1406 = ~n1403 & ~n1404;
  assign n1407 = n1405 & n1406;
  assign n1408 = ~n1400 & n1407;
  assign n1409 = ~n1397 & ~n1408;
  assign n1410 = n1382 & ~n1409;
  assign n1411 = ~n1380 & ~n1410;
  assign n1412 = ~n1320 & ~n1411;
  assign n1413 = ~n1317 & ~n1412;
  assign n1414 = n1201 & ~n1203;
  assign n1415 = ~n1204 & ~n1414;
  assign n1416 = ~n1413 & n1415;
  assign n1417 = n1413 & ~n1415;
  assign n1418 = ~n1416 & ~n1417;
  assign n1419 = n1291 & ~n1293;
  assign n1420 = ~n1294 & ~n1419;
  assign n1421 = n1418 & n1420;
  assign n1422 = ~n1416 & ~n1421;
  assign n1423 = ~n1311 & ~n1422;
  assign n1424 = ~n61 & ~n680;
  assign n1425 = n693 & ~n1424;
  assign n1426 = ~n636 & n1358;
  assign n1427 = ~n643 & n1357;
  assign n1428 = ~n636 & ~n1357;
  assign n1429 = n1018 & ~n1428;
  assign n1430 = ~n1426 & ~n1427;
  assign n1431 = ~n1429 & n1430;
  assign n1432 = n1425 & n1431;
  assign n1433 = ~n72 & n682;
  assign n1434 = n57 & n525;
  assign n1435 = ~n1186 & ~n1434;
  assign n1436 = ~n680 & ~n1435;
  assign n1437 = n72 & n694;
  assign n1438 = ~n1433 & ~n1436;
  assign n1439 = ~n1437 & n1438;
  assign n1440 = n1432 & n1439;
  assign n1441 = n895 & n907;
  assign n1442 = n705 & ~n774;
  assign n1443 = ~n895 & n910;
  assign n1444 = n774 & n912;
  assign n1445 = ~n1441 & ~n1442;
  assign n1446 = ~n1443 & ~n1444;
  assign n1447 = n1445 & n1446;
  assign n1448 = n631 & ~n1023;
  assign n1449 = n638 & n1023;
  assign n1450 = ~n57 & n645;
  assign n1451 = n57 & n649;
  assign n1452 = ~n1448 & ~n1449;
  assign n1453 = ~n1450 & ~n1451;
  assign n1454 = n1452 & n1453;
  assign n1455 = n1447 & ~n1454;
  assign n1456 = ~n1447 & n1454;
  assign n1457 = ~n1455 & ~n1456;
  assign n1458 = ~n532 & n1140;
  assign n1459 = n532 & n1142;
  assign n1460 = ~n474 & n1144;
  assign n1461 = n474 & n1146;
  assign n1462 = ~n1458 & ~n1459;
  assign n1463 = ~n1460 & ~n1461;
  assign n1464 = n1462 & n1463;
  assign n1465 = ~n1457 & n1464;
  assign n1466 = n1447 & n1454;
  assign n1467 = ~n1465 & ~n1466;
  assign n1468 = ~n1432 & ~n1439;
  assign n1469 = ~n1440 & ~n1468;
  assign n1470 = ~n1467 & n1469;
  assign n1471 = ~n1440 & ~n1470;
  assign n1472 = ~n1239 & ~n1250;
  assign n1473 = ~n1251 & ~n1472;
  assign n1474 = ~n1471 & n1473;
  assign n1475 = n1280 & n1287;
  assign n1476 = ~n1280 & ~n1287;
  assign n1477 = ~n1475 & ~n1476;
  assign n1478 = n1471 & ~n1473;
  assign n1479 = ~n1474 & ~n1478;
  assign n1480 = ~n1477 & n1479;
  assign n1481 = ~n1474 & ~n1480;
  assign n1482 = ~n1262 & n1289;
  assign n1483 = ~n1290 & ~n1482;
  assign n1484 = ~n1481 & n1483;
  assign n1485 = n1320 & ~n1411;
  assign n1486 = ~n1320 & n1411;
  assign n1487 = ~n1485 & ~n1486;
  assign n1488 = n1481 & ~n1483;
  assign n1489 = ~n1484 & ~n1488;
  assign n1490 = ~n1487 & n1489;
  assign n1491 = ~n1484 & ~n1490;
  assign n1492 = ~n1418 & ~n1420;
  assign n1493 = ~n1421 & ~n1492;
  assign n1494 = ~n1491 & n1493;
  assign n1495 = ~n1382 & n1409;
  assign n1496 = ~n1410 & ~n1495;
  assign n1497 = ~n1363 & ~n1370;
  assign n1498 = ~n1371 & ~n1497;
  assign n1499 = ~n687 & n1240;
  assign n1500 = n687 & n1242;
  assign n1501 = ~n656 & n1244;
  assign n1502 = n656 & n1246;
  assign n1503 = ~n1499 & ~n1500;
  assign n1504 = ~n1501 & ~n1502;
  assign n1505 = n1503 & n1504;
  assign n1506 = ~n61 & n682;
  assign n1507 = n72 & n525;
  assign n1508 = ~n1236 & ~n1507;
  assign n1509 = ~n680 & ~n1508;
  assign n1510 = n61 & n694;
  assign n1511 = ~n1506 & ~n1509;
  assign n1512 = ~n1510 & n1511;
  assign n1513 = n1505 & n1512;
  assign n1514 = ~n1425 & ~n1431;
  assign n1515 = ~n1432 & ~n1514;
  assign n1516 = ~n1505 & ~n1512;
  assign n1517 = n1515 & ~n1516;
  assign n1518 = ~n1513 & ~n1517;
  assign n1519 = n1498 & ~n1518;
  assign n1520 = ~n1498 & n1518;
  assign n1521 = n1400 & n1407;
  assign n1522 = ~n1400 & ~n1407;
  assign n1523 = ~n1521 & ~n1522;
  assign n1524 = ~n1520 & ~n1523;
  assign n1525 = ~n1519 & ~n1524;
  assign n1526 = n1496 & ~n1525;
  assign n1527 = ~n1496 & n1525;
  assign n1528 = ~n1526 & ~n1527;
  assign n1529 = n1477 & ~n1479;
  assign n1530 = ~n1480 & ~n1529;
  assign n1531 = n1528 & n1530;
  assign n1532 = ~n1526 & ~n1531;
  assign n1533 = n1487 & ~n1489;
  assign n1534 = ~n1490 & ~n1533;
  assign n1535 = ~n1532 & n1534;
  assign n1536 = ~n61 & ~n593;
  assign n1537 = n648 & ~n1536;
  assign n1538 = ~n687 & n1358;
  assign n1539 = ~n656 & n1357;
  assign n1540 = ~n687 & ~n1357;
  assign n1541 = n1018 & ~n1540;
  assign n1542 = ~n1538 & ~n1539;
  assign n1543 = ~n1541 & n1542;
  assign n1544 = n1537 & n1543;
  assign n1545 = ~n474 & n1140;
  assign n1546 = n474 & n1142;
  assign n1547 = ~n895 & n1144;
  assign n1548 = n895 & n1146;
  assign n1549 = ~n1545 & ~n1546;
  assign n1550 = ~n1547 & ~n1548;
  assign n1551 = n1549 & n1550;
  assign n1552 = n774 & n907;
  assign n1553 = n705 & ~n1023;
  assign n1554 = ~n774 & n910;
  assign n1555 = n912 & n1023;
  assign n1556 = ~n1552 & ~n1553;
  assign n1557 = ~n1554 & ~n1555;
  assign n1558 = n1556 & n1557;
  assign n1559 = n1551 & ~n1558;
  assign n1560 = ~n1551 & n1558;
  assign n1561 = ~n1559 & ~n1560;
  assign n1562 = n1544 & ~n1561;
  assign n1563 = n1551 & n1558;
  assign n1564 = ~n1562 & ~n1563;
  assign n1565 = ~n643 & n1358;
  assign n1566 = ~n687 & n1357;
  assign n1567 = ~n643 & ~n1357;
  assign n1568 = n1018 & ~n1567;
  assign n1569 = ~n1565 & ~n1566;
  assign n1570 = ~n1568 & n1569;
  assign n1571 = ~n656 & n1240;
  assign n1572 = n656 & n1242;
  assign n1573 = ~n532 & n1244;
  assign n1574 = n532 & n1246;
  assign n1575 = ~n1571 & ~n1572;
  assign n1576 = ~n1573 & ~n1574;
  assign n1577 = n1575 & n1576;
  assign n1578 = n1570 & ~n1577;
  assign n1579 = ~n1570 & n1577;
  assign n1580 = ~n1578 & ~n1579;
  assign n1581 = ~n57 & n631;
  assign n1582 = n57 & n638;
  assign n1583 = ~n72 & n645;
  assign n1584 = n72 & n649;
  assign n1585 = ~n1581 & ~n1582;
  assign n1586 = ~n1583 & ~n1584;
  assign n1587 = n1585 & n1586;
  assign n1588 = ~n1580 & n1587;
  assign n1589 = n1570 & n1577;
  assign n1590 = ~n1588 & ~n1589;
  assign n1591 = ~n1564 & ~n1590;
  assign n1592 = ~n1564 & n1590;
  assign n1593 = n1564 & ~n1590;
  assign n1594 = ~n1592 & ~n1593;
  assign n1595 = n1457 & n1464;
  assign n1596 = ~n1457 & ~n1464;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n1594 & ~n1597;
  assign n1599 = ~n1591 & ~n1598;
  assign n1600 = n1467 & ~n1469;
  assign n1601 = ~n1470 & ~n1600;
  assign n1602 = ~n1599 & n1601;
  assign n1603 = n1599 & ~n1601;
  assign n1604 = ~n1602 & ~n1603;
  assign n1605 = ~n1519 & ~n1520;
  assign n1606 = ~n1523 & n1605;
  assign n1607 = n1523 & ~n1605;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = n1604 & n1608;
  assign n1610 = ~n1602 & ~n1609;
  assign n1611 = ~n1528 & ~n1530;
  assign n1612 = ~n1531 & ~n1611;
  assign n1613 = ~n1610 & n1612;
  assign n1614 = n1610 & ~n1612;
  assign n1615 = ~n1613 & ~n1614;
  assign n1616 = ~n532 & n1240;
  assign n1617 = n532 & n1242;
  assign n1618 = ~n474 & n1244;
  assign n1619 = n474 & n1246;
  assign n1620 = ~n1616 & ~n1617;
  assign n1621 = ~n1618 & ~n1619;
  assign n1622 = n1620 & n1621;
  assign n1623 = n907 & n1023;
  assign n1624 = ~n57 & n705;
  assign n1625 = n910 & ~n1023;
  assign n1626 = n57 & n912;
  assign n1627 = ~n1623 & ~n1624;
  assign n1628 = ~n1625 & ~n1626;
  assign n1629 = n1627 & n1628;
  assign n1630 = n1622 & ~n1629;
  assign n1631 = ~n1622 & n1629;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = ~n895 & n1140;
  assign n1634 = n895 & n1142;
  assign n1635 = ~n774 & n1144;
  assign n1636 = n774 & n1146;
  assign n1637 = ~n1633 & ~n1634;
  assign n1638 = ~n1635 & ~n1636;
  assign n1639 = n1637 & n1638;
  assign n1640 = ~n1632 & n1639;
  assign n1641 = n1622 & n1629;
  assign n1642 = ~n1640 & ~n1641;
  assign n1643 = n1424 & ~n1642;
  assign n1644 = ~n1544 & n1561;
  assign n1645 = ~n1562 & ~n1644;
  assign n1646 = ~n1424 & n1642;
  assign n1647 = ~n1643 & ~n1646;
  assign n1648 = n1645 & n1647;
  assign n1649 = ~n1643 & ~n1648;
  assign n1650 = ~n1513 & ~n1516;
  assign n1651 = n1515 & ~n1650;
  assign n1652 = ~n1515 & n1650;
  assign n1653 = ~n1651 & ~n1652;
  assign n1654 = ~n1649 & ~n1653;
  assign n1655 = n1649 & n1653;
  assign n1656 = ~n1654 & ~n1655;
  assign n1657 = n1594 & n1597;
  assign n1658 = ~n1598 & ~n1657;
  assign n1659 = n1656 & n1658;
  assign n1660 = ~n1654 & ~n1659;
  assign n1661 = ~n1604 & ~n1608;
  assign n1662 = ~n1609 & ~n1661;
  assign n1663 = ~n1660 & n1662;
  assign n1664 = n1660 & ~n1662;
  assign n1665 = ~n656 & n1358;
  assign n1666 = ~n532 & n1357;
  assign n1667 = ~n656 & ~n1357;
  assign n1668 = n1018 & ~n1667;
  assign n1669 = ~n1665 & ~n1666;
  assign n1670 = ~n1668 & n1669;
  assign n1671 = ~n474 & n1240;
  assign n1672 = n474 & n1242;
  assign n1673 = ~n895 & n1244;
  assign n1674 = n895 & n1246;
  assign n1675 = ~n1671 & ~n1672;
  assign n1676 = ~n1673 & ~n1674;
  assign n1677 = n1675 & n1676;
  assign n1678 = n1670 & n1677;
  assign n1679 = n1670 & ~n1677;
  assign n1680 = ~n1670 & n1677;
  assign n1681 = ~n1679 & ~n1680;
  assign n1682 = ~n774 & n1140;
  assign n1683 = n774 & n1142;
  assign n1684 = ~n1023 & n1144;
  assign n1685 = n1023 & n1146;
  assign n1686 = ~n1682 & ~n1683;
  assign n1687 = ~n1684 & ~n1685;
  assign n1688 = n1686 & n1687;
  assign n1689 = ~n1681 & n1688;
  assign n1690 = ~n1678 & ~n1689;
  assign n1691 = ~n1537 & ~n1543;
  assign n1692 = ~n1544 & ~n1691;
  assign n1693 = ~n72 & n631;
  assign n1694 = n72 & n638;
  assign n1695 = ~n61 & n645;
  assign n1696 = n61 & n649;
  assign n1697 = ~n1693 & ~n1694;
  assign n1698 = ~n1695 & ~n1696;
  assign n1699 = n1697 & n1698;
  assign n1700 = ~n1692 & n1699;
  assign n1701 = n1692 & ~n1699;
  assign n1702 = ~n1700 & ~n1701;
  assign n1703 = ~n1690 & ~n1702;
  assign n1704 = n1692 & n1699;
  assign n1705 = ~n1703 & ~n1704;
  assign n1706 = n1580 & n1587;
  assign n1707 = ~n1580 & ~n1587;
  assign n1708 = ~n1706 & ~n1707;
  assign n1709 = ~n1705 & ~n1708;
  assign n1710 = ~n1645 & ~n1647;
  assign n1711 = ~n1648 & ~n1710;
  assign n1712 = n1705 & n1708;
  assign n1713 = ~n1709 & ~n1712;
  assign n1714 = n1711 & n1713;
  assign n1715 = ~n1709 & ~n1714;
  assign n1716 = ~n61 & ~n701;
  assign n1717 = n470 & ~n1716;
  assign n1718 = ~n532 & n1358;
  assign n1719 = ~n474 & n1357;
  assign n1720 = ~n532 & ~n1357;
  assign n1721 = n1018 & ~n1720;
  assign n1722 = ~n1718 & ~n1719;
  assign n1723 = ~n1721 & n1722;
  assign n1724 = n1717 & n1723;
  assign n1725 = n57 & n907;
  assign n1726 = ~n72 & n705;
  assign n1727 = ~n57 & n910;
  assign n1728 = n72 & n912;
  assign n1729 = ~n1725 & ~n1726;
  assign n1730 = ~n1727 & ~n1728;
  assign n1731 = n1729 & n1730;
  assign n1732 = n1724 & ~n1731;
  assign n1733 = ~n1724 & n1731;
  assign n1734 = ~n1732 & ~n1733;
  assign n1735 = n1536 & ~n1734;
  assign n1736 = n1724 & n1731;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = n1632 & ~n1639;
  assign n1739 = ~n1640 & ~n1738;
  assign n1740 = ~n1737 & n1739;
  assign n1741 = n1737 & ~n1739;
  assign n1742 = ~n1740 & ~n1741;
  assign n1743 = n1690 & n1702;
  assign n1744 = ~n1703 & ~n1743;
  assign n1745 = n1742 & n1744;
  assign n1746 = ~n1740 & ~n1745;
  assign n1747 = ~n895 & n1240;
  assign n1748 = n895 & n1242;
  assign n1749 = ~n774 & n1244;
  assign n1750 = n774 & n1246;
  assign n1751 = ~n1747 & ~n1748;
  assign n1752 = ~n1749 & ~n1750;
  assign n1753 = n1751 & n1752;
  assign n1754 = ~n1023 & n1140;
  assign n1755 = n1023 & n1142;
  assign n1756 = ~n57 & n1144;
  assign n1757 = n57 & n1146;
  assign n1758 = ~n1754 & ~n1755;
  assign n1759 = ~n1756 & ~n1757;
  assign n1760 = n1758 & n1759;
  assign n1761 = n1753 & ~n1760;
  assign n1762 = ~n1753 & n1760;
  assign n1763 = ~n1761 & ~n1762;
  assign n1764 = ~n72 & n910;
  assign n1765 = ~n61 & n705;
  assign n1766 = n61 & n912;
  assign n1767 = n72 & n907;
  assign n1768 = ~n1764 & ~n1765;
  assign n1769 = ~n1766 & ~n1767;
  assign n1770 = n1768 & n1769;
  assign n1771 = ~n1763 & n1770;
  assign n1772 = n1753 & n1760;
  assign n1773 = ~n1771 & ~n1772;
  assign n1774 = n1681 & ~n1688;
  assign n1775 = ~n1689 & ~n1774;
  assign n1776 = ~n1773 & n1775;
  assign n1777 = ~n1536 & n1734;
  assign n1778 = ~n1735 & ~n1777;
  assign n1779 = n1773 & ~n1775;
  assign n1780 = ~n1776 & ~n1779;
  assign n1781 = n1778 & n1780;
  assign n1782 = ~n1776 & ~n1781;
  assign n1783 = ~n1717 & ~n1723;
  assign n1784 = ~n1724 & ~n1783;
  assign n1785 = ~n774 & n1240;
  assign n1786 = n774 & n1242;
  assign n1787 = ~n1023 & n1244;
  assign n1788 = n1023 & n1246;
  assign n1789 = ~n1785 & ~n1786;
  assign n1790 = ~n1787 & ~n1788;
  assign n1791 = n1789 & n1790;
  assign n1792 = ~n474 & n1358;
  assign n1793 = ~n895 & n1357;
  assign n1794 = ~n474 & ~n1357;
  assign n1795 = n1018 & ~n1794;
  assign n1796 = ~n1792 & ~n1793;
  assign n1797 = ~n1795 & n1796;
  assign n1798 = ~n1791 & n1797;
  assign n1799 = n1791 & ~n1797;
  assign n1800 = ~n1798 & ~n1799;
  assign n1801 = ~n57 & n1140;
  assign n1802 = n57 & n1142;
  assign n1803 = ~n72 & n1144;
  assign n1804 = n72 & n1146;
  assign n1805 = ~n1801 & ~n1802;
  assign n1806 = ~n1803 & ~n1804;
  assign n1807 = n1805 & n1806;
  assign n1808 = ~n1800 & n1807;
  assign n1809 = n1791 & n1797;
  assign n1810 = ~n1808 & ~n1809;
  assign n1811 = n1784 & ~n1810;
  assign n1812 = n1763 & n1770;
  assign n1813 = ~n1763 & ~n1770;
  assign n1814 = ~n1812 & ~n1813;
  assign n1815 = ~n1784 & n1810;
  assign n1816 = ~n1811 & ~n1815;
  assign n1817 = ~n1814 & n1816;
  assign n1818 = ~n1811 & ~n1817;
  assign n1819 = ~n61 & ~n1082;
  assign n1820 = n888 & ~n1819;
  assign n1821 = ~n895 & n1358;
  assign n1822 = ~n774 & n1357;
  assign n1823 = ~n895 & ~n1357;
  assign n1824 = n1018 & ~n1823;
  assign n1825 = ~n1821 & ~n1822;
  assign n1826 = ~n1824 & n1825;
  assign n1827 = n1820 & n1826;
  assign n1828 = n1716 & n1827;
  assign n1829 = ~n1716 & n1827;
  assign n1830 = n1716 & ~n1827;
  assign n1831 = ~n1829 & ~n1830;
  assign n1832 = ~n1023 & n1240;
  assign n1833 = n1023 & n1242;
  assign n1834 = ~n57 & n1244;
  assign n1835 = n57 & n1246;
  assign n1836 = ~n1832 & ~n1833;
  assign n1837 = ~n1834 & ~n1835;
  assign n1838 = n1836 & n1837;
  assign n1839 = ~n72 & n1140;
  assign n1840 = n72 & n1142;
  assign n1841 = ~n61 & n1144;
  assign n1842 = n61 & n1146;
  assign n1843 = ~n1839 & ~n1840;
  assign n1844 = ~n1841 & ~n1842;
  assign n1845 = n1843 & n1844;
  assign n1846 = n1838 & n1845;
  assign n1847 = ~n1820 & ~n1826;
  assign n1848 = ~n1827 & ~n1847;
  assign n1849 = ~n1838 & ~n1845;
  assign n1850 = n1848 & ~n1849;
  assign n1851 = ~n1846 & ~n1850;
  assign n1852 = ~n1831 & ~n1851;
  assign n1853 = ~n1828 & ~n1852;
  assign n1854 = n1831 & n1851;
  assign n1855 = ~n1852 & ~n1854;
  assign n1856 = ~n1846 & ~n1849;
  assign n1857 = n1848 & ~n1856;
  assign n1858 = ~n1848 & n1856;
  assign n1859 = ~n1857 & ~n1858;
  assign n1860 = ~n61 & ~n1193;
  assign n1861 = n1191 & ~n1860;
  assign n1862 = n57 & ~n1018;
  assign n1863 = n1357 & ~n1862;
  assign n1864 = ~n1018 & n1023;
  assign n1865 = ~n1023 & ~n1358;
  assign n1866 = ~n1864 & ~n1865;
  assign n1867 = ~n1863 & ~n1866;
  assign n1868 = n1861 & n1867;
  assign n1869 = n1357 & ~n1864;
  assign n1870 = ~n774 & n1358;
  assign n1871 = n774 & n1018;
  assign n1872 = ~n1869 & ~n1871;
  assign n1873 = ~n1870 & n1872;
  assign n1874 = ~n57 & n1240;
  assign n1875 = n57 & n1242;
  assign n1876 = ~n72 & n1244;
  assign n1877 = n72 & n1246;
  assign n1878 = ~n1874 & ~n1875;
  assign n1879 = ~n1876 & ~n1877;
  assign n1880 = n1878 & n1879;
  assign n1881 = n1873 & ~n1880;
  assign n1882 = ~n1873 & n1880;
  assign n1883 = ~n1881 & ~n1882;
  assign n1884 = n1868 & ~n1883;
  assign n1885 = n1873 & n1880;
  assign n1886 = ~n1884 & ~n1885;
  assign n1887 = n1859 & n1886;
  assign n1888 = ~n1859 & ~n1886;
  assign n1889 = ~n72 & ~n1357;
  assign n1890 = n61 & ~n1018;
  assign n1891 = ~n1889 & n1890;
  assign n1892 = n72 & ~n1018;
  assign n1893 = n1357 & ~n1892;
  assign n1894 = ~n57 & n1018;
  assign n1895 = ~n1357 & ~n1862;
  assign n1896 = ~n1894 & n1895;
  assign n1897 = ~n1893 & ~n1896;
  assign n1898 = n1860 & n1897;
  assign n1899 = ~n1891 & ~n1898;
  assign n1900 = ~n1860 & ~n1897;
  assign n1901 = ~n1899 & ~n1900;
  assign n1902 = ~n1861 & ~n1867;
  assign n1903 = ~n1868 & ~n1902;
  assign n1904 = ~n72 & n1240;
  assign n1905 = n72 & n1242;
  assign n1906 = ~n61 & n1244;
  assign n1907 = n61 & n1246;
  assign n1908 = ~n1904 & ~n1905;
  assign n1909 = ~n1906 & ~n1907;
  assign n1910 = n1908 & n1909;
  assign n1911 = n1903 & n1910;
  assign n1912 = ~n1901 & ~n1911;
  assign n1913 = ~n1903 & ~n1910;
  assign n1914 = ~n1912 & ~n1913;
  assign n1915 = ~n1868 & n1883;
  assign n1916 = ~n1884 & ~n1915;
  assign n1917 = n1819 & n1916;
  assign n1918 = ~n1914 & ~n1917;
  assign n1919 = ~n1819 & ~n1916;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = ~n1888 & ~n1920;
  assign n1922 = ~n1887 & ~n1921;
  assign n1923 = n1855 & n1922;
  assign n1924 = ~n1855 & ~n1922;
  assign n1925 = n1800 & ~n1807;
  assign n1926 = ~n1808 & ~n1925;
  assign n1927 = ~n1924 & n1926;
  assign n1928 = ~n1923 & ~n1927;
  assign n1929 = ~n1853 & ~n1928;
  assign n1930 = n1853 & n1928;
  assign n1931 = n1814 & ~n1816;
  assign n1932 = ~n1817 & ~n1931;
  assign n1933 = ~n1930 & n1932;
  assign n1934 = ~n1929 & ~n1933;
  assign n1935 = ~n1818 & ~n1934;
  assign n1936 = n1818 & n1934;
  assign n1937 = ~n1778 & ~n1780;
  assign n1938 = ~n1781 & ~n1937;
  assign n1939 = ~n1936 & n1938;
  assign n1940 = ~n1935 & ~n1939;
  assign n1941 = ~n1782 & ~n1940;
  assign n1942 = n1782 & n1940;
  assign n1943 = ~n1742 & ~n1744;
  assign n1944 = ~n1745 & ~n1943;
  assign n1945 = ~n1942 & n1944;
  assign n1946 = ~n1941 & ~n1945;
  assign n1947 = ~n1746 & ~n1946;
  assign n1948 = n1746 & n1946;
  assign n1949 = ~n1711 & ~n1713;
  assign n1950 = ~n1714 & ~n1949;
  assign n1951 = ~n1948 & n1950;
  assign n1952 = ~n1947 & ~n1951;
  assign n1953 = ~n1715 & ~n1952;
  assign n1954 = n1715 & n1952;
  assign n1955 = ~n1656 & ~n1658;
  assign n1956 = ~n1659 & ~n1955;
  assign n1957 = ~n1954 & n1956;
  assign n1958 = ~n1953 & ~n1957;
  assign n1959 = ~n1664 & ~n1958;
  assign n1960 = ~n1663 & ~n1959;
  assign n1961 = n1615 & ~n1960;
  assign n1962 = ~n1613 & ~n1961;
  assign n1963 = n1532 & ~n1534;
  assign n1964 = ~n1535 & ~n1963;
  assign n1965 = ~n1962 & n1964;
  assign n1966 = ~n1535 & ~n1965;
  assign n1967 = n1491 & ~n1493;
  assign n1968 = ~n1494 & ~n1967;
  assign n1969 = ~n1966 & n1968;
  assign n1970 = ~n1494 & ~n1969;
  assign n1971 = n1311 & n1422;
  assign n1972 = ~n1423 & ~n1971;
  assign n1973 = ~n1970 & n1972;
  assign n1974 = ~n1423 & ~n1973;
  assign n1975 = n1303 & n1307;
  assign n1976 = ~n1308 & ~n1975;
  assign n1977 = ~n1974 & n1976;
  assign n1978 = ~n1308 & ~n1977;
  assign n1979 = ~n1122 & ~n1172;
  assign n1980 = ~n1173 & ~n1979;
  assign n1981 = ~n1978 & n1980;
  assign n1982 = ~n1173 & ~n1981;
  assign n1983 = n1117 & ~n1119;
  assign n1984 = ~n1120 & ~n1983;
  assign n1985 = ~n1982 & n1984;
  assign n1986 = ~n1120 & ~n1985;
  assign n1987 = n949 & n952;
  assign n1988 = ~n953 & ~n1987;
  assign n1989 = ~n1986 & n1988;
  assign n1990 = ~n953 & ~n1989;
  assign n1991 = n748 & ~n769;
  assign n1992 = ~n770 & ~n1991;
  assign n1993 = ~n1990 & n1992;
  assign n1994 = ~n770 & ~n1993;
  assign n1995 = ~n758 & ~n767;
  assign n1996 = ~n761 & ~n764;
  assign n1997 = ~n636 & n680;
  assign n1998 = ~n693 & ~n1997;
  assign n1999 = ~n636 & n682;
  assign n2000 = ~n1998 & ~n1999;
  assign n2001 = ~n737 & n2000;
  assign n2002 = n737 & ~n2000;
  assign n2003 = ~n2001 & ~n2002;
  assign n2004 = ~n1996 & n2003;
  assign n2005 = n1996 & ~n2003;
  assign n2006 = ~n2004 & ~n2005;
  assign n2007 = ~n1995 & n2006;
  assign n2008 = n1995 & ~n2006;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = ~n1994 & n2009;
  assign n2011 = n1994 & ~n2009;
  assign n2012 = ~n2010 & ~n2011;
  assign n2013 = ~n129 & ~n193;
  assign n2014 = ~n358 & n2013;
  assign n2015 = n560 & n2014;
  assign n2016 = ~n252 & ~n546;
  assign n2017 = n841 & n2016;
  assign n2018 = n235 & ~n355;
  assign n2019 = n406 & n2018;
  assign n2020 = n160 & n867;
  assign n2021 = n986 & n2017;
  assign n2022 = n2020 & n2021;
  assign n2023 = n2015 & n2019;
  assign n2024 = n2022 & n2023;
  assign n2025 = ~n241 & ~n320;
  assign n2026 = ~n332 & ~n347;
  assign n2027 = ~n391 & ~n434;
  assign n2028 = n2026 & n2027;
  assign n2029 = n2025 & n2028;
  assign n2030 = n295 & n2029;
  assign n2031 = ~n268 & ~n346;
  assign n2032 = ~n356 & ~n377;
  assign n2033 = ~n563 & n2032;
  assign n2034 = n2031 & n2033;
  assign n2035 = ~n133 & ~n162;
  assign n2036 = ~n167 & ~n240;
  assign n2037 = ~n319 & ~n328;
  assign n2038 = ~n818 & n2037;
  assign n2039 = n2035 & n2036;
  assign n2040 = n238 & n2039;
  assign n2041 = n2038 & n2040;
  assign n2042 = n2034 & n2041;
  assign n2043 = ~n199 & ~n299;
  assign n2044 = ~n594 & n2043;
  assign n2045 = ~n138 & ~n245;
  assign n2046 = ~n284 & ~n404;
  assign n2047 = n2045 & n2046;
  assign n2048 = n256 & n341;
  assign n2049 = n351 & n481;
  assign n2050 = n2048 & n2049;
  assign n2051 = n2044 & n2047;
  assign n2052 = n2050 & n2051;
  assign n2053 = n225 & n2052;
  assign n2054 = n2030 & n2053;
  assign n2055 = n2024 & n2042;
  assign n2056 = n2054 & n2055;
  assign n2057 = ~n2012 & ~n2056;
  assign n2058 = n1990 & ~n1992;
  assign n2059 = ~n1993 & ~n2058;
  assign n2060 = ~n129 & ~n220;
  assign n2061 = ~n228 & ~n320;
  assign n2062 = ~n377 & n2061;
  assign n2063 = n359 & n2060;
  assign n2064 = n439 & n552;
  assign n2065 = n2063 & n2064;
  assign n2066 = n171 & n2062;
  assign n2067 = n306 & n799;
  assign n2068 = n2066 & n2067;
  assign n2069 = n2065 & n2068;
  assign n2070 = n574 & n855;
  assign n2071 = n2069 & n2070;
  assign n2072 = n996 & n2071;
  assign n2073 = ~n2059 & ~n2072;
  assign n2074 = n1986 & ~n1988;
  assign n2075 = ~n1989 & ~n2074;
  assign n2076 = ~n267 & ~n475;
  assign n2077 = ~n172 & ~n392;
  assign n2078 = ~n284 & ~n356;
  assign n2079 = ~n497 & n2078;
  assign n2080 = ~n133 & ~n342;
  assign n2081 = n318 & n2080;
  assign n2082 = n552 & n2076;
  assign n2083 = n2077 & n2082;
  assign n2084 = n2017 & n2081;
  assign n2085 = n2044 & n2079;
  assign n2086 = n2084 & n2085;
  assign n2087 = n453 & n2083;
  assign n2088 = n2086 & n2087;
  assign n2089 = ~n360 & ~n405;
  assign n2090 = ~n168 & ~n362;
  assign n2091 = ~n144 & ~n216;
  assign n2092 = ~n241 & ~n268;
  assign n2093 = ~n304 & n2092;
  assign n2094 = n792 & n2091;
  assign n2095 = n2093 & n2094;
  assign n2096 = ~n162 & ~n296;
  assign n2097 = n2090 & n2096;
  assign n2098 = n562 & n2097;
  assign n2099 = n433 & n2098;
  assign n2100 = n2095 & n2099;
  assign n2101 = ~n177 & ~n214;
  assign n2102 = ~n300 & n2101;
  assign n2103 = ~n217 & ~n229;
  assign n2104 = ~n273 & n2103;
  assign n2105 = ~n339 & n436;
  assign n2106 = n549 & n597;
  assign n2107 = n2089 & n2106;
  assign n2108 = n2102 & n2105;
  assign n2109 = n2104 & n2108;
  assign n2110 = n428 & n2107;
  assign n2111 = n2109 & n2110;
  assign n2112 = n2088 & n2111;
  assign n2113 = n2100 & n2112;
  assign n2114 = ~n2075 & ~n2113;
  assign n2115 = n1982 & ~n1984;
  assign n2116 = ~n1985 & ~n2115;
  assign n2117 = ~n201 & ~n404;
  assign n2118 = ~n565 & ~n657;
  assign n2119 = n2117 & n2118;
  assign n2120 = n344 & n2119;
  assign n2121 = n483 & n613;
  assign n2122 = n2102 & n2121;
  assign n2123 = n2120 & n2122;
  assign n2124 = ~n255 & ~n350;
  assign n2125 = ~n378 & n2124;
  assign n2126 = n2088 & n2125;
  assign n2127 = ~n216 & ~n228;
  assign n2128 = ~n230 & n2127;
  assign n2129 = ~n167 & ~n423;
  assign n2130 = ~n217 & ~n303;
  assign n2131 = n2129 & n2130;
  assign n2132 = n823 & n861;
  assign n2133 = n2131 & n2132;
  assign n2134 = n1324 & n2128;
  assign n2135 = n2133 & n2134;
  assign n2136 = n2030 & n2135;
  assign n2137 = n2123 & n2136;
  assign n2138 = n2126 & n2137;
  assign n2139 = ~n2116 & ~n2138;
  assign n2140 = n1978 & ~n1980;
  assign n2141 = ~n1981 & ~n2140;
  assign n2142 = ~n200 & ~n285;
  assign n2143 = ~n179 & ~n216;
  assign n2144 = ~n292 & ~n320;
  assign n2145 = n435 & n2144;
  assign n2146 = n549 & n977;
  assign n2147 = n2142 & n2143;
  assign n2148 = n2146 & n2147;
  assign n2149 = n2145 & n2148;
  assign n2150 = n829 & n2149;
  assign n2151 = ~n158 & ~n245;
  assign n2152 = ~n253 & ~n315;
  assign n2153 = ~n429 & n2152;
  assign n2154 = n2151 & n2153;
  assign n2155 = ~n142 & ~n346;
  assign n2156 = n817 & n2155;
  assign n2157 = ~n220 & ~n246;
  assign n2158 = n1340 & n2157;
  assign n2159 = n848 & n2090;
  assign n2160 = n2158 & n2159;
  assign n2161 = ~n199 & ~n227;
  assign n2162 = ~n229 & ~n234;
  assign n2163 = ~n284 & ~n353;
  assign n2164 = n2162 & n2163;
  assign n2165 = n612 & n2161;
  assign n2166 = n2164 & n2165;
  assign n2167 = n2154 & n2166;
  assign n2168 = n2160 & n2167;
  assign n2169 = n2150 & n2168;
  assign n2170 = n2156 & n2169;
  assign n2171 = ~n2141 & ~n2170;
  assign n2172 = n1974 & ~n1976;
  assign n2173 = ~n1977 & ~n2172;
  assign n2174 = ~n346 & ~n429;
  assign n2175 = n668 & n2174;
  assign n2176 = n782 & n808;
  assign n2177 = n2175 & n2176;
  assign n2178 = n257 & n2177;
  assign n2179 = ~n246 & ~n315;
  assign n2180 = ~n162 & ~n195;
  assign n2181 = ~n548 & n2180;
  assign n2182 = n667 & n2181;
  assign n2183 = ~n142 & ~n144;
  assign n2184 = ~n244 & n2183;
  assign n2185 = ~n158 & ~n175;
  assign n2186 = ~n337 & ~n350;
  assign n2187 = n2185 & n2186;
  assign n2188 = n354 & n476;
  assign n2189 = n564 & n979;
  assign n2190 = n2179 & n2189;
  assign n2191 = n2187 & n2188;
  assign n2192 = n2184 & n2191;
  assign n2193 = n781 & n2190;
  assign n2194 = n2182 & n2193;
  assign n2195 = n2178 & n2192;
  assign n2196 = n2194 & n2195;
  assign n2197 = n875 & n2196;
  assign n2198 = ~n2173 & ~n2197;
  assign n2199 = n1970 & ~n1972;
  assign n2200 = ~n1973 & ~n2199;
  assign n2201 = ~n228 & ~n353;
  assign n2202 = ~n405 & ~n456;
  assign n2203 = ~n497 & n2202;
  assign n2204 = ~n156 & ~n180;
  assign n2205 = ~n239 & ~n480;
  assign n2206 = n2204 & n2205;
  assign n2207 = n357 & n2201;
  assign n2208 = n2206 & n2207;
  assign n2209 = n2203 & n2208;
  assign n2210 = n796 & n2209;
  assign n2211 = n145 & n213;
  assign n2212 = ~n286 & ~n404;
  assign n2213 = n2142 & n2212;
  assign n2214 = ~n289 & ~n297;
  assign n2215 = ~n315 & ~n396;
  assign n2216 = n2214 & n2215;
  assign n2217 = n567 & n2216;
  assign n2218 = n2213 & n2217;
  assign n2219 = n453 & n1043;
  assign n2220 = n2218 & n2219;
  assign n2221 = ~n243 & n436;
  assign n2222 = n2220 & n2221;
  assign n2223 = ~n172 & ~n296;
  assign n2224 = ~n391 & ~n616;
  assign n2225 = n2223 & n2224;
  assign n2226 = n435 & n801;
  assign n2227 = n2225 & n2226;
  assign n2228 = ~n215 & ~n2211;
  assign n2229 = ~n167 & n2228;
  assign n2230 = ~n237 & ~n292;
  assign n2231 = ~n475 & n2230;
  assign n2232 = n235 & n2229;
  assign n2233 = n2231 & n2232;
  assign n2234 = n2227 & n2233;
  assign n2235 = n2210 & n2234;
  assign n2236 = n2222 & n2235;
  assign n2237 = ~n2200 & ~n2236;
  assign n2238 = n1966 & ~n1968;
  assign n2239 = ~n1969 & ~n2238;
  assign n2240 = ~n245 & ~n328;
  assign n2241 = ~n234 & ~n404;
  assign n2242 = n498 & n2241;
  assign n2243 = n596 & n978;
  assign n2244 = n2242 & n2243;
  assign n2245 = ~n289 & ~n346;
  assign n2246 = ~n424 & ~n430;
  assign n2247 = n2245 & n2246;
  assign n2248 = n792 & n2247;
  assign n2249 = n412 & n504;
  assign n2250 = n2104 & n2249;
  assign n2251 = n2248 & n2250;
  assign n2252 = ~n199 & ~n317;
  assign n2253 = ~n339 & ~n378;
  assign n2254 = ~n392 & ~n405;
  assign n2255 = ~n563 & n2254;
  assign n2256 = n2252 & n2253;
  assign n2257 = n316 & n454;
  assign n2258 = n2240 & n2257;
  assign n2259 = n2255 & n2256;
  assign n2260 = n867 & n2259;
  assign n2261 = n2244 & n2258;
  assign n2262 = n2260 & n2261;
  assign n2263 = n192 & n2262;
  assign n2264 = n2251 & n2263;
  assign n2265 = ~n2239 & ~n2264;
  assign n2266 = n1962 & ~n1964;
  assign n2267 = ~n1965 & ~n2266;
  assign n2268 = ~n138 & ~n174;
  assign n2269 = ~n201 & ~n237;
  assign n2270 = ~n378 & ~n456;
  assign n2271 = ~n391 & ~n565;
  assign n2272 = ~n304 & ~n327;
  assign n2273 = ~n657 & n2272;
  assign n2274 = n2271 & n2273;
  assign n2275 = ~n289 & ~n377;
  assign n2276 = n567 & n2275;
  assign n2277 = n843 & n2269;
  assign n2278 = n2270 & n2277;
  assign n2279 = n777 & n2276;
  assign n2280 = n2128 & n2279;
  assign n2281 = n2182 & n2278;
  assign n2282 = n2274 & n2281;
  assign n2283 = n2280 & n2282;
  assign n2284 = ~n144 & ~n232;
  assign n2285 = ~n271 & ~n284;
  assign n2286 = ~n424 & n2285;
  assign n2287 = n333 & n2284;
  assign n2288 = n482 & n823;
  assign n2289 = n2268 & n2288;
  assign n2290 = n2286 & n2287;
  assign n2291 = n2289 & n2290;
  assign n2292 = n864 & n2244;
  assign n2293 = n2291 & n2292;
  assign n2294 = n804 & n2293;
  assign n2295 = n446 & n2294;
  assign n2296 = n2283 & n2295;
  assign n2297 = ~n2267 & ~n2296;
  assign n2298 = ~n1615 & n1960;
  assign n2299 = ~n1961 & ~n2298;
  assign n2300 = ~n299 & ~n478;
  assign n2301 = ~n292 & ~n349;
  assign n2302 = ~n405 & n2301;
  assign n2303 = n1005 & n2302;
  assign n2304 = ~n233 & ~n286;
  assign n2305 = ~n303 & ~n492;
  assign n2306 = ~n546 & n2305;
  assign n2307 = n2304 & n2306;
  assign n2308 = n137 & n140;
  assign n2309 = ~n201 & ~n2308;
  assign n2310 = ~n320 & ~n455;
  assign n2311 = n2309 & n2310;
  assign n2312 = n2303 & n2311;
  assign n2313 = n2307 & n2312;
  assign n2314 = ~n168 & ~n179;
  assign n2315 = ~n229 & ~n347;
  assign n2316 = ~n450 & ~n616;
  assign n2317 = n2315 & n2316;
  assign n2318 = n359 & n2314;
  assign n2319 = n538 & n2270;
  assign n2320 = n2300 & n2319;
  assign n2321 = n2317 & n2318;
  assign n2322 = n331 & n2321;
  assign n2323 = n2320 & n2322;
  assign n2324 = n2178 & n2323;
  assign n2325 = n2313 & n2324;
  assign n2326 = ~n2299 & ~n2325;
  assign n2327 = ~n1663 & ~n1664;
  assign n2328 = ~n1958 & n2327;
  assign n2329 = n1958 & ~n2327;
  assign n2330 = ~n2328 & ~n2329;
  assign n2331 = ~n296 & ~n377;
  assign n2332 = ~n450 & ~n565;
  assign n2333 = ~n818 & n2332;
  assign n2334 = n567 & n2331;
  assign n2335 = n2333 & n2334;
  assign n2336 = n171 & n270;
  assign n2337 = n984 & n2336;
  assign n2338 = n807 & n2335;
  assign n2339 = n2337 & n2338;
  assign n2340 = n2024 & n2339;
  assign n2341 = n2251 & n2340;
  assign n2342 = n2330 & n2341;
  assign n2343 = n2299 & n2325;
  assign n2344 = ~n2326 & ~n2343;
  assign n2345 = ~n2342 & n2344;
  assign n2346 = ~n2326 & ~n2345;
  assign n2347 = n2267 & n2296;
  assign n2348 = ~n2297 & ~n2347;
  assign n2349 = ~n2346 & n2348;
  assign n2350 = ~n2297 & ~n2349;
  assign n2351 = n2239 & n2264;
  assign n2352 = ~n2265 & ~n2351;
  assign n2353 = ~n2350 & n2352;
  assign n2354 = ~n2265 & ~n2353;
  assign n2355 = n2200 & n2236;
  assign n2356 = ~n2237 & ~n2355;
  assign n2357 = ~n2354 & n2356;
  assign n2358 = ~n2237 & ~n2357;
  assign n2359 = n2173 & n2197;
  assign n2360 = ~n2198 & ~n2359;
  assign n2361 = ~n2358 & n2360;
  assign n2362 = ~n2198 & ~n2361;
  assign n2363 = n2141 & n2170;
  assign n2364 = ~n2171 & ~n2363;
  assign n2365 = ~n2362 & n2364;
  assign n2366 = ~n2171 & ~n2365;
  assign n2367 = n2116 & n2138;
  assign n2368 = ~n2139 & ~n2367;
  assign n2369 = ~n2366 & n2368;
  assign n2370 = ~n2139 & ~n2369;
  assign n2371 = n2075 & n2113;
  assign n2372 = ~n2114 & ~n2371;
  assign n2373 = ~n2370 & n2372;
  assign n2374 = ~n2114 & ~n2373;
  assign n2375 = n2059 & n2072;
  assign n2376 = ~n2073 & ~n2375;
  assign n2377 = ~n2374 & n2376;
  assign n2378 = ~n2073 & ~n2377;
  assign n2379 = n2012 & n2056;
  assign n2380 = ~n2057 & ~n2379;
  assign n2381 = ~n2378 & n2380;
  assign n2382 = ~n2057 & ~n2381;
  assign n2383 = ~n239 & ~n339;
  assign n2384 = ~n657 & n2383;
  assign n2385 = n860 & n2384;
  assign n2386 = ~n195 & ~n348;
  assign n2387 = ~n220 & ~n346;
  assign n2388 = ~n480 & n2387;
  assign n2389 = n2079 & n2388;
  assign n2390 = ~n232 & ~n317;
  assign n2391 = n564 & n609;
  assign n2392 = n823 & n2300;
  assign n2393 = n2386 & n2390;
  assign n2394 = n2392 & n2393;
  assign n2395 = n2391 & n2394;
  assign n2396 = n2385 & n2389;
  assign n2397 = n2395 & n2396;
  assign n2398 = n804 & n1004;
  assign n2399 = n2397 & n2398;
  assign n2400 = n2222 & n2399;
  assign n2401 = n636 & n643;
  assign n2402 = ~n636 & ~n643;
  assign n2403 = ~n2401 & ~n2402;
  assign n2404 = ~n692 & ~n2403;
  assign n2405 = n692 & n2403;
  assign n2406 = ~n2404 & ~n2405;
  assign n2407 = ~n525 & ~n2406;
  assign n2408 = ~n2007 & ~n2010;
  assign n2409 = ~n2001 & ~n2004;
  assign n2410 = n2408 & ~n2409;
  assign n2411 = ~n2408 & n2409;
  assign n2412 = ~n2410 & ~n2411;
  assign n2413 = n2407 & n2412;
  assign n2414 = ~n2407 & ~n2412;
  assign n2415 = ~n2413 & ~n2414;
  assign n2416 = ~n2400 & ~n2415;
  assign n2417 = n2400 & n2415;
  assign n2418 = ~n2416 & ~n2417;
  assign n2419 = ~n2382 & n2418;
  assign n2420 = n2382 & ~n2418;
  assign n2421 = ~n2419 & ~n2420;
  assign n2422 = n76 & n2421;
  assign n2423 = n57 & n72;
  assign n2424 = ~n57 & ~n72;
  assign n2425 = ~n2423 & ~n2424;
  assign n2426 = n68 & n2425;
  assign n2427 = n2378 & ~n2380;
  assign n2428 = ~n2381 & ~n2427;
  assign n2429 = n2421 & n2428;
  assign n2430 = n2374 & ~n2376;
  assign n2431 = ~n2377 & ~n2430;
  assign n2432 = n2428 & n2431;
  assign n2433 = n2370 & ~n2372;
  assign n2434 = ~n2373 & ~n2433;
  assign n2435 = n2431 & n2434;
  assign n2436 = n2366 & ~n2368;
  assign n2437 = ~n2369 & ~n2436;
  assign n2438 = n2434 & n2437;
  assign n2439 = n2362 & ~n2364;
  assign n2440 = ~n2365 & ~n2439;
  assign n2441 = n2437 & n2440;
  assign n2442 = n2358 & ~n2360;
  assign n2443 = ~n2361 & ~n2442;
  assign n2444 = n2440 & n2443;
  assign n2445 = n2354 & ~n2356;
  assign n2446 = ~n2357 & ~n2445;
  assign n2447 = n2443 & n2446;
  assign n2448 = n2350 & ~n2352;
  assign n2449 = ~n2353 & ~n2448;
  assign n2450 = n2446 & n2449;
  assign n2451 = n2346 & ~n2348;
  assign n2452 = ~n2349 & ~n2451;
  assign n2453 = n2449 & n2452;
  assign n2454 = ~n2449 & ~n2452;
  assign n2455 = ~n2453 & ~n2454;
  assign n2456 = ~n2330 & ~n2341;
  assign n2457 = ~n2342 & ~n2456;
  assign n2458 = ~n2452 & n2457;
  assign n2459 = n2342 & ~n2344;
  assign n2460 = ~n2345 & ~n2459;
  assign n2461 = ~n2458 & n2460;
  assign n2462 = n2455 & n2461;
  assign n2463 = ~n2453 & ~n2462;
  assign n2464 = ~n2446 & ~n2449;
  assign n2465 = ~n2450 & ~n2464;
  assign n2466 = ~n2463 & n2465;
  assign n2467 = ~n2450 & ~n2466;
  assign n2468 = ~n2443 & ~n2446;
  assign n2469 = ~n2447 & ~n2468;
  assign n2470 = ~n2467 & n2469;
  assign n2471 = ~n2447 & ~n2470;
  assign n2472 = ~n2440 & ~n2443;
  assign n2473 = ~n2444 & ~n2472;
  assign n2474 = ~n2471 & n2473;
  assign n2475 = ~n2444 & ~n2474;
  assign n2476 = ~n2437 & ~n2440;
  assign n2477 = ~n2441 & ~n2476;
  assign n2478 = ~n2475 & n2477;
  assign n2479 = ~n2441 & ~n2478;
  assign n2480 = ~n2434 & ~n2437;
  assign n2481 = ~n2438 & ~n2480;
  assign n2482 = ~n2479 & n2481;
  assign n2483 = ~n2438 & ~n2482;
  assign n2484 = ~n2431 & ~n2434;
  assign n2485 = ~n2435 & ~n2484;
  assign n2486 = ~n2483 & n2485;
  assign n2487 = ~n2435 & ~n2486;
  assign n2488 = ~n2428 & ~n2431;
  assign n2489 = ~n2432 & ~n2488;
  assign n2490 = ~n2487 & n2489;
  assign n2491 = ~n2432 & ~n2490;
  assign n2492 = ~n2421 & ~n2428;
  assign n2493 = ~n2429 & ~n2492;
  assign n2494 = ~n2491 & n2493;
  assign n2495 = ~n2429 & ~n2494;
  assign n2496 = ~n2416 & ~n2419;
  assign n2497 = ~n200 & ~n227;
  assign n2498 = ~n239 & ~n362;
  assign n2499 = ~n396 & n2498;
  assign n2500 = n2497 & n2499;
  assign n2501 = n302 & n2500;
  assign n2502 = ~n230 & ~n289;
  assign n2503 = ~n332 & ~n405;
  assign n2504 = n2502 & n2503;
  assign n2505 = n316 & n597;
  assign n2506 = n819 & n2505;
  assign n2507 = n986 & n2504;
  assign n2508 = n2506 & n2507;
  assign n2509 = n543 & n2508;
  assign n2510 = n2178 & n2501;
  assign n2511 = n2509 & n2510;
  assign n2512 = n1333 & n2511;
  assign n2513 = n2496 & n2512;
  assign n2514 = ~n2496 & ~n2512;
  assign n2515 = ~n2513 & ~n2514;
  assign n2516 = n2421 & ~n2515;
  assign n2517 = ~n2421 & n2515;
  assign n2518 = ~n2516 & ~n2517;
  assign n2519 = ~n2495 & n2518;
  assign n2520 = n2495 & ~n2518;
  assign n2521 = ~n2519 & ~n2520;
  assign n2522 = n2426 & n2521;
  assign n2523 = ~n68 & ~n75;
  assign n2524 = n2425 & n2523;
  assign n2525 = n2428 & n2524;
  assign n2526 = n68 & ~n2425;
  assign n2527 = ~n2515 & n2526;
  assign n2528 = ~n2422 & ~n2525;
  assign n2529 = ~n2527 & n2528;
  assign n2530 = ~n2522 & n2529;
  assign n2531 = ~n57 & ~n2530;
  assign n2532 = n57 & n2530;
  assign n2533 = ~n2531 & ~n2532;
  assign n2534 = n474 & n532;
  assign n2535 = ~n474 & ~n532;
  assign n2536 = ~n2534 & ~n2535;
  assign n2537 = n474 & n895;
  assign n2538 = ~n474 & ~n895;
  assign n2539 = ~n2537 & ~n2538;
  assign n2540 = n532 & n656;
  assign n2541 = ~n532 & ~n656;
  assign n2542 = ~n2540 & ~n2541;
  assign n2543 = ~n2536 & ~n2539;
  assign n2544 = n2542 & n2543;
  assign n2545 = n2452 & n2544;
  assign n2546 = n2539 & n2542;
  assign n2547 = n2463 & ~n2465;
  assign n2548 = ~n2466 & ~n2547;
  assign n2549 = n2546 & n2548;
  assign n2550 = n2536 & ~n2539;
  assign n2551 = n2449 & n2550;
  assign n2552 = n2539 & ~n2542;
  assign n2553 = n2446 & n2552;
  assign n2554 = ~n2545 & ~n2551;
  assign n2555 = ~n2553 & n2554;
  assign n2556 = ~n2549 & n2555;
  assign n2557 = n656 & n2556;
  assign n2558 = ~n656 & ~n2556;
  assign n2559 = ~n2557 & ~n2558;
  assign n2560 = n656 & n687;
  assign n2561 = ~n656 & ~n687;
  assign n2562 = ~n2560 & ~n2561;
  assign n2563 = n643 & n687;
  assign n2564 = ~n643 & ~n687;
  assign n2565 = ~n2563 & ~n2564;
  assign n2566 = ~n2562 & n2565;
  assign n2567 = ~n2457 & n2566;
  assign n2568 = ~n2403 & n2562;
  assign n2569 = n2460 & n2568;
  assign n2570 = ~n2457 & ~n2460;
  assign n2571 = ~n2344 & n2457;
  assign n2572 = ~n2570 & ~n2571;
  assign n2573 = n2403 & n2562;
  assign n2574 = ~n2572 & n2573;
  assign n2575 = ~n2567 & ~n2569;
  assign n2576 = ~n2574 & n2575;
  assign n2577 = ~n636 & ~n2457;
  assign n2578 = n2562 & n2577;
  assign n2579 = ~n2576 & n2578;
  assign n2580 = n2576 & ~n2578;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = n2559 & n2581;
  assign n2583 = ~n2457 & n2562;
  assign n2584 = ~n2457 & n2539;
  assign n2585 = ~n2457 & n2550;
  assign n2586 = n2460 & n2552;
  assign n2587 = n2546 & ~n2572;
  assign n2588 = ~n2585 & ~n2586;
  assign n2589 = ~n2587 & n2588;
  assign n2590 = ~n656 & ~n2584;
  assign n2591 = n2589 & n2590;
  assign n2592 = ~n2457 & n2544;
  assign n2593 = n2452 & ~n2571;
  assign n2594 = ~n2452 & n2571;
  assign n2595 = ~n2593 & ~n2594;
  assign n2596 = n2546 & ~n2595;
  assign n2597 = n2460 & n2550;
  assign n2598 = n2452 & n2552;
  assign n2599 = ~n2592 & ~n2597;
  assign n2600 = ~n2598 & n2599;
  assign n2601 = ~n2596 & n2600;
  assign n2602 = n2591 & n2601;
  assign n2603 = n2583 & n2602;
  assign n2604 = ~n2583 & n2602;
  assign n2605 = n2583 & ~n2602;
  assign n2606 = ~n2604 & ~n2605;
  assign n2607 = n2452 & n2550;
  assign n2608 = ~n2455 & ~n2461;
  assign n2609 = ~n2462 & ~n2608;
  assign n2610 = n2546 & n2609;
  assign n2611 = n2460 & n2544;
  assign n2612 = n2449 & n2552;
  assign n2613 = ~n2607 & ~n2611;
  assign n2614 = ~n2612 & n2613;
  assign n2615 = ~n2610 & n2614;
  assign n2616 = ~n656 & ~n2615;
  assign n2617 = n656 & n2615;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = ~n2606 & n2618;
  assign n2620 = ~n2603 & ~n2619;
  assign n2621 = ~n2559 & ~n2581;
  assign n2622 = ~n2582 & ~n2621;
  assign n2623 = ~n2620 & n2622;
  assign n2624 = ~n2582 & ~n2623;
  assign n2625 = n2449 & n2544;
  assign n2626 = n2467 & ~n2469;
  assign n2627 = ~n2470 & ~n2626;
  assign n2628 = n2546 & n2627;
  assign n2629 = n2446 & n2550;
  assign n2630 = n2443 & n2552;
  assign n2631 = ~n2625 & ~n2629;
  assign n2632 = ~n2630 & n2631;
  assign n2633 = ~n2628 & n2632;
  assign n2634 = ~n656 & ~n2633;
  assign n2635 = n656 & n2633;
  assign n2636 = ~n2634 & ~n2635;
  assign n2637 = ~n2562 & ~n2565;
  assign n2638 = n2403 & n2637;
  assign n2639 = ~n2457 & n2638;
  assign n2640 = n2573 & ~n2595;
  assign n2641 = n2460 & n2566;
  assign n2642 = n2452 & n2568;
  assign n2643 = ~n2639 & ~n2641;
  assign n2644 = ~n2642 & n2643;
  assign n2645 = ~n2640 & n2644;
  assign n2646 = n2576 & ~n2583;
  assign n2647 = ~n636 & ~n2646;
  assign n2648 = ~n2645 & n2647;
  assign n2649 = n2645 & ~n2647;
  assign n2650 = ~n2648 & ~n2649;
  assign n2651 = n2636 & n2650;
  assign n2652 = ~n2636 & ~n2650;
  assign n2653 = ~n2651 & ~n2652;
  assign n2654 = n2624 & ~n2653;
  assign n2655 = ~n2624 & n2653;
  assign n2656 = ~n2654 & ~n2655;
  assign n2657 = n774 & n1023;
  assign n2658 = ~n774 & ~n1023;
  assign n2659 = ~n2657 & ~n2658;
  assign n2660 = n57 & n1023;
  assign n2661 = ~n57 & ~n1023;
  assign n2662 = ~n2660 & ~n2661;
  assign n2663 = n2659 & ~n2662;
  assign n2664 = n2437 & n2663;
  assign n2665 = n774 & n895;
  assign n2666 = ~n774 & ~n895;
  assign n2667 = ~n2665 & ~n2666;
  assign n2668 = n2662 & n2667;
  assign n2669 = n2479 & ~n2481;
  assign n2670 = ~n2482 & ~n2669;
  assign n2671 = n2668 & n2670;
  assign n2672 = ~n2659 & ~n2662;
  assign n2673 = n2667 & n2672;
  assign n2674 = n2440 & n2673;
  assign n2675 = n2662 & ~n2667;
  assign n2676 = n2434 & n2675;
  assign n2677 = ~n2664 & ~n2674;
  assign n2678 = ~n2676 & n2677;
  assign n2679 = ~n2671 & n2678;
  assign n2680 = n895 & n2679;
  assign n2681 = ~n895 & ~n2679;
  assign n2682 = ~n2680 & ~n2681;
  assign n2683 = n2656 & n2682;
  assign n2684 = ~n2656 & ~n2682;
  assign n2685 = ~n2683 & ~n2684;
  assign n2686 = n2443 & n2673;
  assign n2687 = n2475 & ~n2477;
  assign n2688 = ~n2478 & ~n2687;
  assign n2689 = n2668 & n2688;
  assign n2690 = n2440 & n2663;
  assign n2691 = n2437 & n2675;
  assign n2692 = ~n2686 & ~n2690;
  assign n2693 = ~n2691 & n2692;
  assign n2694 = ~n2689 & n2693;
  assign n2695 = n895 & ~n2694;
  assign n2696 = ~n895 & n2694;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = n2620 & ~n2622;
  assign n2699 = ~n2623 & ~n2698;
  assign n2700 = n2697 & ~n2699;
  assign n2701 = ~n2697 & n2699;
  assign n2702 = ~n2606 & ~n2618;
  assign n2703 = n2606 & n2618;
  assign n2704 = ~n2702 & ~n2703;
  assign n2705 = n2446 & n2673;
  assign n2706 = n2471 & ~n2473;
  assign n2707 = ~n2474 & ~n2706;
  assign n2708 = n2668 & n2707;
  assign n2709 = n2443 & n2663;
  assign n2710 = n2440 & n2675;
  assign n2711 = ~n2705 & ~n2709;
  assign n2712 = ~n2710 & n2711;
  assign n2713 = ~n2708 & n2712;
  assign n2714 = n895 & n2713;
  assign n2715 = ~n895 & ~n2713;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = ~n2704 & n2716;
  assign n2718 = ~n2704 & ~n2716;
  assign n2719 = n2704 & n2716;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = n2449 & n2673;
  assign n2722 = n2627 & n2668;
  assign n2723 = n2446 & n2663;
  assign n2724 = n2443 & n2675;
  assign n2725 = ~n2721 & ~n2723;
  assign n2726 = ~n2724 & n2725;
  assign n2727 = ~n2722 & n2726;
  assign n2728 = n895 & ~n2727;
  assign n2729 = ~n895 & n2727;
  assign n2730 = ~n2728 & ~n2729;
  assign n2731 = ~n656 & ~n2591;
  assign n2732 = ~n2601 & n2731;
  assign n2733 = n2601 & ~n2731;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = n2730 & ~n2734;
  assign n2736 = ~n2730 & n2734;
  assign n2737 = n2452 & n2673;
  assign n2738 = n2548 & n2668;
  assign n2739 = n2449 & n2663;
  assign n2740 = n2446 & n2675;
  assign n2741 = ~n2737 & ~n2739;
  assign n2742 = ~n2740 & n2741;
  assign n2743 = ~n2738 & n2742;
  assign n2744 = n895 & n2743;
  assign n2745 = ~n895 & ~n2743;
  assign n2746 = ~n2744 & ~n2745;
  assign n2747 = ~n656 & n2584;
  assign n2748 = ~n2589 & n2747;
  assign n2749 = n2589 & ~n2747;
  assign n2750 = ~n2748 & ~n2749;
  assign n2751 = n2746 & n2750;
  assign n2752 = ~n2457 & n2662;
  assign n2753 = ~n2457 & n2663;
  assign n2754 = n2460 & n2675;
  assign n2755 = ~n2572 & n2668;
  assign n2756 = ~n2753 & ~n2754;
  assign n2757 = ~n2755 & n2756;
  assign n2758 = ~n895 & ~n2752;
  assign n2759 = n2757 & n2758;
  assign n2760 = ~n2457 & n2673;
  assign n2761 = ~n2595 & n2668;
  assign n2762 = n2460 & n2663;
  assign n2763 = n2452 & n2675;
  assign n2764 = ~n2760 & ~n2762;
  assign n2765 = ~n2763 & n2764;
  assign n2766 = ~n2761 & n2765;
  assign n2767 = n2759 & n2766;
  assign n2768 = n2584 & n2767;
  assign n2769 = ~n2584 & n2767;
  assign n2770 = n2584 & ~n2767;
  assign n2771 = ~n2769 & ~n2770;
  assign n2772 = n2452 & n2663;
  assign n2773 = n2609 & n2668;
  assign n2774 = n2460 & n2673;
  assign n2775 = n2449 & n2675;
  assign n2776 = ~n2772 & ~n2774;
  assign n2777 = ~n2775 & n2776;
  assign n2778 = ~n2773 & n2777;
  assign n2779 = ~n895 & n2778;
  assign n2780 = n895 & ~n2778;
  assign n2781 = ~n2779 & ~n2780;
  assign n2782 = ~n2771 & ~n2781;
  assign n2783 = ~n2768 & ~n2782;
  assign n2784 = ~n2746 & ~n2750;
  assign n2785 = ~n2751 & ~n2784;
  assign n2786 = ~n2783 & n2785;
  assign n2787 = ~n2751 & ~n2786;
  assign n2788 = ~n2736 & n2787;
  assign n2789 = ~n2735 & ~n2788;
  assign n2790 = ~n2720 & n2789;
  assign n2791 = ~n2717 & ~n2790;
  assign n2792 = ~n2701 & n2791;
  assign n2793 = ~n2700 & ~n2792;
  assign n2794 = n2685 & n2793;
  assign n2795 = ~n2683 & ~n2794;
  assign n2796 = ~n2651 & ~n2655;
  assign n2797 = n2446 & n2544;
  assign n2798 = n2546 & n2707;
  assign n2799 = n2443 & n2550;
  assign n2800 = n2440 & n2552;
  assign n2801 = ~n2797 & ~n2799;
  assign n2802 = ~n2800 & n2801;
  assign n2803 = ~n2798 & n2802;
  assign n2804 = ~n656 & ~n2803;
  assign n2805 = n656 & n2803;
  assign n2806 = ~n2804 & ~n2805;
  assign n2807 = n2452 & n2566;
  assign n2808 = n2573 & n2609;
  assign n2809 = n2460 & n2638;
  assign n2810 = n2449 & n2568;
  assign n2811 = ~n2807 & ~n2809;
  assign n2812 = ~n2810 & n2811;
  assign n2813 = ~n2808 & n2812;
  assign n2814 = n636 & ~n2813;
  assign n2815 = ~n636 & n2813;
  assign n2816 = ~n2814 & ~n2815;
  assign n2817 = ~n636 & n2646;
  assign n2818 = n2645 & n2817;
  assign n2819 = ~n2577 & ~n2818;
  assign n2820 = ~n2457 & n2818;
  assign n2821 = ~n2819 & ~n2820;
  assign n2822 = ~n2816 & n2821;
  assign n2823 = n2816 & ~n2821;
  assign n2824 = ~n2822 & ~n2823;
  assign n2825 = n2806 & n2824;
  assign n2826 = ~n2806 & ~n2824;
  assign n2827 = ~n2825 & ~n2826;
  assign n2828 = n2796 & ~n2827;
  assign n2829 = ~n2796 & n2827;
  assign n2830 = ~n2828 & ~n2829;
  assign n2831 = n2437 & n2673;
  assign n2832 = n2483 & ~n2485;
  assign n2833 = ~n2486 & ~n2832;
  assign n2834 = n2668 & n2833;
  assign n2835 = n2434 & n2663;
  assign n2836 = n2431 & n2675;
  assign n2837 = ~n2831 & ~n2835;
  assign n2838 = ~n2836 & n2837;
  assign n2839 = ~n2834 & n2838;
  assign n2840 = n895 & n2839;
  assign n2841 = ~n895 & ~n2839;
  assign n2842 = ~n2840 & ~n2841;
  assign n2843 = n2830 & n2842;
  assign n2844 = ~n2830 & ~n2842;
  assign n2845 = ~n2843 & ~n2844;
  assign n2846 = ~n2795 & n2845;
  assign n2847 = n2795 & ~n2845;
  assign n2848 = ~n2846 & ~n2847;
  assign n2849 = n2533 & n2848;
  assign n2850 = n2431 & n2524;
  assign n2851 = n2491 & ~n2493;
  assign n2852 = ~n2494 & ~n2851;
  assign n2853 = n2426 & n2852;
  assign n2854 = n76 & n2428;
  assign n2855 = n2421 & n2526;
  assign n2856 = ~n2850 & ~n2854;
  assign n2857 = ~n2855 & n2856;
  assign n2858 = ~n2853 & n2857;
  assign n2859 = ~n57 & ~n2858;
  assign n2860 = n57 & n2858;
  assign n2861 = ~n2859 & ~n2860;
  assign n2862 = ~n2685 & ~n2793;
  assign n2863 = ~n2794 & ~n2862;
  assign n2864 = n2861 & n2863;
  assign n2865 = n76 & n2431;
  assign n2866 = n2487 & ~n2489;
  assign n2867 = ~n2490 & ~n2866;
  assign n2868 = n2426 & n2867;
  assign n2869 = n2434 & n2524;
  assign n2870 = n2428 & n2526;
  assign n2871 = ~n2865 & ~n2869;
  assign n2872 = ~n2870 & n2871;
  assign n2873 = ~n2868 & n2872;
  assign n2874 = n57 & n2873;
  assign n2875 = ~n57 & ~n2873;
  assign n2876 = ~n2874 & ~n2875;
  assign n2877 = ~n2700 & ~n2701;
  assign n2878 = n2791 & n2877;
  assign n2879 = ~n2791 & ~n2877;
  assign n2880 = ~n2878 & ~n2879;
  assign n2881 = n2876 & ~n2880;
  assign n2882 = n2720 & n2789;
  assign n2883 = ~n2720 & ~n2789;
  assign n2884 = ~n2882 & ~n2883;
  assign n2885 = n2437 & n2524;
  assign n2886 = n2426 & n2833;
  assign n2887 = n76 & n2434;
  assign n2888 = n2431 & n2526;
  assign n2889 = ~n2885 & ~n2887;
  assign n2890 = ~n2888 & n2889;
  assign n2891 = ~n2886 & n2890;
  assign n2892 = n57 & n2891;
  assign n2893 = ~n57 & ~n2891;
  assign n2894 = ~n2892 & ~n2893;
  assign n2895 = ~n2884 & n2894;
  assign n2896 = n76 & n2437;
  assign n2897 = n2426 & n2670;
  assign n2898 = n2440 & n2524;
  assign n2899 = n2434 & n2526;
  assign n2900 = ~n2896 & ~n2898;
  assign n2901 = ~n2899 & n2900;
  assign n2902 = ~n2897 & n2901;
  assign n2903 = n57 & n2902;
  assign n2904 = ~n57 & ~n2902;
  assign n2905 = ~n2903 & ~n2904;
  assign n2906 = ~n2735 & ~n2736;
  assign n2907 = n2787 & n2906;
  assign n2908 = ~n2787 & ~n2906;
  assign n2909 = ~n2907 & ~n2908;
  assign n2910 = n2905 & ~n2909;
  assign n2911 = n2443 & n2524;
  assign n2912 = n2426 & n2688;
  assign n2913 = n76 & n2440;
  assign n2914 = n2437 & n2526;
  assign n2915 = ~n2911 & ~n2913;
  assign n2916 = ~n2914 & n2915;
  assign n2917 = ~n2912 & n2916;
  assign n2918 = ~n57 & ~n2917;
  assign n2919 = n57 & n2917;
  assign n2920 = ~n2918 & ~n2919;
  assign n2921 = n2783 & ~n2785;
  assign n2922 = ~n2786 & ~n2921;
  assign n2923 = n2920 & n2922;
  assign n2924 = n2446 & n2524;
  assign n2925 = n2426 & n2707;
  assign n2926 = n76 & n2443;
  assign n2927 = n2440 & n2526;
  assign n2928 = ~n2924 & ~n2926;
  assign n2929 = ~n2927 & n2928;
  assign n2930 = ~n2925 & n2929;
  assign n2931 = n57 & n2930;
  assign n2932 = ~n57 & ~n2930;
  assign n2933 = ~n2931 & ~n2932;
  assign n2934 = n2771 & n2781;
  assign n2935 = ~n2782 & ~n2934;
  assign n2936 = n2933 & n2935;
  assign n2937 = n2449 & n2524;
  assign n2938 = n2426 & n2627;
  assign n2939 = n76 & n2446;
  assign n2940 = n2443 & n2526;
  assign n2941 = ~n2937 & ~n2939;
  assign n2942 = ~n2940 & n2941;
  assign n2943 = ~n2938 & n2942;
  assign n2944 = ~n57 & ~n2943;
  assign n2945 = n57 & n2943;
  assign n2946 = ~n2944 & ~n2945;
  assign n2947 = ~n895 & ~n2759;
  assign n2948 = ~n2766 & n2947;
  assign n2949 = n2766 & ~n2947;
  assign n2950 = ~n2948 & ~n2949;
  assign n2951 = n2946 & n2950;
  assign n2952 = n2452 & n2524;
  assign n2953 = n2426 & n2548;
  assign n2954 = n76 & n2449;
  assign n2955 = n2446 & n2526;
  assign n2956 = ~n2952 & ~n2954;
  assign n2957 = ~n2955 & n2956;
  assign n2958 = ~n2953 & n2957;
  assign n2959 = n57 & n2958;
  assign n2960 = ~n57 & ~n2958;
  assign n2961 = ~n2959 & ~n2960;
  assign n2962 = ~n895 & n2752;
  assign n2963 = ~n2757 & n2962;
  assign n2964 = n2757 & ~n2962;
  assign n2965 = ~n2963 & ~n2964;
  assign n2966 = n2961 & n2965;
  assign n2967 = n68 & ~n2457;
  assign n2968 = n76 & ~n2457;
  assign n2969 = n2460 & n2526;
  assign n2970 = n2426 & ~n2572;
  assign n2971 = ~n2968 & ~n2969;
  assign n2972 = ~n2970 & n2971;
  assign n2973 = ~n57 & ~n2967;
  assign n2974 = n2972 & n2973;
  assign n2975 = ~n2457 & n2524;
  assign n2976 = n2426 & ~n2595;
  assign n2977 = n76 & n2460;
  assign n2978 = n2452 & n2526;
  assign n2979 = ~n2975 & ~n2977;
  assign n2980 = ~n2978 & n2979;
  assign n2981 = ~n2976 & n2980;
  assign n2982 = n2974 & n2981;
  assign n2983 = n2752 & n2982;
  assign n2984 = ~n2752 & n2982;
  assign n2985 = n2752 & ~n2982;
  assign n2986 = ~n2984 & ~n2985;
  assign n2987 = n76 & n2452;
  assign n2988 = n2426 & n2609;
  assign n2989 = n2460 & n2524;
  assign n2990 = n2449 & n2526;
  assign n2991 = ~n2987 & ~n2989;
  assign n2992 = ~n2990 & n2991;
  assign n2993 = ~n2988 & n2992;
  assign n2994 = ~n57 & ~n2993;
  assign n2995 = n57 & n2993;
  assign n2996 = ~n2994 & ~n2995;
  assign n2997 = ~n2986 & n2996;
  assign n2998 = ~n2983 & ~n2997;
  assign n2999 = ~n2961 & ~n2965;
  assign n3000 = ~n2966 & ~n2999;
  assign n3001 = ~n2998 & n3000;
  assign n3002 = ~n2966 & ~n3001;
  assign n3003 = ~n2946 & ~n2950;
  assign n3004 = ~n2951 & ~n3003;
  assign n3005 = ~n3002 & n3004;
  assign n3006 = ~n2951 & ~n3005;
  assign n3007 = ~n2933 & ~n2935;
  assign n3008 = ~n2936 & ~n3007;
  assign n3009 = ~n3006 & n3008;
  assign n3010 = ~n2936 & ~n3009;
  assign n3011 = ~n2920 & ~n2922;
  assign n3012 = ~n2923 & ~n3011;
  assign n3013 = ~n3010 & n3012;
  assign n3014 = ~n2923 & ~n3013;
  assign n3015 = ~n2905 & n2909;
  assign n3016 = ~n2910 & ~n3015;
  assign n3017 = ~n3014 & n3016;
  assign n3018 = ~n2910 & ~n3017;
  assign n3019 = ~n2884 & ~n2894;
  assign n3020 = n2884 & n2894;
  assign n3021 = ~n3019 & ~n3020;
  assign n3022 = ~n3018 & ~n3021;
  assign n3023 = ~n2895 & ~n3022;
  assign n3024 = ~n2876 & n2880;
  assign n3025 = ~n2881 & ~n3024;
  assign n3026 = ~n3023 & n3025;
  assign n3027 = ~n2881 & ~n3026;
  assign n3028 = ~n2861 & ~n2863;
  assign n3029 = ~n2864 & ~n3028;
  assign n3030 = ~n3027 & n3029;
  assign n3031 = ~n2864 & ~n3030;
  assign n3032 = ~n2533 & ~n2848;
  assign n3033 = ~n2849 & ~n3032;
  assign n3034 = ~n3031 & n3033;
  assign n3035 = ~n2849 & ~n3034;
  assign n3036 = n2421 & n2524;
  assign n3037 = ~n2516 & ~n2519;
  assign n3038 = ~n133 & ~n478;
  assign n3039 = ~n479 & n3038;
  assign n3040 = ~n563 & ~n657;
  assign n3041 = ~n266 & ~n346;
  assign n3042 = n341 & n3041;
  assign n3043 = ~n156 & ~n336;
  assign n3044 = ~n353 & ~n450;
  assign n3045 = ~n818 & n3044;
  assign n3046 = n3043 & n3045;
  assign n3047 = ~n142 & ~n430;
  assign n3048 = ~n193 & ~n216;
  assign n3049 = ~n286 & ~n328;
  assign n3050 = ~n377 & ~n548;
  assign n3051 = n3049 & n3050;
  assign n3052 = n3040 & n3048;
  assign n3053 = n3047 & n3052;
  assign n3054 = n2044 & n3051;
  assign n3055 = n3042 & n3054;
  assign n3056 = n3046 & n3053;
  assign n3057 = n3055 & n3056;
  assign n3058 = ~n291 & ~n348;
  assign n3059 = ~n303 & ~n327;
  assign n3060 = ~n362 & ~n420;
  assign n3061 = ~n546 & ~n566;
  assign n3062 = n3060 & n3061;
  assign n3063 = n436 & n3059;
  assign n3064 = n3058 & n3063;
  assign n3065 = n2203 & n3062;
  assign n3066 = n3039 & n3065;
  assign n3067 = n185 & n3064;
  assign n3068 = n3066 & n3067;
  assign n3069 = n265 & n3068;
  assign n3070 = n3057 & n3069;
  assign n3071 = ~n2513 & n3070;
  assign n3072 = n2513 & ~n3070;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = ~n2515 & n3073;
  assign n3075 = n2515 & n3070;
  assign n3076 = ~n3074 & ~n3075;
  assign n3077 = ~n3037 & n3076;
  assign n3078 = n3037 & ~n3076;
  assign n3079 = ~n3077 & ~n3078;
  assign n3080 = n2426 & n3079;
  assign n3081 = n76 & ~n2515;
  assign n3082 = n2526 & n3073;
  assign n3083 = ~n3036 & ~n3081;
  assign n3084 = ~n3082 & n3083;
  assign n3085 = ~n3080 & n3084;
  assign n3086 = ~n57 & ~n3085;
  assign n3087 = n57 & n3085;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = ~n2843 & ~n2846;
  assign n3090 = n2431 & n2663;
  assign n3091 = n2668 & n2867;
  assign n3092 = n2434 & n2673;
  assign n3093 = n2428 & n2675;
  assign n3094 = ~n3090 & ~n3092;
  assign n3095 = ~n3093 & n3094;
  assign n3096 = ~n3091 & n3095;
  assign n3097 = n895 & n3096;
  assign n3098 = ~n895 & ~n3096;
  assign n3099 = ~n3097 & ~n3098;
  assign n3100 = ~n2825 & ~n2829;
  assign n3101 = n2443 & n2544;
  assign n3102 = n2546 & n2688;
  assign n3103 = n2440 & n2550;
  assign n3104 = n2437 & n2552;
  assign n3105 = ~n3101 & ~n3103;
  assign n3106 = ~n3104 & n3105;
  assign n3107 = ~n3102 & n3106;
  assign n3108 = ~n656 & ~n3107;
  assign n3109 = n656 & n3107;
  assign n3110 = ~n3108 & ~n3109;
  assign n3111 = ~n2820 & ~n2822;
  assign n3112 = n2452 & n2638;
  assign n3113 = n2548 & n2573;
  assign n3114 = n2449 & n2566;
  assign n3115 = n2446 & n2568;
  assign n3116 = ~n3112 & ~n3114;
  assign n3117 = ~n3115 & n3116;
  assign n3118 = ~n3113 & n3117;
  assign n3119 = ~n636 & ~n2460;
  assign n3120 = ~n3118 & n3119;
  assign n3121 = n3118 & ~n3119;
  assign n3122 = ~n3120 & ~n3121;
  assign n3123 = ~n3111 & n3122;
  assign n3124 = n3111 & ~n3122;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = n3110 & n3125;
  assign n3127 = ~n3110 & ~n3125;
  assign n3128 = ~n3126 & ~n3127;
  assign n3129 = ~n3100 & n3128;
  assign n3130 = n3100 & ~n3128;
  assign n3131 = ~n3129 & ~n3130;
  assign n3132 = n3099 & n3131;
  assign n3133 = ~n3099 & ~n3131;
  assign n3134 = ~n3132 & ~n3133;
  assign n3135 = ~n3089 & n3134;
  assign n3136 = n3089 & ~n3134;
  assign n3137 = ~n3135 & ~n3136;
  assign n3138 = n3088 & n3137;
  assign n3139 = ~n3088 & ~n3137;
  assign n3140 = ~n3138 & ~n3139;
  assign n3141 = ~n3035 & n3140;
  assign n3142 = n3035 & ~n3140;
  assign n3143 = ~n3141 & ~n3142;
  assign n3144 = n2513 & n3070;
  assign n3145 = ~n129 & ~n138;
  assign n3146 = ~n228 & ~n236;
  assign n3147 = ~n317 & ~n822;
  assign n3148 = n3146 & n3147;
  assign n3149 = n321 & n3145;
  assign n3150 = n856 & n2271;
  assign n3151 = n3149 & n3150;
  assign n3152 = n3148 & n3151;
  assign n3153 = n2095 & n2182;
  assign n3154 = n3152 & n3153;
  assign n3155 = n604 & n3154;
  assign n3156 = n521 & n3155;
  assign n3157 = n3144 & n3156;
  assign n3158 = ~n3144 & ~n3156;
  assign n3159 = ~n3157 & ~n3158;
  assign n3160 = pi2  & n50;
  assign n3161 = ~n3159 & n3160;
  assign n3162 = pi0  & ~pi22 ;
  assign n3163 = pi1  & ~n3162;
  assign n3164 = ~pi1  & n3162;
  assign n3165 = ~n3163 & ~n3164;
  assign n3166 = n65 & n3165;
  assign n3167 = ~n65 & ~n3165;
  assign n3168 = ~n3166 & ~n3167;
  assign n3169 = pi0  & n3168;
  assign n3170 = ~n272 & ~n299;
  assign n3171 = n481 & n609;
  assign n3172 = n3170 & n3171;
  assign n3173 = n477 & n1063;
  assign n3174 = n3172 & n3173;
  assign n3175 = n496 & n615;
  assign n3176 = n3174 & n3175;
  assign n3177 = n514 & n604;
  assign n3178 = n664 & n3177;
  assign n3179 = n3176 & n3178;
  assign n3180 = ~n3157 & n3179;
  assign n3181 = n3157 & ~n3179;
  assign n3182 = ~n3180 & ~n3181;
  assign n3183 = ~n3159 & n3182;
  assign n3184 = n3073 & ~n3159;
  assign n3185 = ~n3074 & ~n3077;
  assign n3186 = ~n3073 & n3156;
  assign n3187 = ~n3184 & ~n3186;
  assign n3188 = ~n3185 & n3187;
  assign n3189 = ~n3184 & ~n3188;
  assign n3190 = n3159 & n3179;
  assign n3191 = ~n3183 & ~n3190;
  assign n3192 = ~n3189 & n3191;
  assign n3193 = ~n3183 & ~n3192;
  assign n3194 = n3157 & n3179;
  assign n3195 = ~n244 & n665;
  assign n3196 = ~n198 & ~n616;
  assign n3197 = n489 & n3196;
  assign n3198 = n507 & n604;
  assign n3199 = n673 & n3198;
  assign n3200 = n3197 & n3199;
  assign n3201 = n3195 & n3200;
  assign n3202 = ~n3194 & ~n3201;
  assign n3203 = n3194 & n3201;
  assign n3204 = ~n3202 & ~n3203;
  assign n3205 = n3182 & ~n3204;
  assign n3206 = ~n3182 & n3201;
  assign n3207 = ~n3205 & ~n3206;
  assign n3208 = ~n3193 & n3207;
  assign n3209 = n3193 & ~n3207;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = n3169 & n3210;
  assign n3212 = ~pi0  & ~n3165;
  assign n3213 = n3182 & n3212;
  assign n3214 = pi0  & ~n3168;
  assign n3215 = ~n3204 & n3214;
  assign n3216 = ~n3161 & ~n3213;
  assign n3217 = ~n3215 & n3216;
  assign n3218 = ~n3211 & n3217;
  assign n3219 = n65 & n3218;
  assign n3220 = ~n65 & ~n3218;
  assign n3221 = ~n3219 & ~n3220;
  assign n3222 = n3143 & n3221;
  assign n3223 = n3031 & ~n3033;
  assign n3224 = ~n3034 & ~n3223;
  assign n3225 = n3073 & n3160;
  assign n3226 = n3189 & ~n3191;
  assign n3227 = ~n3192 & ~n3226;
  assign n3228 = n3169 & n3227;
  assign n3229 = ~n3159 & n3212;
  assign n3230 = n3182 & n3214;
  assign n3231 = ~n3225 & ~n3229;
  assign n3232 = ~n3230 & n3231;
  assign n3233 = ~n3228 & n3232;
  assign n3234 = n65 & n3233;
  assign n3235 = ~n65 & ~n3233;
  assign n3236 = ~n3234 & ~n3235;
  assign n3237 = n3224 & n3236;
  assign n3238 = n3027 & ~n3029;
  assign n3239 = ~n3030 & ~n3238;
  assign n3240 = ~n2515 & n3160;
  assign n3241 = n3185 & ~n3187;
  assign n3242 = ~n3188 & ~n3241;
  assign n3243 = n3169 & n3242;
  assign n3244 = n3073 & n3212;
  assign n3245 = ~n3159 & n3214;
  assign n3246 = ~n3240 & ~n3244;
  assign n3247 = ~n3245 & n3246;
  assign n3248 = ~n3243 & n3247;
  assign n3249 = n65 & n3248;
  assign n3250 = ~n65 & ~n3248;
  assign n3251 = ~n3249 & ~n3250;
  assign n3252 = n3239 & n3251;
  assign n3253 = ~n3239 & ~n3251;
  assign n3254 = ~n3252 & ~n3253;
  assign n3255 = n3023 & ~n3025;
  assign n3256 = ~n3026 & ~n3255;
  assign n3257 = n3018 & n3021;
  assign n3258 = ~n3022 & ~n3257;
  assign n3259 = n3014 & ~n3016;
  assign n3260 = ~n3017 & ~n3259;
  assign n3261 = n3010 & ~n3012;
  assign n3262 = ~n3013 & ~n3261;
  assign n3263 = n3006 & ~n3008;
  assign n3264 = ~n3009 & ~n3263;
  assign n3265 = n3002 & ~n3004;
  assign n3266 = ~n3005 & ~n3265;
  assign n3267 = n2998 & ~n3000;
  assign n3268 = ~n3001 & ~n3267;
  assign n3269 = n2446 & n3160;
  assign n3270 = n2707 & n3169;
  assign n3271 = n2443 & n3212;
  assign n3272 = n2440 & n3214;
  assign n3273 = ~n3269 & ~n3271;
  assign n3274 = ~n3272 & n3273;
  assign n3275 = ~n3270 & n3274;
  assign n3276 = n65 & ~n3275;
  assign n3277 = ~n65 & n3275;
  assign n3278 = ~n3276 & ~n3277;
  assign n3279 = ~n57 & ~n2974;
  assign n3280 = ~n2981 & n3279;
  assign n3281 = n2981 & ~n3279;
  assign n3282 = ~n3280 & ~n3281;
  assign n3283 = ~n57 & n2967;
  assign n3284 = ~n2972 & n3283;
  assign n3285 = n2972 & ~n3283;
  assign n3286 = ~n3284 & ~n3285;
  assign n3287 = ~n50 & ~n2457;
  assign n3288 = ~n2457 & n3160;
  assign n3289 = n2460 & n3212;
  assign n3290 = n2452 & n3214;
  assign n3291 = ~n3288 & ~n3289;
  assign n3292 = ~n3290 & n3291;
  assign n3293 = ~n65 & ~n3292;
  assign n3294 = ~n2452 & n2572;
  assign n3295 = ~n65 & n3169;
  assign n3296 = ~n3294 & n3295;
  assign n3297 = n2460 & n3214;
  assign n3298 = ~n65 & ~n3287;
  assign n3299 = ~n3297 & n3298;
  assign n3300 = ~n3296 & n3299;
  assign n3301 = ~n3293 & n3300;
  assign n3302 = n2967 & n3301;
  assign n3303 = ~n2967 & ~n3301;
  assign n3304 = n2452 & n3212;
  assign n3305 = n2609 & n3169;
  assign n3306 = n2449 & n3214;
  assign n3307 = ~n3304 & ~n3306;
  assign n3308 = ~n3305 & n3307;
  assign n3309 = n65 & ~n3308;
  assign n3310 = n50 & n2460;
  assign n3311 = ~n65 & ~n3310;
  assign n3312 = n3308 & n3311;
  assign n3313 = ~n3309 & ~n3312;
  assign n3314 = ~n3303 & ~n3313;
  assign n3315 = ~n3302 & ~n3314;
  assign n3316 = n3286 & ~n3315;
  assign n3317 = ~n3286 & n3315;
  assign n3318 = n2452 & n3160;
  assign n3319 = n2548 & n3169;
  assign n3320 = n2449 & n3212;
  assign n3321 = n2446 & n3214;
  assign n3322 = ~n3318 & ~n3320;
  assign n3323 = ~n3321 & n3322;
  assign n3324 = ~n3319 & n3323;
  assign n3325 = ~n65 & ~n3324;
  assign n3326 = n65 & n3324;
  assign n3327 = ~n3325 & ~n3326;
  assign n3328 = ~n3317 & n3327;
  assign n3329 = ~n3316 & ~n3328;
  assign n3330 = ~n3282 & n3329;
  assign n3331 = n3282 & ~n3329;
  assign n3332 = n2449 & n3160;
  assign n3333 = n2627 & n3169;
  assign n3334 = n2446 & n3212;
  assign n3335 = n2443 & n3214;
  assign n3336 = ~n3332 & ~n3334;
  assign n3337 = ~n3335 & n3336;
  assign n3338 = ~n3333 & n3337;
  assign n3339 = n65 & ~n3338;
  assign n3340 = ~n65 & n3338;
  assign n3341 = ~n3339 & ~n3340;
  assign n3342 = ~n3331 & n3341;
  assign n3343 = ~n3330 & ~n3342;
  assign n3344 = ~n3278 & n3343;
  assign n3345 = n3278 & ~n3343;
  assign n3346 = n2986 & ~n2996;
  assign n3347 = ~n2997 & ~n3346;
  assign n3348 = ~n3345 & n3347;
  assign n3349 = ~n3344 & ~n3348;
  assign n3350 = ~n3268 & n3349;
  assign n3351 = n3268 & ~n3349;
  assign n3352 = n2443 & n3160;
  assign n3353 = n2688 & n3169;
  assign n3354 = n2440 & n3212;
  assign n3355 = n2437 & n3214;
  assign n3356 = ~n3352 & ~n3354;
  assign n3357 = ~n3355 & n3356;
  assign n3358 = ~n3353 & n3357;
  assign n3359 = n65 & ~n3358;
  assign n3360 = ~n65 & n3358;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 = ~n3351 & n3361;
  assign n3363 = ~n3350 & ~n3362;
  assign n3364 = n3266 & n3363;
  assign n3365 = ~n3266 & ~n3363;
  assign n3366 = n2434 & n3214;
  assign n3367 = n2670 & n3169;
  assign n3368 = n2437 & n3212;
  assign n3369 = ~n3366 & ~n3368;
  assign n3370 = ~n3367 & n3369;
  assign n3371 = n65 & ~n3370;
  assign n3372 = n2440 & n3160;
  assign n3373 = ~n65 & ~n3372;
  assign n3374 = n3370 & n3373;
  assign n3375 = ~n3371 & ~n3374;
  assign n3376 = ~n3365 & ~n3375;
  assign n3377 = ~n3364 & ~n3376;
  assign n3378 = n3264 & ~n3377;
  assign n3379 = ~n3264 & n3377;
  assign n3380 = n2437 & n3160;
  assign n3381 = n2833 & n3169;
  assign n3382 = n2434 & n3212;
  assign n3383 = n2431 & n3214;
  assign n3384 = ~n3380 & ~n3382;
  assign n3385 = ~n3383 & n3384;
  assign n3386 = ~n3381 & n3385;
  assign n3387 = ~n65 & ~n3386;
  assign n3388 = n65 & n3386;
  assign n3389 = ~n3387 & ~n3388;
  assign n3390 = ~n3379 & n3389;
  assign n3391 = ~n3378 & ~n3390;
  assign n3392 = n3262 & ~n3391;
  assign n3393 = ~n3262 & n3391;
  assign n3394 = n2428 & n3214;
  assign n3395 = n2867 & n3169;
  assign n3396 = n2431 & n3212;
  assign n3397 = ~n3394 & ~n3396;
  assign n3398 = ~n3395 & n3397;
  assign n3399 = n65 & ~n3398;
  assign n3400 = n2434 & n3160;
  assign n3401 = ~n65 & ~n3400;
  assign n3402 = n3398 & n3401;
  assign n3403 = ~n3399 & ~n3402;
  assign n3404 = ~n3393 & ~n3403;
  assign n3405 = ~n3392 & ~n3404;
  assign n3406 = ~n3260 & n3405;
  assign n3407 = n3260 & ~n3405;
  assign n3408 = n2431 & n3160;
  assign n3409 = n2852 & n3169;
  assign n3410 = n2428 & n3212;
  assign n3411 = n2421 & n3214;
  assign n3412 = ~n3408 & ~n3410;
  assign n3413 = ~n3411 & n3412;
  assign n3414 = ~n3409 & n3413;
  assign n3415 = n65 & ~n3414;
  assign n3416 = ~n65 & n3414;
  assign n3417 = ~n3415 & ~n3416;
  assign n3418 = ~n3407 & n3417;
  assign n3419 = ~n3406 & ~n3418;
  assign n3420 = n3258 & n3419;
  assign n3421 = ~n3258 & ~n3419;
  assign n3422 = ~n2515 & n3214;
  assign n3423 = n2521 & n3169;
  assign n3424 = n2421 & n3212;
  assign n3425 = ~n3422 & ~n3424;
  assign n3426 = ~n3423 & n3425;
  assign n3427 = n65 & ~n3426;
  assign n3428 = n2428 & n3160;
  assign n3429 = ~n65 & ~n3428;
  assign n3430 = n3426 & n3429;
  assign n3431 = ~n3427 & ~n3430;
  assign n3432 = ~n3421 & ~n3431;
  assign n3433 = ~n3420 & ~n3432;
  assign n3434 = ~n3256 & n3433;
  assign n3435 = n3256 & ~n3433;
  assign n3436 = n2421 & n3160;
  assign n3437 = n3079 & n3169;
  assign n3438 = ~n2515 & n3212;
  assign n3439 = n3073 & n3214;
  assign n3440 = ~n3436 & ~n3438;
  assign n3441 = ~n3439 & n3440;
  assign n3442 = ~n3437 & n3441;
  assign n3443 = n65 & ~n3442;
  assign n3444 = ~n65 & n3442;
  assign n3445 = ~n3443 & ~n3444;
  assign n3446 = ~n3435 & n3445;
  assign n3447 = ~n3434 & ~n3446;
  assign n3448 = n3254 & n3447;
  assign n3449 = ~n3252 & ~n3448;
  assign n3450 = ~n3224 & ~n3236;
  assign n3451 = ~n3237 & ~n3450;
  assign n3452 = ~n3449 & n3451;
  assign n3453 = ~n3237 & ~n3452;
  assign n3454 = ~n3143 & ~n3221;
  assign n3455 = ~n3222 & ~n3454;
  assign n3456 = ~n3453 & n3455;
  assign n3457 = ~n3222 & ~n3456;
  assign n3458 = n3160 & n3182;
  assign n3459 = ~n3205 & ~n3208;
  assign n3460 = ~n144 & ~n228;
  assign n3461 = ~n168 & ~n243;
  assign n3462 = ~n429 & ~n479;
  assign n3463 = n3461 & n3462;
  assign n3464 = n454 & n2103;
  assign n3465 = n3460 & n3464;
  assign n3466 = n3463 & n3465;
  assign n3467 = ~n194 & ~n233;
  assign n3468 = ~n253 & ~n254;
  assign n3469 = ~n289 & n3468;
  assign n3470 = n971 & n3467;
  assign n3471 = n2089 & n2271;
  assign n3472 = n3470 & n3471;
  assign n3473 = n452 & n3469;
  assign n3474 = n3472 & n3473;
  assign n3475 = n2389 & n3474;
  assign n3476 = n3466 & n3475;
  assign n3477 = n1060 & n3476;
  assign n3478 = ~n3203 & n3477;
  assign n3479 = n3203 & ~n3477;
  assign n3480 = ~n3478 & ~n3479;
  assign n3481 = ~n3204 & n3480;
  assign n3482 = n3204 & n3477;
  assign n3483 = ~n3481 & ~n3482;
  assign n3484 = ~n3459 & n3483;
  assign n3485 = n3459 & ~n3483;
  assign n3486 = ~n3484 & ~n3485;
  assign n3487 = n3169 & n3486;
  assign n3488 = ~n3204 & n3212;
  assign n3489 = n3214 & n3480;
  assign n3490 = ~n3458 & ~n3488;
  assign n3491 = ~n3489 & n3490;
  assign n3492 = ~n3487 & n3491;
  assign n3493 = n65 & ~n3492;
  assign n3494 = ~n65 & n3492;
  assign n3495 = ~n3493 & ~n3494;
  assign n3496 = ~n3138 & ~n3141;
  assign n3497 = ~n3132 & ~n3135;
  assign n3498 = n2431 & n2673;
  assign n3499 = n2668 & n2852;
  assign n3500 = n2428 & n2663;
  assign n3501 = n2421 & n2675;
  assign n3502 = ~n3498 & ~n3500;
  assign n3503 = ~n3501 & n3502;
  assign n3504 = ~n3499 & n3503;
  assign n3505 = n895 & ~n3504;
  assign n3506 = ~n895 & n3504;
  assign n3507 = ~n3505 & ~n3506;
  assign n3508 = ~n3126 & ~n3129;
  assign n3509 = ~n636 & ~n2452;
  assign n3510 = n2449 & n2638;
  assign n3511 = n2573 & n2627;
  assign n3512 = n2446 & n2566;
  assign n3513 = n2443 & n2568;
  assign n3514 = ~n3510 & ~n3512;
  assign n3515 = ~n3513 & n3514;
  assign n3516 = ~n3511 & n3515;
  assign n3517 = n3509 & ~n3516;
  assign n3518 = ~n3509 & n3516;
  assign n3519 = ~n3517 & ~n3518;
  assign n3520 = ~n636 & n2460;
  assign n3521 = n3118 & n3520;
  assign n3522 = ~n3123 & ~n3521;
  assign n3523 = n3519 & ~n3522;
  assign n3524 = ~n3519 & n3522;
  assign n3525 = ~n3523 & ~n3524;
  assign n3526 = n2437 & n2550;
  assign n3527 = n2546 & n2670;
  assign n3528 = n2440 & n2544;
  assign n3529 = n2434 & n2552;
  assign n3530 = ~n3526 & ~n3528;
  assign n3531 = ~n3529 & n3530;
  assign n3532 = ~n3527 & n3531;
  assign n3533 = n656 & n3532;
  assign n3534 = ~n656 & ~n3532;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = n3525 & n3535;
  assign n3537 = ~n3525 & ~n3535;
  assign n3538 = ~n3536 & ~n3537;
  assign n3539 = ~n3508 & n3538;
  assign n3540 = n3508 & ~n3538;
  assign n3541 = ~n3539 & ~n3540;
  assign n3542 = ~n3507 & n3541;
  assign n3543 = n3507 & ~n3541;
  assign n3544 = ~n3542 & ~n3543;
  assign n3545 = n3497 & ~n3544;
  assign n3546 = ~n3497 & n3544;
  assign n3547 = ~n3545 & ~n3546;
  assign n3548 = ~n2515 & n2524;
  assign n3549 = n2426 & n3242;
  assign n3550 = n76 & n3073;
  assign n3551 = n2526 & ~n3159;
  assign n3552 = ~n3548 & ~n3550;
  assign n3553 = ~n3551 & n3552;
  assign n3554 = ~n3549 & n3553;
  assign n3555 = n57 & n3554;
  assign n3556 = ~n57 & ~n3554;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = n3547 & n3557;
  assign n3559 = ~n3547 & ~n3557;
  assign n3560 = ~n3558 & ~n3559;
  assign n3561 = ~n3496 & n3560;
  assign n3562 = n3496 & ~n3560;
  assign n3563 = ~n3561 & ~n3562;
  assign n3564 = ~n3495 & n3563;
  assign n3565 = n3495 & ~n3563;
  assign n3566 = ~n3564 & ~n3565;
  assign n3567 = n3457 & ~n3566;
  assign n3568 = ~n3457 & n3566;
  assign n3569 = ~n3567 & ~n3568;
  assign n3570 = ~n195 & ~n241;
  assign n3571 = ~n497 & n3570;
  assign n3572 = n333 & n3460;
  assign n3573 = n3571 & n3572;
  assign n3574 = n988 & n1324;
  assign n3575 = n3039 & n3574;
  assign n3576 = n557 & n3573;
  assign n3577 = n3575 & n3576;
  assign n3578 = n374 & n3577;
  assign n3579 = n2150 & n3578;
  assign n3580 = ~n3569 & n3579;
  assign n3581 = n3569 & ~n3579;
  assign n3582 = ~n3580 & ~n3581;
  assign n3583 = n3453 & ~n3455;
  assign n3584 = ~n3456 & ~n3583;
  assign n3585 = ~n167 & ~n204;
  assign n3586 = n508 & n3585;
  assign n3587 = n402 & n3586;
  assign n3588 = n3046 & n3587;
  assign n3589 = ~n236 & ~n548;
  assign n3590 = ~n267 & ~n289;
  assign n3591 = ~n362 & ~n616;
  assign n3592 = n3590 & n3591;
  assign n3593 = n2240 & n3592;
  assign n3594 = ~n199 & ~n240;
  assign n3595 = ~n194 & ~n255;
  assign n3596 = ~n420 & ~n475;
  assign n3597 = n3595 & n3596;
  assign n3598 = n449 & n2077;
  assign n3599 = n3460 & n3594;
  assign n3600 = n3598 & n3599;
  assign n3601 = n3597 & n3600;
  assign n3602 = n3593 & n3601;
  assign n3603 = ~n253 & ~n271;
  assign n3604 = n3589 & n3603;
  assign n3605 = n3602 & n3604;
  assign n3606 = ~n337 & n3039;
  assign n3607 = ~n168 & ~n285;
  assign n3608 = ~n304 & ~n343;
  assign n3609 = n3607 & n3608;
  assign n3610 = n538 & n2390;
  assign n3611 = n3047 & n3610;
  assign n3612 = n3609 & n3611;
  assign n3613 = n3606 & n3612;
  assign n3614 = n446 & n3613;
  assign n3615 = n3588 & n3614;
  assign n3616 = n3605 & n3615;
  assign n3617 = ~n3584 & n3616;
  assign n3618 = n3584 & ~n3616;
  assign n3619 = n3449 & ~n3451;
  assign n3620 = ~n3452 & ~n3619;
  assign n3621 = ~n162 & ~n177;
  assign n3622 = ~n355 & ~n378;
  assign n3623 = ~n430 & n3622;
  assign n3624 = n3621 & n3623;
  assign n3625 = ~n150 & ~n201;
  assign n3626 = ~n217 & ~n252;
  assign n3627 = n3625 & n3626;
  assign n3628 = n298 & n333;
  assign n3629 = n3058 & n3628;
  assign n3630 = n3627 & n3629;
  assign n3631 = n3624 & n3630;
  assign n3632 = ~n214 & ~n229;
  assign n3633 = ~n255 & ~n391;
  assign n3634 = ~n497 & n3633;
  assign n3635 = n2185 & n3632;
  assign n3636 = n345 & n3635;
  assign n3637 = n2213 & n3634;
  assign n3638 = n3636 & n3637;
  assign n3639 = n1029 & n3638;
  assign n3640 = ~n234 & ~n296;
  assign n3641 = n331 & n3640;
  assign n3642 = n3639 & n3641;
  assign n3643 = ~n129 & ~n202;
  assign n3644 = ~n212 & ~n268;
  assign n3645 = ~n315 & n3644;
  assign n3646 = n840 & n3643;
  assign n3647 = n861 & n3040;
  assign n3648 = n3646 & n3647;
  assign n3649 = n3645 & n3648;
  assign n3650 = n2303 & n3649;
  assign n3651 = n3631 & n3650;
  assign n3652 = n3642 & n3651;
  assign n3653 = ~n3620 & n3652;
  assign n3654 = n3620 & ~n3652;
  assign n3655 = ~n212 & ~n352;
  assign n3656 = n325 & n3655;
  assign n3657 = n2385 & n3656;
  assign n3658 = ~n180 & ~n327;
  assign n3659 = ~n340 & ~n358;
  assign n3660 = n3658 & n3659;
  assign n3661 = n481 & n3660;
  assign n3662 = n2128 & n3661;
  assign n3663 = n2160 & n3662;
  assign n3664 = ~n193 & ~n273;
  assign n3665 = ~n348 & ~n360;
  assign n3666 = ~n396 & n3665;
  assign n3667 = n564 & n3664;
  assign n3668 = n608 & n2268;
  assign n3669 = n2270 & n3594;
  assign n3670 = n3668 & n3669;
  assign n3671 = n3666 & n3667;
  assign n3672 = n3670 & n3671;
  assign n3673 = n2227 & n3672;
  assign n3674 = n3657 & n3673;
  assign n3675 = n3663 & n3674;
  assign n3676 = ~n3254 & ~n3447;
  assign n3677 = ~n3448 & ~n3675;
  assign n3678 = ~n3676 & n3677;
  assign n3679 = ~n3654 & ~n3678;
  assign n3680 = ~n3653 & ~n3679;
  assign n3681 = ~n3618 & ~n3680;
  assign n3682 = ~n3617 & ~n3681;
  assign n3683 = n3582 & n3682;
  assign n3684 = ~n3582 & ~n3682;
  assign n3685 = ~n3683 & ~n3684;
  assign n3686 = ~n3617 & ~n3618;
  assign n3687 = n3680 & ~n3686;
  assign n3688 = ~n3680 & n3686;
  assign n3689 = ~n3687 & ~n3688;
  assign n3690 = n3685 & n3689;
  assign n3691 = ~n3685 & ~n3689;
  assign po0  = n3690 | n3691;
  assign n3693 = ~n3581 & ~n3683;
  assign n3694 = ~n3564 & ~n3568;
  assign n3695 = n3160 & ~n3204;
  assign n3696 = ~n3481 & ~n3484;
  assign n3697 = ~n204 & ~n337;
  assign n3698 = n235 & n3697;
  assign n3699 = n398 & n2077;
  assign n3700 = n2268 & n3699;
  assign n3701 = n3698 & n3700;
  assign n3702 = n620 & n3701;
  assign n3703 = ~n175 & ~n202;
  assign n3704 = ~n346 & ~n404;
  assign n3705 = n3703 & n3704;
  assign n3706 = n406 & n797;
  assign n3707 = n856 & n3706;
  assign n3708 = n3705 & n3707;
  assign n3709 = n326 & n3708;
  assign n3710 = n1347 & n3709;
  assign n3711 = n3702 & n3710;
  assign n3712 = n2283 & n3711;
  assign n3713 = ~n3480 & ~n3712;
  assign n3714 = n3203 & n3477;
  assign n3715 = n3712 & ~n3714;
  assign n3716 = ~n3712 & n3714;
  assign n3717 = ~n3715 & ~n3716;
  assign n3718 = n3480 & ~n3717;
  assign n3719 = ~n3713 & ~n3718;
  assign n3720 = ~n3696 & ~n3719;
  assign n3721 = n3696 & n3719;
  assign n3722 = ~n3720 & ~n3721;
  assign n3723 = n3169 & n3722;
  assign n3724 = n3212 & n3480;
  assign n3725 = n3214 & n3717;
  assign n3726 = ~n3695 & ~n3724;
  assign n3727 = ~n3725 & n3726;
  assign n3728 = ~n3723 & n3727;
  assign n3729 = n65 & ~n3728;
  assign n3730 = ~n65 & n3728;
  assign n3731 = ~n3729 & ~n3730;
  assign n3732 = ~n3558 & ~n3561;
  assign n3733 = ~n3542 & ~n3546;
  assign n3734 = n2421 & n2663;
  assign n3735 = n2521 & n2668;
  assign n3736 = n2428 & n2673;
  assign n3737 = ~n2515 & n2675;
  assign n3738 = ~n3734 & ~n3736;
  assign n3739 = ~n3737 & n3738;
  assign n3740 = ~n3735 & n3739;
  assign n3741 = n895 & ~n3740;
  assign n3742 = ~n895 & n3740;
  assign n3743 = ~n3741 & ~n3742;
  assign n3744 = ~n3536 & ~n3539;
  assign n3745 = ~n636 & ~n2449;
  assign n3746 = n2446 & n2638;
  assign n3747 = n2573 & n2707;
  assign n3748 = n2443 & n2566;
  assign n3749 = n2440 & n2568;
  assign n3750 = ~n3746 & ~n3748;
  assign n3751 = ~n3749 & n3750;
  assign n3752 = ~n3747 & n3751;
  assign n3753 = n3745 & ~n3752;
  assign n3754 = ~n3745 & n3752;
  assign n3755 = ~n3753 & ~n3754;
  assign n3756 = ~n636 & n2452;
  assign n3757 = n3516 & n3756;
  assign n3758 = ~n3523 & ~n3757;
  assign n3759 = ~n3755 & ~n3758;
  assign n3760 = n3755 & n3758;
  assign n3761 = ~n3759 & ~n3760;
  assign n3762 = n2437 & n2544;
  assign n3763 = n2546 & n2833;
  assign n3764 = n2434 & n2550;
  assign n3765 = n2431 & n2552;
  assign n3766 = ~n3762 & ~n3764;
  assign n3767 = ~n3765 & n3766;
  assign n3768 = ~n3763 & n3767;
  assign n3769 = n656 & n3768;
  assign n3770 = ~n656 & ~n3768;
  assign n3771 = ~n3769 & ~n3770;
  assign n3772 = ~n3761 & ~n3771;
  assign n3773 = n3761 & n3771;
  assign n3774 = ~n3772 & ~n3773;
  assign n3775 = ~n3744 & n3774;
  assign n3776 = n3744 & ~n3774;
  assign n3777 = ~n3775 & ~n3776;
  assign n3778 = ~n3743 & ~n3777;
  assign n3779 = n3743 & n3777;
  assign n3780 = ~n3778 & ~n3779;
  assign n3781 = n3733 & ~n3780;
  assign n3782 = ~n3733 & n3780;
  assign n3783 = ~n3781 & ~n3782;
  assign n3784 = n2524 & n3073;
  assign n3785 = n2426 & n3227;
  assign n3786 = n76 & ~n3159;
  assign n3787 = n2526 & n3182;
  assign n3788 = ~n3784 & ~n3786;
  assign n3789 = ~n3787 & n3788;
  assign n3790 = ~n3785 & n3789;
  assign n3791 = n57 & n3790;
  assign n3792 = ~n57 & ~n3790;
  assign n3793 = ~n3791 & ~n3792;
  assign n3794 = n3783 & n3793;
  assign n3795 = ~n3783 & ~n3793;
  assign n3796 = ~n3794 & ~n3795;
  assign n3797 = ~n3732 & n3796;
  assign n3798 = n3732 & ~n3796;
  assign n3799 = ~n3797 & ~n3798;
  assign n3800 = ~n3731 & n3799;
  assign n3801 = n3731 & ~n3799;
  assign n3802 = ~n3800 & ~n3801;
  assign n3803 = n3694 & ~n3802;
  assign n3804 = ~n3694 & n3802;
  assign n3805 = ~n3803 & ~n3804;
  assign n3806 = ~n272 & ~n434;
  assign n3807 = n1322 & n3806;
  assign n3808 = ~n156 & ~n229;
  assign n3809 = ~n334 & ~n352;
  assign n3810 = ~n480 & n3809;
  assign n3811 = n235 & n3808;
  assign n3812 = n552 & n2179;
  assign n3813 = n3811 & n3812;
  assign n3814 = n3042 & n3810;
  assign n3815 = n3807 & n3814;
  assign n3816 = n3606 & n3813;
  assign n3817 = n3815 & n3816;
  assign n3818 = n2123 & n3817;
  assign n3819 = n3602 & n3818;
  assign n3820 = ~n3805 & n3819;
  assign n3821 = n3805 & ~n3819;
  assign n3822 = ~n3820 & ~n3821;
  assign n3823 = ~n3693 & n3822;
  assign n3824 = n3693 & ~n3822;
  assign n3825 = ~n3823 & ~n3824;
  assign n3826 = pi22  & ~pi23 ;
  assign n3827 = ~pi22  & pi23 ;
  assign n3828 = ~n3826 & ~n3827;
  assign n3829 = po0  & ~n3828;
  assign n3830 = ~n3825 & n3829;
  assign n3831 = n3685 & ~n3689;
  assign n3832 = n3825 & n3831;
  assign n3833 = ~n3825 & ~n3831;
  assign n3834 = ~n3832 & ~n3833;
  assign n3835 = ~n3829 & n3834;
  assign po1  = n3830 | n3835;
  assign n3837 = ~n3821 & ~n3823;
  assign n3838 = ~n3800 & ~n3804;
  assign n3839 = n3160 & n3480;
  assign n3840 = n3212 & n3717;
  assign n3841 = ~n3717 & n3720;
  assign n3842 = ~n3480 & ~n3484;
  assign n3843 = n3717 & n3842;
  assign n3844 = ~n3841 & ~n3843;
  assign n3845 = n3169 & ~n3844;
  assign n3846 = ~n3839 & ~n3840;
  assign n3847 = ~n3845 & n3846;
  assign n3848 = n65 & ~n3847;
  assign n3849 = ~n65 & n3847;
  assign n3850 = ~n3848 & ~n3849;
  assign n3851 = ~n3794 & ~n3797;
  assign n3852 = ~n3778 & ~n3782;
  assign n3853 = n2421 & n2673;
  assign n3854 = n2668 & n3079;
  assign n3855 = ~n2515 & n2663;
  assign n3856 = n2675 & n3073;
  assign n3857 = ~n3853 & ~n3855;
  assign n3858 = ~n3856 & n3857;
  assign n3859 = ~n3854 & n3858;
  assign n3860 = n895 & ~n3859;
  assign n3861 = ~n895 & n3859;
  assign n3862 = ~n3860 & ~n3861;
  assign n3863 = ~n3761 & n3771;
  assign n3864 = ~n3744 & ~n3774;
  assign n3865 = ~n3863 & ~n3864;
  assign n3866 = ~n636 & ~n2446;
  assign n3867 = n2443 & n2638;
  assign n3868 = n2573 & n2688;
  assign n3869 = n2440 & n2566;
  assign n3870 = n2437 & n2568;
  assign n3871 = ~n3867 & ~n3869;
  assign n3872 = ~n3870 & n3871;
  assign n3873 = ~n3868 & n3872;
  assign n3874 = n3866 & ~n3873;
  assign n3875 = ~n3866 & n3873;
  assign n3876 = ~n3874 & ~n3875;
  assign n3877 = n3755 & ~n3758;
  assign n3878 = ~n636 & n2449;
  assign n3879 = n3752 & n3878;
  assign n3880 = ~n3877 & ~n3879;
  assign n3881 = ~n3876 & ~n3880;
  assign n3882 = n3876 & n3880;
  assign n3883 = ~n3881 & ~n3882;
  assign n3884 = n2431 & n2550;
  assign n3885 = n2546 & n2867;
  assign n3886 = n2434 & n2544;
  assign n3887 = n2428 & n2552;
  assign n3888 = ~n3884 & ~n3886;
  assign n3889 = ~n3887 & n3888;
  assign n3890 = ~n3885 & n3889;
  assign n3891 = n656 & n3890;
  assign n3892 = ~n656 & ~n3890;
  assign n3893 = ~n3891 & ~n3892;
  assign n3894 = ~n3883 & ~n3893;
  assign n3895 = n3883 & n3893;
  assign n3896 = ~n3894 & ~n3895;
  assign n3897 = ~n3865 & n3896;
  assign n3898 = n3865 & ~n3896;
  assign n3899 = ~n3897 & ~n3898;
  assign n3900 = ~n3862 & ~n3899;
  assign n3901 = n3862 & n3899;
  assign n3902 = ~n3900 & ~n3901;
  assign n3903 = n3852 & ~n3902;
  assign n3904 = ~n3852 & n3902;
  assign n3905 = ~n3903 & ~n3904;
  assign n3906 = n2524 & ~n3159;
  assign n3907 = n2426 & n3210;
  assign n3908 = n76 & n3182;
  assign n3909 = n2526 & ~n3204;
  assign n3910 = ~n3906 & ~n3908;
  assign n3911 = ~n3909 & n3910;
  assign n3912 = ~n3907 & n3911;
  assign n3913 = n57 & n3912;
  assign n3914 = ~n57 & ~n3912;
  assign n3915 = ~n3913 & ~n3914;
  assign n3916 = n3905 & n3915;
  assign n3917 = ~n3905 & ~n3915;
  assign n3918 = ~n3916 & ~n3917;
  assign n3919 = ~n3851 & n3918;
  assign n3920 = n3851 & ~n3918;
  assign n3921 = ~n3919 & ~n3920;
  assign n3922 = ~n3850 & n3921;
  assign n3923 = n3850 & ~n3921;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = ~n3838 & n3924;
  assign n3926 = n3838 & ~n3924;
  assign n3927 = ~n3925 & ~n3926;
  assign n3928 = ~n233 & ~n245;
  assign n3929 = ~n343 & n3928;
  assign n3930 = n1061 & n2386;
  assign n3931 = n3929 & n3930;
  assign n3932 = ~n138 & ~n217;
  assign n3933 = ~n315 & ~n320;
  assign n3934 = ~n346 & n3933;
  assign n3935 = n498 & n3932;
  assign n3936 = n568 & n3935;
  assign n3937 = n559 & n3934;
  assign n3938 = n3936 & n3937;
  assign n3939 = n3931 & n3938;
  assign n3940 = n314 & n3939;
  assign n3941 = n3663 & n3940;
  assign n3942 = n3927 & ~n3941;
  assign n3943 = ~n3927 & n3941;
  assign n3944 = ~n3942 & ~n3943;
  assign n3945 = ~n3837 & n3944;
  assign n3946 = n3837 & ~n3944;
  assign n3947 = ~n3945 & ~n3946;
  assign n3948 = ~n3832 & ~n3947;
  assign n3949 = n3832 & n3947;
  assign n3950 = ~n3948 & ~n3949;
  assign n3951 = ~po0  & ~n3834;
  assign n3952 = ~n3828 & ~n3951;
  assign n3953 = n3950 & ~n3952;
  assign n3954 = ~n3950 & n3952;
  assign po2  = n3953 | n3954;
  assign n3956 = ~n3950 & n3951;
  assign n3957 = ~n3828 & ~n3956;
  assign n3958 = ~n3942 & ~n3945;
  assign n3959 = ~n3922 & ~n3925;
  assign n3960 = ~n3916 & ~n3919;
  assign n3961 = n3169 & ~n3842;
  assign n3962 = ~n3160 & ~n3961;
  assign n3963 = n3717 & ~n3962;
  assign n3964 = n65 & n3963;
  assign n3965 = ~n65 & ~n3963;
  assign n3966 = ~n3964 & ~n3965;
  assign n3967 = ~n3900 & ~n3904;
  assign n3968 = ~n2515 & n2673;
  assign n3969 = n2668 & n3242;
  assign n3970 = n2663 & n3073;
  assign n3971 = n2675 & ~n3159;
  assign n3972 = ~n3968 & ~n3970;
  assign n3973 = ~n3971 & n3972;
  assign n3974 = ~n3969 & n3973;
  assign n3975 = n895 & ~n3974;
  assign n3976 = ~n895 & n3974;
  assign n3977 = ~n3975 & ~n3976;
  assign n3978 = ~n3883 & n3893;
  assign n3979 = ~n3865 & ~n3896;
  assign n3980 = ~n3978 & ~n3979;
  assign n3981 = ~n636 & ~n2443;
  assign n3982 = n2437 & n2566;
  assign n3983 = n2573 & n2670;
  assign n3984 = n2440 & n2638;
  assign n3985 = n2434 & n2568;
  assign n3986 = ~n3982 & ~n3984;
  assign n3987 = ~n3985 & n3986;
  assign n3988 = ~n3983 & n3987;
  assign n3989 = n3981 & ~n3988;
  assign n3990 = ~n3981 & n3988;
  assign n3991 = ~n3989 & ~n3990;
  assign n3992 = n3876 & ~n3880;
  assign n3993 = ~n636 & n2446;
  assign n3994 = n3873 & n3993;
  assign n3995 = ~n3992 & ~n3994;
  assign n3996 = ~n3991 & ~n3995;
  assign n3997 = n3991 & n3995;
  assign n3998 = ~n3996 & ~n3997;
  assign n3999 = n2431 & n2544;
  assign n4000 = n2546 & n2852;
  assign n4001 = n2428 & n2550;
  assign n4002 = n2421 & n2552;
  assign n4003 = ~n3999 & ~n4001;
  assign n4004 = ~n4002 & n4003;
  assign n4005 = ~n4000 & n4004;
  assign n4006 = n656 & n4005;
  assign n4007 = ~n656 & ~n4005;
  assign n4008 = ~n4006 & ~n4007;
  assign n4009 = ~n3998 & n4008;
  assign n4010 = n3998 & ~n4008;
  assign n4011 = ~n4009 & ~n4010;
  assign n4012 = ~n3980 & n4011;
  assign n4013 = n3980 & ~n4011;
  assign n4014 = ~n4012 & ~n4013;
  assign n4015 = ~n3977 & n4014;
  assign n4016 = n3977 & ~n4014;
  assign n4017 = ~n4015 & ~n4016;
  assign n4018 = n3967 & ~n4017;
  assign n4019 = ~n3967 & n4017;
  assign n4020 = ~n4018 & ~n4019;
  assign n4021 = n2524 & n3182;
  assign n4022 = n2426 & n3486;
  assign n4023 = n76 & ~n3204;
  assign n4024 = n2526 & n3480;
  assign n4025 = ~n4021 & ~n4023;
  assign n4026 = ~n4024 & n4025;
  assign n4027 = ~n4022 & n4026;
  assign n4028 = n57 & n4027;
  assign n4029 = ~n57 & ~n4027;
  assign n4030 = ~n4028 & ~n4029;
  assign n4031 = n4020 & n4030;
  assign n4032 = ~n4020 & ~n4030;
  assign n4033 = ~n4031 & ~n4032;
  assign n4034 = ~n3966 & n4033;
  assign n4035 = n3966 & ~n4033;
  assign n4036 = ~n4034 & ~n4035;
  assign n4037 = ~n3960 & n4036;
  assign n4038 = n3960 & ~n4036;
  assign n4039 = ~n4037 & ~n4038;
  assign n4040 = ~n3959 & n4039;
  assign n4041 = n3959 & ~n4039;
  assign n4042 = ~n4040 & ~n4041;
  assign n4043 = ~n144 & ~n286;
  assign n4044 = ~n304 & ~n317;
  assign n4045 = ~n334 & ~n360;
  assign n4046 = n4044 & n4045;
  assign n4047 = n481 & n4043;
  assign n4048 = n2179 & n4047;
  assign n4049 = n820 & n4046;
  assign n4050 = n4048 & n4049;
  assign n4051 = n210 & n453;
  assign n4052 = n3624 & n4051;
  assign n4053 = n2030 & n4050;
  assign n4054 = n4052 & n4053;
  assign n4055 = n1333 & n4054;
  assign n4056 = n4042 & ~n4055;
  assign n4057 = ~n4042 & n4055;
  assign n4058 = ~n4056 & ~n4057;
  assign n4059 = ~n3958 & n4058;
  assign n4060 = n3958 & ~n4058;
  assign n4061 = ~n4059 & ~n4060;
  assign n4062 = n3949 & n4061;
  assign n4063 = ~n3949 & ~n4061;
  assign n4064 = ~n4062 & ~n4063;
  assign n4065 = n3957 & n4064;
  assign n4066 = ~n3957 & ~n4064;
  assign po3  = ~n4065 & ~n4066;
  assign n4068 = ~n4056 & ~n4059;
  assign n4069 = ~n4037 & ~n4040;
  assign n4070 = ~n4031 & ~n4034;
  assign n4071 = ~n4015 & ~n4019;
  assign n4072 = ~n4009 & ~n4012;
  assign n4073 = n2437 & n2638;
  assign n4074 = n2573 & n2833;
  assign n4075 = n2434 & n2566;
  assign n4076 = n2431 & n2568;
  assign n4077 = ~n4073 & ~n4075;
  assign n4078 = ~n4076 & n4077;
  assign n4079 = ~n4074 & n4078;
  assign n4080 = n636 & ~n4079;
  assign n4081 = ~n636 & n4079;
  assign n4082 = ~n4080 & ~n4081;
  assign n4083 = ~n636 & n2440;
  assign n4084 = ~n65 & n4083;
  assign n4085 = n65 & ~n4083;
  assign n4086 = ~n4084 & ~n4085;
  assign n4087 = ~n4082 & n4086;
  assign n4088 = n4082 & ~n4086;
  assign n4089 = ~n4087 & ~n4088;
  assign n4090 = n3991 & ~n3995;
  assign n4091 = ~n636 & n2443;
  assign n4092 = n3988 & n4091;
  assign n4093 = ~n4090 & ~n4092;
  assign n4094 = ~n4089 & ~n4093;
  assign n4095 = n4089 & n4093;
  assign n4096 = ~n4094 & ~n4095;
  assign n4097 = n2421 & n2550;
  assign n4098 = n2521 & n2546;
  assign n4099 = n2428 & n2544;
  assign n4100 = ~n2515 & n2552;
  assign n4101 = ~n4097 & ~n4099;
  assign n4102 = ~n4100 & n4101;
  assign n4103 = ~n4098 & n4102;
  assign n4104 = ~n656 & ~n4103;
  assign n4105 = n656 & n4103;
  assign n4106 = ~n4104 & ~n4105;
  assign n4107 = ~n4096 & ~n4106;
  assign n4108 = n4096 & n4106;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = ~n4072 & n4109;
  assign n4111 = n4072 & ~n4109;
  assign n4112 = ~n4110 & ~n4111;
  assign n4113 = n2673 & n3073;
  assign n4114 = n2668 & n3227;
  assign n4115 = n2663 & ~n3159;
  assign n4116 = n2675 & n3182;
  assign n4117 = ~n4113 & ~n4115;
  assign n4118 = ~n4116 & n4117;
  assign n4119 = ~n4114 & n4118;
  assign n4120 = ~n895 & n4119;
  assign n4121 = n895 & ~n4119;
  assign n4122 = ~n4120 & ~n4121;
  assign n4123 = ~n4112 & ~n4122;
  assign n4124 = n4112 & n4122;
  assign n4125 = ~n4123 & ~n4124;
  assign n4126 = ~n4071 & n4125;
  assign n4127 = n4071 & ~n4125;
  assign n4128 = ~n4126 & ~n4127;
  assign n4129 = n2524 & ~n3204;
  assign n4130 = n2426 & n3722;
  assign n4131 = n76 & n3480;
  assign n4132 = n2526 & n3717;
  assign n4133 = ~n4129 & ~n4131;
  assign n4134 = ~n4132 & n4133;
  assign n4135 = ~n4130 & n4134;
  assign n4136 = ~n57 & ~n4135;
  assign n4137 = n57 & n4135;
  assign n4138 = ~n4136 & ~n4137;
  assign n4139 = n4128 & n4138;
  assign n4140 = ~n4128 & ~n4138;
  assign n4141 = ~n4139 & ~n4140;
  assign n4142 = ~n4070 & n4141;
  assign n4143 = n4070 & ~n4141;
  assign n4144 = ~n4142 & ~n4143;
  assign n4145 = n4069 & ~n4144;
  assign n4146 = ~n4069 & n4144;
  assign n4147 = ~n4145 & ~n4146;
  assign n4148 = ~n300 & ~n319;
  assign n4149 = ~n353 & n4148;
  assign n4150 = n318 & n549;
  assign n4151 = n658 & n2271;
  assign n4152 = n2386 & n4151;
  assign n4153 = n4149 & n4150;
  assign n4154 = n4152 & n4153;
  assign n4155 = n847 & n4154;
  assign n4156 = n192 & n4155;
  assign n4157 = n2313 & n4156;
  assign n4158 = ~n4147 & n4157;
  assign n4159 = n4147 & ~n4157;
  assign n4160 = ~n4158 & ~n4159;
  assign n4161 = ~n4068 & n4160;
  assign n4162 = n4068 & ~n4160;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = ~n4062 & ~n4163;
  assign n4165 = n4062 & n4163;
  assign n4166 = ~n4164 & ~n4165;
  assign n4167 = n3956 & ~n4064;
  assign n4168 = ~n3828 & ~n4167;
  assign n4169 = n4166 & ~n4168;
  assign n4170 = ~n4166 & n4168;
  assign po4  = n4169 | n4170;
  assign n4172 = ~n4159 & ~n4161;
  assign n4173 = ~n4142 & ~n4146;
  assign n4174 = ~n4126 & ~n4139;
  assign n4175 = n2524 & n3480;
  assign n4176 = n76 & n3717;
  assign n4177 = n2426 & ~n3844;
  assign n4178 = ~n4175 & ~n4176;
  assign n4179 = ~n4177 & n4178;
  assign n4180 = ~n57 & ~n4179;
  assign n4181 = n57 & n4179;
  assign n4182 = ~n4180 & ~n4181;
  assign n4183 = ~n4072 & ~n4109;
  assign n4184 = ~n4123 & ~n4183;
  assign n4185 = n2673 & ~n3159;
  assign n4186 = n2668 & n3210;
  assign n4187 = n2663 & n3182;
  assign n4188 = n2675 & ~n3204;
  assign n4189 = ~n4185 & ~n4187;
  assign n4190 = ~n4188 & n4189;
  assign n4191 = ~n4186 & n4190;
  assign n4192 = n895 & ~n4191;
  assign n4193 = ~n895 & n4191;
  assign n4194 = ~n4192 & ~n4193;
  assign n4195 = ~n4096 & n4106;
  assign n4196 = n4089 & ~n4093;
  assign n4197 = ~n4195 & ~n4196;
  assign n4198 = n2421 & n2544;
  assign n4199 = n2546 & n3079;
  assign n4200 = ~n2515 & n2550;
  assign n4201 = n2552 & n3073;
  assign n4202 = ~n4198 & ~n4200;
  assign n4203 = ~n4201 & n4202;
  assign n4204 = ~n4199 & n4203;
  assign n4205 = ~n656 & ~n4204;
  assign n4206 = n656 & n4204;
  assign n4207 = ~n4205 & ~n4206;
  assign n4208 = n2431 & n2566;
  assign n4209 = n2573 & n2867;
  assign n4210 = n2434 & n2638;
  assign n4211 = n2428 & n2568;
  assign n4212 = ~n4208 & ~n4210;
  assign n4213 = ~n4211 & n4212;
  assign n4214 = ~n4209 & n4213;
  assign n4215 = n636 & n4214;
  assign n4216 = ~n636 & ~n4214;
  assign n4217 = ~n4215 & ~n4216;
  assign n4218 = ~n4084 & ~n4087;
  assign n4219 = ~n636 & n2437;
  assign n4220 = ~n65 & n4219;
  assign n4221 = n65 & ~n4219;
  assign n4222 = ~n4220 & ~n4221;
  assign n4223 = ~n4218 & n4222;
  assign n4224 = n4218 & ~n4222;
  assign n4225 = ~n4223 & ~n4224;
  assign n4226 = n4217 & n4225;
  assign n4227 = ~n4217 & ~n4225;
  assign n4228 = ~n4226 & ~n4227;
  assign n4229 = n4207 & n4228;
  assign n4230 = ~n4207 & ~n4228;
  assign n4231 = ~n4229 & ~n4230;
  assign n4232 = ~n4197 & n4231;
  assign n4233 = n4197 & ~n4231;
  assign n4234 = ~n4232 & ~n4233;
  assign n4235 = ~n4194 & n4234;
  assign n4236 = n4194 & ~n4234;
  assign n4237 = ~n4235 & ~n4236;
  assign n4238 = ~n4184 & n4237;
  assign n4239 = n4184 & ~n4237;
  assign n4240 = ~n4238 & ~n4239;
  assign n4241 = n4182 & n4240;
  assign n4242 = ~n4182 & ~n4240;
  assign n4243 = ~n4241 & ~n4242;
  assign n4244 = ~n4174 & n4243;
  assign n4245 = n4174 & ~n4243;
  assign n4246 = ~n4244 & ~n4245;
  assign n4247 = ~n4173 & n4246;
  assign n4248 = n4173 & ~n4246;
  assign n4249 = ~n4247 & ~n4248;
  assign n4250 = ~n360 & n2269;
  assign n4251 = n508 & n2142;
  assign n4252 = ~n228 & ~n296;
  assign n4253 = ~n300 & ~n332;
  assign n4254 = n4252 & n4253;
  assign n4255 = n335 & n476;
  assign n4256 = n4254 & n4255;
  assign n4257 = n3807 & n4250;
  assign n4258 = n4251 & n4257;
  assign n4259 = n2154 & n4256;
  assign n4260 = n4258 & n4259;
  assign n4261 = n3057 & n4260;
  assign n4262 = n3702 & n4261;
  assign n4263 = ~n4249 & n4262;
  assign n4264 = n4249 & ~n4262;
  assign n4265 = ~n4263 & ~n4264;
  assign n4266 = ~n4172 & n4265;
  assign n4267 = n4172 & ~n4265;
  assign n4268 = ~n4266 & ~n4267;
  assign n4269 = ~n4165 & ~n4268;
  assign n4270 = n4165 & n4268;
  assign n4271 = ~n4269 & ~n4270;
  assign n4272 = ~n4166 & n4167;
  assign n4273 = ~n3828 & ~n4272;
  assign n4274 = n4271 & ~n4273;
  assign n4275 = ~n4271 & n4273;
  assign po5  = n4274 | n4275;
  assign n4277 = ~n4264 & ~n4266;
  assign n4278 = ~n4244 & ~n4247;
  assign n4279 = ~n4238 & ~n4241;
  assign n4280 = ~n4232 & ~n4235;
  assign n4281 = n2426 & ~n3842;
  assign n4282 = ~n2524 & ~n4281;
  assign n4283 = n3717 & ~n4282;
  assign n4284 = n57 & n4283;
  assign n4285 = ~n57 & ~n4283;
  assign n4286 = ~n4284 & ~n4285;
  assign n4287 = ~n4280 & ~n4286;
  assign n4288 = n4280 & n4286;
  assign n4289 = ~n4287 & ~n4288;
  assign n4290 = n2673 & n3182;
  assign n4291 = n2668 & n3486;
  assign n4292 = n2663 & ~n3204;
  assign n4293 = n2675 & n3480;
  assign n4294 = ~n4290 & ~n4292;
  assign n4295 = ~n4293 & n4294;
  assign n4296 = ~n4291 & n4295;
  assign n4297 = n895 & ~n4296;
  assign n4298 = ~n895 & n4296;
  assign n4299 = ~n4297 & ~n4298;
  assign n4300 = ~n4226 & ~n4229;
  assign n4301 = ~n2515 & n2544;
  assign n4302 = n2546 & n3242;
  assign n4303 = n2550 & n3073;
  assign n4304 = n2552 & ~n3159;
  assign n4305 = ~n4301 & ~n4303;
  assign n4306 = ~n4304 & n4305;
  assign n4307 = ~n4302 & n4306;
  assign n4308 = ~n656 & ~n4307;
  assign n4309 = n656 & n4307;
  assign n4310 = ~n4308 & ~n4309;
  assign n4311 = n2431 & n2638;
  assign n4312 = n2573 & n2852;
  assign n4313 = n2428 & n2566;
  assign n4314 = n2421 & n2568;
  assign n4315 = ~n4311 & ~n4313;
  assign n4316 = ~n4314 & n4315;
  assign n4317 = ~n4312 & n4316;
  assign n4318 = n636 & n4317;
  assign n4319 = ~n636 & ~n4317;
  assign n4320 = ~n4318 & ~n4319;
  assign n4321 = ~n4220 & ~n4223;
  assign n4322 = ~n636 & n2434;
  assign n4323 = ~n65 & n4322;
  assign n4324 = n65 & ~n4322;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = ~n4321 & n4325;
  assign n4327 = n4321 & ~n4325;
  assign n4328 = ~n4326 & ~n4327;
  assign n4329 = n4320 & n4328;
  assign n4330 = ~n4320 & ~n4328;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = n4310 & n4331;
  assign n4333 = ~n4310 & ~n4331;
  assign n4334 = ~n4332 & ~n4333;
  assign n4335 = ~n4300 & n4334;
  assign n4336 = n4300 & ~n4334;
  assign n4337 = ~n4335 & ~n4336;
  assign n4338 = ~n4299 & n4337;
  assign n4339 = n4299 & ~n4337;
  assign n4340 = ~n4338 & ~n4339;
  assign n4341 = n4289 & n4340;
  assign n4342 = ~n4289 & ~n4340;
  assign n4343 = ~n4341 & ~n4342;
  assign n4344 = ~n4279 & n4343;
  assign n4345 = n4279 & ~n4343;
  assign n4346 = ~n4344 & ~n4345;
  assign n4347 = ~n4278 & n4346;
  assign n4348 = n4278 & ~n4346;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = ~n347 & n436;
  assign n4351 = n797 & n856;
  assign n4352 = n1005 & n2142;
  assign n4353 = n2179 & n4352;
  assign n4354 = n4350 & n4351;
  assign n4355 = n461 & n4354;
  assign n4356 = n2274 & n4353;
  assign n4357 = n4355 & n4356;
  assign n4358 = ~n152 & ~n241;
  assign n4359 = ~n290 & ~n348;
  assign n4360 = n4358 & n4359;
  assign n4361 = n843 & n2143;
  assign n4362 = n3170 & n4361;
  assign n4363 = n4360 & n4362;
  assign n4364 = n2307 & n4363;
  assign n4365 = n4357 & n4364;
  assign n4366 = n3605 & n4365;
  assign n4367 = ~n4349 & n4366;
  assign n4368 = n4349 & ~n4366;
  assign n4369 = ~n4367 & ~n4368;
  assign n4370 = ~n4277 & n4369;
  assign n4371 = n4277 & ~n4369;
  assign n4372 = ~n4370 & ~n4371;
  assign n4373 = ~n4270 & ~n4372;
  assign n4374 = n4270 & n4372;
  assign n4375 = ~n4373 & ~n4374;
  assign n4376 = ~n4271 & n4272;
  assign n4377 = ~n3828 & ~n4376;
  assign n4378 = n4375 & ~n4377;
  assign n4379 = ~n4375 & n4377;
  assign po6  = n4378 | n4379;
  assign n4381 = ~n4368 & ~n4370;
  assign n4382 = ~n4344 & ~n4347;
  assign n4383 = ~n4287 & ~n4341;
  assign n4384 = ~n4335 & ~n4338;
  assign n4385 = n2673 & ~n3204;
  assign n4386 = n2668 & n3722;
  assign n4387 = n2663 & n3480;
  assign n4388 = n2675 & n3717;
  assign n4389 = ~n4385 & ~n4387;
  assign n4390 = ~n4388 & n4389;
  assign n4391 = ~n4386 & n4390;
  assign n4392 = n895 & n4391;
  assign n4393 = ~n895 & ~n4391;
  assign n4394 = ~n4392 & ~n4393;
  assign n4395 = ~n4384 & n4394;
  assign n4396 = n4384 & ~n4394;
  assign n4397 = ~n4395 & ~n4396;
  assign n4398 = ~n4329 & ~n4332;
  assign n4399 = n2544 & n3073;
  assign n4400 = n2546 & n3227;
  assign n4401 = n2550 & ~n3159;
  assign n4402 = n2552 & n3182;
  assign n4403 = ~n4399 & ~n4401;
  assign n4404 = ~n4402 & n4403;
  assign n4405 = ~n4400 & n4404;
  assign n4406 = n656 & n4405;
  assign n4407 = ~n656 & ~n4405;
  assign n4408 = ~n4406 & ~n4407;
  assign n4409 = ~n4323 & ~n4326;
  assign n4410 = n2421 & n2566;
  assign n4411 = n2521 & n2573;
  assign n4412 = n2428 & n2638;
  assign n4413 = ~n2515 & n2568;
  assign n4414 = ~n4410 & ~n4412;
  assign n4415 = ~n4413 & n4414;
  assign n4416 = ~n4411 & n4415;
  assign n4417 = n636 & ~n4416;
  assign n4418 = ~n636 & n4416;
  assign n4419 = ~n4417 & ~n4418;
  assign n4420 = ~n636 & n2431;
  assign n4421 = n57 & n65;
  assign n4422 = ~n57 & ~n65;
  assign n4423 = ~n4421 & ~n4422;
  assign n4424 = n4420 & n4423;
  assign n4425 = ~n4420 & ~n4423;
  assign n4426 = ~n4424 & ~n4425;
  assign n4427 = ~n4419 & ~n4426;
  assign n4428 = n4419 & n4426;
  assign n4429 = ~n4427 & ~n4428;
  assign n4430 = ~n4409 & ~n4429;
  assign n4431 = n4409 & n4429;
  assign n4432 = ~n4430 & ~n4431;
  assign n4433 = n4408 & n4432;
  assign n4434 = ~n4408 & ~n4432;
  assign n4435 = ~n4433 & ~n4434;
  assign n4436 = ~n4398 & n4435;
  assign n4437 = n4398 & ~n4435;
  assign n4438 = ~n4436 & ~n4437;
  assign n4439 = n4397 & n4438;
  assign n4440 = ~n4397 & ~n4438;
  assign n4441 = ~n4439 & ~n4440;
  assign n4442 = ~n4383 & n4441;
  assign n4443 = n4383 & ~n4441;
  assign n4444 = ~n4442 & ~n4443;
  assign n4445 = n4382 & ~n4444;
  assign n4446 = ~n4382 & n4444;
  assign n4447 = ~n4445 & ~n4446;
  assign n4448 = ~n240 & ~n353;
  assign n4449 = ~n212 & ~n220;
  assign n4450 = ~n229 & ~n343;
  assign n4451 = n4449 & n4450;
  assign n4452 = n321 & n782;
  assign n4453 = n985 & n4448;
  assign n4454 = n4452 & n4453;
  assign n4455 = n4250 & n4451;
  assign n4456 = n4454 & n4455;
  assign n4457 = n4357 & n4456;
  assign n4458 = n2126 & n4457;
  assign n4459 = n4447 & ~n4458;
  assign n4460 = ~n4447 & n4458;
  assign n4461 = ~n4459 & ~n4460;
  assign n4462 = ~n4381 & n4461;
  assign n4463 = n4381 & ~n4461;
  assign n4464 = ~n4462 & ~n4463;
  assign n4465 = n4374 & n4464;
  assign n4466 = ~n4374 & ~n4464;
  assign n4467 = ~n4465 & ~n4466;
  assign n4468 = ~n4375 & n4376;
  assign n4469 = ~n3828 & ~n4468;
  assign n4470 = n4467 & ~n4469;
  assign n4471 = ~n4467 & n4469;
  assign po7  = n4470 | n4471;
  assign n4473 = ~n4459 & ~n4462;
  assign n4474 = ~n4442 & ~n4446;
  assign n4475 = ~n4395 & ~n4439;
  assign n4476 = n2673 & n3480;
  assign n4477 = n2663 & n3717;
  assign n4478 = n2668 & ~n3844;
  assign n4479 = ~n4476 & ~n4477;
  assign n4480 = ~n4478 & n4479;
  assign n4481 = n895 & ~n4480;
  assign n4482 = ~n895 & n4480;
  assign n4483 = ~n4481 & ~n4482;
  assign n4484 = ~n4433 & ~n4436;
  assign n4485 = n2544 & ~n3159;
  assign n4486 = n2546 & n3210;
  assign n4487 = n2550 & n3182;
  assign n4488 = n2552 & ~n3204;
  assign n4489 = ~n4485 & ~n4487;
  assign n4490 = ~n4488 & n4489;
  assign n4491 = ~n4486 & n4490;
  assign n4492 = ~n656 & ~n4491;
  assign n4493 = n656 & n4491;
  assign n4494 = ~n4492 & ~n4493;
  assign n4495 = ~n4419 & n4426;
  assign n4496 = ~n4430 & ~n4495;
  assign n4497 = ~n636 & n2428;
  assign n4498 = ~n4421 & ~n4424;
  assign n4499 = ~n4497 & n4498;
  assign n4500 = n4497 & ~n4498;
  assign n4501 = ~n4499 & ~n4500;
  assign n4502 = n2421 & n2638;
  assign n4503 = n2573 & n3079;
  assign n4504 = ~n2515 & n2566;
  assign n4505 = n2568 & n3073;
  assign n4506 = ~n4502 & ~n4504;
  assign n4507 = ~n4505 & n4506;
  assign n4508 = ~n4503 & n4507;
  assign n4509 = n636 & n4508;
  assign n4510 = ~n636 & ~n4508;
  assign n4511 = ~n4509 & ~n4510;
  assign n4512 = ~n4501 & n4511;
  assign n4513 = n4501 & ~n4511;
  assign n4514 = ~n4512 & ~n4513;
  assign n4515 = ~n4496 & n4514;
  assign n4516 = n4496 & ~n4514;
  assign n4517 = ~n4515 & ~n4516;
  assign n4518 = n4494 & n4517;
  assign n4519 = ~n4494 & ~n4517;
  assign n4520 = ~n4518 & ~n4519;
  assign n4521 = ~n4484 & n4520;
  assign n4522 = n4484 & ~n4520;
  assign n4523 = ~n4521 & ~n4522;
  assign n4524 = ~n4483 & n4523;
  assign n4525 = n4483 & ~n4523;
  assign n4526 = ~n4524 & ~n4525;
  assign n4527 = ~n4475 & n4526;
  assign n4528 = n4475 & ~n4526;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = ~n4474 & n4529;
  assign n4531 = n4474 & ~n4529;
  assign n4532 = ~n4530 & ~n4531;
  assign n4533 = ~n167 & ~n199;
  assign n4534 = ~n253 & n4533;
  assign n4535 = n361 & n610;
  assign n4536 = n2076 & n4535;
  assign n4537 = n4534 & n4536;
  assign n4538 = n2015 & n4537;
  assign n4539 = n446 & n4538;
  assign n4540 = ~n227 & ~n232;
  assign n4541 = ~n479 & ~n546;
  assign n4542 = ~n616 & n4541;
  assign n4543 = n2174 & n4540;
  assign n4544 = n4542 & n4543;
  assign n4545 = n850 & n2184;
  assign n4546 = n4544 & n4545;
  assign n4547 = n859 & n4546;
  assign n4548 = n3642 & n4547;
  assign n4549 = n4539 & n4548;
  assign n4550 = ~n4532 & n4549;
  assign n4551 = n4532 & ~n4549;
  assign n4552 = ~n4550 & ~n4551;
  assign n4553 = ~n4473 & n4552;
  assign n4554 = n4473 & ~n4552;
  assign n4555 = ~n4553 & ~n4554;
  assign n4556 = ~n4465 & ~n4555;
  assign n4557 = n4465 & n4555;
  assign n4558 = ~n4556 & ~n4557;
  assign n4559 = ~n4467 & n4468;
  assign n4560 = ~n3828 & ~n4559;
  assign n4561 = n4558 & ~n4560;
  assign n4562 = ~n4558 & n4560;
  assign po8  = n4561 | n4562;
  assign n4564 = ~n4551 & ~n4553;
  assign n4565 = ~n4527 & ~n4530;
  assign n4566 = ~n4521 & ~n4524;
  assign n4567 = ~n4515 & ~n4518;
  assign n4568 = n2668 & ~n3842;
  assign n4569 = ~n2673 & ~n4568;
  assign n4570 = n3717 & ~n4569;
  assign n4571 = ~n895 & ~n4570;
  assign n4572 = n895 & n4570;
  assign n4573 = ~n4571 & ~n4572;
  assign n4574 = ~n4567 & ~n4573;
  assign n4575 = n4567 & n4573;
  assign n4576 = ~n4574 & ~n4575;
  assign n4577 = n2544 & n3182;
  assign n4578 = n2546 & n3486;
  assign n4579 = n2550 & ~n3204;
  assign n4580 = n2552 & n3480;
  assign n4581 = ~n4577 & ~n4579;
  assign n4582 = ~n4580 & n4581;
  assign n4583 = ~n4578 & n4582;
  assign n4584 = ~n656 & ~n4583;
  assign n4585 = n656 & n4583;
  assign n4586 = ~n4584 & ~n4585;
  assign n4587 = ~n4497 & ~n4498;
  assign n4588 = ~n4512 & ~n4587;
  assign n4589 = ~n2515 & n2638;
  assign n4590 = n2573 & n3242;
  assign n4591 = n2566 & n3073;
  assign n4592 = n2568 & ~n3159;
  assign n4593 = ~n4589 & ~n4591;
  assign n4594 = ~n4592 & n4593;
  assign n4595 = ~n4590 & n4594;
  assign n4596 = n636 & ~n4595;
  assign n4597 = ~n636 & n4595;
  assign n4598 = ~n4596 & ~n4597;
  assign n4599 = ~n636 & n2493;
  assign n4600 = ~n4598 & ~n4599;
  assign n4601 = n4598 & n4599;
  assign n4602 = ~n4600 & ~n4601;
  assign n4603 = ~n4588 & n4602;
  assign n4604 = n4588 & ~n4602;
  assign n4605 = ~n4603 & ~n4604;
  assign n4606 = n4586 & n4605;
  assign n4607 = ~n4586 & ~n4605;
  assign n4608 = ~n4606 & ~n4607;
  assign n4609 = n4576 & n4608;
  assign n4610 = ~n4576 & ~n4608;
  assign n4611 = ~n4609 & ~n4610;
  assign n4612 = ~n4566 & n4611;
  assign n4613 = n4566 & ~n4611;
  assign n4614 = ~n4612 & ~n4613;
  assign n4615 = n4565 & ~n4614;
  assign n4616 = ~n4565 & n4614;
  assign n4617 = ~n4615 & ~n4616;
  assign n4618 = ~n165 & ~n179;
  assign n4619 = ~n267 & ~n297;
  assign n4620 = ~n358 & ~n392;
  assign n4621 = ~n480 & n4620;
  assign n4622 = n4618 & n4619;
  assign n4623 = n321 & n3170;
  assign n4624 = n4622 & n4623;
  assign n4625 = n3042 & n4621;
  assign n4626 = n4624 & n4625;
  assign n4627 = n251 & n4626;
  assign n4628 = n3588 & n4627;
  assign n4629 = n2283 & n4628;
  assign n4630 = ~n4617 & n4629;
  assign n4631 = n4617 & ~n4629;
  assign n4632 = ~n4630 & ~n4631;
  assign n4633 = ~n4564 & n4632;
  assign n4634 = n4564 & ~n4632;
  assign n4635 = ~n4633 & ~n4634;
  assign n4636 = ~n4557 & ~n4635;
  assign n4637 = n4557 & n4635;
  assign n4638 = ~n4636 & ~n4637;
  assign n4639 = ~n4558 & n4559;
  assign n4640 = ~n3828 & ~n4639;
  assign n4641 = n4638 & ~n4640;
  assign n4642 = ~n4638 & n4640;
  assign po9  = n4641 | n4642;
  assign n4644 = ~n4631 & ~n4633;
  assign n4645 = ~n4612 & ~n4616;
  assign n4646 = ~n4574 & ~n4609;
  assign n4647 = ~n4603 & ~n4606;
  assign n4648 = n2544 & ~n3204;
  assign n4649 = n2546 & n3722;
  assign n4650 = n2550 & n3480;
  assign n4651 = n2552 & n3717;
  assign n4652 = ~n4648 & ~n4650;
  assign n4653 = ~n4651 & n4652;
  assign n4654 = ~n4649 & n4653;
  assign n4655 = n656 & n4654;
  assign n4656 = ~n656 & ~n4654;
  assign n4657 = ~n4655 & ~n4656;
  assign n4658 = ~n4647 & n4657;
  assign n4659 = n4647 & ~n4657;
  assign n4660 = ~n4658 & ~n4659;
  assign n4661 = n2638 & n3073;
  assign n4662 = n2573 & n3227;
  assign n4663 = n2566 & ~n3159;
  assign n4664 = n2568 & n3182;
  assign n4665 = ~n4661 & ~n4663;
  assign n4666 = ~n4664 & n4665;
  assign n4667 = ~n4662 & n4666;
  assign n4668 = ~n636 & n4667;
  assign n4669 = n636 & ~n4667;
  assign n4670 = ~n4668 & ~n4669;
  assign n4671 = ~n636 & ~n2515;
  assign n4672 = n895 & n4671;
  assign n4673 = ~n895 & ~n4671;
  assign n4674 = ~n4672 & ~n4673;
  assign n4675 = n4497 & ~n4674;
  assign n4676 = ~n4497 & n4674;
  assign n4677 = ~n4675 & ~n4676;
  assign n4678 = ~n636 & ~n2428;
  assign n4679 = n2421 & n4678;
  assign n4680 = ~n4600 & ~n4679;
  assign n4681 = ~n4677 & ~n4680;
  assign n4682 = n4677 & n4680;
  assign n4683 = ~n4681 & ~n4682;
  assign n4684 = n4670 & ~n4683;
  assign n4685 = ~n4670 & n4683;
  assign n4686 = ~n4684 & ~n4685;
  assign n4687 = n4660 & n4686;
  assign n4688 = ~n4660 & ~n4686;
  assign n4689 = ~n4687 & ~n4688;
  assign n4690 = ~n4646 & n4689;
  assign n4691 = n4646 & ~n4689;
  assign n4692 = ~n4690 & ~n4691;
  assign n4693 = ~n4645 & n4692;
  assign n4694 = n4645 & ~n4692;
  assign n4695 = ~n4693 & ~n4694;
  assign n4696 = ~n218 & ~n450;
  assign n4697 = ~n492 & n4696;
  assign n4698 = n345 & n2390;
  assign n4699 = n3170 & n4698;
  assign n4700 = n160 & n4697;
  assign n4701 = n857 & n3039;
  assign n4702 = n4700 & n4701;
  assign n4703 = n4699 & n4702;
  assign n4704 = n545 & n4703;
  assign n4705 = n996 & n3631;
  assign n4706 = n4704 & n4705;
  assign n4707 = ~n4695 & n4706;
  assign n4708 = n4695 & ~n4706;
  assign n4709 = ~n4707 & ~n4708;
  assign n4710 = ~n4644 & n4709;
  assign n4711 = n4644 & ~n4709;
  assign n4712 = ~n4710 & ~n4711;
  assign n4713 = ~n4637 & ~n4712;
  assign n4714 = n4637 & n4712;
  assign n4715 = ~n4713 & ~n4714;
  assign n4716 = ~n4638 & n4639;
  assign n4717 = ~n3828 & ~n4716;
  assign n4718 = n4715 & ~n4717;
  assign n4719 = ~n4715 & n4717;
  assign po10  = n4718 | n4719;
  assign n4721 = ~n4708 & ~n4710;
  assign n4722 = ~n4690 & ~n4693;
  assign n4723 = ~n4658 & ~n4687;
  assign n4724 = n2544 & n3480;
  assign n4725 = n2550 & n3717;
  assign n4726 = n2546 & ~n3844;
  assign n4727 = ~n4724 & ~n4725;
  assign n4728 = ~n4726 & n4727;
  assign n4729 = ~n656 & ~n4728;
  assign n4730 = n656 & n4728;
  assign n4731 = ~n4729 & ~n4730;
  assign n4732 = n2638 & ~n3159;
  assign n4733 = n2573 & n3210;
  assign n4734 = n2566 & n3182;
  assign n4735 = n2568 & ~n3204;
  assign n4736 = ~n4732 & ~n4734;
  assign n4737 = ~n4735 & n4736;
  assign n4738 = ~n4733 & n4737;
  assign n4739 = n636 & n4738;
  assign n4740 = ~n636 & ~n4738;
  assign n4741 = ~n4739 & ~n4740;
  assign n4742 = ~n636 & n3073;
  assign n4743 = ~n4497 & ~n4672;
  assign n4744 = ~n4673 & ~n4743;
  assign n4745 = ~n4742 & n4744;
  assign n4746 = n4742 & ~n4744;
  assign n4747 = ~n4745 & ~n4746;
  assign n4748 = n4741 & n4747;
  assign n4749 = ~n4741 & ~n4747;
  assign n4750 = ~n4748 & ~n4749;
  assign n4751 = n4670 & ~n4681;
  assign n4752 = ~n4682 & ~n4751;
  assign n4753 = n4750 & n4752;
  assign n4754 = ~n4750 & ~n4752;
  assign n4755 = ~n4753 & ~n4754;
  assign n4756 = n4731 & n4755;
  assign n4757 = ~n4731 & ~n4755;
  assign n4758 = ~n4756 & ~n4757;
  assign n4759 = ~n4723 & n4758;
  assign n4760 = n4723 & ~n4758;
  assign n4761 = ~n4759 & ~n4760;
  assign n4762 = ~n4722 & n4761;
  assign n4763 = n4722 & ~n4761;
  assign n4764 = ~n4762 & ~n4763;
  assign n4765 = ~n339 & n805;
  assign n4766 = n842 & n4765;
  assign n4767 = n615 & n4766;
  assign n4768 = n661 & n4767;
  assign n4769 = n3466 & n4768;
  assign n4770 = n582 & n4769;
  assign n4771 = ~n4764 & n4770;
  assign n4772 = n4764 & ~n4770;
  assign n4773 = ~n4771 & ~n4772;
  assign n4774 = ~n4721 & n4773;
  assign n4775 = n4721 & ~n4773;
  assign n4776 = ~n4774 & ~n4775;
  assign n4777 = ~n4714 & ~n4776;
  assign n4778 = n4714 & n4776;
  assign n4779 = ~n4777 & ~n4778;
  assign n4780 = ~n4715 & n4716;
  assign n4781 = ~n3828 & ~n4780;
  assign n4782 = n4779 & ~n4781;
  assign n4783 = ~n4779 & n4781;
  assign po11  = n4782 | n4783;
  assign n4785 = ~n4772 & ~n4774;
  assign n4786 = ~n4759 & ~n4762;
  assign n4787 = ~n4753 & ~n4756;
  assign n4788 = ~n4745 & ~n4748;
  assign n4789 = ~n636 & ~n3159;
  assign n4790 = ~n3073 & n4789;
  assign n4791 = n3159 & n4742;
  assign n4792 = ~n4790 & ~n4791;
  assign n4793 = ~n4788 & n4792;
  assign n4794 = n4788 & ~n4792;
  assign n4795 = ~n4793 & ~n4794;
  assign n4796 = n2638 & n3182;
  assign n4797 = n2573 & n3486;
  assign n4798 = n2566 & ~n3204;
  assign n4799 = n2568 & n3480;
  assign n4800 = ~n4796 & ~n4798;
  assign n4801 = ~n4799 & n4800;
  assign n4802 = ~n4797 & n4801;
  assign n4803 = ~n636 & n4802;
  assign n4804 = n636 & ~n4802;
  assign n4805 = ~n4803 & ~n4804;
  assign n4806 = n2546 & ~n3842;
  assign n4807 = ~n2544 & ~n4806;
  assign n4808 = n3717 & ~n4807;
  assign n4809 = n656 & n4808;
  assign n4810 = ~n656 & ~n4808;
  assign n4811 = ~n4809 & ~n4810;
  assign n4812 = ~n4805 & ~n4811;
  assign n4813 = n4805 & n4811;
  assign n4814 = ~n4812 & ~n4813;
  assign n4815 = n4795 & n4814;
  assign n4816 = ~n4795 & ~n4814;
  assign n4817 = ~n4815 & ~n4816;
  assign n4818 = ~n4787 & n4817;
  assign n4819 = n4787 & ~n4817;
  assign n4820 = ~n4818 & ~n4819;
  assign n4821 = ~n4786 & n4820;
  assign n4822 = n4786 & ~n4820;
  assign n4823 = ~n4821 & ~n4822;
  assign n4824 = ~n254 & ~n291;
  assign n4825 = ~n392 & ~n479;
  assign n4826 = ~n657 & n4825;
  assign n4827 = n4824 & n4826;
  assign n4828 = ~n149 & ~n253;
  assign n4829 = n2201 & n4828;
  assign n4830 = n820 & n4829;
  assign n4831 = n3931 & n4830;
  assign n4832 = n4827 & n4831;
  assign n4833 = n2100 & n4832;
  assign n4834 = n2220 & n4833;
  assign n4835 = ~n4823 & n4834;
  assign n4836 = n4823 & ~n4834;
  assign n4837 = ~n4835 & ~n4836;
  assign n4838 = ~n4785 & n4837;
  assign n4839 = n4785 & ~n4837;
  assign n4840 = ~n4838 & ~n4839;
  assign n4841 = ~n4778 & ~n4840;
  assign n4842 = n4778 & n4840;
  assign n4843 = ~n4841 & ~n4842;
  assign n4844 = ~n4779 & n4780;
  assign n4845 = ~n3828 & ~n4844;
  assign n4846 = n4843 & ~n4845;
  assign n4847 = ~n4843 & n4845;
  assign po12  = n4846 | n4847;
  assign n4849 = ~n4836 & ~n4838;
  assign n4850 = ~n4818 & ~n4821;
  assign n4851 = ~n4812 & ~n4815;
  assign n4852 = ~n4791 & ~n4793;
  assign n4853 = n2638 & ~n3204;
  assign n4854 = n2573 & n3722;
  assign n4855 = n2566 & n3480;
  assign n4856 = n2568 & n3717;
  assign n4857 = ~n4853 & ~n4855;
  assign n4858 = ~n4856 & n4857;
  assign n4859 = ~n4854 & n4858;
  assign n4860 = n636 & ~n4859;
  assign n4861 = ~n636 & n4859;
  assign n4862 = ~n4860 & ~n4861;
  assign n4863 = n656 & n4789;
  assign n4864 = ~n656 & ~n4789;
  assign n4865 = ~n4863 & ~n4864;
  assign n4866 = ~n636 & n3182;
  assign n4867 = n4865 & n4866;
  assign n4868 = ~n4865 & ~n4866;
  assign n4869 = ~n4867 & ~n4868;
  assign n4870 = ~n4862 & ~n4869;
  assign n4871 = n4862 & n4869;
  assign n4872 = ~n4870 & ~n4871;
  assign n4873 = ~n4852 & ~n4872;
  assign n4874 = n4852 & n4872;
  assign n4875 = ~n4873 & ~n4874;
  assign n4876 = ~n4851 & n4875;
  assign n4877 = n4851 & ~n4875;
  assign n4878 = ~n4876 & ~n4877;
  assign n4879 = ~n4850 & n4878;
  assign n4880 = n4850 & ~n4878;
  assign n4881 = ~n4879 & ~n4880;
  assign n4882 = ~n337 & ~n342;
  assign n4883 = ~n353 & ~n424;
  assign n4884 = ~n497 & n4883;
  assign n4885 = n4882 & n4884;
  assign n4886 = ~n174 & ~n202;
  assign n4887 = ~n232 & ~n252;
  assign n4888 = ~n455 & n4887;
  assign n4889 = n436 & n4886;
  assign n4890 = n861 & n1025;
  assign n4891 = n4889 & n4890;
  assign n4892 = n3807 & n4888;
  assign n4893 = n4891 & n4892;
  assign n4894 = n4885 & n4893;
  assign n4895 = n1004 & n4894;
  assign n4896 = n2042 & n3663;
  assign n4897 = n4895 & n4896;
  assign n4898 = n4881 & ~n4897;
  assign n4899 = ~n4881 & n4897;
  assign n4900 = ~n4898 & ~n4899;
  assign n4901 = ~n4849 & n4900;
  assign n4902 = n4849 & ~n4900;
  assign n4903 = ~n4901 & ~n4902;
  assign n4904 = ~n4842 & ~n4903;
  assign n4905 = n4842 & n4903;
  assign n4906 = ~n4904 & ~n4905;
  assign n4907 = ~n4843 & n4844;
  assign n4908 = ~n3828 & ~n4907;
  assign n4909 = n4906 & ~n4908;
  assign n4910 = ~n4906 & n4908;
  assign po13  = n4909 | n4910;
  assign n4912 = ~n4898 & ~n4901;
  assign n4913 = ~n4876 & ~n4879;
  assign n4914 = ~n4862 & n4869;
  assign n4915 = ~n4873 & ~n4914;
  assign n4916 = ~n636 & ~n3204;
  assign n4917 = ~n4863 & ~n4867;
  assign n4918 = ~n4916 & n4917;
  assign n4919 = n4916 & ~n4917;
  assign n4920 = ~n4918 & ~n4919;
  assign n4921 = n2638 & n3480;
  assign n4922 = n2566 & n3717;
  assign n4923 = n2573 & ~n3844;
  assign n4924 = ~n4921 & ~n4922;
  assign n4925 = ~n4923 & n4924;
  assign n4926 = n636 & n4925;
  assign n4927 = ~n636 & ~n4925;
  assign n4928 = ~n4926 & ~n4927;
  assign n4929 = ~n4920 & n4928;
  assign n4930 = n4920 & ~n4928;
  assign n4931 = ~n4929 & ~n4930;
  assign n4932 = ~n4915 & n4931;
  assign n4933 = n4915 & ~n4931;
  assign n4934 = ~n4932 & ~n4933;
  assign n4935 = ~n4913 & n4934;
  assign n4936 = n4913 & ~n4934;
  assign n4937 = ~n4935 & ~n4936;
  assign n4938 = ~n177 & ~n246;
  assign n4939 = ~n303 & ~n339;
  assign n4940 = ~n455 & n4939;
  assign n4941 = n287 & n4938;
  assign n4942 = n596 & n2201;
  assign n4943 = n2268 & n3170;
  assign n4944 = n4942 & n4943;
  assign n4945 = n4940 & n4941;
  assign n4946 = n4944 & n4945;
  assign n4947 = n864 & n4946;
  assign n4948 = n855 & n1339;
  assign n4949 = n4947 & n4948;
  assign n4950 = n2024 & n4949;
  assign n4951 = ~n4937 & n4950;
  assign n4952 = n4937 & ~n4950;
  assign n4953 = ~n4951 & ~n4952;
  assign n4954 = ~n4912 & n4953;
  assign n4955 = n4912 & ~n4953;
  assign n4956 = ~n4954 & ~n4955;
  assign n4957 = ~n4905 & ~n4956;
  assign n4958 = n4905 & n4956;
  assign n4959 = ~n4957 & ~n4958;
  assign n4960 = ~n4906 & n4907;
  assign n4961 = ~n3828 & ~n4960;
  assign n4962 = n4959 & ~n4961;
  assign n4963 = ~n4959 & n4961;
  assign po14  = n4962 | n4963;
  assign n4965 = ~n4952 & ~n4954;
  assign n4966 = n2573 & ~n3842;
  assign n4967 = ~n2638 & ~n4966;
  assign n4968 = n3717 & ~n4967;
  assign n4969 = n636 & n4968;
  assign n4970 = ~n636 & ~n4968;
  assign n4971 = ~n4969 & ~n4970;
  assign n4972 = ~n636 & n3483;
  assign n4973 = n4971 & ~n4972;
  assign n4974 = n3483 & n4970;
  assign n4975 = ~n4973 & ~n4974;
  assign n4976 = ~n4916 & ~n4917;
  assign n4977 = ~n4929 & ~n4976;
  assign n4978 = n4975 & n4977;
  assign n4979 = ~n4975 & ~n4977;
  assign n4980 = ~n4978 & ~n4979;
  assign n4981 = ~n4932 & ~n4935;
  assign n4982 = ~n4980 & n4981;
  assign n4983 = n4980 & ~n4981;
  assign n4984 = ~n4982 & ~n4983;
  assign n4985 = ~n179 & ~n268;
  assign n4986 = ~n284 & n4985;
  assign n4987 = n1039 & n4986;
  assign n4988 = ~n158 & ~n285;
  assign n4989 = ~n328 & ~n358;
  assign n4990 = n4988 & n4989;
  assign n4991 = n564 & n843;
  assign n4992 = n3621 & n4991;
  assign n4993 = n4990 & n4992;
  assign n4994 = n4827 & n4993;
  assign n4995 = n976 & n4994;
  assign n4996 = n2210 & n4995;
  assign n4997 = n4987 & n4996;
  assign n4998 = n4984 & ~n4997;
  assign n4999 = ~n4984 & n4997;
  assign n5000 = ~n4998 & ~n4999;
  assign n5001 = ~n4965 & n5000;
  assign n5002 = n4965 & ~n5000;
  assign n5003 = ~n5001 & ~n5002;
  assign n5004 = ~n4958 & ~n5003;
  assign n5005 = n4958 & n5003;
  assign n5006 = ~n5004 & ~n5005;
  assign n5007 = ~n4959 & n4960;
  assign n5008 = ~n3828 & ~n5007;
  assign n5009 = n5006 & ~n5008;
  assign n5010 = ~n5006 & n5008;
  assign po15  = n5009 | n5010;
  assign n5012 = ~n4998 & ~n5001;
  assign n5013 = ~n216 & ~n327;
  assign n5014 = ~n478 & n5013;
  assign n5015 = n159 & n551;
  assign n5016 = n5014 & n5015;
  assign n5017 = n2102 & n5016;
  assign n5018 = n3593 & n4885;
  assign n5019 = n5017 & n5018;
  assign n5020 = n3657 & n5019;
  assign n5021 = n2156 & n5020;
  assign n5022 = ~n4971 & ~n4972;
  assign n5023 = ~n636 & n3480;
  assign n5024 = ~n4916 & n5023;
  assign n5025 = ~n5022 & ~n5024;
  assign n5026 = ~n4979 & ~n4983;
  assign n5027 = ~n3717 & n4916;
  assign n5028 = n3204 & ~n3712;
  assign n5029 = ~n636 & ~n5028;
  assign n5030 = ~n5027 & n5029;
  assign n5031 = n5026 & ~n5030;
  assign n5032 = ~n5026 & n5030;
  assign n5033 = ~n5031 & ~n5032;
  assign n5034 = n5025 & n5033;
  assign n5035 = ~n5025 & ~n5033;
  assign n5036 = ~n5034 & ~n5035;
  assign n5037 = n5021 & ~n5036;
  assign n5038 = ~n5021 & n5036;
  assign n5039 = ~n5037 & ~n5038;
  assign n5040 = n5012 & n5039;
  assign n5041 = ~n5012 & ~n5039;
  assign n5042 = ~n5040 & ~n5041;
  assign n5043 = ~n5005 & n5042;
  assign n5044 = n5005 & ~n5042;
  assign n5045 = ~n5043 & ~n5044;
  assign n5046 = ~n5006 & n5007;
  assign n5047 = ~n3828 & ~n5046;
  assign n5048 = n5045 & ~n5047;
  assign n5049 = ~n5045 & n5047;
  assign po16  = n5048 | n5049;
  assign n5051 = ~n5045 & n5046;
  assign n5052 = ~n3828 & ~n5051;
  assign n5053 = n5012 & ~n5038;
  assign n5054 = ~n5037 & ~n5053;
  assign n5055 = ~n129 & ~n150;
  assign n5056 = ~n200 & ~n255;
  assign n5057 = ~n479 & n5056;
  assign n5058 = n792 & n5055;
  assign n5059 = n861 & n2390;
  assign n5060 = n5058 & n5059;
  assign n5061 = n275 & n5057;
  assign n5062 = n5060 & n5061;
  assign n5063 = n438 & n5062;
  assign n5064 = n419 & n5063;
  assign n5065 = n3057 & n5064;
  assign n5066 = n5054 & ~n5065;
  assign n5067 = ~n5054 & n5065;
  assign n5068 = ~n5066 & ~n5067;
  assign n5069 = n5044 & n5068;
  assign n5070 = ~n5044 & ~n5068;
  assign n5071 = ~n5069 & ~n5070;
  assign n5072 = n5052 & n5071;
  assign n5073 = ~n5052 & ~n5071;
  assign po17  = ~n5072 & ~n5073;
  assign n5075 = n5051 & ~n5071;
  assign n5076 = ~n3828 & ~n5075;
  assign n5077 = ~n5066 & ~n5069;
  assign n5078 = ~n144 & ~n303;
  assign n5079 = ~n347 & ~n362;
  assign n5080 = ~n479 & n5079;
  assign n5081 = n5078 & n5080;
  assign n5082 = n559 & n867;
  assign n5083 = n5081 & n5082;
  assign n5084 = n981 & n2034;
  assign n5085 = n5083 & n5084;
  assign n5086 = n1050 & n5085;
  assign n5087 = n3639 & n5086;
  assign n5088 = n448 & n5087;
  assign n5089 = ~n5077 & n5088;
  assign n5090 = n5077 & ~n5088;
  assign n5091 = ~n5089 & ~n5090;
  assign n5092 = n5076 & n5091;
  assign n5093 = ~n5076 & ~n5091;
  assign po18  = n5092 | n5093;
  assign n5095 = n5066 & ~n5088;
  assign n5096 = ~n340 & ~n350;
  assign n5097 = ~n234 & ~n434;
  assign n5098 = ~n566 & n5097;
  assign n5099 = n3038 & n5096;
  assign n5100 = n567 & n5099;
  assign n5101 = n4250 & n5098;
  assign n5102 = n5100 & n5101;
  assign n5103 = n2501 & n5102;
  assign n5104 = n789 & n5103;
  assign n5105 = n4987 & n5104;
  assign n5106 = ~n5095 & n5105;
  assign n5107 = n5095 & ~n5105;
  assign n5108 = ~n5106 & ~n5107;
  assign n5109 = n5069 & ~n5088;
  assign n5110 = ~n5108 & ~n5109;
  assign n5111 = n5108 & n5109;
  assign n5112 = ~n5110 & ~n5111;
  assign n5113 = n5075 & n5091;
  assign n5114 = ~n3828 & ~n5113;
  assign n5115 = n5112 & ~n5114;
  assign n5116 = ~n5112 & n5114;
  assign po19  = n5115 | n5116;
  assign n5118 = ~n5112 & n5113;
  assign n5119 = ~n3828 & ~n5118;
  assign n5120 = ~n5107 & ~n5111;
  assign n5121 = ~n405 & n493;
  assign n5122 = n611 & n3589;
  assign n5123 = n4448 & n5122;
  assign n5124 = n4251 & n5121;
  assign n5125 = n5123 & n5124;
  assign n5126 = n664 & n5125;
  assign n5127 = n878 & n5126;
  assign n5128 = n4539 & n5127;
  assign n5129 = ~n5120 & n5128;
  assign n5130 = n5120 & ~n5128;
  assign n5131 = ~n5129 & ~n5130;
  assign n5132 = n5119 & n5131;
  assign n5133 = ~n5119 & ~n5131;
  assign po20  = n5132 | n5133;
  assign n5135 = n5107 & ~n5128;
  assign n5136 = ~n423 & n607;
  assign n5137 = n3195 & n5136;
  assign n5138 = n525 & n5137;
  assign n5139 = ~n5135 & n5138;
  assign n5140 = n5135 & ~n5138;
  assign n5141 = ~n5139 & ~n5140;
  assign n5142 = n5111 & ~n5128;
  assign n5143 = ~n5141 & ~n5142;
  assign n5144 = n5141 & n5142;
  assign n5145 = ~n5143 & ~n5144;
  assign n5146 = n5118 & n5131;
  assign n5147 = ~n3828 & ~n5146;
  assign n5148 = n5145 & ~n5147;
  assign n5149 = ~n5145 & n5147;
  assign po21  = n5148 | n5149;
  assign n5151 = ~n5145 & n5146;
  assign n5152 = ~n3828 & ~n5151;
  assign n5153 = n525 & n676;
  assign n5154 = ~n5140 & ~n5144;
  assign n5155 = n5153 & ~n5154;
  assign n5156 = ~n5153 & n5154;
  assign n5157 = ~n5155 & ~n5156;
  assign n5158 = n5152 & n5157;
  assign n5159 = ~n5152 & ~n5157;
  assign po22  = n5158 | n5159;
  assign n5161 = ~pi22  & n118;
  assign n5162 = n5151 & n5157;
  assign n5163 = ~n3828 & ~n5162;
  assign n5164 = ~n5153 & ~n5154;
  assign n5165 = n5140 & n5144;
  assign n5166 = n5164 & ~n5165;
  assign n5167 = n5163 & ~n5166;
  assign n5168 = ~n5163 & n5166;
  assign n5169 = ~n5161 & ~n5167;
  assign po23  = n5168 | ~n5169;
  assign n5171 = ~n5153 & n5165;
  assign n5172 = ~n5162 & ~n5171;
  assign n5173 = n5151 & n5164;
  assign n5174 = ~n5161 & ~n5173;
  assign n5175 = ~n5172 & n5174;
  assign po24  = ~n3828 & ~n5175;
endmodule
