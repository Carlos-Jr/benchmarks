module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 ,
    pi7 , pi8 , pi9 , pi10 , pi11 , pi12 ,
    pi13 , pi14 , pi15 , pi16 , pi17 , pi18 ,
    pi19 , pi20 , pi21 , pi22 , pi23 , pi24 ,
    pi25 , pi26 , pi27 , pi28 , pi29 , pi30 ,
    pi31 , pi32 , pi33 , pi34 , pi35 , pi36 ,
    pi37 , pi38 , pi39 , pi40 , pi41 , pi42 ,
    pi43 , pi44 , pi45 , pi46 , pi47 , pi48 ,
    pi49 , pi50 , pi51 , pi52 , pi53 , pi54 ,
    pi55 , pi56 , pi57 , pi58 , pi59 , pi60 ,
    pi61 , pi62 , pi63 , pi64 , pi65 , pi66 ,
    pi67 , pi68 , pi69 , pi70 , pi71 , pi72 ,
    pi73 , pi74 , pi75 , pi76 , pi77 , pi78 ,
    pi79 , pi80 , pi81 , pi82 , pi83 , pi84 ,
    pi85 , pi86 , pi87 , pi88 , pi89 , pi90 ,
    pi91 , pi92 , pi93 , pi94 , pi95 , pi96 ,
    pi97 , pi98 , pi99 , pi100 , pi101 , pi102 ,
    pi103 , pi104 , pi105 , pi106 , pi107 , pi108 ,
    pi109 , pi110 , pi111 , pi112 , pi113 , pi114 ,
    pi115 , pi116 , pi117 , pi118 , pi119 , pi120 ,
    pi121 , pi122 , pi123 , pi124 , pi125 , pi126 ,
    pi127 , pi128 , pi129 , pi130 , pi131 , pi132 , pi133 ,
    pi134 , pi135 , pi136 , pi137 , pi138 , pi139 ,
    pi140 , pi141 , pi142 , pi143 , pi144 , pi145 ,
    pi146 , pi147 , pi148 , pi149 , pi150 , pi151 ,
    pi152 , pi153 , pi154 , pi155 , pi156 , pi157 ,
    pi158 , pi159 , pi160 , pi161 , pi162 , pi163 ,
    pi164 , pi165 , pi166 , pi167 , pi168 , pi169 ,
    pi170 , pi171 , pi172 , pi173 , pi174 , pi175 ,
    pi176 , pi177 , pi178 , pi179 , pi180 , pi181 ,
    pi182 , pi183 , pi184 , pi185 , pi186 , pi187 ,
    pi188 , pi189 , pi190 , pi191 , pi192 , pi193 ,
    pi194 , pi195 , pi196 , pi197 , pi198 , pi199 ,
    pi200 , pi201 , pi202 , pi203 , pi204 , pi205 ,
    pi206 , pi207 , pi208 , pi209 , pi210 , pi211 ,
    pi212 , pi213 , pi214 , pi215 , pi216 , pi217 ,
    pi218 , pi219 , pi220 , pi221 , pi222 , pi223 ,
    pi224 , pi225 , pi226 , pi227 , pi228 , pi229 ,
    pi230 , pi231 , pi232 , pi233 , pi234 , pi235 ,
    pi236 , pi237 , pi238 , pi239 , pi240 , pi241 ,
    pi242 , pi243 , pi244 , pi245 , pi246 , pi247 ,
    pi248 , pi249 , pi250 , pi251 , pi252 , pi253 ,
    pi254 , pi255 , pi256 , pi257 , pi258 , pi259 ,
    pi260 , pi261 , pi262 , pi263 , pi264 , pi265 , pi266 ,
    pi267 , pi268 , pi269 , pi270 , pi271 , pi272 ,
    pi273 , pi274 , pi275 , pi276 , pi277 , pi278 ,
    pi279 , pi280 , pi281 , pi282 , pi283 , pi284 ,
    pi285 , pi286 , pi287 , pi288 , pi289 , pi290 ,
    pi291 , pi292 , pi293 , pi294 , pi295 , pi296 ,
    pi297 , pi298 , pi299 , pi300 , pi301 , pi302 ,
    pi303 , pi304 , pi305 , pi306 , pi307 , pi308 ,
    pi309 , pi310 , pi311 , pi312 , pi313 , pi314 ,
    pi315 , pi316 , pi317 , pi318 , pi319 , pi320 ,
    pi321 , pi322 , pi323 , pi324 , pi325 , pi326 ,
    pi327 , pi328 , pi329 , pi330 , pi331 , pi332 ,
    pi333 , pi334 , pi335 , pi336 , pi337 , pi338 ,
    pi339 , pi340 , pi341 , pi342 , pi343 , pi344 ,
    pi345 , pi346 , pi347 , pi348 , pi349 , pi350 ,
    pi351 , pi352 , pi353 , pi354 , pi355 , pi356 ,
    pi357 , pi358 , pi359 , pi360 , pi361 , pi362 ,
    pi363 , pi364 , pi365 , pi366 , pi367 , pi368 ,
    pi369 , pi370 , pi371 , pi372 , pi373 , pi374 ,
    pi375 , pi376 , pi377 , pi378 , pi379 , pi380 ,
    pi381 , pi382 , pi383 , pi384 , pi385 , pi386 ,
    pi387 , pi388 , pi389 , pi390 , pi391 , pi392 , pi393 ,
    pi394 , pi395 , pi396 , pi397 , pi398 , pi399 ,
    pi400 , pi401 , pi402 , pi403 , pi404 , pi405 ,
    pi406 , pi407 , pi408 , pi409 , pi410 , pi411 ,
    pi412 , pi413 , pi414 , pi415 , pi416 , pi417 ,
    pi418 , pi419 , pi420 , pi421 , pi422 , pi423 ,
    pi424 , pi425 , pi426 , pi427 , pi428 , pi429 ,
    pi430 , pi431 , pi432 , pi433 , pi434 , pi435 ,
    pi436 , pi437 , pi438 , pi439 , pi440 , pi441 ,
    pi442 , pi443 , pi444 , pi445 , pi446 , pi447 ,
    pi448 , pi449 , pi450 , pi451 , pi452 , pi453 ,
    pi454 , pi455 , pi456 , pi457 , pi458 , pi459 ,
    pi460 , pi461 , pi462 , pi463 , pi464 , pi465 ,
    pi466 , pi467 , pi468 , pi469 , pi470 , pi471 ,
    pi472 , pi473 , pi474 , pi475 , pi476 , pi477 ,
    pi478 , pi479 , pi480 , pi481 , pi482 , pi483 ,
    pi484 , pi485 , pi486 , pi487 , pi488 , pi489 ,
    pi490 , pi491 , pi492 , pi493 , pi494 , pi495 ,
    pi496 , pi497 , pi498 , pi499 , pi500 , pi501 ,
    pi502 , pi503 , pi504 , pi505 , pi506 , pi507 ,
    pi508 , pi509 , pi510 , pi511 ,
    po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ,
    po128 , po129   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 ,
    pi6 , pi7 , pi8 , pi9 , pi10 , pi11 ,
    pi12 , pi13 , pi14 , pi15 , pi16 , pi17 ,
    pi18 , pi19 , pi20 , pi21 , pi22 , pi23 ,
    pi24 , pi25 , pi26 , pi27 , pi28 , pi29 ,
    pi30 , pi31 , pi32 , pi33 , pi34 , pi35 ,
    pi36 , pi37 , pi38 , pi39 , pi40 , pi41 ,
    pi42 , pi43 , pi44 , pi45 , pi46 , pi47 ,
    pi48 , pi49 , pi50 , pi51 , pi52 , pi53 ,
    pi54 , pi55 , pi56 , pi57 , pi58 , pi59 ,
    pi60 , pi61 , pi62 , pi63 , pi64 , pi65 ,
    pi66 , pi67 , pi68 , pi69 , pi70 , pi71 ,
    pi72 , pi73 , pi74 , pi75 , pi76 , pi77 ,
    pi78 , pi79 , pi80 , pi81 , pi82 , pi83 ,
    pi84 , pi85 , pi86 , pi87 , pi88 , pi89 ,
    pi90 , pi91 , pi92 , pi93 , pi94 , pi95 ,
    pi96 , pi97 , pi98 , pi99 , pi100 , pi101 ,
    pi102 , pi103 , pi104 , pi105 , pi106 , pi107 ,
    pi108 , pi109 , pi110 , pi111 , pi112 , pi113 ,
    pi114 , pi115 , pi116 , pi117 , pi118 , pi119 ,
    pi120 , pi121 , pi122 , pi123 , pi124 , pi125 ,
    pi126 , pi127 , pi128 , pi129 , pi130 , pi131 ,
    pi132 , pi133 , pi134 , pi135 , pi136 , pi137 , pi138 ,
    pi139 , pi140 , pi141 , pi142 , pi143 , pi144 ,
    pi145 , pi146 , pi147 , pi148 , pi149 , pi150 ,
    pi151 , pi152 , pi153 , pi154 , pi155 , pi156 ,
    pi157 , pi158 , pi159 , pi160 , pi161 , pi162 ,
    pi163 , pi164 , pi165 , pi166 , pi167 , pi168 ,
    pi169 , pi170 , pi171 , pi172 , pi173 , pi174 ,
    pi175 , pi176 , pi177 , pi178 , pi179 , pi180 ,
    pi181 , pi182 , pi183 , pi184 , pi185 , pi186 ,
    pi187 , pi188 , pi189 , pi190 , pi191 , pi192 ,
    pi193 , pi194 , pi195 , pi196 , pi197 , pi198 ,
    pi199 , pi200 , pi201 , pi202 , pi203 , pi204 ,
    pi205 , pi206 , pi207 , pi208 , pi209 , pi210 ,
    pi211 , pi212 , pi213 , pi214 , pi215 , pi216 ,
    pi217 , pi218 , pi219 , pi220 , pi221 , pi222 ,
    pi223 , pi224 , pi225 , pi226 , pi227 , pi228 ,
    pi229 , pi230 , pi231 , pi232 , pi233 , pi234 ,
    pi235 , pi236 , pi237 , pi238 , pi239 , pi240 ,
    pi241 , pi242 , pi243 , pi244 , pi245 , pi246 ,
    pi247 , pi248 , pi249 , pi250 , pi251 , pi252 ,
    pi253 , pi254 , pi255 , pi256 , pi257 , pi258 ,
    pi259 , pi260 , pi261 , pi262 , pi263 , pi264 , pi265 ,
    pi266 , pi267 , pi268 , pi269 , pi270 , pi271 ,
    pi272 , pi273 , pi274 , pi275 , pi276 , pi277 ,
    pi278 , pi279 , pi280 , pi281 , pi282 , pi283 ,
    pi284 , pi285 , pi286 , pi287 , pi288 , pi289 ,
    pi290 , pi291 , pi292 , pi293 , pi294 , pi295 ,
    pi296 , pi297 , pi298 , pi299 , pi300 , pi301 ,
    pi302 , pi303 , pi304 , pi305 , pi306 , pi307 ,
    pi308 , pi309 , pi310 , pi311 , pi312 , pi313 ,
    pi314 , pi315 , pi316 , pi317 , pi318 , pi319 ,
    pi320 , pi321 , pi322 , pi323 , pi324 , pi325 ,
    pi326 , pi327 , pi328 , pi329 , pi330 , pi331 ,
    pi332 , pi333 , pi334 , pi335 , pi336 , pi337 ,
    pi338 , pi339 , pi340 , pi341 , pi342 , pi343 ,
    pi344 , pi345 , pi346 , pi347 , pi348 , pi349 ,
    pi350 , pi351 , pi352 , pi353 , pi354 , pi355 ,
    pi356 , pi357 , pi358 , pi359 , pi360 , pi361 ,
    pi362 , pi363 , pi364 , pi365 , pi366 , pi367 ,
    pi368 , pi369 , pi370 , pi371 , pi372 , pi373 ,
    pi374 , pi375 , pi376 , pi377 , pi378 , pi379 ,
    pi380 , pi381 , pi382 , pi383 , pi384 , pi385 ,
    pi386 , pi387 , pi388 , pi389 , pi390 , pi391 , pi392 ,
    pi393 , pi394 , pi395 , pi396 , pi397 , pi398 ,
    pi399 , pi400 , pi401 , pi402 , pi403 , pi404 ,
    pi405 , pi406 , pi407 , pi408 , pi409 , pi410 ,
    pi411 , pi412 , pi413 , pi414 , pi415 , pi416 ,
    pi417 , pi418 , pi419 , pi420 , pi421 , pi422 ,
    pi423 , pi424 , pi425 , pi426 , pi427 , pi428 ,
    pi429 , pi430 , pi431 , pi432 , pi433 , pi434 ,
    pi435 , pi436 , pi437 , pi438 , pi439 , pi440 ,
    pi441 , pi442 , pi443 , pi444 , pi445 , pi446 ,
    pi447 , pi448 , pi449 , pi450 , pi451 , pi452 ,
    pi453 , pi454 , pi455 , pi456 , pi457 , pi458 ,
    pi459 , pi460 , pi461 , pi462 , pi463 , pi464 ,
    pi465 , pi466 , pi467 , pi468 , pi469 , pi470 ,
    pi471 , pi472 , pi473 , pi474 , pi475 , pi476 ,
    pi477 , pi478 , pi479 , pi480 , pi481 , pi482 ,
    pi483 , pi484 , pi485 , pi486 , pi487 , pi488 ,
    pi489 , pi490 , pi491 , pi492 , pi493 , pi494 ,
    pi495 , pi496 , pi497 , pi498 , pi499 , pi500 ,
    pi501 , pi502 , pi503 , pi504 , pi505 , pi506 ,
    pi507 , pi508 , pi509 , pi510 , pi511 ;
  output po0 , po1 , po2 , po3 , po4 ,
    po5 , po6 , po7 , po8 , po9 ,
    po10 , po11 , po12 , po13 , po14 ,
    po15 , po16 , po17 , po18 , po19 ,
    po20 , po21 , po22 , po23 , po24 ,
    po25 , po26 , po27 , po28 , po29 ,
    po30 , po31 , po32 , po33 , po34 ,
    po35 , po36 , po37 , po38 , po39 ,
    po40 , po41 , po42 , po43 , po44 ,
    po45 , po46 , po47 , po48 , po49 ,
    po50 , po51 , po52 , po53 , po54 ,
    po55 , po56 , po57 , po58 , po59 ,
    po60 , po61 , po62 , po63 , po64 ,
    po65 , po66 , po67 , po68 , po69 ,
    po70 , po71 , po72 , po73 , po74 ,
    po75 , po76 , po77 , po78 , po79 ,
    po80 , po81 , po82 , po83 , po84 ,
    po85 , po86 , po87 , po88 , po89 ,
    po90 , po91 , po92 , po93 , po94 ,
    po95 , po96 , po97 , po98 , po99 ,
    po100 , po101 , po102 , po103 ,
    po104 , po105 , po106 , po107 ,
    po108 , po109 , po110 , po111 ,
    po112 , po113 , po114 , po115 ,
    po116 , po117 , po118 , po119 ,
    po120 , po121 , po122 , po123 ,
    po124 , po125 , po126 , po127 ,
    po128 , po129 ;
  wire n643, n644, n645, n646, n647, n648, n649,
    n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663,
    n664, n665, n666, n667, n668, n669, n670,
    n671, n672, n673, n674, n675, n676, n677,
    n678, n679, n680, n681, n682, n683, n684,
    n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698,
    n699, n700, n701, n702, n703, n704, n705,
    n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719,
    n720, n721, n722, n723, n724, n725, n726,
    n727, n728, n729, n730, n731, n732, n733,
    n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n743, n744, n745, n746, n747,
    n748, n749, n750, n751, n752, n753, n754,
    n755, n756, n757, n758, n759, n760, n761,
    n762, n763, n764, n765, n766, n767, n768,
    n769, n770, n771, n772, n773, n774, n775,
    n776, n777, n778, n779, n780, n781, n782,
    n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803,
    n804, n805, n806, n807, n808, n809, n810,
    n811, n812, n813, n814, n815, n816, n817,
    n818, n819, n820, n821, n822, n823, n824,
    n825, n826, n827, n828, n829, n830, n831,
    n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n851, n852,
    n853, n854, n855, n856, n857, n858, n859,
    n860, n861, n862, n863, n864, n865, n866,
    n867, n868, n869, n870, n871, n872, n873,
    n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887,
    n888, n889, n890, n891, n892, n893, n894,
    n895, n896, n897, n898, n899, n900, n901,
    n902, n903, n904, n905, n906, n907, n908,
    n909, n910, n911, n912, n913, n914, n915,
    n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929,
    n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943,
    n944, n945, n946, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978,
    n979, n980, n981, n982, n983, n984, n985,
    n986, n987, n988, n989, n990, n991, n992,
    n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011,
    n1012, n1013, n1014, n1015, n1016, n1017,
    n1018, n1019, n1020, n1021, n1022, n1023,
    n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1044, n1045, n1046, n1047,
    n1048, n1049, n1050, n1051, n1052, n1053,
    n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065,
    n1066, n1067, n1068, n1069, n1070, n1071,
    n1072, n1073, n1074, n1075, n1076, n1077,
    n1078, n1079, n1080, n1081, n1082, n1083,
    n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1107,
    n1108, n1109, n1110, n1111, n1112, n1113,
    n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125,
    n1126, n1127, n1128, n1129, n1130, n1131,
    n1132, n1133, n1134, n1135, n1136, n1137,
    n1138, n1139, n1140, n1141, n1142, n1143,
    n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155,
    n1156, n1157, n1158, n1159, n1160, n1161,
    n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173,
    n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185,
    n1186, n1187, n1188, n1189, n1190, n1191,
    n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203,
    n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215,
    n1216, n1217, n1218, n1219, n1220, n1221,
    n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233,
    n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245,
    n1246, n1247, n1248, n1249, n1250, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257,
    n1258, n1259, n1260, n1261, n1262, n1263,
    n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275,
    n1276, n1277, n1278, n1279, n1280, n1281,
    n1282, n1283, n1284, n1285, n1286, n1287,
    n1288, n1289, n1290, n1291, n1292, n1293,
    n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305,
    n1306, n1307, n1308, n1309, n1310, n1311,
    n1312, n1313, n1314, n1315, n1316, n1317,
    n1318, n1319, n1320, n1321, n1322, n1323,
    n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1344, n1345, n1346, n1347,
    n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365,
    n1366, n1367, n1368, n1369, n1370, n1371,
    n1372, n1373, n1374, n1375, n1376, n1377,
    n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395,
    n1396, n1397, n1398, n1399, n1400, n1401,
    n1402, n1403, n1404, n1405, n1406, n1407,
    n1408, n1409, n1410, n1411, n1412, n1413,
    n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425,
    n1426, n1427, n1428, n1429, n1430, n1431,
    n1432, n1433, n1434, n1435, n1436, n1437,
    n1438, n1439, n1440, n1441, n1442, n1443,
    n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461,
    n1462, n1463, n1464, n1465, n1466, n1467,
    n1468, n1469, n1470, n1471, n1472, n1473,
    n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497,
    n1498, n1499, n1500, n1501, n1502, n1503,
    n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527,
    n1528, n1529, n1530, n1531, n1532, n1533,
    n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1556, n1557,
    n1558, n1559, n1560, n1561, n1562, n1563,
    n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581,
    n1582, n1583, n1584, n1585, n1586, n1587,
    n1588, n1589, n1590, n1591, n1592, n1593,
    n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605,
    n1606, n1607, n1608, n1609, n1610, n1611,
    n1612, n1613, n1614, n1615, n1616, n1617,
    n1618, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635,
    n1636, n1637, n1638, n1639, n1640, n1641,
    n1642, n1643, n1644, n1645, n1646, n1647,
    n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665,
    n1666, n1667, n1668, n1669, n1670, n1671,
    n1672, n1673, n1674, n1675, n1676, n1677,
    n1678, n1679, n1680, n1681, n1682, n1683,
    n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695,
    n1696, n1697, n1698, n1699, n1700, n1701,
    n1702, n1703, n1704, n1705, n1706, n1707,
    n1708, n1709, n1710, n1711, n1712, n1713,
    n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731,
    n1732, n1733, n1734, n1735, n1736, n1737,
    n1738, n1739, n1740, n1741, n1742, n1743,
    n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1759, n1760, n1761,
    n1762, n1763, n1764, n1765, n1766, n1767,
    n1768, n1769, n1770, n1771, n1772, n1773,
    n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785,
    n1786, n1787, n1788, n1789, n1790, n1791,
    n1792, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803,
    n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815,
    n1816, n1817, n1818, n1819, n1820, n1821,
    n1822, n1823, n1824, n1825, n1826, n1827,
    n1828, n1829, n1830, n1831, n1832, n1833,
    n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845,
    n1846, n1847, n1848, n1849, n1850, n1851,
    n1852, n1853, n1854, n1855, n1856, n1857,
    n1858, n1859, n1860, n1861, n1862, n1863,
    n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875,
    n1876, n1877, n1878, n1879, n1880, n1881,
    n1882, n1883, n1884, n1885, n1886, n1887,
    n1888, n1889, n1890, n1891, n1892, n1893,
    n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905,
    n1906, n1907, n1908, n1909, n1910, n1911,
    n1912, n1913, n1914, n1915, n1916, n1917,
    n1918, n1919, n1920, n1921, n1922, n1923,
    n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935,
    n1936, n1937, n1938, n1939, n1940, n1941,
    n1942, n1943, n1944, n1945, n1946, n1947,
    n1948, n1949, n1950, n1951, n1952, n1953,
    n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965,
    n1966, n1967, n1968, n1969, n1970, n1971,
    n1972, n1973, n1974, n1975, n1976, n1977,
    n1978, n1979, n1980, n1981, n1982, n1983,
    n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995,
    n1996, n1997, n1998, n1999, n2000, n2001,
    n2002, n2003, n2004, n2005, n2006, n2007,
    n2008, n2009, n2010, n2011, n2012, n2013,
    n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025,
    n2026, n2027, n2028, n2029, n2030, n2031,
    n2032, n2033, n2034, n2035, n2036, n2037,
    n2038, n2039, n2040, n2041, n2042, n2043,
    n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055,
    n2056, n2057, n2058, n2059, n2060, n2061,
    n2062, n2063, n2064, n2065, n2066, n2067,
    n2068, n2069, n2070, n2071, n2072, n2073,
    n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085,
    n2086, n2087, n2088, n2089, n2090, n2091,
    n2092, n2093, n2094, n2095, n2096, n2097,
    n2098, n2099, n2100, n2101, n2102, n2103,
    n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115,
    n2116, n2117, n2118, n2119, n2120, n2121,
    n2122, n2123, n2124, n2125, n2126, n2127,
    n2128, n2129, n2130, n2131, n2132, n2133,
    n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145,
    n2146, n2147, n2148, n2149, n2150, n2151,
    n2152, n2153, n2154, n2155, n2156, n2157,
    n2158, n2159, n2160, n2161, n2162, n2163,
    n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175,
    n2176, n2177, n2178, n2179, n2180, n2181,
    n2182, n2183, n2184, n2185, n2186, n2187,
    n2188, n2189, n2190, n2191, n2192, n2193,
    n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205,
    n2206, n2207, n2208, n2209, n2210, n2211,
    n2212, n2213, n2214, n2215, n2216, n2217,
    n2218, n2219, n2220, n2221, n2222, n2223,
    n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235,
    n2236, n2237, n2238, n2239, n2240, n2241,
    n2242, n2243, n2244, n2245, n2246, n2247,
    n2248, n2249, n2250, n2251, n2252, n2253,
    n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265,
    n2266, n2267, n2268, n2269, n2270, n2271,
    n2272, n2273, n2274, n2275, n2276, n2277,
    n2278, n2279, n2280, n2281, n2282, n2283,
    n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295,
    n2296, n2297, n2298, n2299, n2300, n2301,
    n2302, n2303, n2304, n2305, n2306, n2307,
    n2308, n2309, n2310, n2311, n2312, n2313,
    n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325,
    n2326, n2327, n2328, n2329, n2330, n2331,
    n2332, n2333, n2334, n2335, n2336, n2337,
    n2338, n2339, n2340, n2341, n2342, n2343,
    n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355,
    n2356, n2357, n2358, n2359, n2360, n2361,
    n2362, n2363, n2364, n2365, n2366, n2367,
    n2368, n2369, n2370, n2371, n2372, n2373,
    n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385,
    n2386, n2387, n2388, n2389, n2390, n2391,
    n2392, n2393, n2394, n2395, n2396, n2397,
    n2398, n2399, n2400, n2401, n2402, n2403,
    n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415,
    n2416, n2417, n2418, n2419, n2420, n2421,
    n2422, n2423, n2424, n2425, n2426, n2427,
    n2428, n2429, n2430, n2431, n2432, n2433,
    n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445,
    n2446, n2447, n2448, n2449, n2450, n2451,
    n2452, n2453, n2454, n2455, n2456, n2457,
    n2458, n2459, n2460, n2461, n2462, n2463,
    n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475,
    n2476, n2477, n2478, n2479, n2480, n2481,
    n2482, n2483, n2484, n2485, n2486, n2487,
    n2488, n2489, n2490, n2491, n2492, n2493,
    n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505,
    n2506, n2507, n2508, n2509, n2510, n2511,
    n2512, n2513, n2514, n2515, n2516, n2517,
    n2518, n2519, n2520, n2521, n2522, n2523,
    n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535,
    n2536, n2537, n2538, n2539, n2540, n2541,
    n2542, n2543, n2544, n2545, n2546, n2547,
    n2548, n2549, n2550, n2551, n2552, n2553,
    n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565,
    n2566, n2567, n2568, n2569, n2570, n2571,
    n2572, n2573, n2574, n2575, n2576, n2577,
    n2578, n2579, n2580, n2581, n2582, n2583,
    n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595,
    n2596, n2597, n2598, n2599, n2600, n2601,
    n2602, n2603, n2604, n2605, n2606, n2607,
    n2608, n2609, n2610, n2611, n2612, n2613,
    n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625,
    n2626, n2627, n2628, n2629, n2630, n2631,
    n2632, n2633, n2634, n2635, n2636, n2637,
    n2638, n2639, n2640, n2641, n2642, n2643,
    n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655,
    n2656, n2657, n2658, n2659, n2660, n2661,
    n2662, n2663, n2664, n2665, n2666, n2667,
    n2668, n2669, n2670, n2671, n2672, n2673,
    n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685,
    n2686, n2687, n2688, n2689, n2690, n2691,
    n2692, n2693, n2694, n2695, n2696, n2697,
    n2698, n2699, n2700, n2701, n2702, n2703,
    n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715,
    n2716, n2717, n2718, n2719, n2720, n2721,
    n2722, n2723, n2724, n2725, n2726, n2727,
    n2728, n2729, n2730, n2731, n2732, n2733,
    n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745,
    n2746, n2747, n2748, n2749, n2750, n2751,
    n2752, n2753, n2754, n2755, n2756, n2757,
    n2758, n2759, n2760, n2761, n2762, n2763,
    n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775,
    n2776, n2777, n2778, n2779, n2780, n2781,
    n2782, n2783, n2784, n2785, n2786, n2787,
    n2788, n2789, n2790, n2791, n2792, n2793,
    n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805,
    n2806, n2807, n2808, n2809, n2810, n2811,
    n2812, n2813, n2814, n2815, n2816, n2817,
    n2818, n2819, n2820, n2821, n2822, n2823,
    n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835,
    n2836, n2837, n2838, n2839, n2840, n2841,
    n2842, n2843, n2844, n2845, n2846, n2847,
    n2848, n2849, n2850, n2851, n2852, n2853,
    n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865,
    n2866, n2867, n2868, n2869, n2870, n2871,
    n2872, n2873, n2874, n2875, n2876, n2877,
    n2878, n2879, n2880, n2881, n2882, n2883,
    n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895,
    n2896, n2897, n2898, n2899, n2900, n2901,
    n2902, n2903, n2904, n2905, n2906, n2907,
    n2908, n2909, n2910, n2911, n2912, n2913,
    n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925,
    n2926, n2927, n2928, n2929, n2930, n2931,
    n2932, n2933, n2934, n2935, n2936, n2937,
    n2938, n2939, n2940, n2941, n2942, n2943,
    n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955,
    n2956, n2957, n2958, n2959, n2960, n2961,
    n2962, n2963, n2964, n2965, n2966, n2967,
    n2968, n2969, n2970, n2971, n2972, n2973,
    n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985,
    n2986, n2987, n2988, n2989, n2990, n2991,
    n2992, n2993, n2994, n2995, n2996, n2997,
    n2998, n2999, n3000, n3001, n3002, n3003,
    n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015,
    n3016, n3017, n3018, n3019, n3020, n3021,
    n3022, n3023, n3024, n3025, n3026, n3027,
    n3028, n3029, n3030, n3031, n3032, n3033,
    n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045,
    n3046, n3047, n3048, n3049, n3050, n3051,
    n3052, n3053, n3054, n3055, n3056, n3057,
    n3058, n3059, n3060, n3061, n3062, n3063,
    n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075,
    n3076, n3077, n3078, n3079, n3080, n3081,
    n3082, n3083, n3084, n3085, n3086, n3087,
    n3088, n3089, n3090, n3091, n3092, n3093,
    n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105,
    n3106, n3107, n3108, n3109, n3110, n3111,
    n3112, n3113, n3114, n3115, n3116, n3117,
    n3118, n3119, n3120, n3121, n3122, n3123,
    n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135,
    n3136, n3137, n3138, n3139, n3140, n3141,
    n3142, n3143, n3144, n3145, n3146, n3147,
    n3148, n3149, n3150, n3151, n3152, n3153,
    n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165,
    n3166, n3167, n3168, n3169, n3170, n3171,
    n3172, n3173, n3174, n3175, n3176, n3177,
    n3178, n3179, n3180, n3181, n3182, n3183,
    n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195,
    n3196, n3197, n3198, n3199, n3200, n3201,
    n3202, n3203, n3204, n3205, n3206, n3207,
    n3208, n3209, n3210, n3211, n3212, n3213,
    n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225,
    n3226, n3227, n3228, n3229, n3230, n3231,
    n3232, n3233, n3234, n3235, n3236, n3237,
    n3238, n3239, n3240, n3241, n3242, n3243,
    n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255,
    n3256, n3257, n3258, n3259, n3260, n3261,
    n3262, n3263, n3264, n3265, n3266, n3267,
    n3268, n3269, n3270, n3271, n3272, n3273,
    n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285,
    n3286, n3287, n3288, n3289, n3290, n3291,
    n3292, n3293, n3294, n3295, n3296, n3297,
    n3298, n3299, n3300, n3301, n3302, n3303,
    n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315,
    n3316, n3317, n3318, n3319, n3320, n3321,
    n3322, n3323, n3324, n3325, n3326, n3327,
    n3328, n3329, n3330, n3331, n3332, n3333,
    n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345,
    n3346, n3347, n3348, n3349, n3350, n3351,
    n3352, n3353, n3354, n3355, n3356, n3357,
    n3358, n3359, n3360, n3361, n3362, n3363,
    n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375,
    n3376, n3377, n3378, n3379, n3380, n3381,
    n3382, n3383, n3384, n3385, n3386, n3387,
    n3388, n3389, n3390, n3391, n3392, n3393,
    n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405,
    n3406, n3407, n3408, n3409, n3410, n3411,
    n3412, n3413, n3414, n3415, n3416, n3417,
    n3418, n3419, n3420, n3421, n3422, n3423,
    n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435,
    n3436, n3437, n3438, n3439, n3440, n3441,
    n3442, n3443, n3444, n3445, n3446, n3447,
    n3448, n3449, n3450, n3451, n3452, n3453,
    n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465,
    n3466, n3467, n3468, n3469, n3470, n3471,
    n3472, n3473, n3474, n3475, n3476, n3477,
    n3478, n3479, n3480, n3481, n3482, n3483,
    n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495,
    n3496, n3497, n3498, n3499, n3500, n3501,
    n3502, n3503, n3504, n3505, n3506, n3507,
    n3508, n3509, n3510, n3511, n3512, n3513,
    n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525,
    n3526, n3527, n3528, n3529, n3530, n3531,
    n3532, n3533, n3534, n3535, n3536, n3537,
    n3538, n3539, n3540, n3541, n3542, n3543,
    n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555,
    n3556, n3557, n3558, n3559, n3560, n3561,
    n3562, n3563, n3564, n3565, n3566, n3567,
    n3568, n3569, n3570, n3571, n3572, n3573,
    n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585,
    n3586, n3587, n3588, n3589, n3590, n3591,
    n3592, n3593, n3594, n3595, n3596, n3597,
    n3598, n3599, n3600, n3601, n3602, n3603,
    n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615,
    n3616, n3617, n3618, n3619, n3620, n3621,
    n3622, n3623, n3624, n3625, n3626, n3627,
    n3628, n3629, n3630, n3631, n3632, n3633,
    n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645,
    n3646, n3647, n3648, n3649, n3650, n3651,
    n3652, n3653, n3654, n3655, n3656, n3657,
    n3658, n3659, n3660, n3661, n3662, n3663,
    n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675,
    n3676, n3677, n3678, n3679, n3680, n3681,
    n3682, n3683, n3684, n3685, n3686, n3687,
    n3688, n3689, n3690, n3691, n3692, n3693,
    n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705,
    n3706, n3707, n3708, n3709, n3710, n3711,
    n3712, n3713, n3714, n3715, n3716, n3717,
    n3718, n3719, n3720, n3721, n3722, n3723,
    n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735,
    n3736, n3737, n3738, n3739, n3740, n3741,
    n3742, n3743, n3744, n3745, n3746, n3747,
    n3748, n3749, n3750, n3751, n3752, n3753,
    n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765,
    n3766, n3767, n3768, n3769, n3770, n3771,
    n3772, n3773, n3774, n3775, n3776, n3777,
    n3778, n3779, n3780, n3781, n3782, n3783,
    n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795,
    n3796, n3797, n3798, n3799, n3800, n3801,
    n3802, n3803, n3804, n3805, n3806, n3807,
    n3808, n3809, n3810, n3811, n3812, n3813,
    n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825,
    n3826, n3827, n3828, n3829, n3830, n3831,
    n3832, n3833, n3834, n3835, n3836, n3837,
    n3838, n3839, n3840, n3841, n3842, n3843,
    n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855,
    n3856, n3857, n3858, n3859, n3860, n3861,
    n3862, n3863, n3864, n3865, n3866, n3867,
    n3868, n3869, n3870, n3871, n3872, n3873,
    n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885,
    n3886, n3887, n3888, n3889, n3890, n3891,
    n3892, n3893, n3894, n3895, n3896, n3897,
    n3898, n3899, n3900, n3901, n3902, n3903,
    n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915,
    n3916, n3917, n3918, n3919, n3920, n3921,
    n3922, n3923, n3924, n3925, n3926, n3927,
    n3928, n3929, n3930, n3931, n3932, n3933,
    n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945,
    n3946, n3947, n3948, n3949, n3950, n3951,
    n3952, n3953, n3954, n3955, n3956, n3957,
    n3958, n3959, n3960, n3961, n3962, n3963,
    n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975,
    n3976, n3977, n3978, n3979, n3980, n3981,
    n3982, n3983, n3984, n3985, n3986, n3987,
    n3988, n3989, n3990, n3991, n3992, n3993,
    n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005,
    n4006, n4007, n4008, n4009, n4010, n4011,
    n4012, n4013, n4014, n4015, n4016, n4017,
    n4018, n4019, n4020, n4021, n4022, n4023,
    n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035,
    n4036, n4037, n4038, n4039, n4040, n4041,
    n4042, n4043, n4044, n4045, n4046, n4047,
    n4048, n4049, n4050, n4051, n4052, n4053,
    n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065,
    n4066, n4067, n4068, n4069, n4070, n4071,
    n4072, n4073, n4074, n4075, n4076, n4077,
    n4078, n4079, n4080, n4081, n4082, n4083,
    n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095,
    n4096, n4097, n4098, n4099, n4100, n4101,
    n4102, n4103, n4104, n4105, n4106, n4107,
    n4108, n4109, n4110, n4111, n4112, n4113,
    n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125,
    n4126, n4127, n4128, n4129, n4130, n4131,
    n4132, n4133, n4134, n4135, n4136, n4137,
    n4138, n4139, n4140, n4141, n4142, n4143,
    n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155,
    n4156, n4157, n4158, n4159, n4160, n4161,
    n4162, n4163, n4164, n4165, n4166, n4167,
    n4168, n4169, n4170, n4171, n4172, n4173,
    n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185,
    n4186, n4187, n4188, n4189, n4190, n4191,
    n4192, n4193, n4194, n4195, n4196, n4197,
    n4198, n4199, n4200, n4201, n4202, n4203,
    n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215,
    n4216, n4217, n4218, n4219, n4220, n4221,
    n4222, n4223, n4224, n4225, n4226, n4227,
    n4228, n4229, n4230, n4231, n4232, n4233,
    n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245,
    n4246, n4247, n4248, n4249, n4250, n4251,
    n4252, n4253, n4254, n4255, n4256, n4257,
    n4258, n4259, n4260, n4261, n4262, n4263,
    n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275,
    n4276, n4277, n4278, n4279, n4280, n4281,
    n4282, n4283, n4284, n4285, n4286, n4287,
    n4288, n4289, n4290, n4291, n4292, n4293,
    n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305,
    n4306, n4307, n4308, n4309, n4310, n4311,
    n4312, n4313, n4314, n4315, n4316, n4317,
    n4318, n4319, n4320, n4321, n4322, n4323,
    n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335,
    n4336, n4337, n4338, n4339, n4340, n4341,
    n4342, n4343, n4344, n4345, n4346, n4347,
    n4348, n4349, n4350, n4351, n4352, n4353,
    n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365,
    n4366, n4367, n4368, n4369, n4370, n4371,
    n4372, n4373, n4374, n4375, n4376, n4377,
    n4378, n4379, n4380, n4381, n4382, n4383,
    n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395,
    n4396, n4397, n4398, n4399, n4400, n4401,
    n4402, n4403, n4404, n4405, n4406, n4407,
    n4408, n4409, n4410, n4411, n4412, n4413,
    n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425,
    n4426, n4427, n4428, n4429, n4430, n4431,
    n4432, n4433, n4434, n4435, n4436, n4437,
    n4438, n4439, n4440, n4441, n4442, n4443,
    n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4455,
    n4456, n4457, n4458, n4459, n4460, n4461,
    n4462, n4463, n4464, n4465, n4466, n4467,
    n4468, n4469, n4470, n4471, n4472, n4473,
    n4474, n4475, n4476, n4477, n4478, n4479,
    n4480, n4481, n4482, n4483, n4484, n4485,
    n4486, n4487, n4488, n4489, n4490, n4491,
    n4492, n4493, n4494, n4495, n4496, n4497,
    n4498, n4499, n4500, n4501, n4502, n4503,
    n4504, n4505, n4506, n4507, n4508, n4509,
    n4510, n4511, n4512, n4513, n4514, n4515,
    n4516, n4517, n4518, n4519, n4520, n4521,
    n4522, n4523, n4524, n4525, n4526, n4527,
    n4528, n4529, n4530, n4531, n4532, n4533,
    n4534, n4535, n4536, n4537, n4538, n4539,
    n4540, n4541, n4542, n4543, n4544, n4545,
    n4546, n4547, n4548, n4549, n4550, n4551,
    n4552, n4553, n4554, n4555, n4556, n4557,
    n4558, n4559, n4560, n4561, n4562, n4563,
    n4564, n4565, n4566, n4567, n4568, n4569,
    n4570, n4571, n4572, n4573, n4574, n4575,
    n4576, n4577, n4578, n4579, n4580, n4581,
    n4582, n4583, n4584, n4585, n4586, n4587,
    n4588, n4589, n4590, n4591, n4592, n4593,
    n4594, n4595, n4596, n4597, n4598, n4599,
    n4600, n4601, n4602, n4603, n4604, n4605,
    n4606, n4607, n4608, n4609, n4610, n4611,
    n4612, n4613, n4614, n4615, n4616, n4617,
    n4618, n4619, n4620, n4621, n4622, n4623,
    n4624, n4625, n4626, n4627, n4628, n4629,
    n4630, n4631, n4632, n4633, n4634, n4635,
    n4636, n4637, n4638, n4639, n4640, n4641,
    n4642, n4643, n4644, n4645, n4646, n4647,
    n4648, n4649, n4650, n4651, n4652, n4653,
    n4654, n4655, n4656, n4657, n4658, n4659,
    n4660, n4661, n4662, n4663, n4664, n4665,
    n4666, n4667, n4668, n4669, n4670, n4671,
    n4672, n4673, n4674, n4675, n4676, n4677,
    n4678, n4679, n4680, n4681, n4682, n4683,
    n4684, n4685, n4686, n4687, n4688, n4689,
    n4690, n4691, n4692, n4693, n4694, n4695,
    n4696, n4697, n4698, n4699, n4700, n4701,
    n4702, n4703, n4704, n4705, n4706, n4707,
    n4708, n4709, n4710, n4711, n4712, n4713,
    n4714, n4715, n4716, n4717, n4718, n4719,
    n4720, n4721, n4722, n4723, n4724, n4725,
    n4726, n4727, n4728, n4729, n4730, n4731,
    n4732, n4733, n4734, n4735, n4736, n4737,
    n4738, n4739, n4740, n4741, n4742, n4743,
    n4744, n4745, n4746, n4747, n4748, n4749,
    n4750, n4751, n4752, n4753, n4754, n4755,
    n4756, n4757, n4758, n4759, n4760, n4761,
    n4762, n4763, n4764, n4765, n4766, n4767,
    n4768, n4769, n4770, n4771, n4772, n4773,
    n4774, n4775, n4776, n4777, n4778, n4779,
    n4780, n4781, n4782, n4783, n4784, n4785,
    n4786, n4787, n4788, n4789, n4790, n4791,
    n4792, n4793, n4794, n4795, n4796, n4797,
    n4798, n4799, n4800, n4801, n4802, n4803,
    n4804, n4805, n4806, n4807, n4808, n4809,
    n4810, n4811, n4812, n4813, n4814, n4815,
    n4816, n4817, n4818, n4819, n4820, n4821,
    n4822, n4823, n4824, n4825, n4826, n4827,
    n4828, n4829, n4830, n4831, n4832, n4833,
    n4834, n4835, n4836, n4837, n4838, n4839,
    n4840, n4841, n4842, n4843, n4844, n4845,
    n4846, n4847, n4848, n4849, n4850, n4851,
    n4852, n4853, n4854, n4855, n4856, n4857,
    n4858, n4859, n4860, n4861, n4862, n4863,
    n4864, n4865, n4866, n4867, n4868, n4869,
    n4870, n4871, n4872, n4873, n4874, n4875,
    n4876, n4877, n4878, n4879, n4880, n4881,
    n4882, n4883, n4884, n4885, n4886, n4887,
    n4888, n4889, n4890, n4891, n4892, n4893,
    n4894, n4895, n4896, n4897, n4898, n4899,
    n4900, n4901, n4902, n4903, n4904, n4905,
    n4906, n4907, n4908, n4909, n4910, n4911,
    n4912, n4913, n4914, n4915, n4916, n4917,
    n4918, n4919, n4920, n4921, n4922, n4923,
    n4924, n4925, n4926, n4927, n4928, n4929,
    n4930, n4931, n4932, n4933, n4934, n4935,
    n4936, n4937, n4938, n4943;
  assign n643 = ~pi26  & pi154 ;
  assign n644 = pi25  & ~pi153 ;
  assign n645 = ~pi25  & pi153 ;
  assign n646 = pi24  & ~pi152 ;
  assign n647 = ~pi24  & pi152 ;
  assign n648 = pi23  & ~pi151 ;
  assign n649 = ~pi23  & pi151 ;
  assign n650 = pi22  & ~pi150 ;
  assign n651 = ~pi22  & pi150 ;
  assign n652 = pi21  & ~pi149 ;
  assign n653 = ~pi21  & pi149 ;
  assign n654 = pi20  & ~pi148 ;
  assign n655 = ~pi20  & pi148 ;
  assign n656 = pi19  & ~pi147 ;
  assign n657 = ~pi19  & pi147 ;
  assign n658 = pi18  & ~pi146 ;
  assign n659 = ~pi18  & pi146 ;
  assign n660 = pi17  & ~pi145 ;
  assign n661 = ~pi17  & pi145 ;
  assign n662 = pi16  & ~pi144 ;
  assign n663 = ~pi16  & pi144 ;
  assign n664 = pi15  & ~pi143 ;
  assign n665 = ~pi15  & pi143 ;
  assign n666 = pi14  & ~pi142 ;
  assign n667 = ~pi14  & pi142 ;
  assign n668 = pi13  & ~pi141 ;
  assign n669 = ~pi13  & pi141 ;
  assign n670 = pi12  & ~pi140 ;
  assign n671 = ~pi12  & pi140 ;
  assign n672 = pi11  & ~pi139 ;
  assign n673 = ~pi11  & pi139 ;
  assign n674 = pi10  & ~pi138 ;
  assign n675 = ~pi10  & pi138 ;
  assign n676 = pi9  & ~pi137 ;
  assign n677 = ~pi9  & pi137 ;
  assign n678 = pi8  & ~pi136 ;
  assign n679 = ~pi8  & pi136 ;
  assign n680 = pi7  & ~pi135 ;
  assign n681 = ~pi7  & pi135 ;
  assign n682 = pi6  & ~pi134 ;
  assign n683 = ~pi6  & pi134 ;
  assign n684 = pi5  & ~pi133 ;
  assign n685 = ~pi5  & pi133 ;
  assign n686 = pi4  & ~pi132 ;
  assign n687 = ~pi4  & pi132 ;
  assign n688 = pi3  & ~pi131 ;
  assign n689 = ~pi3  & pi131 ;
  assign n690 = pi2  & ~pi130 ;
  assign n691 = pi1  & ~pi129 ;
  assign n692 = pi0  & ~pi128 ;
  assign n693 = ~n691 & ~n692;
  assign n694 = ~pi2  & pi130 ;
  assign n695 = ~pi1  & pi129 ;
  assign n696 = ~n694 & ~n695;
  assign n697 = n692 & ~n695;
  assign n698 = ~n691 & ~n697;
  assign n699 = ~n694 & ~n698;
  assign n700 = ~n693 & n696;
  assign n701 = ~n690 & ~n4684;
  assign n702 = ~n689 & ~n701;
  assign n703 = ~n688 & ~n702;
  assign n704 = ~n687 & ~n703;
  assign n705 = ~pi4  & n703;
  assign n706 = ~pi132  & ~n705;
  assign n707 = pi4  & ~n703;
  assign n708 = ~n706 & ~n707;
  assign n709 = ~n686 & ~n704;
  assign n710 = ~n685 & ~n4685;
  assign n711 = ~pi5  & n4685;
  assign n712 = ~pi133  & ~n711;
  assign n713 = pi5  & ~n4685;
  assign n714 = ~n712 & ~n713;
  assign n715 = ~n684 & ~n710;
  assign n716 = ~n683 & ~n4686;
  assign n717 = ~n682 & ~n716;
  assign n718 = ~n681 & ~n717;
  assign n719 = ~n680 & ~n718;
  assign n720 = ~n679 & ~n719;
  assign n721 = ~pi8  & n719;
  assign n722 = ~pi136  & ~n721;
  assign n723 = pi8  & ~n719;
  assign n724 = ~n722 & ~n723;
  assign n725 = ~n678 & ~n720;
  assign n726 = ~n677 & ~n4687;
  assign n727 = ~pi9  & n4687;
  assign n728 = ~pi137  & ~n727;
  assign n729 = pi9  & ~n4687;
  assign n730 = ~n728 & ~n729;
  assign n731 = ~n676 & ~n726;
  assign n732 = ~n675 & ~n4688;
  assign n733 = ~n674 & ~n732;
  assign n734 = ~n673 & ~n733;
  assign n735 = ~n672 & ~n734;
  assign n736 = ~n671 & ~n735;
  assign n737 = ~n670 & ~n736;
  assign n738 = ~n669 & ~n737;
  assign n739 = ~n668 & ~n738;
  assign n740 = ~n667 & ~n739;
  assign n741 = ~n666 & ~n740;
  assign n742 = ~n665 & ~n741;
  assign n743 = ~n664 & ~n742;
  assign n744 = ~n663 & ~n743;
  assign n745 = ~pi16  & n743;
  assign n746 = ~pi144  & ~n745;
  assign n747 = pi16  & ~n743;
  assign n748 = ~n746 & ~n747;
  assign n749 = ~n662 & ~n744;
  assign n750 = ~n661 & ~n4689;
  assign n751 = ~pi17  & n4689;
  assign n752 = ~pi145  & ~n751;
  assign n753 = pi17  & ~n4689;
  assign n754 = ~n752 & ~n753;
  assign n755 = ~n660 & ~n750;
  assign n756 = ~n659 & ~n4690;
  assign n757 = ~n658 & ~n756;
  assign n758 = ~n657 & ~n757;
  assign n759 = ~n656 & ~n758;
  assign n760 = ~n655 & ~n759;
  assign n761 = ~n654 & ~n760;
  assign n762 = ~n653 & ~n761;
  assign n763 = ~n652 & ~n762;
  assign n764 = ~n651 & ~n763;
  assign n765 = ~n650 & ~n764;
  assign n766 = ~n649 & ~n765;
  assign n767 = ~n648 & ~n766;
  assign n768 = ~n647 & ~n767;
  assign n769 = ~pi24  & n767;
  assign n770 = ~pi152  & ~n769;
  assign n771 = pi24  & ~n767;
  assign n772 = ~n770 & ~n771;
  assign n773 = ~n646 & ~n768;
  assign n774 = ~n645 & ~n4691;
  assign n775 = ~pi25  & n4691;
  assign n776 = ~pi153  & ~n775;
  assign n777 = pi25  & ~n4691;
  assign n778 = ~n776 & ~n777;
  assign n779 = ~n644 & ~n774;
  assign n780 = ~n643 & ~n4692;
  assign n781 = pi26  & ~pi154 ;
  assign n782 = pi27  & ~pi155 ;
  assign n783 = ~n781 & ~n782;
  assign n784 = ~n780 & n783;
  assign n785 = ~pi27  & pi155 ;
  assign n786 = ~pi28  & pi156 ;
  assign n787 = ~n785 & ~n786;
  assign n788 = ~n780 & ~n781;
  assign n789 = ~n785 & ~n788;
  assign n790 = ~n782 & ~n789;
  assign n791 = ~n786 & ~n790;
  assign n792 = ~n784 & n787;
  assign n793 = pi28  & ~pi156 ;
  assign n794 = pi29  & ~pi157 ;
  assign n795 = ~n793 & ~n794;
  assign n796 = ~n4693 & n795;
  assign n797 = ~pi29  & pi157 ;
  assign n798 = ~pi30  & pi158 ;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~n4693 & ~n793;
  assign n801 = ~n797 & ~n800;
  assign n802 = ~n794 & ~n801;
  assign n803 = ~n798 & ~n802;
  assign n804 = ~n796 & n799;
  assign n805 = pi30  & ~pi158 ;
  assign n806 = pi31  & ~pi159 ;
  assign n807 = ~n805 & ~n806;
  assign n808 = ~n4694 & n807;
  assign n809 = ~pi37  & pi165 ;
  assign n810 = ~pi36  & pi164 ;
  assign n811 = ~pi164  & ~n809;
  assign n812 = pi36  & ~n809;
  assign n813 = ~n811 & ~n812;
  assign n814 = ~n809 & ~n810;
  assign n815 = ~pi33  & pi161 ;
  assign n816 = ~pi31  & pi159 ;
  assign n817 = ~pi32  & pi160 ;
  assign n818 = ~n816 & ~n817;
  assign n819 = ~n815 & ~n816;
  assign n820 = ~n817 & n819;
  assign n821 = ~n815 & n818;
  assign n822 = ~pi35  & pi163 ;
  assign n823 = ~pi34  & pi162 ;
  assign n824 = ~n822 & ~n823;
  assign n825 = ~pi39  & pi167 ;
  assign n826 = ~pi38  & pi166 ;
  assign n827 = ~n825 & ~n826;
  assign n828 = n824 & n827;
  assign n829 = n4696 & n828;
  assign n830 = ~n4695 & n827;
  assign n831 = n4696 & n824;
  assign n832 = n830 & n831;
  assign n833 = ~n4695 & n829;
  assign n834 = ~n4694 & ~n805;
  assign n835 = ~n816 & ~n834;
  assign n836 = ~n806 & ~n835;
  assign n837 = ~n815 & n824;
  assign n838 = n830 & n837;
  assign n839 = ~n836 & n838;
  assign n840 = ~n817 & n839;
  assign n841 = ~n815 & ~n817;
  assign n842 = n824 & n841;
  assign n843 = n830 & n842;
  assign n844 = ~n836 & n843;
  assign n845 = ~n808 & n4697;
  assign n846 = pi35  & ~pi163 ;
  assign n847 = pi32  & ~pi160 ;
  assign n848 = ~pi160  & ~n815;
  assign n849 = pi32  & n848;
  assign n850 = ~n815 & n847;
  assign n851 = pi33  & ~pi161 ;
  assign n852 = pi34  & ~pi162 ;
  assign n853 = ~n851 & ~n852;
  assign n854 = ~n4699 & ~n851;
  assign n855 = ~n852 & n854;
  assign n856 = ~n4699 & n853;
  assign n857 = n824 & ~n4700;
  assign n858 = ~n846 & ~n857;
  assign n859 = n830 & ~n858;
  assign n860 = pi36  & ~pi164 ;
  assign n861 = pi36  & n811;
  assign n862 = ~n809 & n860;
  assign n863 = pi37  & ~pi165 ;
  assign n864 = ~n4701 & ~n863;
  assign n865 = n827 & ~n864;
  assign n866 = pi39  & ~pi167 ;
  assign n867 = pi38  & ~pi166 ;
  assign n868 = ~pi166  & ~n825;
  assign n869 = pi38  & n868;
  assign n870 = ~n825 & n867;
  assign n871 = ~n866 & ~n4702;
  assign n872 = ~n863 & ~n867;
  assign n873 = ~n4701 & n872;
  assign n874 = n827 & ~n873;
  assign n875 = ~n866 & ~n874;
  assign n876 = ~n865 & n871;
  assign n877 = ~n4695 & ~n858;
  assign n878 = n873 & ~n877;
  assign n879 = ~n859 & ~n4702;
  assign n880 = ~n865 & n879;
  assign n881 = n827 & ~n878;
  assign n882 = ~n866 & n4704;
  assign n883 = ~n859 & n4703;
  assign n884 = ~n4698 & n4705;
  assign n885 = ~pi45  & pi173 ;
  assign n886 = ~pi44  & pi172 ;
  assign n887 = ~pi172  & ~n885;
  assign n888 = pi44  & ~n885;
  assign n889 = ~n887 & ~n888;
  assign n890 = ~n885 & ~n886;
  assign n891 = ~pi47  & pi175 ;
  assign n892 = ~pi46  & pi174 ;
  assign n893 = ~n891 & ~n892;
  assign n894 = ~n4706 & n893;
  assign n895 = ~pi43  & pi171 ;
  assign n896 = ~pi42  & pi170 ;
  assign n897 = ~n895 & ~n896;
  assign n898 = ~pi40  & pi168 ;
  assign n899 = ~pi41  & pi169 ;
  assign n900 = ~n898 & ~n899;
  assign n901 = n897 & n900;
  assign n902 = n893 & n900;
  assign n903 = n897 & n902;
  assign n904 = ~n4706 & n903;
  assign n905 = n894 & n901;
  assign n906 = ~n884 & n4707;
  assign n907 = pi43  & ~pi171 ;
  assign n908 = pi40  & ~pi168 ;
  assign n909 = ~n899 & n908;
  assign n910 = pi41  & ~pi169 ;
  assign n911 = pi42  & ~pi170 ;
  assign n912 = ~n910 & ~n911;
  assign n913 = ~n909 & ~n910;
  assign n914 = ~n911 & n913;
  assign n915 = ~n909 & n912;
  assign n916 = n897 & ~n4708;
  assign n917 = ~n907 & ~n916;
  assign n918 = n894 & ~n917;
  assign n919 = pi44  & ~pi172 ;
  assign n920 = pi44  & n887;
  assign n921 = ~n885 & n919;
  assign n922 = pi45  & ~pi173 ;
  assign n923 = ~n4709 & ~n922;
  assign n924 = n893 & ~n923;
  assign n925 = pi47  & ~pi175 ;
  assign n926 = pi46  & ~pi174 ;
  assign n927 = ~pi174  & ~n891;
  assign n928 = pi46  & n927;
  assign n929 = ~n891 & n926;
  assign n930 = ~n925 & ~n4710;
  assign n931 = ~n922 & ~n926;
  assign n932 = ~n4709 & n931;
  assign n933 = n893 & ~n932;
  assign n934 = ~n925 & ~n933;
  assign n935 = ~n924 & n930;
  assign n936 = ~n4706 & ~n917;
  assign n937 = n932 & ~n936;
  assign n938 = n893 & ~n937;
  assign n939 = ~n925 & ~n938;
  assign n940 = ~n918 & n4711;
  assign n941 = ~n906 & ~n4710;
  assign n942 = ~n924 & n941;
  assign n943 = ~n918 & n942;
  assign n944 = ~n925 & n943;
  assign n945 = ~n906 & n4712;
  assign n946 = ~pi53  & pi181 ;
  assign n947 = ~pi52  & pi180 ;
  assign n948 = ~pi180  & ~n946;
  assign n949 = pi52  & ~n946;
  assign n950 = ~n948 & ~n949;
  assign n951 = ~n946 & ~n947;
  assign n952 = ~pi55  & pi183 ;
  assign n953 = ~pi54  & pi182 ;
  assign n954 = ~n952 & ~n953;
  assign n955 = ~n4714 & n954;
  assign n956 = ~pi51  & pi179 ;
  assign n957 = ~pi50  & pi178 ;
  assign n958 = ~n956 & ~n957;
  assign n959 = ~pi49  & pi177 ;
  assign n960 = ~pi48  & pi176 ;
  assign n961 = ~n959 & ~n960;
  assign n962 = n958 & n961;
  assign n963 = n954 & n961;
  assign n964 = n958 & n963;
  assign n965 = ~n4714 & n964;
  assign n966 = n958 & ~n959;
  assign n967 = n955 & n966;
  assign n968 = ~n960 & n967;
  assign n969 = n955 & n962;
  assign n970 = ~n4713 & n4715;
  assign n971 = pi51  & ~pi179 ;
  assign n972 = pi48  & ~pi176 ;
  assign n973 = ~pi176  & ~n959;
  assign n974 = pi48  & n973;
  assign n975 = ~n959 & n972;
  assign n976 = pi49  & ~pi177 ;
  assign n977 = pi50  & ~pi178 ;
  assign n978 = ~n976 & ~n977;
  assign n979 = ~n4716 & ~n976;
  assign n980 = ~n977 & n979;
  assign n981 = ~n4716 & n978;
  assign n982 = n958 & ~n4717;
  assign n983 = ~n971 & ~n982;
  assign n984 = n955 & ~n983;
  assign n985 = pi55  & ~pi183 ;
  assign n986 = pi52  & ~pi180 ;
  assign n987 = pi52  & n948;
  assign n988 = ~n946 & n986;
  assign n989 = pi53  & ~pi181 ;
  assign n990 = pi54  & ~pi182 ;
  assign n991 = ~n989 & ~n990;
  assign n992 = ~n4718 & ~n989;
  assign n993 = ~n990 & n992;
  assign n994 = ~n4718 & n991;
  assign n995 = n954 & ~n4719;
  assign n996 = ~n985 & ~n995;
  assign n997 = ~n4714 & ~n983;
  assign n998 = n4719 & ~n997;
  assign n999 = n954 & ~n998;
  assign n1000 = ~n984 & ~n995;
  assign n1001 = ~n985 & ~n4720;
  assign n1002 = ~n984 & n996;
  assign n1003 = ~n970 & n4721;
  assign n1004 = ~pi61  & pi189 ;
  assign n1005 = ~pi60  & pi188 ;
  assign n1006 = ~pi188  & ~n1004;
  assign n1007 = pi60  & ~n1004;
  assign n1008 = ~n1006 & ~n1007;
  assign n1009 = ~n1004 & ~n1005;
  assign n1010 = ~pi63  & pi191 ;
  assign n1011 = ~pi62  & pi190 ;
  assign n1012 = ~n1010 & ~n1011;
  assign n1013 = ~n4722 & n1012;
  assign n1014 = ~pi59  & pi187 ;
  assign n1015 = ~pi58  & pi186 ;
  assign n1016 = ~n1014 & ~n1015;
  assign n1017 = ~pi56  & pi184 ;
  assign n1018 = ~pi57  & pi185 ;
  assign n1019 = ~n1017 & ~n1018;
  assign n1020 = n1016 & n1019;
  assign n1021 = n1012 & n1019;
  assign n1022 = n1016 & n1021;
  assign n1023 = ~n4722 & n1022;
  assign n1024 = n1013 & n1019;
  assign n1025 = n1016 & n1024;
  assign n1026 = n1013 & n1020;
  assign n1027 = ~n1003 & n4723;
  assign n1028 = pi59  & ~pi187 ;
  assign n1029 = pi56  & ~pi184 ;
  assign n1030 = ~n1018 & n1029;
  assign n1031 = pi57  & ~pi185 ;
  assign n1032 = pi58  & ~pi186 ;
  assign n1033 = ~n1031 & ~n1032;
  assign n1034 = ~n1030 & ~n1031;
  assign n1035 = ~n1032 & n1034;
  assign n1036 = ~n1030 & n1033;
  assign n1037 = n1016 & ~n4724;
  assign n1038 = ~n1028 & ~n1037;
  assign n1039 = n1013 & ~n1038;
  assign n1040 = pi60  & ~pi188 ;
  assign n1041 = pi60  & n1006;
  assign n1042 = ~n1004 & n1040;
  assign n1043 = pi61  & ~pi189 ;
  assign n1044 = ~n4725 & ~n1043;
  assign n1045 = n1012 & ~n1044;
  assign n1046 = pi63  & ~pi191 ;
  assign n1047 = pi62  & ~pi190 ;
  assign n1048 = ~pi190  & ~n1010;
  assign n1049 = pi62  & n1048;
  assign n1050 = ~n1010 & n1047;
  assign n1051 = ~n1046 & ~n4726;
  assign n1052 = ~n1043 & ~n1047;
  assign n1053 = ~n4725 & n1052;
  assign n1054 = n1012 & ~n1053;
  assign n1055 = ~n1046 & ~n1054;
  assign n1056 = ~n1045 & n1051;
  assign n1057 = ~n4722 & ~n1038;
  assign n1058 = n1053 & ~n1057;
  assign n1059 = n1012 & ~n1058;
  assign n1060 = ~n1046 & ~n1059;
  assign n1061 = ~n1039 & n4727;
  assign n1062 = ~n1027 & ~n4726;
  assign n1063 = ~n1045 & n1062;
  assign n1064 = ~n1039 & n1063;
  assign n1065 = ~n1046 & n1064;
  assign n1066 = ~n1027 & n4728;
  assign n1067 = ~pi67  & pi195 ;
  assign n1068 = ~pi66  & pi194 ;
  assign n1069 = ~n1067 & ~n1068;
  assign n1070 = ~pi65  & pi193 ;
  assign n1071 = ~pi64  & pi192 ;
  assign n1072 = ~n1070 & ~n1071;
  assign n1073 = n1069 & n1072;
  assign n1074 = ~n4729 & ~n1071;
  assign n1075 = ~n1070 & n1074;
  assign n1076 = n1069 & n1075;
  assign n1077 = ~n4729 & n1073;
  assign n1078 = pi67  & ~pi195 ;
  assign n1079 = pi64  & ~pi192 ;
  assign n1080 = ~n1070 & n1079;
  assign n1081 = pi65  & ~pi193 ;
  assign n1082 = pi66  & ~pi194 ;
  assign n1083 = ~n1081 & ~n1082;
  assign n1084 = ~n1080 & ~n1081;
  assign n1085 = ~n1082 & n1084;
  assign n1086 = ~n1080 & n1083;
  assign n1087 = n1069 & ~n4731;
  assign n1088 = ~n1078 & ~n1087;
  assign n1089 = ~n4730 & n1088;
  assign n1090 = ~pi71  & pi199 ;
  assign n1091 = ~pi70  & pi198 ;
  assign n1092 = ~n1090 & ~n1091;
  assign n1093 = ~pi69  & pi197 ;
  assign n1094 = ~pi68  & pi196 ;
  assign n1095 = ~n1093 & ~n1094;
  assign n1096 = n1092 & n1095;
  assign n1097 = ~n1089 & n1096;
  assign n1098 = pi71  & ~pi199 ;
  assign n1099 = pi68  & ~pi196 ;
  assign n1100 = ~n1093 & n1099;
  assign n1101 = pi70  & ~pi198 ;
  assign n1102 = pi69  & ~pi197 ;
  assign n1103 = ~n1101 & ~n1102;
  assign n1104 = ~n1100 & n1103;
  assign n1105 = n1092 & ~n1104;
  assign n1106 = ~n1100 & ~n1102;
  assign n1107 = n1092 & ~n1106;
  assign n1108 = ~pi198  & ~n1090;
  assign n1109 = pi70  & n1108;
  assign n1110 = ~n1090 & n1101;
  assign n1111 = ~n1098 & ~n4732;
  assign n1112 = ~n1107 & n1111;
  assign n1113 = ~n1098 & ~n1105;
  assign n1114 = ~n1097 & ~n4732;
  assign n1115 = ~n1107 & n1114;
  assign n1116 = ~n1098 & n1115;
  assign n1117 = ~n1097 & n4733;
  assign n1118 = ~pi75  & pi203 ;
  assign n1119 = ~pi74  & pi202 ;
  assign n1120 = ~n1118 & ~n1119;
  assign n1121 = ~pi73  & pi201 ;
  assign n1122 = ~pi72  & pi200 ;
  assign n1123 = ~n1121 & ~n1122;
  assign n1124 = n1120 & n1123;
  assign n1125 = ~n4734 & n1124;
  assign n1126 = pi75  & ~pi203 ;
  assign n1127 = pi72  & ~pi200 ;
  assign n1128 = ~n1121 & n1127;
  assign n1129 = pi73  & ~pi201 ;
  assign n1130 = pi74  & ~pi202 ;
  assign n1131 = ~n1129 & ~n1130;
  assign n1132 = ~n1128 & ~n1129;
  assign n1133 = ~n1130 & n1132;
  assign n1134 = ~n1128 & n1131;
  assign n1135 = n1120 & ~n4735;
  assign n1136 = ~n1126 & ~n1135;
  assign n1137 = ~n1125 & n1136;
  assign n1138 = ~pi79  & pi207 ;
  assign n1139 = ~pi78  & pi206 ;
  assign n1140 = ~n1138 & ~n1139;
  assign n1141 = ~pi77  & pi205 ;
  assign n1142 = ~pi76  & pi204 ;
  assign n1143 = ~n1141 & ~n1142;
  assign n1144 = n1140 & n1143;
  assign n1145 = ~n1137 & n1144;
  assign n1146 = pi79  & ~pi207 ;
  assign n1147 = pi76  & ~pi204 ;
  assign n1148 = ~n1141 & n1147;
  assign n1149 = pi78  & ~pi206 ;
  assign n1150 = pi77  & ~pi205 ;
  assign n1151 = ~n1149 & ~n1150;
  assign n1152 = ~n1148 & n1151;
  assign n1153 = n1140 & ~n1152;
  assign n1154 = ~n1148 & ~n1150;
  assign n1155 = n1140 & ~n1154;
  assign n1156 = ~pi206  & ~n1138;
  assign n1157 = pi78  & n1156;
  assign n1158 = ~n1138 & n1149;
  assign n1159 = ~n1146 & ~n4736;
  assign n1160 = ~n1155 & n1159;
  assign n1161 = ~n1146 & ~n1153;
  assign n1162 = ~n1145 & ~n4736;
  assign n1163 = ~n1155 & n1162;
  assign n1164 = ~n1146 & n1163;
  assign n1165 = ~n1145 & n4737;
  assign n1166 = ~pi83  & pi211 ;
  assign n1167 = ~pi82  & pi210 ;
  assign n1168 = ~n1166 & ~n1167;
  assign n1169 = ~pi81  & pi209 ;
  assign n1170 = ~pi80  & pi208 ;
  assign n1171 = ~n1169 & ~n1170;
  assign n1172 = n1168 & n1171;
  assign n1173 = ~n4738 & ~n1169;
  assign n1174 = n1168 & n1173;
  assign n1175 = ~n1170 & n1174;
  assign n1176 = ~n4738 & n1172;
  assign n1177 = pi83  & ~pi211 ;
  assign n1178 = pi80  & ~pi208 ;
  assign n1179 = ~pi208  & ~n1169;
  assign n1180 = pi80  & n1179;
  assign n1181 = ~n1169 & n1178;
  assign n1182 = pi81  & ~pi209 ;
  assign n1183 = pi82  & ~pi210 ;
  assign n1184 = ~n1182 & ~n1183;
  assign n1185 = ~n4740 & ~n1182;
  assign n1186 = ~n1183 & n1185;
  assign n1187 = ~n4740 & n1184;
  assign n1188 = n1168 & ~n4741;
  assign n1189 = ~n1177 & ~n1188;
  assign n1190 = ~n4739 & n1189;
  assign n1191 = ~pi87  & pi215 ;
  assign n1192 = ~pi86  & pi214 ;
  assign n1193 = ~n1191 & ~n1192;
  assign n1194 = ~pi85  & pi213 ;
  assign n1195 = ~pi84  & pi212 ;
  assign n1196 = ~n1194 & ~n1195;
  assign n1197 = n1193 & n1196;
  assign n1198 = ~n1190 & n1197;
  assign n1199 = pi87  & ~pi215 ;
  assign n1200 = pi84  & ~pi212 ;
  assign n1201 = ~n1194 & n1200;
  assign n1202 = pi86  & ~pi214 ;
  assign n1203 = pi85  & ~pi213 ;
  assign n1204 = ~n1202 & ~n1203;
  assign n1205 = ~n1201 & n1204;
  assign n1206 = n1193 & ~n1205;
  assign n1207 = ~n1201 & ~n1203;
  assign n1208 = n1193 & ~n1207;
  assign n1209 = ~pi214  & ~n1191;
  assign n1210 = pi86  & n1209;
  assign n1211 = ~n1191 & n1202;
  assign n1212 = ~n1199 & ~n4742;
  assign n1213 = ~n1208 & n1212;
  assign n1214 = ~n1199 & ~n1206;
  assign n1215 = ~n1198 & ~n4742;
  assign n1216 = ~n1208 & n1215;
  assign n1217 = ~n1199 & n1216;
  assign n1218 = ~n1198 & n4743;
  assign n1219 = ~pi91  & pi219 ;
  assign n1220 = ~pi90  & pi218 ;
  assign n1221 = ~n1219 & ~n1220;
  assign n1222 = ~pi89  & pi217 ;
  assign n1223 = ~pi88  & pi216 ;
  assign n1224 = ~n1222 & ~n1223;
  assign n1225 = n1221 & n1224;
  assign n1226 = ~n4744 & n1225;
  assign n1227 = pi91  & ~pi219 ;
  assign n1228 = pi88  & ~pi216 ;
  assign n1229 = ~n1222 & n1228;
  assign n1230 = pi89  & ~pi217 ;
  assign n1231 = pi90  & ~pi218 ;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = ~n1229 & ~n1230;
  assign n1234 = ~n1231 & n1233;
  assign n1235 = ~n1229 & n1232;
  assign n1236 = n1221 & ~n4745;
  assign n1237 = ~n1227 & ~n1236;
  assign n1238 = ~n1226 & n1237;
  assign n1239 = ~pi95  & pi223 ;
  assign n1240 = ~pi94  & pi222 ;
  assign n1241 = ~n1239 & ~n1240;
  assign n1242 = ~pi93  & pi221 ;
  assign n1243 = ~pi92  & pi220 ;
  assign n1244 = ~n1242 & ~n1243;
  assign n1245 = n1241 & n1244;
  assign n1246 = ~n1238 & n1245;
  assign n1247 = pi95  & ~pi223 ;
  assign n1248 = pi92  & ~pi220 ;
  assign n1249 = ~n1242 & n1248;
  assign n1250 = pi94  & ~pi222 ;
  assign n1251 = pi93  & ~pi221 ;
  assign n1252 = ~n1250 & ~n1251;
  assign n1253 = ~n1249 & n1252;
  assign n1254 = n1241 & ~n1253;
  assign n1255 = ~n1249 & ~n1251;
  assign n1256 = n1241 & ~n1255;
  assign n1257 = ~pi222  & ~n1239;
  assign n1258 = pi94  & n1257;
  assign n1259 = ~n1239 & n1250;
  assign n1260 = ~n1247 & ~n4746;
  assign n1261 = ~n1256 & n1260;
  assign n1262 = ~n1247 & ~n1254;
  assign n1263 = ~n1246 & ~n4746;
  assign n1264 = ~n1256 & n1263;
  assign n1265 = ~n1247 & n1264;
  assign n1266 = ~n1246 & n4747;
  assign n1267 = ~pi99  & pi227 ;
  assign n1268 = ~pi98  & pi226 ;
  assign n1269 = ~n1267 & ~n1268;
  assign n1270 = ~pi97  & pi225 ;
  assign n1271 = ~pi96  & pi224 ;
  assign n1272 = ~n1270 & ~n1271;
  assign n1273 = n1269 & n1272;
  assign n1274 = ~n4748 & ~n1270;
  assign n1275 = n1269 & n1274;
  assign n1276 = ~n1271 & n1275;
  assign n1277 = ~n4748 & n1273;
  assign n1278 = pi99  & ~pi227 ;
  assign n1279 = pi96  & ~pi224 ;
  assign n1280 = ~pi224  & ~n1270;
  assign n1281 = pi96  & n1280;
  assign n1282 = ~n1270 & n1279;
  assign n1283 = pi97  & ~pi225 ;
  assign n1284 = pi98  & ~pi226 ;
  assign n1285 = ~n1283 & ~n1284;
  assign n1286 = ~n4750 & ~n1283;
  assign n1287 = ~n1284 & n1286;
  assign n1288 = ~n4750 & n1285;
  assign n1289 = n1269 & ~n4751;
  assign n1290 = ~n1278 & ~n1289;
  assign n1291 = ~n4749 & n1290;
  assign n1292 = ~pi103  & pi231 ;
  assign n1293 = ~pi102  & pi230 ;
  assign n1294 = ~n1292 & ~n1293;
  assign n1295 = ~pi101  & pi229 ;
  assign n1296 = ~pi100  & pi228 ;
  assign n1297 = ~n1295 & ~n1296;
  assign n1298 = n1294 & n1297;
  assign n1299 = ~n1291 & n1298;
  assign n1300 = pi103  & ~pi231 ;
  assign n1301 = pi100  & ~pi228 ;
  assign n1302 = ~n1295 & n1301;
  assign n1303 = pi102  & ~pi230 ;
  assign n1304 = pi101  & ~pi229 ;
  assign n1305 = ~n1303 & ~n1304;
  assign n1306 = ~n1302 & n1305;
  assign n1307 = n1294 & ~n1306;
  assign n1308 = ~n1302 & ~n1304;
  assign n1309 = n1294 & ~n1308;
  assign n1310 = ~pi230  & ~n1292;
  assign n1311 = pi102  & n1310;
  assign n1312 = ~n1292 & n1303;
  assign n1313 = ~n1300 & ~n4752;
  assign n1314 = ~n1309 & n1313;
  assign n1315 = ~n1300 & ~n1307;
  assign n1316 = ~n1299 & ~n4752;
  assign n1317 = ~n1309 & n1316;
  assign n1318 = ~n1300 & n1317;
  assign n1319 = ~n1299 & n4753;
  assign n1320 = ~pi107  & pi235 ;
  assign n1321 = ~pi106  & pi234 ;
  assign n1322 = ~n1320 & ~n1321;
  assign n1323 = ~pi105  & pi233 ;
  assign n1324 = ~pi104  & pi232 ;
  assign n1325 = ~n1323 & ~n1324;
  assign n1326 = n1322 & n1325;
  assign n1327 = ~n4754 & n1326;
  assign n1328 = pi107  & ~pi235 ;
  assign n1329 = pi104  & ~pi232 ;
  assign n1330 = ~n1323 & n1329;
  assign n1331 = pi105  & ~pi233 ;
  assign n1332 = pi106  & ~pi234 ;
  assign n1333 = ~n1331 & ~n1332;
  assign n1334 = ~n1330 & ~n1331;
  assign n1335 = ~n1332 & n1334;
  assign n1336 = ~n1330 & n1333;
  assign n1337 = n1322 & ~n4755;
  assign n1338 = ~n1328 & ~n1337;
  assign n1339 = ~n1327 & n1338;
  assign n1340 = ~pi111  & pi239 ;
  assign n1341 = ~pi110  & pi238 ;
  assign n1342 = ~n1340 & ~n1341;
  assign n1343 = ~pi109  & pi237 ;
  assign n1344 = ~pi108  & pi236 ;
  assign n1345 = ~n1343 & ~n1344;
  assign n1346 = n1342 & n1345;
  assign n1347 = ~n1339 & n1346;
  assign n1348 = pi111  & ~pi239 ;
  assign n1349 = pi108  & ~pi236 ;
  assign n1350 = ~n1343 & n1349;
  assign n1351 = pi110  & ~pi238 ;
  assign n1352 = pi109  & ~pi237 ;
  assign n1353 = ~n1351 & ~n1352;
  assign n1354 = ~n1350 & n1353;
  assign n1355 = n1342 & ~n1354;
  assign n1356 = ~n1350 & ~n1352;
  assign n1357 = n1342 & ~n1356;
  assign n1358 = ~pi238  & ~n1340;
  assign n1359 = pi110  & n1358;
  assign n1360 = ~n1340 & n1351;
  assign n1361 = ~n1348 & ~n4756;
  assign n1362 = ~n1357 & n1361;
  assign n1363 = ~n1348 & ~n1355;
  assign n1364 = ~n1347 & ~n4756;
  assign n1365 = ~n1357 & n1364;
  assign n1366 = ~n1348 & n1365;
  assign n1367 = ~n1347 & n4757;
  assign n1368 = ~pi115  & pi243 ;
  assign n1369 = ~pi114  & pi242 ;
  assign n1370 = ~n1368 & ~n1369;
  assign n1371 = ~pi113  & pi241 ;
  assign n1372 = ~pi112  & pi240 ;
  assign n1373 = ~n1371 & ~n1372;
  assign n1374 = n1370 & n1373;
  assign n1375 = ~n4758 & ~n1371;
  assign n1376 = n1370 & n1375;
  assign n1377 = ~n1372 & n1376;
  assign n1378 = ~n4758 & n1374;
  assign n1379 = pi115  & ~pi243 ;
  assign n1380 = pi112  & ~pi240 ;
  assign n1381 = ~pi240  & ~n1371;
  assign n1382 = pi112  & n1381;
  assign n1383 = ~n1371 & n1380;
  assign n1384 = pi113  & ~pi241 ;
  assign n1385 = pi114  & ~pi242 ;
  assign n1386 = ~n1384 & ~n1385;
  assign n1387 = ~n4760 & ~n1384;
  assign n1388 = ~n1385 & n1387;
  assign n1389 = ~n4760 & n1386;
  assign n1390 = n1370 & ~n4761;
  assign n1391 = ~n1379 & ~n1390;
  assign n1392 = ~n4759 & n1391;
  assign n1393 = ~pi119  & pi247 ;
  assign n1394 = ~pi118  & pi246 ;
  assign n1395 = ~n1393 & ~n1394;
  assign n1396 = ~pi117  & pi245 ;
  assign n1397 = ~pi116  & pi244 ;
  assign n1398 = ~n1396 & ~n1397;
  assign n1399 = n1395 & n1398;
  assign n1400 = ~n1392 & n1399;
  assign n1401 = pi119  & ~pi247 ;
  assign n1402 = pi116  & ~pi244 ;
  assign n1403 = ~n1396 & n1402;
  assign n1404 = pi118  & ~pi246 ;
  assign n1405 = pi117  & ~pi245 ;
  assign n1406 = ~n1404 & ~n1405;
  assign n1407 = ~n1403 & n1406;
  assign n1408 = n1395 & ~n1407;
  assign n1409 = ~n1403 & ~n1405;
  assign n1410 = n1395 & ~n1409;
  assign n1411 = ~pi246  & ~n1393;
  assign n1412 = pi118  & n1411;
  assign n1413 = ~n1393 & n1404;
  assign n1414 = ~n1401 & ~n4762;
  assign n1415 = ~n1410 & n1414;
  assign n1416 = ~n1401 & ~n1408;
  assign n1417 = ~n1400 & ~n4762;
  assign n1418 = ~n1410 & n1417;
  assign n1419 = ~n1401 & n1418;
  assign n1420 = ~n1400 & n4763;
  assign n1421 = ~pi123  & pi251 ;
  assign n1422 = ~pi122  & pi250 ;
  assign n1423 = ~n1421 & ~n1422;
  assign n1424 = ~pi121  & pi249 ;
  assign n1425 = ~pi120  & pi248 ;
  assign n1426 = ~n1424 & ~n1425;
  assign n1427 = n1423 & n1426;
  assign n1428 = ~n4764 & n1427;
  assign n1429 = pi123  & ~pi251 ;
  assign n1430 = pi120  & ~pi248 ;
  assign n1431 = ~n1424 & n1430;
  assign n1432 = pi121  & ~pi249 ;
  assign n1433 = pi122  & ~pi250 ;
  assign n1434 = ~n1432 & ~n1433;
  assign n1435 = ~n1431 & ~n1432;
  assign n1436 = ~n1433 & n1435;
  assign n1437 = ~n1431 & n1434;
  assign n1438 = n1423 & ~n4765;
  assign n1439 = ~n1429 & ~n1438;
  assign n1440 = ~n1428 & n1439;
  assign n1441 = ~pi126  & pi254 ;
  assign n1442 = ~pi125  & pi253 ;
  assign n1443 = ~n1441 & ~n1442;
  assign n1444 = pi127  & ~pi255 ;
  assign n1445 = ~pi124  & pi252 ;
  assign n1446 = ~n1444 & ~n1445;
  assign n1447 = n1443 & ~n1444;
  assign n1448 = ~n1445 & n1447;
  assign n1449 = n1443 & n1446;
  assign n1450 = ~n1440 & n4766;
  assign n1451 = pi124  & ~pi252 ;
  assign n1452 = pi125  & ~pi253 ;
  assign n1453 = ~n1451 & ~n1452;
  assign n1454 = n1443 & ~n1453;
  assign n1455 = pi126  & ~pi254 ;
  assign n1456 = ~n1454 & ~n1455;
  assign n1457 = ~n1444 & ~n1456;
  assign n1458 = ~pi127  & pi255 ;
  assign n1459 = ~n1457 & ~n1458;
  assign n1460 = ~n1450 & ~n1457;
  assign n1461 = ~n1458 & n1460;
  assign n1462 = ~n1450 & n1459;
  assign n1463 = pi28  & ~n4767;
  assign n1464 = pi156  & n4767;
  assign n1465 = ~n1463 & ~n1464;
  assign n1466 = ~pi282  & pi410 ;
  assign n1467 = pi281  & ~pi409 ;
  assign n1468 = ~pi281  & pi409 ;
  assign n1469 = pi280  & ~pi408 ;
  assign n1470 = ~pi280  & pi408 ;
  assign n1471 = pi279  & ~pi407 ;
  assign n1472 = ~pi279  & pi407 ;
  assign n1473 = pi278  & ~pi406 ;
  assign n1474 = ~pi278  & pi406 ;
  assign n1475 = pi277  & ~pi405 ;
  assign n1476 = ~pi277  & pi405 ;
  assign n1477 = pi276  & ~pi404 ;
  assign n1478 = ~pi276  & pi404 ;
  assign n1479 = pi275  & ~pi403 ;
  assign n1480 = ~pi275  & pi403 ;
  assign n1481 = pi274  & ~pi402 ;
  assign n1482 = ~pi274  & pi402 ;
  assign n1483 = pi273  & ~pi401 ;
  assign n1484 = ~pi273  & pi401 ;
  assign n1485 = pi272  & ~pi400 ;
  assign n1486 = ~pi272  & pi400 ;
  assign n1487 = pi271  & ~pi399 ;
  assign n1488 = ~pi271  & pi399 ;
  assign n1489 = pi270  & ~pi398 ;
  assign n1490 = ~pi270  & pi398 ;
  assign n1491 = pi269  & ~pi397 ;
  assign n1492 = ~pi269  & pi397 ;
  assign n1493 = pi268  & ~pi396 ;
  assign n1494 = ~pi268  & pi396 ;
  assign n1495 = pi267  & ~pi395 ;
  assign n1496 = ~pi267  & pi395 ;
  assign n1497 = pi266  & ~pi394 ;
  assign n1498 = ~pi266  & pi394 ;
  assign n1499 = pi265  & ~pi393 ;
  assign n1500 = ~pi265  & pi393 ;
  assign n1501 = pi264  & ~pi392 ;
  assign n1502 = ~pi264  & pi392 ;
  assign n1503 = pi263  & ~pi391 ;
  assign n1504 = ~pi263  & pi391 ;
  assign n1505 = pi262  & ~pi390 ;
  assign n1506 = ~pi262  & pi390 ;
  assign n1507 = pi261  & ~pi389 ;
  assign n1508 = ~pi261  & pi389 ;
  assign n1509 = pi260  & ~pi388 ;
  assign n1510 = ~pi260  & pi388 ;
  assign n1511 = pi259  & ~pi387 ;
  assign n1512 = ~pi259  & pi387 ;
  assign n1513 = pi258  & ~pi386 ;
  assign n1514 = ~pi258  & pi386 ;
  assign n1515 = pi257  & ~pi385 ;
  assign n1516 = ~pi257  & pi385 ;
  assign n1517 = pi256  & ~pi384 ;
  assign n1518 = ~n1516 & n1517;
  assign n1519 = ~n1515 & ~n1518;
  assign n1520 = pi257  & n1517;
  assign n1521 = pi385  & ~n1520;
  assign n1522 = ~pi257  & ~n1517;
  assign n1523 = ~n1514 & ~n1522;
  assign n1524 = ~n1521 & n1523;
  assign n1525 = ~n1514 & ~n1519;
  assign n1526 = ~n1513 & ~n4768;
  assign n1527 = ~n1512 & ~n1526;
  assign n1528 = ~n1511 & ~n1527;
  assign n1529 = ~n1510 & ~n1528;
  assign n1530 = ~pi260  & n1528;
  assign n1531 = ~pi388  & ~n1530;
  assign n1532 = pi260  & ~n1528;
  assign n1533 = ~n1531 & ~n1532;
  assign n1534 = ~n1509 & ~n1529;
  assign n1535 = ~n1508 & ~n4769;
  assign n1536 = ~pi261  & n4769;
  assign n1537 = ~pi389  & ~n1536;
  assign n1538 = pi261  & ~n4769;
  assign n1539 = ~n1537 & ~n1538;
  assign n1540 = ~n1507 & ~n1535;
  assign n1541 = ~n1506 & ~n4770;
  assign n1542 = ~n1505 & ~n1541;
  assign n1543 = ~n1504 & ~n1542;
  assign n1544 = ~n1503 & ~n1543;
  assign n1545 = ~n1502 & ~n1544;
  assign n1546 = ~pi264  & n1544;
  assign n1547 = ~pi392  & ~n1546;
  assign n1548 = pi264  & ~n1544;
  assign n1549 = ~n1547 & ~n1548;
  assign n1550 = ~n1501 & ~n1545;
  assign n1551 = ~n1500 & ~n4771;
  assign n1552 = ~pi265  & n4771;
  assign n1553 = ~pi393  & ~n1552;
  assign n1554 = pi265  & ~n4771;
  assign n1555 = ~n1553 & ~n1554;
  assign n1556 = ~n1499 & ~n1551;
  assign n1557 = ~n1498 & ~n4772;
  assign n1558 = ~n1497 & ~n1557;
  assign n1559 = ~n1496 & ~n1558;
  assign n1560 = ~n1495 & ~n1559;
  assign n1561 = ~n1494 & ~n1560;
  assign n1562 = ~n1493 & ~n1561;
  assign n1563 = ~n1492 & ~n1562;
  assign n1564 = ~n1491 & ~n1563;
  assign n1565 = ~n1490 & ~n1564;
  assign n1566 = ~n1489 & ~n1565;
  assign n1567 = ~n1488 & ~n1566;
  assign n1568 = ~n1487 & ~n1567;
  assign n1569 = ~n1486 & ~n1568;
  assign n1570 = ~pi272  & n1568;
  assign n1571 = ~pi400  & ~n1570;
  assign n1572 = pi272  & ~n1568;
  assign n1573 = ~n1571 & ~n1572;
  assign n1574 = ~n1485 & ~n1569;
  assign n1575 = ~n1484 & ~n4773;
  assign n1576 = ~pi273  & n4773;
  assign n1577 = ~pi401  & ~n1576;
  assign n1578 = pi273  & ~n4773;
  assign n1579 = ~n1577 & ~n1578;
  assign n1580 = ~n1483 & ~n1575;
  assign n1581 = ~n1482 & ~n4774;
  assign n1582 = ~n1481 & ~n1581;
  assign n1583 = ~n1480 & ~n1582;
  assign n1584 = ~n1479 & ~n1583;
  assign n1585 = ~n1478 & ~n1584;
  assign n1586 = ~n1477 & ~n1585;
  assign n1587 = ~n1476 & ~n1586;
  assign n1588 = ~n1475 & ~n1587;
  assign n1589 = ~n1474 & ~n1588;
  assign n1590 = ~n1473 & ~n1589;
  assign n1591 = ~n1472 & ~n1590;
  assign n1592 = ~n1471 & ~n1591;
  assign n1593 = ~n1470 & ~n1592;
  assign n1594 = ~pi280  & n1592;
  assign n1595 = ~pi408  & ~n1594;
  assign n1596 = pi280  & ~n1592;
  assign n1597 = ~n1595 & ~n1596;
  assign n1598 = ~n1469 & ~n1593;
  assign n1599 = ~n1468 & ~n4775;
  assign n1600 = ~pi281  & n4775;
  assign n1601 = ~pi409  & ~n1600;
  assign n1602 = pi281  & ~n4775;
  assign n1603 = ~n1601 & ~n1602;
  assign n1604 = ~n1467 & ~n1599;
  assign n1605 = ~n1466 & ~n4776;
  assign n1606 = pi282  & ~pi410 ;
  assign n1607 = pi283  & ~pi411 ;
  assign n1608 = ~n1606 & ~n1607;
  assign n1609 = ~n1605 & n1608;
  assign n1610 = ~pi283  & pi411 ;
  assign n1611 = ~pi284  & pi412 ;
  assign n1612 = ~n1610 & ~n1611;
  assign n1613 = ~n1605 & ~n1606;
  assign n1614 = ~n1610 & ~n1613;
  assign n1615 = ~n1607 & ~n1614;
  assign n1616 = ~n1611 & ~n1615;
  assign n1617 = ~n1609 & n1612;
  assign n1618 = pi284  & ~pi412 ;
  assign n1619 = pi285  & ~pi413 ;
  assign n1620 = ~n1618 & ~n1619;
  assign n1621 = ~n4777 & n1620;
  assign n1622 = ~pi285  & pi413 ;
  assign n1623 = ~pi286  & pi414 ;
  assign n1624 = ~n1622 & ~n1623;
  assign n1625 = ~n4777 & ~n1618;
  assign n1626 = ~n1622 & ~n1625;
  assign n1627 = ~n1619 & ~n1626;
  assign n1628 = ~n1623 & ~n1627;
  assign n1629 = ~n1621 & n1624;
  assign n1630 = pi286  & ~pi414 ;
  assign n1631 = pi287  & ~pi415 ;
  assign n1632 = ~n1630 & ~n1631;
  assign n1633 = ~n4778 & n1632;
  assign n1634 = ~pi293  & pi421 ;
  assign n1635 = ~pi292  & pi420 ;
  assign n1636 = ~pi420  & ~n1634;
  assign n1637 = pi292  & ~n1634;
  assign n1638 = ~n1636 & ~n1637;
  assign n1639 = ~n1634 & ~n1635;
  assign n1640 = ~pi289  & pi417 ;
  assign n1641 = ~pi287  & pi415 ;
  assign n1642 = ~pi288  & pi416 ;
  assign n1643 = ~n1641 & ~n1642;
  assign n1644 = ~n1640 & ~n1641;
  assign n1645 = ~n1642 & n1644;
  assign n1646 = ~n1640 & n1643;
  assign n1647 = ~pi291  & pi419 ;
  assign n1648 = ~pi290  & pi418 ;
  assign n1649 = ~n1647 & ~n1648;
  assign n1650 = ~pi295  & pi423 ;
  assign n1651 = ~pi294  & pi422 ;
  assign n1652 = ~n1650 & ~n1651;
  assign n1653 = n1649 & n1652;
  assign n1654 = n4780 & n1653;
  assign n1655 = ~n4779 & n1652;
  assign n1656 = n4780 & n1649;
  assign n1657 = n1655 & n1656;
  assign n1658 = ~n4779 & n1654;
  assign n1659 = ~n4778 & ~n1630;
  assign n1660 = ~n1641 & ~n1659;
  assign n1661 = ~n1631 & ~n1660;
  assign n1662 = ~n1640 & n1649;
  assign n1663 = n1655 & n1662;
  assign n1664 = ~n1661 & n1663;
  assign n1665 = ~n1642 & n1664;
  assign n1666 = ~n1640 & ~n1642;
  assign n1667 = n1649 & n1666;
  assign n1668 = n1655 & n1667;
  assign n1669 = ~n1661 & n1668;
  assign n1670 = ~n1633 & n4781;
  assign n1671 = pi291  & ~pi419 ;
  assign n1672 = pi288  & ~pi416 ;
  assign n1673 = ~pi416  & ~n1640;
  assign n1674 = pi288  & n1673;
  assign n1675 = ~n1640 & n1672;
  assign n1676 = pi289  & ~pi417 ;
  assign n1677 = pi290  & ~pi418 ;
  assign n1678 = ~n1676 & ~n1677;
  assign n1679 = ~n4783 & ~n1676;
  assign n1680 = ~n1677 & n1679;
  assign n1681 = ~n4783 & n1678;
  assign n1682 = n1649 & ~n4784;
  assign n1683 = ~n1671 & ~n1682;
  assign n1684 = n1655 & ~n1683;
  assign n1685 = pi292  & ~pi420 ;
  assign n1686 = pi292  & n1636;
  assign n1687 = ~n1634 & n1685;
  assign n1688 = pi293  & ~pi421 ;
  assign n1689 = ~n4785 & ~n1688;
  assign n1690 = n1652 & ~n1689;
  assign n1691 = pi295  & ~pi423 ;
  assign n1692 = pi294  & ~pi422 ;
  assign n1693 = ~pi422  & ~n1650;
  assign n1694 = pi294  & n1693;
  assign n1695 = ~n1650 & n1692;
  assign n1696 = ~n1691 & ~n4786;
  assign n1697 = ~n1688 & ~n1692;
  assign n1698 = ~n4785 & n1697;
  assign n1699 = n1652 & ~n1698;
  assign n1700 = ~n1691 & ~n1699;
  assign n1701 = ~n1690 & n1696;
  assign n1702 = ~n4779 & ~n1683;
  assign n1703 = n1698 & ~n1702;
  assign n1704 = ~n1684 & ~n4786;
  assign n1705 = ~n1690 & n1704;
  assign n1706 = n1652 & ~n1703;
  assign n1707 = ~n1691 & n4788;
  assign n1708 = ~n1684 & n4787;
  assign n1709 = ~n4782 & n4789;
  assign n1710 = ~pi301  & pi429 ;
  assign n1711 = ~pi300  & pi428 ;
  assign n1712 = ~pi428  & ~n1710;
  assign n1713 = pi300  & ~n1710;
  assign n1714 = ~n1712 & ~n1713;
  assign n1715 = ~n1710 & ~n1711;
  assign n1716 = ~pi303  & pi431 ;
  assign n1717 = ~pi302  & pi430 ;
  assign n1718 = ~n1716 & ~n1717;
  assign n1719 = ~n4790 & n1718;
  assign n1720 = ~pi299  & pi427 ;
  assign n1721 = ~pi298  & pi426 ;
  assign n1722 = ~n1720 & ~n1721;
  assign n1723 = ~pi296  & pi424 ;
  assign n1724 = ~pi297  & pi425 ;
  assign n1725 = ~n1723 & ~n1724;
  assign n1726 = n1722 & n1725;
  assign n1727 = n1718 & n1725;
  assign n1728 = n1722 & n1727;
  assign n1729 = ~n4790 & n1728;
  assign n1730 = n1719 & n1726;
  assign n1731 = ~n1709 & n4791;
  assign n1732 = pi299  & ~pi427 ;
  assign n1733 = pi296  & ~pi424 ;
  assign n1734 = ~n1724 & n1733;
  assign n1735 = pi297  & ~pi425 ;
  assign n1736 = pi298  & ~pi426 ;
  assign n1737 = ~n1735 & ~n1736;
  assign n1738 = ~n1734 & ~n1735;
  assign n1739 = ~n1736 & n1738;
  assign n1740 = ~n1734 & n1737;
  assign n1741 = n1722 & ~n4792;
  assign n1742 = ~n1732 & ~n1741;
  assign n1743 = n1719 & ~n1742;
  assign n1744 = pi300  & ~pi428 ;
  assign n1745 = pi300  & n1712;
  assign n1746 = ~n1710 & n1744;
  assign n1747 = pi301  & ~pi429 ;
  assign n1748 = ~n4793 & ~n1747;
  assign n1749 = n1718 & ~n1748;
  assign n1750 = pi303  & ~pi431 ;
  assign n1751 = pi302  & ~pi430 ;
  assign n1752 = ~pi430  & ~n1716;
  assign n1753 = pi302  & n1752;
  assign n1754 = ~n1716 & n1751;
  assign n1755 = ~n1750 & ~n4794;
  assign n1756 = ~n1747 & ~n1751;
  assign n1757 = ~n4793 & n1756;
  assign n1758 = n1718 & ~n1757;
  assign n1759 = ~n1750 & ~n1758;
  assign n1760 = ~n1749 & n1755;
  assign n1761 = ~n4790 & ~n1742;
  assign n1762 = n1757 & ~n1761;
  assign n1763 = n1718 & ~n1762;
  assign n1764 = ~n1750 & ~n1763;
  assign n1765 = ~n1743 & n4795;
  assign n1766 = ~n1731 & ~n4794;
  assign n1767 = ~n1749 & n1766;
  assign n1768 = ~n1743 & n1767;
  assign n1769 = ~n1750 & n1768;
  assign n1770 = ~n1731 & n4796;
  assign n1771 = ~pi309  & pi437 ;
  assign n1772 = ~pi308  & pi436 ;
  assign n1773 = ~pi436  & ~n1771;
  assign n1774 = pi308  & ~n1771;
  assign n1775 = ~n1773 & ~n1774;
  assign n1776 = ~n1771 & ~n1772;
  assign n1777 = ~pi311  & pi439 ;
  assign n1778 = ~pi310  & pi438 ;
  assign n1779 = ~n1777 & ~n1778;
  assign n1780 = ~n4798 & n1779;
  assign n1781 = ~pi307  & pi435 ;
  assign n1782 = ~pi306  & pi434 ;
  assign n1783 = ~n1781 & ~n1782;
  assign n1784 = ~pi305  & pi433 ;
  assign n1785 = ~pi304  & pi432 ;
  assign n1786 = ~n1784 & ~n1785;
  assign n1787 = n1783 & n1786;
  assign n1788 = n1779 & n1786;
  assign n1789 = n1783 & n1788;
  assign n1790 = ~n4798 & n1789;
  assign n1791 = n1783 & ~n1784;
  assign n1792 = n1780 & n1791;
  assign n1793 = ~n1785 & n1792;
  assign n1794 = n1780 & n1787;
  assign n1795 = ~n4797 & n4799;
  assign n1796 = pi307  & ~pi435 ;
  assign n1797 = pi304  & ~pi432 ;
  assign n1798 = ~pi432  & ~n1784;
  assign n1799 = pi304  & n1798;
  assign n1800 = ~n1784 & n1797;
  assign n1801 = pi305  & ~pi433 ;
  assign n1802 = pi306  & ~pi434 ;
  assign n1803 = ~n1801 & ~n1802;
  assign n1804 = ~n4800 & ~n1801;
  assign n1805 = ~n1802 & n1804;
  assign n1806 = ~n4800 & n1803;
  assign n1807 = n1783 & ~n4801;
  assign n1808 = ~n1796 & ~n1807;
  assign n1809 = n1780 & ~n1808;
  assign n1810 = pi311  & ~pi439 ;
  assign n1811 = pi308  & ~pi436 ;
  assign n1812 = pi308  & n1773;
  assign n1813 = ~n1771 & n1811;
  assign n1814 = pi309  & ~pi437 ;
  assign n1815 = pi310  & ~pi438 ;
  assign n1816 = ~n1814 & ~n1815;
  assign n1817 = ~n4802 & ~n1814;
  assign n1818 = ~n1815 & n1817;
  assign n1819 = ~n4802 & n1816;
  assign n1820 = n1779 & ~n4803;
  assign n1821 = ~n1810 & ~n1820;
  assign n1822 = ~n4798 & ~n1808;
  assign n1823 = n4803 & ~n1822;
  assign n1824 = n1779 & ~n1823;
  assign n1825 = ~n1809 & ~n1820;
  assign n1826 = ~n1810 & ~n4804;
  assign n1827 = ~n1809 & n1821;
  assign n1828 = ~n1795 & n4805;
  assign n1829 = ~pi317  & pi445 ;
  assign n1830 = ~pi316  & pi444 ;
  assign n1831 = ~pi444  & ~n1829;
  assign n1832 = pi316  & ~n1829;
  assign n1833 = ~n1831 & ~n1832;
  assign n1834 = ~n1829 & ~n1830;
  assign n1835 = ~pi319  & pi447 ;
  assign n1836 = ~pi318  & pi446 ;
  assign n1837 = ~n1835 & ~n1836;
  assign n1838 = ~n4806 & n1837;
  assign n1839 = ~pi315  & pi443 ;
  assign n1840 = ~pi314  & pi442 ;
  assign n1841 = ~n1839 & ~n1840;
  assign n1842 = ~pi312  & pi440 ;
  assign n1843 = ~pi313  & pi441 ;
  assign n1844 = ~n1842 & ~n1843;
  assign n1845 = n1841 & n1844;
  assign n1846 = n1837 & n1844;
  assign n1847 = n1841 & n1846;
  assign n1848 = ~n4806 & n1847;
  assign n1849 = n1838 & n1844;
  assign n1850 = n1841 & n1849;
  assign n1851 = n1838 & n1845;
  assign n1852 = ~n1828 & n4807;
  assign n1853 = pi315  & ~pi443 ;
  assign n1854 = pi312  & ~pi440 ;
  assign n1855 = ~n1843 & n1854;
  assign n1856 = pi313  & ~pi441 ;
  assign n1857 = pi314  & ~pi442 ;
  assign n1858 = ~n1856 & ~n1857;
  assign n1859 = ~n1855 & ~n1856;
  assign n1860 = ~n1857 & n1859;
  assign n1861 = ~n1855 & n1858;
  assign n1862 = n1841 & ~n4808;
  assign n1863 = ~n1853 & ~n1862;
  assign n1864 = n1838 & ~n1863;
  assign n1865 = pi316  & ~pi444 ;
  assign n1866 = pi316  & n1831;
  assign n1867 = ~n1829 & n1865;
  assign n1868 = pi317  & ~pi445 ;
  assign n1869 = ~n4809 & ~n1868;
  assign n1870 = n1837 & ~n1869;
  assign n1871 = pi319  & ~pi447 ;
  assign n1872 = pi318  & ~pi446 ;
  assign n1873 = ~pi446  & ~n1835;
  assign n1874 = pi318  & n1873;
  assign n1875 = ~n1835 & n1872;
  assign n1876 = ~n1871 & ~n4810;
  assign n1877 = ~n1868 & ~n1872;
  assign n1878 = ~n4809 & n1877;
  assign n1879 = n1837 & ~n1878;
  assign n1880 = ~n1871 & ~n1879;
  assign n1881 = ~n1870 & n1876;
  assign n1882 = ~n4806 & ~n1863;
  assign n1883 = n1878 & ~n1882;
  assign n1884 = n1837 & ~n1883;
  assign n1885 = ~n1871 & ~n1884;
  assign n1886 = ~n1864 & n4811;
  assign n1887 = ~n1852 & ~n4810;
  assign n1888 = ~n1870 & n1887;
  assign n1889 = ~n1864 & n1888;
  assign n1890 = ~n1871 & n1889;
  assign n1891 = ~n1852 & n4812;
  assign n1892 = ~pi323  & pi451 ;
  assign n1893 = ~pi322  & pi450 ;
  assign n1894 = ~n1892 & ~n1893;
  assign n1895 = ~pi321  & pi449 ;
  assign n1896 = ~pi320  & pi448 ;
  assign n1897 = ~n1895 & ~n1896;
  assign n1898 = n1894 & n1897;
  assign n1899 = ~n4813 & ~n1896;
  assign n1900 = ~n1895 & n1899;
  assign n1901 = n1894 & n1900;
  assign n1902 = ~n4813 & n1898;
  assign n1903 = pi323  & ~pi451 ;
  assign n1904 = pi320  & ~pi448 ;
  assign n1905 = ~n1895 & n1904;
  assign n1906 = pi321  & ~pi449 ;
  assign n1907 = pi322  & ~pi450 ;
  assign n1908 = ~n1906 & ~n1907;
  assign n1909 = ~n1905 & ~n1906;
  assign n1910 = ~n1907 & n1909;
  assign n1911 = ~n1905 & n1908;
  assign n1912 = n1894 & ~n4815;
  assign n1913 = ~n1903 & ~n1912;
  assign n1914 = ~n4814 & n1913;
  assign n1915 = ~pi327  & pi455 ;
  assign n1916 = ~pi326  & pi454 ;
  assign n1917 = ~n1915 & ~n1916;
  assign n1918 = ~pi325  & pi453 ;
  assign n1919 = ~pi324  & pi452 ;
  assign n1920 = ~n1918 & ~n1919;
  assign n1921 = n1917 & n1920;
  assign n1922 = ~n1914 & n1921;
  assign n1923 = pi327  & ~pi455 ;
  assign n1924 = pi324  & ~pi452 ;
  assign n1925 = ~n1918 & n1924;
  assign n1926 = pi326  & ~pi454 ;
  assign n1927 = pi325  & ~pi453 ;
  assign n1928 = ~n1926 & ~n1927;
  assign n1929 = ~n1925 & n1928;
  assign n1930 = n1917 & ~n1929;
  assign n1931 = ~n1925 & ~n1927;
  assign n1932 = n1917 & ~n1931;
  assign n1933 = ~pi454  & ~n1915;
  assign n1934 = pi326  & n1933;
  assign n1935 = ~n1915 & n1926;
  assign n1936 = ~n1923 & ~n4816;
  assign n1937 = ~n1932 & n1936;
  assign n1938 = ~n1923 & ~n1930;
  assign n1939 = ~n1922 & ~n4816;
  assign n1940 = ~n1932 & n1939;
  assign n1941 = ~n1923 & n1940;
  assign n1942 = ~n1922 & n4817;
  assign n1943 = ~pi331  & pi459 ;
  assign n1944 = ~pi330  & pi458 ;
  assign n1945 = ~n1943 & ~n1944;
  assign n1946 = ~pi329  & pi457 ;
  assign n1947 = ~pi328  & pi456 ;
  assign n1948 = ~n1946 & ~n1947;
  assign n1949 = n1945 & n1948;
  assign n1950 = ~n4818 & n1949;
  assign n1951 = pi331  & ~pi459 ;
  assign n1952 = pi328  & ~pi456 ;
  assign n1953 = ~n1946 & n1952;
  assign n1954 = pi329  & ~pi457 ;
  assign n1955 = pi330  & ~pi458 ;
  assign n1956 = ~n1954 & ~n1955;
  assign n1957 = ~n1953 & ~n1954;
  assign n1958 = ~n1955 & n1957;
  assign n1959 = ~n1953 & n1956;
  assign n1960 = n1945 & ~n4819;
  assign n1961 = ~n1951 & ~n1960;
  assign n1962 = ~n1950 & n1961;
  assign n1963 = ~pi335  & pi463 ;
  assign n1964 = ~pi334  & pi462 ;
  assign n1965 = ~n1963 & ~n1964;
  assign n1966 = ~pi333  & pi461 ;
  assign n1967 = ~pi332  & pi460 ;
  assign n1968 = ~n1966 & ~n1967;
  assign n1969 = n1965 & n1968;
  assign n1970 = ~n1962 & n1969;
  assign n1971 = pi335  & ~pi463 ;
  assign n1972 = pi332  & ~pi460 ;
  assign n1973 = ~n1966 & n1972;
  assign n1974 = pi334  & ~pi462 ;
  assign n1975 = pi333  & ~pi461 ;
  assign n1976 = ~n1974 & ~n1975;
  assign n1977 = ~n1973 & n1976;
  assign n1978 = n1965 & ~n1977;
  assign n1979 = ~n1973 & ~n1975;
  assign n1980 = n1965 & ~n1979;
  assign n1981 = ~pi462  & ~n1963;
  assign n1982 = pi334  & n1981;
  assign n1983 = ~n1963 & n1974;
  assign n1984 = ~n1971 & ~n4820;
  assign n1985 = ~n1980 & n1984;
  assign n1986 = ~n1971 & ~n1978;
  assign n1987 = ~n1970 & ~n4820;
  assign n1988 = ~n1980 & n1987;
  assign n1989 = ~n1971 & n1988;
  assign n1990 = ~n1970 & n4821;
  assign n1991 = ~pi339  & pi467 ;
  assign n1992 = ~pi338  & pi466 ;
  assign n1993 = ~n1991 & ~n1992;
  assign n1994 = ~pi337  & pi465 ;
  assign n1995 = ~pi336  & pi464 ;
  assign n1996 = ~n1994 & ~n1995;
  assign n1997 = n1993 & n1996;
  assign n1998 = ~n4822 & ~n1994;
  assign n1999 = n1993 & n1998;
  assign n2000 = ~n1995 & n1999;
  assign n2001 = ~n4822 & n1997;
  assign n2002 = pi339  & ~pi467 ;
  assign n2003 = pi336  & ~pi464 ;
  assign n2004 = ~pi464  & ~n1994;
  assign n2005 = pi336  & n2004;
  assign n2006 = ~n1994 & n2003;
  assign n2007 = pi337  & ~pi465 ;
  assign n2008 = pi338  & ~pi466 ;
  assign n2009 = ~n2007 & ~n2008;
  assign n2010 = ~n4824 & ~n2007;
  assign n2011 = ~n2008 & n2010;
  assign n2012 = ~n4824 & n2009;
  assign n2013 = n1993 & ~n4825;
  assign n2014 = ~n2002 & ~n2013;
  assign n2015 = ~n4823 & n2014;
  assign n2016 = ~pi343  & pi471 ;
  assign n2017 = ~pi342  & pi470 ;
  assign n2018 = ~n2016 & ~n2017;
  assign n2019 = ~pi341  & pi469 ;
  assign n2020 = ~pi340  & pi468 ;
  assign n2021 = ~n2019 & ~n2020;
  assign n2022 = n2018 & n2021;
  assign n2023 = ~n2015 & n2022;
  assign n2024 = pi343  & ~pi471 ;
  assign n2025 = pi340  & ~pi468 ;
  assign n2026 = ~n2019 & n2025;
  assign n2027 = pi342  & ~pi470 ;
  assign n2028 = pi341  & ~pi469 ;
  assign n2029 = ~n2027 & ~n2028;
  assign n2030 = ~n2026 & n2029;
  assign n2031 = n2018 & ~n2030;
  assign n2032 = ~n2026 & ~n2028;
  assign n2033 = n2018 & ~n2032;
  assign n2034 = ~pi470  & ~n2016;
  assign n2035 = pi342  & n2034;
  assign n2036 = ~n2016 & n2027;
  assign n2037 = ~n2024 & ~n4826;
  assign n2038 = ~n2033 & n2037;
  assign n2039 = ~n2024 & ~n2031;
  assign n2040 = ~n2023 & ~n4826;
  assign n2041 = ~n2033 & n2040;
  assign n2042 = ~n2024 & n2041;
  assign n2043 = ~n2023 & n4827;
  assign n2044 = ~pi347  & pi475 ;
  assign n2045 = ~pi346  & pi474 ;
  assign n2046 = ~n2044 & ~n2045;
  assign n2047 = ~pi345  & pi473 ;
  assign n2048 = ~pi344  & pi472 ;
  assign n2049 = ~n2047 & ~n2048;
  assign n2050 = n2046 & n2049;
  assign n2051 = ~n4828 & n2050;
  assign n2052 = pi347  & ~pi475 ;
  assign n2053 = pi344  & ~pi472 ;
  assign n2054 = ~n2047 & n2053;
  assign n2055 = pi345  & ~pi473 ;
  assign n2056 = pi346  & ~pi474 ;
  assign n2057 = ~n2055 & ~n2056;
  assign n2058 = ~n2054 & ~n2055;
  assign n2059 = ~n2056 & n2058;
  assign n2060 = ~n2054 & n2057;
  assign n2061 = n2046 & ~n4829;
  assign n2062 = ~n2052 & ~n2061;
  assign n2063 = ~n2051 & n2062;
  assign n2064 = ~pi351  & pi479 ;
  assign n2065 = ~pi350  & pi478 ;
  assign n2066 = ~n2064 & ~n2065;
  assign n2067 = ~pi349  & pi477 ;
  assign n2068 = ~pi348  & pi476 ;
  assign n2069 = ~n2067 & ~n2068;
  assign n2070 = n2066 & n2069;
  assign n2071 = ~n2063 & n2070;
  assign n2072 = pi351  & ~pi479 ;
  assign n2073 = pi348  & ~pi476 ;
  assign n2074 = ~n2067 & n2073;
  assign n2075 = pi350  & ~pi478 ;
  assign n2076 = pi349  & ~pi477 ;
  assign n2077 = ~n2075 & ~n2076;
  assign n2078 = ~n2074 & n2077;
  assign n2079 = n2066 & ~n2078;
  assign n2080 = ~n2074 & ~n2076;
  assign n2081 = n2066 & ~n2080;
  assign n2082 = ~pi478  & ~n2064;
  assign n2083 = pi350  & n2082;
  assign n2084 = ~n2064 & n2075;
  assign n2085 = ~n2072 & ~n4830;
  assign n2086 = ~n2081 & n2085;
  assign n2087 = ~n2072 & ~n2079;
  assign n2088 = ~n2071 & ~n4830;
  assign n2089 = ~n2081 & n2088;
  assign n2090 = ~n2072 & n2089;
  assign n2091 = ~n2071 & n4831;
  assign n2092 = ~pi355  & pi483 ;
  assign n2093 = ~pi354  & pi482 ;
  assign n2094 = ~n2092 & ~n2093;
  assign n2095 = ~pi353  & pi481 ;
  assign n2096 = ~pi352  & pi480 ;
  assign n2097 = ~n2095 & ~n2096;
  assign n2098 = n2094 & n2097;
  assign n2099 = ~n4832 & ~n2095;
  assign n2100 = n2094 & n2099;
  assign n2101 = ~n2096 & n2100;
  assign n2102 = ~n4832 & n2098;
  assign n2103 = pi355  & ~pi483 ;
  assign n2104 = pi352  & ~pi480 ;
  assign n2105 = ~pi480  & ~n2095;
  assign n2106 = pi352  & n2105;
  assign n2107 = ~n2095 & n2104;
  assign n2108 = pi353  & ~pi481 ;
  assign n2109 = pi354  & ~pi482 ;
  assign n2110 = ~n2108 & ~n2109;
  assign n2111 = ~n4834 & ~n2108;
  assign n2112 = ~n2109 & n2111;
  assign n2113 = ~n4834 & n2110;
  assign n2114 = n2094 & ~n4835;
  assign n2115 = ~n2103 & ~n2114;
  assign n2116 = ~n4833 & n2115;
  assign n2117 = ~pi359  & pi487 ;
  assign n2118 = ~pi358  & pi486 ;
  assign n2119 = ~n2117 & ~n2118;
  assign n2120 = ~pi357  & pi485 ;
  assign n2121 = ~pi356  & pi484 ;
  assign n2122 = ~n2120 & ~n2121;
  assign n2123 = n2119 & n2122;
  assign n2124 = ~n2116 & n2123;
  assign n2125 = pi359  & ~pi487 ;
  assign n2126 = pi356  & ~pi484 ;
  assign n2127 = ~n2120 & n2126;
  assign n2128 = pi358  & ~pi486 ;
  assign n2129 = pi357  & ~pi485 ;
  assign n2130 = ~n2128 & ~n2129;
  assign n2131 = ~n2127 & n2130;
  assign n2132 = n2119 & ~n2131;
  assign n2133 = ~n2127 & ~n2129;
  assign n2134 = n2119 & ~n2133;
  assign n2135 = ~pi486  & ~n2117;
  assign n2136 = pi358  & n2135;
  assign n2137 = ~n2117 & n2128;
  assign n2138 = ~n2125 & ~n4836;
  assign n2139 = ~n2134 & n2138;
  assign n2140 = ~n2125 & ~n2132;
  assign n2141 = ~n2124 & ~n4836;
  assign n2142 = ~n2134 & n2141;
  assign n2143 = ~n2125 & n2142;
  assign n2144 = ~n2124 & n4837;
  assign n2145 = ~pi363  & pi491 ;
  assign n2146 = ~pi362  & pi490 ;
  assign n2147 = ~n2145 & ~n2146;
  assign n2148 = ~pi361  & pi489 ;
  assign n2149 = ~pi360  & pi488 ;
  assign n2150 = ~n2148 & ~n2149;
  assign n2151 = n2147 & n2150;
  assign n2152 = ~n4838 & n2151;
  assign n2153 = pi363  & ~pi491 ;
  assign n2154 = pi360  & ~pi488 ;
  assign n2155 = ~n2148 & n2154;
  assign n2156 = pi361  & ~pi489 ;
  assign n2157 = pi362  & ~pi490 ;
  assign n2158 = ~n2156 & ~n2157;
  assign n2159 = ~n2155 & ~n2156;
  assign n2160 = ~n2157 & n2159;
  assign n2161 = ~n2155 & n2158;
  assign n2162 = n2147 & ~n4839;
  assign n2163 = ~n2153 & ~n2162;
  assign n2164 = ~n2152 & n2163;
  assign n2165 = ~pi367  & pi495 ;
  assign n2166 = ~pi366  & pi494 ;
  assign n2167 = ~n2165 & ~n2166;
  assign n2168 = ~pi365  & pi493 ;
  assign n2169 = ~pi364  & pi492 ;
  assign n2170 = ~n2168 & ~n2169;
  assign n2171 = n2167 & n2170;
  assign n2172 = ~n2164 & n2171;
  assign n2173 = pi367  & ~pi495 ;
  assign n2174 = pi364  & ~pi492 ;
  assign n2175 = ~n2168 & n2174;
  assign n2176 = pi366  & ~pi494 ;
  assign n2177 = pi365  & ~pi493 ;
  assign n2178 = ~n2176 & ~n2177;
  assign n2179 = ~n2175 & n2178;
  assign n2180 = n2167 & ~n2179;
  assign n2181 = ~n2175 & ~n2177;
  assign n2182 = n2167 & ~n2181;
  assign n2183 = ~pi494  & ~n2165;
  assign n2184 = pi366  & n2183;
  assign n2185 = ~n2165 & n2176;
  assign n2186 = ~n2173 & ~n4840;
  assign n2187 = ~n2182 & n2186;
  assign n2188 = ~n2173 & ~n2180;
  assign n2189 = ~n2172 & ~n4840;
  assign n2190 = ~n2182 & n2189;
  assign n2191 = ~n2173 & n2190;
  assign n2192 = ~n2172 & n4841;
  assign n2193 = ~pi371  & pi499 ;
  assign n2194 = ~pi370  & pi498 ;
  assign n2195 = ~n2193 & ~n2194;
  assign n2196 = ~pi369  & pi497 ;
  assign n2197 = ~pi368  & pi496 ;
  assign n2198 = ~n2196 & ~n2197;
  assign n2199 = n2195 & n2198;
  assign n2200 = ~n4842 & ~n2196;
  assign n2201 = n2195 & n2200;
  assign n2202 = ~n2197 & n2201;
  assign n2203 = ~n4842 & n2199;
  assign n2204 = pi371  & ~pi499 ;
  assign n2205 = pi368  & ~pi496 ;
  assign n2206 = ~pi496  & ~n2196;
  assign n2207 = pi368  & n2206;
  assign n2208 = ~n2196 & n2205;
  assign n2209 = pi369  & ~pi497 ;
  assign n2210 = pi370  & ~pi498 ;
  assign n2211 = ~n2209 & ~n2210;
  assign n2212 = ~n4844 & ~n2209;
  assign n2213 = ~n2210 & n2212;
  assign n2214 = ~n4844 & n2211;
  assign n2215 = n2195 & ~n4845;
  assign n2216 = ~n2204 & ~n2215;
  assign n2217 = ~n4843 & n2216;
  assign n2218 = ~pi375  & pi503 ;
  assign n2219 = ~pi374  & pi502 ;
  assign n2220 = ~n2218 & ~n2219;
  assign n2221 = ~pi373  & pi501 ;
  assign n2222 = ~pi372  & pi500 ;
  assign n2223 = ~n2221 & ~n2222;
  assign n2224 = n2220 & n2223;
  assign n2225 = ~n2217 & n2224;
  assign n2226 = pi375  & ~pi503 ;
  assign n2227 = pi372  & ~pi500 ;
  assign n2228 = ~n2221 & n2227;
  assign n2229 = pi374  & ~pi502 ;
  assign n2230 = pi373  & ~pi501 ;
  assign n2231 = ~n2229 & ~n2230;
  assign n2232 = ~n2228 & n2231;
  assign n2233 = n2220 & ~n2232;
  assign n2234 = ~n2228 & ~n2230;
  assign n2235 = n2220 & ~n2234;
  assign n2236 = ~pi502  & ~n2218;
  assign n2237 = pi374  & n2236;
  assign n2238 = ~n2218 & n2229;
  assign n2239 = ~n2226 & ~n4846;
  assign n2240 = ~n2235 & n2239;
  assign n2241 = ~n2226 & ~n2233;
  assign n2242 = ~n2225 & ~n4846;
  assign n2243 = ~n2235 & n2242;
  assign n2244 = ~n2226 & n2243;
  assign n2245 = ~n2225 & n4847;
  assign n2246 = ~pi379  & pi507 ;
  assign n2247 = ~pi378  & pi506 ;
  assign n2248 = ~n2246 & ~n2247;
  assign n2249 = ~pi377  & pi505 ;
  assign n2250 = ~pi376  & pi504 ;
  assign n2251 = ~n2249 & ~n2250;
  assign n2252 = n2248 & n2251;
  assign n2253 = ~n4848 & n2252;
  assign n2254 = pi379  & ~pi507 ;
  assign n2255 = pi376  & ~pi504 ;
  assign n2256 = ~n2249 & n2255;
  assign n2257 = pi377  & ~pi505 ;
  assign n2258 = pi378  & ~pi506 ;
  assign n2259 = ~n2257 & ~n2258;
  assign n2260 = ~n2256 & ~n2257;
  assign n2261 = ~n2258 & n2260;
  assign n2262 = ~n2256 & n2259;
  assign n2263 = n2248 & ~n4849;
  assign n2264 = ~n2254 & ~n2263;
  assign n2265 = ~n2253 & n2264;
  assign n2266 = ~pi382  & pi510 ;
  assign n2267 = ~pi381  & pi509 ;
  assign n2268 = ~n2266 & ~n2267;
  assign n2269 = pi383  & ~pi511 ;
  assign n2270 = ~pi380  & pi508 ;
  assign n2271 = ~n2269 & ~n2270;
  assign n2272 = n2268 & ~n2269;
  assign n2273 = ~n2270 & n2272;
  assign n2274 = n2268 & n2271;
  assign n2275 = ~n2265 & n4850;
  assign n2276 = pi380  & ~pi508 ;
  assign n2277 = pi381  & ~pi509 ;
  assign n2278 = ~n2276 & ~n2277;
  assign n2279 = n2268 & ~n2278;
  assign n2280 = pi382  & ~pi510 ;
  assign n2281 = ~n2279 & ~n2280;
  assign n2282 = ~n2269 & ~n2281;
  assign n2283 = ~pi383  & pi511 ;
  assign n2284 = ~n2282 & ~n2283;
  assign n2285 = ~n2275 & ~n2282;
  assign n2286 = ~n2283 & n2285;
  assign n2287 = ~n2275 & n2284;
  assign n2288 = pi284  & ~n4851;
  assign n2289 = pi412  & n4851;
  assign n2290 = ~n2288 & ~n2289;
  assign n2291 = n1465 & ~n2290;
  assign n2292 = pi27  & ~n4767;
  assign n2293 = pi155  & n4767;
  assign n2294 = ~n2292 & ~n2293;
  assign n2295 = pi283  & ~n4851;
  assign n2296 = pi411  & n4851;
  assign n2297 = ~n2295 & ~n2296;
  assign n2298 = ~n2294 & n2297;
  assign n2299 = pi26  & ~n4767;
  assign n2300 = pi154  & n4767;
  assign n2301 = ~n2299 & ~n2300;
  assign n2302 = pi25  & ~n4767;
  assign n2303 = pi153  & n4767;
  assign n2304 = ~n2302 & ~n2303;
  assign n2305 = pi281  & ~n4851;
  assign n2306 = pi409  & n4851;
  assign n2307 = ~n2305 & ~n2306;
  assign n2308 = ~n2304 & n2307;
  assign n2309 = pi20  & ~n4767;
  assign n2310 = pi148  & n4767;
  assign n2311 = ~n2309 & ~n2310;
  assign n2312 = pi19  & ~n4767;
  assign n2313 = pi147  & n4767;
  assign n2314 = ~n2312 & ~n2313;
  assign n2315 = pi275  & ~n4851;
  assign n2316 = pi403  & n4851;
  assign n2317 = ~n2315 & ~n2316;
  assign n2318 = ~n2314 & n2317;
  assign n2319 = pi18  & ~n4767;
  assign n2320 = pi146  & n4767;
  assign n2321 = ~n2319 & ~n2320;
  assign n2322 = pi17  & ~n4767;
  assign n2323 = pi145  & n4767;
  assign n2324 = ~n2322 & ~n2323;
  assign n2325 = pi273  & ~n4851;
  assign n2326 = pi401  & n4851;
  assign n2327 = ~n2325 & ~n2326;
  assign n2328 = ~n2324 & n2327;
  assign n2329 = pi13  & ~n4767;
  assign n2330 = pi141  & n4767;
  assign n2331 = ~n2329 & ~n2330;
  assign n2332 = pi269  & ~n4851;
  assign n2333 = pi397  & n4851;
  assign n2334 = ~n2332 & ~n2333;
  assign n2335 = n2331 & ~n2334;
  assign n2336 = pi12  & ~n4767;
  assign n2337 = pi140  & n4767;
  assign n2338 = ~n2336 & ~n2337;
  assign n2339 = pi268  & ~n4851;
  assign n2340 = pi396  & n4851;
  assign n2341 = ~n2339 & ~n2340;
  assign n2342 = ~n2338 & n2341;
  assign n2343 = pi11  & ~n4767;
  assign n2344 = pi139  & n4767;
  assign n2345 = ~n2343 & ~n2344;
  assign n2346 = pi10  & ~n4767;
  assign n2347 = pi138  & n4767;
  assign n2348 = ~n2346 & ~n2347;
  assign n2349 = pi266  & ~n4851;
  assign n2350 = pi394  & n4851;
  assign n2351 = ~n2349 & ~n2350;
  assign n2352 = ~n2348 & n2351;
  assign n2353 = pi262  & ~n4851;
  assign n2354 = pi390  & n4851;
  assign n2355 = ~n2353 & ~n2354;
  assign n2356 = pi6  & ~n4767;
  assign n2357 = pi134  & n4767;
  assign n2358 = ~n2356 & ~n2357;
  assign n2359 = ~n2355 & n2358;
  assign n2360 = pi4  & ~n4767;
  assign n2361 = pi132  & n4767;
  assign n2362 = ~n2360 & ~n2361;
  assign n2363 = pi3  & ~n4767;
  assign n2364 = pi131  & n4767;
  assign n2365 = ~n2363 & ~n2364;
  assign n2366 = pi259  & ~n4851;
  assign n2367 = pi387  & n4851;
  assign n2368 = ~n2366 & ~n2367;
  assign n2369 = ~n2365 & n2368;
  assign n2370 = n2365 & ~n2368;
  assign n2371 = pi2  & ~n4767;
  assign n2372 = pi130  & n4767;
  assign n2373 = ~n2371 & ~n2372;
  assign n2374 = pi258  & ~n4851;
  assign n2375 = pi386  & n4851;
  assign n2376 = ~n2374 & ~n2375;
  assign n2377 = ~n2373 & n2376;
  assign n2378 = n2373 & ~n2376;
  assign n2379 = pi1  & ~n4767;
  assign n2380 = pi129  & n4767;
  assign n2381 = ~n2379 & ~n2380;
  assign n2382 = pi257  & ~n4851;
  assign n2383 = pi385  & n4851;
  assign n2384 = ~n2382 & ~n2383;
  assign n2385 = n2381 & ~n2384;
  assign n2386 = pi256  & ~n4851;
  assign n2387 = pi384  & n4851;
  assign n2388 = ~n2386 & ~n2387;
  assign n2389 = pi0  & ~n4767;
  assign n2390 = pi128  & n4767;
  assign n2391 = ~n2389 & ~n2390;
  assign n2392 = n2388 & ~n2391;
  assign n2393 = ~n2385 & n2392;
  assign n2394 = ~n2381 & n2384;
  assign n2395 = ~n2392 & ~n2394;
  assign n2396 = ~n2385 & ~n2395;
  assign n2397 = ~n2393 & ~n2394;
  assign n2398 = n2384 & n2392;
  assign n2399 = n2381 & ~n2398;
  assign n2400 = ~n2384 & ~n2392;
  assign n2401 = ~n2378 & ~n2400;
  assign n2402 = ~n2399 & n2401;
  assign n2403 = ~n2378 & n4852;
  assign n2404 = n2381 & ~n2392;
  assign n2405 = n2384 & ~n2404;
  assign n2406 = ~n2381 & n2392;
  assign n2407 = ~n2377 & ~n2406;
  assign n2408 = ~n2377 & ~n4852;
  assign n2409 = ~n2405 & n2407;
  assign n2410 = ~n2378 & ~n4854;
  assign n2411 = ~n2377 & ~n4853;
  assign n2412 = ~n2370 & n4855;
  assign n2413 = ~n2369 & ~n4855;
  assign n2414 = ~n2370 & ~n2413;
  assign n2415 = ~n2369 & ~n2412;
  assign n2416 = pi260  & ~n4851;
  assign n2417 = pi388  & n4851;
  assign n2418 = ~n2416 & ~n2417;
  assign n2419 = n4856 & n2418;
  assign n2420 = n2362 & ~n2419;
  assign n2421 = ~n4856 & ~n2418;
  assign n2422 = pi5  & ~n4767;
  assign n2423 = pi133  & n4767;
  assign n2424 = ~n2422 & ~n2423;
  assign n2425 = pi261  & ~n4851;
  assign n2426 = pi389  & n4851;
  assign n2427 = ~n2425 & ~n2426;
  assign n2428 = n2424 & ~n2427;
  assign n2429 = ~n2421 & ~n2428;
  assign n2430 = ~n2420 & n2429;
  assign n2431 = ~n2424 & n2427;
  assign n2432 = n2362 & ~n4856;
  assign n2433 = n2418 & ~n2432;
  assign n2434 = ~n2362 & n4856;
  assign n2435 = ~n2420 & ~n2421;
  assign n2436 = ~n2433 & ~n2434;
  assign n2437 = n2427 & n4857;
  assign n2438 = n2424 & ~n2437;
  assign n2439 = ~n2427 & ~n4857;
  assign n2440 = ~n2438 & ~n2439;
  assign n2441 = n2424 & ~n4857;
  assign n2442 = n2427 & ~n2441;
  assign n2443 = ~n2424 & n4857;
  assign n2444 = ~n2442 & ~n2443;
  assign n2445 = ~n2430 & ~n2431;
  assign n2446 = ~n2359 & n4858;
  assign n2447 = n2355 & ~n2358;
  assign n2448 = pi7  & ~n4767;
  assign n2449 = pi135  & n4767;
  assign n2450 = ~n2448 & ~n2449;
  assign n2451 = pi263  & ~n4851;
  assign n2452 = pi391  & n4851;
  assign n2453 = ~n2451 & ~n2452;
  assign n2454 = ~n2450 & n2453;
  assign n2455 = ~n2447 & ~n2454;
  assign n2456 = n2358 & ~n4858;
  assign n2457 = n2355 & ~n2456;
  assign n2458 = ~n2358 & n4858;
  assign n2459 = ~n2355 & ~n4858;
  assign n2460 = n2355 & n4858;
  assign n2461 = n2358 & ~n2460;
  assign n2462 = ~n2459 & ~n2461;
  assign n2463 = ~n2457 & ~n2458;
  assign n2464 = ~n2454 & ~n4859;
  assign n2465 = ~n2446 & n2455;
  assign n2466 = pi8  & ~n4767;
  assign n2467 = pi136  & n4767;
  assign n2468 = ~n2466 & ~n2467;
  assign n2469 = pi264  & ~n4851;
  assign n2470 = pi392  & n4851;
  assign n2471 = ~n2469 & ~n2470;
  assign n2472 = n2468 & ~n2471;
  assign n2473 = n2450 & ~n2453;
  assign n2474 = ~n2472 & ~n2473;
  assign n2475 = ~n4860 & n2474;
  assign n2476 = ~n2468 & n2471;
  assign n2477 = pi9  & ~n4767;
  assign n2478 = pi137  & n4767;
  assign n2479 = ~n2477 & ~n2478;
  assign n2480 = pi265  & ~n4851;
  assign n2481 = pi393  & n4851;
  assign n2482 = ~n2480 & ~n2481;
  assign n2483 = ~n2479 & n2482;
  assign n2484 = ~n2476 & ~n2483;
  assign n2485 = ~n2475 & n2484;
  assign n2486 = n2348 & ~n2351;
  assign n2487 = n2479 & ~n2482;
  assign n2488 = ~n2486 & ~n2487;
  assign n2489 = n4859 & ~n2473;
  assign n2490 = ~n2454 & ~n2476;
  assign n2491 = ~n2489 & n2490;
  assign n2492 = ~n2454 & ~n2489;
  assign n2493 = n2468 & n2492;
  assign n2494 = n2471 & ~n2493;
  assign n2495 = ~n2468 & ~n2492;
  assign n2496 = ~n2494 & ~n2495;
  assign n2497 = ~n2472 & ~n2491;
  assign n2498 = n2479 & n4861;
  assign n2499 = n2482 & ~n2498;
  assign n2500 = ~n2479 & ~n4861;
  assign n2501 = ~n2499 & ~n2500;
  assign n2502 = ~n2486 & ~n2501;
  assign n2503 = ~n2485 & n2488;
  assign n2504 = ~n2352 & ~n4862;
  assign n2505 = pi267  & ~n4851;
  assign n2506 = pi395  & n4851;
  assign n2507 = ~n2505 & ~n2506;
  assign n2508 = ~n2504 & n2507;
  assign n2509 = n2345 & ~n2508;
  assign n2510 = n2338 & ~n2341;
  assign n2511 = n2504 & ~n2507;
  assign n2512 = ~n2510 & ~n2511;
  assign n2513 = n2345 & ~n2507;
  assign n2514 = ~n2504 & ~n2513;
  assign n2515 = ~n2345 & n2507;
  assign n2516 = ~n2514 & ~n2515;
  assign n2517 = ~n2510 & ~n2516;
  assign n2518 = ~n2509 & n2512;
  assign n2519 = ~n2342 & ~n4863;
  assign n2520 = ~n2335 & ~n2519;
  assign n2521 = ~n2331 & n2334;
  assign n2522 = pi14  & ~n4767;
  assign n2523 = pi142  & n4767;
  assign n2524 = ~n2522 & ~n2523;
  assign n2525 = pi270  & ~n4851;
  assign n2526 = pi398  & n4851;
  assign n2527 = ~n2525 & ~n2526;
  assign n2528 = ~n2524 & n2527;
  assign n2529 = ~n2521 & ~n2528;
  assign n2530 = ~n2520 & n2529;
  assign n2531 = n2524 & ~n2527;
  assign n2532 = pi15  & ~n4767;
  assign n2533 = pi143  & n4767;
  assign n2534 = ~n2532 & ~n2533;
  assign n2535 = pi271  & ~n4851;
  assign n2536 = pi399  & n4851;
  assign n2537 = ~n2535 & ~n2536;
  assign n2538 = n2534 & ~n2537;
  assign n2539 = ~n2531 & ~n2538;
  assign n2540 = ~n2520 & ~n2521;
  assign n2541 = ~n2531 & ~n2540;
  assign n2542 = ~n2528 & ~n2541;
  assign n2543 = ~n2538 & ~n2542;
  assign n2544 = ~n2530 & n2539;
  assign n2545 = ~n2534 & n2537;
  assign n2546 = pi16  & ~n4767;
  assign n2547 = pi144  & n4767;
  assign n2548 = ~n2546 & ~n2547;
  assign n2549 = pi272  & ~n4851;
  assign n2550 = pi400  & n4851;
  assign n2551 = ~n2549 & ~n2550;
  assign n2552 = ~n2548 & n2551;
  assign n2553 = ~n2545 & ~n2552;
  assign n2554 = ~n4864 & n2553;
  assign n2555 = n2548 & ~n2551;
  assign n2556 = n2324 & ~n2327;
  assign n2557 = ~n2555 & ~n2556;
  assign n2558 = ~n2554 & n2557;
  assign n2559 = ~n4864 & ~n2545;
  assign n2560 = n2548 & n2559;
  assign n2561 = n2551 & ~n2560;
  assign n2562 = ~n2548 & ~n2559;
  assign n2563 = ~n2561 & ~n2562;
  assign n2564 = ~n2554 & ~n2555;
  assign n2565 = n2324 & n4865;
  assign n2566 = n2327 & ~n2565;
  assign n2567 = ~n2324 & ~n4865;
  assign n2568 = ~n2566 & ~n2567;
  assign n2569 = ~n2328 & ~n2558;
  assign n2570 = pi274  & ~n4851;
  assign n2571 = pi402  & n4851;
  assign n2572 = ~n2570 & ~n2571;
  assign n2573 = ~n4866 & n2572;
  assign n2574 = n2321 & ~n2573;
  assign n2575 = n2314 & ~n2317;
  assign n2576 = n4866 & ~n2572;
  assign n2577 = ~n2575 & ~n2576;
  assign n2578 = n2321 & ~n2572;
  assign n2579 = ~n4866 & ~n2578;
  assign n2580 = ~n2321 & n2572;
  assign n2581 = ~n2579 & ~n2580;
  assign n2582 = ~n2575 & ~n2581;
  assign n2583 = ~n2574 & n2577;
  assign n2584 = ~n2318 & ~n4867;
  assign n2585 = pi276  & ~n4851;
  assign n2586 = pi404  & n4851;
  assign n2587 = ~n2585 & ~n2586;
  assign n2588 = ~n2584 & n2587;
  assign n2589 = n2311 & ~n2588;
  assign n2590 = pi21  & ~n4767;
  assign n2591 = pi149  & n4767;
  assign n2592 = ~n2590 & ~n2591;
  assign n2593 = pi277  & ~n4851;
  assign n2594 = pi405  & n4851;
  assign n2595 = ~n2593 & ~n2594;
  assign n2596 = n2592 & ~n2595;
  assign n2597 = n2584 & ~n2587;
  assign n2598 = ~n2596 & ~n2597;
  assign n2599 = n2311 & ~n2587;
  assign n2600 = ~n2584 & ~n2599;
  assign n2601 = ~n2311 & n2587;
  assign n2602 = ~n2600 & ~n2601;
  assign n2603 = ~n2596 & ~n2602;
  assign n2604 = ~n2589 & n2598;
  assign n2605 = ~n2592 & n2595;
  assign n2606 = pi22  & ~n4767;
  assign n2607 = pi150  & n4767;
  assign n2608 = ~n2606 & ~n2607;
  assign n2609 = pi278  & ~n4851;
  assign n2610 = pi406  & n4851;
  assign n2611 = ~n2609 & ~n2610;
  assign n2612 = ~n2608 & n2611;
  assign n2613 = ~n2605 & ~n2612;
  assign n2614 = ~n4868 & n2613;
  assign n2615 = n2608 & ~n2611;
  assign n2616 = pi23  & ~n4767;
  assign n2617 = pi151  & n4767;
  assign n2618 = ~n2616 & ~n2617;
  assign n2619 = pi279  & ~n4851;
  assign n2620 = pi407  & n4851;
  assign n2621 = ~n2619 & ~n2620;
  assign n2622 = n2618 & ~n2621;
  assign n2623 = ~n2615 & ~n2622;
  assign n2624 = ~n4868 & ~n2605;
  assign n2625 = ~n2615 & ~n2624;
  assign n2626 = ~n2612 & ~n2625;
  assign n2627 = ~n2622 & ~n2626;
  assign n2628 = ~n2614 & n2623;
  assign n2629 = ~n2618 & n2621;
  assign n2630 = pi24  & ~n4767;
  assign n2631 = pi152  & n4767;
  assign n2632 = ~n2630 & ~n2631;
  assign n2633 = pi280  & ~n4851;
  assign n2634 = pi408  & n4851;
  assign n2635 = ~n2633 & ~n2634;
  assign n2636 = ~n2632 & n2635;
  assign n2637 = ~n2629 & ~n2636;
  assign n2638 = ~n4869 & n2637;
  assign n2639 = n2632 & ~n2635;
  assign n2640 = n2304 & ~n2307;
  assign n2641 = ~n2639 & ~n2640;
  assign n2642 = ~n2638 & n2641;
  assign n2643 = ~n4869 & ~n2629;
  assign n2644 = n2632 & n2643;
  assign n2645 = n2635 & ~n2644;
  assign n2646 = ~n2632 & ~n2643;
  assign n2647 = ~n2645 & ~n2646;
  assign n2648 = ~n2638 & ~n2639;
  assign n2649 = n2304 & n4870;
  assign n2650 = n2307 & ~n2649;
  assign n2651 = ~n2304 & ~n4870;
  assign n2652 = ~n2650 & ~n2651;
  assign n2653 = ~n2308 & ~n2642;
  assign n2654 = pi282  & ~n4851;
  assign n2655 = pi410  & n4851;
  assign n2656 = ~n2654 & ~n2655;
  assign n2657 = ~n4871 & n2656;
  assign n2658 = n2301 & ~n2657;
  assign n2659 = n2294 & ~n2297;
  assign n2660 = n4871 & ~n2656;
  assign n2661 = ~n2659 & ~n2660;
  assign n2662 = n2301 & ~n2656;
  assign n2663 = ~n4871 & ~n2662;
  assign n2664 = ~n2301 & n2656;
  assign n2665 = ~n2663 & ~n2664;
  assign n2666 = ~n2659 & ~n2665;
  assign n2667 = ~n2658 & n2661;
  assign n2668 = ~n2298 & ~n4872;
  assign n2669 = ~n2291 & ~n2668;
  assign n2670 = ~n1465 & n2290;
  assign n2671 = pi29  & ~n4767;
  assign n2672 = pi157  & n4767;
  assign n2673 = ~n2671 & ~n2672;
  assign n2674 = pi285  & ~n4851;
  assign n2675 = pi413  & n4851;
  assign n2676 = ~n2674 & ~n2675;
  assign n2677 = ~n2673 & n2676;
  assign n2678 = ~n2670 & ~n2677;
  assign n2679 = ~n2669 & n2678;
  assign n2680 = n2673 & ~n2676;
  assign n2681 = pi30  & ~n4767;
  assign n2682 = pi158  & n4767;
  assign n2683 = ~n2681 & ~n2682;
  assign n2684 = pi286  & ~n4851;
  assign n2685 = pi414  & n4851;
  assign n2686 = ~n2684 & ~n2685;
  assign n2687 = n2683 & ~n2686;
  assign n2688 = ~n2680 & ~n2687;
  assign n2689 = ~n2669 & ~n2670;
  assign n2690 = ~n2680 & ~n2689;
  assign n2691 = ~n2677 & ~n2690;
  assign n2692 = ~n2687 & ~n2691;
  assign n2693 = ~n2679 & n2688;
  assign n2694 = ~n2683 & n2686;
  assign n2695 = pi31  & ~n4767;
  assign n2696 = pi159  & n4767;
  assign n2697 = ~n2695 & ~n2696;
  assign n2698 = pi287  & ~n4851;
  assign n2699 = pi415  & n4851;
  assign n2700 = ~n2698 & ~n2699;
  assign n2701 = ~n2697 & n2700;
  assign n2702 = ~n2694 & ~n2701;
  assign n2703 = ~n4873 & n2702;
  assign n2704 = pi294  & ~n4851;
  assign n2705 = pi422  & n4851;
  assign n2706 = ~n2704 & ~n2705;
  assign n2707 = pi38  & ~n4767;
  assign n2708 = pi166  & n4767;
  assign n2709 = ~n2707 & ~n2708;
  assign n2710 = ~n2706 & n2709;
  assign n2711 = pi37  & ~n4767;
  assign n2712 = pi165  & n4767;
  assign n2713 = ~n2711 & ~n2712;
  assign n2714 = pi293  & ~n4851;
  assign n2715 = pi421  & n4851;
  assign n2716 = ~n2714 & ~n2715;
  assign n2717 = n2713 & ~n2716;
  assign n2718 = pi39  & ~n4767;
  assign n2719 = pi167  & n4767;
  assign n2720 = ~n2718 & ~n2719;
  assign n2721 = pi295  & ~n4851;
  assign n2722 = pi423  & n4851;
  assign n2723 = ~n2721 & ~n2722;
  assign n2724 = n2720 & ~n2723;
  assign n2725 = ~n2717 & ~n2724;
  assign n2726 = ~n2710 & ~n2717;
  assign n2727 = ~n2724 & n2726;
  assign n2728 = ~n2710 & n2725;
  assign n2729 = pi290  & ~n4851;
  assign n2730 = pi418  & n4851;
  assign n2731 = ~n2729 & ~n2730;
  assign n2732 = pi34  & ~n4767;
  assign n2733 = pi162  & n4767;
  assign n2734 = ~n2732 & ~n2733;
  assign n2735 = ~n2731 & n2734;
  assign n2736 = pi33  & ~n4767;
  assign n2737 = pi161  & n4767;
  assign n2738 = ~n2736 & ~n2737;
  assign n2739 = pi289  & ~n4851;
  assign n2740 = pi417  & n4851;
  assign n2741 = ~n2739 & ~n2740;
  assign n2742 = n2738 & ~n2741;
  assign n2743 = pi35  & ~n4767;
  assign n2744 = pi163  & n4767;
  assign n2745 = ~n2743 & ~n2744;
  assign n2746 = pi291  & ~n4851;
  assign n2747 = pi419  & n4851;
  assign n2748 = ~n2746 & ~n2747;
  assign n2749 = n2745 & ~n2748;
  assign n2750 = ~n2742 & ~n2749;
  assign n2751 = ~n2735 & ~n2749;
  assign n2752 = ~n2742 & n2751;
  assign n2753 = ~n2735 & n2750;
  assign n2754 = pi288  & ~n4851;
  assign n2755 = pi416  & n4851;
  assign n2756 = ~n2754 & ~n2755;
  assign n2757 = pi32  & ~n4767;
  assign n2758 = pi160  & n4767;
  assign n2759 = ~n2757 & ~n2758;
  assign n2760 = ~n2756 & n2759;
  assign n2761 = pi36  & ~n4767;
  assign n2762 = pi164  & n4767;
  assign n2763 = ~n2761 & ~n2762;
  assign n2764 = pi292  & ~n4851;
  assign n2765 = pi420  & n4851;
  assign n2766 = ~n2764 & ~n2765;
  assign n2767 = n2763 & ~n2766;
  assign n2768 = n2697 & ~n2700;
  assign n2769 = ~n2767 & ~n2768;
  assign n2770 = ~n2760 & n2769;
  assign n2771 = n4875 & n2770;
  assign n2772 = n4874 & n2770;
  assign n2773 = n4875 & n2772;
  assign n2774 = ~n2710 & ~n2724;
  assign n2775 = ~n2717 & ~n2767;
  assign n2776 = n4874 & ~n2767;
  assign n2777 = n2774 & n2775;
  assign n2778 = ~n2760 & ~n2768;
  assign n2779 = n4875 & n2778;
  assign n2780 = n4877 & n2779;
  assign n2781 = n4874 & n2771;
  assign n2782 = ~n4873 & ~n2694;
  assign n2783 = ~n2768 & ~n2782;
  assign n2784 = ~n2701 & ~n2783;
  assign n2785 = n4875 & n4877;
  assign n2786 = ~n2784 & n2785;
  assign n2787 = ~n2760 & n2786;
  assign n2788 = ~n2760 & n4877;
  assign n2789 = n4875 & n2788;
  assign n2790 = ~n2784 & n2789;
  assign n2791 = ~n2703 & n4876;
  assign n2792 = n2756 & ~n2759;
  assign n2793 = ~n2738 & n2741;
  assign n2794 = ~n2792 & ~n2793;
  assign n2795 = n4875 & ~n2794;
  assign n2796 = n2731 & ~n2734;
  assign n2797 = n2731 & ~n2749;
  assign n2798 = ~n2734 & n2797;
  assign n2799 = ~n2749 & n2796;
  assign n2800 = ~n2745 & n2748;
  assign n2801 = ~n4879 & ~n2800;
  assign n2802 = ~n2795 & ~n4879;
  assign n2803 = ~n2800 & n2802;
  assign n2804 = ~n2795 & n2801;
  assign n2805 = n4877 & ~n4880;
  assign n2806 = n2706 & ~n2709;
  assign n2807 = n2706 & ~n2724;
  assign n2808 = ~n2709 & n2807;
  assign n2809 = ~n2724 & n2806;
  assign n2810 = ~n2720 & n2723;
  assign n2811 = ~n4881 & ~n2810;
  assign n2812 = ~n2713 & n2716;
  assign n2813 = ~n2763 & n2766;
  assign n2814 = ~n2717 & n2813;
  assign n2815 = ~n2812 & ~n2814;
  assign n2816 = ~n2812 & ~n2813;
  assign n2817 = n4874 & ~n2816;
  assign n2818 = n2774 & ~n2815;
  assign n2819 = n2811 & ~n4882;
  assign n2820 = ~n2767 & ~n4880;
  assign n2821 = n2816 & ~n2820;
  assign n2822 = n4874 & ~n2821;
  assign n2823 = n2811 & ~n2822;
  assign n2824 = ~n2805 & ~n4881;
  assign n2825 = ~n4882 & n2824;
  assign n2826 = ~n2810 & n2825;
  assign n2827 = ~n2805 & n2819;
  assign n2828 = ~n4878 & n4883;
  assign n2829 = pi302  & ~n4851;
  assign n2830 = pi430  & n4851;
  assign n2831 = ~n2829 & ~n2830;
  assign n2832 = pi46  & ~n4767;
  assign n2833 = pi174  & n4767;
  assign n2834 = ~n2832 & ~n2833;
  assign n2835 = ~n2831 & n2834;
  assign n2836 = pi47  & ~n4767;
  assign n2837 = pi175  & n4767;
  assign n2838 = ~n2836 & ~n2837;
  assign n2839 = pi303  & ~n4851;
  assign n2840 = pi431  & n4851;
  assign n2841 = ~n2839 & ~n2840;
  assign n2842 = n2838 & ~n2841;
  assign n2843 = ~n2835 & ~n2842;
  assign n2844 = pi45  & ~n4767;
  assign n2845 = pi173  & n4767;
  assign n2846 = ~n2844 & ~n2845;
  assign n2847 = pi301  & ~n4851;
  assign n2848 = pi429  & n4851;
  assign n2849 = ~n2847 & ~n2848;
  assign n2850 = n2846 & ~n2849;
  assign n2851 = pi44  & ~n4767;
  assign n2852 = pi172  & n4767;
  assign n2853 = ~n2851 & ~n2852;
  assign n2854 = pi300  & ~n4851;
  assign n2855 = pi428  & n4851;
  assign n2856 = ~n2854 & ~n2855;
  assign n2857 = n2853 & ~n2856;
  assign n2858 = ~n2850 & ~n2857;
  assign n2859 = ~n2842 & ~n2850;
  assign n2860 = ~n2835 & ~n2850;
  assign n2861 = ~n2842 & n2860;
  assign n2862 = ~n2835 & n2859;
  assign n2863 = ~n2857 & n4884;
  assign n2864 = n2843 & n2858;
  assign n2865 = pi43  & ~n4767;
  assign n2866 = pi171  & n4767;
  assign n2867 = ~n2865 & ~n2866;
  assign n2868 = pi299  & ~n4851;
  assign n2869 = pi427  & n4851;
  assign n2870 = ~n2868 & ~n2869;
  assign n2871 = n2867 & ~n2870;
  assign n2872 = pi42  & ~n4767;
  assign n2873 = pi170  & n4767;
  assign n2874 = ~n2872 & ~n2873;
  assign n2875 = pi298  & ~n4851;
  assign n2876 = pi426  & n4851;
  assign n2877 = ~n2875 & ~n2876;
  assign n2878 = n2874 & ~n2877;
  assign n2879 = ~n2871 & ~n2878;
  assign n2880 = pi41  & ~n4767;
  assign n2881 = pi169  & n4767;
  assign n2882 = ~n2880 & ~n2881;
  assign n2883 = pi297  & ~n4851;
  assign n2884 = pi425  & n4851;
  assign n2885 = ~n2883 & ~n2884;
  assign n2886 = n2882 & ~n2885;
  assign n2887 = pi40  & ~n4767;
  assign n2888 = pi168  & n4767;
  assign n2889 = ~n2887 & ~n2888;
  assign n2890 = pi296  & ~n4851;
  assign n2891 = pi424  & n4851;
  assign n2892 = ~n2890 & ~n2891;
  assign n2893 = n2889 & ~n2892;
  assign n2894 = ~n2886 & ~n2893;
  assign n2895 = n2879 & n2894;
  assign n2896 = ~n2857 & ~n2893;
  assign n2897 = ~n2886 & n2896;
  assign n2898 = n2879 & n2897;
  assign n2899 = n4884 & n2898;
  assign n2900 = n4885 & n2895;
  assign n2901 = ~n2828 & n4886;
  assign n2902 = ~n2867 & n2870;
  assign n2903 = ~n2889 & n2892;
  assign n2904 = ~n2886 & n2903;
  assign n2905 = ~n2874 & n2877;
  assign n2906 = ~n2882 & n2885;
  assign n2907 = ~n2905 & ~n2906;
  assign n2908 = ~n2904 & ~n2906;
  assign n2909 = ~n2905 & n2908;
  assign n2910 = ~n2904 & n2907;
  assign n2911 = n2879 & ~n4887;
  assign n2912 = ~n2902 & ~n2911;
  assign n2913 = n4885 & ~n2912;
  assign n2914 = n2831 & ~n2834;
  assign n2915 = ~n2842 & n2914;
  assign n2916 = ~n2838 & n2841;
  assign n2917 = ~n2915 & ~n2916;
  assign n2918 = ~n2846 & n2849;
  assign n2919 = ~n2853 & n2856;
  assign n2920 = ~n2850 & n2919;
  assign n2921 = ~n2918 & ~n2920;
  assign n2922 = ~n2918 & ~n2919;
  assign n2923 = n4884 & ~n2922;
  assign n2924 = n2843 & ~n2921;
  assign n2925 = n2917 & ~n4888;
  assign n2926 = ~n2857 & ~n2912;
  assign n2927 = n2922 & ~n2926;
  assign n2928 = n4884 & ~n2927;
  assign n2929 = n2917 & ~n2928;
  assign n2930 = ~n2913 & n2925;
  assign n2931 = ~n2901 & ~n2915;
  assign n2932 = ~n4888 & n2931;
  assign n2933 = ~n2913 & n2932;
  assign n2934 = ~n2916 & n2933;
  assign n2935 = ~n2901 & n4889;
  assign n2936 = pi55  & ~n4767;
  assign n2937 = pi183  & n4767;
  assign n2938 = ~n2936 & ~n2937;
  assign n2939 = pi311  & ~n4851;
  assign n2940 = pi439  & n4851;
  assign n2941 = ~n2939 & ~n2940;
  assign n2942 = n2938 & ~n2941;
  assign n2943 = pi310  & ~n4851;
  assign n2944 = pi438  & n4851;
  assign n2945 = ~n2943 & ~n2944;
  assign n2946 = pi54  & ~n4767;
  assign n2947 = pi182  & n4767;
  assign n2948 = ~n2946 & ~n2947;
  assign n2949 = ~n2945 & n2948;
  assign n2950 = ~n2942 & ~n2949;
  assign n2951 = pi53  & ~n4767;
  assign n2952 = pi181  & n4767;
  assign n2953 = ~n2951 & ~n2952;
  assign n2954 = pi309  & ~n4851;
  assign n2955 = pi437  & n4851;
  assign n2956 = ~n2954 & ~n2955;
  assign n2957 = n2953 & ~n2956;
  assign n2958 = pi308  & ~n4851;
  assign n2959 = pi436  & n4851;
  assign n2960 = ~n2958 & ~n2959;
  assign n2961 = pi52  & ~n4767;
  assign n2962 = pi180  & n4767;
  assign n2963 = ~n2961 & ~n2962;
  assign n2964 = ~n2960 & n2963;
  assign n2965 = ~n2957 & ~n2964;
  assign n2966 = n2950 & n2965;
  assign n2967 = pi306  & ~n4851;
  assign n2968 = pi434  & n4851;
  assign n2969 = ~n2967 & ~n2968;
  assign n2970 = pi50  & ~n4767;
  assign n2971 = pi178  & n4767;
  assign n2972 = ~n2970 & ~n2971;
  assign n2973 = ~n2969 & n2972;
  assign n2974 = pi49  & ~n4767;
  assign n2975 = pi177  & n4767;
  assign n2976 = ~n2974 & ~n2975;
  assign n2977 = pi305  & ~n4851;
  assign n2978 = pi433  & n4851;
  assign n2979 = ~n2977 & ~n2978;
  assign n2980 = n2976 & ~n2979;
  assign n2981 = pi51  & ~n4767;
  assign n2982 = pi179  & n4767;
  assign n2983 = ~n2981 & ~n2982;
  assign n2984 = pi307  & ~n4851;
  assign n2985 = pi435  & n4851;
  assign n2986 = ~n2984 & ~n2985;
  assign n2987 = n2983 & ~n2986;
  assign n2988 = ~n2980 & ~n2987;
  assign n2989 = ~n2973 & ~n2987;
  assign n2990 = ~n2980 & n2989;
  assign n2991 = ~n2973 & n2988;
  assign n2992 = pi304  & ~n4851;
  assign n2993 = pi432  & n4851;
  assign n2994 = ~n2992 & ~n2993;
  assign n2995 = pi48  & ~n4767;
  assign n2996 = pi176  & n4767;
  assign n2997 = ~n2995 & ~n2996;
  assign n2998 = ~n2994 & n2997;
  assign n2999 = n4891 & ~n2998;
  assign n3000 = n2966 & n4891;
  assign n3001 = ~n2998 & n3000;
  assign n3002 = n2966 & ~n2998;
  assign n3003 = n4891 & n3002;
  assign n3004 = n2966 & n2999;
  assign n3005 = ~n4890 & n4892;
  assign n3006 = n2994 & ~n2997;
  assign n3007 = ~n2976 & n2979;
  assign n3008 = ~n3006 & ~n3007;
  assign n3009 = n4891 & ~n3008;
  assign n3010 = ~n2983 & n2986;
  assign n3011 = n2969 & ~n2972;
  assign n3012 = n2969 & ~n2987;
  assign n3013 = ~n2972 & n3012;
  assign n3014 = ~n2987 & n3011;
  assign n3015 = ~n3010 & ~n4893;
  assign n3016 = ~n3009 & ~n4893;
  assign n3017 = ~n3010 & n3016;
  assign n3018 = ~n3009 & n3015;
  assign n3019 = n2966 & ~n4894;
  assign n3020 = ~n2938 & n2941;
  assign n3021 = n2960 & ~n2963;
  assign n3022 = ~n2957 & n3021;
  assign n3023 = ~n2953 & n2956;
  assign n3024 = n2945 & ~n2948;
  assign n3025 = ~n3023 & ~n3024;
  assign n3026 = ~n3022 & ~n3023;
  assign n3027 = ~n3024 & n3026;
  assign n3028 = ~n3022 & n3025;
  assign n3029 = n2950 & ~n4895;
  assign n3030 = ~n3020 & ~n3029;
  assign n3031 = ~n3019 & ~n3029;
  assign n3032 = ~n3020 & n3031;
  assign n3033 = ~n3019 & n3030;
  assign n3034 = ~n3005 & n4896;
  assign n3035 = pi318  & ~n4851;
  assign n3036 = pi446  & n4851;
  assign n3037 = ~n3035 & ~n3036;
  assign n3038 = pi62  & ~n4767;
  assign n3039 = pi190  & n4767;
  assign n3040 = ~n3038 & ~n3039;
  assign n3041 = ~n3037 & n3040;
  assign n3042 = pi63  & ~n4767;
  assign n3043 = pi191  & n4767;
  assign n3044 = ~n3042 & ~n3043;
  assign n3045 = pi319  & ~n4851;
  assign n3046 = pi447  & n4851;
  assign n3047 = ~n3045 & ~n3046;
  assign n3048 = n3044 & ~n3047;
  assign n3049 = ~n3041 & ~n3048;
  assign n3050 = pi61  & ~n4767;
  assign n3051 = pi189  & n4767;
  assign n3052 = ~n3050 & ~n3051;
  assign n3053 = pi317  & ~n4851;
  assign n3054 = pi445  & n4851;
  assign n3055 = ~n3053 & ~n3054;
  assign n3056 = n3052 & ~n3055;
  assign n3057 = pi60  & ~n4767;
  assign n3058 = pi188  & n4767;
  assign n3059 = ~n3057 & ~n3058;
  assign n3060 = pi316  & ~n4851;
  assign n3061 = pi444  & n4851;
  assign n3062 = ~n3060 & ~n3061;
  assign n3063 = n3059 & ~n3062;
  assign n3064 = ~n3056 & ~n3063;
  assign n3065 = ~n3048 & ~n3056;
  assign n3066 = ~n3041 & ~n3056;
  assign n3067 = ~n3048 & n3066;
  assign n3068 = ~n3041 & n3065;
  assign n3069 = ~n3063 & n4897;
  assign n3070 = n3049 & n3064;
  assign n3071 = pi59  & ~n4767;
  assign n3072 = pi187  & n4767;
  assign n3073 = ~n3071 & ~n3072;
  assign n3074 = pi315  & ~n4851;
  assign n3075 = pi443  & n4851;
  assign n3076 = ~n3074 & ~n3075;
  assign n3077 = n3073 & ~n3076;
  assign n3078 = pi58  & ~n4767;
  assign n3079 = pi186  & n4767;
  assign n3080 = ~n3078 & ~n3079;
  assign n3081 = pi314  & ~n4851;
  assign n3082 = pi442  & n4851;
  assign n3083 = ~n3081 & ~n3082;
  assign n3084 = n3080 & ~n3083;
  assign n3085 = ~n3077 & ~n3084;
  assign n3086 = pi57  & ~n4767;
  assign n3087 = pi185  & n4767;
  assign n3088 = ~n3086 & ~n3087;
  assign n3089 = pi313  & ~n4851;
  assign n3090 = pi441  & n4851;
  assign n3091 = ~n3089 & ~n3090;
  assign n3092 = n3088 & ~n3091;
  assign n3093 = pi56  & ~n4767;
  assign n3094 = pi184  & n4767;
  assign n3095 = ~n3093 & ~n3094;
  assign n3096 = pi312  & ~n4851;
  assign n3097 = pi440  & n4851;
  assign n3098 = ~n3096 & ~n3097;
  assign n3099 = n3095 & ~n3098;
  assign n3100 = ~n3092 & ~n3099;
  assign n3101 = n3085 & n3100;
  assign n3102 = ~n3063 & ~n3099;
  assign n3103 = ~n3092 & n3102;
  assign n3104 = n3085 & n3103;
  assign n3105 = n4897 & n3104;
  assign n3106 = n4898 & n3100;
  assign n3107 = n3085 & n3106;
  assign n3108 = n4898 & n3101;
  assign n3109 = ~n3034 & n4899;
  assign n3110 = ~n3073 & n3076;
  assign n3111 = ~n3095 & n3098;
  assign n3112 = ~n3092 & n3111;
  assign n3113 = ~n3080 & n3083;
  assign n3114 = ~n3088 & n3091;
  assign n3115 = ~n3113 & ~n3114;
  assign n3116 = ~n3112 & ~n3114;
  assign n3117 = ~n3113 & n3116;
  assign n3118 = ~n3112 & n3115;
  assign n3119 = n3085 & ~n4900;
  assign n3120 = ~n3110 & ~n3119;
  assign n3121 = n4898 & ~n3120;
  assign n3122 = n3037 & ~n3040;
  assign n3123 = ~n3048 & n3122;
  assign n3124 = ~n3044 & n3047;
  assign n3125 = ~n3123 & ~n3124;
  assign n3126 = ~n3052 & n3055;
  assign n3127 = ~n3059 & n3062;
  assign n3128 = ~n3056 & n3127;
  assign n3129 = ~n3126 & ~n3128;
  assign n3130 = ~n3126 & ~n3127;
  assign n3131 = n4897 & ~n3130;
  assign n3132 = n3049 & ~n3129;
  assign n3133 = n3125 & ~n4901;
  assign n3134 = ~n3063 & ~n3120;
  assign n3135 = n3130 & ~n3134;
  assign n3136 = n4897 & ~n3135;
  assign n3137 = n3125 & ~n3136;
  assign n3138 = ~n3121 & n3133;
  assign n3139 = ~n3109 & ~n3123;
  assign n3140 = ~n4901 & n3139;
  assign n3141 = ~n3121 & n3140;
  assign n3142 = ~n3124 & n3141;
  assign n3143 = ~n3109 & n4902;
  assign n3144 = pi67  & ~n4767;
  assign n3145 = pi195  & n4767;
  assign n3146 = ~n3144 & ~n3145;
  assign n3147 = pi323  & ~n4851;
  assign n3148 = pi451  & n4851;
  assign n3149 = ~n3147 & ~n3148;
  assign n3150 = n3146 & ~n3149;
  assign n3151 = pi322  & ~n4851;
  assign n3152 = pi450  & n4851;
  assign n3153 = ~n3151 & ~n3152;
  assign n3154 = pi66  & ~n4767;
  assign n3155 = pi194  & n4767;
  assign n3156 = ~n3154 & ~n3155;
  assign n3157 = ~n3153 & n3156;
  assign n3158 = ~n3150 & ~n3157;
  assign n3159 = pi65  & ~n4767;
  assign n3160 = pi193  & n4767;
  assign n3161 = ~n3159 & ~n3160;
  assign n3162 = pi321  & ~n4851;
  assign n3163 = pi449  & n4851;
  assign n3164 = ~n3162 & ~n3163;
  assign n3165 = n3161 & ~n3164;
  assign n3166 = pi320  & ~n4851;
  assign n3167 = pi448  & n4851;
  assign n3168 = ~n3166 & ~n3167;
  assign n3169 = pi64  & ~n4767;
  assign n3170 = pi192  & n4767;
  assign n3171 = ~n3169 & ~n3170;
  assign n3172 = ~n3168 & n3171;
  assign n3173 = ~n3165 & ~n3172;
  assign n3174 = n3158 & n3173;
  assign n3175 = ~n4903 & ~n3165;
  assign n3176 = ~n3172 & n3175;
  assign n3177 = n3158 & n3176;
  assign n3178 = ~n4903 & n3174;
  assign n3179 = ~n3146 & n3149;
  assign n3180 = n3168 & ~n3171;
  assign n3181 = ~n3165 & n3168;
  assign n3182 = ~n3171 & n3181;
  assign n3183 = ~n3165 & n3180;
  assign n3184 = ~n3161 & n3164;
  assign n3185 = n3153 & ~n3156;
  assign n3186 = ~n3184 & ~n3185;
  assign n3187 = ~n4905 & ~n3184;
  assign n3188 = ~n3185 & n3187;
  assign n3189 = ~n4905 & n3186;
  assign n3190 = n3158 & ~n4906;
  assign n3191 = ~n3179 & ~n3190;
  assign n3192 = ~n4904 & n3191;
  assign n3193 = pi71  & ~n4767;
  assign n3194 = pi199  & n4767;
  assign n3195 = ~n3193 & ~n3194;
  assign n3196 = pi327  & ~n4851;
  assign n3197 = pi455  & n4851;
  assign n3198 = ~n3196 & ~n3197;
  assign n3199 = n3195 & ~n3198;
  assign n3200 = pi326  & ~n4851;
  assign n3201 = pi454  & n4851;
  assign n3202 = ~n3200 & ~n3201;
  assign n3203 = pi70  & ~n4767;
  assign n3204 = pi198  & n4767;
  assign n3205 = ~n3203 & ~n3204;
  assign n3206 = ~n3202 & n3205;
  assign n3207 = ~n3199 & ~n3206;
  assign n3208 = pi69  & ~n4767;
  assign n3209 = pi197  & n4767;
  assign n3210 = ~n3208 & ~n3209;
  assign n3211 = pi325  & ~n4851;
  assign n3212 = pi453  & n4851;
  assign n3213 = ~n3211 & ~n3212;
  assign n3214 = n3210 & ~n3213;
  assign n3215 = pi324  & ~n4851;
  assign n3216 = pi452  & n4851;
  assign n3217 = ~n3215 & ~n3216;
  assign n3218 = pi68  & ~n4767;
  assign n3219 = pi196  & n4767;
  assign n3220 = ~n3218 & ~n3219;
  assign n3221 = ~n3217 & n3220;
  assign n3222 = ~n3214 & ~n3221;
  assign n3223 = n3207 & n3222;
  assign n3224 = ~n3192 & n3223;
  assign n3225 = ~n3195 & n3198;
  assign n3226 = n3217 & ~n3220;
  assign n3227 = ~n3214 & n3226;
  assign n3228 = n3202 & ~n3205;
  assign n3229 = ~n3210 & n3213;
  assign n3230 = ~n3228 & ~n3229;
  assign n3231 = ~n3227 & n3230;
  assign n3232 = n3207 & ~n3231;
  assign n3233 = ~n3227 & ~n3229;
  assign n3234 = n3207 & ~n3233;
  assign n3235 = ~n3199 & n3228;
  assign n3236 = ~n3225 & ~n3235;
  assign n3237 = ~n3234 & n3236;
  assign n3238 = ~n3225 & ~n3232;
  assign n3239 = ~n3224 & ~n3235;
  assign n3240 = ~n3234 & n3239;
  assign n3241 = ~n3225 & n3240;
  assign n3242 = ~n3224 & n4907;
  assign n3243 = pi75  & ~n4767;
  assign n3244 = pi203  & n4767;
  assign n3245 = ~n3243 & ~n3244;
  assign n3246 = pi331  & ~n4851;
  assign n3247 = pi459  & n4851;
  assign n3248 = ~n3246 & ~n3247;
  assign n3249 = n3245 & ~n3248;
  assign n3250 = pi330  & ~n4851;
  assign n3251 = pi458  & n4851;
  assign n3252 = ~n3250 & ~n3251;
  assign n3253 = pi74  & ~n4767;
  assign n3254 = pi202  & n4767;
  assign n3255 = ~n3253 & ~n3254;
  assign n3256 = ~n3252 & n3255;
  assign n3257 = ~n3249 & ~n3256;
  assign n3258 = pi73  & ~n4767;
  assign n3259 = pi201  & n4767;
  assign n3260 = ~n3258 & ~n3259;
  assign n3261 = pi329  & ~n4851;
  assign n3262 = pi457  & n4851;
  assign n3263 = ~n3261 & ~n3262;
  assign n3264 = n3260 & ~n3263;
  assign n3265 = pi328  & ~n4851;
  assign n3266 = pi456  & n4851;
  assign n3267 = ~n3265 & ~n3266;
  assign n3268 = pi72  & ~n4767;
  assign n3269 = pi200  & n4767;
  assign n3270 = ~n3268 & ~n3269;
  assign n3271 = ~n3267 & n3270;
  assign n3272 = ~n3264 & ~n3271;
  assign n3273 = n3257 & n3272;
  assign n3274 = ~n4908 & n3273;
  assign n3275 = ~n3245 & n3248;
  assign n3276 = n3267 & ~n3270;
  assign n3277 = ~n3264 & n3276;
  assign n3278 = ~n3260 & n3263;
  assign n3279 = n3252 & ~n3255;
  assign n3280 = ~n3278 & ~n3279;
  assign n3281 = ~n3277 & ~n3278;
  assign n3282 = ~n3279 & n3281;
  assign n3283 = ~n3277 & n3280;
  assign n3284 = n3257 & ~n4909;
  assign n3285 = ~n3275 & ~n3284;
  assign n3286 = ~n3274 & n3285;
  assign n3287 = pi79  & ~n4767;
  assign n3288 = pi207  & n4767;
  assign n3289 = ~n3287 & ~n3288;
  assign n3290 = pi335  & ~n4851;
  assign n3291 = pi463  & n4851;
  assign n3292 = ~n3290 & ~n3291;
  assign n3293 = n3289 & ~n3292;
  assign n3294 = pi334  & ~n4851;
  assign n3295 = pi462  & n4851;
  assign n3296 = ~n3294 & ~n3295;
  assign n3297 = pi78  & ~n4767;
  assign n3298 = pi206  & n4767;
  assign n3299 = ~n3297 & ~n3298;
  assign n3300 = ~n3296 & n3299;
  assign n3301 = ~n3293 & ~n3300;
  assign n3302 = pi77  & ~n4767;
  assign n3303 = pi205  & n4767;
  assign n3304 = ~n3302 & ~n3303;
  assign n3305 = pi333  & ~n4851;
  assign n3306 = pi461  & n4851;
  assign n3307 = ~n3305 & ~n3306;
  assign n3308 = n3304 & ~n3307;
  assign n3309 = pi332  & ~n4851;
  assign n3310 = pi460  & n4851;
  assign n3311 = ~n3309 & ~n3310;
  assign n3312 = pi76  & ~n4767;
  assign n3313 = pi204  & n4767;
  assign n3314 = ~n3312 & ~n3313;
  assign n3315 = ~n3311 & n3314;
  assign n3316 = ~n3308 & ~n3315;
  assign n3317 = n3301 & n3316;
  assign n3318 = ~n3286 & n3317;
  assign n3319 = ~n3289 & n3292;
  assign n3320 = n3311 & ~n3314;
  assign n3321 = ~n3308 & n3320;
  assign n3322 = n3296 & ~n3299;
  assign n3323 = ~n3304 & n3307;
  assign n3324 = ~n3322 & ~n3323;
  assign n3325 = ~n3321 & n3324;
  assign n3326 = n3301 & ~n3325;
  assign n3327 = ~n3321 & ~n3323;
  assign n3328 = n3301 & ~n3327;
  assign n3329 = ~n3293 & n3322;
  assign n3330 = ~n3319 & ~n3329;
  assign n3331 = ~n3328 & n3330;
  assign n3332 = ~n3319 & ~n3326;
  assign n3333 = ~n3318 & ~n3329;
  assign n3334 = ~n3328 & n3333;
  assign n3335 = ~n3319 & n3334;
  assign n3336 = ~n3318 & n4910;
  assign n3337 = pi83  & ~n4767;
  assign n3338 = pi211  & n4767;
  assign n3339 = ~n3337 & ~n3338;
  assign n3340 = pi339  & ~n4851;
  assign n3341 = pi467  & n4851;
  assign n3342 = ~n3340 & ~n3341;
  assign n3343 = n3339 & ~n3342;
  assign n3344 = pi338  & ~n4851;
  assign n3345 = pi466  & n4851;
  assign n3346 = ~n3344 & ~n3345;
  assign n3347 = pi82  & ~n4767;
  assign n3348 = pi210  & n4767;
  assign n3349 = ~n3347 & ~n3348;
  assign n3350 = ~n3346 & n3349;
  assign n3351 = ~n3343 & ~n3350;
  assign n3352 = pi81  & ~n4767;
  assign n3353 = pi209  & n4767;
  assign n3354 = ~n3352 & ~n3353;
  assign n3355 = pi337  & ~n4851;
  assign n3356 = pi465  & n4851;
  assign n3357 = ~n3355 & ~n3356;
  assign n3358 = n3354 & ~n3357;
  assign n3359 = pi336  & ~n4851;
  assign n3360 = pi464  & n4851;
  assign n3361 = ~n3359 & ~n3360;
  assign n3362 = pi80  & ~n4767;
  assign n3363 = pi208  & n4767;
  assign n3364 = ~n3362 & ~n3363;
  assign n3365 = ~n3361 & n3364;
  assign n3366 = ~n3358 & ~n3365;
  assign n3367 = n3351 & n3366;
  assign n3368 = ~n4911 & ~n3358;
  assign n3369 = n3351 & n3368;
  assign n3370 = ~n3365 & n3369;
  assign n3371 = ~n4911 & n3367;
  assign n3372 = ~n3339 & n3342;
  assign n3373 = n3361 & ~n3364;
  assign n3374 = ~n3358 & n3361;
  assign n3375 = ~n3364 & n3374;
  assign n3376 = ~n3358 & n3373;
  assign n3377 = ~n3354 & n3357;
  assign n3378 = n3346 & ~n3349;
  assign n3379 = ~n3377 & ~n3378;
  assign n3380 = ~n4913 & ~n3377;
  assign n3381 = ~n3378 & n3380;
  assign n3382 = ~n4913 & n3379;
  assign n3383 = n3351 & ~n4914;
  assign n3384 = ~n3372 & ~n3383;
  assign n3385 = ~n4912 & n3384;
  assign n3386 = pi87  & ~n4767;
  assign n3387 = pi215  & n4767;
  assign n3388 = ~n3386 & ~n3387;
  assign n3389 = pi343  & ~n4851;
  assign n3390 = pi471  & n4851;
  assign n3391 = ~n3389 & ~n3390;
  assign n3392 = n3388 & ~n3391;
  assign n3393 = pi342  & ~n4851;
  assign n3394 = pi470  & n4851;
  assign n3395 = ~n3393 & ~n3394;
  assign n3396 = pi86  & ~n4767;
  assign n3397 = pi214  & n4767;
  assign n3398 = ~n3396 & ~n3397;
  assign n3399 = ~n3395 & n3398;
  assign n3400 = ~n3392 & ~n3399;
  assign n3401 = pi85  & ~n4767;
  assign n3402 = pi213  & n4767;
  assign n3403 = ~n3401 & ~n3402;
  assign n3404 = pi341  & ~n4851;
  assign n3405 = pi469  & n4851;
  assign n3406 = ~n3404 & ~n3405;
  assign n3407 = n3403 & ~n3406;
  assign n3408 = pi340  & ~n4851;
  assign n3409 = pi468  & n4851;
  assign n3410 = ~n3408 & ~n3409;
  assign n3411 = pi84  & ~n4767;
  assign n3412 = pi212  & n4767;
  assign n3413 = ~n3411 & ~n3412;
  assign n3414 = ~n3410 & n3413;
  assign n3415 = ~n3407 & ~n3414;
  assign n3416 = n3400 & n3415;
  assign n3417 = ~n3385 & n3416;
  assign n3418 = ~n3388 & n3391;
  assign n3419 = n3410 & ~n3413;
  assign n3420 = ~n3407 & n3419;
  assign n3421 = n3395 & ~n3398;
  assign n3422 = ~n3403 & n3406;
  assign n3423 = ~n3421 & ~n3422;
  assign n3424 = ~n3420 & n3423;
  assign n3425 = n3400 & ~n3424;
  assign n3426 = ~n3420 & ~n3422;
  assign n3427 = n3400 & ~n3426;
  assign n3428 = ~n3392 & n3421;
  assign n3429 = ~n3418 & ~n3428;
  assign n3430 = ~n3427 & n3429;
  assign n3431 = ~n3418 & ~n3425;
  assign n3432 = ~n3417 & ~n3428;
  assign n3433 = ~n3427 & n3432;
  assign n3434 = ~n3418 & n3433;
  assign n3435 = ~n3417 & n4915;
  assign n3436 = pi91  & ~n4767;
  assign n3437 = pi219  & n4767;
  assign n3438 = ~n3436 & ~n3437;
  assign n3439 = pi347  & ~n4851;
  assign n3440 = pi475  & n4851;
  assign n3441 = ~n3439 & ~n3440;
  assign n3442 = n3438 & ~n3441;
  assign n3443 = pi346  & ~n4851;
  assign n3444 = pi474  & n4851;
  assign n3445 = ~n3443 & ~n3444;
  assign n3446 = pi90  & ~n4767;
  assign n3447 = pi218  & n4767;
  assign n3448 = ~n3446 & ~n3447;
  assign n3449 = ~n3445 & n3448;
  assign n3450 = ~n3442 & ~n3449;
  assign n3451 = pi89  & ~n4767;
  assign n3452 = pi217  & n4767;
  assign n3453 = ~n3451 & ~n3452;
  assign n3454 = pi345  & ~n4851;
  assign n3455 = pi473  & n4851;
  assign n3456 = ~n3454 & ~n3455;
  assign n3457 = n3453 & ~n3456;
  assign n3458 = pi344  & ~n4851;
  assign n3459 = pi472  & n4851;
  assign n3460 = ~n3458 & ~n3459;
  assign n3461 = pi88  & ~n4767;
  assign n3462 = pi216  & n4767;
  assign n3463 = ~n3461 & ~n3462;
  assign n3464 = ~n3460 & n3463;
  assign n3465 = ~n3457 & ~n3464;
  assign n3466 = n3450 & n3465;
  assign n3467 = ~n4916 & n3466;
  assign n3468 = ~n3438 & n3441;
  assign n3469 = n3460 & ~n3463;
  assign n3470 = ~n3457 & n3469;
  assign n3471 = ~n3453 & n3456;
  assign n3472 = n3445 & ~n3448;
  assign n3473 = ~n3471 & ~n3472;
  assign n3474 = ~n3470 & ~n3471;
  assign n3475 = ~n3472 & n3474;
  assign n3476 = ~n3470 & n3473;
  assign n3477 = n3450 & ~n4917;
  assign n3478 = ~n3468 & ~n3477;
  assign n3479 = ~n3467 & n3478;
  assign n3480 = pi95  & ~n4767;
  assign n3481 = pi223  & n4767;
  assign n3482 = ~n3480 & ~n3481;
  assign n3483 = pi351  & ~n4851;
  assign n3484 = pi479  & n4851;
  assign n3485 = ~n3483 & ~n3484;
  assign n3486 = n3482 & ~n3485;
  assign n3487 = pi350  & ~n4851;
  assign n3488 = pi478  & n4851;
  assign n3489 = ~n3487 & ~n3488;
  assign n3490 = pi94  & ~n4767;
  assign n3491 = pi222  & n4767;
  assign n3492 = ~n3490 & ~n3491;
  assign n3493 = ~n3489 & n3492;
  assign n3494 = ~n3486 & ~n3493;
  assign n3495 = pi93  & ~n4767;
  assign n3496 = pi221  & n4767;
  assign n3497 = ~n3495 & ~n3496;
  assign n3498 = pi349  & ~n4851;
  assign n3499 = pi477  & n4851;
  assign n3500 = ~n3498 & ~n3499;
  assign n3501 = n3497 & ~n3500;
  assign n3502 = pi348  & ~n4851;
  assign n3503 = pi476  & n4851;
  assign n3504 = ~n3502 & ~n3503;
  assign n3505 = pi92  & ~n4767;
  assign n3506 = pi220  & n4767;
  assign n3507 = ~n3505 & ~n3506;
  assign n3508 = ~n3504 & n3507;
  assign n3509 = ~n3501 & ~n3508;
  assign n3510 = n3494 & n3509;
  assign n3511 = ~n3479 & n3510;
  assign n3512 = ~n3482 & n3485;
  assign n3513 = n3504 & ~n3507;
  assign n3514 = ~n3501 & n3513;
  assign n3515 = n3489 & ~n3492;
  assign n3516 = ~n3497 & n3500;
  assign n3517 = ~n3515 & ~n3516;
  assign n3518 = ~n3514 & n3517;
  assign n3519 = n3494 & ~n3518;
  assign n3520 = ~n3514 & ~n3516;
  assign n3521 = n3494 & ~n3520;
  assign n3522 = ~n3486 & n3515;
  assign n3523 = ~n3512 & ~n3522;
  assign n3524 = ~n3521 & n3523;
  assign n3525 = ~n3512 & ~n3519;
  assign n3526 = ~n3511 & ~n3522;
  assign n3527 = ~n3521 & n3526;
  assign n3528 = ~n3512 & n3527;
  assign n3529 = ~n3511 & n4918;
  assign n3530 = pi99  & ~n4767;
  assign n3531 = pi227  & n4767;
  assign n3532 = ~n3530 & ~n3531;
  assign n3533 = pi355  & ~n4851;
  assign n3534 = pi483  & n4851;
  assign n3535 = ~n3533 & ~n3534;
  assign n3536 = n3532 & ~n3535;
  assign n3537 = pi354  & ~n4851;
  assign n3538 = pi482  & n4851;
  assign n3539 = ~n3537 & ~n3538;
  assign n3540 = pi98  & ~n4767;
  assign n3541 = pi226  & n4767;
  assign n3542 = ~n3540 & ~n3541;
  assign n3543 = ~n3539 & n3542;
  assign n3544 = ~n3536 & ~n3543;
  assign n3545 = pi97  & ~n4767;
  assign n3546 = pi225  & n4767;
  assign n3547 = ~n3545 & ~n3546;
  assign n3548 = pi353  & ~n4851;
  assign n3549 = pi481  & n4851;
  assign n3550 = ~n3548 & ~n3549;
  assign n3551 = n3547 & ~n3550;
  assign n3552 = pi352  & ~n4851;
  assign n3553 = pi480  & n4851;
  assign n3554 = ~n3552 & ~n3553;
  assign n3555 = pi96  & ~n4767;
  assign n3556 = pi224  & n4767;
  assign n3557 = ~n3555 & ~n3556;
  assign n3558 = ~n3554 & n3557;
  assign n3559 = ~n3551 & ~n3558;
  assign n3560 = n3544 & n3559;
  assign n3561 = ~n4919 & ~n3551;
  assign n3562 = n3544 & n3561;
  assign n3563 = ~n3558 & n3562;
  assign n3564 = ~n4919 & n3560;
  assign n3565 = ~n3532 & n3535;
  assign n3566 = n3554 & ~n3557;
  assign n3567 = ~n3551 & n3554;
  assign n3568 = ~n3557 & n3567;
  assign n3569 = ~n3551 & n3566;
  assign n3570 = ~n3547 & n3550;
  assign n3571 = n3539 & ~n3542;
  assign n3572 = ~n3570 & ~n3571;
  assign n3573 = ~n4921 & ~n3570;
  assign n3574 = ~n3571 & n3573;
  assign n3575 = ~n4921 & n3572;
  assign n3576 = n3544 & ~n4922;
  assign n3577 = ~n3565 & ~n3576;
  assign n3578 = ~n4920 & n3577;
  assign n3579 = pi103  & ~n4767;
  assign n3580 = pi231  & n4767;
  assign n3581 = ~n3579 & ~n3580;
  assign n3582 = pi359  & ~n4851;
  assign n3583 = pi487  & n4851;
  assign n3584 = ~n3582 & ~n3583;
  assign n3585 = n3581 & ~n3584;
  assign n3586 = pi358  & ~n4851;
  assign n3587 = pi486  & n4851;
  assign n3588 = ~n3586 & ~n3587;
  assign n3589 = pi102  & ~n4767;
  assign n3590 = pi230  & n4767;
  assign n3591 = ~n3589 & ~n3590;
  assign n3592 = ~n3588 & n3591;
  assign n3593 = ~n3585 & ~n3592;
  assign n3594 = pi101  & ~n4767;
  assign n3595 = pi229  & n4767;
  assign n3596 = ~n3594 & ~n3595;
  assign n3597 = pi357  & ~n4851;
  assign n3598 = pi485  & n4851;
  assign n3599 = ~n3597 & ~n3598;
  assign n3600 = n3596 & ~n3599;
  assign n3601 = pi356  & ~n4851;
  assign n3602 = pi484  & n4851;
  assign n3603 = ~n3601 & ~n3602;
  assign n3604 = pi100  & ~n4767;
  assign n3605 = pi228  & n4767;
  assign n3606 = ~n3604 & ~n3605;
  assign n3607 = ~n3603 & n3606;
  assign n3608 = ~n3600 & ~n3607;
  assign n3609 = n3593 & n3608;
  assign n3610 = ~n3578 & n3609;
  assign n3611 = ~n3581 & n3584;
  assign n3612 = n3603 & ~n3606;
  assign n3613 = ~n3600 & n3612;
  assign n3614 = n3588 & ~n3591;
  assign n3615 = ~n3596 & n3599;
  assign n3616 = ~n3614 & ~n3615;
  assign n3617 = ~n3613 & n3616;
  assign n3618 = n3593 & ~n3617;
  assign n3619 = ~n3613 & ~n3615;
  assign n3620 = n3593 & ~n3619;
  assign n3621 = ~n3585 & n3614;
  assign n3622 = ~n3611 & ~n3621;
  assign n3623 = ~n3620 & n3622;
  assign n3624 = ~n3611 & ~n3618;
  assign n3625 = ~n3610 & ~n3621;
  assign n3626 = ~n3620 & n3625;
  assign n3627 = ~n3611 & n3626;
  assign n3628 = ~n3610 & n4923;
  assign n3629 = pi107  & ~n4767;
  assign n3630 = pi235  & n4767;
  assign n3631 = ~n3629 & ~n3630;
  assign n3632 = pi363  & ~n4851;
  assign n3633 = pi491  & n4851;
  assign n3634 = ~n3632 & ~n3633;
  assign n3635 = n3631 & ~n3634;
  assign n3636 = pi362  & ~n4851;
  assign n3637 = pi490  & n4851;
  assign n3638 = ~n3636 & ~n3637;
  assign n3639 = pi106  & ~n4767;
  assign n3640 = pi234  & n4767;
  assign n3641 = ~n3639 & ~n3640;
  assign n3642 = ~n3638 & n3641;
  assign n3643 = ~n3635 & ~n3642;
  assign n3644 = pi105  & ~n4767;
  assign n3645 = pi233  & n4767;
  assign n3646 = ~n3644 & ~n3645;
  assign n3647 = pi361  & ~n4851;
  assign n3648 = pi489  & n4851;
  assign n3649 = ~n3647 & ~n3648;
  assign n3650 = n3646 & ~n3649;
  assign n3651 = pi360  & ~n4851;
  assign n3652 = pi488  & n4851;
  assign n3653 = ~n3651 & ~n3652;
  assign n3654 = pi104  & ~n4767;
  assign n3655 = pi232  & n4767;
  assign n3656 = ~n3654 & ~n3655;
  assign n3657 = ~n3653 & n3656;
  assign n3658 = ~n3650 & ~n3657;
  assign n3659 = n3643 & n3658;
  assign n3660 = ~n4924 & n3659;
  assign n3661 = ~n3631 & n3634;
  assign n3662 = n3653 & ~n3656;
  assign n3663 = ~n3650 & n3662;
  assign n3664 = ~n3646 & n3649;
  assign n3665 = n3638 & ~n3641;
  assign n3666 = ~n3664 & ~n3665;
  assign n3667 = ~n3663 & ~n3664;
  assign n3668 = ~n3665 & n3667;
  assign n3669 = ~n3663 & n3666;
  assign n3670 = n3643 & ~n4925;
  assign n3671 = ~n3661 & ~n3670;
  assign n3672 = ~n3660 & n3671;
  assign n3673 = pi111  & ~n4767;
  assign n3674 = pi239  & n4767;
  assign n3675 = ~n3673 & ~n3674;
  assign n3676 = pi367  & ~n4851;
  assign n3677 = pi495  & n4851;
  assign n3678 = ~n3676 & ~n3677;
  assign n3679 = n3675 & ~n3678;
  assign n3680 = pi366  & ~n4851;
  assign n3681 = pi494  & n4851;
  assign n3682 = ~n3680 & ~n3681;
  assign n3683 = pi110  & ~n4767;
  assign n3684 = pi238  & n4767;
  assign n3685 = ~n3683 & ~n3684;
  assign n3686 = ~n3682 & n3685;
  assign n3687 = ~n3679 & ~n3686;
  assign n3688 = pi109  & ~n4767;
  assign n3689 = pi237  & n4767;
  assign n3690 = ~n3688 & ~n3689;
  assign n3691 = pi365  & ~n4851;
  assign n3692 = pi493  & n4851;
  assign n3693 = ~n3691 & ~n3692;
  assign n3694 = n3690 & ~n3693;
  assign n3695 = pi364  & ~n4851;
  assign n3696 = pi492  & n4851;
  assign n3697 = ~n3695 & ~n3696;
  assign n3698 = pi108  & ~n4767;
  assign n3699 = pi236  & n4767;
  assign n3700 = ~n3698 & ~n3699;
  assign n3701 = ~n3697 & n3700;
  assign n3702 = ~n3694 & ~n3701;
  assign n3703 = n3687 & n3702;
  assign n3704 = ~n3672 & n3703;
  assign n3705 = ~n3675 & n3678;
  assign n3706 = n3697 & ~n3700;
  assign n3707 = ~n3694 & n3706;
  assign n3708 = n3682 & ~n3685;
  assign n3709 = ~n3690 & n3693;
  assign n3710 = ~n3708 & ~n3709;
  assign n3711 = ~n3707 & n3710;
  assign n3712 = n3687 & ~n3711;
  assign n3713 = ~n3707 & ~n3709;
  assign n3714 = n3687 & ~n3713;
  assign n3715 = ~n3679 & n3708;
  assign n3716 = ~n3705 & ~n3715;
  assign n3717 = ~n3714 & n3716;
  assign n3718 = ~n3705 & ~n3712;
  assign n3719 = ~n3704 & ~n3715;
  assign n3720 = ~n3714 & n3719;
  assign n3721 = ~n3705 & n3720;
  assign n3722 = ~n3704 & n4926;
  assign n3723 = pi115  & ~n4767;
  assign n3724 = pi243  & n4767;
  assign n3725 = ~n3723 & ~n3724;
  assign n3726 = pi371  & ~n4851;
  assign n3727 = pi499  & n4851;
  assign n3728 = ~n3726 & ~n3727;
  assign n3729 = n3725 & ~n3728;
  assign n3730 = pi370  & ~n4851;
  assign n3731 = pi498  & n4851;
  assign n3732 = ~n3730 & ~n3731;
  assign n3733 = pi114  & ~n4767;
  assign n3734 = pi242  & n4767;
  assign n3735 = ~n3733 & ~n3734;
  assign n3736 = ~n3732 & n3735;
  assign n3737 = ~n3729 & ~n3736;
  assign n3738 = pi113  & ~n4767;
  assign n3739 = pi241  & n4767;
  assign n3740 = ~n3738 & ~n3739;
  assign n3741 = pi369  & ~n4851;
  assign n3742 = pi497  & n4851;
  assign n3743 = ~n3741 & ~n3742;
  assign n3744 = n3740 & ~n3743;
  assign n3745 = pi368  & ~n4851;
  assign n3746 = pi496  & n4851;
  assign n3747 = ~n3745 & ~n3746;
  assign n3748 = pi112  & ~n4767;
  assign n3749 = pi240  & n4767;
  assign n3750 = ~n3748 & ~n3749;
  assign n3751 = ~n3747 & n3750;
  assign n3752 = ~n3744 & ~n3751;
  assign n3753 = n3737 & n3752;
  assign n3754 = ~n4927 & ~n3744;
  assign n3755 = n3737 & n3754;
  assign n3756 = ~n3751 & n3755;
  assign n3757 = ~n4927 & n3753;
  assign n3758 = ~n3725 & n3728;
  assign n3759 = n3747 & ~n3750;
  assign n3760 = ~n3744 & n3747;
  assign n3761 = ~n3750 & n3760;
  assign n3762 = ~n3744 & n3759;
  assign n3763 = ~n3740 & n3743;
  assign n3764 = n3732 & ~n3735;
  assign n3765 = ~n3763 & ~n3764;
  assign n3766 = ~n4929 & ~n3763;
  assign n3767 = ~n3764 & n3766;
  assign n3768 = ~n4929 & n3765;
  assign n3769 = n3737 & ~n4930;
  assign n3770 = ~n3758 & ~n3769;
  assign n3771 = ~n4928 & n3770;
  assign n3772 = pi119  & ~n4767;
  assign n3773 = pi247  & n4767;
  assign n3774 = ~n3772 & ~n3773;
  assign n3775 = pi375  & ~n4851;
  assign n3776 = pi503  & n4851;
  assign n3777 = ~n3775 & ~n3776;
  assign n3778 = n3774 & ~n3777;
  assign n3779 = pi374  & ~n4851;
  assign n3780 = pi502  & n4851;
  assign n3781 = ~n3779 & ~n3780;
  assign n3782 = pi118  & ~n4767;
  assign n3783 = pi246  & n4767;
  assign n3784 = ~n3782 & ~n3783;
  assign n3785 = ~n3781 & n3784;
  assign n3786 = ~n3778 & ~n3785;
  assign n3787 = pi117  & ~n4767;
  assign n3788 = pi245  & n4767;
  assign n3789 = ~n3787 & ~n3788;
  assign n3790 = pi373  & ~n4851;
  assign n3791 = pi501  & n4851;
  assign n3792 = ~n3790 & ~n3791;
  assign n3793 = n3789 & ~n3792;
  assign n3794 = pi372  & ~n4851;
  assign n3795 = pi500  & n4851;
  assign n3796 = ~n3794 & ~n3795;
  assign n3797 = pi116  & ~n4767;
  assign n3798 = pi244  & n4767;
  assign n3799 = ~n3797 & ~n3798;
  assign n3800 = ~n3796 & n3799;
  assign n3801 = ~n3793 & ~n3800;
  assign n3802 = n3786 & n3801;
  assign n3803 = ~n3771 & n3802;
  assign n3804 = ~n3774 & n3777;
  assign n3805 = n3796 & ~n3799;
  assign n3806 = ~n3793 & n3796;
  assign n3807 = ~n3799 & n3806;
  assign n3808 = ~n3793 & n3805;
  assign n3809 = n3781 & ~n3784;
  assign n3810 = ~n3789 & n3792;
  assign n3811 = ~n3809 & ~n3810;
  assign n3812 = ~n4931 & n3811;
  assign n3813 = n3786 & ~n3812;
  assign n3814 = ~n4931 & ~n3810;
  assign n3815 = n3786 & ~n3814;
  assign n3816 = ~n3778 & n3809;
  assign n3817 = ~n3804 & ~n3816;
  assign n3818 = ~n3815 & n3817;
  assign n3819 = ~n3804 & ~n3813;
  assign n3820 = ~n3803 & ~n3816;
  assign n3821 = ~n3815 & n3820;
  assign n3822 = ~n3804 & n3821;
  assign n3823 = ~n3803 & n4932;
  assign n3824 = pi123  & ~n4767;
  assign n3825 = pi251  & n4767;
  assign n3826 = ~n3824 & ~n3825;
  assign n3827 = pi379  & ~n4851;
  assign n3828 = pi507  & n4851;
  assign n3829 = ~n3827 & ~n3828;
  assign n3830 = n3826 & ~n3829;
  assign n3831 = pi378  & ~n4851;
  assign n3832 = pi506  & n4851;
  assign n3833 = ~n3831 & ~n3832;
  assign n3834 = pi122  & ~n4767;
  assign n3835 = pi250  & n4767;
  assign n3836 = ~n3834 & ~n3835;
  assign n3837 = ~n3833 & n3836;
  assign n3838 = ~n3830 & ~n3837;
  assign n3839 = pi121  & ~n4767;
  assign n3840 = pi249  & n4767;
  assign n3841 = ~n3839 & ~n3840;
  assign n3842 = pi377  & ~n4851;
  assign n3843 = pi505  & n4851;
  assign n3844 = ~n3842 & ~n3843;
  assign n3845 = n3841 & ~n3844;
  assign n3846 = pi376  & ~n4851;
  assign n3847 = pi504  & n4851;
  assign n3848 = ~n3846 & ~n3847;
  assign n3849 = pi120  & ~n4767;
  assign n3850 = pi248  & n4767;
  assign n3851 = ~n3849 & ~n3850;
  assign n3852 = ~n3848 & n3851;
  assign n3853 = ~n3845 & ~n3852;
  assign n3854 = n3838 & n3853;
  assign n3855 = ~n4933 & n3854;
  assign n3856 = ~n3826 & n3829;
  assign n3857 = n3848 & ~n3851;
  assign n3858 = ~n3845 & n3848;
  assign n3859 = ~n3851 & n3858;
  assign n3860 = ~n3845 & n3857;
  assign n3861 = ~n3841 & n3844;
  assign n3862 = n3833 & ~n3836;
  assign n3863 = ~n3861 & ~n3862;
  assign n3864 = ~n4934 & ~n3861;
  assign n3865 = ~n3862 & n3864;
  assign n3866 = ~n4934 & n3863;
  assign n3867 = n3838 & ~n4935;
  assign n3868 = ~n3856 & ~n3867;
  assign n3869 = ~n3855 & n3868;
  assign n3870 = pi126  & ~n4767;
  assign n3871 = pi254  & n4767;
  assign n3872 = ~n3870 & ~n3871;
  assign n3873 = pi382  & ~n4851;
  assign n3874 = pi510  & n4851;
  assign n3875 = ~n3873 & ~n3874;
  assign n3876 = n3872 & ~n3875;
  assign n3877 = pi125  & ~n4767;
  assign n3878 = pi253  & n4767;
  assign n3879 = ~n3877 & ~n3878;
  assign n3880 = pi381  & ~n4851;
  assign n3881 = pi509  & n4851;
  assign n3882 = ~n3880 & ~n3881;
  assign n3883 = n3879 & ~n3882;
  assign n3884 = ~n3876 & ~n3883;
  assign n3885 = ~pi511  & ~n2275;
  assign n3886 = pi383  & ~n3885;
  assign n3887 = ~pi511  & n2285;
  assign n3888 = pi383  & ~n3887;
  assign n3889 = pi383  & pi511 ;
  assign n3890 = ~pi255  & ~n1450;
  assign n3891 = pi127  & ~n3890;
  assign n3892 = ~pi255  & n1460;
  assign n3893 = pi127  & ~n3892;
  assign n3894 = pi127  & pi255 ;
  assign n3895 = ~n4936 & n4937;
  assign n3896 = pi124  & ~n4767;
  assign n3897 = pi252  & n4767;
  assign n3898 = ~n3896 & ~n3897;
  assign n3899 = pi380  & ~n4851;
  assign n3900 = pi508  & n4851;
  assign n3901 = ~n3899 & ~n3900;
  assign n3902 = n3898 & ~n3901;
  assign n3903 = ~n3895 & ~n3902;
  assign n3904 = n3884 & ~n3895;
  assign n3905 = ~n3902 & n3904;
  assign n3906 = n3884 & n3903;
  assign n3907 = ~n3869 & n4938;
  assign n3908 = ~n3898 & n3901;
  assign n3909 = ~n3879 & n3882;
  assign n3910 = ~n3908 & ~n3909;
  assign n3911 = n3884 & ~n3910;
  assign n3912 = n4936 & ~n4937;
  assign n3913 = ~n3872 & n3875;
  assign n3914 = ~n3912 & ~n3913;
  assign n3915 = ~n3911 & n3914;
  assign n3916 = ~n3895 & ~n3915;
  assign n3917 = ~n3911 & ~n3913;
  assign n3918 = ~n3895 & ~n3917;
  assign n3919 = ~n3907 & ~n3918;
  assign n3920 = ~n3912 & n3919;
  assign n3921 = ~n3907 & ~n3916;
  assign n3922 = ~n2388 & po129 ;
  assign n3923 = ~n2391 & ~po129 ;
  assign n3924 = ~n3922 & ~n3923;
  assign n3925 = ~n2381 & ~po129 ;
  assign n3926 = ~n2384 & po129 ;
  assign n3927 = n2381 & ~po129 ;
  assign n3928 = n2384 & po129 ;
  assign n3929 = ~n3927 & ~n3928;
  assign n3930 = ~n3925 & ~n3926;
  assign n3931 = ~n2376 & po129 ;
  assign n3932 = ~n2373 & ~po129 ;
  assign n3933 = n2373 & ~po129 ;
  assign n3934 = n2376 & po129 ;
  assign n3935 = ~n3933 & ~n3934;
  assign n3936 = ~n3931 & ~n3932;
  assign n3937 = ~n2368 & po129 ;
  assign n3938 = ~n2365 & ~po129 ;
  assign n3939 = n2365 & ~po129 ;
  assign n3940 = n2368 & po129 ;
  assign n3941 = ~n3939 & ~n3940;
  assign n3942 = ~n3937 & ~n3938;
  assign n3943 = ~n2418 & po129 ;
  assign n3944 = ~n2362 & ~po129 ;
  assign n3945 = ~n3943 & ~n3944;
  assign n3946 = ~n2427 & po129 ;
  assign n3947 = ~n2424 & ~po129 ;
  assign n3948 = ~n3946 & ~n3947;
  assign n3949 = n2358 & ~po129 ;
  assign n3950 = n2355 & po129 ;
  assign n3951 = ~n2355 & po129 ;
  assign n3952 = ~n2358 & ~po129 ;
  assign n3953 = ~n3951 & ~n3952;
  assign n3954 = ~n3949 & ~n3950;
  assign n3955 = ~n2453 & po129 ;
  assign n3956 = ~n2450 & ~po129 ;
  assign n3957 = n2450 & ~po129 ;
  assign n3958 = n2453 & po129 ;
  assign n3959 = ~n3957 & ~n3958;
  assign n3960 = ~n3955 & ~n3956;
  assign n3961 = ~n2471 & po129 ;
  assign n3962 = ~n2468 & ~po129 ;
  assign n3963 = n2468 & ~po129 ;
  assign n3964 = n2471 & po129 ;
  assign n3965 = ~n3963 & ~n3964;
  assign n3966 = ~n3961 & ~n3962;
  assign n3967 = ~n2482 & po129 ;
  assign n3968 = ~n2479 & ~po129 ;
  assign n3969 = n2479 & ~po129 ;
  assign n3970 = n2482 & po129 ;
  assign n3971 = ~n3969 & ~n3970;
  assign n3972 = ~n3967 & ~n3968;
  assign n3973 = ~n2351 & po129 ;
  assign n3974 = ~n2348 & ~po129 ;
  assign n3975 = n2348 & ~po129 ;
  assign n3976 = n2351 & po129 ;
  assign n3977 = ~n3975 & ~n3976;
  assign n3978 = ~n3973 & ~n3974;
  assign n3979 = ~n2507 & po129 ;
  assign n3980 = ~n2345 & ~po129 ;
  assign n3981 = n2345 & ~po129 ;
  assign n3982 = n2507 & po129 ;
  assign n3983 = ~n3981 & ~n3982;
  assign n3984 = ~n3979 & ~n3980;
  assign n3985 = ~n2341 & po129 ;
  assign n3986 = ~n2338 & ~po129 ;
  assign n3987 = n2338 & ~po129 ;
  assign n3988 = n2341 & po129 ;
  assign n3989 = ~n3987 & ~n3988;
  assign n3990 = ~n3985 & ~n3986;
  assign n3991 = ~n2334 & po129 ;
  assign n3992 = ~n2331 & ~po129 ;
  assign n3993 = n2331 & ~po129 ;
  assign n3994 = n2334 & po129 ;
  assign n3995 = ~n3993 & ~n3994;
  assign n3996 = ~n3991 & ~n3992;
  assign n3997 = ~n2527 & po129 ;
  assign n3998 = ~n2524 & ~po129 ;
  assign n3999 = n2524 & ~po129 ;
  assign n4000 = n2527 & po129 ;
  assign n4001 = ~n3999 & ~n4000;
  assign n4002 = ~n3997 & ~n3998;
  assign n4003 = ~n2537 & po129 ;
  assign n4004 = ~n2534 & ~po129 ;
  assign n4005 = n2534 & ~po129 ;
  assign n4006 = n2537 & po129 ;
  assign n4007 = ~n4005 & ~n4006;
  assign n4008 = ~n4003 & ~n4004;
  assign n4009 = ~n2551 & po129 ;
  assign n4010 = ~n2548 & ~po129 ;
  assign n4011 = n2548 & ~po129 ;
  assign n4012 = n2551 & po129 ;
  assign n4013 = ~n4011 & ~n4012;
  assign n4014 = ~n4009 & ~n4010;
  assign n4015 = ~n2327 & po129 ;
  assign n4016 = ~n2324 & ~po129 ;
  assign n4017 = n2324 & ~po129 ;
  assign n4018 = n2327 & po129 ;
  assign n4019 = ~n4017 & ~n4018;
  assign n4020 = ~n4015 & ~n4016;
  assign n4021 = ~n2572 & po129 ;
  assign n4022 = ~n2321 & ~po129 ;
  assign n4023 = n2321 & ~po129 ;
  assign n4024 = n2572 & po129 ;
  assign n4025 = ~n4023 & ~n4024;
  assign n4026 = ~n4021 & ~n4022;
  assign n4027 = ~n2317 & po129 ;
  assign n4028 = ~n2314 & ~po129 ;
  assign n4029 = n2314 & ~po129 ;
  assign n4030 = n2317 & po129 ;
  assign n4031 = ~n4029 & ~n4030;
  assign n4032 = ~n4027 & ~n4028;
  assign n4033 = ~n2587 & po129 ;
  assign n4034 = ~n2311 & ~po129 ;
  assign n4035 = n2311 & ~po129 ;
  assign n4036 = n2587 & po129 ;
  assign n4037 = ~n4035 & ~n4036;
  assign n4038 = ~n4033 & ~n4034;
  assign n4039 = ~n2595 & po129 ;
  assign n4040 = ~n2592 & ~po129 ;
  assign n4041 = n2592 & ~po129 ;
  assign n4042 = n2595 & po129 ;
  assign n4043 = ~n4041 & ~n4042;
  assign n4044 = ~n4039 & ~n4040;
  assign n4045 = ~n2611 & po129 ;
  assign n4046 = ~n2608 & ~po129 ;
  assign n4047 = n2608 & ~po129 ;
  assign n4048 = n2611 & po129 ;
  assign n4049 = ~n4047 & ~n4048;
  assign n4050 = ~n4045 & ~n4046;
  assign n4051 = ~n2621 & po129 ;
  assign n4052 = ~n2618 & ~po129 ;
  assign n4053 = n2618 & ~po129 ;
  assign n4054 = n2621 & po129 ;
  assign n4055 = ~n4053 & ~n4054;
  assign n4056 = ~n4051 & ~n4052;
  assign n4057 = ~n2635 & po129 ;
  assign n4058 = ~n2632 & ~po129 ;
  assign n4059 = n2632 & ~po129 ;
  assign n4060 = n2635 & po129 ;
  assign n4061 = ~n4059 & ~n4060;
  assign n4062 = ~n4057 & ~n4058;
  assign n4063 = ~n2307 & po129 ;
  assign n4064 = ~n2304 & ~po129 ;
  assign n4065 = n2304 & ~po129 ;
  assign n4066 = n2307 & po129 ;
  assign n4067 = ~n4065 & ~n4066;
  assign n4068 = ~n4063 & ~n4064;
  assign n4069 = ~n2656 & po129 ;
  assign n4070 = ~n2301 & ~po129 ;
  assign n4071 = n2301 & ~po129 ;
  assign n4072 = n2656 & po129 ;
  assign n4073 = ~n4071 & ~n4072;
  assign n4074 = ~n4069 & ~n4070;
  assign n4075 = ~n2297 & po129 ;
  assign n4076 = ~n2294 & ~po129 ;
  assign n4077 = n2294 & ~po129 ;
  assign n4078 = n2297 & po129 ;
  assign n4079 = ~n4077 & ~n4078;
  assign n4080 = ~n4075 & ~n4076;
  assign n4081 = ~n2290 & po129 ;
  assign n4082 = ~n1465 & ~po129 ;
  assign n4083 = n1465 & ~po129 ;
  assign n4084 = n2290 & po129 ;
  assign n4085 = ~n4083 & ~n4084;
  assign n4086 = ~n4081 & ~n4082;
  assign n4087 = ~n2676 & po129 ;
  assign n4088 = ~n2673 & ~po129 ;
  assign n4089 = n2673 & ~po129 ;
  assign n4090 = n2676 & po129 ;
  assign n4091 = ~n4089 & ~n4090;
  assign n4092 = ~n4087 & ~n4088;
  assign n4093 = ~n2686 & po129 ;
  assign n4094 = ~n2683 & ~po129 ;
  assign n4095 = n2683 & ~po129 ;
  assign n4096 = n2686 & po129 ;
  assign n4097 = ~n4095 & ~n4096;
  assign n4098 = ~n4093 & ~n4094;
  assign n4099 = ~n2700 & po129 ;
  assign n4100 = ~n2697 & ~po129 ;
  assign n4101 = n2697 & ~po129 ;
  assign n4102 = n2700 & po129 ;
  assign n4103 = ~n4101 & ~n4102;
  assign n4104 = ~n4099 & ~n4100;
  assign n4105 = ~n2756 & po129 ;
  assign n4106 = ~n2759 & ~po129 ;
  assign n4107 = n2759 & ~po129 ;
  assign n4108 = n2756 & po129 ;
  assign n4109 = ~n4107 & ~n4108;
  assign n4110 = ~n4105 & ~n4106;
  assign n4111 = ~n2741 & po129 ;
  assign n4112 = ~n2738 & ~po129 ;
  assign n4113 = n2738 & ~po129 ;
  assign n4114 = n2741 & po129 ;
  assign n4115 = ~n4113 & ~n4114;
  assign n4116 = ~n4111 & ~n4112;
  assign n4117 = ~n2731 & po129 ;
  assign n4118 = ~n2734 & ~po129 ;
  assign n4119 = n2734 & ~po129 ;
  assign n4120 = n2731 & po129 ;
  assign n4121 = ~n4119 & ~n4120;
  assign n4122 = ~n4117 & ~n4118;
  assign n4123 = ~n2748 & po129 ;
  assign n4124 = ~n2745 & ~po129 ;
  assign n4125 = n2745 & ~po129 ;
  assign n4126 = n2748 & po129 ;
  assign n4127 = ~n4125 & ~n4126;
  assign n4128 = ~n4123 & ~n4124;
  assign n4129 = ~n2766 & po129 ;
  assign n4130 = ~n2763 & ~po129 ;
  assign n4131 = n2763 & ~po129 ;
  assign n4132 = n2766 & po129 ;
  assign n4133 = ~n4131 & ~n4132;
  assign n4134 = ~n4129 & ~n4130;
  assign n4135 = ~n2716 & po129 ;
  assign n4136 = ~n2713 & ~po129 ;
  assign n4137 = n2713 & ~po129 ;
  assign n4138 = n2716 & po129 ;
  assign n4139 = ~n4137 & ~n4138;
  assign n4140 = ~n4135 & ~n4136;
  assign n4141 = ~n2706 & po129 ;
  assign n4142 = ~n2709 & ~po129 ;
  assign n4143 = n2709 & ~po129 ;
  assign n4144 = n2706 & po129 ;
  assign n4145 = ~n4143 & ~n4144;
  assign n4146 = ~n4141 & ~n4142;
  assign n4147 = ~n2723 & po129 ;
  assign n4148 = ~n2720 & ~po129 ;
  assign n4149 = n2720 & ~po129 ;
  assign n4150 = n2723 & po129 ;
  assign n4151 = ~n4149 & ~n4150;
  assign n4152 = ~n4147 & ~n4148;
  assign n4153 = ~n2892 & po129 ;
  assign n4154 = ~n2889 & ~po129 ;
  assign n4155 = n2889 & ~po129 ;
  assign n4156 = n2892 & po129 ;
  assign n4157 = ~n4155 & ~n4156;
  assign n4158 = ~n4153 & ~n4154;
  assign n4159 = ~n2885 & po129 ;
  assign n4160 = ~n2882 & ~po129 ;
  assign n4161 = n2882 & ~po129 ;
  assign n4162 = n2885 & po129 ;
  assign n4163 = ~n4161 & ~n4162;
  assign n4164 = ~n4159 & ~n4160;
  assign n4165 = ~n2877 & po129 ;
  assign n4166 = ~n2874 & ~po129 ;
  assign n4167 = n2874 & ~po129 ;
  assign n4168 = n2877 & po129 ;
  assign n4169 = ~n4167 & ~n4168;
  assign n4170 = ~n4165 & ~n4166;
  assign n4171 = ~n2870 & po129 ;
  assign n4172 = ~n2867 & ~po129 ;
  assign n4173 = n2867 & ~po129 ;
  assign n4174 = n2870 & po129 ;
  assign n4175 = ~n4173 & ~n4174;
  assign n4176 = ~n4171 & ~n4172;
  assign n4177 = ~n2856 & po129 ;
  assign n4178 = ~n2853 & ~po129 ;
  assign n4179 = n2853 & ~po129 ;
  assign n4180 = n2856 & po129 ;
  assign n4181 = ~n4179 & ~n4180;
  assign n4182 = ~n4177 & ~n4178;
  assign n4183 = ~n2849 & po129 ;
  assign n4184 = ~n2846 & ~po129 ;
  assign n4185 = n2846 & ~po129 ;
  assign n4186 = n2849 & po129 ;
  assign n4187 = ~n4185 & ~n4186;
  assign n4188 = ~n4183 & ~n4184;
  assign n4189 = ~n2831 & po129 ;
  assign n4190 = ~n2834 & ~po129 ;
  assign n4191 = n2834 & ~po129 ;
  assign n4192 = n2831 & po129 ;
  assign n4193 = ~n4191 & ~n4192;
  assign n4194 = ~n4189 & ~n4190;
  assign n4195 = ~n2841 & po129 ;
  assign n4196 = ~n2838 & ~po129 ;
  assign n4197 = n2838 & ~po129 ;
  assign n4198 = n2841 & po129 ;
  assign n4199 = ~n4197 & ~n4198;
  assign n4200 = ~n4195 & ~n4196;
  assign n4201 = ~n2994 & po129 ;
  assign n4202 = ~n2997 & ~po129 ;
  assign n4203 = n2997 & ~po129 ;
  assign n4204 = n2994 & po129 ;
  assign n4205 = ~n4203 & ~n4204;
  assign n4206 = ~n4201 & ~n4202;
  assign n4207 = ~n2979 & po129 ;
  assign n4208 = ~n2976 & ~po129 ;
  assign n4209 = n2976 & ~po129 ;
  assign n4210 = n2979 & po129 ;
  assign n4211 = ~n4209 & ~n4210;
  assign n4212 = ~n4207 & ~n4208;
  assign n4213 = ~n2969 & po129 ;
  assign n4214 = ~n2972 & ~po129 ;
  assign n4215 = n2972 & ~po129 ;
  assign n4216 = n2969 & po129 ;
  assign n4217 = ~n4215 & ~n4216;
  assign n4218 = ~n4213 & ~n4214;
  assign n4219 = ~n2986 & po129 ;
  assign n4220 = ~n2983 & ~po129 ;
  assign n4221 = n2983 & ~po129 ;
  assign n4222 = n2986 & po129 ;
  assign n4223 = ~n4221 & ~n4222;
  assign n4224 = ~n4219 & ~n4220;
  assign n4225 = ~n2960 & po129 ;
  assign n4226 = ~n2963 & ~po129 ;
  assign n4227 = n2963 & ~po129 ;
  assign n4228 = n2960 & po129 ;
  assign n4229 = ~n4227 & ~n4228;
  assign n4230 = ~n4225 & ~n4226;
  assign n4231 = ~n2956 & po129 ;
  assign n4232 = ~n2953 & ~po129 ;
  assign n4233 = n2953 & ~po129 ;
  assign n4234 = n2956 & po129 ;
  assign n4235 = ~n4233 & ~n4234;
  assign n4236 = ~n4231 & ~n4232;
  assign n4237 = ~n2945 & po129 ;
  assign n4238 = ~n2948 & ~po129 ;
  assign n4239 = n2948 & ~po129 ;
  assign n4240 = n2945 & po129 ;
  assign n4241 = ~n4239 & ~n4240;
  assign n4242 = ~n4237 & ~n4238;
  assign n4243 = ~n2941 & po129 ;
  assign n4244 = ~n2938 & ~po129 ;
  assign n4245 = n2938 & ~po129 ;
  assign n4246 = n2941 & po129 ;
  assign n4247 = ~n4245 & ~n4246;
  assign n4248 = ~n4243 & ~n4244;
  assign n4249 = ~n3098 & po129 ;
  assign n4250 = ~n3095 & ~po129 ;
  assign n4251 = n3095 & ~po129 ;
  assign n4252 = n3098 & po129 ;
  assign n4253 = ~n4251 & ~n4252;
  assign n4254 = ~n4249 & ~n4250;
  assign n4255 = ~n3091 & po129 ;
  assign n4256 = ~n3088 & ~po129 ;
  assign n4257 = n3088 & ~po129 ;
  assign n4258 = n3091 & po129 ;
  assign n4259 = ~n4257 & ~n4258;
  assign n4260 = ~n4255 & ~n4256;
  assign n4261 = ~n3083 & po129 ;
  assign n4262 = ~n3080 & ~po129 ;
  assign n4263 = n3080 & ~po129 ;
  assign n4264 = n3083 & po129 ;
  assign n4265 = ~n4263 & ~n4264;
  assign n4266 = ~n4261 & ~n4262;
  assign n4267 = ~n3076 & po129 ;
  assign n4268 = ~n3073 & ~po129 ;
  assign n4269 = n3073 & ~po129 ;
  assign n4270 = n3076 & po129 ;
  assign n4271 = ~n4269 & ~n4270;
  assign n4272 = ~n4267 & ~n4268;
  assign n4273 = ~n3062 & po129 ;
  assign n4274 = ~n3059 & ~po129 ;
  assign n4275 = n3059 & ~po129 ;
  assign n4276 = n3062 & po129 ;
  assign n4277 = ~n4275 & ~n4276;
  assign n4278 = ~n4273 & ~n4274;
  assign n4279 = ~n3055 & po129 ;
  assign n4280 = ~n3052 & ~po129 ;
  assign n4281 = n3052 & ~po129 ;
  assign n4282 = n3055 & po129 ;
  assign n4283 = ~n4281 & ~n4282;
  assign n4284 = ~n4279 & ~n4280;
  assign n4285 = ~n3037 & po129 ;
  assign n4286 = ~n3040 & ~po129 ;
  assign n4287 = n3040 & ~po129 ;
  assign n4288 = n3037 & po129 ;
  assign n4289 = ~n4287 & ~n4288;
  assign n4290 = ~n4285 & ~n4286;
  assign n4291 = ~n3047 & po129 ;
  assign n4292 = ~n3044 & ~po129 ;
  assign n4293 = n3044 & ~po129 ;
  assign n4294 = n3047 & po129 ;
  assign n4295 = ~n4293 & ~n4294;
  assign n4296 = ~n4291 & ~n4292;
  assign n4297 = ~n3168 & po129 ;
  assign n4298 = ~n3171 & ~po129 ;
  assign n4299 = n3171 & ~po129 ;
  assign n4300 = n3168 & po129 ;
  assign n4301 = ~n4299 & ~n4300;
  assign n4302 = ~n4297 & ~n4298;
  assign n4303 = ~n3164 & po129 ;
  assign n4304 = ~n3161 & ~po129 ;
  assign n4305 = n3161 & ~po129 ;
  assign n4306 = n3164 & po129 ;
  assign n4307 = ~n4305 & ~n4306;
  assign n4308 = ~n4303 & ~n4304;
  assign n4309 = ~n3153 & po129 ;
  assign n4310 = ~n3156 & ~po129 ;
  assign n4311 = n3156 & ~po129 ;
  assign n4312 = n3153 & po129 ;
  assign n4313 = ~n4311 & ~n4312;
  assign n4314 = ~n4309 & ~n4310;
  assign n4315 = ~n3149 & po129 ;
  assign n4316 = ~n3146 & ~po129 ;
  assign n4317 = n3146 & ~po129 ;
  assign n4318 = n3149 & po129 ;
  assign n4319 = ~n4317 & ~n4318;
  assign n4320 = ~n4315 & ~n4316;
  assign n4321 = ~n3217 & po129 ;
  assign n4322 = ~n3220 & ~po129 ;
  assign n4323 = n3220 & ~po129 ;
  assign n4324 = n3217 & po129 ;
  assign n4325 = ~n4323 & ~n4324;
  assign n4326 = ~n4321 & ~n4322;
  assign n4327 = ~n3213 & po129 ;
  assign n4328 = ~n3210 & ~po129 ;
  assign n4329 = n3210 & ~po129 ;
  assign n4330 = n3213 & po129 ;
  assign n4331 = ~n4329 & ~n4330;
  assign n4332 = ~n4327 & ~n4328;
  assign n4333 = ~n3202 & po129 ;
  assign n4334 = ~n3205 & ~po129 ;
  assign n4335 = n3205 & ~po129 ;
  assign n4336 = n3202 & po129 ;
  assign n4337 = ~n4335 & ~n4336;
  assign n4338 = ~n4333 & ~n4334;
  assign n4339 = ~n3198 & po129 ;
  assign n4340 = ~n3195 & ~po129 ;
  assign n4341 = n3195 & ~po129 ;
  assign n4342 = n3198 & po129 ;
  assign n4343 = ~n4341 & ~n4342;
  assign n4344 = ~n4339 & ~n4340;
  assign n4345 = ~n3267 & po129 ;
  assign n4346 = ~n3270 & ~po129 ;
  assign n4347 = n3270 & ~po129 ;
  assign n4348 = n3267 & po129 ;
  assign n4349 = ~n4347 & ~n4348;
  assign n4350 = ~n4345 & ~n4346;
  assign n4351 = ~n3263 & po129 ;
  assign n4352 = ~n3260 & ~po129 ;
  assign n4353 = n3260 & ~po129 ;
  assign n4354 = n3263 & po129 ;
  assign n4355 = ~n4353 & ~n4354;
  assign n4356 = ~n4351 & ~n4352;
  assign n4357 = ~n3252 & po129 ;
  assign n4358 = ~n3255 & ~po129 ;
  assign n4359 = n3255 & ~po129 ;
  assign n4360 = n3252 & po129 ;
  assign n4361 = ~n4359 & ~n4360;
  assign n4362 = ~n4357 & ~n4358;
  assign n4363 = ~n3248 & po129 ;
  assign n4364 = ~n3245 & ~po129 ;
  assign n4365 = n3245 & ~po129 ;
  assign n4366 = n3248 & po129 ;
  assign n4367 = ~n4365 & ~n4366;
  assign n4368 = ~n4363 & ~n4364;
  assign n4369 = ~n3311 & po129 ;
  assign n4370 = ~n3314 & ~po129 ;
  assign n4371 = n3314 & ~po129 ;
  assign n4372 = n3311 & po129 ;
  assign n4373 = ~n4371 & ~n4372;
  assign n4374 = ~n4369 & ~n4370;
  assign n4375 = ~n3307 & po129 ;
  assign n4376 = ~n3304 & ~po129 ;
  assign n4377 = n3304 & ~po129 ;
  assign n4378 = n3307 & po129 ;
  assign n4379 = ~n4377 & ~n4378;
  assign n4380 = ~n4375 & ~n4376;
  assign n4381 = ~n3296 & po129 ;
  assign n4382 = ~n3299 & ~po129 ;
  assign n4383 = n3299 & ~po129 ;
  assign n4384 = n3296 & po129 ;
  assign n4385 = ~n4383 & ~n4384;
  assign n4386 = ~n4381 & ~n4382;
  assign n4387 = ~n3292 & po129 ;
  assign n4388 = ~n3289 & ~po129 ;
  assign n4389 = n3289 & ~po129 ;
  assign n4390 = n3292 & po129 ;
  assign n4391 = ~n4389 & ~n4390;
  assign n4392 = ~n4387 & ~n4388;
  assign n4393 = ~n3361 & po129 ;
  assign n4394 = ~n3364 & ~po129 ;
  assign n4395 = n3364 & ~po129 ;
  assign n4396 = n3361 & po129 ;
  assign n4397 = ~n4395 & ~n4396;
  assign n4398 = ~n4393 & ~n4394;
  assign n4399 = ~n3357 & po129 ;
  assign n4400 = ~n3354 & ~po129 ;
  assign n4401 = n3354 & ~po129 ;
  assign n4402 = n3357 & po129 ;
  assign n4403 = ~n4401 & ~n4402;
  assign n4404 = ~n4399 & ~n4400;
  assign n4405 = ~n3346 & po129 ;
  assign n4406 = ~n3349 & ~po129 ;
  assign n4407 = n3349 & ~po129 ;
  assign n4408 = n3346 & po129 ;
  assign n4409 = ~n4407 & ~n4408;
  assign n4410 = ~n4405 & ~n4406;
  assign n4411 = ~n3342 & po129 ;
  assign n4412 = ~n3339 & ~po129 ;
  assign n4413 = n3339 & ~po129 ;
  assign n4414 = n3342 & po129 ;
  assign n4415 = ~n4413 & ~n4414;
  assign n4416 = ~n4411 & ~n4412;
  assign n4417 = ~n3410 & po129 ;
  assign n4418 = ~n3413 & ~po129 ;
  assign n4419 = n3413 & ~po129 ;
  assign n4420 = n3410 & po129 ;
  assign n4421 = ~n4419 & ~n4420;
  assign n4422 = ~n4417 & ~n4418;
  assign n4423 = ~n3406 & po129 ;
  assign n4424 = ~n3403 & ~po129 ;
  assign n4425 = n3403 & ~po129 ;
  assign n4426 = n3406 & po129 ;
  assign n4427 = ~n4425 & ~n4426;
  assign n4428 = ~n4423 & ~n4424;
  assign n4429 = ~n3395 & po129 ;
  assign n4430 = ~n3398 & ~po129 ;
  assign n4431 = n3398 & ~po129 ;
  assign n4432 = n3395 & po129 ;
  assign n4433 = ~n4431 & ~n4432;
  assign n4434 = ~n4429 & ~n4430;
  assign n4435 = ~n3391 & po129 ;
  assign n4436 = ~n3388 & ~po129 ;
  assign n4437 = n3388 & ~po129 ;
  assign n4438 = n3391 & po129 ;
  assign n4439 = ~n4437 & ~n4438;
  assign n4440 = ~n4435 & ~n4436;
  assign n4441 = ~n3460 & po129 ;
  assign n4442 = ~n3463 & ~po129 ;
  assign n4443 = n3463 & ~po129 ;
  assign n4444 = n3460 & po129 ;
  assign n4445 = ~n4443 & ~n4444;
  assign n4446 = ~n4441 & ~n4442;
  assign n4447 = ~n3456 & po129 ;
  assign n4448 = ~n3453 & ~po129 ;
  assign n4449 = n3453 & ~po129 ;
  assign n4450 = n3456 & po129 ;
  assign n4451 = ~n4449 & ~n4450;
  assign n4452 = ~n4447 & ~n4448;
  assign n4453 = ~n3445 & po129 ;
  assign n4454 = ~n3448 & ~po129 ;
  assign n4455 = n3448 & ~po129 ;
  assign n4456 = n3445 & po129 ;
  assign n4457 = ~n4455 & ~n4456;
  assign n4458 = ~n4453 & ~n4454;
  assign n4459 = ~n3441 & po129 ;
  assign n4460 = ~n3438 & ~po129 ;
  assign n4461 = n3438 & ~po129 ;
  assign n4462 = n3441 & po129 ;
  assign n4463 = ~n4461 & ~n4462;
  assign n4464 = ~n4459 & ~n4460;
  assign n4465 = ~n3504 & po129 ;
  assign n4466 = ~n3507 & ~po129 ;
  assign n4467 = n3507 & ~po129 ;
  assign n4468 = n3504 & po129 ;
  assign n4469 = ~n4467 & ~n4468;
  assign n4470 = ~n4465 & ~n4466;
  assign n4471 = ~n3500 & po129 ;
  assign n4472 = ~n3497 & ~po129 ;
  assign n4473 = n3497 & ~po129 ;
  assign n4474 = n3500 & po129 ;
  assign n4475 = ~n4473 & ~n4474;
  assign n4476 = ~n4471 & ~n4472;
  assign n4477 = ~n3489 & po129 ;
  assign n4478 = ~n3492 & ~po129 ;
  assign n4479 = n3492 & ~po129 ;
  assign n4480 = n3489 & po129 ;
  assign n4481 = ~n4479 & ~n4480;
  assign n4482 = ~n4477 & ~n4478;
  assign n4483 = ~n3485 & po129 ;
  assign n4484 = ~n3482 & ~po129 ;
  assign n4485 = n3482 & ~po129 ;
  assign n4486 = n3485 & po129 ;
  assign n4487 = ~n4485 & ~n4486;
  assign n4488 = ~n4483 & ~n4484;
  assign n4489 = ~n3554 & po129 ;
  assign n4490 = ~n3557 & ~po129 ;
  assign n4491 = n3557 & ~po129 ;
  assign n4492 = n3554 & po129 ;
  assign n4493 = ~n4491 & ~n4492;
  assign n4494 = ~n4489 & ~n4490;
  assign n4495 = ~n3550 & po129 ;
  assign n4496 = ~n3547 & ~po129 ;
  assign n4497 = n3547 & ~po129 ;
  assign n4498 = n3550 & po129 ;
  assign n4499 = ~n4497 & ~n4498;
  assign n4500 = ~n4495 & ~n4496;
  assign n4501 = ~n3539 & po129 ;
  assign n4502 = ~n3542 & ~po129 ;
  assign n4503 = n3542 & ~po129 ;
  assign n4504 = n3539 & po129 ;
  assign n4505 = ~n4503 & ~n4504;
  assign n4506 = ~n4501 & ~n4502;
  assign n4507 = ~n3535 & po129 ;
  assign n4508 = ~n3532 & ~po129 ;
  assign n4509 = n3532 & ~po129 ;
  assign n4510 = n3535 & po129 ;
  assign n4511 = ~n4509 & ~n4510;
  assign n4512 = ~n4507 & ~n4508;
  assign n4513 = ~n3603 & po129 ;
  assign n4514 = ~n3606 & ~po129 ;
  assign n4515 = n3606 & ~po129 ;
  assign n4516 = n3603 & po129 ;
  assign n4517 = ~n4515 & ~n4516;
  assign n4518 = ~n4513 & ~n4514;
  assign n4519 = ~n3599 & po129 ;
  assign n4520 = ~n3596 & ~po129 ;
  assign n4521 = n3596 & ~po129 ;
  assign n4522 = n3599 & po129 ;
  assign n4523 = ~n4521 & ~n4522;
  assign n4524 = ~n4519 & ~n4520;
  assign n4525 = ~n3588 & po129 ;
  assign n4526 = ~n3591 & ~po129 ;
  assign n4527 = n3591 & ~po129 ;
  assign n4528 = n3588 & po129 ;
  assign n4529 = ~n4527 & ~n4528;
  assign n4530 = ~n4525 & ~n4526;
  assign n4531 = ~n3584 & po129 ;
  assign n4532 = ~n3581 & ~po129 ;
  assign n4533 = n3581 & ~po129 ;
  assign n4534 = n3584 & po129 ;
  assign n4535 = ~n4533 & ~n4534;
  assign n4536 = ~n4531 & ~n4532;
  assign n4537 = ~n3653 & po129 ;
  assign n4538 = ~n3656 & ~po129 ;
  assign n4539 = n3656 & ~po129 ;
  assign n4540 = n3653 & po129 ;
  assign n4541 = ~n4539 & ~n4540;
  assign n4542 = ~n4537 & ~n4538;
  assign n4543 = ~n3649 & po129 ;
  assign n4544 = ~n3646 & ~po129 ;
  assign n4545 = n3646 & ~po129 ;
  assign n4546 = n3649 & po129 ;
  assign n4547 = ~n4545 & ~n4546;
  assign n4548 = ~n4543 & ~n4544;
  assign n4549 = ~n3638 & po129 ;
  assign n4550 = ~n3641 & ~po129 ;
  assign n4551 = n3641 & ~po129 ;
  assign n4552 = n3638 & po129 ;
  assign n4553 = ~n4551 & ~n4552;
  assign n4554 = ~n4549 & ~n4550;
  assign n4555 = ~n3634 & po129 ;
  assign n4556 = ~n3631 & ~po129 ;
  assign n4557 = n3631 & ~po129 ;
  assign n4558 = n3634 & po129 ;
  assign n4559 = ~n4557 & ~n4558;
  assign n4560 = ~n4555 & ~n4556;
  assign n4561 = ~n3697 & po129 ;
  assign n4562 = ~n3700 & ~po129 ;
  assign n4563 = n3700 & ~po129 ;
  assign n4564 = n3697 & po129 ;
  assign n4565 = ~n4563 & ~n4564;
  assign n4566 = ~n4561 & ~n4562;
  assign n4567 = ~n3693 & po129 ;
  assign n4568 = ~n3690 & ~po129 ;
  assign n4569 = n3690 & ~po129 ;
  assign n4570 = n3693 & po129 ;
  assign n4571 = ~n4569 & ~n4570;
  assign n4572 = ~n4567 & ~n4568;
  assign n4573 = ~n3682 & po129 ;
  assign n4574 = ~n3685 & ~po129 ;
  assign n4575 = n3685 & ~po129 ;
  assign n4576 = n3682 & po129 ;
  assign n4577 = ~n4575 & ~n4576;
  assign n4578 = ~n4573 & ~n4574;
  assign n4579 = ~n3678 & po129 ;
  assign n4580 = ~n3675 & ~po129 ;
  assign n4581 = n3675 & ~po129 ;
  assign n4582 = n3678 & po129 ;
  assign n4583 = ~n4581 & ~n4582;
  assign n4584 = ~n4579 & ~n4580;
  assign n4585 = ~n3747 & po129 ;
  assign n4586 = ~n3750 & ~po129 ;
  assign n4587 = n3750 & ~po129 ;
  assign n4588 = n3747 & po129 ;
  assign n4589 = ~n4587 & ~n4588;
  assign n4590 = ~n4585 & ~n4586;
  assign n4591 = ~n3743 & po129 ;
  assign n4592 = ~n3740 & ~po129 ;
  assign n4593 = n3740 & ~po129 ;
  assign n4594 = n3743 & po129 ;
  assign n4595 = ~n4593 & ~n4594;
  assign n4596 = ~n4591 & ~n4592;
  assign n4597 = ~n3732 & po129 ;
  assign n4598 = ~n3735 & ~po129 ;
  assign n4599 = n3735 & ~po129 ;
  assign n4600 = n3732 & po129 ;
  assign n4601 = ~n4599 & ~n4600;
  assign n4602 = ~n4597 & ~n4598;
  assign n4603 = ~n3728 & po129 ;
  assign n4604 = ~n3725 & ~po129 ;
  assign n4605 = n3725 & ~po129 ;
  assign n4606 = n3728 & po129 ;
  assign n4607 = ~n4605 & ~n4606;
  assign n4608 = ~n4603 & ~n4604;
  assign n4609 = ~n3796 & po129 ;
  assign n4610 = ~n3799 & ~po129 ;
  assign n4611 = n3799 & ~po129 ;
  assign n4612 = n3796 & po129 ;
  assign n4613 = ~n4611 & ~n4612;
  assign n4614 = ~n4609 & ~n4610;
  assign n4615 = ~n3792 & po129 ;
  assign n4616 = ~n3789 & ~po129 ;
  assign n4617 = n3789 & ~po129 ;
  assign n4618 = n3792 & po129 ;
  assign n4619 = ~n4617 & ~n4618;
  assign n4620 = ~n4615 & ~n4616;
  assign n4621 = ~n3781 & po129 ;
  assign n4622 = ~n3784 & ~po129 ;
  assign n4623 = n3784 & ~po129 ;
  assign n4624 = n3781 & po129 ;
  assign n4625 = ~n4623 & ~n4624;
  assign n4626 = ~n4621 & ~n4622;
  assign n4627 = ~n3777 & po129 ;
  assign n4628 = ~n3774 & ~po129 ;
  assign n4629 = n3774 & ~po129 ;
  assign n4630 = n3777 & po129 ;
  assign n4631 = ~n4629 & ~n4630;
  assign n4632 = ~n4627 & ~n4628;
  assign n4633 = ~n3848 & po129 ;
  assign n4634 = ~n3851 & ~po129 ;
  assign n4635 = n3851 & ~po129 ;
  assign n4636 = n3848 & po129 ;
  assign n4637 = ~n4635 & ~n4636;
  assign n4638 = ~n4633 & ~n4634;
  assign n4639 = ~n3844 & po129 ;
  assign n4640 = ~n3841 & ~po129 ;
  assign n4641 = n3841 & ~po129 ;
  assign n4642 = n3844 & po129 ;
  assign n4643 = ~n4641 & ~n4642;
  assign n4644 = ~n4639 & ~n4640;
  assign n4645 = ~n3833 & po129 ;
  assign n4646 = ~n3836 & ~po129 ;
  assign n4647 = n3836 & ~po129 ;
  assign n4648 = n3833 & po129 ;
  assign n4649 = ~n4647 & ~n4648;
  assign n4650 = ~n4645 & ~n4646;
  assign n4651 = ~n3829 & po129 ;
  assign n4652 = ~n3826 & ~po129 ;
  assign n4653 = n3826 & ~po129 ;
  assign n4654 = n3829 & po129 ;
  assign n4655 = ~n4653 & ~n4654;
  assign n4656 = ~n4651 & ~n4652;
  assign n4657 = ~n3901 & po129 ;
  assign n4658 = ~n3898 & ~po129 ;
  assign n4659 = n3898 & ~po129 ;
  assign n4660 = n3901 & po129 ;
  assign n4661 = ~n4659 & ~n4660;
  assign n4662 = ~n4657 & ~n4658;
  assign n4663 = ~n3882 & po129 ;
  assign n4664 = ~n3879 & ~po129 ;
  assign n4665 = n3879 & ~po129 ;
  assign n4666 = n3882 & po129 ;
  assign n4667 = ~n4665 & ~n4666;
  assign n4668 = ~n4663 & ~n4664;
  assign n4669 = ~n3875 & po129 ;
  assign n4670 = ~n3872 & ~po129 ;
  assign n4671 = n3872 & ~po129 ;
  assign n4672 = n3875 & po129 ;
  assign n4673 = ~n4671 & ~n4672;
  assign n4674 = ~n4669 & ~n4670;
  assign n4675 = n4767 & ~po129 ;
  assign n4676 = n4851 & po129 ;
  assign n4677 = ~n4851 & po129 ;
  assign n4678 = ~n4767 & ~po129 ;
  assign n4679 = ~n4677 & ~n4678;
  assign n4680 = ~n4675 & ~n4676;
  assign n4681 = ~n4936 & n3919;
  assign n4682 = n4937 & ~n4681;
  assign n4683 = n4936 & n4937;
  assign n4684 = n699 | n700;
  assign n4685 = n708 | n709;
  assign n4686 = n714 | n715;
  assign n4687 = n724 | n725;
  assign n4688 = n730 | n731;
  assign n4689 = n748 | n749;
  assign n4690 = n754 | n755;
  assign n4691 = n772 | n773;
  assign n4692 = n778 | n779;
  assign n4693 = n791 | n792;
  assign n4694 = n803 | n804;
  assign n4695 = n813 | ~n814;
  assign n4696 = n820 | n821;
  assign n4697 = n832 | n833;
  assign n4698 = n845 | n840 | n844;
  assign n4699 = n849 | n850;
  assign n4700 = n855 | n856;
  assign n4701 = n861 | n862;
  assign n4702 = n869 | n870;
  assign n4703 = n875 | n876;
  assign n4704 = n880 | ~n881;
  assign n4705 = n882 | n883;
  assign n4706 = n889 | ~n890;
  assign n4707 = n904 | n905;
  assign n4708 = n914 | n915;
  assign n4709 = n920 | n921;
  assign n4710 = n928 | n929;
  assign n4711 = n934 | n935;
  assign n4712 = n939 | n940;
  assign n4713 = n944 | n945;
  assign n4714 = n950 | ~n951;
  assign n4715 = n969 | n965 | n968;
  assign n4716 = n974 | n975;
  assign n4717 = n980 | n981;
  assign n4718 = n987 | n988;
  assign n4719 = n993 | n994;
  assign n4720 = n999 | ~n1000;
  assign n4721 = n1001 | n1002;
  assign n4722 = n1008 | ~n1009;
  assign n4723 = n1026 | n1023 | n1025;
  assign n4724 = n1035 | n1036;
  assign n4725 = n1041 | n1042;
  assign n4726 = n1049 | n1050;
  assign n4727 = n1055 | n1056;
  assign n4728 = n1060 | n1061;
  assign n4729 = n1065 | n1066;
  assign n4730 = n1076 | n1077;
  assign n4731 = n1085 | n1086;
  assign n4732 = n1109 | n1110;
  assign n4733 = n1112 | n1113;
  assign n4734 = n1116 | n1117;
  assign n4735 = n1133 | n1134;
  assign n4736 = n1157 | n1158;
  assign n4737 = n1160 | n1161;
  assign n4738 = n1164 | n1165;
  assign n4739 = n1175 | n1176;
  assign n4740 = n1180 | n1181;
  assign n4741 = n1186 | n1187;
  assign n4742 = n1210 | n1211;
  assign n4743 = n1213 | n1214;
  assign n4744 = n1217 | n1218;
  assign n4745 = n1234 | n1235;
  assign n4746 = n1258 | n1259;
  assign n4747 = n1261 | n1262;
  assign n4748 = n1265 | n1266;
  assign n4749 = n1276 | n1277;
  assign n4750 = n1281 | n1282;
  assign n4751 = n1287 | n1288;
  assign n4752 = n1311 | n1312;
  assign n4753 = n1314 | n1315;
  assign n4754 = n1318 | n1319;
  assign n4755 = n1335 | n1336;
  assign n4756 = n1359 | n1360;
  assign n4757 = n1362 | n1363;
  assign n4758 = n1366 | n1367;
  assign n4759 = n1377 | n1378;
  assign n4760 = n1382 | n1383;
  assign n4761 = n1388 | n1389;
  assign n4762 = n1412 | n1413;
  assign n4763 = n1415 | n1416;
  assign n4764 = n1419 | n1420;
  assign n4765 = n1436 | n1437;
  assign n4766 = n1448 | n1449;
  assign n4767 = n1461 | n1462;
  assign n4768 = n1524 | n1525;
  assign n4769 = n1533 | n1534;
  assign n4770 = n1539 | n1540;
  assign n4771 = n1549 | n1550;
  assign n4772 = n1555 | n1556;
  assign n4773 = n1573 | n1574;
  assign n4774 = n1579 | n1580;
  assign n4775 = n1597 | n1598;
  assign n4776 = n1603 | n1604;
  assign n4777 = n1616 | n1617;
  assign n4778 = n1628 | n1629;
  assign n4779 = n1638 | ~n1639;
  assign n4780 = n1645 | n1646;
  assign n4781 = n1657 | n1658;
  assign n4782 = n1670 | n1665 | n1669;
  assign n4783 = n1674 | n1675;
  assign n4784 = n1680 | n1681;
  assign n4785 = n1686 | n1687;
  assign n4786 = n1694 | n1695;
  assign n4787 = n1700 | n1701;
  assign n4788 = n1705 | ~n1706;
  assign n4789 = n1707 | n1708;
  assign n4790 = n1714 | ~n1715;
  assign n4791 = n1729 | n1730;
  assign n4792 = n1739 | n1740;
  assign n4793 = n1745 | n1746;
  assign n4794 = n1753 | n1754;
  assign n4795 = n1759 | n1760;
  assign n4796 = n1764 | n1765;
  assign n4797 = n1769 | n1770;
  assign n4798 = n1775 | ~n1776;
  assign n4799 = n1794 | n1790 | n1793;
  assign n4800 = n1799 | n1800;
  assign n4801 = n1805 | n1806;
  assign n4802 = n1812 | n1813;
  assign n4803 = n1818 | n1819;
  assign n4804 = n1824 | ~n1825;
  assign n4805 = n1826 | n1827;
  assign n4806 = n1833 | ~n1834;
  assign n4807 = n1851 | n1848 | n1850;
  assign n4808 = n1860 | n1861;
  assign n4809 = n1866 | n1867;
  assign n4810 = n1874 | n1875;
  assign n4811 = n1880 | n1881;
  assign n4812 = n1885 | n1886;
  assign n4813 = n1890 | n1891;
  assign n4814 = n1901 | n1902;
  assign n4815 = n1910 | n1911;
  assign n4816 = n1934 | n1935;
  assign n4817 = n1937 | n1938;
  assign n4818 = n1941 | n1942;
  assign n4819 = n1958 | n1959;
  assign n4820 = n1982 | n1983;
  assign n4821 = n1985 | n1986;
  assign n4822 = n1989 | n1990;
  assign n4823 = n2000 | n2001;
  assign n4824 = n2005 | n2006;
  assign n4825 = n2011 | n2012;
  assign n4826 = n2035 | n2036;
  assign n4827 = n2038 | n2039;
  assign n4828 = n2042 | n2043;
  assign n4829 = n2059 | n2060;
  assign n4830 = n2083 | n2084;
  assign n4831 = n2086 | n2087;
  assign n4832 = n2090 | n2091;
  assign n4833 = n2101 | n2102;
  assign n4834 = n2106 | n2107;
  assign n4835 = n2112 | n2113;
  assign n4836 = n2136 | n2137;
  assign n4837 = n2139 | n2140;
  assign n4838 = n2143 | n2144;
  assign n4839 = n2160 | n2161;
  assign n4840 = n2184 | n2185;
  assign n4841 = n2187 | n2188;
  assign n4842 = n2191 | n2192;
  assign n4843 = n2202 | n2203;
  assign n4844 = n2207 | n2208;
  assign n4845 = n2213 | n2214;
  assign n4846 = n2237 | n2238;
  assign n4847 = n2240 | n2241;
  assign n4848 = n2244 | n2245;
  assign n4849 = n2261 | n2262;
  assign n4850 = n2273 | n2274;
  assign n4851 = n2286 | n2287;
  assign n4852 = n2396 | ~n2397;
  assign n4853 = n2402 | n2403;
  assign n4854 = n2408 | n2409;
  assign n4855 = n2410 | ~n2411;
  assign n4856 = n2414 | ~n2415;
  assign n4857 = n2435 | ~n2436;
  assign n4858 = ~n2445 | n2440 | ~n2444;
  assign n4859 = n2462 | ~n2463;
  assign n4860 = n2464 | n2465;
  assign n4861 = n2496 | ~n2497;
  assign n4862 = n2502 | n2503;
  assign n4863 = n2517 | n2518;
  assign n4864 = n2543 | n2544;
  assign n4865 = n2563 | ~n2564;
  assign n4866 = n2568 | n2569;
  assign n4867 = n2582 | n2583;
  assign n4868 = n2603 | n2604;
  assign n4869 = n2627 | n2628;
  assign n4870 = n2647 | ~n2648;
  assign n4871 = n2652 | n2653;
  assign n4872 = n2666 | n2667;
  assign n4873 = n2692 | n2693;
  assign n4874 = n2727 | n2728;
  assign n4875 = n2752 | n2753;
  assign n4876 = n2781 | n2773 | n2780;
  assign n4877 = n2776 | n2777;
  assign n4878 = n2791 | n2787 | n2790;
  assign n4879 = n2798 | n2799;
  assign n4880 = n2803 | n2804;
  assign n4881 = n2808 | n2809;
  assign n4882 = n2817 | n2818;
  assign n4883 = n2827 | n2823 | n2826;
  assign n4884 = n2861 | n2862;
  assign n4885 = n2863 | n2864;
  assign n4886 = n2899 | n2900;
  assign n4887 = n2909 | n2910;
  assign n4888 = n2923 | n2924;
  assign n4889 = n2929 | n2930;
  assign n4890 = n2934 | n2935;
  assign n4891 = n2990 | n2991;
  assign n4892 = n3004 | n3001 | n3003;
  assign n4893 = n3013 | n3014;
  assign n4894 = n3017 | n3018;
  assign n4895 = n3027 | n3028;
  assign n4896 = n3032 | n3033;
  assign n4897 = n3067 | n3068;
  assign n4898 = n3069 | n3070;
  assign n4899 = n3108 | n3105 | n3107;
  assign n4900 = n3117 | n3118;
  assign n4901 = n3131 | n3132;
  assign n4902 = n3137 | n3138;
  assign n4903 = n3142 | n3143;
  assign n4904 = n3177 | n3178;
  assign n4905 = n3182 | n3183;
  assign n4906 = n3188 | n3189;
  assign n4907 = n3237 | n3238;
  assign n4908 = n3241 | n3242;
  assign n4909 = n3282 | n3283;
  assign n4910 = n3331 | n3332;
  assign n4911 = n3335 | n3336;
  assign n4912 = n3370 | n3371;
  assign n4913 = n3375 | n3376;
  assign n4914 = n3381 | n3382;
  assign n4915 = n3430 | n3431;
  assign n4916 = n3434 | n3435;
  assign n4917 = n3475 | n3476;
  assign n4918 = n3524 | n3525;
  assign n4919 = n3528 | n3529;
  assign n4920 = n3563 | n3564;
  assign n4921 = n3568 | n3569;
  assign n4922 = n3574 | n3575;
  assign n4923 = n3623 | n3624;
  assign n4924 = n3627 | n3628;
  assign n4925 = n3668 | n3669;
  assign n4926 = n3717 | n3718;
  assign n4927 = n3721 | n3722;
  assign n4928 = n3756 | n3757;
  assign n4929 = n3761 | n3762;
  assign n4930 = n3767 | n3768;
  assign n4931 = n3807 | n3808;
  assign n4932 = n3818 | n3819;
  assign n4933 = n3822 | n3823;
  assign n4934 = n3859 | n3860;
  assign n4935 = n3865 | n3866;
  assign n4936 = n3889 | n3886 | n3888;
  assign n4937 = n3894 | n3891 | n3893;
  assign n4938 = n3905 | n3906;
  assign po129  = n3920 | n3921;
  assign po1  = n3929 | ~n3930;
  assign po2  = n3935 | ~n3936;
  assign po3  = n3941 | ~n3942;
  assign n4943 = n3953 | ~n3954;
  assign po7  = n3959 | ~n3960;
  assign po8  = n3965 | ~n3966;
  assign po9  = n3971 | ~n3972;
  assign po10  = n3977 | ~n3978;
  assign po11  = n3983 | ~n3984;
  assign po12  = n3989 | ~n3990;
  assign po13  = n3995 | ~n3996;
  assign po14  = n4001 | ~n4002;
  assign po15  = n4007 | ~n4008;
  assign po16  = n4013 | ~n4014;
  assign po17  = n4019 | ~n4020;
  assign po18  = n4025 | ~n4026;
  assign po19  = n4031 | ~n4032;
  assign po20  = n4037 | ~n4038;
  assign po21  = n4043 | ~n4044;
  assign po22  = n4049 | ~n4050;
  assign po23  = n4055 | ~n4056;
  assign po24  = n4061 | ~n4062;
  assign po25  = n4067 | ~n4068;
  assign po26  = n4073 | ~n4074;
  assign po27  = n4079 | ~n4080;
  assign po28  = n4085 | ~n4086;
  assign po29  = n4091 | ~n4092;
  assign po30  = n4097 | ~n4098;
  assign po31  = n4103 | ~n4104;
  assign po32  = n4109 | ~n4110;
  assign po33  = n4115 | ~n4116;
  assign po34  = n4121 | ~n4122;
  assign po35  = n4127 | ~n4128;
  assign po36  = n4133 | ~n4134;
  assign po37  = n4139 | ~n4140;
  assign po38  = n4145 | ~n4146;
  assign po39  = n4151 | ~n4152;
  assign po40  = n4157 | ~n4158;
  assign po41  = n4163 | ~n4164;
  assign po42  = n4169 | ~n4170;
  assign po43  = n4175 | ~n4176;
  assign po44  = n4181 | ~n4182;
  assign po45  = n4187 | ~n4188;
  assign po46  = n4193 | ~n4194;
  assign po47  = n4199 | ~n4200;
  assign po48  = n4205 | ~n4206;
  assign po49  = n4211 | ~n4212;
  assign po50  = n4217 | ~n4218;
  assign po51  = n4223 | ~n4224;
  assign po52  = n4229 | ~n4230;
  assign po53  = n4235 | ~n4236;
  assign po54  = n4241 | ~n4242;
  assign po55  = n4247 | ~n4248;
  assign po56  = n4253 | ~n4254;
  assign po57  = n4259 | ~n4260;
  assign po58  = n4265 | ~n4266;
  assign po59  = n4271 | ~n4272;
  assign po60  = n4277 | ~n4278;
  assign po61  = n4283 | ~n4284;
  assign po62  = n4289 | ~n4290;
  assign po63  = n4295 | ~n4296;
  assign po64  = n4301 | ~n4302;
  assign po65  = n4307 | ~n4308;
  assign po66  = n4313 | ~n4314;
  assign po67  = n4319 | ~n4320;
  assign po68  = n4325 | ~n4326;
  assign po69  = n4331 | ~n4332;
  assign po70  = n4337 | ~n4338;
  assign po71  = n4343 | ~n4344;
  assign po72  = n4349 | ~n4350;
  assign po73  = n4355 | ~n4356;
  assign po74  = n4361 | ~n4362;
  assign po75  = n4367 | ~n4368;
  assign po76  = n4373 | ~n4374;
  assign po77  = n4379 | ~n4380;
  assign po78  = n4385 | ~n4386;
  assign po79  = n4391 | ~n4392;
  assign po80  = n4397 | ~n4398;
  assign po81  = n4403 | ~n4404;
  assign po82  = n4409 | ~n4410;
  assign po83  = n4415 | ~n4416;
  assign po84  = n4421 | ~n4422;
  assign po85  = n4427 | ~n4428;
  assign po86  = n4433 | ~n4434;
  assign po87  = n4439 | ~n4440;
  assign po88  = n4445 | ~n4446;
  assign po89  = n4451 | ~n4452;
  assign po90  = n4457 | ~n4458;
  assign po91  = n4463 | ~n4464;
  assign po92  = n4469 | ~n4470;
  assign po93  = n4475 | ~n4476;
  assign po94  = n4481 | ~n4482;
  assign po95  = n4487 | ~n4488;
  assign po96  = n4493 | ~n4494;
  assign po97  = n4499 | ~n4500;
  assign po98  = n4505 | ~n4506;
  assign po99  = n4511 | ~n4512;
  assign po100  = n4517 | ~n4518;
  assign po101  = n4523 | ~n4524;
  assign po102  = n4529 | ~n4530;
  assign po103  = n4535 | ~n4536;
  assign po104  = n4541 | ~n4542;
  assign po105  = n4547 | ~n4548;
  assign po106  = n4553 | ~n4554;
  assign po107  = n4559 | ~n4560;
  assign po108  = n4565 | ~n4566;
  assign po109  = n4571 | ~n4572;
  assign po110  = n4577 | ~n4578;
  assign po111  = n4583 | ~n4584;
  assign po112  = n4589 | ~n4590;
  assign po113  = n4595 | ~n4596;
  assign po114  = n4601 | ~n4602;
  assign po115  = n4607 | ~n4608;
  assign po116  = n4613 | ~n4614;
  assign po117  = n4619 | ~n4620;
  assign po118  = n4625 | ~n4626;
  assign po119  = n4631 | ~n4632;
  assign po120  = n4637 | ~n4638;
  assign po121  = n4643 | ~n4644;
  assign po122  = n4649 | ~n4650;
  assign po123  = n4655 | ~n4656;
  assign po124  = n4661 | ~n4662;
  assign po125  = n4667 | ~n4668;
  assign po126  = n4673 | ~n4674;
  assign po128  = n4679 | ~n4680;
  assign po127  = n4682 | n4683;
  assign po0  = ~n3924;
  assign po4  = ~n3945;
  assign po5  = ~n3948;
  assign po6  = ~n4943;
endmodule
