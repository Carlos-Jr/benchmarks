module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n367, n368,
    n369, n370, n371, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404,
    n406, n407, n408, n409, n410, n411, n412,
    n413, n414, n415, n416, n418, n419, n420,
    n421, n422, n423, n424, n425, n426, n427,
    n429, n430, n431, n432, n433, n434, n435,
    n436, n437, n438, n439, n441, n442, n443,
    n444, n445, n446, n447, n448, n450, n451,
    n452, n453, n454, n455, n457, n458, n459,
    n460, n461, n462, n463, n465, n466, n467,
    n468, n469, n470, n471, n472, n473, n474,
    n476, n477, n478, n479, n480, n481, n482,
    n484, n485, n486, n487, n488, n489, n490,
    n491, n493, n494, n495, n496, n497, n499,
    n500, n501, n502, n503, n504, n505, n507,
    n508, n509, n510, n511, n512, n513, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529,
    n530, n531, n532, n533, n534, n535, n536,
    n537, n538, n539, n541, n542, n543, n544,
    n545, n546, n548, n549, n550, n551, n552,
    n553, n554, n555, n556, n557, n559, n560,
    n561, n562, n563, n564, n566, n567, n568,
    n569, n570, n572, n573, n574, n575, n576,
    n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n591,
    n592, n593, n594, n595, n596, n597, n599,
    n600, n601, n602, n603, n604, n605, n606,
    n608, n609, n611, n612, n613, n614, n615,
    n616, n617, n618, n619, n620, n621, n622,
    n623, n624, n625, n626, n627, n628, n630,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651,
    n652, n653, n654, n655, n656, n657, n658,
    n659, n660, n661, n662, n663, n664, n665,
    n666, n667, n668, n669, n670, n671, n672,
    n673, n675, n676, n677, n678, n679, n680,
    n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n692, n693, n694, n695, n696,
    n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n710,
    n711, n712, n713, n714, n715, n716, n717,
    n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n732,
    n733, n734, n735, n736, n737, n738, n739,
    n740, n741, n742, n743, n744, n745, n746,
    n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n761,
    n762, n763, n764, n765, n766, n768, n769,
    n770, n771, n772, n773, n775, n776, n777,
    n778, n779, n780, n782, n783, n784, n785,
    n786, n787, n789, n790, n791, n792, n793,
    n794, n796, n797, n798, n799, n800, n801,
    n803, n804, n805, n806, n807, n808, n810,
    n811, n812, n813, n814, n815, n817, n818,
    n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839,
    n841, n842, n843, n844, n845, n846, n848,
    n849, n850, n851, n852, n853, n854, n855,
    n856, n857, n858, n859, n860, n861, n862,
    n863, n865, n866, n867, n868, n869, n870,
    n871, n872, n873, n874, n875, n876, n877,
    n879, n880, n881, n882, n883, n884, n885,
    n886, n887, n888, n889, n890, n892, n893,
    n894, n895, n896, n897, n898, n899, n900,
    n901, n902, n903, n904, n905, n906, n907,
    n909, n910, n911, n912, n913, n914, n916,
    n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n927, n928, n929, n931,
    n932, n933, n934, n935, n936, n937, n938,
    n939, n940, n942, n943, n944, n945, n946,
    n947, n948, n949, n950, n951, n952, n953,
    n954, n956, n957, n958, n959, n960, n961,
    n962, n963, n964, n965, n966, n967, n968,
    n969, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983,
    n984, n986, n987, n988, n989, n990, n991,
    n992, n993, n994, n995, n996, n997, n998,
    n1000, n1001, n1002, n1004, n1005, n1006,
    n1008, n1009, n1010, n1011, n1012, n1013,
    n1014, n1015, n1016, n1018, n1019, n1020,
    n1023, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1038, n1039, n1040, n1041,
    n1042, n1043, n1045, n1046, n1047, n1048,
    n1049, n1050, n1051, n1052, n1053, n1054,
    n1055, n1056, n1057, n1058, n1060, n1061,
    n1062, n1063, n1064, n1065, n1067, n1068,
    n1069, n1070, n1071, n1072, n1073, n1074,
    n1075, n1076, n1077, n1078, n1079, n1080,
    n1081, n1082, n1083, n1084, n1086, n1087,
    n1088, n1090, n1091, n1093, n1094, n1095,
    n1096, n1097, n1098, n1099, n1100, n1102,
    n1103, n1104, n1106, n1107, n1108, n1110,
    n1111, n1112, n1114, n1115, n1116, n1117,
    n1118, n1120, n1121, n1122, n1124, n1125,
    n1126, n1128, n1129, n1130, n1132, n1133,
    n1134, n1136, n1137, n1138, n1140, n1141,
    n1142, n1144, n1145, n1146, n1148, n1149,
    n1150, n1152, n1153, n1154, n1156, n1157,
    n1158, n1160, n1161, n1162, n1164, n1165,
    n1166, n1167, n1168, n1170, n1171, n1172,
    n1174, n1175, n1176, n1178, n1179, n1180,
    n1182, n1183, n1184, n1186, n1187, n1188,
    n1189, n1190, n1191, n1192, n1193, n1194,
    n1195, n1196, n1197, n1198, n1199, n1200,
    n1201, n1202, n1203, n1205, n1206, n1207,
    n1209, n1210, n1211, n1212, n1214, n1215,
    n1216, n1218, n1219, n1220, n1222, n1223,
    n1224, n1225, n1226, n1228, n1229, n1230,
    n1232, n1233, n1234, n1236, n1237, n1238,
    n1240, n1241, n1242, n1244, n1245, n1246,
    n1248, n1249, n1250, n1251, n1252, n1253,
    n1255, n1256, n1257, n1258, n1259, n1260,
    n1262, n1263, n1264, n1266, n1267, n1268,
    n1270, n1271, n1272, n1274, n1275, n1276,
    n1278, n1279, n1280, n1282, n1283, n1284,
    n1285, n1286, n1287, n1288, n1289, n1290,
    n1291, n1292, n1293, n1294, n1295, n1296,
    n1297, n1298, n1300, n1301, n1302, n1303,
    n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1315, n1316,
    n1317, n1318, n1319, n1320, n1321, n1322,
    n1323, n1324, n1325, n1326, n1327, n1328,
    n1330, n1331, n1332, n1333, n1334, n1335,
    n1336, n1337, n1338, n1339, n1340, n1341,
    n1342, n1343, n1345, n1346, n1347, n1348,
    n1349, n1350, n1351, n1352, n1353, n1354,
    n1355, n1356, n1357, n1358, n1359, n1360,
    n1361, n1363, n1364, n1365, n1367, n1368,
    n1369, n1370, n1371, n1372, n1373, n1374,
    n1375, n1376, n1377, n1378, n1379, n1380,
    n1381, n1382, n1383, n1385, n1386, n1387,
    n1388, n1389, n1390, n1391, n1392, n1393,
    n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1403, n1404, n1406, n1407,
    n1409, n1410, n1411, n1412, n1414, n1415,
    n1416, n1418, n1419, n1420, n1421, n1423,
    n1424, n1425, n1427, n1428, n1429, n1430,
    n1433, n1434, n1435, n1436, n1439, n1440,
    n1442, n1447, n1448, n1450;
  assign n291 = ~pi7 & ~pi13;
  assign n292 = ~pi9 & ~pi11;
  assign n293 = ~pi14 & ~pi22;
  assign n294 = ~pi17 & ~pi21;
  assign n295 = ~pi8 & n294;
  assign n296 = ~pi4 & ~pi19;
  assign n297 = ~pi18 & n296;
  assign n298 = ~pi16 & n297;
  assign n299 = ~pi6 & ~pi12;
  assign n300 = ~pi5 & n299;
  assign n301 = n291 & n292;
  assign n302 = n293 & n301;
  assign n303 = n295 & n300;
  assign n304 = n302 & n303;
  assign n305 = n298 & n304;
  assign n306 = pi54 & ~n305;
  assign n307 = ~pi0 & ~n306;
  assign n308 = ~pi5 & ~pi22;
  assign n309 = ~pi56 & ~n308;
  assign n310 = ~pi8 & ~pi21;
  assign n311 = n291 & n310;
  assign n312 = ~pi14 & n311;
  assign n313 = ~pi10 & n312;
  assign n314 = ~pi7 & n310;
  assign n315 = pi8 & pi21;
  assign n316 = pi7 & ~n310;
  assign n317 = ~pi13 & ~n315;
  assign n318 = ~n316 & n317;
  assign n319 = ~n314 & ~n318;
  assign n320 = ~pi14 & ~n319;
  assign n321 = ~n311 & ~n320;
  assign n322 = ~pi10 & ~n321;
  assign n323 = ~n312 & ~n322;
  assign n324 = ~pi17 & n299;
  assign n325 = n308 & n324;
  assign n326 = n298 & n325;
  assign n327 = ~n313 & n326;
  assign n328 = ~n323 & n327;
  assign n329 = ~n309 & ~n328;
  assign n330 = n292 & ~n329;
  assign n331 = ~pi56 & ~n292;
  assign n332 = n308 & n331;
  assign n333 = ~n330 & ~n332;
  assign n334 = pi54 & ~n333;
  assign n335 = ~n307 & ~n334;
  assign n336 = ~pi3 & ~pi129;
  assign po15 = n335 | ~n336;
  assign n338 = ~pi17 & pi54;
  assign n339 = ~pi5 & ~pi6;
  assign n340 = n291 & n339;
  assign n341 = ~pi11 & ~pi12;
  assign n342 = ~pi10 & ~pi22;
  assign n343 = ~pi14 & n310;
  assign n344 = n341 & n342;
  assign n345 = n343 & n344;
  assign n346 = n340 & n345;
  assign n347 = n298 & n346;
  assign n348 = n338 & ~n347;
  assign n349 = ~pi1 & ~n348;
  assign n350 = ~pi8 & ~pi11;
  assign n351 = n294 & n350;
  assign n352 = ~pi10 & pi54;
  assign n353 = n293 & n352;
  assign n354 = pi5 & pi6;
  assign n355 = pi12 & ~n339;
  assign n356 = ~pi7 & ~n354;
  assign n357 = ~n355 & n356;
  assign n358 = ~n300 & ~n357;
  assign n359 = ~pi13 & ~n358;
  assign n360 = ~pi5 & ~pi7;
  assign n361 = n299 & n360;
  assign n362 = ~n359 & ~n361;
  assign n363 = ~pi9 & ~n362;
  assign n364 = n291 & n300;
  assign n365 = ~n363 & ~n364;
  assign n366 = ~pi9 & n364;
  assign n367 = n351 & n353;
  assign n368 = n298 & n367;
  assign n369 = ~n366 & n368;
  assign n370 = ~n365 & n369;
  assign n371 = ~n349 & ~n370;
  assign po16 = ~n336 | n371;
  assign n373 = ~pi15 & ~pi20;
  assign n374 = ~pi24 & ~pi49;
  assign n375 = ~pi45 & n373;
  assign n376 = n374 & n375;
  assign n377 = ~pi41 & ~pi43;
  assign n378 = ~pi42 & ~pi44;
  assign n379 = ~pi38 & ~pi50;
  assign n380 = ~pi46 & n379;
  assign n381 = ~pi40 & n380;
  assign n382 = n378 & n381;
  assign n383 = n377 & n382;
  assign n384 = ~pi47 & n383;
  assign n385 = ~pi48 & n384;
  assign n386 = pi82 & n376;
  assign n387 = n385 & n386;
  assign n388 = pi122 & pi127;
  assign n389 = ~pi82 & ~n388;
  assign n390 = pi2 & ~n389;
  assign n391 = ~n387 & n390;
  assign n392 = ~pi40 & n378;
  assign n393 = ~pi41 & ~pi46;
  assign n394 = n379 & n393;
  assign n395 = ~pi43 & ~pi47;
  assign n396 = ~pi48 & n395;
  assign n397 = ~pi2 & n396;
  assign n398 = n376 & n397;
  assign n399 = n394 & n398;
  assign n400 = n392 & n399;
  assign n401 = pi82 & ~n400;
  assign n402 = ~pi65 & ~n388;
  assign n403 = ~n401 & n402;
  assign n404 = ~n391 & ~n403;
  assign po17 = ~pi129 & ~n404;
  assign n406 = pi0 & ~pi113;
  assign n407 = ~pi123 & n406;
  assign n408 = ~pi9 & ~pi14;
  assign n409 = n342 & n408;
  assign n410 = n340 & n409;
  assign n411 = ~pi12 & n351;
  assign n412 = n298 & n410;
  assign n413 = n411 & n412;
  assign n414 = ~pi61 & ~pi118;
  assign n415 = ~n413 & n414;
  assign n416 = ~n407 & ~n415;
  assign po18 = ~pi129 & ~n416;
  assign n418 = pi4 & ~pi54;
  assign n419 = ~pi16 & pi54;
  assign n420 = n296 & n419;
  assign n421 = ~pi18 & n420;
  assign n422 = n294 & n421;
  assign n423 = n350 & n422;
  assign n424 = pi10 & n293;
  assign n425 = n366 & n424;
  assign n426 = n423 & n425;
  assign n427 = ~n418 & ~n426;
  assign po19 = n336 & ~n427;
  assign n429 = pi5 & ~pi54;
  assign n430 = ~pi7 & ~pi29;
  assign n431 = ~pi13 & n409;
  assign n432 = ~pi59 & n351;
  assign n433 = n431 & n432;
  assign n434 = ~pi25 & pi28;
  assign n435 = n430 & n434;
  assign n436 = n300 & n435;
  assign n437 = n421 & n436;
  assign n438 = n433 & n437;
  assign n439 = ~n429 & ~n438;
  assign po20 = n336 & ~n439;
  assign n441 = pi6 & ~pi54;
  assign n442 = pi25 & ~pi28;
  assign n443 = ~pi29 & n442;
  assign n444 = n419 & n443;
  assign n445 = n297 & n361;
  assign n446 = n444 & n445;
  assign n447 = n433 & n446;
  assign n448 = ~n441 & ~n447;
  assign po21 = n336 & ~n448;
  assign n450 = pi7 & ~pi54;
  assign n451 = n361 & n431;
  assign n452 = pi8 & ~pi11;
  assign n453 = n422 & n452;
  assign n454 = n451 & n453;
  assign n455 = ~n450 & ~n454;
  assign po22 = n336 & ~n455;
  assign n457 = pi8 & ~pi54;
  assign n458 = ~pi17 & ~pi18;
  assign n459 = n350 & n458;
  assign n460 = pi21 & n420;
  assign n461 = n459 & n460;
  assign n462 = n451 & n461;
  assign n463 = ~n457 & ~n462;
  assign po23 = n336 & ~n463;
  assign n465 = pi9 & ~pi54;
  assign n466 = ~pi18 & n295;
  assign n467 = ~pi9 & n466;
  assign n468 = n342 & n467;
  assign n469 = pi11 & ~pi13;
  assign n470 = ~pi14 & n469;
  assign n471 = n361 & n470;
  assign n472 = n420 & n471;
  assign n473 = n468 & n472;
  assign n474 = ~n465 & ~n473;
  assign po24 = n336 & ~n474;
  assign n476 = pi10 & ~pi54;
  assign n477 = ~pi11 & n361;
  assign n478 = ~pi13 & pi14;
  assign n479 = n420 & n478;
  assign n480 = n477 & n479;
  assign n481 = n468 & n480;
  assign n482 = ~n476 & ~n481;
  assign po25 = n336 & ~n482;
  assign n484 = pi11 & ~pi54;
  assign n485 = ~pi10 & ~pi11;
  assign n486 = pi22 & n485;
  assign n487 = n408 & n486;
  assign n488 = n420 & n487;
  assign n489 = n364 & n466;
  assign n490 = n488 & n489;
  assign n491 = ~n484 & ~n490;
  assign po26 = n336 & ~n491;
  assign n493 = pi12 & ~pi54;
  assign n494 = pi18 & n420;
  assign n495 = n410 & n494;
  assign n496 = n411 & n495;
  assign n497 = ~n493 & ~n496;
  assign po27 = n336 & ~n497;
  assign n499 = pi13 & ~pi54;
  assign n500 = ~pi25 & ~pi28;
  assign n501 = pi29 & n500;
  assign n502 = ~pi59 & n501;
  assign n503 = n451 & n502;
  assign n504 = n423 & n503;
  assign n505 = ~n499 & ~n504;
  assign po28 = n336 & ~n505;
  assign n507 = pi14 & ~pi54;
  assign n508 = pi13 & ~pi16;
  assign n509 = n296 & n508;
  assign n510 = n353 & n509;
  assign n511 = n477 & n510;
  assign n512 = n467 & n511;
  assign n513 = ~n507 & ~n512;
  assign po29 = n336 & ~n513;
  assign n515 = ~pi82 & n388;
  assign n516 = pi15 & n515;
  assign n517 = ~pi45 & n374;
  assign n518 = n392 & n394;
  assign n519 = n396 & n517;
  assign n520 = n518 & n519;
  assign n521 = pi15 & ~n520;
  assign n522 = ~pi47 & ~pi48;
  assign n523 = ~pi45 & n522;
  assign n524 = ~pi2 & ~pi20;
  assign n525 = ~pi15 & n374;
  assign n526 = n523 & ~n524;
  assign n527 = n525 & n526;
  assign n528 = n383 & n527;
  assign n529 = ~n521 & ~n528;
  assign n530 = pi82 & ~n529;
  assign n531 = ~pi15 & n377;
  assign n532 = n522 & n531;
  assign n533 = n517 & n532;
  assign n534 = n382 & n533;
  assign n535 = pi82 & ~n534;
  assign n536 = ~pi70 & ~n388;
  assign n537 = ~n535 & n536;
  assign n538 = ~n516 & ~n537;
  assign n539 = ~n530 & n538;
  assign po30 = ~pi129 & ~n539;
  assign n541 = pi16 & ~pi54;
  assign n542 = pi6 & ~pi12;
  assign n543 = n360 & n542;
  assign n544 = n431 & n543;
  assign n545 = n423 & n544;
  assign n546 = ~n541 & ~n545;
  assign po31 = n336 & ~n546;
  assign n548 = pi17 & ~pi54;
  assign n549 = ~pi11 & n310;
  assign n550 = pi59 & n338;
  assign n551 = n430 & n500;
  assign n552 = n550 & n551;
  assign n553 = n300 & n549;
  assign n554 = n552 & n553;
  assign n555 = n298 & n431;
  assign n556 = n554 & n555;
  assign n557 = ~n548 & ~n556;
  assign po32 = n336 & ~n557;
  assign n559 = pi18 & ~pi54;
  assign n560 = n297 & n451;
  assign n561 = pi16 & pi54;
  assign n562 = n351 & n561;
  assign n563 = n560 & n562;
  assign n564 = ~n559 & ~n563;
  assign po33 = n336 & ~n564;
  assign n566 = pi19 & ~pi54;
  assign n567 = pi17 & n419;
  assign n568 = n549 & n567;
  assign n569 = n560 & n568;
  assign n570 = ~n566 & ~n569;
  assign po34 = n336 & ~n570;
  assign n572 = pi20 & n515;
  assign n573 = n377 & n523;
  assign n574 = ~pi38 & n392;
  assign n575 = ~pi50 & n574;
  assign n576 = ~pi46 & n575;
  assign n577 = n573 & n576;
  assign n578 = n374 & n577;
  assign n579 = n373 & n578;
  assign n580 = pi2 & n579;
  assign n581 = ~pi15 & n578;
  assign n582 = pi20 & ~n581;
  assign n583 = ~n580 & ~n582;
  assign n584 = pi82 & ~n583;
  assign n585 = pi82 & ~n579;
  assign n586 = ~pi71 & ~n388;
  assign n587 = ~n585 & n586;
  assign n588 = ~n572 & ~n587;
  assign n589 = ~n584 & n588;
  assign po35 = ~pi129 & ~n589;
  assign n591 = pi21 & ~pi54;
  assign n592 = ~pi4 & pi19;
  assign n593 = ~pi21 & n592;
  assign n594 = n419 & n593;
  assign n595 = n459 & n594;
  assign n596 = n451 & n595;
  assign n597 = ~n591 & ~n596;
  assign po36 = n336 & ~n597;
  assign n599 = pi22 & ~pi54;
  assign n600 = pi5 & ~pi6;
  assign n601 = ~pi14 & n600;
  assign n602 = n291 & n341;
  assign n603 = n601 & n602;
  assign n604 = n420 & n603;
  assign n605 = n468 & n604;
  assign n606 = ~n599 & ~n605;
  assign po37 = n336 & ~n606;
  assign n608 = ~pi23 & pi55;
  assign n609 = pi61 & ~pi129;
  assign po38 = ~n608 & n609;
  assign n611 = ~pi2 & n373;
  assign n612 = ~pi49 & n611;
  assign n613 = pi82 & ~n612;
  assign n614 = n388 & ~n613;
  assign n615 = n382 & n573;
  assign n616 = pi82 & ~n615;
  assign n617 = ~n614 & ~n616;
  assign n618 = ~pi24 & ~n617;
  assign n619 = pi24 & pi82;
  assign n620 = n577 & n619;
  assign n621 = ~pi45 & ~pi49;
  assign n622 = n611 & n621;
  assign n623 = n385 & n622;
  assign n624 = pi82 & ~n623;
  assign n625 = pi63 & ~n388;
  assign n626 = ~n624 & n625;
  assign n627 = ~pi129 & ~n620;
  assign n628 = ~n618 & n627;
  assign po39 = ~n626 & n628;
  assign n630 = ~pi53 & ~pi58;
  assign n631 = pi25 & ~pi116;
  assign n632 = ~pi27 & ~pi85;
  assign n633 = ~pi26 & n631;
  assign n634 = n632 & n633;
  assign n635 = ~n630 & ~n634;
  assign n636 = ~pi53 & pi58;
  assign n637 = pi53 & ~pi58;
  assign n638 = ~n636 & ~n637;
  assign n639 = pi85 & pi116;
  assign n640 = ~pi85 & ~pi110;
  assign n641 = ~pi96 & n640;
  assign n642 = ~n639 & ~n641;
  assign n643 = pi100 & ~n642;
  assign n644 = pi85 & ~pi116;
  assign n645 = pi25 & n644;
  assign n646 = ~n643 & ~n645;
  assign n647 = ~pi26 & ~n646;
  assign n648 = ~pi39 & ~pi52;
  assign n649 = ~pi51 & n648;
  assign n650 = pi116 & n649;
  assign n651 = ~pi85 & ~n650;
  assign n652 = pi26 & n651;
  assign n653 = ~pi25 & ~pi116;
  assign n654 = n652 & ~n653;
  assign n655 = ~n647 & ~n654;
  assign n656 = ~pi27 & ~n655;
  assign n657 = ~n631 & ~n650;
  assign n658 = pi27 & ~n657;
  assign n659 = ~pi95 & ~pi100;
  assign n660 = ~pi97 & n659;
  assign n661 = ~pi110 & ~n660;
  assign n662 = ~pi51 & ~pi52;
  assign n663 = ~pi39 & n662;
  assign n664 = pi27 & ~n663;
  assign n665 = pi25 & ~n661;
  assign n666 = ~n664 & n665;
  assign n667 = ~n658 & ~n666;
  assign n668 = ~pi26 & ~pi85;
  assign n669 = ~n667 & n668;
  assign n670 = ~n656 & ~n669;
  assign n671 = ~pi53 & ~n670;
  assign n672 = n638 & ~n671;
  assign n673 = n336 & ~n635;
  assign po40 = ~n672 & n673;
  assign n675 = ~pi27 & ~pi53;
  assign n676 = ~pi58 & n675;
  assign n677 = pi26 & pi116;
  assign n678 = n643 & ~n677;
  assign n679 = ~n652 & ~n678;
  assign n680 = n336 & n676;
  assign po41 = ~n679 & n680;
  assign n682 = ~pi26 & n336;
  assign n683 = pi27 & n651;
  assign n684 = pi95 & ~pi96;
  assign n685 = n640 & n684;
  assign n686 = ~n639 & ~n685;
  assign n687 = ~pi27 & ~pi100;
  assign n688 = ~n686 & n687;
  assign n689 = ~n683 & ~n688;
  assign n690 = n630 & n682;
  assign po42 = ~n689 & n690;
  assign n692 = ~pi26 & ~pi27;
  assign n693 = ~pi28 & ~pi116;
  assign n694 = pi100 & pi116;
  assign n695 = n692 & ~n693;
  assign n696 = ~n694 & n695;
  assign n697 = pi85 & ~n696;
  assign n698 = n649 & n677;
  assign n699 = ~pi26 & ~pi100;
  assign n700 = ~pi110 & n699;
  assign n701 = n684 & n700;
  assign n702 = ~n698 & ~n701;
  assign n703 = ~pi27 & ~n702;
  assign n704 = ~pi26 & ~n663;
  assign n705 = ~pi27 & n649;
  assign n706 = ~n704 & ~n705;
  assign n707 = ~n661 & ~n706;
  assign n708 = pi26 & pi27;
  assign n709 = ~n692 & ~n708;
  assign n710 = ~pi116 & n709;
  assign n711 = ~n707 & ~n710;
  assign n712 = pi28 & ~n711;
  assign n713 = ~pi26 & n664;
  assign n714 = pi116 & n713;
  assign n715 = ~pi85 & ~n703;
  assign n716 = ~n714 & n715;
  assign n717 = ~n712 & n716;
  assign n718 = ~pi53 & ~n697;
  assign n719 = ~n717 & n718;
  assign n720 = ~pi27 & pi28;
  assign n721 = ~pi116 & n720;
  assign n722 = pi53 & n668;
  assign n723 = n721 & n722;
  assign n724 = ~n719 & ~n723;
  assign n725 = ~pi58 & ~n724;
  assign n726 = ~pi26 & ~pi53;
  assign n727 = ~pi85 & n726;
  assign n728 = pi58 & n721;
  assign n729 = n727 & n728;
  assign n730 = ~n725 & ~n729;
  assign po43 = n336 & ~n730;
  assign n732 = pi29 & ~pi116;
  assign n733 = pi97 & pi116;
  assign n734 = pi58 & ~n732;
  assign n735 = ~n733 & n734;
  assign n736 = ~pi96 & ~pi110;
  assign n737 = pi97 & n659;
  assign n738 = n736 & n737;
  assign n739 = pi29 & ~n661;
  assign n740 = ~pi58 & ~n738;
  assign n741 = ~n739 & n740;
  assign n742 = ~pi53 & ~n735;
  assign n743 = ~n741 & n742;
  assign n744 = n637 & n732;
  assign n745 = ~n743 & ~n744;
  assign n746 = ~pi27 & ~n745;
  assign n747 = pi27 & n630;
  assign n748 = n732 & n747;
  assign n749 = ~n746 & ~n748;
  assign n750 = ~pi85 & ~n749;
  assign n751 = pi85 & n732;
  assign n752 = n676 & n751;
  assign n753 = ~n750 & ~n752;
  assign n754 = ~pi26 & ~n753;
  assign n755 = pi26 & ~pi27;
  assign n756 = ~pi85 & n630;
  assign n757 = n755 & n756;
  assign n758 = n732 & n757;
  assign n759 = ~n754 & ~n758;
  assign po44 = n336 & ~n759;
  assign n761 = ~pi88 & pi106;
  assign n762 = ~pi30 & ~pi109;
  assign n763 = ~pi60 & pi109;
  assign n764 = ~n762 & ~n763;
  assign n765 = ~pi106 & ~n764;
  assign n766 = ~pi129 & ~n761;
  assign po45 = ~n765 & n766;
  assign n768 = ~pi89 & pi106;
  assign n769 = ~pi31 & ~pi109;
  assign n770 = ~pi30 & pi109;
  assign n771 = ~n769 & ~n770;
  assign n772 = ~pi106 & ~n771;
  assign n773 = ~pi129 & ~n768;
  assign po46 = ~n772 & n773;
  assign n775 = ~pi99 & pi106;
  assign n776 = ~pi32 & ~pi109;
  assign n777 = ~pi31 & pi109;
  assign n778 = ~n776 & ~n777;
  assign n779 = ~pi106 & ~n778;
  assign n780 = ~pi129 & ~n775;
  assign po47 = ~n779 & n780;
  assign n782 = ~pi90 & pi106;
  assign n783 = ~pi33 & ~pi109;
  assign n784 = ~pi32 & pi109;
  assign n785 = ~n783 & ~n784;
  assign n786 = ~pi106 & ~n785;
  assign n787 = ~pi129 & ~n782;
  assign po48 = ~n786 & n787;
  assign n789 = ~pi91 & pi106;
  assign n790 = ~pi34 & ~pi109;
  assign n791 = ~pi33 & pi109;
  assign n792 = ~n790 & ~n791;
  assign n793 = ~pi106 & ~n792;
  assign n794 = ~pi129 & ~n789;
  assign po49 = ~n793 & n794;
  assign n796 = ~pi92 & pi106;
  assign n797 = ~pi35 & ~pi109;
  assign n798 = ~pi34 & pi109;
  assign n799 = ~n797 & ~n798;
  assign n800 = ~pi106 & ~n799;
  assign n801 = ~pi129 & ~n796;
  assign po50 = ~n800 & n801;
  assign n803 = ~pi98 & pi106;
  assign n804 = ~pi36 & ~pi109;
  assign n805 = ~pi35 & pi109;
  assign n806 = ~n804 & ~n805;
  assign n807 = ~pi106 & ~n806;
  assign n808 = ~pi129 & ~n803;
  assign po51 = ~n807 & n808;
  assign n810 = ~pi93 & pi106;
  assign n811 = ~pi37 & ~pi109;
  assign n812 = ~pi36 & pi109;
  assign n813 = ~n811 & ~n812;
  assign n814 = ~pi106 & ~n813;
  assign n815 = ~pi129 & ~n810;
  assign po52 = ~n814 & n815;
  assign n817 = ~pi40 & ~pi42;
  assign n818 = ~pi44 & pi82;
  assign n819 = pi38 & n817;
  assign n820 = n818 & n819;
  assign n821 = n517 & n611;
  assign n822 = ~pi48 & n821;
  assign n823 = n393 & n395;
  assign n824 = ~pi50 & n823;
  assign n825 = n822 & n824;
  assign n826 = n392 & n825;
  assign n827 = pi82 & ~n826;
  assign n828 = pi74 & ~n388;
  assign n829 = ~n827 & n828;
  assign n830 = pi82 & ~n392;
  assign n831 = n393 & n396;
  assign n832 = ~pi50 & n821;
  assign n833 = n831 & n832;
  assign n834 = pi82 & ~n833;
  assign n835 = n388 & ~n834;
  assign n836 = ~n830 & ~n835;
  assign n837 = ~pi38 & ~n836;
  assign n838 = ~pi129 & ~n820;
  assign n839 = ~n829 & n838;
  assign po53 = ~n837 & n839;
  assign n841 = pi109 & n662;
  assign n842 = pi39 & ~n841;
  assign n843 = ~pi51 & pi109;
  assign n844 = n648 & n843;
  assign n845 = ~pi106 & ~n844;
  assign n846 = ~n842 & n845;
  assign po54 = ~pi129 & ~n846;
  assign n848 = ~pi42 & n818;
  assign n849 = pi40 & n848;
  assign n850 = pi82 & ~n378;
  assign n851 = pi82 & ~n399;
  assign n852 = n388 & ~n851;
  assign n853 = ~n850 & ~n852;
  assign n854 = ~pi40 & ~n853;
  assign n855 = n522 & n821;
  assign n856 = n377 & n855;
  assign n857 = n380 & n856;
  assign n858 = n378 & n857;
  assign n859 = pi82 & ~n858;
  assign n860 = pi73 & ~n388;
  assign n861 = ~n859 & n860;
  assign n862 = ~pi129 & ~n849;
  assign n863 = ~n854 & n862;
  assign po55 = ~n861 & n863;
  assign n865 = pi41 & n848;
  assign n866 = n381 & n865;
  assign n867 = pi82 & ~n382;
  assign n868 = pi82 & ~n398;
  assign n869 = n388 & ~n868;
  assign n870 = ~n867 & ~n869;
  assign n871 = ~pi41 & ~n870;
  assign n872 = n398 & n576;
  assign n873 = pi82 & ~n872;
  assign n874 = pi76 & ~n388;
  assign n875 = ~n873 & n874;
  assign n876 = ~pi129 & ~n866;
  assign n877 = ~n871 & n876;
  assign po56 = ~n875 & n877;
  assign n879 = pi42 & n818;
  assign n880 = n817 & n857;
  assign n881 = ~n389 & ~n880;
  assign n882 = pi72 & ~n881;
  assign n883 = pi44 & pi82;
  assign n884 = ~pi40 & n857;
  assign n885 = pi82 & ~n884;
  assign n886 = n388 & ~n885;
  assign n887 = ~n883 & ~n886;
  assign n888 = ~pi42 & ~n887;
  assign n889 = ~pi129 & ~n879;
  assign n890 = ~n882 & n889;
  assign po57 = ~n888 & n890;
  assign n892 = n817 & n818;
  assign n893 = n394 & n892;
  assign n894 = pi43 & n893;
  assign n895 = pi82 & ~n518;
  assign n896 = n524 & n525;
  assign n897 = n523 & n896;
  assign n898 = pi82 & ~n897;
  assign n899 = n388 & ~n898;
  assign n900 = ~n895 & ~n899;
  assign n901 = ~pi43 & ~n900;
  assign n902 = n518 & n855;
  assign n903 = pi82 & ~n902;
  assign n904 = pi77 & ~n388;
  assign n905 = ~n903 & n904;
  assign n906 = ~pi129 & ~n894;
  assign n907 = ~n905 & n906;
  assign po58 = ~n901 & n907;
  assign n909 = pi82 & ~n880;
  assign n910 = ~pi67 & ~n388;
  assign n911 = pi44 & n388;
  assign n912 = ~n910 & ~n911;
  assign n913 = ~n909 & n912;
  assign n914 = ~pi129 & ~n883;
  assign po59 = ~n913 & n914;
  assign n916 = n575 & n831;
  assign n917 = pi45 & pi82;
  assign n918 = n916 & n917;
  assign n919 = pi82 & ~n896;
  assign n920 = n388 & ~n919;
  assign n921 = pi82 & ~n916;
  assign n922 = ~n920 & ~n921;
  assign n923 = ~pi45 & ~n922;
  assign n924 = n385 & n896;
  assign n925 = pi82 & ~n924;
  assign n926 = pi68 & ~n388;
  assign n927 = ~n925 & n926;
  assign n928 = ~pi129 & ~n918;
  assign n929 = ~n923 & n928;
  assign po60 = ~n927 & n929;
  assign n931 = ~pi75 & n389;
  assign n932 = ~pi75 & ~n388;
  assign n933 = pi82 & ~n856;
  assign n934 = ~n932 & ~n933;
  assign n935 = n576 & ~n934;
  assign n936 = pi82 & n575;
  assign n937 = pi46 & ~n389;
  assign n938 = ~n936 & n937;
  assign n939 = ~n931 & ~n938;
  assign n940 = ~n935 & n939;
  assign po61 = ~pi129 & ~n940;
  assign n942 = ~pi43 & pi47;
  assign n943 = n893 & n942;
  assign n944 = pi82 & ~n383;
  assign n945 = pi82 & ~n822;
  assign n946 = n388 & ~n945;
  assign n947 = ~n944 & ~n946;
  assign n948 = ~pi47 & ~n947;
  assign n949 = n383 & n822;
  assign n950 = pi82 & ~n949;
  assign n951 = pi64 & ~n388;
  assign n952 = ~n950 & n951;
  assign n953 = ~pi129 & ~n943;
  assign n954 = ~n948 & n953;
  assign po62 = ~n952 & n954;
  assign n956 = pi48 & n395;
  assign n957 = n893 & n956;
  assign n958 = pi82 & ~n821;
  assign n959 = n388 & ~n958;
  assign n960 = n575 & n823;
  assign n961 = pi82 & ~n960;
  assign n962 = ~n959 & ~n961;
  assign n963 = ~pi48 & ~n962;
  assign n964 = n384 & n821;
  assign n965 = pi82 & ~n964;
  assign n966 = pi62 & ~n388;
  assign n967 = ~n965 & n966;
  assign n968 = ~pi129 & ~n957;
  assign n969 = ~n963 & n968;
  assign po63 = ~n967 & n969;
  assign n971 = ~pi24 & ~pi40;
  assign n972 = n378 & n971;
  assign n973 = n380 & n972;
  assign n974 = n573 & n973;
  assign n975 = pi49 & ~n974;
  assign n976 = n578 & ~n611;
  assign n977 = ~n975 & ~n976;
  assign n978 = pi82 & ~n977;
  assign n979 = pi49 & n515;
  assign n980 = pi82 & ~n578;
  assign n981 = ~pi69 & ~n388;
  assign n982 = ~n980 & n981;
  assign n983 = ~n979 & ~n982;
  assign n984 = ~n978 & n983;
  assign po64 = ~pi129 & ~n984;
  assign n986 = pi50 & pi82;
  assign n987 = n574 & n986;
  assign n988 = pi82 & ~n574;
  assign n989 = n393 & n398;
  assign n990 = pi82 & ~n989;
  assign n991 = n388 & ~n990;
  assign n992 = ~n988 & ~n991;
  assign n993 = ~pi50 & ~n992;
  assign n994 = pi82 & ~n825;
  assign n995 = pi66 & ~n388;
  assign n996 = ~n994 & n995;
  assign n997 = ~pi129 & ~n987;
  assign n998 = ~n996 & n997;
  assign po65 = ~n993 & n998;
  assign n1000 = pi51 & ~pi109;
  assign n1001 = ~pi106 & ~n843;
  assign n1002 = ~n1000 & n1001;
  assign po66 = ~pi129 & ~n1002;
  assign n1004 = pi52 & ~n843;
  assign n1005 = ~pi106 & ~n841;
  assign n1006 = ~n1004 & n1005;
  assign po67 = ~pi129 & ~n1006;
  assign n1008 = ~pi116 & n637;
  assign n1009 = pi58 & pi116;
  assign n1010 = ~pi58 & n659;
  assign n1011 = n736 & n1010;
  assign n1012 = ~n1009 & ~n1011;
  assign n1013 = ~pi53 & pi97;
  assign n1014 = ~n1012 & n1013;
  assign n1015 = ~n1008 & ~n1014;
  assign n1016 = n632 & n682;
  assign po68 = ~n1015 & n1016;
  assign n1018 = ~n388 & n896;
  assign n1019 = n615 & n1018;
  assign n1020 = ~pi129 & ~n389;
  assign po69 = n1019 | ~n1020;
  assign po129 = pi123 | pi129;
  assign n1023 = pi114 & ~pi122;
  assign po70 = ~po129 & n1023;
  assign n1025 = ~pi26 & pi58;
  assign n1026 = ~pi58 & n677;
  assign n1027 = ~n1025 & ~n1026;
  assign n1028 = pi94 & ~n1027;
  assign n1029 = pi58 & ~pi116;
  assign n1030 = pi37 & ~pi116;
  assign n1031 = ~n1025 & ~n1030;
  assign n1032 = ~n1029 & ~n1031;
  assign n1033 = ~n1028 & ~n1032;
  assign n1034 = ~pi53 & ~n1033;
  assign n1035 = ~pi26 & pi37;
  assign n1036 = ~pi58 & n1035;
  assign n1037 = ~n1034 & ~n1036;
  assign n1038 = ~pi85 & ~n1037;
  assign n1039 = n630 & n1035;
  assign n1040 = ~n1038 & ~n1039;
  assign n1041 = ~pi27 & ~n1040;
  assign n1042 = n756 & n1035;
  assign n1043 = ~n1041 & ~n1042;
  assign po71 = n336 & ~n1043;
  assign n1045 = ~pi116 & n727;
  assign n1046 = pi85 & ~n726;
  assign n1047 = pi26 & pi53;
  assign n1048 = ~pi58 & ~n1047;
  assign n1049 = ~n1046 & n1048;
  assign n1050 = ~n1045 & ~n1049;
  assign n1051 = pi57 & ~n1050;
  assign n1052 = pi60 & n1009;
  assign n1053 = n727 & n1052;
  assign n1054 = ~n1051 & ~n1053;
  assign n1055 = ~pi27 & ~n1054;
  assign n1056 = pi57 & ~pi58;
  assign n1057 = n727 & n1056;
  assign n1058 = ~n1055 & ~n1057;
  assign po72 = n336 & ~n1058;
  assign n1060 = n692 & n1029;
  assign n1061 = ~pi58 & n709;
  assign n1062 = n650 & n1061;
  assign n1063 = ~n1060 & ~n1062;
  assign n1064 = ~pi53 & ~pi85;
  assign n1065 = n336 & n1064;
  assign po73 = ~n1063 & n1065;
  assign n1067 = ~pi59 & ~n661;
  assign n1068 = ~pi96 & n661;
  assign n1069 = n630 & ~n1067;
  assign n1070 = ~n1068 & n1069;
  assign n1071 = pi59 & ~pi116;
  assign n1072 = ~n638 & n1071;
  assign n1073 = ~n1070 & ~n1072;
  assign n1074 = ~pi85 & ~n1073;
  assign n1075 = pi85 & n630;
  assign n1076 = n1071 & n1075;
  assign n1077 = ~n1074 & ~n1076;
  assign n1078 = ~pi27 & ~n1077;
  assign n1079 = pi27 & n1071;
  assign n1080 = n756 & n1079;
  assign n1081 = ~n1078 & ~n1080;
  assign n1082 = ~pi26 & ~n1081;
  assign n1083 = n757 & n1071;
  assign n1084 = ~n1082 & ~n1083;
  assign po74 = n336 & ~n1084;
  assign n1086 = ~pi117 & ~pi122;
  assign n1087 = pi60 & ~n1086;
  assign n1088 = pi123 & n1086;
  assign po75 = n1087 | n1088;
  assign n1090 = ~pi114 & ~pi122;
  assign n1091 = pi123 & ~pi129;
  assign po76 = n1090 & n1091;
  assign n1093 = pi136 & ~pi137;
  assign n1094 = pi131 & pi132;
  assign n1095 = pi133 & n1094;
  assign n1096 = ~pi138 & n1095;
  assign n1097 = n1093 & n1096;
  assign n1098 = ~pi62 & ~n1097;
  assign n1099 = pi140 & n1097;
  assign n1100 = ~pi129 & ~n1098;
  assign po77 = n1099 | ~n1100;
  assign n1102 = ~pi63 & ~n1097;
  assign n1103 = pi142 & n1097;
  assign n1104 = ~pi129 & ~n1102;
  assign po78 = n1103 | ~n1104;
  assign n1106 = ~pi64 & ~n1097;
  assign n1107 = pi139 & n1097;
  assign n1108 = ~pi129 & ~n1106;
  assign po79 = n1107 | ~n1108;
  assign n1110 = ~pi65 & ~n1097;
  assign n1111 = pi146 & n1097;
  assign n1112 = ~pi129 & ~n1110;
  assign po80 = n1111 | ~n1112;
  assign n1114 = ~pi136 & ~pi137;
  assign n1115 = n1096 & n1114;
  assign n1116 = ~pi66 & ~n1115;
  assign n1117 = pi143 & n1115;
  assign n1118 = ~pi129 & ~n1116;
  assign po81 = n1117 | ~n1118;
  assign n1120 = ~pi67 & ~n1115;
  assign n1121 = pi139 & n1115;
  assign n1122 = ~pi129 & ~n1120;
  assign po82 = n1121 | ~n1122;
  assign n1124 = ~pi68 & ~n1097;
  assign n1125 = pi141 & n1097;
  assign n1126 = ~pi129 & ~n1124;
  assign po83 = n1125 | ~n1126;
  assign n1128 = ~pi69 & ~n1097;
  assign n1129 = pi143 & n1097;
  assign n1130 = ~pi129 & ~n1128;
  assign po84 = n1129 | ~n1130;
  assign n1132 = ~pi70 & ~n1097;
  assign n1133 = pi144 & n1097;
  assign n1134 = ~pi129 & ~n1132;
  assign po85 = n1133 | ~n1134;
  assign n1136 = ~pi71 & ~n1097;
  assign n1137 = pi145 & n1097;
  assign n1138 = ~pi129 & ~n1136;
  assign po86 = n1137 | ~n1138;
  assign n1140 = ~pi72 & ~n1115;
  assign n1141 = pi140 & n1115;
  assign n1142 = ~pi129 & ~n1140;
  assign po87 = n1141 | ~n1142;
  assign n1144 = ~pi73 & ~n1115;
  assign n1145 = pi141 & n1115;
  assign n1146 = ~pi129 & ~n1144;
  assign po88 = n1145 | ~n1146;
  assign n1148 = ~pi74 & ~n1115;
  assign n1149 = pi142 & n1115;
  assign n1150 = ~pi129 & ~n1148;
  assign po89 = n1149 | ~n1150;
  assign n1152 = ~pi75 & ~n1115;
  assign n1153 = pi144 & n1115;
  assign n1154 = ~pi129 & ~n1152;
  assign po90 = n1153 | ~n1154;
  assign n1156 = ~pi76 & ~n1115;
  assign n1157 = pi145 & n1115;
  assign n1158 = ~pi129 & ~n1156;
  assign po91 = n1157 | ~n1158;
  assign n1160 = ~pi77 & ~n1115;
  assign n1161 = pi146 & n1115;
  assign n1162 = ~pi129 & ~n1160;
  assign po92 = n1161 | ~n1162;
  assign n1164 = ~pi136 & pi137;
  assign n1165 = n1096 & n1164;
  assign n1166 = ~pi78 & ~n1165;
  assign n1167 = ~pi142 & n1165;
  assign n1168 = ~pi129 & ~n1166;
  assign po93 = ~n1167 & n1168;
  assign n1170 = ~pi79 & ~n1165;
  assign n1171 = ~pi143 & n1165;
  assign n1172 = ~pi129 & ~n1170;
  assign po94 = ~n1171 & n1172;
  assign n1174 = ~pi80 & ~n1165;
  assign n1175 = ~pi144 & n1165;
  assign n1176 = ~pi129 & ~n1174;
  assign po95 = ~n1175 & n1176;
  assign n1178 = ~pi81 & ~n1165;
  assign n1179 = ~pi145 & n1165;
  assign n1180 = ~pi129 & ~n1178;
  assign po96 = ~n1179 & n1180;
  assign n1182 = ~pi82 & ~n1165;
  assign n1183 = ~pi146 & n1165;
  assign n1184 = ~pi129 & ~n1182;
  assign po97 = ~n1183 & n1184;
  assign n1186 = pi136 & ~pi138;
  assign n1187 = pi31 & n1186;
  assign n1188 = ~pi87 & ~pi138;
  assign n1189 = pi115 & pi138;
  assign n1190 = ~pi136 & ~n1188;
  assign n1191 = ~n1189 & n1190;
  assign n1192 = ~n1187 & ~n1191;
  assign n1193 = pi137 & ~n1192;
  assign n1194 = ~pi89 & pi138;
  assign n1195 = pi62 & ~pi138;
  assign n1196 = pi136 & ~n1194;
  assign n1197 = ~n1195 & n1196;
  assign n1198 = ~pi119 & pi138;
  assign n1199 = pi72 & ~pi138;
  assign n1200 = ~pi136 & ~n1198;
  assign n1201 = ~n1199 & n1200;
  assign n1202 = ~n1197 & ~n1201;
  assign n1203 = ~pi137 & ~n1202;
  assign po98 = n1193 | n1203;
  assign n1205 = ~pi84 & ~n1165;
  assign n1206 = ~pi141 & n1165;
  assign n1207 = ~pi129 & ~n1205;
  assign po99 = ~n1206 & n1207;
  assign n1209 = n640 & ~n660;
  assign n1210 = pi96 & n1209;
  assign n1211 = ~n644 & ~n1210;
  assign n1212 = n676 & n682;
  assign po100 = ~n1211 & n1212;
  assign n1214 = ~pi86 & ~n1165;
  assign n1215 = ~pi139 & n1165;
  assign n1216 = ~pi129 & ~n1214;
  assign po101 = ~n1215 & n1216;
  assign n1218 = ~pi87 & ~n1165;
  assign n1219 = ~pi140 & n1165;
  assign n1220 = ~pi129 & ~n1218;
  assign po102 = ~n1219 & n1220;
  assign n1222 = pi137 & n1186;
  assign n1223 = n1095 & n1222;
  assign n1224 = ~pi88 & ~n1223;
  assign n1225 = ~pi139 & n1223;
  assign n1226 = ~pi129 & ~n1224;
  assign po103 = ~n1225 & n1226;
  assign n1228 = ~pi89 & ~n1223;
  assign n1229 = ~pi140 & n1223;
  assign n1230 = ~pi129 & ~n1228;
  assign po104 = ~n1229 & n1230;
  assign n1232 = ~pi90 & ~n1223;
  assign n1233 = ~pi142 & n1223;
  assign n1234 = ~pi129 & ~n1232;
  assign po105 = ~n1233 & n1234;
  assign n1236 = ~pi91 & ~n1223;
  assign n1237 = ~pi143 & n1223;
  assign n1238 = ~pi129 & ~n1236;
  assign po106 = ~n1237 & n1238;
  assign n1240 = ~pi92 & ~n1223;
  assign n1241 = ~pi144 & n1223;
  assign n1242 = ~pi129 & ~n1240;
  assign po107 = ~n1241 & n1242;
  assign n1244 = ~pi93 & ~n1223;
  assign n1245 = ~pi146 & n1223;
  assign n1246 = ~pi129 & ~n1244;
  assign po108 = ~n1245 & n1246;
  assign n1248 = pi82 & pi138;
  assign n1249 = n1114 & n1248;
  assign n1250 = n1095 & n1249;
  assign n1251 = ~pi94 & ~n1250;
  assign n1252 = ~pi142 & n1250;
  assign n1253 = ~pi129 & ~n1251;
  assign po109 = ~n1252 & n1253;
  assign n1255 = ~pi3 & ~pi110;
  assign n1256 = ~n1095 & ~n1255;
  assign n1257 = ~n1250 & ~n1256;
  assign n1258 = pi95 & n1257;
  assign n1259 = pi143 & n1250;
  assign n1260 = ~n1258 & ~n1259;
  assign po110 = ~pi129 & ~n1260;
  assign n1262 = pi96 & n1257;
  assign n1263 = pi146 & n1250;
  assign n1264 = ~n1262 & ~n1263;
  assign po111 = ~pi129 & ~n1264;
  assign n1266 = pi97 & n1257;
  assign n1267 = pi145 & n1250;
  assign n1268 = ~n1266 & ~n1267;
  assign po112 = ~pi129 & ~n1268;
  assign n1270 = ~pi98 & ~n1223;
  assign n1271 = ~pi145 & n1223;
  assign n1272 = ~pi129 & ~n1270;
  assign po113 = ~n1271 & n1272;
  assign n1274 = ~pi99 & ~n1223;
  assign n1275 = ~pi141 & n1223;
  assign n1276 = ~pi129 & ~n1274;
  assign po114 = ~n1275 & n1276;
  assign n1278 = pi100 & n1257;
  assign n1279 = pi144 & n1250;
  assign n1280 = ~n1278 & ~n1279;
  assign po115 = ~pi129 & ~n1280;
  assign n1282 = pi37 & n1186;
  assign n1283 = ~pi82 & ~pi138;
  assign n1284 = ~pi96 & pi138;
  assign n1285 = ~pi136 & ~n1283;
  assign n1286 = ~n1284 & n1285;
  assign n1287 = ~n1282 & ~n1286;
  assign n1288 = pi137 & ~n1287;
  assign n1289 = ~pi93 & pi138;
  assign n1290 = pi65 & ~pi138;
  assign n1291 = pi136 & ~n1289;
  assign n1292 = ~n1290 & n1291;
  assign n1293 = ~pi124 & pi138;
  assign n1294 = pi77 & ~pi138;
  assign n1295 = ~pi136 & ~n1293;
  assign n1296 = ~n1294 & n1295;
  assign n1297 = ~n1292 & ~n1296;
  assign n1298 = ~pi137 & ~n1297;
  assign po116 = n1288 | n1298;
  assign n1300 = pi91 & n1093;
  assign n1301 = pi95 & n1164;
  assign n1302 = ~n1300 & ~n1301;
  assign n1303 = pi138 & ~n1302;
  assign n1304 = ~pi79 & ~pi136;
  assign n1305 = ~pi34 & pi136;
  assign n1306 = pi137 & ~n1304;
  assign n1307 = ~n1305 & n1306;
  assign n1308 = pi66 & ~pi136;
  assign n1309 = pi69 & pi136;
  assign n1310 = ~pi137 & ~n1308;
  assign n1311 = ~n1309 & n1310;
  assign n1312 = ~n1307 & ~n1311;
  assign n1313 = ~pi138 & ~n1312;
  assign po117 = n1303 | n1313;
  assign n1315 = pi90 & n1093;
  assign n1316 = pi94 & n1164;
  assign n1317 = ~n1315 & ~n1316;
  assign n1318 = pi138 & ~n1317;
  assign n1319 = ~pi78 & ~pi136;
  assign n1320 = ~pi33 & pi136;
  assign n1321 = pi137 & ~n1319;
  assign n1322 = ~n1320 & n1321;
  assign n1323 = pi74 & ~pi136;
  assign n1324 = pi63 & pi136;
  assign n1325 = ~pi137 & ~n1323;
  assign n1326 = ~n1324 & n1325;
  assign n1327 = ~n1322 & ~n1326;
  assign n1328 = ~pi138 & ~n1327;
  assign po118 = n1318 | n1328;
  assign n1330 = pi99 & n1093;
  assign n1331 = ~pi112 & n1164;
  assign n1332 = ~n1330 & ~n1331;
  assign n1333 = pi138 & ~n1332;
  assign n1334 = ~pi84 & ~pi136;
  assign n1335 = ~pi32 & pi136;
  assign n1336 = pi137 & ~n1334;
  assign n1337 = ~n1335 & n1336;
  assign n1338 = pi73 & ~pi136;
  assign n1339 = pi68 & pi136;
  assign n1340 = ~pi137 & ~n1338;
  assign n1341 = ~n1339 & n1340;
  assign n1342 = ~n1337 & ~n1341;
  assign n1343 = ~pi138 & ~n1342;
  assign po119 = n1333 | n1343;
  assign n1345 = pi35 & n1186;
  assign n1346 = ~pi80 & ~pi138;
  assign n1347 = ~pi100 & pi138;
  assign n1348 = ~pi136 & ~n1346;
  assign n1349 = ~n1347 & n1348;
  assign n1350 = ~n1345 & ~n1349;
  assign n1351 = pi137 & ~n1350;
  assign n1352 = ~pi92 & pi138;
  assign n1353 = pi70 & ~pi138;
  assign n1354 = pi136 & ~n1352;
  assign n1355 = ~n1353 & n1354;
  assign n1356 = ~pi125 & pi138;
  assign n1357 = pi75 & ~pi138;
  assign n1358 = ~pi136 & ~n1356;
  assign n1359 = ~n1357 & n1358;
  assign n1360 = ~n1355 & ~n1359;
  assign n1361 = ~pi137 & ~n1360;
  assign po120 = n1351 | n1361;
  assign n1363 = ~pi26 & n676;
  assign n1364 = n1209 & n1363;
  assign n1365 = ~n639 & ~n1364;
  assign po121 = n336 & ~n1365;
  assign n1367 = pi36 & n1186;
  assign n1368 = ~pi81 & ~pi138;
  assign n1369 = ~pi97 & pi138;
  assign n1370 = ~pi136 & ~n1368;
  assign n1371 = ~n1369 & n1370;
  assign n1372 = ~n1367 & ~n1371;
  assign n1373 = pi137 & ~n1372;
  assign n1374 = ~pi98 & pi138;
  assign n1375 = pi71 & ~pi138;
  assign n1376 = pi136 & ~n1374;
  assign n1377 = ~n1375 & n1376;
  assign n1378 = ~pi23 & pi138;
  assign n1379 = pi76 & ~pi138;
  assign n1380 = ~pi136 & ~n1378;
  assign n1381 = ~n1379 & n1380;
  assign n1382 = ~n1377 & ~n1381;
  assign n1383 = ~pi137 & ~n1382;
  assign po122 = n1373 | n1383;
  assign n1385 = pi30 & n1186;
  assign n1386 = ~pi86 & ~pi138;
  assign n1387 = ~pi111 & pi138;
  assign n1388 = ~pi136 & ~n1386;
  assign n1389 = ~n1387 & n1388;
  assign n1390 = ~n1385 & ~n1389;
  assign n1391 = pi137 & ~n1390;
  assign n1392 = ~pi88 & pi138;
  assign n1393 = pi64 & ~pi138;
  assign n1394 = pi136 & ~n1392;
  assign n1395 = ~n1393 & n1394;
  assign n1396 = ~pi120 & pi138;
  assign n1397 = pi67 & ~pi138;
  assign n1398 = ~pi136 & ~n1396;
  assign n1399 = ~n1397 & n1398;
  assign n1400 = ~n1395 & ~n1399;
  assign n1401 = ~pi137 & ~n1400;
  assign po123 = n1391 | n1401;
  assign n1403 = ~n713 & ~n755;
  assign n1404 = pi116 & n336;
  assign po124 = ~n1403 & n1404;
  assign n1406 = ~pi97 & n636;
  assign n1407 = ~n637 & ~n1406;
  assign po125 = n1404 & ~n1407;
  assign n1409 = ~pi129 & n1095;
  assign n1410 = ~pi111 & ~n1249;
  assign n1411 = ~pi139 & n1249;
  assign n1412 = n1409 & ~n1410;
  assign po126 = ~n1411 & n1412;
  assign n1414 = ~pi141 & n1249;
  assign n1415 = pi112 & ~n1249;
  assign n1416 = n1409 & ~n1414;
  assign po127 = ~n1415 & n1416;
  assign n1418 = ~pi54 & pi113;
  assign n1419 = ~pi11 & ~pi22;
  assign n1420 = pi54 & n1419;
  assign n1421 = n336 & ~n1418;
  assign po128 = ~n1420 & n1421;
  assign n1423 = ~pi140 & n1249;
  assign n1424 = pi115 & ~n1249;
  assign n1425 = n1409 & ~n1423;
  assign po130 = ~n1424 & n1425;
  assign n1427 = ~pi4 & ~pi7;
  assign n1428 = ~pi9 & ~pi12;
  assign n1429 = n1427 & n1428;
  assign n1430 = pi54 & n336;
  assign po131 = ~n1429 & n1430;
  assign po132 = ~pi122 | pi129;
  assign n1433 = ~pi54 & pi118;
  assign n1434 = pi54 & ~pi59;
  assign n1435 = n501 & n1434;
  assign n1436 = ~n1433 & ~n1435;
  assign po133 = ~pi129 & ~n1436;
  assign po134 = ~pi129 & ~n659;
  assign n1439 = ~pi120 & n1255;
  assign n1440 = ~pi111 & ~pi129;
  assign po135 = ~n1439 & n1440;
  assign n1442 = pi81 & pi120;
  assign po136 = ~pi129 & n1442;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi57 & ~pi129;
  assign n1447 = ~pi96 & pi125;
  assign n1448 = ~pi3 & ~n1447;
  assign po140 = ~pi129 & ~n1448;
  assign n1450 = ~pi126 & pi132;
  assign po141 = pi133 & n1450;
  assign po12 = 1'b1;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
endmodule
