module top ( 
    pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 , pi8 ,
    pi9 , pi10 ,
    po0 , po1 , po2 , po3 , po4 , po5 , po6   );
  input  pi0 , pi1 , pi2 , pi3 , pi4 , pi5 , pi6 , pi7 ,
    pi8 , pi9 , pi10 ;
  output po0 , po1 , po2 , po3 , po4 , po5 , po6 ;
  wire n19, n20, n21, n22, n23, n24, n25,
    n26, n27, n28, n29, n30, n31, n32, n33,
    n34, n35, n36, n37, n38, n39, n40, n41,
    n42, n43, n44, n45, n46, n47, n48, n49,
    n50, n51, n52, n53, n54, n55, n56, n57,
    n58, n59, n60, n61, n62, n63, n64, n65,
    n66, n67, n68, n69, n70, n71, n72, n73,
    n74, n75, n76, n77, n79, n80, n81, n82,
    n83, n84, n85, n86, n87, n88, n89, n90,
    n91, n92, n93, n94, n95, n96, n97, n98,
    n99, n100, n101, n102, n103, n104, n105,
    n106, n107, n108, n109, n110, n111, n112,
    n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126,
    n127, n128, n129, n130, n131, n132, n133,
    n134, n135, n137, n138, n139, n140, n141,
    n142, n143, n144, n145, n146, n147, n148,
    n149, n150, n151, n152, n153, n154, n155,
    n156, n157, n158, n159, n160, n161, n162,
    n163, n164, n165, n166, n167, n168, n169,
    n170, n171, n172, n173, n174, n175, n176,
    n177, n178, n179, n180, n181, n182, n183,
    n184, n186, n187, n188, n189, n190, n191,
    n192, n193, n194, n195, n197, n198, n199,
    n200, n201, n202, n203, n204, n205, n206,
    n207, n208, n209, n210, n211, n212, n213,
    n214, n216, n217, n218, n219, n220, n221,
    n222, n223, n224, n225;
  assign n19 = ~pi6  & pi7 ;
  assign n20 = pi10  & n19;
  assign n21 = ~pi8  & ~pi9 ;
  assign n22 = ~pi2  & pi3 ;
  assign n23 = pi3  & ~pi8 ;
  assign n24 = ~pi2  & ~pi3 ;
  assign n25 = ~n23 & ~n24;
  assign n26 = ~n22 & ~n25;
  assign n27 = n21 & ~n26;
  assign n28 = ~pi10  & ~n27;
  assign n29 = ~pi7  & ~n28;
  assign n30 = pi8  & pi10 ;
  assign n31 = pi9  & n30;
  assign n32 = ~n29 & ~n31;
  assign n33 = pi6  & ~n32;
  assign n34 = ~pi5  & pi6 ;
  assign n35 = pi9  & n34;
  assign n36 = pi5  & ~pi6 ;
  assign n37 = ~pi7  & ~pi8 ;
  assign n38 = ~pi1  & pi2 ;
  assign n39 = n37 & n38;
  assign n40 = ~pi4  & pi7 ;
  assign n41 = pi3  & pi4 ;
  assign n42 = pi4  & pi8 ;
  assign n43 = pi1  & ~pi2 ;
  assign n44 = ~n40 & n43;
  assign n45 = ~n41 & ~n42;
  assign n46 = n44 & n45;
  assign n47 = ~pi9  & ~n39;
  assign n48 = ~n46 & n47;
  assign n49 = n36 & ~n48;
  assign n50 = ~pi2  & ~pi7 ;
  assign n51 = pi1  & pi5 ;
  assign n52 = n50 & n51;
  assign n53 = ~n40 & ~n52;
  assign n54 = pi3  & ~n53;
  assign n55 = ~pi3  & pi4 ;
  assign n56 = pi7  & n55;
  assign n57 = ~n54 & ~n56;
  assign n58 = ~pi8  & ~n57;
  assign n59 = ~pi4  & pi5 ;
  assign n60 = pi8  & n59;
  assign n61 = pi1  & pi4 ;
  assign n62 = ~pi4  & pi8 ;
  assign n63 = ~n61 & ~n62;
  assign n64 = pi0  & ~n63;
  assign n65 = ~pi0  & ~n61;
  assign n66 = ~pi6  & ~pi7 ;
  assign n67 = ~n65 & n66;
  assign n68 = ~n64 & n67;
  assign n69 = ~n42 & ~n68;
  assign n70 = ~pi5  & ~n69;
  assign n71 = ~n58 & ~n60;
  assign n72 = ~n70 & n71;
  assign n73 = ~pi9  & ~n72;
  assign n74 = ~n35 & ~n49;
  assign n75 = ~n73 & n74;
  assign n76 = ~pi10  & ~n75;
  assign n77 = ~n20 & ~n33;
  assign po0  = n76 | ~n77;
  assign n79 = pi6  & pi7 ;
  assign n80 = ~pi9  & n79;
  assign n81 = n30 & n80;
  assign n82 = ~pi7  & pi9 ;
  assign n83 = ~pi9  & n62;
  assign n84 = ~n82 & ~n83;
  assign n85 = ~pi6  & ~n84;
  assign n86 = ~pi4  & ~pi6 ;
  assign n87 = pi1  & pi2 ;
  assign n88 = ~pi7  & n87;
  assign n89 = n86 & n88;
  assign n90 = ~pi4  & ~pi9 ;
  assign n91 = ~n50 & ~n90;
  assign n92 = n21 & ~n39;
  assign n93 = n91 & n92;
  assign n94 = ~n89 & ~n93;
  assign n95 = pi3  & ~n94;
  assign n96 = pi6  & ~n21;
  assign n97 = n84 & n96;
  assign n98 = ~n95 & ~n97;
  assign n99 = pi5  & ~n98;
  assign n100 = ~pi1  & ~n91;
  assign n101 = pi8  & ~pi9 ;
  assign n102 = ~pi0  & pi2 ;
  assign n103 = pi0  & ~n87;
  assign n104 = pi4  & ~pi7 ;
  assign n105 = ~n102 & n104;
  assign n106 = ~n103 & n105;
  assign n107 = ~n100 & ~n101;
  assign n108 = ~n106 & n107;
  assign n109 = ~pi6  & ~n108;
  assign n110 = pi7  & n21;
  assign n111 = ~n41 & n110;
  assign n112 = ~n82 & ~n111;
  assign n113 = ~n109 & n112;
  assign n114 = ~pi5  & ~n113;
  assign n115 = ~n85 & ~n99;
  assign n116 = ~n114 & n115;
  assign n117 = ~pi10  & ~n116;
  assign n118 = pi6  & ~pi9 ;
  assign n119 = ~pi4  & n118;
  assign n120 = ~pi3  & pi5 ;
  assign n121 = ~pi6  & n120;
  assign n122 = ~n119 & ~n121;
  assign n123 = ~pi2  & ~n122;
  assign n124 = pi2  & n41;
  assign n125 = n118 & n124;
  assign n126 = ~pi1  & n36;
  assign n127 = ~n119 & ~n126;
  assign n128 = ~pi3  & ~n127;
  assign n129 = ~n123 & ~n125;
  assign n130 = ~n128 & n129;
  assign n131 = ~pi7  & ~n130;
  assign n132 = ~pi10  & ~n131;
  assign n133 = ~pi8  & ~n79;
  assign n134 = ~n132 & n133;
  assign n135 = ~n81 & ~n134;
  assign po1  = ~n117 & n135;
  assign n137 = pi4  & pi5 ;
  assign n138 = n79 & ~n137;
  assign n139 = pi3  & n19;
  assign n140 = pi6  & ~pi7 ;
  assign n141 = ~pi2  & n140;
  assign n142 = ~n139 & ~n141;
  assign n143 = n137 & ~n142;
  assign n144 = pi5  & pi6 ;
  assign n145 = ~n41 & n144;
  assign n146 = pi2  & n34;
  assign n147 = ~n126 & ~n146;
  assign n148 = n41 & ~n147;
  assign n149 = pi3  & n59;
  assign n150 = pi0  & ~pi6 ;
  assign n151 = n55 & n150;
  assign n152 = ~n149 & ~n151;
  assign n153 = pi1  & ~n152;
  assign n154 = pi0  & pi1 ;
  assign n155 = n41 & ~n154;
  assign n156 = ~n86 & ~n155;
  assign n157 = ~pi5  & ~n156;
  assign n158 = ~n153 & ~n157;
  assign n159 = pi2  & ~n158;
  assign n160 = ~pi6  & n22;
  assign n161 = ~n120 & ~n160;
  assign n162 = pi4  & ~n161;
  assign n163 = ~n159 & ~n162;
  assign n164 = ~pi7  & ~n163;
  assign n165 = ~n145 & ~n148;
  assign n166 = ~n164 & n165;
  assign n167 = ~pi8  & ~n166;
  assign n168 = ~n138 & ~n143;
  assign n169 = ~n167 & n168;
  assign n170 = ~pi9  & ~n169;
  assign n171 = n137 & n140;
  assign n172 = ~n19 & ~n171;
  assign n173 = pi8  & ~n172;
  assign n174 = ~n170 & ~n173;
  assign n175 = ~pi10  & ~n174;
  assign n176 = pi5  & ~pi8 ;
  assign n177 = pi9  & n176;
  assign n178 = ~n30 & ~n177;
  assign n179 = n79 & ~n178;
  assign n180 = pi5  & pi7 ;
  assign n181 = pi8  & ~n180;
  assign n182 = ~pi10  & ~n181;
  assign n183 = pi9  & ~n182;
  assign n184 = ~n179 & ~n183;
  assign po2  = n175 | ~n184;
  assign n186 = ~pi9  & ~pi10 ;
  assign n187 = pi7  & n144;
  assign n188 = ~pi2  & n42;
  assign n189 = n187 & n188;
  assign n190 = ~pi5  & ~pi6 ;
  assign n191 = ~pi4  & ~pi7 ;
  assign n192 = ~pi8  & n191;
  assign n193 = n190 & n192;
  assign n194 = ~n189 & ~n193;
  assign n195 = ~pi3  & n186;
  assign po3  = n194 | ~n195;
  assign n197 = pi8  & n187;
  assign n198 = pi9  & ~n197;
  assign n199 = ~n88 & ~n144;
  assign n200 = pi3  & ~n199;
  assign n201 = ~pi5  & ~pi7 ;
  assign n202 = ~n200 & ~n201;
  assign n203 = pi4  & ~n202;
  assign n204 = ~n140 & ~n203;
  assign n205 = n154 & n190;
  assign n206 = ~n171 & ~n205;
  assign n207 = pi2  & pi3 ;
  assign n208 = ~n206 & n207;
  assign n209 = ~n204 & ~n208;
  assign n210 = ~pi8  & ~n209;
  assign n211 = n25 & n137;
  assign n212 = n80 & n211;
  assign n213 = ~n198 & ~n212;
  assign n214 = ~n210 & n213;
  assign po4  = pi10  | n214;
  assign n216 = n124 & n144;
  assign n217 = n37 & ~n216;
  assign n218 = ~n190 & n217;
  assign n219 = ~n24 & n197;
  assign n220 = pi2  & n23;
  assign n221 = n154 & n201;
  assign n222 = n220 & n221;
  assign n223 = ~n219 & ~n222;
  assign n224 = pi4  & ~n223;
  assign n225 = n186 & ~n218;
  assign po5  = n224 | ~n225;
  assign po6  = ~n186 | ~n217;
endmodule
