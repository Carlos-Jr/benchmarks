module i2c ( 
    pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8, pi9,
    pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18, pi19,
    pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28, pi29,
    pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38, pi39,
    pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48, pi49,
    pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58, pi59,
    pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68, pi69,
    pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78, pi79,
    pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88, pi89,
    pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98, pi99,
    pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108, pi109,
    pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118, pi119,
    pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128, pi129,
    pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138, pi139,
    pi140, pi141, pi142, pi143, pi144, pi145, pi146,
    po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141  );
  input  pi0, pi1, pi2, pi3, pi4, pi5, pi6, pi7, pi8,
    pi9, pi10, pi11, pi12, pi13, pi14, pi15, pi16, pi17, pi18,
    pi19, pi20, pi21, pi22, pi23, pi24, pi25, pi26, pi27, pi28,
    pi29, pi30, pi31, pi32, pi33, pi34, pi35, pi36, pi37, pi38,
    pi39, pi40, pi41, pi42, pi43, pi44, pi45, pi46, pi47, pi48,
    pi49, pi50, pi51, pi52, pi53, pi54, pi55, pi56, pi57, pi58,
    pi59, pi60, pi61, pi62, pi63, pi64, pi65, pi66, pi67, pi68,
    pi69, pi70, pi71, pi72, pi73, pi74, pi75, pi76, pi77, pi78,
    pi79, pi80, pi81, pi82, pi83, pi84, pi85, pi86, pi87, pi88,
    pi89, pi90, pi91, pi92, pi93, pi94, pi95, pi96, pi97, pi98,
    pi99, pi100, pi101, pi102, pi103, pi104, pi105, pi106, pi107, pi108,
    pi109, pi110, pi111, pi112, pi113, pi114, pi115, pi116, pi117, pi118,
    pi119, pi120, pi121, pi122, pi123, pi124, pi125, pi126, pi127, pi128,
    pi129, pi130, pi131, pi132, pi133, pi134, pi135, pi136, pi137, pi138,
    pi139, pi140, pi141, pi142, pi143, pi144, pi145, pi146;
  output po0, po1, po2, po3, po4, po5, po6, po7, po8, po9,
    po10, po11, po12, po13, po14, po15, po16, po17, po18, po19,
    po20, po21, po22, po23, po24, po25, po26, po27, po28, po29,
    po30, po31, po32, po33, po34, po35, po36, po37, po38, po39,
    po40, po41, po42, po43, po44, po45, po46, po47, po48, po49,
    po50, po51, po52, po53, po54, po55, po56, po57, po58, po59,
    po60, po61, po62, po63, po64, po65, po66, po67, po68, po69,
    po70, po71, po72, po73, po74, po75, po76, po77, po78, po79,
    po80, po81, po82, po83, po84, po85, po86, po87, po88, po89,
    po90, po91, po92, po93, po94, po95, po96, po97, po98, po99,
    po100, po101, po102, po103, po104, po105, po106, po107, po108, po109,
    po110, po111, po112, po113, po114, po115, po116, po117, po118, po119,
    po120, po121, po122, po123, po124, po125, po126, po127, po128, po129,
    po130, po131, po132, po133, po134, po135, po136, po137, po138, po139,
    po140, po141;
  wire n291, n292, n293, n294, n295, n296, n297,
    n298, n299, n300, n301, n302, n303, n304,
    n305, n306, n307, n308, n309, n310, n311,
    n312, n313, n314, n315, n316, n317, n318,
    n319, n320, n321, n322, n323, n324, n325,
    n326, n327, n328, n329, n330, n331, n332,
    n333, n334, n335, n336, n337, n339, n340,
    n341, n342, n343, n344, n345, n346, n347,
    n348, n349, n350, n351, n352, n353, n354,
    n355, n356, n357, n358, n359, n360, n361,
    n362, n363, n364, n365, n366, n368, n369,
    n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383,
    n384, n385, n386, n387, n388, n389, n390,
    n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n403, n404, n405,
    n406, n407, n408, n409, n410, n411, n412,
    n414, n415, n416, n417, n418, n419, n420,
    n422, n423, n424, n425, n426, n427, n428,
    n429, n430, n431, n432, n433, n434, n436,
    n437, n438, n439, n440, n441, n442, n444,
    n445, n446, n447, n448, n449, n450, n451,
    n453, n454, n455, n456, n457, n458, n459,
    n460, n461, n462, n463, n465, n466, n467,
    n468, n469, n470, n472, n473, n474, n475,
    n476, n477, n479, n480, n481, n482, n483,
    n484, n485, n486, n488, n489, n490, n491,
    n492, n494, n495, n496, n497, n498, n499,
    n500, n502, n503, n504, n505, n507, n508,
    n509, n510, n511, n512, n513, n514, n515,
    n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n529, n530,
    n531, n532, n533, n534, n536, n537, n538,
    n539, n540, n541, n542, n543, n544, n546,
    n547, n548, n549, n550, n552, n553, n554,
    n555, n556, n558, n559, n560, n561, n562,
    n563, n564, n565, n566, n567, n568, n570,
    n571, n572, n573, n574, n575, n577, n578,
    n579, n580, n582, n583, n585, n586, n587,
    n588, n589, n590, n591, n592, n593, n594,
    n595, n596, n597, n598, n599, n601, n602,
    n603, n604, n605, n606, n607, n608, n609,
    n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623,
    n624, n625, n626, n627, n628, n629, n630,
    n631, n632, n633, n634, n635, n636, n637,
    n638, n640, n641, n642, n643, n644, n645,
    n646, n648, n649, n650, n651, n652, n653,
    n654, n655, n656, n658, n659, n660, n661,
    n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675,
    n676, n677, n678, n679, n680, n681, n682,
    n683, n684, n685, n686, n687, n688, n689,
    n691, n692, n693, n694, n695, n696, n697,
    n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711,
    n712, n713, n714, n715, n716, n717, n719,
    n720, n721, n722, n723, n724, n726, n727,
    n728, n729, n730, n731, n733, n734, n735,
    n736, n737, n738, n740, n741, n742, n743,
    n744, n745, n747, n748, n749, n750, n751,
    n752, n754, n755, n756, n757, n758, n759,
    n761, n762, n763, n764, n765, n766, n768,
    n769, n770, n771, n772, n773, n775, n776,
    n777, n778, n779, n780, n781, n782, n783,
    n784, n785, n786, n787, n788, n789, n790,
    n791, n792, n793, n794, n796, n797, n798,
    n799, n800, n801, n802, n804, n805, n806,
    n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n821,
    n822, n823, n824, n825, n826, n827, n828,
    n829, n830, n831, n832, n833, n835, n836,
    n837, n838, n839, n840, n841, n842, n844,
    n845, n846, n847, n848, n849, n850, n851,
    n853, n854, n855, n856, n857, n858, n859,
    n861, n862, n863, n864, n865, n866, n867,
    n869, n870, n871, n872, n873, n874, n875,
    n877, n878, n879, n880, n881, n882, n883,
    n884, n886, n887, n888, n889, n890, n891,
    n892, n893, n895, n896, n897, n898, n899,
    n900, n901, n902, n903, n905, n906, n907,
    n908, n909, n911, n912, n913, n915, n916,
    n917, n919, n920, n921, n925, n927, n928,
    n929, n930, n931, n932, n933, n934, n935,
    n936, n937, n938, n939, n940, n941, n942,
    n943, n944, n945, n947, n948, n949, n950,
    n951, n952, n953, n954, n955, n956, n957,
    n958, n959, n960, n962, n963, n964, n965,
    n966, n967, n968, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980,
    n981, n982, n983, n984, n985, n987, n988,
    n989, n991, n992, n994, n995, n996, n997,
    n998, n999, n1000, n1001, n1003, n1004,
    n1005, n1007, n1008, n1009, n1011, n1012,
    n1013, n1015, n1016, n1017, n1018, n1019,
    n1021, n1022, n1023, n1025, n1026, n1027,
    n1029, n1030, n1031, n1033, n1034, n1035,
    n1037, n1038, n1039, n1041, n1042, n1043,
    n1045, n1046, n1047, n1049, n1050, n1051,
    n1053, n1054, n1055, n1057, n1058, n1059,
    n1061, n1062, n1063, n1065, n1066, n1067,
    n1068, n1069, n1071, n1072, n1073, n1075,
    n1076, n1077, n1079, n1080, n1081, n1083,
    n1084, n1085, n1087, n1088, n1089, n1090,
    n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102,
    n1103, n1104, n1106, n1107, n1108, n1110,
    n1111, n1112, n1114, n1115, n1116, n1118,
    n1119, n1120, n1122, n1123, n1124, n1125,
    n1126, n1128, n1129, n1130, n1132, n1133,
    n1134, n1136, n1137, n1138, n1140, n1141,
    n1142, n1144, n1145, n1146, n1148, n1149,
    n1150, n1151, n1152, n1153, n1155, n1156,
    n1157, n1158, n1159, n1160, n1162, n1163,
    n1164, n1166, n1167, n1168, n1170, n1171,
    n1172, n1174, n1175, n1176, n1178, n1179,
    n1180, n1182, n1183, n1184, n1185, n1186,
    n1187, n1188, n1189, n1190, n1191, n1192,
    n1193, n1194, n1195, n1196, n1197, n1198,
    n1200, n1201, n1202, n1203, n1204, n1205,
    n1206, n1207, n1208, n1209, n1210, n1211,
    n1212, n1213, n1215, n1216, n1217, n1218,
    n1219, n1220, n1221, n1222, n1223, n1224,
    n1225, n1226, n1227, n1228, n1230, n1231,
    n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1240, n1241, n1242, n1243,
    n1245, n1246, n1247, n1248, n1249, n1250,
    n1251, n1252, n1253, n1254, n1255, n1256,
    n1257, n1258, n1259, n1260, n1261, n1263,
    n1264, n1265, n1267, n1268, n1269, n1270,
    n1271, n1272, n1273, n1274, n1275, n1276,
    n1277, n1278, n1279, n1280, n1281, n1282,
    n1283, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295,
    n1296, n1297, n1298, n1299, n1300, n1301,
    n1303, n1304, n1305, n1307, n1308, n1310,
    n1311, n1312, n1313, n1315, n1316, n1317,
    n1319, n1320, n1321, n1322, n1324, n1325,
    n1326, n1328, n1329, n1330, n1333, n1334,
    n1335, n1336, n1339, n1340, n1342, n1347,
    n1348, n1350;
  assign n291 = ~pi4 & ~pi19;
  assign n292 = ~pi18 & n291;
  assign n293 = ~pi16 & n292;
  assign n294 = ~pi8 & ~pi21;
  assign n295 = ~pi11 & n294;
  assign n296 = ~pi17 & n295;
  assign n297 = ~pi6 & ~pi9;
  assign n298 = n296 & n297;
  assign n299 = ~pi5 & ~pi22;
  assign n300 = ~pi7 & ~pi12;
  assign n301 = ~pi13 & ~pi14;
  assign n302 = n299 & n301;
  assign n303 = n300 & n302;
  assign n304 = n293 & n303;
  assign n305 = n298 & n304;
  assign n306 = pi54 & ~n305;
  assign n307 = ~pi0 & ~n306;
  assign n308 = ~pi9 & ~pi11;
  assign n309 = ~pi56 & ~n299;
  assign n310 = ~pi7 & ~pi13;
  assign n311 = n294 & n310;
  assign n312 = ~pi10 & n311;
  assign n313 = pi14 & ~n312;
  assign n314 = ~pi14 & n312;
  assign n315 = ~pi7 & n294;
  assign n316 = pi8 & pi21;
  assign n317 = pi7 & ~n294;
  assign n318 = ~pi13 & ~n316;
  assign n319 = ~n317 & n318;
  assign n320 = ~n315 & ~n319;
  assign n321 = ~pi10 & ~n320;
  assign n322 = ~n311 & ~n321;
  assign n323 = ~pi6 & ~pi12;
  assign n324 = ~pi17 & n299;
  assign n325 = n323 & n324;
  assign n326 = n293 & n325;
  assign n327 = ~n313 & n326;
  assign n328 = ~n314 & n327;
  assign n329 = ~n322 & n328;
  assign n330 = ~n309 & ~n329;
  assign n331 = n308 & ~n330;
  assign n332 = ~pi56 & n299;
  assign n333 = ~n308 & n332;
  assign n334 = ~n331 & ~n333;
  assign n335 = pi54 & ~n334;
  assign n336 = ~n307 & ~n335;
  assign n337 = ~pi3 & ~pi129;
  assign po15 = n336 | ~n337;
  assign n339 = ~pi17 & pi54;
  assign n340 = ~pi10 & ~pi22;
  assign n341 = ~pi14 & n340;
  assign n342 = n293 & n341;
  assign n343 = ~pi5 & ~pi7;
  assign n344 = n323 & n343;
  assign n345 = ~pi13 & n344;
  assign n346 = n295 & n345;
  assign n347 = n342 & n346;
  assign n348 = n339 & ~n347;
  assign n349 = ~pi1 & ~n348;
  assign n350 = pi6 & ~n300;
  assign n351 = ~pi5 & ~pi12;
  assign n352 = pi7 & ~n351;
  assign n353 = ~n323 & ~n343;
  assign n354 = ~pi13 & ~n344;
  assign n355 = ~n350 & ~n352;
  assign n356 = ~n353 & n355;
  assign n357 = n354 & n356;
  assign n358 = pi13 & n344;
  assign n359 = ~pi9 & ~n358;
  assign n360 = ~n357 & n359;
  assign n361 = pi9 & ~n345;
  assign n362 = pi54 & n342;
  assign n363 = n296 & ~n361;
  assign n364 = n362 & n363;
  assign n365 = ~n360 & n364;
  assign n366 = ~n349 & ~n365;
  assign po16 = ~n337 | n366;
  assign n368 = ~pi47 & ~pi48;
  assign n369 = ~pi42 & ~pi44;
  assign n370 = ~pi40 & n369;
  assign n371 = ~pi38 & ~pi50;
  assign n372 = ~pi41 & ~pi46;
  assign n373 = n371 & n372;
  assign n374 = n370 & n373;
  assign n375 = ~pi43 & n374;
  assign n376 = n368 & n375;
  assign n377 = pi82 & ~n376;
  assign n378 = pi122 & pi127;
  assign n379 = ~pi24 & ~pi49;
  assign n380 = ~pi15 & ~pi20;
  assign n381 = ~pi2 & n380;
  assign n382 = n379 & n381;
  assign n383 = pi82 & ~n382;
  assign n384 = n378 & ~n383;
  assign n385 = ~n377 & ~n384;
  assign n386 = ~pi45 & n382;
  assign n387 = n368 & n386;
  assign n388 = pi82 & ~n387;
  assign n389 = n385 & ~n388;
  assign n390 = ~pi65 & n389;
  assign n391 = ~pi82 & n378;
  assign n392 = pi82 & ~n375;
  assign n393 = ~n391 & ~n392;
  assign n394 = ~pi15 & n379;
  assign n395 = ~pi45 & n368;
  assign n396 = n394 & n395;
  assign n397 = ~pi20 & n396;
  assign n398 = pi82 & ~n397;
  assign n399 = n393 & ~n398;
  assign n400 = pi2 & ~n399;
  assign n401 = ~n390 & ~n400;
  assign po17 = ~pi129 & ~n401;
  assign n403 = pi0 & ~pi113;
  assign n404 = ~pi123 & n403;
  assign n405 = ~pi17 & ~pi18;
  assign n406 = n294 & n405;
  assign n407 = ~pi9 & n340;
  assign n408 = n406 & n407;
  assign n409 = n347 & n408;
  assign n410 = ~pi61 & ~pi118;
  assign n411 = ~n409 & n410;
  assign n412 = ~n404 & ~n411;
  assign po18 = ~pi129 & ~n412;
  assign n414 = pi4 & ~pi54;
  assign n415 = ~pi16 & pi54;
  assign n416 = n292 & n415;
  assign n417 = pi10 & n303;
  assign n418 = n416 & n417;
  assign n419 = n298 & n418;
  assign n420 = ~n414 & ~n419;
  assign po19 = n337 & ~n420;
  assign n422 = pi5 & ~pi54;
  assign n423 = ~pi59 & n296;
  assign n424 = ~pi9 & ~pi14;
  assign n425 = n340 & n424;
  assign n426 = ~pi13 & n425;
  assign n427 = n423 & n426;
  assign n428 = n344 & n415;
  assign n429 = ~pi25 & pi28;
  assign n430 = ~pi29 & n429;
  assign n431 = n292 & n430;
  assign n432 = n428 & n431;
  assign n433 = n427 & n432;
  assign n434 = ~n422 & ~n433;
  assign po20 = n337 & ~n434;
  assign n436 = pi6 & ~pi54;
  assign n437 = ~pi28 & ~pi29;
  assign n438 = pi25 & n437;
  assign n439 = n292 & n438;
  assign n440 = n428 & n439;
  assign n441 = n427 & n440;
  assign n442 = ~n436 & ~n441;
  assign po21 = n337 & ~n442;
  assign n444 = pi7 & ~pi54;
  assign n445 = ~pi11 & n344;
  assign n446 = pi8 & ~pi17;
  assign n447 = ~pi21 & n446;
  assign n448 = n416 & n447;
  assign n449 = n426 & n445;
  assign n450 = n448 & n449;
  assign n451 = ~n444 & ~n450;
  assign po22 = n337 & ~n451;
  assign n453 = pi8 & ~pi54;
  assign n454 = n344 & n426;
  assign n455 = n291 & n415;
  assign n456 = ~pi4 & ~pi8;
  assign n457 = ~pi11 & ~pi16;
  assign n458 = n456 & n457;
  assign n459 = n405 & n458;
  assign n460 = pi21 & n455;
  assign n461 = n459 & n460;
  assign n462 = n454 & n461;
  assign n463 = ~n453 & ~n462;
  assign po23 = n337 & ~n463;
  assign n465 = pi9 & ~pi54;
  assign n466 = pi11 & n291;
  assign n467 = n406 & n466;
  assign n468 = n426 & n467;
  assign n469 = n428 & n468;
  assign n470 = ~n465 & ~n469;
  assign po24 = n337 & ~n470;
  assign n472 = pi10 & ~pi54;
  assign n473 = ~pi13 & pi14;
  assign n474 = n455 & n473;
  assign n475 = n408 & n474;
  assign n476 = n445 & n475;
  assign n477 = ~n472 & ~n476;
  assign po25 = n337 & ~n477;
  assign n479 = pi11 & ~pi54;
  assign n480 = n406 & n455;
  assign n481 = n345 & n480;
  assign n482 = ~pi10 & ~pi11;
  assign n483 = pi22 & n482;
  assign n484 = n424 & n483;
  assign n485 = n481 & n484;
  assign n486 = ~n479 & ~n485;
  assign po26 = n337 & ~n486;
  assign n488 = pi12 & ~pi54;
  assign n489 = n296 & n454;
  assign n490 = pi18 & n455;
  assign n491 = n489 & n490;
  assign n492 = ~n488 & ~n491;
  assign po27 = n337 & ~n492;
  assign n494 = pi13 & ~pi54;
  assign n495 = ~pi25 & ~pi28;
  assign n496 = pi29 & n495;
  assign n497 = n425 & n496;
  assign n498 = n423 & n497;
  assign n499 = n481 & n498;
  assign n500 = ~n494 & ~n499;
  assign po28 = n337 & ~n500;
  assign n502 = pi14 & ~pi54;
  assign n503 = n298 & n358;
  assign n504 = n362 & n503;
  assign n505 = ~n502 & ~n504;
  assign po29 = n337 & ~n505;
  assign n507 = pi15 & n391;
  assign n508 = n370 & n371;
  assign n509 = ~pi46 & n508;
  assign n510 = ~pi41 & ~pi43;
  assign n511 = ~pi45 & ~pi47;
  assign n512 = ~pi48 & n511;
  assign n513 = n510 & n512;
  assign n514 = n509 & n513;
  assign n515 = ~pi24 & n514;
  assign n516 = ~pi49 & n515;
  assign n517 = pi15 & ~n516;
  assign n518 = ~n382 & n396;
  assign n519 = n375 & n518;
  assign n520 = ~n517 & ~n519;
  assign n521 = pi82 & ~n520;
  assign n522 = n394 & n514;
  assign n523 = pi82 & ~n522;
  assign n524 = ~pi70 & ~n378;
  assign n525 = ~n523 & n524;
  assign n526 = ~n507 & ~n525;
  assign n527 = ~n521 & n526;
  assign po30 = ~pi129 & ~n527;
  assign n529 = pi16 & ~pi54;
  assign n530 = ~pi11 & n425;
  assign n531 = n480 & n530;
  assign n532 = pi6 & n531;
  assign n533 = n357 & n532;
  assign n534 = ~n529 & ~n533;
  assign po31 = n337 & ~n534;
  assign n536 = pi17 & ~pi54;
  assign n537 = ~pi25 & pi59;
  assign n538 = n339 & n537;
  assign n539 = n437 & n538;
  assign n540 = n295 & n344;
  assign n541 = n539 & n540;
  assign n542 = n293 & n426;
  assign n543 = n541 & n542;
  assign n544 = ~n536 & ~n543;
  assign po32 = n337 & ~n544;
  assign n546 = pi18 & ~pi54;
  assign n547 = pi16 & pi54;
  assign n548 = n292 & n547;
  assign n549 = n489 & n548;
  assign n550 = ~n546 & ~n549;
  assign po33 = n337 & ~n550;
  assign n552 = pi19 & ~pi54;
  assign n553 = pi17 & n295;
  assign n554 = n416 & n553;
  assign n555 = n454 & n554;
  assign n556 = ~n552 & ~n555;
  assign po34 = n337 & ~n556;
  assign n558 = pi20 & n391;
  assign n559 = pi20 & ~n522;
  assign n560 = n380 & n516;
  assign n561 = pi2 & n560;
  assign n562 = ~n559 & ~n561;
  assign n563 = pi82 & ~n562;
  assign n564 = pi82 & ~n560;
  assign n565 = ~pi71 & ~n378;
  assign n566 = ~n564 & n565;
  assign n567 = ~n558 & ~n566;
  assign n568 = ~n563 & n567;
  assign po35 = ~pi129 & ~n568;
  assign n570 = pi21 & ~pi54;
  assign n571 = pi19 & ~pi21;
  assign n572 = pi54 & n571;
  assign n573 = n459 & n572;
  assign n574 = n454 & n573;
  assign n575 = ~n570 & ~n574;
  assign po36 = n337 & ~n575;
  assign n577 = pi22 & ~pi54;
  assign n578 = pi5 & n531;
  assign n579 = n357 & n578;
  assign n580 = ~n577 & ~n579;
  assign po37 = n337 & ~n580;
  assign n582 = ~pi23 & pi55;
  assign n583 = pi61 & ~pi129;
  assign po38 = ~n582 & n583;
  assign n585 = ~pi49 & n381;
  assign n586 = pi82 & ~n585;
  assign n587 = n378 & ~n586;
  assign n588 = pi82 & ~n514;
  assign n589 = ~n587 & ~n588;
  assign n590 = ~pi24 & ~n589;
  assign n591 = pi24 & pi82;
  assign n592 = n514 & n591;
  assign n593 = ~pi45 & n585;
  assign n594 = n376 & n593;
  assign n595 = pi82 & ~n594;
  assign n596 = pi63 & ~n378;
  assign n597 = ~n595 & n596;
  assign n598 = ~pi129 & ~n592;
  assign n599 = ~n590 & n598;
  assign po39 = ~n597 & n599;
  assign n601 = pi25 & ~pi116;
  assign n602 = ~pi39 & ~pi52;
  assign n603 = ~pi51 & n602;
  assign n604 = pi116 & n603;
  assign n605 = ~n601 & ~n604;
  assign n606 = ~pi26 & ~n605;
  assign n607 = pi27 & ~n606;
  assign n608 = ~pi26 & ~pi27;
  assign n609 = pi85 & ~n608;
  assign n610 = pi116 & ~n603;
  assign n611 = pi26 & ~n601;
  assign n612 = ~n610 & n611;
  assign n613 = pi85 & pi116;
  assign n614 = ~pi85 & ~pi110;
  assign n615 = ~pi96 & n614;
  assign n616 = ~n613 & ~n615;
  assign n617 = pi100 & ~n616;
  assign n618 = pi85 & ~n601;
  assign n619 = ~pi27 & ~pi85;
  assign n620 = ~pi95 & ~pi100;
  assign n621 = ~pi97 & n620;
  assign n622 = ~pi110 & ~n621;
  assign n623 = pi25 & ~n622;
  assign n624 = ~pi26 & n619;
  assign n625 = ~n623 & n624;
  assign n626 = ~n618 & ~n625;
  assign n627 = ~n617 & ~n626;
  assign n628 = ~pi53 & ~pi58;
  assign n629 = ~n609 & n628;
  assign n630 = ~n612 & n629;
  assign n631 = ~n607 & n630;
  assign n632 = ~n627 & n631;
  assign n633 = ~pi53 & pi58;
  assign n634 = pi53 & ~pi58;
  assign n635 = ~n633 & ~n634;
  assign n636 = n601 & n624;
  assign n637 = ~n635 & n636;
  assign n638 = ~n632 & ~n637;
  assign po40 = n337 & ~n638;
  assign n640 = ~pi27 & n628;
  assign n641 = ~pi85 & ~n604;
  assign n642 = pi26 & n641;
  assign n643 = pi26 & pi116;
  assign n644 = n617 & ~n643;
  assign n645 = ~n642 & ~n644;
  assign n646 = n337 & n640;
  assign po41 = ~n645 & n646;
  assign n648 = ~pi26 & n337;
  assign n649 = pi27 & n641;
  assign n650 = pi95 & ~pi96;
  assign n651 = n614 & n650;
  assign n652 = ~n613 & ~n651;
  assign n653 = ~pi27 & ~pi100;
  assign n654 = ~n652 & n653;
  assign n655 = ~n649 & ~n654;
  assign n656 = n628 & n648;
  assign po42 = ~n655 & n656;
  assign n658 = ~pi27 & pi28;
  assign n659 = ~pi116 & n658;
  assign n660 = ~pi26 & pi53;
  assign n661 = ~pi85 & n660;
  assign n662 = n659 & n661;
  assign n663 = pi28 & ~pi116;
  assign n664 = ~pi100 & pi116;
  assign n665 = ~n663 & ~n664;
  assign n666 = n608 & ~n665;
  assign n667 = pi85 & ~n666;
  assign n668 = ~n604 & ~n663;
  assign n669 = ~pi27 & ~n668;
  assign n670 = pi26 & ~n669;
  assign n671 = ~pi100 & ~pi110;
  assign n672 = n650 & n671;
  assign n673 = pi28 & ~n622;
  assign n674 = n608 & ~n672;
  assign n675 = ~n673 & n674;
  assign n676 = pi27 & ~n663;
  assign n677 = ~n610 & n676;
  assign n678 = ~n675 & ~n677;
  assign n679 = ~n670 & n678;
  assign n680 = ~pi85 & ~n679;
  assign n681 = ~pi53 & ~n667;
  assign n682 = ~n680 & n681;
  assign n683 = ~n662 & ~n682;
  assign n684 = ~pi58 & ~n683;
  assign n685 = ~pi26 & ~pi53;
  assign n686 = ~pi85 & n685;
  assign n687 = pi58 & n659;
  assign n688 = n686 & n687;
  assign n689 = ~n684 & ~n688;
  assign po43 = n337 & ~n689;
  assign n691 = ~pi116 & ~n635;
  assign n692 = ~n622 & n628;
  assign n693 = ~n691 & ~n692;
  assign n694 = pi29 & ~n693;
  assign n695 = pi58 & pi116;
  assign n696 = ~pi58 & ~pi96;
  assign n697 = ~pi110 & n696;
  assign n698 = n620 & n697;
  assign n699 = ~n695 & ~n698;
  assign n700 = ~pi53 & pi97;
  assign n701 = ~n699 & n700;
  assign n702 = ~n694 & ~n701;
  assign n703 = ~pi27 & ~n702;
  assign n704 = pi29 & ~pi116;
  assign n705 = pi27 & n628;
  assign n706 = n704 & n705;
  assign n707 = ~n703 & ~n706;
  assign n708 = ~pi85 & ~n707;
  assign n709 = pi85 & n704;
  assign n710 = n640 & n709;
  assign n711 = ~n708 & ~n710;
  assign n712 = ~pi26 & ~n711;
  assign n713 = pi26 & ~pi27;
  assign n714 = ~pi85 & n628;
  assign n715 = n713 & n714;
  assign n716 = n704 & n715;
  assign n717 = ~n712 & ~n716;
  assign po44 = n337 & ~n717;
  assign n719 = ~pi88 & pi106;
  assign n720 = ~pi30 & ~pi109;
  assign n721 = ~pi60 & pi109;
  assign n722 = ~n720 & ~n721;
  assign n723 = ~pi106 & ~n722;
  assign n724 = ~pi129 & ~n719;
  assign po45 = ~n723 & n724;
  assign n726 = ~pi89 & pi106;
  assign n727 = ~pi31 & ~pi109;
  assign n728 = ~pi30 & pi109;
  assign n729 = ~n727 & ~n728;
  assign n730 = ~pi106 & ~n729;
  assign n731 = ~pi129 & ~n726;
  assign po46 = ~n730 & n731;
  assign n733 = ~pi99 & pi106;
  assign n734 = ~pi32 & ~pi109;
  assign n735 = ~pi31 & pi109;
  assign n736 = ~n734 & ~n735;
  assign n737 = ~pi106 & ~n736;
  assign n738 = ~pi129 & ~n733;
  assign po47 = ~n737 & n738;
  assign n740 = ~pi90 & pi106;
  assign n741 = ~pi33 & ~pi109;
  assign n742 = ~pi32 & pi109;
  assign n743 = ~n741 & ~n742;
  assign n744 = ~pi106 & ~n743;
  assign n745 = ~pi129 & ~n740;
  assign po48 = ~n744 & n745;
  assign n747 = ~pi91 & pi106;
  assign n748 = ~pi34 & ~pi109;
  assign n749 = ~pi33 & pi109;
  assign n750 = ~n748 & ~n749;
  assign n751 = ~pi106 & ~n750;
  assign n752 = ~pi129 & ~n747;
  assign po49 = ~n751 & n752;
  assign n754 = ~pi92 & pi106;
  assign n755 = ~pi35 & ~pi109;
  assign n756 = ~pi34 & pi109;
  assign n757 = ~n755 & ~n756;
  assign n758 = ~pi106 & ~n757;
  assign n759 = ~pi129 & ~n754;
  assign po50 = ~n758 & n759;
  assign n761 = ~pi98 & pi106;
  assign n762 = ~pi36 & ~pi109;
  assign n763 = ~pi35 & pi109;
  assign n764 = ~n762 & ~n763;
  assign n765 = ~pi106 & ~n764;
  assign n766 = ~pi129 & ~n761;
  assign po51 = ~n765 & n766;
  assign n768 = ~pi93 & pi106;
  assign n769 = ~pi37 & ~pi109;
  assign n770 = ~pi36 & pi109;
  assign n771 = ~n769 & ~n770;
  assign n772 = ~pi106 & ~n771;
  assign n773 = ~pi129 & ~n768;
  assign po52 = ~n772 & n773;
  assign n775 = pi38 & pi82;
  assign n776 = n370 & n775;
  assign n777 = n382 & n513;
  assign n778 = ~pi46 & n777;
  assign n779 = ~pi50 & n370;
  assign n780 = n778 & n779;
  assign n781 = pi82 & ~n780;
  assign n782 = pi74 & ~n378;
  assign n783 = ~n781 & n782;
  assign n784 = ~pi38 & n370;
  assign n785 = pi82 & ~n784;
  assign n786 = pi82 & ~n778;
  assign n787 = n378 & ~n786;
  assign n788 = ~n785 & ~n787;
  assign n789 = pi82 & ~n508;
  assign n790 = n784 & n789;
  assign n791 = ~pi38 & ~n790;
  assign n792 = ~n788 & n791;
  assign n793 = ~pi129 & ~n776;
  assign n794 = ~n783 & n793;
  assign po53 = ~n792 & n794;
  assign n796 = ~pi51 & ~pi52;
  assign n797 = pi109 & n796;
  assign n798 = pi39 & ~n797;
  assign n799 = ~pi51 & pi109;
  assign n800 = n602 & n799;
  assign n801 = ~pi106 & ~n800;
  assign n802 = ~n798 & n801;
  assign po54 = ~pi129 & ~n802;
  assign n804 = pi82 & ~n369;
  assign n805 = ~pi43 & n387;
  assign n806 = n373 & n805;
  assign n807 = ~pi40 & n806;
  assign n808 = pi82 & ~n807;
  assign n809 = n378 & ~n808;
  assign n810 = ~n804 & ~n809;
  assign n811 = ~pi40 & ~n810;
  assign n812 = pi82 & n369;
  assign n813 = ~n370 & n812;
  assign n814 = pi82 & ~n806;
  assign n815 = pi73 & ~n378;
  assign n816 = ~n804 & n815;
  assign n817 = ~n814 & n816;
  assign n818 = ~pi129 & ~n813;
  assign n819 = ~n817 & n818;
  assign po55 = ~n811 & n819;
  assign n821 = pi82 & ~n374;
  assign n822 = n509 & n821;
  assign n823 = n509 & n805;
  assign n824 = pi82 & ~n823;
  assign n825 = pi76 & ~n378;
  assign n826 = ~n824 & n825;
  assign n827 = pi82 & ~n509;
  assign n828 = pi82 & ~n777;
  assign n829 = n378 & ~n828;
  assign n830 = ~n827 & ~n829;
  assign n831 = ~pi41 & ~n830;
  assign n832 = ~pi129 & ~n822;
  assign n833 = ~n831 & n832;
  assign po56 = ~n826 & n833;
  assign n835 = ~pi44 & n804;
  assign n836 = pi44 & pi82;
  assign n837 = ~n809 & ~n836;
  assign n838 = ~pi42 & ~n837;
  assign n839 = pi72 & ~n808;
  assign n840 = n837 & n839;
  assign n841 = ~pi129 & ~n835;
  assign n842 = ~n838 & n841;
  assign po57 = ~n840 & n842;
  assign n844 = n374 & n392;
  assign n845 = n378 & ~n388;
  assign n846 = ~n821 & ~n845;
  assign n847 = pi77 & ~n388;
  assign n848 = n846 & n847;
  assign n849 = ~pi43 & ~n846;
  assign n850 = ~pi129 & ~n844;
  assign n851 = ~n848 & n850;
  assign po58 = ~n849 & n851;
  assign n853 = ~pi42 & n807;
  assign n854 = pi82 & ~n853;
  assign n855 = ~pi67 & ~n378;
  assign n856 = pi44 & n378;
  assign n857 = ~n855 & ~n856;
  assign n858 = ~n854 & n857;
  assign n859 = ~pi129 & ~n836;
  assign po59 = ~n858 & n859;
  assign n861 = pi68 & ~n383;
  assign n862 = n385 & n861;
  assign n863 = ~pi45 & ~n385;
  assign n864 = pi45 & pi82;
  assign n865 = n376 & n864;
  assign n866 = ~pi129 & ~n865;
  assign n867 = ~n862 & n866;
  assign po60 = ~n863 & n867;
  assign n869 = n508 & n827;
  assign n870 = ~n789 & ~n829;
  assign n871 = pi75 & ~n828;
  assign n872 = n870 & n871;
  assign n873 = ~pi46 & ~n870;
  assign n874 = ~pi129 & ~n869;
  assign n875 = ~n872 & n874;
  assign po61 = ~n873 & n875;
  assign n877 = ~pi47 & n375;
  assign n878 = n814 & n877;
  assign n879 = pi47 & ~n393;
  assign n880 = pi82 & ~n877;
  assign n881 = ~n378 & ~n880;
  assign n882 = ~pi64 & n881;
  assign n883 = ~n879 & ~n882;
  assign n884 = ~n878 & n883;
  assign po62 = ~pi129 & ~n884;
  assign n886 = n377 & n877;
  assign n887 = ~pi48 & ~n865;
  assign n888 = ~n385 & n887;
  assign n889 = pi82 & ~n386;
  assign n890 = pi62 & ~n889;
  assign n891 = n881 & n890;
  assign n892 = ~pi129 & ~n886;
  assign n893 = ~n888 & n892;
  assign po63 = ~n891 & n893;
  assign n895 = pi49 & n391;
  assign n896 = pi49 & ~n515;
  assign n897 = ~n516 & ~n896;
  assign n898 = n586 & ~n897;
  assign n899 = pi82 & ~n516;
  assign n900 = ~pi69 & ~n378;
  assign n901 = ~n899 & n900;
  assign n902 = ~n895 & ~n898;
  assign n903 = ~n901 & n902;
  assign po64 = ~pi129 & ~n903;
  assign n905 = pi66 & ~n786;
  assign n906 = n788 & n905;
  assign n907 = ~pi50 & ~n788;
  assign n908 = ~pi129 & ~n790;
  assign n909 = ~n906 & n908;
  assign po65 = ~n907 & n909;
  assign n911 = pi51 & ~pi109;
  assign n912 = ~pi106 & ~n799;
  assign n913 = ~n911 & n912;
  assign po66 = ~pi129 & ~n913;
  assign n915 = pi52 & ~n799;
  assign n916 = ~pi106 & ~n797;
  assign n917 = ~n915 & n916;
  assign po67 = ~pi129 & ~n917;
  assign n919 = ~pi116 & n634;
  assign n920 = ~n701 & ~n919;
  assign n921 = n619 & n648;
  assign po68 = ~n920 & n921;
  assign po69 = pi129 | n389;
  assign po129 = pi123 | pi129;
  assign n925 = pi114 & ~pi122;
  assign po70 = ~po129 & n925;
  assign n927 = ~pi26 & pi58;
  assign n928 = ~pi58 & n643;
  assign n929 = ~n927 & ~n928;
  assign n930 = pi94 & ~n929;
  assign n931 = pi58 & ~pi116;
  assign n932 = pi37 & ~pi116;
  assign n933 = ~n927 & ~n932;
  assign n934 = ~n931 & ~n933;
  assign n935 = ~n930 & ~n934;
  assign n936 = ~pi53 & ~n935;
  assign n937 = ~pi26 & pi37;
  assign n938 = ~pi58 & n937;
  assign n939 = ~n936 & ~n938;
  assign n940 = ~pi85 & ~n939;
  assign n941 = n628 & n937;
  assign n942 = ~n940 & ~n941;
  assign n943 = ~pi27 & ~n942;
  assign n944 = n714 & n937;
  assign n945 = ~n943 & ~n944;
  assign po71 = n337 & ~n945;
  assign n947 = ~pi116 & n686;
  assign n948 = ~pi53 & ~pi85;
  assign n949 = ~n685 & ~n948;
  assign n950 = ~n661 & n949;
  assign n951 = ~pi58 & ~n950;
  assign n952 = ~n947 & ~n951;
  assign n953 = pi57 & ~n952;
  assign n954 = pi60 & n695;
  assign n955 = n686 & n954;
  assign n956 = ~n953 & ~n955;
  assign n957 = ~pi27 & ~n956;
  assign n958 = pi57 & ~pi58;
  assign n959 = n686 & n958;
  assign n960 = ~n957 & ~n959;
  assign po72 = n337 & ~n960;
  assign n962 = n608 & n931;
  assign n963 = ~pi26 & pi27;
  assign n964 = ~n713 & ~n963;
  assign n965 = ~pi58 & ~n964;
  assign n966 = n604 & n965;
  assign n967 = ~n962 & ~n966;
  assign n968 = n337 & n948;
  assign po73 = ~n967 & n968;
  assign n970 = pi59 & ~n693;
  assign n971 = pi96 & n628;
  assign n972 = n622 & n971;
  assign n973 = ~n970 & ~n972;
  assign n974 = ~pi85 & ~n973;
  assign n975 = pi59 & ~pi116;
  assign n976 = pi85 & n628;
  assign n977 = n975 & n976;
  assign n978 = ~n974 & ~n977;
  assign n979 = ~pi27 & ~n978;
  assign n980 = pi27 & n975;
  assign n981 = n714 & n980;
  assign n982 = ~n979 & ~n981;
  assign n983 = ~pi26 & ~n982;
  assign n984 = n715 & n975;
  assign n985 = ~n983 & ~n984;
  assign po74 = n337 & ~n985;
  assign n987 = ~pi117 & ~pi122;
  assign n988 = pi60 & ~n987;
  assign n989 = pi123 & n987;
  assign po75 = n988 | n989;
  assign n991 = ~pi114 & ~pi122;
  assign n992 = pi123 & ~pi129;
  assign po76 = n991 & n992;
  assign n994 = pi136 & ~pi137;
  assign n995 = pi131 & pi132;
  assign n996 = pi133 & n995;
  assign n997 = ~pi138 & n996;
  assign n998 = n994 & n997;
  assign n999 = ~pi62 & ~n998;
  assign n1000 = pi140 & n998;
  assign n1001 = ~pi129 & ~n999;
  assign po77 = n1000 | ~n1001;
  assign n1003 = ~pi63 & ~n998;
  assign n1004 = pi142 & n998;
  assign n1005 = ~pi129 & ~n1003;
  assign po78 = n1004 | ~n1005;
  assign n1007 = ~pi64 & ~n998;
  assign n1008 = pi139 & n998;
  assign n1009 = ~pi129 & ~n1007;
  assign po79 = n1008 | ~n1009;
  assign n1011 = ~pi65 & ~n998;
  assign n1012 = pi146 & n998;
  assign n1013 = ~pi129 & ~n1011;
  assign po80 = n1012 | ~n1013;
  assign n1015 = ~pi136 & ~pi137;
  assign n1016 = n997 & n1015;
  assign n1017 = ~pi66 & ~n1016;
  assign n1018 = pi143 & n1016;
  assign n1019 = ~pi129 & ~n1017;
  assign po81 = n1018 | ~n1019;
  assign n1021 = ~pi67 & ~n1016;
  assign n1022 = pi139 & n1016;
  assign n1023 = ~pi129 & ~n1021;
  assign po82 = n1022 | ~n1023;
  assign n1025 = ~pi68 & ~n998;
  assign n1026 = pi141 & n998;
  assign n1027 = ~pi129 & ~n1025;
  assign po83 = n1026 | ~n1027;
  assign n1029 = ~pi69 & ~n998;
  assign n1030 = pi143 & n998;
  assign n1031 = ~pi129 & ~n1029;
  assign po84 = n1030 | ~n1031;
  assign n1033 = ~pi70 & ~n998;
  assign n1034 = pi144 & n998;
  assign n1035 = ~pi129 & ~n1033;
  assign po85 = n1034 | ~n1035;
  assign n1037 = ~pi71 & ~n998;
  assign n1038 = pi145 & n998;
  assign n1039 = ~pi129 & ~n1037;
  assign po86 = n1038 | ~n1039;
  assign n1041 = ~pi72 & ~n1016;
  assign n1042 = pi140 & n1016;
  assign n1043 = ~pi129 & ~n1041;
  assign po87 = n1042 | ~n1043;
  assign n1045 = ~pi73 & ~n1016;
  assign n1046 = pi141 & n1016;
  assign n1047 = ~pi129 & ~n1045;
  assign po88 = n1046 | ~n1047;
  assign n1049 = ~pi74 & ~n1016;
  assign n1050 = pi142 & n1016;
  assign n1051 = ~pi129 & ~n1049;
  assign po89 = n1050 | ~n1051;
  assign n1053 = ~pi75 & ~n1016;
  assign n1054 = pi144 & n1016;
  assign n1055 = ~pi129 & ~n1053;
  assign po90 = n1054 | ~n1055;
  assign n1057 = ~pi76 & ~n1016;
  assign n1058 = pi145 & n1016;
  assign n1059 = ~pi129 & ~n1057;
  assign po91 = n1058 | ~n1059;
  assign n1061 = ~pi77 & ~n1016;
  assign n1062 = pi146 & n1016;
  assign n1063 = ~pi129 & ~n1061;
  assign po92 = n1062 | ~n1063;
  assign n1065 = ~pi136 & pi137;
  assign n1066 = n997 & n1065;
  assign n1067 = ~pi78 & ~n1066;
  assign n1068 = ~pi142 & n1066;
  assign n1069 = ~pi129 & ~n1067;
  assign po93 = ~n1068 & n1069;
  assign n1071 = ~pi79 & ~n1066;
  assign n1072 = ~pi143 & n1066;
  assign n1073 = ~pi129 & ~n1071;
  assign po94 = ~n1072 & n1073;
  assign n1075 = ~pi80 & ~n1066;
  assign n1076 = ~pi144 & n1066;
  assign n1077 = ~pi129 & ~n1075;
  assign po95 = ~n1076 & n1077;
  assign n1079 = ~pi81 & ~n1066;
  assign n1080 = ~pi145 & n1066;
  assign n1081 = ~pi129 & ~n1079;
  assign po96 = ~n1080 & n1081;
  assign n1083 = ~pi82 & ~n1066;
  assign n1084 = ~pi146 & n1066;
  assign n1085 = ~pi129 & ~n1083;
  assign po97 = ~n1084 & n1085;
  assign n1087 = pi136 & ~pi138;
  assign n1088 = pi31 & n1087;
  assign n1089 = ~pi87 & ~pi138;
  assign n1090 = pi115 & pi138;
  assign n1091 = ~pi136 & ~n1089;
  assign n1092 = ~n1090 & n1091;
  assign n1093 = ~n1088 & ~n1092;
  assign n1094 = pi137 & ~n1093;
  assign n1095 = ~pi89 & pi138;
  assign n1096 = pi62 & ~pi138;
  assign n1097 = pi136 & ~n1095;
  assign n1098 = ~n1096 & n1097;
  assign n1099 = ~pi119 & pi138;
  assign n1100 = pi72 & ~pi138;
  assign n1101 = ~pi136 & ~n1099;
  assign n1102 = ~n1100 & n1101;
  assign n1103 = ~n1098 & ~n1102;
  assign n1104 = ~pi137 & ~n1103;
  assign po98 = n1094 | n1104;
  assign n1106 = ~pi84 & ~n1066;
  assign n1107 = ~pi141 & n1066;
  assign n1108 = ~pi129 & ~n1106;
  assign po99 = ~n1107 & n1108;
  assign n1110 = ~pi85 & ~n622;
  assign n1111 = n640 & n648;
  assign n1112 = n616 & n1111;
  assign po100 = ~n1110 & n1112;
  assign n1114 = ~pi86 & ~n1066;
  assign n1115 = ~pi139 & n1066;
  assign n1116 = ~pi129 & ~n1114;
  assign po101 = ~n1115 & n1116;
  assign n1118 = ~pi87 & ~n1066;
  assign n1119 = ~pi140 & n1066;
  assign n1120 = ~pi129 & ~n1118;
  assign po102 = ~n1119 & n1120;
  assign n1122 = pi137 & n1087;
  assign n1123 = n996 & n1122;
  assign n1124 = ~pi88 & ~n1123;
  assign n1125 = ~pi139 & n1123;
  assign n1126 = ~pi129 & ~n1124;
  assign po103 = ~n1125 & n1126;
  assign n1128 = ~pi89 & ~n1123;
  assign n1129 = ~pi140 & n1123;
  assign n1130 = ~pi129 & ~n1128;
  assign po104 = ~n1129 & n1130;
  assign n1132 = ~pi90 & ~n1123;
  assign n1133 = ~pi142 & n1123;
  assign n1134 = ~pi129 & ~n1132;
  assign po105 = ~n1133 & n1134;
  assign n1136 = ~pi91 & ~n1123;
  assign n1137 = ~pi143 & n1123;
  assign n1138 = ~pi129 & ~n1136;
  assign po106 = ~n1137 & n1138;
  assign n1140 = ~pi92 & ~n1123;
  assign n1141 = ~pi144 & n1123;
  assign n1142 = ~pi129 & ~n1140;
  assign po107 = ~n1141 & n1142;
  assign n1144 = ~pi93 & ~n1123;
  assign n1145 = ~pi146 & n1123;
  assign n1146 = ~pi129 & ~n1144;
  assign po108 = ~n1145 & n1146;
  assign n1148 = pi82 & pi138;
  assign n1149 = n1015 & n1148;
  assign n1150 = n996 & n1149;
  assign n1151 = ~pi94 & ~n1150;
  assign n1152 = ~pi142 & n1150;
  assign n1153 = ~pi129 & ~n1151;
  assign po109 = ~n1152 & n1153;
  assign n1155 = ~pi3 & ~pi110;
  assign n1156 = ~n996 & ~n1155;
  assign n1157 = ~n1150 & ~n1156;
  assign n1158 = pi95 & n1157;
  assign n1159 = pi143 & n1150;
  assign n1160 = ~n1158 & ~n1159;
  assign po110 = ~pi129 & ~n1160;
  assign n1162 = pi96 & n1157;
  assign n1163 = pi146 & n1150;
  assign n1164 = ~n1162 & ~n1163;
  assign po111 = ~pi129 & ~n1164;
  assign n1166 = pi97 & n1157;
  assign n1167 = pi145 & n1150;
  assign n1168 = ~n1166 & ~n1167;
  assign po112 = ~pi129 & ~n1168;
  assign n1170 = ~pi98 & ~n1123;
  assign n1171 = ~pi145 & n1123;
  assign n1172 = ~pi129 & ~n1170;
  assign po113 = ~n1171 & n1172;
  assign n1174 = ~pi99 & ~n1123;
  assign n1175 = ~pi141 & n1123;
  assign n1176 = ~pi129 & ~n1174;
  assign po114 = ~n1175 & n1176;
  assign n1178 = pi100 & n1157;
  assign n1179 = pi144 & n1150;
  assign n1180 = ~n1178 & ~n1179;
  assign po115 = ~pi129 & ~n1180;
  assign n1182 = pi37 & n1087;
  assign n1183 = ~pi82 & ~pi138;
  assign n1184 = ~pi96 & pi138;
  assign n1185 = ~pi136 & ~n1183;
  assign n1186 = ~n1184 & n1185;
  assign n1187 = ~n1182 & ~n1186;
  assign n1188 = pi137 & ~n1187;
  assign n1189 = ~pi93 & pi138;
  assign n1190 = pi65 & ~pi138;
  assign n1191 = pi136 & ~n1189;
  assign n1192 = ~n1190 & n1191;
  assign n1193 = ~pi124 & pi138;
  assign n1194 = pi77 & ~pi138;
  assign n1195 = ~pi136 & ~n1193;
  assign n1196 = ~n1194 & n1195;
  assign n1197 = ~n1192 & ~n1196;
  assign n1198 = ~pi137 & ~n1197;
  assign po116 = n1188 | n1198;
  assign n1200 = pi91 & n994;
  assign n1201 = pi95 & n1065;
  assign n1202 = ~n1200 & ~n1201;
  assign n1203 = pi138 & ~n1202;
  assign n1204 = ~pi79 & ~pi136;
  assign n1205 = ~pi34 & pi136;
  assign n1206 = pi137 & ~n1204;
  assign n1207 = ~n1205 & n1206;
  assign n1208 = pi66 & ~pi136;
  assign n1209 = pi69 & pi136;
  assign n1210 = ~pi137 & ~n1208;
  assign n1211 = ~n1209 & n1210;
  assign n1212 = ~n1207 & ~n1211;
  assign n1213 = ~pi138 & ~n1212;
  assign po117 = n1203 | n1213;
  assign n1215 = pi90 & n994;
  assign n1216 = pi94 & n1065;
  assign n1217 = ~n1215 & ~n1216;
  assign n1218 = pi138 & ~n1217;
  assign n1219 = ~pi78 & ~pi136;
  assign n1220 = ~pi33 & pi136;
  assign n1221 = pi137 & ~n1219;
  assign n1222 = ~n1220 & n1221;
  assign n1223 = pi74 & ~pi136;
  assign n1224 = pi63 & pi136;
  assign n1225 = ~pi137 & ~n1223;
  assign n1226 = ~n1224 & n1225;
  assign n1227 = ~n1222 & ~n1226;
  assign n1228 = ~pi138 & ~n1227;
  assign po118 = n1218 | n1228;
  assign n1230 = pi99 & n994;
  assign n1231 = ~pi112 & n1065;
  assign n1232 = ~n1230 & ~n1231;
  assign n1233 = pi138 & ~n1232;
  assign n1234 = ~pi84 & ~pi136;
  assign n1235 = ~pi32 & pi136;
  assign n1236 = pi137 & ~n1234;
  assign n1237 = ~n1235 & n1236;
  assign n1238 = pi73 & ~pi136;
  assign n1239 = pi68 & pi136;
  assign n1240 = ~pi137 & ~n1238;
  assign n1241 = ~n1239 & n1240;
  assign n1242 = ~n1237 & ~n1241;
  assign n1243 = ~pi138 & ~n1242;
  assign po119 = n1233 | n1243;
  assign n1245 = pi35 & n1087;
  assign n1246 = ~pi80 & ~pi138;
  assign n1247 = ~pi100 & pi138;
  assign n1248 = ~pi136 & ~n1246;
  assign n1249 = ~n1247 & n1248;
  assign n1250 = ~n1245 & ~n1249;
  assign n1251 = pi137 & ~n1250;
  assign n1252 = ~pi92 & pi138;
  assign n1253 = pi70 & ~pi138;
  assign n1254 = pi136 & ~n1252;
  assign n1255 = ~n1253 & n1254;
  assign n1256 = ~pi125 & pi138;
  assign n1257 = pi75 & ~pi138;
  assign n1258 = ~pi136 & ~n1256;
  assign n1259 = ~n1257 & n1258;
  assign n1260 = ~n1255 & ~n1259;
  assign n1261 = ~pi137 & ~n1260;
  assign po120 = n1251 | n1261;
  assign n1263 = n608 & n714;
  assign n1264 = n622 & n1263;
  assign n1265 = ~n613 & ~n1264;
  assign po121 = n337 & ~n1265;
  assign n1267 = pi36 & n1087;
  assign n1268 = ~pi81 & ~pi138;
  assign n1269 = ~pi97 & pi138;
  assign n1270 = ~pi136 & ~n1268;
  assign n1271 = ~n1269 & n1270;
  assign n1272 = ~n1267 & ~n1271;
  assign n1273 = pi137 & ~n1272;
  assign n1274 = ~pi98 & pi138;
  assign n1275 = pi71 & ~pi138;
  assign n1276 = pi136 & ~n1274;
  assign n1277 = ~n1275 & n1276;
  assign n1278 = ~pi23 & pi138;
  assign n1279 = pi76 & ~pi138;
  assign n1280 = ~pi136 & ~n1278;
  assign n1281 = ~n1279 & n1280;
  assign n1282 = ~n1277 & ~n1281;
  assign n1283 = ~pi137 & ~n1282;
  assign po122 = n1273 | n1283;
  assign n1285 = pi30 & n1087;
  assign n1286 = ~pi86 & ~pi138;
  assign n1287 = ~pi111 & pi138;
  assign n1288 = ~pi136 & ~n1286;
  assign n1289 = ~n1287 & n1288;
  assign n1290 = ~n1285 & ~n1289;
  assign n1291 = pi137 & ~n1290;
  assign n1292 = ~pi88 & pi138;
  assign n1293 = pi64 & ~pi138;
  assign n1294 = pi136 & ~n1292;
  assign n1295 = ~n1293 & n1294;
  assign n1296 = ~pi120 & pi138;
  assign n1297 = pi67 & ~pi138;
  assign n1298 = ~pi136 & ~n1296;
  assign n1299 = ~n1297 & n1298;
  assign n1300 = ~n1295 & ~n1299;
  assign n1301 = ~pi137 & ~n1300;
  assign po123 = n1291 | n1301;
  assign n1303 = pi116 & n337;
  assign n1304 = pi27 & n603;
  assign n1305 = ~n964 & n1303;
  assign po124 = ~n1304 & n1305;
  assign n1307 = ~pi97 & n633;
  assign n1308 = ~n634 & ~n1307;
  assign po125 = n1303 & ~n1308;
  assign n1310 = ~pi129 & n996;
  assign n1311 = ~pi111 & ~n1149;
  assign n1312 = ~pi139 & n1149;
  assign n1313 = n1310 & ~n1311;
  assign po126 = ~n1312 & n1313;
  assign n1315 = ~pi141 & n1149;
  assign n1316 = pi112 & ~n1149;
  assign n1317 = n1310 & ~n1315;
  assign po127 = ~n1316 & n1317;
  assign n1319 = ~pi54 & pi113;
  assign n1320 = ~pi11 & ~pi22;
  assign n1321 = pi54 & n1320;
  assign n1322 = n337 & ~n1319;
  assign po128 = ~n1321 & n1322;
  assign n1324 = ~pi140 & n1149;
  assign n1325 = pi115 & ~n1149;
  assign n1326 = n1310 & ~n1324;
  assign po130 = ~n1325 & n1326;
  assign n1328 = ~pi4 & ~pi9;
  assign n1329 = n300 & n1328;
  assign n1330 = pi54 & n337;
  assign po131 = ~n1329 & n1330;
  assign po132 = ~pi122 | pi129;
  assign n1333 = ~pi54 & pi118;
  assign n1334 = pi54 & ~pi59;
  assign n1335 = n496 & n1334;
  assign n1336 = ~n1333 & ~n1335;
  assign po133 = ~pi129 & ~n1336;
  assign po134 = ~pi129 & ~n620;
  assign n1339 = ~pi120 & n1155;
  assign n1340 = ~pi111 & ~pi129;
  assign po135 = ~n1339 & n1340;
  assign n1342 = pi81 & pi120;
  assign po136 = ~pi129 & n1342;
  assign po137 = pi129 | pi134;
  assign po138 = pi129 | pi135;
  assign po139 = pi57 & ~pi129;
  assign n1347 = ~pi96 & pi125;
  assign n1348 = ~pi3 & ~n1347;
  assign po140 = ~pi129 & ~n1348;
  assign n1350 = ~pi126 & pi132;
  assign po141 = pi133 & n1350;
  assign po12 = 1'b1;
  assign po0 = pi108;
  assign po1 = pi83;
  assign po2 = pi104;
  assign po3 = pi103;
  assign po4 = pi102;
  assign po5 = pi105;
  assign po6 = pi107;
  assign po7 = pi101;
  assign po8 = pi126;
  assign po9 = pi121;
  assign po10 = pi1;
  assign po11 = pi0;
  assign po13 = pi130;
  assign po14 = pi128;
endmodule
